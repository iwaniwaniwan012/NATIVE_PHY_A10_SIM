// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 01:23:56 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oUE9ejpSRb1hPHZXXFsXq/gs/RiGVaekChk5S2CbvmLeKY5sMP/3lvBSoGxFRpuc
jLWm3YF8oqK7SkKrylUYwA8R+hU1lFtNDtl2N/sAlDUs28fmyDULIdBiUAAnw+MM
VZ/sIolw0yMs+CV8v5mQwEHXLg5xXwf4CmWlvkspkOI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2992)
VzPFoWlipyCdJqDPFa/nX9RKodltEVb0ntmofyxkRnoIaIff+n14ncq+5vGxVM+0
MeEq3FTGYPnOo+MWo+7MUtKFhZMB1whPW5AI5mGFBRZUI1S2boB4OOuYty0yLXzE
fHR0s5Wq3UJLM7hlLNSTv0Urkh4BgcLvbvaKX9FSnnhhuKIPneDmvMYhFGIxPvBm
RXtad38CWGwvQnpD9svpIGKfzyygpWlTJv+QxA2AgI3S/IJmV4ivUccEonWMN8vM
kb4Xdv++EGaayQXsGMHtogDYgbK7gr50681Y5Az0C8pXxPvDGh0f9qeA8uHxYu5G
ajV1dDdi7/FnKc41n2hTxZ8mGFSrEatA6eANhXPqyB9TX+XHIbUukSHTxfeImJCa
rrAE3sI/gevyrvv82jChBCjL+red6mtl3RjY+IbhcRXGR8g3yVmwGTEpNN8FkFLR
9cDvHe2Rx6aqyB+iDq+WOVQ+iEbNBZ1qlexR3tERWPybm2osA5Bl8YTSPt/acnrR
kfj+kcDyz1fSk1tFHAwe5DQCznc62VSVGG37RuunEZaPFI20SrFxJ6V9FtjffN6/
IcQyorgDCM18FVMbDfpdXhqYT/QDS3eP3Qp6irS7sWmZDoJNNYTWaSODDqf+y9hh
pAo7ws8RRC3S8Lu+qsZw4jwISLfli9sWhEcSOkgk2j6kbyAe1N5d6lzflc5Gk2pL
tgG8OGVCiUVxzOxjSE/vNnTpiuwRopnGFAIEK/i28tAllTwXWWaOX+j88wAGE+gr
qXR8uXKe+PbpPFBjxDvCp5hwUvQMSf0eoZ/wXAqJ+wBkKgS03tdg402oO7rfSUTN
0hrvLyhFUrkX3+k+nQnDOJRzZFSLGvR5Ox5LbDvcU9ps2iuMfG9g/Am/SiRtGIE+
eAF05XLr4X2t04n9Y5cArMRLlVSXdOud/BefmWS8miKEssT4ERBU4aXMeZq1Mk+u
obp5Kyb3tmqnp8bF4GgoBxAPjPIZgoKONwqwsJkD5sXKoI8CDSqMUXS59I2UaWUM
+/SJcq6UoU2RSQoqMM6xBm+uPCANRViFgEobXqGOCcHsaxGj+bRsavaciZABii6Z
vVcIwJ9dWC7KSNtqzB+XQQCAeu2KO5w2t/V0hi99lIfLhdZDLgOyQ8ERstn0aCr0
KikjsHn/spiJdrEjfAuKKQVJ/I71AUxWQ8cMhWjT+IahLPOZMGxSITm7gCwbqEC1
8Rn/XOS1K3g5dY7je881kF6nmLnY+Hy7R48o5mAaN2ovp5pkS+isdTaGFw+hawEE
NjYUPzJQumgUyhkFPJBBjSG1YYzfbDyRaN1Yutr5/xi77BIFk8Wv4Sy292PKWrmu
e1BD++e6tDIMMPiC6CHJbBXPwIQesBKvR2tl9fIIcok1cKGLPLgFoeO81EU1z6d5
uD1JnrE3zTjvnWmcxld0vWmkzzw09RZ+EJfRmzxfc0XQvoVbxdQL+pDJiYC5Vp0a
42E9egGr+VNf3jy3dLsOgiDkeulp6xptl1jTssGEPuhYP+8ft+7wGTMsum9pk1UU
nnhmfekp/EYTWLzyx3nF6Y2jkXE4boPwRuZ7/2DeNQEvq7cqj78fCcDWGiGyKyEy
08Q/deGlBLrSLRnoKV0S3v9tZWUV5h1UhG4uSkMRbxJB0yvv/Gx/8aRxRPYMXvil
Fck9R7CbHzBWyPt1ZcEpPsGfejC/3NxrFGWZd0X8JoN00SoB6lEX+cAQ7JlyfWxM
JKNv977zoMRhKAMRdGHbLdMLh8F451ziOEeARvIm4Dyq8waMReIWEoKTexHjE6T7
iqrHD+pmLlgJgkzdhq9HHmVOJoR/0MD1MI/IOL+UIwmJ5sWfwdLgAbTfX83jBFCC
D+zTdOBlvnyc38EUezDWUmkhbc+v/+NE4uxfyNuXAhECc9nDJcgqUmwyGJhJqd9l
t9Nt7xRmJdv4NN2H5ZXnelMnT3OxMvxu0UT8S4EXG6uG632zrX3xZd6tUQfYfWQY
ZGmUHG5k25azHIyWep3AhLX8TnR2+zK1FJO9bIEHp5Wudb0f/b38y+wwQHSkq5iz
NaMl5b68RZo/ZrCEfqQ5LCmYbK1yYXdwsfFHPuslqHr2hwvsZlpDJOuiYM7DMROs
yp4KRJPfuJ8oLm+XnaxlMFnZC9CKRuwgFxJwgkuPxUvj0fwU9U+TXbezaDBkDfiN
s3LLdaqcRdmmORzHj//6nOfH4/tL5EQcb6iemIRaGQTaF4FLtOtb08y4yfS5vif7
jJzxq8PM8n9oylp4DfZd9dW7kKSR7D44WbMhrUYz3K0m6BxSqNV7WkSAOUgJxAjC
HiMtq99SaX50s2zmqWHiad8EubUaJ7az5giP2+616jUNyTgZcQbT0rVs8xGAlYcb
iW2LSg73GuE9nrH+ElfeAN40ur75SbGEQBxO79ZBccim67Mn2mY1HL1V5xPq26dG
EkhsSQJyJbzY6HzYZbffJualBaxhJU7d3ul9i/LLHmuKJdbT9D2rLY0y0PI6HfGZ
C2zQgOMHymBA+3piktzJh7MQYL0SnqK92MIpH2ZxpQMQqMyXy/Nrx/eYhWK/ggqh
cM3tpzNHv7Lszi+jE/aK6exFQAyIHpR6R98GsndO+n+swxnkTcNds6P7lA9n+n+V
15J4NCHsGSkeRR5R8lH/y6nQrRNUTBYfHzfHL1IK+2UKzl/r0WMF1yRaOmZRQEO/
tE9eMWugO5jZ+k4dk5ETULuxeGSMPcNom9EH41LI4Nnx1RwgP4hTfk1iyz1j+q2A
VvXiFnXdDma5IV5ye+yMUaHN/BiWktkxeQS9T+74qDMk3punwX1zhK9r09Rin0XC
kp0T0piVfJB5xd/mDgOF24WHQvEEbHt1IOEnNe8q1UwgZpdkGQYuX97oYYLZvLfF
5VagILWhLQlqs5xnMNi7q49ObuKmPZJfb4wTV+D5eInsvI6JQQXqh4k+mh7/+c5u
qqSMwl1fA1umcYuE51Eco76RiXCAAUq6ANR90kfPd575ClzpFk04llr6lFAzvgfs
msEDEpH5thRwRK991omm2TzvBIQBnVJRtTdeOtucrDJsxxks315gfbLMpM8LZ26E
f2NsDugnjeB7NwSX1iMiDeWVW4yfGbUmtepjkDzRHBS8Kaf0aWxB56AKItcYPPOA
SWtQqHIv+0PA+UoFOHzPWOU7cS1vRQpbDQQY0ctn6vWi6wZjvFbWpcNDCCorRoEq
05sg1J2uuZ9rPG/nwuU866j5xt4AIGUGTTA5l3auIWaYI94WSHF5Pg0u59OTtJD1
nINEhrvpINOFP5O0vrKaCdYKfDBxAUg9L7UUU24yKYHK/hm9THTbfP8/xzrlDPHZ
J/kB+wskT9HfpnXfpiReXDBOFiNsVA0jEUxfYBHqh0zngJelmjAyeVrK1lrD36Sh
R9n2es5rJD8LocCSgbom6BIzhDBuFlUBDOZdwvNXdxv0v4I2uYu17TF9RKqC0QsY
D7FEdYX4TryJwRsdXh+BFBJg7qdChixBHCmmvnmp75H5o4wvMMatQz3r3Hz0j6rC
RwQ7T+jLCfymWifS0IrE8dfWnndfu5DDLFxxhuDVDi6H4XpEpB5HhevIkvERXJYE
yIxRbVDcWVnPFMtjMqgJ7P9J3JgkvFllDmQ32R2LjBDQJWvAkuvMIZvGoejSgt9W
tgxdBdAnHuo32aHV99Rh9rtOrrcE6Zvqot9pZjpdsqDtiFruo7VRgTK6bli8ZS24
8Ie7XequUojE9jKoXcjMpdmS032wCQE9WCRU8wErroS9Bzxo1jsVOx+LWz2ugjng
Ku9658443xhah7V7Rkbq4GRtxLCQbAPGi5BWE99a7GOC/cmTPrpXav/5pQ53utFV
gTwlHcn+mDSbgPs53pA3SLhQ4ZPopgmqPoUQJYdXfIut48+24XsYMhUvjCGsLUOK
MTYMTSgS0DixWe4GnrszTLR3Ba2WqZHQXFEN74ghbFKrjpz93L/44VwdqbphfgQ2
54TO/j9yN7ru50q+PRqWhA==
`pragma protect end_protected
