// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 01:23:58 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Pur2+bq6qU37x/CoWHxMfSLL3OfMCHntamuThIwiLAOmEMtfcryqK1yTfdaD9N3v
HLqCxbUGTUqhD+RfEMIAqAevTzbN+trkbkLOR9sWubiQNZlTSdIJBLDBx83v4z6B
92QJfdw3HX56E/4digGPohHR5AAwq5O+TBKgIGqbe7A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34464)
5WVmIMvuvs43dsw+yJkfnnGNUq7nVJv2DcYI99jYhQh06Q3mbOI4sRAI9AJ11NAP
x8eDA80YaktKsFUrzomC9jbH8VXFl2RiaspvalUUWvxOiqWIZjGzBWwJphFGsbk8
hsfMw3js/nLMMWd9rX1a96tNBnaOYlbbZ/V3WDjMn70bcTO+0w8AUHcemVkzkTTJ
3hbxNrb6IHXsp9WW17wSThdNvOTb8lJbfglM6dEBnsLf9TFvw5VJBE/nLFxzYN0d
au4MDEERF9rwgNwamWZU28/FWz7GT5xXbskNFt9h6+NHyIY1yBSLVHlxxh+iZIlh
YpmODI9swmPyM3Y/1fkF9l4MiferVvAa3eNMJsByYzau3nTB/lU0VUkvL72LnDvZ
bk9iJ//gXm8T3Zf8o0qBXahEnMNHslM/Iw6USeFAc6z9J1qJ5tYKYhlpMji2BSJX
wrNd2fu9UVJ7poB7xPD8+2J9kaXY1ye+8zA2olbQTu+7BkhV6zvJjhW6pS2ynv39
L+0Hr1Si1FKsP1d2oYha5Z4xrHKZzcOJ1P9prR6W11A9KamfMOMlJsvP2amI2e9z
6XLJVnZMpQpQnFJGpkrWWNu3HDIO/6VFv5c4hJMpe2ZDbAUWau9Fv8AHTu1GdYgK
UGE3B+3bRuHFkXcRFSeXSoBv7XOSUBxBGE4+dp0DUtbHDFlMj7P9B70sfvwgGX9j
iwkixauMDaQ1A+ZVKTpeR7keKmKXv2gjzNaFNLDHp8hYfyscWYzTAQf6BxRl1aXl
q32YXhql8Df3eCFT7mztAIHhzjjL7151j/PNs0/sdgLrUM8NzO7uZvU12mu9Fu8L
6p0jqF3X9uX84cY0NPAxk/NaA0VxHR+/R8fBSgSxCaOhpfjnwnIMJgTPq1ckrtNC
rVA1tWS5ZOZ7xeZ82rvjQtkb7EVeepskZlFp8LgToUH7M1niQEwtewP2NX4gSbIP
moGOdqWQ93ZEx6lkv0S2FFs5VL/8UROdFF8JHvK0ZZNOqJOoRufbNggkillBDzJA
ennkuF3VX9B+A8tE5ztotxLREuA3UFe+b4K07lXx7GqilN27t8VTvdmUU41KSiP+
kePjSL8acHWlgi46JazZgb8K2Z+Fq2QoTylrNcp1go6cYbbnhHRWa8gWwcBPPqcV
+vaHNcDOnkEX+xXAGmJaCkGN63fh8wX3YQ/PrRX/dWGAUXuaSn3iCpbcmspFnj1T
diQNvdUmiZSK+6bzuWs6XxeVZw2cLvAee7q9xJvwpVW51BWAWKs4BdVhXQSTjPl3
ehjLu7TzsqLVyz2uY9jbPNcYam7FBE3D6VgyPWLvQB/rpUfjC9pkEU30xzH6/vFJ
Jy8LDLSUtkAnrDzNlgAJNiCzHfVzvkFf7FPzbsUGFU+z7Tu/O3fwtJCMqGDnWXuA
Qe1B9KvvK3CWdvJoJCv1PTmHXUptKeNdnlZud48mSpS4G/u+djtBVERRTpFwWH8G
Kv6P7vNLqbn0QD/6hmLUAA/pudlI3aKccQn9rNIlCicmgYVUUO+kjsER0NPgXxrT
nMKFQ1jxqmBM0iLHZq1cE9RoCszWy0Y3yDAPN6MHtVmiEhWHRLhc8ExQrx/X5H1U
W1IcMqRdyhHu1WZkpXj8htISF05O06B7ukd2IX2FER8alaND18ibjfWr14dg8sM0
8+NvGy507oLjyJBA0enIScuTrreBZ1kCVuv27Jpn8+H2FH2YNloow+xlet/WD35j
G8fImBx1A7kxXw3grPEXZjHvg9xVZLYwZep4fmHD86YG7A7wxDI7KHbIJiZwOk1W
bmMhQBykrBOIO70FqnUC4OliJvEL7U1ARd8yeSrr6/z1vA2qwwqkKot6rgVUdYrE
ru1OtAGedXKLKIPfnqRy3EBly6FhwUrueA1w1DLuG0xWhFW9FzGjqY2w0f4d3Uxu
AA1E//g0AEHFicZWwfueyRVfxBRVC2RToDz8heI764HzDEfQkfb7RGDIfJ2CgOse
R88OXKEFtIp2f4w7rldlFkEa8yBBEjv7TTlKA9CQUIvj5j0x+vlTE+k/7p8/BxGS
ns+dc6TcmJPS4b2XFvjemBgjzNUEfOC9Kh7lJ9UVqPyGZ3RFpEZj0y1rM/OU3dP0
+vuRKIoaEkDBxlZmNUrLuAyiCLA7Z3b0YUO1VGTxCrhQXDQ7L8tP/JCo0NNR3cf7
YyL1JQUKOSNX3I3+SRsGruUqHPMsGZmVTdhWnzt3trcYhb3JgDH8Ksbwz2YsrYCd
aO3gumE+n99pfb1g5VqfC+qMRxjj21iCSbPb+VluQ+iExyb7a1bwxHgGCIMjHVAe
QekUJ3BypArCZdPkYG17fHWNI6NLfnPkJSgcWpYFBaqtvSs+KZnzoZVChZKYw2qw
aAbdBJ9u56iJOOXS3Ci3JK54BOKX0MDBJVguwuY8J1Ywx4dOOysPbCiz0YAOYGeu
WnbT9GhM8luWY0cUk1C5O1srHxAHesNbDfL2e2K4hIXbnVksZZYL950B2eZkMq7I
+Up/KZ08ik8fR0oHdoLoOkhKVArFO2vY9RLg23iGNVVGk/WWNNjJT1YOGKOgI4ZU
Lu2uoi05FU+6IUy35p4Al3cxetcPC8nkR+f4PWLq6CeMiporrppURMh/RAWenm8B
p8ei6roV+2ElH0UTYZCnOvCPSFvw7+HErwjIs6lvAKTOxd4JYMfKAJupbQtfWbCZ
Zx+Ht3fKnmU7XIzw1zHSF4c318EZL0WBGynM1qk31udFajRKVJGak/8NWBagjjfx
JyE1oz66qOZTapBq7dSs4gDq+HKDjkXSUaBwY0Fc2iaLwVGGyj7Wm/9fj9+EMJrO
FxuhvZ8eMFZoVmuoj5Cz5aW/8nZ47ZG69JUrhNL+fjJxZvGDrKTDpwu1a8dVLlQm
iRy7woO0vKUwr0UvZar+yoX7idl9i5yg4nOZw7VTwH7h6cXi68Hi0PKl9aEnrfoB
fNktY+PcjTfugC5dfRTGhjzENsFSMc2b0snCj8KuTfOqQlt2E4Ky0f4RooHecAd4
73vzJ/leUVkIdicxpgyA8Y28O+ZaDfJZfq50O9IGEUW0RHL/7F3b+BkyfBuGji2X
dZEEW20+BqtfxslGcQzXzyD6trt7Zs9LO1+SJ3c/L0ZuGou1Evezx//uPXURCmFy
iiDOgVTMzwAFrH+XiJEJ1YmOjDP9BcnpX0L5ldVYBhpbWeGLiSMuFySIZtX171GV
2kWyekbyGgl3wPchT7vXeeMzI5A1Szd1C5m48QTeyBTAntWO4imh7VWk8PG/gQJZ
0AdypCWYybs+HP9XnMLogUT8ah/WUAfH11CT3YnC0p42Hi7ktuVYkk5cgxyyvbfs
1GHmIPnhw9fIebpdV6lJ2646BaZNPsKZ/wkIpOptz3xfE0Gl8NOUNEg/7Jrm6Xvq
JngzklgN0Rodv19OZSwX3cBP2dx3AxUoxSlY8bNrdTWsS5zsYviJlyN4SEdYdvsa
zLdMu16xwmG1gCtaNrW7avGSQQR9pNHTAaoDKhXoq12XrvmzTqyV/5oLqZ7u4ggH
LSVvCdao7Sxq0R0MiD2bTL5nkbmR5eOU4XKsSbBIc+/UJUgRBpx7CS3jPIb/3Ak0
msw0x9oKFM4Bx8lDYqfzlySUT1O6mNA2/6BpRahYA90y9zPSYQhvrtelZI7BEdNC
pHX6zbAcSly0LBvTyhzwKzMKNPxA7PVepdh3/kgxHZKnyBqVS/KXG/T2lm0up+JU
Cu7vu00XBF2WI3St9SQxO9axrERN8Qr2K/DzTqv5McV4+9rwFQugN/k/UCH2s6qt
PWv4Wk83Dt26+cNlbl2qpWcLgobgr3KpPQhWGTPUpsxFVO1eOAaWkakeFOtKb8wa
v0xsGGVUv6bdnNZa89jncX/B3h95+7RODm39HWLtKyBtchEJJwlZvb6a+Qa7efYw
9uXARu2q0Vn/3E4PA8kJISY+8bm7QLGS0r/LLbPoRbUquP2zxYnOJbg+AmqIKhPE
L9CqNeYuUCdvY3qqM9uy8abR6s5/w8aBCXKFTfOE4HDVOrI6JGGSM4vv5O+HOllS
jRfTY5OU2nLxk7XA+sjlAG0lR8yZBXBiJyZywi3AUbTlNNJKwAhfYK9tMP2FfEDR
dPD3g2YzYjmChoAY74JmtaNeFyuGrczcZksA6k9RVfQuubErQYx8QkJITBhtTqYr
i3YaoUzAZ5NnZuy99hHvyJFv8sOf4g5eJ2hprRTmE4s6FNnvc6PMQXAE3RWb5yhP
5TiTxp2GCsjqpmfUNZgXkCP0XLPfSe6OWthpvU2kBVlqbY8cJylt5IdwFizWQstE
vxAXG/LPSRfcQ+ICEyKUZG+CPJvycJAeiIRE+KxLbpkPzZJVoFqFw5ILDq+C2D4b
c0z5/sPdWZ+F9GVniZJU/TwFc1/mIa/fGdlJ/t/halxJ19YOXEBOZ6R2GZEw02zF
8Dl+aixVOnxeqUFoggqqLVDLAFSUHqv4YXSv8aBd4PjuxaFHOGbthsGPoCZWuYBy
S56V7A4d7ze3e/a+33WqCf+Ne7NDUgSWcMVQioAlSy9b3JMxhVIpCnNZjIwQORNr
xYhTAj1VuxkFzt1rmBDKBw2DM22EFCXsUi5DD9Ybil3sX2dFklCxYiEB8MVCCd5p
HXsxbvBtrM17CC8RkwQ6NjFz0dDCKPuvpdlcOkTJEbuNugjvFQgtIoUD22jTVyPx
1GXTLiBja0DWcNWi4ayOckFId/b0Kh3spzt8rdKG4118SOQ1kdV0EfLUs3YuqFQv
nPqlaV75b8uTn37qSMiRSbucSR1/jTlroh/vH4z5N8HWN9fsuvz70FEQ2XhX28ij
t5Rp5g8AjoovzMek1uQYvEIh7e6TU19apv5y8h0+8BAvgrt+QfsyYi2FUmrzjzen
Evkm+ZLy8EwldcQ5MiDEJQMNVb5CgadL8F1i+5KmPJpUEnZBzXH8VDQDw5SU28U9
ByChYTbjo9GGnb/EH6lO13DFd/mtHb6yrs0bzW0Zp/MMAWhYh0brrdyo7f8e7zkP
tRUZZBKw+yVMpCc3AVhbmuaHn0K2ZFb6jUqAuRpKfnl734ER7klJ3JTIjIb7MBhb
emFZGgHUnZDCwBxqwEJ3PFyyZ3zX2+oBsYk/H1Pat3SBj+HQ6hhzJeQ00QMXYKp3
rNNvR0Cl5AOgKwo49GH3+EkuJ8k3S749x9wqIpkW32GoA5eeCxPEQyBN3jsjMfoH
zLThUXRr5sZ7aTuptJSnFOe/6/x7cjOMZ+oeJ3N6kFSrbPp9/VKe/45IEzy+ccrG
5v2BKATN6ONv2jNFGd7T8ixQn5KtfI1YYLfYbTOMrOX2mjsIZblHuDz8aT007IbK
dY08V0idYf1JCMdh+q4t5c/pPxEBofiDv9k+bZR9BDkzpsboTFMWC2N0tQHkd0Hb
YzdI4vRBW9RBsTI9idS5dgR5biEw3PAxFpJ6yqfCNcmR4S5czH6uF0F8EBkDrddr
rHL1dczUiIhOzwF63QoOF3KsZEqvTjNkN7qD/WIzJYaocfzrXu7/I0WqZR+Dk6Tx
McCrdTN8MVpfeNtzwZDbk2dR8JIjEud+4cknf6rGqtwXUCeLP4H+qDzS+0WLVmbp
JJ8M5wkGmvL7Tmd+pT9hc/ZQSdys6e+QRax/cpoo3wk5Y9/rjAtS9b6CdL7kZCmA
fGm1iLHyhrgsxgRG0uE6vwnF89Tm40GUDs7rb0eHMQ5Tcxqy5Rw9ax8pBPFHlPVq
CLXfB11Fqcj+1nfHFPdv8WeUbGKW5b+0K3qwbglWQnmTxNf7Oxnfa2lZ6A7n89UY
fCu4DFASi3Yu8Ix7n9/wR8Gm6WJlaOpPesRt+bTXrLrvQTV5rsRnkYMonP3Y2AeM
JAsYhRCA3tEQUTqdMhAebIZEUoRTqWWiIzw0usTglEzzTqx202kvC82fiJvaR1O1
pxf2GCT1deJ4+DNsz2DQwxadd7pqpDBWBFmk/iC2loKcdquYavgPh9++suKNj9Jy
OKqdT9TE54otJcP8yNDbKa8KQW909yvuoNXORJYoBm3IVkNvWaPin/GqFQDPSueu
xY3Tu6+7v8XHrksqCSpF2jSCQ1cS0v5Jj2edCVuGxupC9kaCkiZn62R8babsrwuJ
Qi4E6PsAHt40lOHJRxI1blw6Q0d7r6CAKQPGC3UKoJLXQS3ucowyArj7Ladi+Coo
SkEbhHgLdtnQAZXpifsVjuNGcMdPvebwAOTxQFQqh4APy4K/A8fFDuk1XyUtgam5
+yFiA2XF8ucsez4OmzUP/Gu44uA33CzbZ4U00fU5aaEEhP/vbSc2eJnHkNKHgbbt
y3K0fd0wgAFZRiBlbkyvQVrVv3LQmhX/BvPELyT1ZzxG/xjsQKxg/f+gsVXxCfBn
1jSdMKPJ2W/3KMRCgi55EHMnNSPZ2xtOOrtqZIZCaM6+oRLs/mCtUu2ytV6+x8Wi
/cWiD+2HK/roNrT//LpjoddYzmA62gJtl9Kd5NBZjoNnNAkY/m0EGpQdJfbZN1m8
3jG9OikjjENt/ciVisYr0FNVL2IuRa33wwV2FLSCugmWy1kQvGVNxfrXXeFKCqVU
MqmyUZiuc5HZAIvoLHEJZP2SHs541MgDNnlYhfdj5BeE30Pm54KvmD1dprH64Umv
oKVBvLnpNWncNvAT1PGdOVG2PrVhwJ2I/wxooifXMN+QCFVPNLh9uA1Gdp6Vg9ux
AQiMKsy7yz41ginC3HqH/6sqXKBF1/QaMXq9MgWaXiJhl53+YzNv7lDDn3R8AtDE
7FAt3+oV/aEoKLVaQ3nOKcxIFakxW/rz1O+IPele/OiN/DL5L2DYWzKEOg4XZNII
YBDJQ/z/y4+Md5Cqecs9N0Y5m315x6WD/9AWXNv3sioo60JjYTimCLOM7UM7LFbF
GLpv2HaQDpdbfezVqaSfC5Le2DmusmFMOFl90WtVfdwCv5oW8acKqt3Ij6ApqQvS
e9A3TZILg/W3/GLTSoPgZ/FYscfTX9PX+fZqiZH1r2x0d0L99r01M6sXkXvF8x4B
ooi7t497oMgaKoZtwgFYrqlTnimJyqjMpk0gIeANPIMeWMsOePBHpKJgzpo6PM1/
JI7FbJORzlY4AWrEjWhADIqnfl1OQXFnuGbX4BPkSOT/vvTvrY24xy9T0HZKFt/1
JTy1sywACqzIG4Px8n8DmmjaCgA1X09VrBgJW1lDRKLCI5l5aSdfchTbQzXPcHqj
cMo+7h2ke5tpNU1sqFv9mnEuKlUWJuraaNfuIChxKlG4pO0BVGJVbP1nyzEz3DKM
hSDRYKuhnCfoXK3Eio/P1UwqbUt/G4ukqKfu43qxbBZcx7wbaehpRuFDp9DuK8EO
XKh5d5/YtQVpInkBdGH/zXGLQNPba2OS5q3u/BFYbMs1flNVO1LEFBrIcLQjGoLO
1Dx3wULrlC90oyGZE1D7u/KwOaCgJr4yZVx7XWgVqCJufBC91YnM5wK095ppVRjA
pdnPdTUdQaR2zXgHE1UFADyhchGxapEYIemERQytMcoXKDSiAY1gxu1/oJuYbCky
/mwfdKoghHc0w4JInNuWGq1uQr8PFsEjrRZvGEq9crcpAAiIqpSr6JCsfvbhgVKJ
9W3qplnW+YaBA2OSfu3L3EY2wycjImzJFYfp0TowzTm5RC4eviueYQ5rqReyD16D
MfNb8rLJ6r9oTk3qopQIWHDWU+PCXL1hE80WPf1qmH2ZIKgPo14YiDfVyT3+LlhA
wBBCpUDsNlFjoGkh6djHocBDJZV4feFKB5Nwf/9VR4Z6nXrpi6qfhhsNdWDwslyE
g4b4aJE1xSc8/B91+1k+FNBPGRWwGuLraZOOBUbuIWSfadtYz2cta2dMPz4fz1ww
IjMNMBvLJ/w7Kxk9DLj65Z6Obi9wKfHKnRaGScU0OpClr1G0LOMQkT70uwuRvL3k
p16W9asbApQbxQn1HqQQ9AwpuIPH6tly1oWW40v5ZU2rVP0B2AlRJKJVT5CeVSx+
ylWcselgAK9pDvpAQMlzjuwRBX4bMLJd+lCdKujyGuuzD9RTQzEqJfDVkxum3Ty+
/zEKNGW4bitHfC1ZerzIIZuuVkWTAB2CUPvHxN9duJ+mcjWiofXxM9BX057ABNY7
VfFgtSrJAnSWjVSjJ3xwM/ajTLdf6gCwItrd/rJUjVz7ZLn8BRpe63kKDU66qh3s
cp2wxvVRpGMylf0QAB5cP7fSQaYk7bB6yd75tkpK+rxZSGpnPWL0vRgzAhGf/xl2
Dw2tvo99Q+2VRkBkI0lX4YWUUiSjZifsF7M0x2wD9Fp8iPyquHLH88SxUht1CH0l
hNlc60xTPsP2ilQhwGtXd38PX3ble8P8uKk2MUKSgLfX6R64RBTy5NObVvj9etCK
SGP0fcpvmlCbjnpMbOINUhpCC35mu1uBAvur6iVD5qqd6nPN7DYEm7KUBfFsA4J0
aIA6YNh5RHRscQE65m8mNYWta6OldQFcs2UP/mbS/tWJ7XXbtSrFKeeJ63jJ4MgM
aNhyPv+P+gXFZLzO1PS/TbLJD2n0xA/lS2+77KICdN9F/wNyzUS00O/arh5z7uxw
yZm7IuHEu5WNxmqQNVT2HWdnBJ1nyQu2yc4dQ4OzvNOk1cxzmWMaQB26dfBBrCom
byI/Lt3532DEiSxhRyS5tm8s3CYeRi4dO9sl26FALjGG6zDlbVZmQCzvsqNIFKkj
sUS2A6q9/KEi24joqJjPtB/GeTsxJxZpS2Dhwguv/M/CMfDLUdMrQ8h3V4763Kup
Mvo+IffCIONwusXXl5/NjH1TTR8iv0PAps7J7x4G6VJFz/Km5pkfqdHBU8q7av6t
xU6L5kwBZfShYL3mZCEjmutorXe9qNay4YABmGMPZfaxY5TvzoQd+2oRkp12hHuC
Jg0/OE+gxFL4sz4xM48dQYoalXwh18cpitEA7HIOMPyVFAUKzGG6aVC0wG5Cm9F3
L9GfczOsQwiWJotqjfNPDiVdc/5rkUgJGrMzlqs2VJLNd/uo8fWdJ6qetWnKsage
tutqL943J77FMHjxcInzqJOz03jc9uRke2y3sNQ4DfRaWIRDPUHzrZHeEGHkiavB
tDeOP6+zn4ysc0xMUi6O2MBYUXp6r4hqabpjeH71TbqGD2v65WqGpWykAp3A6ca/
qA3dTmmZ5eTH+jo439VZc5vXJvWODDjSYk928CtqAV5Tvsfifatm6Rq6Uhv67QVw
vi+ItmhkuSuCMwmPc8Z1Mh3T5+5gHMYSCCJxhhPLYltlw224+ETFVOXqHKycmXqk
0Z/9E2/JmlcgtnF6ZrYDpO5UJDrqiVBjgSU0DWvgXx77iCZCF5R3sswIEjzicl3Y
Ac2tzhMvySpyq1XOb6APffL5IAPTFVagkBtX1KkQjtsq+3WtUST6nxDPmjvpY5pB
tXUIOOFNABA34jPN/aG6HgoeWmG/wtGMZEAQyqv5DpuT8o5v9ag4O91LjGi4OL8s
M1nLQ/zt48X8PdOGbBpolrr7lVjb+BXa40GVxZTCKNfh/2Rx6mscjVmt3rXqziz6
fzV1IDOzFtnw5p7VktQiUT7E3JqAvoHTq1LWI7hm2lm8vM8wLCARBSW3HiQ2vKQH
gI/mgm+wpZFJ43IzCgTwZ6iozVmfFVo7sn2huz/xB67aJD4mJJePOEjS+2zVL8nu
1+VIrCDgmnUM6ibBadz2zAWoB53Zym08wC4dL06tWOaxo7HbUcivYe0hlCsxn1Em
AXJHercxEkNW1XVkSIqrfi5BCyUbI9JR5kyPCggAzs+1+tegZ0yiGoJgUd8+vhnP
hqzWtbr0/nriWDJelTI1bNGUy961vW2yblSD1tjc/8nouaxtx0WH+bHxLWuSKU02
CtRyAFNV8CtcDXw53d+o0wKMiCq7EG46R+dmBBkQVNM0bTTFX1AYnIA4p9rZiQ0a
mS9tDEkox/0iN8ekQvGSSff/l/CJEHuhFek97xLgQTg8inNKe3ona7+Ew/hxjhoc
vA0KpMJBiCLVwLEb4DkuvPbJ+/hg9c9HtaDxtMhZjeTz6sQ6JKwQf2NvswmPA+Fo
EpMkX1nSD0S6hnBdsvD1woHmtwtTzodPyjtCtkNt62yp6wFV4ebcnROHwZ/22nBd
y4y2aCKkejaj61CiLl8qse1V4MvlEP+QT5a8oP9ucHZbmWWHAXsiQgP76D+V5KlK
7TEyiUjY16Ho3L7GsTlMek3yopLbcMEwBaxx2/8FkH78rnKTH7YJV8BaAZiJFFdE
KKqi4FFofuR0h5TpEEMb2W6gqHCFH+Y4o8TqaLue/gy9Io3stpB7RhWNAy6R5UNw
T4kqCUy0W95lv/56qvAb647Oj1MrSh3OqXpW2V7cvXYaF6XST01kVIFncT7cwquj
FYrEhdmr/91DaIATXO24mugWV/798OmhtIdbry3F9zcEB/EvZ0PzXXXHrBhcWvwz
D9C9v7vuEgbemT+HMGdrfysa0FhUWcNvbhKc+hIeVCqW1zhszQjIXL1Y4llqEf6T
WCfIJnPlbRxpy1t4Zfb1B8LDdpAhw4E3pC6tjSJB72tyf1WHD9XhWNbZYsPdRtig
RhD8EOvOfX5Bh7hF7N7kVxrYEMZRjRE28YC+NPR/oCoJI3g018385VHSMXnATUJZ
D49LCiaiQ5KEDedMmnSKUyv/mS0MQ32jQpQ3MbG8bA784ZEnATLIdFJ6it87R+n1
+5xBThz39k7zEK6HxMxC2Z4w6eefssoKEO3CD1YY7MMndPxWO+Qu75gxn8e5NpBE
sX8eREX7F4DPaES13ItXKQVGBecOB+UgIyjoGHT4yDAJEYAfHRgsHZog3Aj4Y+uU
GBE04NU27Z9Fp+PLxELUQyNWnT39nfNvh2MHA7kbaYduu0L0r3RMmMerLDtJKicF
UYc+QqRdWFedFBChy5tWm7Oo1EF7cBTEVp21hxQFQJar1PEZ5osHQdVGPvdI5Eor
342gdo3lbqwdZJl3a4RPZKe9Rn2Ypdlj0DsgtrxS2y66qr80c1fvp7vCTL5IvDks
no1sIFci7JMyawjolRvxUNiCx6hnZn/nw+1KSffooR+ehamCTQ/RVgjbFDmXXTd8
FN3v0KuKbBWr4vKEEe/HaxLbt77BCr2//xC9/QcvyrqXO52LSQzjoq6bxOFXIJa2
ttNroIqmICBW7s6OD8NFquRkkCBL+11BM6MtwXLBpq8lpl4v1PJNKXvVL4yfUWx7
0ppK6nvgVwG4IfMuZWQAWxLe5u2RVVTnLjJuioiAB0s3REgVSzVgeCvR9NPLCJUP
kS0qSEh7dN4GkAqljcRZLm8U7PoWotgxAMbhDIoXA41UCIrpdWbpSuJr2IiLJz2r
9B2nanZgnDvlrC6UjrRUTYMfK143Z6wnBvFsIfOZeDKYInDjl3vzDUg3c+aU/Hj9
kpJmvWQ7RshQ4tsg0FIuyiRTBuf0MyHXsptpL2YfKHfFI+vHAkcjJAUjhLwNmnmc
zqkNdk6oY0YL69bnXo6r+H39684voLC/XWSh/yCvjH+m2LmmFXEdIymGf4pcCwp9
8OKjcwRmSBLKvm6ONlyydIEiu4CwiQJqUo6DeX81wUGbYkKS2neUfTVqunT21ih/
sAMpkTWC7X83EuY9TcOm5tKVjtzFCYiMG1NDOdeg1uMj10H5DtyOtxdGb6JujpP6
eagR0UVWCtCBnXVqSkCC10Zkro4/qo/RPoM8DSMTqkcbVEiITv28T2CeCjNUPUol
kS9PBcop0N72eku3w4J5VVq6hRcwmWdt26hIAXbWMU0eVgE6aPu4DnrFBkuIRl8i
uileznsIuFY26A7AKYqU4xCOulbDCOLJ/YWt0iUQyRYOgBeLy9xBz6tZ25WxnJae
eNBcBvxOLgTKv/K+Zk6PTVaTmjzEs+MGNbompmdHlDkz5wmXBCnMZ2F1ZijZJvSM
5M3KAvFBtYM1kicUfro+8VXtY82UZEZIxyXVZuVjf+31puzQVGNoIsIj+4QXLx9N
hTfnXGz+QqOirh+Qc8bKgxbhZtRqh5KPTbGd9dvYCcfnU2b0TbTV+m49LEYz7D/d
331TZ8Na1CojDlOZObvAWFEtyeBfAX1Vevy6ej9e7CifhInOvqm9X+4ohOuavphY
iDzCKXjRuaU5XCMV/AodXvZ4+7fPgGZAWNiONZkrwKq/T8/RnsRrib/5lE+OzEbw
nYqUk6xniMZQXN8Xhgoyms9iNc3JdB9Ux21MSDM+h2p4uAE8acGWr6NUHT88vgZX
0L9De2nQ6I7rcg0AWVWQmKVuQS3wMnlPKGYHYiDCI6Ixn9aI7zUTwbhB85kDP57i
gukP/4bExlL7UAWhQ2t/MO/bE/4PHtdIrBlIorF7XKNhmlmQlVl9sg9U5yNnBDWG
Gey7iCZWmTh/reQbXCJQViu+eTIrK0RRtWxvofPtRDUwbCdKCiyZPUVjvChKLjqb
UFxJ8YMMYPwkEzVgSD41Uc8ODKv4IgIyrpXqpLwSqaYLiCZ/7E8R5JVTci232HER
/FaBJHx32tiducUhzphteXDRrFzHH8g3KCfvShZj1c70wUjjgCn6zOJGPz4qRhg4
vyvbaIOj6svepZcAPEBks76P05PZ7t17ycH5Wsy5iq3o8Nj8XqKuwarNWk4uWJd8
sObyLdU4uarHvN3rNO8Y1GSRKp9qZ5pyB+GbN+AxavNYatDXzbMaYgeEoxYnwCoy
CcOMvPZkaKjEA0sPV1XIa81izHlAka4lBcZMlKdPyCp4rUfHg/Po5E7ZCKaW1Rt1
0FVtYyLroH4qbWDwypSMje1tHWnhZko8nfwa5tZy5d+w/N7SgYu8TFfjs2Sou+Te
Q9uPwLru2VILKX6itWbe1aZM4+8SJaRCrWkz+8+d0Lb2UjeeGgI9TtT10a2vIgby
OQN299MY9C0mdX0HO9kvicRRb08GTj/XcvM1GzQXOd8Lk6kzweoze8JTistNRhZb
bi0PVPQcpJt48mkLKK0Eq1AWfEABsuvExwDaJk96CVd+51+dGGFQdovx9BJbJjrQ
FCcNoNwO1R3xMGa4eC1nFpgorAMqektL0akTBY5BSchiErQhjYBKVq7F9wyVo7eQ
b/ZkeHQmEk3q/hVkx/R7NuFEQejmCQH713dGQ3k+/li739o+S525v/+/K1+uKF3+
hlAkOUELLCM8hnFM9b+mXVoM6GbQWqbc9noL5r/d3dQ/vkMGMCdnzjHN9xn9pUYJ
UpKeCH63xfrVMA0T+j9hwe5gChWAt8QdptLNRp1/Sbi7kp8YX+o39SFUVMDnzMuM
aQ1wuZQjjvBiIT1U1XrZzXab8acMt5quFtOc9zaxGddXrHEvw8zep1W61jdCUbz1
2WTR73/iVBDCFyDh556sNEUN/7W2APwdr/j/Psu55e6hfzn+bLyS8GXqOsAl5f1l
iqOhR4sHxyPcRKuVfDTECR1OcLxk/O8SXSLtkPf5SyJ8BPJ8fvNOVAKxPQoljPbR
PZwLCK9BFo2X8Wpe86VNnZsCjw+pJELDlzvhLcATfr8+Bt6Wy6h8d9B+NPwa8mut
a+22NEc70Xpi8TgXNzbW2zRKjgmJvBQ+bazugndaiC6ZE2x8b92k32UEdzlOUlyR
nhNhIE5s/3H+DfOBr6yQp4Pmz4p6zkiW2HWtjxVpVjs7h3rvrVO8tdNaRUBlfPQQ
spJECvJg3SyVGwz+LqrxBgynlQEdlRzoA11qofnwSCoF/6e4v9uhwQvsNhJxPaql
GwW2kNC/oKCGUzAdTy9peg0XFRIYjXe/M4PhLrOkdvOAs/xdp3RQkpR5MUFfn5kk
nD51h2Por28l6F5kQfUijWfPrplZId67ULZxwXFagqbs8/8i9XmawMMmxb0biAiY
HM0ptpveeIJttE+EF0R0uZovuzYWqO7b6WFSTnvq0Bu8iNfGvcIA7q1U8i9vqVpN
uk+JOFwgbYkyk4K5bY3DunphJpnF4EGiWd0+LA+fagakePddvQ6lBDvHUu5Zpkm7
mHx+/jZjK2MyUW2hR1z57g1Zuod1S851opfJXE7eK5tEqEuqf5X7/2zs9FUcMTBk
0vV6wJRkZSJaElM7Z60nTL5GBYo4L1RKeYnMNffZnHjCE0C/mNlFmHCukanoXDfb
z1lT0s/AVrkTZ0FLmn3+jXJh1SXP6nEcqyRst28ilk3r+5DvI54yHBzLich5zqMY
o5oW1DDdzw+EmijUuqRVFOTFRXPeTC9zG43jq6Zm02mrQmZHSMcWjSgnaliMg+ZQ
VpS51jzquU+H0zQjoCc5NMjnOAS+0Mo+Zn/8K8MMiXbES+6XUE4jD/zVGi+M4jmK
WA0p0Djsugi66Qa+EwQ9BeGkmVu40p3zzn+ItoYgaPiQmHc1qKAxS6vpWjwPVLKK
emo1BZpyzWO4fohHoxSIn4g6/8nej9V4c+5HuYNn40ZiSWLbRVNJnh0Y8b3q619M
BYEzVihUxQLsFsaY7bxTrSGpQKu7Zft2F+PyPDF8uQ+BjC2rfocxpbY78qi/XJeO
9a3CHIGfXP9DAfyKBvZslr6bVfsdzJy+ltn0DmKyAsxe2xZb6jnSjM3jWXVSPckp
TI+wOt3XzSoQGbAnUPPRGE+UBcKWPGFeChD0x81c/PW6wIEyX40keaMb071E/dyj
B3c3ZDyh7GUyuhbM2w5C3WziMecAYeFSjRd+u0aC6Le9Y79aVSG7W7LH1GUvQOEB
a+Fnp2UDpqwNvBxwYc1Maels0BuvS7cUekP3ZshrFXVgrReMnMQjxbk04H5oEUiz
fvxoYrh3aRSYv8kDDzNy/6Dkw/ujfOqhpLwkMalUvrB55tgQqaPsnu6t9/KS8F8j
OOKSnJOXMLPnBoCLc28XZFFVJIYQYFX1E8l1GGZ125pb6AKr/seD/ZytdAeZNuVZ
wvht549N9XgldnKJAXXr2+Bwb0uDP13wlw0ZZPeduBicpFgSafPomXwsmKsVDjVe
PfVVr2lUIG0YzSZyIOSuaCV6iiEjMAoSW5WoEZxdi1UpWP1UV3QCKUNwtcwPYgag
Ns4jpjSw2XdT5neSDLb3Yr38XoiLQW305OCKIt/sNG8I85FymsUMlc3ci/lDfJP3
cJnZau6keCczB8mttoE/gQ0hObYYHQTRr+RDrFJQ8nSUsDMkoeojM6FsrXcgu2Jh
QgpeCxi0YKUbBB8aYS9LxDco8WWUl7eT5y1r+hEsYSmcpXv4ViLJw4CWAqzidnY1
Qpk6nJSEGfDNl+cd+hdHQVlfXQojR87lrNtkmXWQKspwPo6CShJ4LeqlseBf5UTV
mQ3vcCvf6Gjd4sahLaQ1nYj/p8IUnGCq1KZ0Q2QNF6DHSwjQRzCdPUTwoFXg+RRX
945W2R1e+re/KMEW8EVTK0HGjIAuGLboxDJeRnTcnTDrkVQEhM8zQeGprCRyJ4E+
qGaAnxUGCPnQgMrVLTBNbeokz955CWYxJ0pzyhSHBRib91mwCL+BnAPmq6X5gw5k
sJovAXIbQVqLYVKuPbrXeE9cczt+KaOt/ZGCNi7WenM/djO1UBZliiCz5kNIX+NH
sFzLK9qvbVgmtFB4LewK8Z7EsX07k/OXMM1DzuXSBcnLGK6WYU3/RGsPT1Nhs9Xb
r8mCMiOd7DQCkHEJM6fEcBtzQnGDud2Zp3sLM8qS+JMqyDuN3c/6GUhCGsX/ccAE
r7gza5rbqzWoc4yKPU+wx7xG1nSqvFTCJqXHGAxRI9tZBdp3ZRC/4NFES4EpD4ys
40dEc/wfeIwaenGn4chtseFyhIEIY4py6j1Ka31TrOJI3pLBba3nKkmh15zBTDvq
zEfw/1w1iPKIrmX+ZR2qlq88Odlgld0VQa/BriUuR9a5uzUQl84FKyZ7TDD0A7iw
QAlhAb2tIIxRvdAFb6fKf/V/VxFxhvV1Fj+0nLd7dGj4rcW0AkG9O/DiW+u7A0yr
lS+O26Fk9EUQmLMEEP0mEOQArUR5LvGefZPAmVHebeA4bceQYudEJg2/ZVu/Xbzf
ZQLwIephLBBsK6Naq18348xNWHv0b54fctJCa+qKc6cUI5axamflPp0CYCI8nR1a
eGpm0C8ezkG/zFydRABX9UvpgfzJf3fw7zF2LediOhujQgLWJSXzcr/z2XiQVe56
1tTSyUgB7kw/AFCtW4RFvggQaQG9rP/4649BC33iPIAw9hTnb9jj6bLKhaqf+7o6
S6n3SJRLpjBchdzDwhpIoUgZ7ZWidxyIa0a+oHL6QPIwKQS5EtSRLoK0etRatKmH
iPK7jGxxhszBpmTe2WRXzCUQAkRggqAykQrwe/Niy/zEE6RQRyELoqB0httJ0AG7
FEVNyVkwCmHFvSbXdpmmD2XtCMyx/e/SpIDx49FvS1oSG8HpzXh2Fuf2TUTbJz1r
a6SlKBGQ4AudYR5vwetZqdoRXDUhdFrNhtXMpcfJDgftjRADh6g34dhN5JoJMAHA
rO4zWmyv74dzluFKiUKxEMgNkzP0TYRvIO74w7FTgdmm4RUgNebVwgRfhPUKJj2H
5OzHiX/s0PK+6iODgc4bGYXDIN2TqVqAaz2z3VZaGzC+phQP5j/oyE1266bUYk/g
fHjVJVc+igVwZ0pi/biEtPTsBg0BLps1bCx7E1uIGdMa3X46XypGnVDt57OhM+Ov
e5xFtZ8CYA6o/QbfJiT++Ypshp47ClynzajSwmeVzZ/X7G8FHtPJqTQqYojycToc
cfSf26O7YCxyoqt23hrVAmCOOjiPP+Zeya2ejRGFi0v/eRaPP+K8/rVyVN5aJhhd
Q6mE/obr+HXhL8Cg29Jo/vZFCAD8o4zq3oo4FAIrkXAhLLUSTxeNJg8sJftwBqIf
GPCzyNTAFrXKHJ4VN8AhaR3vWuyjxWQUGDFiXgc9YSuZK9OzERYWoOg2sDRQvpdi
tKR+d7toDUn5pfG2TcwCb3FUx4pnDh9PRg0YtXPaJrcnlFHqVQFxKm5IHw3h+T8j
47UHCesls4prp4CYcTfR38qj7Os7EGCWnXi11Hx2GVd2oo8CIW5v5c/hF1V13W4F
H4CoA1+yvuwgGM3uY8gr4HhuXJwsdksDPLlrr+4E9680KNPz1MaBedJvnPm+PJLT
ub3x1HblZDnmCaXlVOPf8UVPvyxKTZBpVQKcxzozhw3JNwhqjDaIu6jjNAycarkS
nsa5GuMF/t4rNCQnKAkaUpA0d0VMYtltu6OfUJFdvLabJ32v/mUIrkLwyekJVmOd
0M3Yf3slzRaFE/cGSKB4bESubP3zZQnd7qg33joPSPA6blvGuGUlZFwJJ8ke/VLH
Fo50W9/OImg6N6nIIkyoBdw+xJqgmxX8tV9ntSnGR0nBAfhNdF5R/p/aFcCwGCHM
PibYHCGjNY/rNMDDT/CQA7lwz5mDoVPVmYxKU8NRffOvRUVXgg0Bwk3WaUdXWFTU
UNZntHDP2fSFS1M88EtKnaEmEaJESf17yZ/6/gAPcu1Ucfzzf58oUtQWnpdVkco/
t+eSkWfGNhhebmblqRnjSfEpaExRfFcjEo0ilNfhzUrzugjbEY8oNCUljdgXZk4e
9xgfz79GcwIBaz5m5C0D0jH4fDrPTBFl/xeJeRXC+X6oxViXTp1AQFVWlz1EHvq0
bZ4BE/uFsL0CSl3Z/qupECY4w02cOxXcesQZaj++HjS54sSly96jH/7LKfPKxSiw
CUgShgE4l/LpXAnGw9zv0sAs6i4VXOYQWoMs2hBXKQFWuVgsafNJLQ2g5ZLGyu3N
vtpmdlR6c8oRIeYgE44o4WyUn+quq32l8Ta/VOpUkdDg4baM3FHMctg0UyK8Ngzh
zOJuKEr2Y7Oce2ejJttWtSD575lYildxfPbKUc6JH0pzlDJxNFiAsOim1a9zbz2P
IOn4sokjuP68mh7/RjiOY/fNVzWFpCah8M5cwkkxTOUMRaB/wxgBTg1TLlVoc8Ny
e5nlbMat3rdLxMlGq/p8az0oGSZEOIp83EGW7EHEfFwVklLQuH7Gsj/aOpd+Tqam
isE3udPllhw9fSE96IGwOumvSUdA3FNfkrTp69pXMkLNtXmcU5mF/zAOUQ4CPRFO
WvcSDvPhJ+dHV2EAmkTIya0O8UqUdRMPU7Ypv08sRg+SOx60vhahvMUhCYPznnbA
jBktssEbf3JwEEj2qGYmpEpXf4iK/EedtZKGbCuYrHMaDTUSQ83F0mIKWUbzNR7C
lid2PGvYUPhD/yy4oskvtaS26LQ13TFbaAMDQLjbdgOE9te3zwBokk7ZPYyXg16l
Pdij81hPzXcp7XY/a+YIWBBYHlmn46wilyteURnIBIZzvWOEMmYxDr1uV3EyJEjg
d+X4u1lsdFg1aDMMwhznC8e/AWzLovDd3fCWua2KPvOl5TzZH38sy52uZpaAUi42
0PEM/+uCVZWYvcYWQ1i3g0IGFeEk03xKS9nft/2gvO+resAwEybfrFVNZRyNQQ7i
PKAxMa3Rat3DmgOYYwSYPdgYxVcK1zuwfRO3NzPHnfMnLP0dBgaI9dARvz2XRQ35
xzfvDDgcL01+td/GWpCEo9AxHKeG8k77XCXumYNe3ENQojSK4rAIYumRBR39y1Fp
7fzdCTkkDXKFBnYUfe4fIOSK6acaOg1OPfHhpSs72+lJTuNn57GschUP1Ww6FXt7
nv8BDoXhpXQDtFpjURA1e+fcQDj+gRDFnQUJQfjjwUPfFo/12NI1LiwprAdzQr4+
oOWdVDGiz368uWoInP4GLMfSKTFFGmS8K1LZQ1AjwdzxX0D6GsFZ5Pb/SI1A5z7X
sDxV3cSI3r6JXNwwlRgswQsWyEXtmzpxsj3iYtnhzYSoNNEpVqxI9dCzWhsk40RC
V9ycUb9SvjiReg3zANNX0DP+Dcot9F3sUvSJc+V55SawXlAduOyJOiCGfypVJGZ0
hkx3aQljHDuHVucQ+Ygp7JNL0SvER/9U/WVm2KCrvYRvkaIuXq4JaDxhrd6b/aYD
On97MZs0SFHr/n7Ni5VBUcT74dOMfZu0P9kSER2Pg0ELGQ88teunxLYJSIKD+k51
Y2UA7bdEpxhiDEEZtil5DQJU61uxtQEgNdIAmvX7nldrt4qfYoHFtlWGz8QoG0Pa
ux38axWYUywXDhMfPp5ZCD9EnFvsnE2h4Sl1PYKDHBQcuzV7FXsJstKoyAaeyUSs
dCXJyNCMH1SCGo9wLYQP8H+umhvaCFWPLCdy2Vr2cgCQjSgr3yqtX0S+BWacenyC
nQdxp9joxZq6vrjY6yG/AG5DypzQ61yOxIvPyhs0VIOOymU3aMbF4O6CoI196B7I
Ez9mhclJzrcWYhP+rvDFOlRtDNorLJezhLEHP6R1yg1PJ1QbNxeXRfIdIYLywmgW
D8csJDo7sweAbe5I1KlIEAUYKFivzjiklpY4TUMWYj0IMm7FQYMFflUuCRLe3hIx
l5sqL6uHxh//zgnl74Q28kr2Xj1y9R/RIv6p6WWedSA7LOg/4ct7bsWR74Xl0u8r
vG2mOAPlwJTBDBaSBrFNVxP7f4/pU4HZzedmufA0pbwNOBZH5knhkdsKJEtcjD1i
cOq0Ts46D5AG/KpKvvb5zu6o+koMCgDL31Ktxgalx2BZ2xjbuF0eLMAZDNjeaCNR
73vjQ9ByPFPBhEnq/uaMJYji1UVrNLYrY6Xt96YD5Eo9T9+89wrkYRO97HrADlIe
L729IP4CRSDx3wqgzpMD7dOSK682gryDKUBsr50RDOV/mORnEeLHZQP5SPrpTq7Z
bX0op4JXyEBMyGPkijmP0LhVful6bq+6cq5C8uhCDcE0rU1mS5ycglhwEJDBh2mB
oFGkIahitDEWcREEGqu3jFS/o2lg3VjrR9U+n2b4p+BTqunDyxGEWNEu28QVei62
Rrm5AmRyKBfkkNJCVlHXkuvnKYzUKMfWHHMXKaEggtxu882YIANxnUKIbS1tsVKL
hu2IDDSfKKb415en3hMa3soxb8cXa46TeH14nr5HLeiJYgOzKjVwhe/yAwt8dzfv
3cpN6/qVmBhQaFt4BSE04hzwQQ+3/OkTPYz6FBBXPDDoCUwQO+g5s0vfUaNOhjNo
qRGuOuBI5+rDtycP68W0ta+lWJvK7gm7LMIqrIoPAfyK8xKD/zWHfmDyeSnAQoPL
3gXe6oDWbzyAK8OWDr/mm4T+X39dne16F49A9hz6ulWiFbc/qjlisc/Ydo+tUcBe
8mQD0MbAgH4cr94ns5vq6UjwPTrDyaH90llxGDTTzAsLrRWxvAA5FBuT+o0lJ9yZ
Fc7isIsSj9HkMtHaBUO/TPEWEvFiae7tp0PB0jJIfpdcHyQ0mPBmJtK+dZD9kdkE
njtkO8actIjeTDVyAcFdaMdyUnivKEvUesHdPhjgrhtrQOTuE+reG1E1EJOy+O4c
e531xACaTSb98H5J7nDJ7f86p//T/dYGwGWWlMragvytPi0kk/kTtYjA28A6WHuJ
xLt4lX1I5gKaATKyDn6BHYs4ayQg8mm2fC15SATudExYXlnv0hHNqWbjdEcoTJ5w
UEex+R9KP7OqtCpnp1xJ93kSmkuyAf+pCosItacFvjqMxHGm8W9+K3tFUVaX6Lav
UHPt1udwF1pVE97A2sQHijd9mGEVThuI1LKRf944hwIPmgZS/jcFiKJB2WYu0dq4
afjGs9bSbifE0ltqUrjWxDmVAtrjB5lBdNrSO9jnxLeA69L0WtY2VYMXSOrVNXqy
UU+HHVE+RE8S6180TG/mfLC0MtDpD1CR8Jy4+1jDsYF5guOaaP+0Xt/AnMFKLFJL
vrh5nhNdPjFAHRIChQtSTOkfBaQLzwERzBkoLYm983FR1ggbT1qM0Ew2teOR95YV
IOemM9b8uV2dceRUd79H1rL0lFXsTCMJjTc79NMCqKwOpiQtdLIXXcxUs5IEdtyy
qisXqaEmWS5SJ4HxxXtA52GztkwZQTVCy/sKieBEONpGm1h7BuR6yD3N9Vykv80L
q45mgVYHFZreUOoaYvOmJKYesbaTZ1BwYiSH0tbMbxm6miHTneSrljIje9Y1BMXm
cuEKIMRMbpN6P0AOHOtbUTQiGmzSRBdz6g5hL5hcflTBmYHBiczt6Mtzs+yEeHfu
kEyOwGlpyAk3RVOx5/pYyf6CAFUUz7JtWp46IbIooMMRFEdw9QeFQ8konEcCrTWl
J/NLNN+lE5jZjvfVgEO3bphemurVFse8aI26/1f3B+z9yqtcy/4ZA/lCdlFaXnLa
sFFmXUUdG4saHV5HWhiPrvDD9lEuErApYudJdqcI84PmYYk1WcSPjyNw6grh8kwM
dCyZwuOu27hwOsuUV3dHYG75cOA/FdmBeRYpdC+ShBoNfVVfXtdXvpoxG+p9yel7
bx+D3adtbbVHAMCeH/7CCdgrlNuk3+Da2K/d2fOFmhHgUnbpJP8c/Qi8P6ldInWP
yCVf55TQAnGCsPN+HZ7YcmdykvjySBXqLUVX11ee67XV2rV7LkxYDgQBDusMzmJ2
Z90VbhXJ/PvmpWLwO285vobn6ffaOU1vnBeVF8MDNSpu69MNJgJ4zjOtRjhq2554
TIQK+SgWok0DXF3m4xk3PV5JGqAhlwFyrG5Z6nbYFeqF0dTRBpTCnYzH6YkPaHUo
xZuldmbWm6f6/aee6oCZC7a2onRoFoSs4qNRtakWbt+XhzN/UfkCcKLPYzxzNyYE
xzDWtzAGBYoAh/+M3IGgC5hUDoOo29yjWqNWFa1KXafVfoHek18qMDTr4DlOkv7C
gmOXlTyeXbjIYGSBQ8H9YtX+a7qMsyzUL328memmtjZwlcv/1T4173ptXp+ojt4/
uZr7NuuQixJ2BlLO3Mmu84AdqjZrM2UXku5rZl/EHVhpoxyOrjg3TyWIi+UhC9Ji
cwvq5nGQ/FH5ZjhE/IVu1ML5Brgh4FG/UcY50q/fYVvvXw3EcaJMfgOSyZ41/5mC
XtE9JPG4AIB/mobDJR5wfxVPKvlEdaW9IcEqvIcNVYA4h5/z5MbmRVRuermVlpB4
Ru8zaVkAyhwSbVyZcG1glNUr9FA7hOfLtg/WSg5lBi+wAPIuRYHNmyk/cp1IsXro
ZEP6nGWww8QJT3BS+a3HmpyQ2JCE98RpEjGeKwmgtIgS31TgoFNejJQzyfn7sn4h
vVzWNZ6ryyTbsbn05oHloKe6uF0t0Fkvb+QnxSmgMPjOrQToReTVDZVBM4ff9UCc
Hhdf4Pb72hlLzsFA/C0xtVWDfgR4GckpPDgoO4lG3LgpPR6alpk4dcLiFfuE7bEg
cbo9WrkwiVj41r32b5AmjmbgUITQptSL5y1WKgINtx4JsjMlHzK8y9ddmDISlFhX
D10c0zcxrFzvaUfYXrBwPIPgBJ3aZ/XgNMnY68yiIoorPa6R9InVBcUKw9cO88a4
VogWjZcjcHNvl4hTB/O2C0f0tplgcb3KZGsZOn8kwOndIz+WRM4JBXyVZ2PfF+g0
gCRousn4Mf6qYjZRh86ii39ob1sXMqollYOrPnsIgoW93PGuWlo+Ev1Ci0rMLfuJ
TglfqB8OocByPeEbChCO/YrEVxXm3lK0NGsrFOG3w2kOCaJ8+MFlRklnjx6kDiOC
pwkV15mvZyqz6z/vZa8zTyXmxbUdcrW4Js7kViRQwJZbIGl4jaISpFU/GzGWFylQ
nL0xC32RYPu/NvMZin4A3evpxhKRhU1rCOL0UDjFjoIP5DB8UgnyJ84pRScEssj3
y1tUVcoV0vD65NN+y3kxu4Hccrdkbg9BY4uvEag52KxYYoH7nzh2VrwWb/zcPJno
4/Ubbf0rhazFiF/FySDBn3vZLXvj/E+LZ3uOottVdpRlREnSicbUlXkGwoxbwGVJ
8IATEEbQmb1rjRvq94mNEJeMrPpyft4C/AqDYRK6oEY6pL9qSFVAk8+pgkZg1n2o
gFOulIuf28kmc4QpxF3rjIGRUGfxCgceum9AdH0YJf+aBiz5HGBENyoex+QBjXcV
I59+xdpM9mAfp4Qd1/Nfg7O8K7amriUBw0LFKTGbsx18CQ41fRJeSxKbCooF0f7L
bzyQf6ThtFrFkJDfDF2Sb/luLTssBj7ukNzaw32vamO7JM9gExEpLcyav+/Wc0pI
h3SfY3gjAkCUKLMhPCFWLTmLszo2JRF6H+xZGJB777O4+C+QGrG5F2Xl9KUz3hyD
9vBRhv2sHCh8dmPrzFy0aUJw3fN7QGi/GrAO+fp9btA17+1tp1gyGyUcp9GtgdzJ
954WCJHzEpwy/V+vPkwM7Ah++HeSwxe/bJAppON5Fvucj6iAjRJUzhyc8IgWQUF+
qqogL++qDidJ5eTFWYvY1+XPzKbqnez3/aqsf7ydgeFFA3ginBdVqxcd8aPvFLrM
GmLGBZJTNiPbv5tLjuq8Z3J2K0dDqwIL4t6QEW2Kbuw4rWrN0bVuXgCYbDGnbR4T
PXerfBb2mfEfl90tlGxrTnzwfmXmUkmekw4mseQQpQfb18puUbwM2Jyk1Kz/WywH
FkCFnPcfLXpupwXnoNFgGMzSk9hSOcJmA6qDrJTLwjF6DUJeKqeqvmEla49A5Ith
qb7wtQuNPFOU0pnt7+KJLwHtin2Nx1ozR5qmny0Mt8QaFH7keo7Z0LfKNPuDesGB
dearvX+Od7v3kWlF/OG6tl0ct2X/iKStnwxbK39ch5D4mZH7UsHOb/uP7dh6trwp
93tTOwTGRl3vDUhekWJ40PADtVwwbFIpfh6neklAUfujbDDn+4PS3uAF9skTCuIL
uGub+9Do11NFquAysvAAhWwilCO9KkJKiPz4UcJVwkOqW66aud/1Bo8RK8j4pnHL
AHrnXM7cPGSkSMUowujFHzo/1iexWuFQKnmfpBfmUyyXM99QyTnMP/MzTDQVBL6L
ZObPTtHBPTZXCYw76bWKS5xnumdJbnDqj9pd5E3apqFDyFA0VUfkf35WA6DvAZy2
TNyvAbRmrjJdaasHe7bkFXmD1POO9FQ/PdAwRM1dKkVoyX/R2CT2USgob1J4WBy1
6Mm9qLurmNzkUf3dD9aqx3531Mqy+XBiw2zRXWaD610Q/rVNn3hjNyor+7yLEvYU
O8TOTaIJ8r3cAnqbkaABELla5WUxz++8kMIBKwGpa2fX3jEJOmP95PucFnMFHoDd
qtTBPuEnFcvMwG9oLSrR1XYQbKArIHtgrzER3dWDWkQYUcWknWiq4ukKWVtmW58q
L2fnSaKNuGoPWcvQAdPhXORqs6clSKl2SmVuxfDKjgNfoiqNwr/BT3kM+4KHdliq
sPInS9g+NmMm3YOU89Ro9Gh9hFYQ03alZHPSsy1/7ZLoMouA9aKYFvPCwCz3fVIz
hkSQxM+46PUViQ9LYN4fFXDt7mcN0TFo3aEOehKRDJYE/fXbM/tMOuJfbo/TeBJ5
DGNmP7fsaz2a0bQ36Jyh2c6mT6LGH7CHakGoUv3qPnvBE/sUP/F0Vhg2FKu52HZy
xWIiT6X0Pmgv0lRBFxYgrT80jpyc8pDlQSNYGmcCoNej7+WxoLMLSGNcU7cHj7fN
zEMRiSCWMEk48O5lQrtU9l/3y0eT5f7FiXJY4PUZxho2FReqeNxwS+zM3zRgueqC
JrVA6YV0nBdoFSdKol/fGsbetd1Az/36YfSjREjCgxv2neqy1OBpAQA1GVP4u/9V
/srYIIibrrMQNvpBmp3iXZsiudI7139M2dMrt417t9I9XR+QMMs5DuO0UDsEHK3l
AdHRs9KTAfTHY3/cc0m7EluUtoYXj4Te96tJY5ATG4KOSK8EcpaqIkqCFrErWJBx
Y2bhVj7TIZQdN41mH09oLvKg5GtzUraWV+jIbaveUhbJ2m1Bmq8pFwkzR9EEKLAT
noAA9a8sJXQEbj7vXDTIvVPP2b7mdtfp6+hAr6zFpYh9a0WCQEmbVlCzloyIKz6v
RktEQzKfFhYLaQOJJzeWQjVmuWTX9FfOd5yvlmmPdszP8RICx0AuJrAYZ0+hr0jN
z9VcbEj/SNWEdpQWw7meL3B9MknV5VkiCn7Jnvf5SaJ6BeMQmhWNsyXGqtF6bC9B
Xae0tloqYSUUUiYr3TpJR+cQqFb5OngiirWpMtpO3VeOwe4fLV/+Sbr7D+bf1zdZ
aLp8FSnaLejeusKOjFkaJjdscXFz4Sla54u0tleYWYBW1euYwCi7VOwYcJrrNj75
KfZPwVSgTb4cKS31gIvqcytWZzKwSDND3b6hUTPL/WkQd4lgQBo/ENxWzxYHjyvO
uysRsG/6/oLO444DakFx0xFrarwob5WPAux7Bt/hqhXBNhtkyqeqXdURsV5BuDu5
EKUWjUGc8tVWYzPVu5ZsqFHf4ec3a7qvw2Yo3/GsB54vPHIaqtikRCL0yhsRKtqf
bb32gXQ3o+Z8ocSAsQFbmWL87iP3BZbkBTYcwxP84zyLS7a3FUCtETBFtjyMUgGz
mYlf1BuexqKwf8B+OFgrFxpOdS/gj64BM/KaFpKcvoVMBoE3ME13+NMQPxYOWVlY
ngNULuXV5NH+6WButiX8l/uVy8rKL2IwmY1R1zaWtEb34TqqZ2suQb9ckvdSD6mT
Bn9ZsPim5hk7/SWo0JeWjMXmwqbhjLXNzOHYV/RA4qjOsIs+ZMlgpOaXzwDwjKW6
+ppnVimJdkANO082Nqv7W1GNPrsrvn0wGivqITtm9t0nlu0+qOa7HdjRQFeIxxdA
vlXEQj2PZ1mv6U6tBz4/K8sIoKkd8rc5QwSAlLjLFpE/YvdsIw3xXyu/R7Qx7CsY
jZURxX82woftrhMIz4y88+WqIqvxxxOkhz3KEMcEJm/HqaCqBJsETPV0iqkLlUWv
7UTJxpoJWc/VmfzbHv+Dr40Iky6rHmJuUuEvKu5A6WFoqIj7QnyFjpmEgc0avAy2
IcjjducuMHPYdNBtzVPRMEMKbIWvo48qWb6BrsJ98mAmTe63s5GwhGJIIlkauP7B
jiPm35appUQjBfroQHzim9kYIwnoPskbfWlEfU4i+qxJtVHJyBNarEqSoSd4D+J2
AMGNQdcStje4g7Hu4d1PRknn/rOZPCq1Ovnz9k4NamJzRhIrLMVAQ4lFiQFW2727
7HJDvvMZ2t5MgIkqEy/Wpj2ePwqe3HV8LBrZzFDy0HVVRdsJXDngkK2vLO/qywTJ
zlk9hsbuL7ZoXZ2QaK78d+aYUtXpj9aCOH4ze3pMjIecN4RGxbxXmjygglsvAtI/
I4ALs17+pS5elMmOMBuCvr7YDXl1o89HYH/pQKWa7/sB9i3HokS2ekP6pbr6x3Wo
LvIpQYwJ0FRUrYoPwpUe8be7uIDLBU9cbqnCCVXp6IsshT9br8Ya4Y+GL1jL69wx
ErOXiJr9C7gd92SfczKqrarR4CQykrhJOPuRNzy6Tz2dVoTLxqUW8Ur9ZDT7KlCD
gCHGsEJ+kpYNxaUt/9UUU9GHORU5RIl3veQpQUOU6p1GRoJTjkhBNV8fl+++VyZj
70yPTz90WYEk1zpVvB9yuPAmLNe+EbEMhOEdzWqTNpf2MhdlIzQJud/hyyLxsMif
JFlFuf/pL1giqprcK6L1M4jbX3fNlhCnSg3N8M3im7gYsEutDSbji2wfNQSV4ZL5
B5KhMCXFStbjwLFe/m3VbZct1BnZERsZ6Q1Yu9r24ZMjUuiHBwFp+ArJ4mxZdXZ0
sASy2zfYxAZwFjDFqTY4HafMPvDbG3UbfOANEnNuPp5cz15jY73pbPgk0s3CoteO
9QOMgjAs5Y67bNHPl6ACQ47RIR7g0yRJyRswwU3k496UIQhfbSl/vZv88eJPjvmX
mougYgWHN7GROgFoHlXqqjI8XGKzy1t1XtpxZSWs/AvW5OYHhxvpO7qN58dL3Irn
L7sNL9wo2eCa8lGmFfqZGjVc/r5H6X7Fjak23P7m/FRV7WyqKw9vlWUowYWBpM7S
Rok4GtluVQnNAY7ibKq1CRO4SIsX8E90sQwAQ850bpsYfbe1B6MVaHxpMDowg30E
xNoBFsrrdUoAjhq2UHEIeqF7Uvks+GudX9qqnqp9dV6xknKRloVM9mZFXkjBcCgs
fXQyJYx+Fjd36o+dCdylo0tTT7abDMFKlQun7SJ3CQBJBezjwUh+GEkuURATcvr0
djrJ4zaEO07I/DKW4FY3Xq1uuczbMB83ALdGNOtqGAPoXsFIC7ArBxtOL/TFpHl+
ua7RwYdHGxkvf1aPsv8rB5Foojf+6Gvh29wouWEEysbYC748HLWjLjWi7K5V/iPN
/1flpelItyn1eIvz+jWxmGkMGKA+MHPcOMQmX2ZMlToeMSb99f5QI56gXhWpeSJd
pVbVzZrVaK9yQCFpeFaGowVRrFWYvnb+2l/GIZ2stPVmMJhH996IjmQnmd4M1KP7
hBGqq5vhervtpoli9WN94XcZ1EJmgnsfEI7fNpdOCzRrjgIgTjC8A5cXXss5fwic
BwOy9zVlw1sAlS48LWNMgtN3DjDFthyw1MYcD+aptac4ASr5D95Evb4D5uKgYyjV
HnItMrBx/4I/MkWJwv8UReK3ywYPvON648BTMu/56oA19iOEGrX6AWh0At8Pb7bs
FEJS6ZMjvhRtH+1eEyFAcj9P+yAPfYS6MY1UBtPhNjENDJfIiGtZcvYMtJYf15zC
GOnYgEDaMkQfLvQyfb9O1B2nl6NGDEY5Mi01nlCSuOIqgN+nOsSCdF6kns4ssAOE
mefISEcrnP35S5Kq5JrN0KmJLxIsYe7WjuDSYHJA08QfyQ6928Goxib+GM+nNWsS
ORu8POxQT46ppZVnI9YJ3mzPjwFvIAt+gOlVzgSkWb1/rl3SwOh04IBCgJiF8vkE
5HwJ/GerpgOpBv7pEvrasoIb9B6ZpMfUdxj61OeXzjBwA+tvWZDVAUB4FyawhiUW
NDoqtLIS9AnWWKuTpaOEI2VWC+lZe7Ck9BZtzAI5kTyI5Jq4LoXem3JvrwMlCg3a
i7zWDgrgT7a+FU51Qd/R4H45KCkcVR/Vpt9sPZW4eWGIVsWz5Q1wrL6JGeVD13lD
Lw+lEd2/5lZznvmjYGOW1rXMFZfPmSijlPDT+nK4G6XJSWGUsTPGvhf5O+6ZhVGa
53J8PKqbbpcKlx9/TFfZAWRzq3YncSSsg52UHt7NsW8Mp6NeMeE7PjpkTM1PvY5o
0f/Up5eCHtSqjyCyktIuxIYMHs56Z0ucogjhLkqRdC0Kurmz8tPE6pAo0Sf5dNFA
S+RIKmA8O76TOFYmbAPYFI7P1FzcMtZymNbuIR0Kqv49xCYP1PGWcTAUBAUa747T
4qSkqH4Wp/RJOLrOEVJL2jBO8u32z+6cL9RxpH9klTpb+I2XEfn18KWVf+GQfN4N
6HuOsrDgpg7fdQ2VkHKlTdcKUwHU0Foup6vmwbw5XBzXotaUrTcezfgLkcrDFADU
PRkg3xf6zRXV0Ycycpa78sjE8XKBkMlFlxhB/yA44g/VJBkgDFc7gteYYx6U0nQL
jnV5BpALB7lK517wlbei05sIz1rQXjmEAYxyks9JRQV+dDnDAn+ubngseoiNZwbE
II3sUtyeALkGTWgvmkAfwRBH/bktUK9F1Kss/5VAAdHn13ZNjuuTaVRVmRCvQLdB
FlfU92KuF/ssW6dFjDUFarCu3VMyhz83j+PtwBy6AQ3n9frgf1RUEX8OAuHHbn16
R86trT+uNhj6SBpAWH2eHJBToV+Xbw7GOZ+V110nUACfuNV33k5BquKjBk+A0Osl
d9SF3kzOQSFDezOh05JiLrDWJunFloAfTtzhgh9uyVj2+5ZERwBXbKiJPnjXTRMa
ccFWWtzldhsEf/L3KmZ8Pm3vmrxbFV2esM98L1ckA62/20+wqoWhgmH4/1D5/FYP
ADWKWGk3Z/D0k3wvUpfutbJD0PR6SJP2EtPXpkq8BTNNQRCO7UrwFPBt0v/mZiHW
mmFEDASGvORlLgLrKkAuq5Go+791akfXIiLyI1LXf7xFhlxi+w2E3FBy1AXrMT2z
Ur/uae9d5S3rKEED7Nxdi59B3URTMz9zOZU6YksZyXuoWTe4xZik59ubXB/mJv14
hETv0aQqd/Gh+HGeu9M+TZzxE6AQiVtL5W74kwQ0aoy3FKytnhTYE7mYUzw10sRF
Qs/UQGJlyJEZBHIkKmLgJR7O72dxoMfD+MM4RQfhEBLsLJa35lwHDVT65jBvwFsn
51sbFaKxwlOb4LhFU0ZWDu+dyB+RUWPH9dgFqI4c26ousT0Yj7ZcPg+RjSus4ZVs
IcY4hT2CaPZhzHuGVVrbRhlUmcFrk1k9fa7h/HQtaUt3SdB5WxTbfhmscMrbO+s4
maG9pLKeYDhGfrS03jl6U/fDjb/Qj+IdKf7ld1ZpGT3xkDiXhsSPis+j2dRJcKzY
WFE+pqiLnb4jDMDN59OaosoeMca/IDG8FGhI3RlMfgZJ+CauBh9ALtxQZBQN2uO1
rCM5wK0836ssYQvfIX6Eugc5PwmA7/yt1sPWoVAQooFyCtLyKkTBPwMxadrVEYE7
Z+iBhnjWmOXY0XakQyL2UWYNYM/bcYtcHHalEI85asjCC9jrTdVyJoUilr07HrbA
JzQj0rChJC0pJhE8RMt79jjDQ9dNgx7P3MxzAtdYk1RnvA8JMU30UQDGaVyMAtiW
pXsnIc1bjL9Ei5IChXCFDBSsEKD0L0lnPOXr8z9HOM4eZAr44Wuq0Lmt+K8OSUmk
B1tAZvK1ElndfZntSKx1qAPfrYAprAbMfLlNT/vMqIjEU98we9UE9wyO4iwbedSB
Fd2LU8rR0ivp+Kgwx6CEC5AySZk5OVC6Eu1fdtv62UPTp8jCtmiUZg8PEJfAj/gQ
Lbx+R2UDN8a/qKzDmkA/j/oK3UW5IXzS0ipHvmrgKTDR3PuT2u77q8URElGkXdC4
CxmKCgFbHHp7Us3Tz43IKL4WkXG4VDXa5E+FUtwzEAoPRdmQkTkR6xOP5aqXMDSx
PWsm64fxQUScvgSVQVeMxREIpWDxQlQNV2dpQo0oMM8qmYymBMYD1WIFmV9GoJy0
FgnkPdrgiA2BdgBhrhHCF/DBbx+DEaUZ5mqSImqISMyPs6/WrWShA3vvl84ce83x
LWVjL2H8XK9CQqCQDHfMyw+QJ1P2j8Do+36pnlcE0wgsJHbL324uh8ooW0R+2ufV
Q/4gzdjGp37M+LAfWBqBd8pCOrPUgrtarEoq6gbn16ac8oNzyxnuzSmkUgZB+70L
tVwx+fdwAyN0WZSTWLCdPzICJXdj8fs5Sy3lueKqM2rDEKdN47zxe4rxnz8jiGJP
VuGVy6Ckn0wAYs7SlebBWY26eM/0+kgX4SuyRsCawP/aDT5dsuTaR1VjRjqq84kM
x5ohc9iN08IgUoubdpy1nOQ1uY88BhvPDjga9JCMfYrh74yVBnEycNkFPOQPeKEs
54ACidVdyKEeakIkyC5pKtovvUgBCd7ggRkki3DANtbPOelI2+a9Vwp6tkDOxFgl
ug3m5+G6RRHiu4fTansS9VTJSISnofC4aFrOypjb8ysKjbanBWK15gtDfWap9pC2
eX6ovmJ38dzowyZKMy34cYIU0Qm0vf5pA4Q+7CW75YvVxI+n0OWJBRFbJ4u6pUuG
w/eFzPkgiSjBpzz192wkv1k73fgvX3QIP8U7kCAlSbBYkGLt1VIGxK9DgKiZd//b
wSyJAaBXt73m28bLsjZ2IJOYT4AA/JkGvNICH6q5z8/3lSiSZ6jCRXDfHOTOA63H
jH0n8Awi787ajCFmA9rMVf3KxM+iMsr+c/jAuEpZCZQVms8qafjPxUQxzC/yFwft
UaP516FXjbhyrWi+ocFxo/zARO5NP4xE5OEJa5r3Cx+2faC6xmfDeR0e1D5irFyu
6yd3oVH9PpeKZTxyMbwhKPVSrl9DyusCfg0xdNwpL1w1+VMgEQ5cUm9R3z2Y4qav
dZwoBXJn770ksQwUqTg7+C27UdtSPLwQjpuGeGmZGdNv9iQwPFqMgmzWUNqJUFRy
puqWAvqdG0yqHiVSSUjee8saB0vxNXMCWlZeuAjdCBhQvcYp5sM6Dzyrh62xWzFN
ujR/WdwRlZt4pGym6hug/ukmA0QAMu/yrenU5Lrzwsyc5nZwYjIGXMxNXvcKKkTe
q0ZEOID45XdV15vqUO56PfbA8mHvYXe+Ry9ECsaPIHxiyR5hXJRvP7wJbG3bPzb9
jsdyVJBNZLDSGH8WQFub7V7qdsXxkNN5ik6b8x6MFyubpb7005vCp4CezsmslNpg
aXC8m+10llsoCHxQuITMFGmPSJvJy7wswTZZ8EN7ZLo6osKIs6Cv2fRzY3EJTQsw
9TKDlBC7ygo+Hhck99CGCHhYrctCFQnrs1g8izQ0dbcTZCRmDK1L0/xWRgGHqmYn
v3+diK9LznygJ6nOC3vSKBgHdeBtxCR/1da+YghaOf9gC+QmL+aVODwX2sutu9nT
jmNU/n1V1GwLJzCq+CYss1opgJXc6+8Sl8++28IdO35tpRAMSuT5cmtXE/m3oDQZ
gUH2sRQh+UH+YiJWu8k5M5a3dxcdeGOyF8y/8mVwNRJOszT49ROUnGasN1Hj+jBD
Mu+eUcnaHhKlWqClrljD7eeNQlOl/jkGqJWntNbgl4Udbt3jVhOgYwzipFPsXg3j
z21gpoWqGlrGLQgDGHRJrZOwat6bq1NcJ3Hf0ZnPUz2yQ5WiO5a78ishKYld6GKH
J7j3HhIZmvNfR2+yu6Lrc6+/W6Q03fy+HlJzlolh0OQnNaMb30ET2pOtN93jGfe/
dBtLUdBAnGykctCqAfrBaxtjNAUJPkTUKO1MnpYXM1YU4ajsfgkZRCz4hcD+0t5P
+dezN2N/vI2NsppZuDeirA4SLixFFQuJy6vGC6SRxhDp/UznRp1bSfpXQRKbZt2Z
Ed2Zvjt6JXBMzQfmVgux6FfE4tzUB1ydjD9fBlIH7UNMcA75SumlVdUicaiXOQ+w
U1NRpDQRzmE1/zCwfOwTWcZb1frFF/tVLOWCpw5WANu/czRGOOBjmvszAwaeBpa4
xtsnOElUE3xBXU1TrJrTaZnFZmlpbB4dhFCvyAx/3Sw1kH4ot1sO5MGqUdJRhWfy
/gXpMbKXxY195TVSewyl/mUCFOGHlYgNOvyHRKZ2S/Fa+RDDtYkC7rPTD1YMR8w3
3tjkSysuZDgZ0cZyiZMIwOhWsNLiMUdlElGUBXrRSD409Sc2kKzbesAxI1KZNQLo
OazN3itLPKCVI9ykkJx/XxrdH8TMdNz3UJ95C6SG8DARcqAMEzW9fVWsiJvDxw28
hlbDWokPtoxSswFToVwtlsZCVF/2ag+pUtTjdTneNR3YPiOwGxdRNp6UIf1+iVdp
Hb298GF8qorxdx4hxjBuegtYqnF8vTZ+V5GHj5Fl82p1vXE3wZSG/bI0JOGldexE
RZS7dsD8Ud69WHfqqyWC8Kl8mSQwfvuCPiH0R0KuEcjImBcoji6H2PhyggymqqAN
v6wP3PC++8n5p5LEuvJQ2hp9t8VpelAracwqWBFWCBdhxhZj5kvw191BQx9msKwq
Ix9rsU2E7RzfwHn2Lzo51bKzL/b9XcdADAJ+c2AaDwoGw3/mohNT5G5uB992Jr9S
/Pewg7SeAdo8cbqkR1FBOif5W8sc8uw1Qnyn3MTqypTMvZn6Gdz+Eb6zvAjTwFj0
+Cia5vm6wYyYR1McW9nu9+nBpJYpqQnWlYyJZJh7VPnBB+UgMIQpo3STTjiA48P9
nWLKHY5aj8J3L6ekXfCRI81yhn2tSJgngR2i1hBHJiiJVQKdHAiUmLNa68p0CRm4
ZzW9hb6IlvuKNae82PDCHzGwAgl0ZEBUu0Uv7Esk1Rn+g0yqEOx6HxGgq1srlmY8
j0FGQWyLFkkTo+LTYAGekMKid90xaKFUHE7klqzrq37RyVKRxOX1H2HA03AI6ZG5
7bU+tFd2BChBW10vmaWA5RU7b665fAI+SnXJZqc0AJK3F3hm3sPn9RgaIwkL0Vkz
Tn/EcTeX7TwEIjhYtt/Dzynk2ivS/k5iV5lpFeBU1AvMav17qRwuKWCqWX7dpMs2
gz44AagVSTfkdCHikd/AVsD14Lf/i3AiQ7t7PWdmWGfM5rujBHRH4PWh454P0j8g
IWZYqJUx4pItplbHEqHRRFZ+yQViF5yEcP4IXf5Vph2d7572tey517SnRu0aj0Js
Zy4FyqS3x/n/O1K8bbnzqh4EJvNpX+zfl2KGoIZtr1zsiVLQaa4U7Wk4hdGHGt2+
7ITjJ3sbnBgCFbkkKpnKAhzrC0SH/H3e4DH6AGX9wKLBcGQdvbfnQZLIDD4rNhjh
4nTMAW7m0vK0YOaSAtzZnVJWCEt1vxe6v0TBn+bwj+3783LI5xQgLVv5uzqciVId
PLRrosbSPd1hredrSAS4H9s4tNbkTcWEd0DxgkXi3nrNan04pGJWPniwklxPWrcU
cDKf1C7FyiVafi6EvIThqFN2LkjzImtW+hwCXEIcqCs2XHXvVKEvl1/L4haGpB8r
hln9R9CKNCUCTfnMgr1t5AieEw5nDBE/lDwXtHU+zi5DPi6owunaR/6xH81oOTg4
9AR7V2JjAkCUHJgwG0kU5pR0Lf6wlOjPEoZrdptmx4duYVLcfUJXM5yEocUoJIcL
YF9Q/LSa7rnTbV59/hdxGmt9Xsbo/tJJFZ11BsvPNROG7ujfuGVH8ratnm5C7FCu
/os5sCChcOXxM6XM08/ox/F5ghlpEIJyAcPaXQ+0MAtV2qdw7u0ZcKWRYcqdsTOP
3n/Hv1T7KcPB4Eai2g/oTWKPfOZphP3QtbiJVNkaFqnBvFY9FD+dIf/O1Ncuc+Uo
zFR2rdI0uKDdqMK508gOQsqfJXp6aVI6CuYgfgAZ2mOfiiBrU6V3imgKxKQ1qge0
bibnjPmR8nGdNkKbYKAVOhBZ/GVekQDoZ5AkDHkwxcxXpvPS2itDo7l3t5beLVnb
cSC1tHqKYyqM9M7kdpOMHF6AKTqqk3zXcK/nxybx4BeF7uA5GNxXZxqSL16aTxrM
gymEy3kDqy/iEFYB82354lkknRtMli1S9oJhU7gbxU7Ra8Rf6IzdZNJquQlgjFz/
wl2y1TEYB+KYbMCxYSJAs2CtoK0nSBM2x3um2r6R3IMFW+BjpaXi/iZYxtbDe8bv
U5TY1fL+dMZPYV3x98SiEdDDxdtl1A8iH2hdrtDHsrXUpdjP+XUaKvFxkyfXmRvS
7UkwxrmaDxVjDPkO9lLRgQyy5UmFtpysm51Rtjt/m+ybBVnnu9ez0mbbfKWLmHjG
Xndfxl+Pa1mByxOXFeVaKfCJZbCEXA2bZqW/pS4CSOdQEbGGPvOgnHYtUj3w7aEh
OxqzUtvsGFO1WM817UZiaBPMxJT8xyy7sB9fCEdY+Ew7uogFXFn0b5TVwBz+A/1s
s0aS5mfbko6I/GqurtK04QvL62GouXcnxNonBPWNl8Cz/aw74XfT4fBmu6AABhiq
z1UfUjAjzpGVDvExaxVIb9gluC4QEspnVTBRe7s0VgVRUKJewnm5HveepYuhjy76
T7lDeC5+q54JzKhnaL+/ZIpEpLQ3GqkpBL/aDFkMy26EfaxwrVJOsPzwooAtyRUF
ADUkuLaGEJAYzbzKjgi6/ovV6aj8obGwCYS8WifZCrbO3+vRUckVO5e4YixDUEte
nCA2NNB4/qrsD8lJX/BhCsU73TMDWKyiZN46PQ6E7aGf3yDcg2Uz3AEQpl4sre+b
J9i83+bSNlg4hjR2yyHAk1cSgZQCswsOjTzwBKtmuCStzLy3jf0SeVxbjKj7rCK/
iaqz6lg6zkVPkcFIFAZngNBxRVBsR+apPLm/hd5w6VtoOLl9jWsV9S8pFDu+KRJM
O03AI56TartxE8EgQOQeaUp+kpz5EcebegW+1Rw8ianTSU1Z+DDZFbnhklNV6P3H
nlL9H0BbbCLcQT4rhtJPI0IQ8584gfuG5JnCCLi1UeW6c5cXc/kW0SZ4B/r85YeM
W9UvWrNwTmALDeh2K0gu+KIP2SYJXnP+RI6+1wdWwXJahaJ5n39UbUuLTgXI7/Hd
iqkaGxys0yZGwgO91eSEZIOwzsFK9TQj0mOACGLnThq/PsItcgDevV0aGnKZ14MW
ILN4LFGDORWEOsgbBYp0DuMWCkjKlTgxKipbyGuBH/HbdRKUHN1NuPRKyq7M75hN
3/h6xiiodSDkV4mXs8oUQdPYCU04hZN72TktEygHaRhUuqz42T3kPtoxpSScpdRb
HLRRC5pDytQ2W1Ydksd28UYKJhvoa9Jq5AysAQ/unb2Umu19LwVyeAEBW8WZhFbk
lWPpas+CrvlDdVr39g/N5PUc7Oo8gKRpXbTdYZE6lZwuP0QjXKUUUNX/ayijkh7W
nbqXWFniQrVWDVw6fUfPNKnL/ITbzN5q5OOv3qMUV4uJJXUSl1DemFTGTQYlNdmA
woGUQ1wQTEiBHBU6Ee974ZsymedmUjH/yWs2rdoCqAPiPWvw5EMgADy3CGxNV0i7
DfmDpIZPeiHe2vzfUagwEelW+8BlzV0pjdVuwm08XrzTUYMZJFZ3NkGHDeQePmFY
r1Bvu2BwRXScyW9Kx1wHw+OlyAh6u1GWaMJzcqDoHDLAwiI0fdHM+ny8WKtW2uda
OHGDhYBghn29qAhYSFCVpNPqrSTbxmS98qR2Shm2E59qe8ZgMFQ58sK+x6OKjCpO
l/UiMigyZ6l5hVkj65wxKL34GwkCKSF1krVAbPza2szGgqC7y0BvT3NTsUq/TCAP
OAvJXosPSMBb0d8oIxYv7XEFkEFtAHUMiaqZAaeovCt7dEKfrZ2YFMtux4fnTR5Q
0IkyCpXtfVGOG8vS0t1Zf4KqrBf25/H1DPuX/hEKhm4tLp2ieUXhD0jlBuCE95qf
/9JWX2PitgZ9XIeaaW1Qn8EmHwLqXhE6TykwM0QNYemY/Ls0MyJu+yfSsUFadhS1
jRKUGXv6QRyUINcaTijJ7b4HWb6M0gn8fqSr4tdOZ00EacIPPTMsZedm+ES3zOQS
fEaLyWGuasUOZW/ZyQFTkGHz2sZNLJTDUY56339fYB1oT9vWnvrPqQhOMBX+2clc
HbIsByA3FvLSNGb7nLA2VV718/bXxOJ9CLHaGLZ5JtyjUNreYVVPrupm5Fw0aODq
RzyU/KnTXy5LXKDHI1zfjqwoewtBRFa47d+wIxhvYETWeyVXX0/eRNxEr/Zy4jN2
qEK7v0CkIwc2ApXlMEJwwJLac9+nWNxgRv8jNZqUbX6pbccEhnJio7eOD0NjJ8iT
R8HJDwYRWDR3SIhf9vwimrbruXzJgTFGdn9N2STyT8Hi5/UJGYzh4ONQ5j1gxIxD
8elXviPXoH0ACFUHzBudltDZvl2j8xzDw6wmIfzGD24bVQbJpLsh5mwYPqIOMy/c
ZqnvpYD/P8b429LjyuRuDGUwCw2+MewEXV3XoR6Ic+4pkPHKhUi7Bpb0LwLPgxEm
Py0cTTgdhdNhPUQE8kcVBXzay19lBUNexz9RzS18WR15udsx3zzQZ0yGb0ioGLZE
ZnOEQQXy4Alt1py7WYEY1pkXq4Pv1USsiHnMV4ClTtaZyCZZuXakBw0rh0NDmUKu
cDU6PuDkW7LeUZ0WmIP1Wrg4ss+jZF9afEBBjyjFc5r4PBAz2rtshd02N+dAdrFZ
r9ObTzzce7EVPhFqdpEjq8r/ISw/UX4NbowYEvC+5enyM/lMRg+cRAqf4HAWf9So
9Yd3I6NxlC7bhofmFAUueoEFD5wVdJZxEglouFDkdyAPOGpvw/H+1FqpXkcjwzdO
H/inpJ1ct7hiLunqeTU5L3aHkUXibgtHkrQEYuRtlhXieOk3osOfE/On+d4QpQ93
SGHs7JQcu7ZfA+xWcQJhpVbpVUFFkXDCa9E+VOszmdeb+jKW7Bl9oqRES9BwkiM7
otcwMTcQn0HhW3hXjNsFqzksp8aA5FqSXqOURCUqHmxUZEqoNjcIJghOLuejtQgY
/1/x5MAZ54EOcsuVJTxxrwHjk9QgAhJ0re9QW8B6PRIv3VpMN2G7obh+IHoXC/DY
hyewnPipG+u6u3Jl6Zzms10dWtG/aMUzLonVtl59irCf0rqXrvBZQoZsh4mnz3RE
mvQ7dRlbpgpOzPo3VkV0Pvhgu5cqmaADbxeo5SII1mljROJEsouyodhdpgiGLfby
oNwDT/CnxBqvUcEs3pulCi3NzczFWUA9ckkrA+35RQRTO9hpnlemhLuU8Z1cH7Xc
2AzplGauJfzNmdhK9BXctk9ErpYhn9mDYZbygR/EWIvGHbj63qOG8sUQ3nPJqjtf
eKRL9Erl0Bj2XDNscXY6XjjGtS4ISEtxmVMsPCpp87cVC3mQtHT1+U8ghmJ3Fe7E
HIegmtLhHKq4fbFagoUQ4pEFPMtoDv/qEZWnw3lzsfXityc/Wvt37698NUj6O4Ny
SFyZ8/YvgIzDCIG1ynBLjzbO2K4HZE3/Sf/CiX41ZNTpSuPfQnSijEV6okaJkMrC
Ddnjv8D+DxWa2DyR9TfvPlXlYvsRkBatH/m1jbsg22tUvZoIYHOBKeP/FibW/hmP
1GtoPb/oVYrUOY8MD+D4//BE7tUOQDWFAxed76TpY5N0lVu3cf20J7h2gy33Kc+4
rW4SiA2n1fCLL+sCKqlqWNqRFd1wBTFSkJlqT61LNEpAgps3q9oV3glNlgW6GEFY
24AaKpP8NjQsGxEcqqMpNBkipOmJ48qP2BO5ZvBes1uDiL51BhPEIl4v1okkWMhS
bOHxYIEtJf667eAI67QyGAbvjpPrd3yjOrXKiTWfBLm8hVHBuT8h9cAZVfC2jpRU
X3kLghHKU7vW/yIh64BOL6GqTI+r5DRgx8VFmWtMepmpQdbmgOJYcAKqDa3TVgbJ
62yJazOzRkkGdF+auJq/yv6+NsGSqrdaPWxwXzAFonjeYLH6c6GRlibYoJft1kaX
NJy+oHLfz4HQOKrvzZv1hcVSQh77bEkf9kjOdfcHNBHeVnP+qwg/KMHetcm3ddJk
JFN8DWdue/4GIib9z7K/+O9ZKj0iECAAVWL0s4twGmePaJuTTCzQp9amc3vhSzJZ
rwPt5114xWHV/Nel53HH/XLI+sn/LuODNa5dqHo7Gu4wABgcJRFA9BgG6xcmDgzn
ma7PhymGqZPgJnaRzwicq7B/gldCIn+7+GzEogj03fnjZuL5Hcg1Jd8Wt0svMtnl
ekgMK2QXKMVr2rTDQsFveE0q+jaxIVY9Jj6My83Unqh6PgcExvnJGfOduBu5As62
zad0/xgFEInxhGyTDZxiKDT7LyCl4cxSqMvqfNjL9QfFk7TML0Eo+Nlk8A+1VWWX
sxzU9XLMq7wKmCW3bIe5miX+6zYueGHpOqidzo3cs49oQOX39BrvOgSjEaRkv2/b
1XjytRHWfXK6IREJFD+KPsOqsqApS2XUnRSH00RqP9OPVbdkdyEwnwB3hFQnNYVe
CLPeinop1qad+G3OzBXZubb5O5K0hrgfk/suvfoWYqsqjhMKud9YL3P2FiR5j12p
8SuiNk4PEQw/LdiM9Tu0jPSAwLko2r9lOUnkGZeFAWp7mQAczcLbReOIUA1m0Ram
YevKOOND+a8XIdqZOpwwpwBkeTBQZDeAUivb5V3Lw8CFp9qykowT5ok0SHiFd7Ws
FKfYoEesY5uL5tmi4mdnVsGX/OYVFo4Qmk6HPrJPadVlH9rWiYOxa0koREBsHkK4
7F34FNGgM7BQIrSLWQtljYB9DKk6AOg24pTvJXgukKbbNA30Q4eqlrIuwYASxCAA
9ZA1pehP9YojdbKysgVAiyBBlD61om57z7goQo6Ma5TCHOKAlVdMNMPHPmqL2rKa
oM7cqZ68gzm2lUTPBSDqlNeaH1l1LgSV129zfOcqxkFFWvhB8aYOqPBQn7Ny+uNd
EuFNldvLhIPwoaqPebcsrdX4ol43Filye9KU7OiPINtY9EFCthkPKt4S75zHoNJ9
jBSwVcVTYNE8JJ+istX1SMDpZypidXuDJ2F9SGQAymb5pvB5T2mfBrn8DXLLJL5D
ho2m+veZcxqjfs/M39yftQQ8isMkm8n+eLw+b21xGg9zzbW9qbTVeEmlvB3YGoV/
N1JsPcid8R3BmqEIVcXBNWA1Atx5xc+I+Lq/bc87YCivihRD7ZwZsdVhf9lFiV1a
QvK29e1v5yyfcQQiz3kzjhrQHmDRSfdcJjJPAfp03fnfX8pn5VkWmze+HgLSxHZh
JtrbaFLSAyRJbYZpP5nF1P+9PYlh+GD/3IdsIYtbTnQYzpypNlNiL7C+ThRMtdv1
nv4gQ1XmuVn+kizbkgMAV6AqXlV4xwb0C5WOtUSY564Ypx7YhaRZyvVGwkMgSD3a
u518rqkG6yNEetmaa3e5lNV+oPiCKQTLI54F5iodMhakHrN2tNEyRqh1rD/4EZuu
+JSPmFqGYhJMHTBjKPof3kmcRoOuyjf0RZmOzDcfWj4kL5AiUYdcAmddF5GuQnNF
albyhg8KIBlRo0JuEz4oTv3eG0tY2QEmjYAiBsURHjsrtAUfBgpBPb9bJ5hkH17Y
i7Q2hLZq6nGPtRkq1BgD8rb3W8wxT/EEEtW0DjhBXihiTkmsrRclPSkLeedXWkBR
2td14u33RGOAvag9wSXvyBec9+gxmEai6esDTxEK7D/t9i1WFjVemFNiPJs4TFAR
tDM1p7zm5trlYAvDWCV0kNCifJijJJY4iydEjXCIfguDlyUl2/1Hb8GQkF6GMxm8
olgZllzr+4yhWnfxIyPg6/JMe9Ec9iJUkWDfHvQsvWiPfUCB1y/R4T3Qn9BshyUK
Na6sv98kBFV1IUfUgYk0Kh5ycYUmZTYjWFGljoVOAbS6DGTv1WnRJwxPp2LtIM02
DiFhCLF9Q6SM1mls2Wowrsrt5n6lPl1Xx84kb3mYrQlqyuHDRjTyAZCz4LmasUXS
zFLM8shuqMFI7QK3THvNld6dGfUJ9LfvK6cbLGdaH05vJBRttpwWkoFIAvLY1xjn
BlBM10eS7N3rXrnpzeThqeGMkdRn6x/seJpoGFkLevgBwSuDNvO8+ttBpKLipvTF
xmepVcpatLN+tgcvt3p3csX/zUs+ppAxE4cAk+pWiBIUTN0EHM/VtvJ8hsBuEbR+
H59DOk3OVccRMnXsBx/9gbsLet2iiT2FYMdMmA64KV2xrHvMKABiLZzTfyofz7gL
W9geYNdyIoK0rbz2Vilb7KE9UkMjZJaiByOT1m2aWSZu1HO75hCHLLtQNtd6O0BF
UrzD0rfTHXnX/oPche6LITpgx1vA3NZOOK2uTwosm+1aoSK1p8bMBti+I6iywYpg
p/6ZUYa1vnbdfctHLncDsXE+hABa4FEg6yWgRzGmmQiAP+stFaD4qFcUxIL/YzEW
Eu9JrQAKOaVFgi/MKcz/lspgmWsvK1Yy1U6uYpb1RG4AylHPMtyz/0kBtxRYaxfG
YLerdD9bPhG9Ofy3Vpz6GrsUkFtFjtFIAxpNvesR4ln8EZLk3In+gHLjphX3Z7jA
RreiQbxOJicW/nPLkl7BoCnASC+sfF1ZGM+YJ2GQFmCco9d+w6my8u60aGzQ1s7g
B2ZD+yRmaVFs+VNkGATtP1llq7AdXSV/9/oFFDG0H+IBEWqr72tX0flK9Yn8gthF
xKthIHuG0otXmahgxlKhaMDD6FEX47lhWBWRZ4FDnPTQZB0fVHwYpacSjR5eOOXs
eNc7SXvvCVrzWiX3CfKcP4C1WljA668z6pvQoWzyF2KNyGRibM9zPudW4Fr+z7+e
myWN69tiG9og0PRIeHd9QdLE0H+fNR8I6zzDkRV/2lmSOvMvTr6xp0qm+WqlI6s0
togCLhIRwM7ZLdpJF16JRyxWWfz6zMptmfUK5o1BeodwysFxLFiuCppmfeaBReMa
MFnZL41FAzGRXPJH0V8HrkpWoktUzeJNRo/yPR1ufSXiZKL1l9Wf6xwwbGTGVwR+
+XXVfzbmGp82tCDlZAEia5VBRuW51zmDO6dtLJTA41VG2voATk+fTf4v5/oiLa+q
u7wf2fO7lD/sEOyIS6z1HWIbyxuOKRIRIRhWGcUqn60NXwmBFbOXwPjhxKlEss+I
QkZzOlotW0PInj/Xhe7cDwCcuOjJ7H/Of26C/cXHisRWEOO8yk7p4soInxBcvWwp
uaJULfnqwHtjKABvt85pLLZloOTehRrSTn5bWqCN9UDaiDa3UkosPb7ZFOenidmG
63hTviW1I7KlJRotMOfpa/flyk6glJnM/zQzv4jB3jo8vsmPSEzop1gwy6cRZxF4
lacDX4tlURtAQnw8Bvl6GD4cJgqLBoV885rVgEVoTlBJHNOw4OyX+n94/NlNrD9f
xwSPFUstigFbnIBw78IFodTHZ/vHs0nXwo1+Kb67xCueJHJ+Um+sGebHJ4O/7Kk+
myf/n/rXJAxdS18Vn1IvWghLNTb/DgGigrTmUeLqdjT6tqEAgOuLaB+xUpZgWX3e
rn8+kr/KDKBP1p4ZAMvqhq/mai4XjV9bao3Q/Yx4alnmy4BHgcCqlJgIsNHsQOvh
3sVLEKg9bVgEwyoSeDSTyKsJb5yGe72p4evgjybstX3pByL6hvQpWlPmelVeKLLz
NtAi+DS5NIcRzdyB9jv3NiI56UM2R4uOHOooPqUnRoEEO8QzDVbZHCQmRH6K5fuQ
PccSvtB/Exf3vNZL4yPFjEI763+9djpVcidhwKnFP96hzF+X0wozzZ1DJcrZ+s12
oE4DJ6gTpBwRbiueS7knR5eWrUwSWtMS3lGG78viP2W1T4CC/hQdbKrvY/sD7VoU
gfP99jhFOOXVNIg9G1qc71giqxWYxkcS8+nySru3bf+r3SA/sF/u30nRftMbjsv6
Ig/hgGsFChe7STJWTBZE0mSrCG1rUHVILH6I8VUHmm5x3SoAf8t2HVyIGe8hBYIq
gWeT78dr0twAUdLq4iVXhL9adsb6lVFNlSlsBMB5yeGixKcrp8xmow72LQjMDIzU
5gkpw/e3c3mqucUIJjO78T0FgDU7T6ypJtj8czHgESXC2Awj0NX3B2ISLMcVAqsR
FE6SSVpqqBPWKatJWllVDAiaY8YnooKOfmI3KMUny6/cOuXZXvjT46t1GO9p4Zk9
RbmtZ7eyftv7gUtPcWlYCU0EnmpwWD8BhMO4kjXrxz/gZrywiQ5cPEgKNbMAsmRE
itJHMFYdjsvWSl4COO6nUvYrdFzHgjuvJxj+Q1p9HQvJ4ONvc/ExIfshouQMYV20
M4FyF5R6VHJvvnEpo+lFkA5qx1L/0USGx7N/rmSBCE7sxoSskBX2mqu9y/LHwwqK
+0lL9BrSeSNGoLhK2ULddVc2XglaSDJ+7bam1mxQ6nlTCU5scLWFXx6TWrPsBOEr
i3+N2tMgbaJK4bZG9BhcmjklhqVaihHirOEVVoZH74+G3yeGgVbdR5uZK5bdA998
6HrkuazTgA05zRnKn7B9aao4xWUddNqoLa0mupNKlOjsfW61GkZiqmlJu2hcZkie
kzfkTr9cb7LqsJSSiU/LdJXUnBIZh8xOxuyba/aeaEWOstuNPyDd+ksaC0IeF/ht
0stcUmN5VmVCvmLhnGbCcui4qcuY0kmxkwoJ13YlebCU9Oyt5/oGbBq+H2+sD3yX
CyxkTdZP+ic9A/omg2DYMDw8W/aUCVR7eHbpIxsKUHazeJNxXx4rX4ne96Sz7CDT
ctvJjoPFNvziF35zyh1cuXWzfx/wdSaWpRBhZQ4yxW4K1u2Y/GpmaCrmXIMdAakd
ydPBJYPvucPLNCoz+69jNV3V6yHqtsoLz9HbvNxpxGsC2PpYGLsdeYMDrJLN+GZN
5CGwNP1FKNH6vtCW8B6YR7+eJ2FCQuQggiiHHirGUZ3KuiB5g9UUOSdGumB27fFv
5aJ49e+DCe6fQ8qR4wpJBDHonMpI6lTguNwFxzr1BjYwVnj0E0bfXTYVL5AVQVwP
7MVh4x5VJK53Sdh7IqKOjrZyxLhXx7ONJ7UKx/ewEtt0VjyrmtHZkpy1tdpVqj0P
Nk+9ceaUMi/EdzxlETD2LE7SuvfRjMqkHroxPBtiKKMBzLD6y5n3OXloEG6mSWbs
HlYIn5Bi3rv4y/1gFyBY9cTaS32EelEpGJxX1J5nu2p6NcAjMHx9RLLGGSp8/U7A
LI9nNIxj9joVxNjKKnaTNFfFjPFKHpFOKzJ4FrtuaitE2CyYSSVfiM9pQOToBU6i
YyjKrLJuLK//YaTXvDp7O0o5G0KADFckr5xoeqCtOxQ08nYff11ze1FbdioG02EI
OGI8jeIS0YU5gT2Tr5APBlKdFj+/fxFvRROYCSa8fv0a0PTWqcShP99x14nvsMy4
lZLRDTvzBdbjisnlGqZWqhv1qaFDcEagI3ZVJGexUSOBH33JrPw9HDLgWqtcejB0
1NyU92rovWWv/b90HWyA+pRdp2Il75i4Gmzw4Jnst3oDqWWVu7SXmXajjKTKwuHr
8gKkZzG2w5Apgk2rgAqEimAgcVXqOxMDjOHiokfsinK/bCzLibloql+Qn1Ssu7aZ
L/to8sBA/L7BYNsmDN7JNj/tvDgeXWmb8FG17TjPyINCAvD6NWpxm6fe3yKVxscK
tZx29b/k7CWHp4kCHhu3sGOBHpWzjuR/EAl99pNf/2pZJTX132Hd2X/VUbvyIA37
xFIHfX5xgAuaZ5QT353RIz7ACKuoPe7WpPuFi/Z9WZhNx72GbT8cs+QSOkl1t0SH
pmuG5GCW2D5AsIUYIVrajSrFmayDG9ARASjvlzrZS4wieWaHelurlX6Y8VGcF43U
lVSGJJ/UQYRfV3/lJSAt1gt8P0l8qNQfH0hVaUtfdZr64wC27oyet1XtKVzvgELb
UobSWl1bl8eClAeoJp/m6UU7kTlb7A/0YWq2YMSeiLgXSchB51TfCQKT2asFTrvK
hqxD9FpNBKtJqsN/CZzMZJ4XwJgjrVnqQtNZd/SOeFr0rofgWWxzhSTWMFzZrINF
SlPlyAOOrK3U7zAPtDlJn84v9S3LDhuNEoTTrZvgIva7ZUXRXxqCJ4SXnd4VVgDp
1Y55oLjOz8Rr83S2t/YMxoDN/5vxG6Aw4a/WGYsR9eN6v9yObrHikNmxqDEfVOZm
8/iGQma9jtFP36dVfPqp1uX/YjH2rm7ZFyPyFou87I/HSUNuNQ55wU2Y4uB/aT1C
+K8m1Uir7D2EaipDalbuA2NDJsyKo/eMuybPmxKNofQIay5GU/q8ArcNZCjgPIji
YjRTu12BS3mKxo7Gz4s/Akv3Cq6G2HTihFL3AEy2OD4TX2gZJ32IZP/pf8A2uZgX
8IDutU3NOXZwAtFkmNsRGwkOojyNuwVGNDJJa1FaOU8JkC7c0/Zm3FrOaki9Rqwk
afkBU5IQ9TR6U3P3zqPpTuWvnFTU0/Bh55iVCKcvQRkojQ5jIX3mIsaa91HQgx3L
iVDGjZ4GrvyF/wmF5W7CmzGX9i9onTgqo7i42GB+sxZXpMWrjVcnAv5BgUGsb9l0
ALO9ZeCoVtBJXyjhp+23jW9+4aVvFS2Jd1+s7pVitAyRGYlaBlHVdjiEr3he4ik8
ZeQfSWOGzHM8AyJWG3YQWhI6lt8wSp989e92SqoFefH+8+ZeODzMhKEcovqg8nn7
JfkL6i00Kaz3ISxiBeBtCi7XLrdsh0QCu+SWHiktDtyN+lawCf/OF++jNd3d7ctb
9WTgz4fFmLMMRQVC9Db4XqCQo9H7DWh0EIeR0Yj6sp3TX5ER4cmqzJUXFa+tqGxs
8e5bCbL2bWBKJoIvozHs0uiRiRt8gvYBDlrplkyfkryoSEZu/N/CWf/BICaq5FM1
NIRP8HrWQ+k856X4pxKq6xHUnyxs6R60HUsEzOmOQZmHcbhIkr6cSJiHtrG26svV
RehGdgopkFInY+Z0Dj98gY5rL6kg3CjECLuCZ4tmD/14WbW2SGqsh95z402644Y0
oW2zmc0ajlkxQ26TusewftdYImIOvqxyUr4XWE5rFQniZNu0jrtjWAXxyq8YnSb/
hjzFipHPYkwB7hFkOaHtwboSL+VyBpPShKp9iwYrHUgb1taJEN2s5jNhiMzFfCEg
73D3JbMfT3rPGBuM6J5y9k+bPDmhIppdOyejOSeEx3SCsyyqGcKHnkCAH/vqD2ST
HsyHotXP9IaMqyHWLwfPfdvvb8gtUPv1SMkVGSm008s4q8PQXJaenwvgeeUglfIF
00koUT4so6bQO8ow/VTXW0M96eb78Arx6xfxBM4TIspilih54D+8fntVZPZBXqRK
GlMDiqqMbRNkAkzItKltT44uYkfWJZMskx1mUbHH4WTIy0s7oi5Ka1hZevt/rm2n
VwpLwjGNvqKrUuLZOsOiOIAYpf8omsC/dfPVp1nQfyJbhYlXYt9SgDw/5qyFjzG0
2KHFxlWhdgLAJ/fySOS4fGeYhyp31mgGONj/Kc+apuPHUr3E3KNJnRE3O2RyJh6s
eocO9e0XB4NDR02QbKZJ87eot1TJw4nBTxVtWTyB2S/hyzgerxpN/I6wsNzzfPMm
ynI2cf0a+9HibiXdMK0/4uV+tryKpkd6JxGiw17kjz6DNm6OMJyjXEYHY8tPMqMo
vX3mvr6mKXA9mbql/gCE8ZG9vH0O3BKATSnJgqDe3EEuvXgZBqnGjI9sZ6uw+g0y
T5SMYC8GFOOzuRrTV8PYtRflq/wCaWgeB7R1kEf6ZszQoOwKg+/2VLADZMa3rrpm
GHMBtaiYj1sLGWAKc0EIq/TgrMigOj73r3CTW8LUsBLrVuxRyrhoQM/eYspjr45q
YoDCPGV/V2jlF4y4Kgb94lFyAvX7Y3hdyHYT0Tcq/v5NjuCC01rsYtoPjHSw7pRI
a0orAXyq/sHilMawI7IQO18RncD8EjHkUS/oA6ONaSRFQmw+BNbGYHm4JHalp7E2
dhZBTPYQxkxIrfaGvh37CCgGUf3rSn5Ff2IuLW8lH+TpaikZqHX9+RSeoNodpGBR
nMY4oOO0BPKDeS3y6nQkpyCO6OZAQifdGNgJ4qFRrZ+cW4lJxy5FD9b9G8peTAVl
nzYArMfC+QsAs95N0lLTkL6YjsvnQdYZaAxJuYkncVoktmKSm2EC9M9EUjg3yMUv
Wib4En1IRcWEquxWyfGa1GkhBfodkQMOGoyQp6wQtfy50BH2ZaXj/CEdazN1jNmC
JgkBSu6eRS8r/6BRpl0rbmrUb+3BwRx21tjjg9XojmB9kIzLv4JBXm3aOF2ru1qg
J1Sgrn9yrGN8Q7YWGTfzdpcsLncRwrPpzhBaysennxlNtQv2TWDfrPuzOhZ3Q0nl
`pragma protect end_protected
