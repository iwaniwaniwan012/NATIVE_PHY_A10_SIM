// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 01:23:58 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VeThdgF3sRnVdVnoPPdZv1RbCGL/uNQSD7DbcDe4lNJtSpPYPk1WLJjI2y+prEYi
7e92WWRh0al+i6n/eNqmo+AL7Um3gjZPuEoAeF944+bGtKsJuErWaeQlVEP51/ni
iuiiiuNk4sO1Xnczi7mdognCroAjzRBCCUFJu9Qoip8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2809888)
Aj6PkDie+X5BjYJ5Jl5DaQO5aG2cTRe7tbJyUQkJlXNW+YXY83JLigBF2zKpTtUw
GLswW1cGRDeJdVBf9fu+c5IWlaCl+qIqoGJUI7AEqtHewuSW++dwgdB+fl9T7Xfw
u25HInIBgh8o9UwJSXJTI/aaX0LXLLUZ/D/nUtNz+iJFhmtsskrA9ndGfGaAFO6s
gO1lc7ExJ9+xnOkKE8TFgTmjGcywlZvoXE0fBC68+x7MPCRlaxYu9rlb7e+0EOl9
SSnleQqZCsRrOzY+0pkkAbH2G3JR/iFMADF1yuaJHzs2anliab48XtuZEfOth7IX
CBoHFP2yhTxgq8Y5jn6SsCTsGIUuLoKYV2GkIz8tXqKN++ryNM7ckZSvm4z38FS3
aHtrqBz2QY+3rHA+CQl4nZicR8M80fNKKkEuiWEQEkE2pT0ZuBLZZthxMvZV9Gs3
dr9CzbBvf8V+O40huV25jCmgbUwf87aYYWnZwSq86nQXZNQDIpwn7f5eXgZ+da1P
aXAkpwVit3uKZwjvzLYtC4QlGYEJwH96/bmCLCWVEmZbLG9Kd25dkmCRWwvFI05w
utV62PCs2/i0zq2TaQzsDepFfacuRUekOIEpBDnp5WjIi7l5Wal6xiAW/BnLNof7
Qcj/K8fGbjWitQF/1b/Okrj0bad8Y3buADdn6UNSzUHAxcC0uJQyu6JgFwwbN4h2
JyqezT0uExk3CRlQZsS5WomXQFiWUEmMsdtIR0jciHpugOiMPs0hYC9elf+xcuGz
4RwmXESn3jljADxlo7I1xWfzgaAQX2OH7bKpVuNf9lbATiiEF6i8dBJpNoLgIm8C
DHeuYj1lem33F4kITZ+PpIHAi9PkKPYW1dRvmNoXFFyKLIMdp9jMalmIb16O16c6
UylbeqsgAGJd0AlRvjjsM6o796s9HkPDkX2+BpQK0zI2avegRTYOzh8C3tIq5tAa
2RTQehpBMp/KRCRO++IEyXkmRdzcU0LOL0Rx0lCNYK2cntJ5Iei7f/6rbUsW+N23
hF/81+G67K8gl59U0eMQnElvues+DGb77pnJrDVyhjfpmaMgewUKG/3pmYf7b0q+
A+XgQxkh8Tkl7Yz+FVvjR0Aeib5Z60mhT6qPyYPw56MK9RFmYDwHaflcAX/TF9Gq
JCEtDBFWqov3gs2oGRScbuX1LJHYuUiu9s+mcDkGdtbMN9PhDIKmxT4jqIuMxRNI
VxEA7EbR+znlvrolb11VfddWtr/fhsuQ1WKyvfgagucjN5Yrm6UZy6YStaebTCVY
p9S12Bhl77coCKOB4k8uS6Z7v0dzxfVFNwncwteaNAcGfQsu/Xof01hYUdDNSTGS
8C2yCeXYr18Nh78ARF20rhQZ3REGDTlAZvU7cInTVjzZVuHyoG2sPQ1kMHApfjpK
r2GDlaO/DiCqEdz2HcUwBuZnQBdam06JZ8NpHDgC9HXTugrvBW1iLbLvCduz5maK
uAcriaz8ijfyWYV9bnALaoBHohvFTGzrgC4qMsliIPx76Iza+XcDHwvnYCvmRv84
ZWhfKUFJAOLq2Z/W03yAO0M/1G784utKHjDWdEfx18bAYi/Cq/vWG73JX9JBncgJ
xcVxhW3+bv58fXJrBJ8JAW98csGDpYg1qQ9GacSJ3XToQqmCmRDdK7RFSGD0lZYj
an7dQZUnI3ZFeiLUhFzMyguRM9Yr/BLtg40e+QviBJGX2WvzM6w382bkEBpGA8Ee
GoyfNlbOO+i3FGqPm7/PNntspmf92vbIqRZmOFLtFul/xX6kHuMOLpNjOMq2MWHg
BKVwmkejgOfdjkFpRIuNa5nK6zUnr4GrFulcwSnEExxU8hVOY9B2UizsFBy8esr8
0f4bN8GFqUbHyZ8hzmUp1FIyqENyd5eaX0lV2HxtwRA0UxiEm3wa7gQvr60BgDBa
63yIWEgW3XJl3ZxMd/Y1vkKZe/WfWILR7YjTzj/OKZqJLRauquA2/+J4bhwlP9da
4ygnF34bnxyAuP9yv92/hvqb2rWFKbmYpAkQTcdQur7AeICEl8LpUeGiUd7DJbwy
ONf1b0ZnkOBPOcIuQ+FCFkyeuS6xdNTTLE60+J1H6k6BnUCPsqCDfCyeF4AQa78S
UFiHuNJYK5VOZwtX28H/KVNLcMkXSyo/L25cH8pzJJ2JgPHSzm5gLvQEvB96dBWC
PdWCAuzhz7ATUXObM08Nj+ICyMABGYWIEGqhya56SwmruB7DJCGtvJdfvrq84dE9
3SjD8qS2Pp6PMwD7X+BKseQJUQMhvMlqTYwl1NsSawBbJazewzi0sOkWcNG8nO3c
EAyfs8wKuBUyYlTQWfKxUfT1JuYJiV9Li80g4o09NQE5QCPX9nl9ehp1N8qKl1Nq
/WuNjQVSfaNSGi4DKccaJwuL+mjmbYcVQFsfFf/IPBl0SsoljGP+t7bZZZS+gvik
Vxn1UsM3t7Lgzx4eXbnYydu9I7MDLl8+sIixGeEZFNUIcqaP5eMyFoOUvb7UewI/
SuBnLkIZi4uDUx6NYd+R0ECmMp5QtOyU4dFwy0m60Qnt4+BLpGvyQbLdmJXHWsTg
pHunv+9CLCw9Djn5AXIA6sfjd+8BO05XPObvy38cFQsdVsR3fDRbZSCQPMt3gqqG
SI181kDdb6xrbVmb2tiy9XSB/SyRLPyKJHFlsORiFv1XLdN2uPtc/ftNHibN0cTW
D0XyzGSC7Ez3TPaARTgtEtcyk0aOjrfc4FYd6wicJMoaATH3/EctDqFhWEXqvtyJ
twR5OTVc5MHH+kNUIdq7UUlT9ecYFHHX60tbz9GNAnguYNL/oLrA6eO75/6BNcH4
5P1lrZKa36eDDaSRLdZCX7D3yqG3yYpXaz5GswdPlzp4WipEn35epSZH8Z+OWVIm
/m6Hf09Z4emvmebIlqgUAZxcjS9wKv21a9gRtf+z2oAIqZvAlpHi7WGlLtSkx5u/
CvpolNc7F319ZoYWkkqZyXuIP5i5S0IP3XLdtvMZPvbLP303KjdBHen9YIwHnELm
aeXoidgG2c43H2IuRHRsTGL7/m5q0cwnAD93gUb+4Pe+L0ylKAklvVqdp01kHJaT
XpLOojaLyV91+l1yATxP1ZN/ulGRQk1iej15+pIF+RgsjjIYNik6tQkZC5vKhAuu
gkiYaxXvtBlxTNPsMkL7tbVDBw4MsifBHyrTFOOArjimG05GXQNgRLBa90/3zIlw
TqTk80PAjKGqxz461caEBnLajOyvVwNpC0Edn0uqkt2HFr6tCrLztmnv/ORhVTun
dOg6K4Q8+lSBc+GUAPk6yJNgtvomQ2IYrujSAnQOnyhxYHUHPMXiiMNBvsYf6fay
odBwmF/4YaHmA43admWBoVkqFVx0P4NHQuZKtY/3pvyZhWwnCdaaNkHj/qIXG+gx
iH1KnJey4s9t8XkexIadngnuMjknSVmzLaHPHGLNaDYW7aGBoierd4OZ9bQ/u/AW
NRexHEz2hFuI8hR+RhGSzz/KA3LlRgw4jtTjLzLWcKr4TbDVL++PyHa+y1qImDvX
/OCcxowLms05MdNXLVuYM5ECj04ggEYseFv9daJjM/mn067M2r0LGmidhedkUkTi
KIB6k0V1zLh3qhK1ZqkFIj8cGArn6EbKrEcSgE3ugR9LLKtJ2krOsd9TbOySWnD6
eue7Yt6dDM+PNi00FMdJm9A/6BinMuagJuzrWduywOWZS0vJny2y0Vj1nOlFPoZK
vtuXpVHxicEqf9/xlahbSLPPkb70FVGN56qgg5EbZ1fCMtqPI/vLxNytYEAJtJ6l
qS2ij0tRdWoDKXffP1t9SZIND6sd8YdbsRPYkXfV/xSG6yvcDV5gF1ADRmCegmy1
Nm8fX+y/sjcDBAF6HKOcCF7xz9zj9NwuJ6I3rq9rC87fpa/+tcima96Y+wWcvVTW
ilJhXME+70UaVB8auujP+wh9+hIWH2mijKVqM+QnUff8UlMMv+CkwT9XhNM7Vg0h
phhn6C3ziumOCJExFAcQNnKufjjLd5SyO+TfmdcWfA9MSWU3hrGGwJIbpxf3R6Us
n20m9xH1Kq4reUtknmzsD1VrZa5K2XPniE6MQjl9VcvdOA2AgNwDm8YLUiZES6gk
ffD5vMh/8Cq/NPie1BnYUsmkpkgd8j1+6mK6tgjVtP+zKAl9pMSieMUZBAnk1i45
alSYhgT58BhkpIu5wSD44pVpF2F868oJHmyd1FyIvu7Ue4xp5MtiGNsq+TzQsGV0
BKy7bltKEU45nLUDS/J1rmYcqB2y8G5uhLqvqdh2uOixVEqnoInExZ3bTfG8H6+p
BfwgMe4QdfdI3KZbE99JL+cXOnF5BpDtfAwsGSlPu4sso0ydw70KMP5plfng7tmd
+1xM7qZ5YXdqgp43iicAzGlBY3FVJu01yWrzl75ZEvRQX1JOaEb+Fve/GadUPL+i
Gih9YVwLE2G+Aq1RLDnHvdNUEBmnzHFzlBkh01PNZX4dfPkdWQvT+I9NYWHXR10w
XfJhQtoxeR1+pdAnxg/e849BUUjI+oBnISwCAr3E6AheXQ7ectcUgP4TGO3fb4xm
ZLCpVIDXE3BpMndnzMZhu5xAqmYnheEhTiv/4eP5lh+Ym23UJDmsiVrFWgmtT4J/
fiJ2p0u+6nvEziIvUkFWxU69ZzLuZKrcILs+mIP5a62b5s5OazTG239YFX4LU/nW
xXD55B+p/gsWJ+LTQM6a5qItlppTPddbOVywlZt32iPhXm2lNMq5YvzCRRllKoM7
fXVXgTkdDXPW58sqbeaLZhP0Q17ioRPsmbzH+SHC/XTxmPTlFe05gHds3fC/eoCC
DMvel7p4fRa9A9Af3kJnDAmmjTe21gg2t6I0tc6h3diYOCaik5638v80PAf5a5JP
L0Vepc905s8/pQ2qkrMwWC1Yw2XL34x7m2X7XxWDcdJCVEnt54k9woNiior46Ziu
Om/UtMzwwbOBCk4IsYghUQVnxVeZSerCxyGgyWYo5hv7CXAntr5lxgXHV9Q//XJW
YxTccaD0ErnvtOr0sOP/S/GNzffXZ56FcH0vjK35bVXW+IgKUFC/lhPIPdDnI9NQ
aV3Jg4QQnKKjjOYtTULZyLlFuuDNRKDj/2T6lm9sgYRxaV3lEbISthIp468QvTGM
aLKFlPRunxfi9B7ZdiWHvbd6k2KIxgvSLA7ilwx0+02+Z56kv+o38N0I+DcAn8RF
si/Ur6Cl63ohKat4r5jtZIpgbiR7P8dB25l5sz7n73UIGA/brwMjrC2AEkUzjbRr
8lIgs9DjXzw921AAxasahZp7qy1uq8q56MjodT86GXbKe47COUcUbYWwaObC8e3B
SnRBdTaoeSRbP8ZrifgAygRVg8YR6lh1GyUOM6z36ycYikByzIHWxH0AM4gCs+MA
svTeniNEpbcgSyovsK0jvnXmqjbMOqrevjCaWT+C9QHgGXYyTXo/o7gZTnLi0tGd
3tUdeVM41kAcwvy5IAOcOXUTC3X72guCS1eqbOoiN7l5YmaoeqzmLH6QMJ/OPU/U
hLVrdK2UwEj1T+7vthHsYx8nzFC1SoYCNLo4YK1wWBXI+oCye4XMJihjtORCujZN
jOsBCbI8wHePqv2GNXFN5SAtH6P8MStArIx/56EXvrbSYCLoaGKPn2m3nOGEizT4
1R9CEeiY7RWtC4TCTEcq+UimeZcOctn/UPZ8EydBPJCXlEraHCQLayowKVmtzIjB
k3pnlTpMf86TqtZ/F0wZu5bUyGFOwNwLZgb7POSiq6iADuDAWhPIbdzSquxFkXeI
SIzWWM1Bq4DerYjQVheXLGOHyNvRf5NY34WRetyoEUSriWOM+HttIk2DuMcVBYos
To/LsHR7kPrI1v44/qdhzKshF1/rlhkVPswiSA91e2SXbLzfPVZVEWZ21ybqbQig
q9VchRmo4WHEx0EGkMHXUKVCPJ9/vpauDIQ8U+yhec6l3rj5dq/n7VAhKvf14iKI
M8rQsr++stqTpS3axRGYyUb3XuegrA9pml4RIOe8j0bdY9mBuE9UIgzTaFGIOAvi
O6OHDWh0d+SpO/gaL1ymXKyWhuu1V1TcaTHECjXu3m/qvFVfutbVpnQitEJ0H6Oo
HDrO0plu7vHtQWsAiBgyl8mN1apaJ/OqZLKkEflrgr2oaExWf6J/6K7ZJdyDoa3F
mUyZkcLa9s9LePFr5cLsLDFH0BobOgmSMIj28X8ZNiK4Uvywl6i0lQdphqaKxLa7
v6Qo4HjJlHjAKndTCb0FP6dV9Lvmdu1PzLuu5Y+ifcxYRT3K4doomDQBcTK1M6sy
oh9tT7eDPOB4rIB8I3kMu8zEkbqM+FERgWUhietkvjnHPmuRhjajtUHjNmjBoZvd
RpcMOhg87mZlcJXcz5FIzlFLcFaDXX0/a13/NJtNmDSy97e0hPjrkmZJgGQr4zUY
cdm2/wEO3YjgMlXjgGuLcEK0zeVMLe8seHsloi7n6THoEKbCySXYjKHa1Lur9sun
aZ0HVXHLm/K00fKHuxau6jmG2dUADt4eQczYDiTUaWlVob9whO85usv13NPtkAcb
zgWYzSKoLJFzEkzI+UqC0eznmfsr1xdAK+mMGAMWNLOVrzYXAH4hV9oUOy3pN2WI
Z4oWjivuYy0EK0MKfOGOywYMTLzm0UL/5+9KBKkoZgk5/eYPCfbgLngpGZWDpSmU
7TvO27BIjRvc2NXO+CooaNwMae2+fgm1jJPrutxoENJDbkIOto0Y47XrIVgVpoSm
KL71hZue1eJBSwT3OOXOax49eqIZQOfJcpX8EpFEwnVcBAiSFdcDSnwQ5tf+R+D0
OFjk/GUezyvSTekseKN8lsilbaXl83Ao/DBVnG3RbEDgLfP/AMnJYqw052uXDlgV
y25Bbc1X0SQOSdLCmK5CpcVzI2ceHrezS/kBwBxPKoZDiI7r1ok1nuDj39P/Hwoh
tf8Erw7ZZ+Ht0hCeMy6/y8fJHXDMnb0D4SeWXFP5tNYpHqtrLvk0DxNsYlzxXt3n
97e67glnwl/aW4VfSSBIke0qLOU9ygnH5C25hLenCF4cQTu6LdFa/Z9YHpRSlkr5
0v/SgtU4NnhMoB6NnJKVzdPrVEwAD/u/cZUqvgfFmRXWNyFgKjEzVzmIBe3pfh5S
PUelmKxxiI7HnFEYv/CB+UDgcoOU6XGsktCNS9uhNdbXqEcbJR1DTQNhsSkQB0Zl
ID7FkTWqHi8Qopev6phfBGWGclwVA2o3MHoPxia6iBEPEtpBQ5dQ5OeRSZtIeNfs
aUmXkxxZwdvmlF+We12qDnS6h/b0A6nzgsqK77njQcmRiASWIsIKY7WT2jlJMYFs
p3wl+C49ybHeB7zb5hZhm/Z7izQGsU4gwmbgwUiDX9Dwf9wAGqzCwWFQcU+zTe3x
t6Q8pFeKxqdcwM+RHMGfMYP/bib4DZW35fEQYfex2e5TXc7gfbTMxUjXeKB+ZGj0
sJbOXgYC/IIJ60fdkQkwk0QspT4v3vQaiM2s/8Kom5QYXq+uO2Zcel+gBn6/eAUO
8+qLMV4CoSk+3x5kUOrZFU1N/W8t4GfDVrmSd8rdts69EPkmnWTCoMUUxBuZgRRZ
tVQIMQ4y0IrOoMIuEjqGDDmNWW/XHjJgjyEsgzPlDJ/yf7mqso/MVtHJqJswFWaT
ysqTtB09rFXm7RlcpfXQgPpZFkXnZPHnhwyDrLK5AHFUMQITf8aslpV3e+FsKBVv
WlAj75CwqCBI9eMathIQu/X+DudwHsbfKvtGcZKKGakQey1d4eHquJDBihyOfIjt
kA4iYL9A8y+vJGVvPjr9IMKN+eqps6vjNQYuqSWywaGI0vXZyIydLNB/sCDt3TB9
yxFzVpPw7ck3yMlQ3O6CZ6LnSfwfvxcoNmYdzHX60mtB8teUhs+uWpGYBg6PSg9Q
xSbMAVZ4DoGWfCtUma24SXllMZaNYTscHaN6G+Kk0E3FRT/GRwttYsD8D5X9mqMs
ZwR9S0tEy/K4DD/37mvOtqo2f5o8FS9JnO7T4ldWXFlRWcecLz0f95TkRBEGwS37
ef0H2zkwJIatHb63UWH/Zg38KoWpXJVD2cZeNaEI/cFJHqo5oG2qZQxBSCLTDvKd
7cP6V9/vbkQe4pMXklte7Q52SHs9QV/jV0I85XAArha0WOstSETN2aiPYaBPZ3ia
ldNDRoIDvHos+EitmXbaYXZqpTQH9lDTFwkecCPOz7J7huyNYfamhDrvXQgrYMHC
/jK0I3wvLfASwM0YDEbbDID1IoWkx9/nzsjbqEJFZw3ATXvca98e8DWhEgEk750e
Ksi1omEIcdIOr5WARG484ZrkNEgBIboKUlhRjg3QSqyYuFFzmr5ETFGEosvdPnhl
0X8o37exrnQFQnyJpAIcm926SmWveUFylYQwTPGfqtJ9P/C0Por/l5haJ0gi3BEY
nHt++GS/Us06sUoeqm7GvvoZh2EAkTPoNBEW05BHswgPG1dI6mRWo99RiNaHplCA
RwtksE/FcNlc6jnPzHjs1R5ZeCkDbmWnrGPuQhiIEHwc/aaVuxcoyvYDZ7q1V4C2
BX8ZT7JU5D6v7hY3lBW73iBekBUC4jEGgusrDZzIJLBWaRMhFgdbEQEtjoBS/5A2
NwG1L9KVz7R9fcdaz7C4IcZSRJbo3CWEvIDvIg6OboAaoTcd4lh1feidtYiDk31K
n2LQkg2uzsQ1IpUX/PtrTs7v7BAPGX35m9FMVTcUUO9pSUzT+lfMO+NUzFP1w0AU
1ne9RiGk/TrncSq6n2kqwyzlVjr/qHnLfeoxL0vD53ckyb6bwOIrmAFRi35f28+M
qUkpOJySWMEi7XQCJl0E5rk01hr06hdmwwI4oMwASoDIheC7WRlV2LeEgGWJaxh3
TF5x0YC2bSbEcfZJV/3wcsIh0sEKgsNa2ITt45BQKN2lSDl1Ycz3YCdYhcxIYM86
wyxACKouZckWfvM64KuYYRdIHA78f5F4Ve6qygUDlDH8AQLy5yEX2m49i9fq2zcd
N6oTr8yJriW089QkN4A/zs2VKQMte0LNhitGSaJHV1iS7Pirzq3QPLnydtKp/jTX
1f7/EikRoqqY4J7U10PEr7Ucwy+dDr0pPuMiF2dP28AHreHyy6OA0+KNwP4FSANd
pidt/9fdeHUOozKfXOnKoCfJ0OYj+GzoWde9/eylsGp9nWrKdYaGYWuzE5HXFbWL
C6mPCC+CdHpV6BYYJQUqSuazMq1w72dCigsRmotUhgrje61FaYUU2CyjayHUiwyB
Pe4157iHepV0qcYg4/OTKKuNmpZ48kb0GVOBgr9Yityd7uObu2S/hmpvt+HdwfYB
R8iSpX9UW2SLiPOh1TZ5RYSI6X/tJdwYVBpYhdb4GZFakbcKeOv5mmYv7JPSW/Zo
R2WYHO499/hJZcorbM+Ur97x32lz0FB24fALEXItwn48uh6y1+R8498YudmgsvAr
iwQp6kRYMWMk0Yj/ELomhzhFtxtTB5eBHWgUV7RUGocaYLNlr/DTvUH2dqwr17IJ
ey1+A/dy4UPF1Ko5LorDnz3owo1GSgvvZ1hMOQYw4N9mNDMdVhEgYuOY++qT3Pm5
q+mPBai4JMuGY18yefoVrvzicW9k3lwZ/V2jlESGdXiUe7DbmgmpQQEGBekyA+6Y
XfrpWyDKiRibHEYETCPaW7fNgiNnOazxH9YHxENAv065Dt9Rk7lvEBlYwqHVdQcV
T46/Foxps5uX/41HENAsOrVsHRmMO58o0/1D/vpztHTA6hCu1QxCE1m9P2NOI9Sz
y+KsES4OENJNxqcUF1M+gUy+eJvPsE2nb4R79KcWBpy3LvguWPRjkUlN9lGU2y6Z
ODyl9+kVH19dkTMrsXYQcN1ZiabgpXkAg5sDEeDXb/C2gMyyRwJCxlKBgWHl2kJk
qFGaA2gs+MLcs9G2Oj4z3KACrIkLVGjZIJilbszZSszP+y2fuMZIAuwlCrR21DvS
+pd9GC4jX/hwkThB5NdVTQTP1+AEm/3srGMPxykefWNcPCgg4m54HFaJXCGstuY8
qiHdVx041pecoOKMyFqaX6/3LJHYvi8tDXsqwyimkCU0AA6PCXrNXOfj9hAUfH3h
vFridDOGPLhMFvmli5d/TOncYdcXuJ7uoVEO91Pl6W3tA1DNzs1h43iPsxnKwowW
g2rvsE8E+4ZpTdcuhIdI3jBrzOBuKcqKIggs2NNHq3R532WPAz+im9stY15JL5q3
Nt+86BHMs2Jb6AFLIEJSf+qGLEhRlf+oN8OLvv3K6ZzHgxsP6LaZFH17TMAMqbD9
WVvw0YCBUoiHe3Zc4tRKFTvCFjGKoVYr0dGBP+/NNzHTxP1B6t8w0QjVl9X7OLbp
C5ICDHcYJdSRCS+N5tWYMhssxL+fzcPY6hwdCRy5+ZklQUFy/8YpEOp0KVdMACph
1KaerbgLb8b8nEEmpId+GvM2eYsV3j8IFqXu+zyjrwIORevZbnzneNgjWH69vaRO
Pfa7j53pE8OSMapWB2ipG+1Qkl0VocNfdOEfXo/qux2v0w9yfdKEF/Af62cuW0/S
wNHo79+2359X9WP4MeWlgtPT9Cy3Kpg+NfBCZKk0PppK90PzMVvBIaBrzYDnQp1W
gz9yBM1o0bT2fpkZYgeAdKa9UR7W3qK26ZpslpR2bYjUBTmV62ijrhiF2mB0TuO7
lpSbyGLxIRTqsY3TvJrfcBJ0XB9/CIMPW8zF0yQCHz89XC6M9KRnRtSRzKbuyyIw
8TdoQHchoOrOvXjBwVSghoGJ/nARRBHa4H/ULBFxlpOS/EVHB8IT7N6dAOOR2Mfl
xoqyKsDaxzU+KRwXODYvvK7AmBHobxUYbwHbIpeytQoRoLK5ct8qohrhi5jrtof7
Uah+Mx7RzIiUxJYKK2YvXSDQaftV4e8knOOo97nkcsRevPQ0oqatOY/3M75eHMHL
mWqKtbzGYJDVB5KQju/hemXx53QWE+lMnhsiDaQAzyp9RRYoTnLpwKFCa3E3BYaF
L3ZoKzleZgSCIRHTITxVkHrIjgfi6/vjIvX1xIQ9dunRq8eet+pt78uPEfvCFX2g
JSAqTanlTc1soADoPvqDEt2KFP5gIDCnxXJay05e6mHcZHWercNpi3X1ihKtDPrB
ivkxqvTg55wFdy3QBPXQcSDYebP41U2dAyzIcVbEDoSUloB1xV355WPNyuW4rdz7
HiGfuOgzl0O5kgwC0MZOokqYQ3tWwgSD+oYsvgkFfxuH9Y5GZYEG2ciiAiZKDzRP
1dCI8t5yoT3OBnEm13keifmC5WFsOESKXU9fQe4aIKG4Nk32ixXKY5svh7iacwWt
N49n3/x8sV/+lI1SBAkg+xwGzEpH46v1OhVjvlkjMI2YjFjOxQEIBuAs5XugpFxX
aNSP8uitqPXs32gdOUnJnxyfRloNfDO1HHoMBA8Py0ZEpv958MWLzOZvkx+F6rnr
jBzReIOEeM9SA3zSywOiw3TQTh6//pYnd/RfRbrjiwlgpfgYWzJ1eBaEYVcsrzq8
Shm/lLFN+1jpt+8RF8ANAP0lIem+71Csi15A3HCbjgkK0QT0EjwUDdyB2p5HAQkD
Cyz3N+w47dQd8VO4B+bcpOv8SJzZ2oH73QHXTRBGGNK1gqhN9vGZ7eon2wtAGRbr
dHZkznjpHKgTOISqcIoxpTxN1jphvbDbjer0xVeOahEZzGF8FOxaWHjyquJwveEq
0lHqj8dYG/j429HH0l+AwYceuEFlyJFDLDWIrRP6NxOQVV3GoSL4Ij8lWBmvcLAT
7dWxAewRCnSY+NSBY2NjeHR6o+2uNgrjUh7mjsXO8gKby/Ged7+neym81oX8CN0H
/lj/iIJezPcHf1BhCxBxzrTGZNVdqFKDCEUAoO7MpAvde2kTTvmCr2oDGY+Drnpx
T+u8stXDANkBXDOtTNde/R6IOCgLkypPMFboZpaJsI8U9gPex4+EDrJmbgFBzWZO
+V05aIbrIBSuCch7EwRGFakqme22WZBADCjnnszvFYiOXSNMdVfYSTbrNFcMr8IU
W4IDugvY+CoTLBe1hmhr+UQ3b62F3cmqJrajQrVYUFO3ptpnM4jNLj394GSweMMF
8qDZuUkRqVh1dZx/bMsJHxhbadzIYNNXvLInyAdXFX7bP/i2xjMFSWXzUkKc4qDa
VnQ41T1/b+uPZbyw7Tw+j8y2Wrpm8P2sElrdzZ3kEMDGg94kd83y/dtmPYsjYWnu
xz90QjXVBat4Th/s4p48XPrvwqECbz9kH+aJwt6nlfsT0UU3cacoxmhsY0LRKSwY
y334NLz5txZ99ai04GxJ0eOOBEQLN5SBfyUBjjOu8hzh5UDAYCYDA41h3e1booYD
bYBLXMsTEG8N6r/ZuDJLiT8piqHst8rcYBF2pIE2KJnuEo8aRyynU+6CuhyQDQ68
hHOVkItIEVfpIXRAi9pbtlZb1+hFVo3Jm9mqW62GlG+3m6OJ/30QIX6jIRbEbgRT
tkkF2MF5eSQhJ6GmKH+jLGQlPA0FgGR1EJFw2Mqu4gHK26vTstD28sOcc6iQAngt
Xx4A47DHPvgkcvWeiW5l9kqtzndd6Zcr5chHqgqkzFtBtzlF2iz+jJ00wsrRPfio
v7FXMZn1iv6+6wjJ98ACcKVuFGlDOpnADXaNkGA1AJU51ATfI3IKvRYSx7n51puS
GBHCssS3+fcZ1dcm3AWXF0T0aPukykU0zmLktp7qvEgFgZVdPTjUxx5QT1BrE7a4
bLimNw/4Gnf+AzNBOLzbjsMeZlfhx0jxlaXvEs2CsNbOZNpnGcBTWIWbGICjJO+D
SQtUamwWz+hGivTDMQtVzNsALGJeFhA0iW9R4xkAintJbLnk1EPRrefCAeur+Jzf
9w8z5s6S70cOvnx2MeBKBqJDkkCKnxEV2YGKb/gZYQ2vTzEIqgioLR4KKx96BAXv
9GFuaye4vXUR1tC5tgae6QrcP2mgCT5XpGH/ubSLIIfZQtLFZgWKqoOQ2xKqoB5V
lIm/kTBWGkP1Ee/L0veD+/RctkkbhPgszfBTTq5+FPNi/DvippH1ZgJdlg3FAq3A
WGvAC15JRNvyCPSF2HR6dCxRJ7zqKk6cVm19BeDSvtd5kGM11VbWu9ppiwMnUVrm
WtcHIfWNaDtk4YLYhx4HHG2SYkzlnuxQjLkse65XYH7hqB8G2z4MB7Q5Z3uAAEzO
D4Z2evNJkh6Cr7rZbDr3CRybrlhfghbISZcy6jlHYvcQCy7lcK0uaAeMJJJbM6OB
Yc9+Qh4oBessv1PaN2J+KIZIDJUv3qA6s+GrSEJGcDVoGyBPZLl3n6a3cYICSm4u
D4+/wiXCp14ivH2MGmsJfYoNM2b8VUiSQUByZjuZC192sRrUh122by4cJT2E1ZJs
vjsLIIfXGeiY7xXmVrGUkUe4GTxZjF0oJZYPc7p8wb22Dm4GPzTBAfWoL1rm7vRX
yJEmakHXA82Mu58i7SYzWCEsWkB/TcwVjSJGE3LfxqFIOzUcmT69yANQIJHqEWDl
13RyzjkTih+zehyFqwzcS0vztNrAPzdG3LYfbbKNpENdzuEhAehkskCFwImRlPpk
xFMySq0FuXSL8K2kPgKVBnG2LxQ+KibccjcJEmFhaZfg0Jn2OXJC89KO5u/G7rNK
5/X36ZTERVgXythv560HlXLGnHk5P64BKIuJNTQsoUR7sop6kKAhk9q12f19xvSA
5IaFuzhUuYQGmrYKUF3zdmG/A74Mb51PlWMhNSepVzxZhzhZfz74wCL8Wgzu3yab
mJmb2hmty9e9BQ1ORNeK1bGZiqxRbCdtpG5vMnOsXiSvlLT618k9ODCYvYeYuL0l
bk8xa35OwPmrItoTHVYdXL1gsBdJ9QiaZwvD3ZvPAYR5SBCvt8QaHIbQhpnj+xD9
WNAs25B6bx/yT4HP9SDltot9kK9Gq9Q/e514r/h0Kc31Kg4FSRM/+qJpbSdjAuWJ
li1UNvRTys0t8uJzlnzYy0xVti+j7YBZzYkmrv/hjhrNe0ObcQDZ64MsbDpkHzRO
SCEZj0Mtzcbc+EPwx8+r3WqSRipZPgQUb/dhbce7S+kyOdh4qcay8OnilSi+Avng
EgbXqcbziXdJDDsbM2wya5fs4YutuJV3OADfOsVp6533Up64E00HAkXqJWCXGbRx
3qEncUHv4JOSqveY58auhxQTY0HhmOqWZ3KR4fKG459bf46W9atL+rRNuyLjGdzc
yCvCsnlrHuSdFAVSivVn4RtKMzZnZukWqkXAzY2m52VD316Vjy4Kr7lU82bDiJRZ
GVkm4EPbhLGZm8r9kQKzHywGv/jeaDEanunDTLTzZM9LHc/cY5GUCSz2aPz6QeIn
nkDemq1aDUZFy+3OtNVD8ESmXSFZrNAF36C1UgHNcV02VgL0MvrjJTHDq/C/SZL6
ZChaRxDrTY9cJwDAL5UVKA7Q86dTSEWvog6a29YL8bJqbC8uY7s4HOzpxez1Gvop
VKQvfMt9vKbzlLjlDC3+jKf2M2AtWfITxkNcGjDvosQzLtab05t+fITPKvGEB9Hv
8ZRZ/ct4UnI5eO5FX3LMhOFubM8/No6MWo/QpaInr2pNiiuKKeoAKtCUWGt+H1Rw
y32XkoDfL/5sXodGBfK8QsyZIJ0Dou5MJnlNuebAL2Ut69MbIR55CIBqwz3zJ/4z
EPjBC27bZabtaJ1x8IrgQddcWwZLxhMvzJky6IwYRwuepShYwgNekdavatzJ/Y8m
O8j4F3s1vB0CpmQmI2KIMIL+RbIZfr0g0KL69QADsLHW1rPM/TZaQsKrCVUPoQXW
n9PBAkembxQu5uhTCNIbrDth67eisCPg+LoMUM28i4xzjIozojGm3G6o7pFlXiaK
6HNzkvSBE1wFEMi6uOwRP1hQxMnbrAGQ3CFA+I0HGY4NJB4JmVJzD21WBV+GHy4z
OWPQfWzA7i70r3URF3bNetojuXVAoqySbtEi8p9WVQt0zbWIa0u2OvqT7jxOhcaU
lZfWn/1ciu2fzFR+5hZjhbSwWv7X0Wh0TBoncQiTLo1ZAiCHsXVdujjoEIF6aLea
g1c7ZVCRqMT5jv/CS76sdu9eE05hyywGNg5Bjyv4rWRtP44AhwPTWPkzfBnvR2Gd
aGknJXPZsgvorFah7z1tiLqQcealpdINWGFY4DN3WLIV6gDLNEx8Qiy+YcBWLJa4
UbGg0YDfW9qb+nFrwSwpzjvwO8VzRajpNS7ufDDkIBOkjUgdGnFn2R4jwNx6f2w/
rBNesf4ruv8qmZtINaO/4orLd1Jaq1C6MIFSs4NJrOMB9SO3nEFw0gtq/IOYojwJ
3HkMSF+9xs+AZFs4emOto7PuebeS1kjwWuWYLsQjDs5UJsqkFvIrpu38eEfKMScg
+4n3FGQ+kod464y6JXiozDAh8FssXG+lsTqOEF5dk6StFsIPghU8Wfgy2agvvbjE
k2B3Wwub9jgYN8uCx+g2+8Yze9snaNj4fcTIZdcSSDLZpcEboyYdC5OPpyo9aMKP
6oLuq/RHtHM+dnMSVoQkmQAnXVrFBCG9utxEMvQ68SJT4X+lTh49Vgzg3/BIj/RG
E32TZhPXNf7zClwBC+43uYUdxh2gCBC4BoTHyr7MSfTlc9lWskg6VZ8Y4mviFdjC
rJi5F/lPQfIV0uLpphVKbbIHJWHSMEV98pNVALn+ZJTFJ8UWsXkGEAzJRIdeuMqT
yt0q5xkjQ+F0MpWB6JKWOB3n1B+ZJB3+hoWWwy/S1WEvJ+mh9KNZcbLIlpgFk35O
Q+TLOzX26ovSOIJIGoClWuO48fjXv0ZyIXTbmGYxWqmUT121O2bC6bMkxSIcqPyU
JFB4MvV8Yhgj5iMFbOR1PubGTotftFoznuZ+3b+R61bdpEuvb2AjsTrn9/lhVqEe
KMqx977ctH/YJJPjmSrn81G5h6MayOfF8ify19Pg8rVurOby4sUXzoDYtoKSaAmR
dB1ejG2S5RvBKxZmdWdbwEOYnEsRF5ya+aoSpgdm3ux3FwAZ7D1bswLMIXtd9zYP
JQ0WyuAyOYDxGB6yShu2swD7jRUIzbePZ3/31U7NSLdPtyhqA4fI6nqCQo+AQSr7
CtMYqHebdbbQBZqP8/LOyWdi6qj4Bo3Oezr0zqcm+wqzQRRa7NGF5jXjn3bISCOg
1tedLa+Qt5ZKJsAqhc8vM3oquOmfbzgi7s5RHCSN7oX4Mb+0yF1Ih9gDFNwfqYTD
+PkgRUcvyFATzeuxqXy4QuikZtG2CTHtnPFtc64ZdlY1yzzk3pM/nS1pun5Jv1tB
TpqX1EbnGSXOoVvSWW5xkAg76uzPRlh1D1Ys6I1ryhOgko1ryPN08m0VIbFx0hxM
+jUKf8nQv5vH7OukBSyKzsnqan3FXGVioD8/N5KbmV7mgjnjvd3C85Umyreb31FK
dAGrkYp1vIWFhfq3iOheVZX7Vyjhd/amI4ZBUx/kX43VpiWynm9cOGhuJBiA/ccd
A5dv6buqxwYTyYBAZ4paxoMsduOraIqihpAGfPRGA3sqOXCmevYmRS6sB3E5PrJ+
SsxekX0E1WJYXoxWwsD8JYuHLcHXVQRcFjV7C1yFCi7669mhS/b5Lxl+XglgvBP1
BuUXdMDArkc8JjwE86do6r1ctFf/T0+blZWIK7FoRAshkxQvsTXdC+z3Nxg1Wfyu
QX2ZwsKogVWLZjbJBzfJQr2UBIf2YpywqkexsXYsxSuBM4fhcjtMLAFDXS93UWb7
4F5cOX49YDR4tmmMZYxOdNORWY/OoLvxA4rXHwMax3qvMXc/Rg7ODbsntloDf/Et
ZUy178Dm/SeehHVYOiog/dcuPxhlZM+yuHSekdwG7/jQWtOZseznA+z7eFXCArxv
buSY3w1rVz6+4ePbqUBKDCEk30st2yg5e6pMxRJaYV+U1pJLRQEse8OSfPnykb6B
GGT41fONk5Fs0dkS5zutpkDn51eXbIzmagwrDYzvsE1SeH1uABvS7ELjxc8kgEW+
UliM9hgdI/8EMV4fvEosNunE5F3BHopJxvQeZW7dPiRBkl0k1MP0862ZoHJNPAS8
g3Wkms7FMoq3wlC3s61IYT9knfIryqn9HhtZKj9q6OC2LTAYskzrhS2SS1UwqMPm
B/IQjFs/InBIwbR6b6R0ApqiGZxp/uTAPMJe0HXDpOIZyBYx8yGXQswqm8enwQuX
QV3Z1mPVOMkJ3ycRMdq6VTHkIf5ZyoqeQFGjng3oJxtFkHwWwlilXLhVym7IU7qY
ljSG8NzuRG8knkmggbkk48Yrf9fbySqUzyKtYbvFtG5yoeXXLLRtA3m5KqOP48nK
dk9zZEwGEXwYjc/Xeb5VvE8GCBdUKKIAff7EgP/Fob+85igAqYjB+/PymdiVB5mt
Sz76xVlyH3rs04+RTqXDq4jKrgHuYGyYsBSlm6FTJWmzj1mUKakdxcFNqzN1Ic61
RSoKmFH0OQUT+vtRaq71wlJAGBaWS3JbOvfVlTKdtvRpb3QcpLdveNEH7LpD5PBf
ESNx7KMlFCdDAI6+uWUardj7pwdWVL/zZeuLogvF9pdRdttN9a70EZRShgmQh7us
eP7ZDU/dSkiKg9V4a7euRgzSwdf/3ql7CDCLM13W3D82YWpusaAHl91bdEotlosI
4OMM622lp/Jm0K6ERof8nPdEuqe0q/9reYtcapJzjlzrGO6id6FHJ8s6QIcYU+T1
scw2PNJyQW9RrSPaHbNSyb3w6XMWPtdSRUp2qbVKBP8iIjQakzfFo2N0SbrouDzx
9r7+NQ62kZurrOTl4kJ9AL9ei1V9RIbmmswznT87k4612WW3NKFmur2UcBiR30wH
N/5dhNwr7e8e5buHzaJ7YkyGwoFhxmHKOQqo+TYWfpYvNzkAo5A4IvJQEA+jQg4A
fD1ogPaFv/PubWrrIYggRC/Rm8O79jZi2eR42r40a//BE7VOg9G0AdoXhKJSa2z6
GnanxOSwohl0mBKNkuvQdfk2CbS33ECJm6lHxxtPDY7bxZp+JA839mGSzfwnZRU3
QTQsHmBqxdOss+Ojh2bGF492KtR5i9K5OPXLEB1IHdnSMxGpT81kp9jdyeYTR6eZ
R1POEFuHIMO0VnUUA0zBNKTFpSnh3lXuRMuaNgEjcEllq9NXmiKixD/rp9zII+hM
5w1v1By/cS9LvUTPDfqaph8LRzptJrhHsPcPkp+8ylKJvRJrQ54wz7bdCPV9jujc
qf7tuBkHHggIH4Lw5otRDRmrgECbYKHaUUFraf2V0T/WQNnQ7Y5tYMnt2pa9Nvgi
NkLW9t4FJPOOpKKKRw+F3ax6gxPr5P9TF0z9umdFTEklCIOIaCFapR+mZJBSFjh+
UruoNPAQTYoTXRsQiSL/N5vwTdedgjQ25V7uBY26SEo/q0eqyihDtIErT16OxShF
o/fz9y86S8vhlesdom+JPKEOdzZeo5IJ/9ZAdvFY3QsNvYsWeC7plohEhTxKqAni
BEmy9cD7BHc/nU6OuqAlcTO/eUNWEY/UkTqkLZxEoOgLN8oCTycUrZhxYb0d/Pte
rlyWNA5ES0lIxtHHBgiiiq8MAH/7VwZ72UZQpCwPfuE5NWmOFiYsv7Ch5il3E976
QofThGzGAUoMQuJDHBPZergqd25bFEiEc2GVeTm0/HMnT7ydc2mF+zNE6FaaqYSt
v2LyDjHSAjCrf0xFrVVJmVvT0CU24HUrvaak4ziQP0aR2/N4HDIHd8gJdAl75a6h
HbGQgV+sZosy8rJ6uPNZODtUUWlRzBmhO0bnKsDudezOBK7DJrWA8HAurB2+VVDs
QblwvvfjXd7pPrZWyYi5GcxF/MjOtinexXJV3tVoekO4DK08bLM5vF5KVtNl8q5c
M3wxEh5x6gNIAMi5vyvV/SfsXtRQ+PDJ33xzYZBPaipfEXbKC9hs2PemeTGEqX88
+sc/uzOUyCG2jJ6e3iCgR8MZybbE8WMAV9DT0WSU27k/PhUbqIsAsXpwAPocaWq7
UxexCrkLsil4hpnMgWAFefwJCx4u1rMXCp7pQ2RPajFIoPSYA6d7LHxWRn0/7MRH
VfmvdK60zNufwOWZXGptpQ4eGtOvyJI8feA7sDHzdYKSV1iJ3oYWkTNmHffHVivS
MOaVw/0yB8bB5xJG0uMJnQ7fKp650zwKU/NDffK9M3crSJYjIA/JUqKBB5QOQ8g9
U9ea4ABzdVri4pUjTEtqvLMNS51hMJOjOx9Fuf6SwhwCd54zFz5moMZp6uaKAip+
dLA4wKekoSLHU+9+jeepJwnbste2lHbYu/bpcB8DYcIH9d2bIhKanAhaauoVwJhS
nvSrlvv7/m1AoOguzOdMZwn70OH7FvspcKpW6zEx+nBQJ8hKzSkBayrJCQ6N7QMo
6Be38VhqRjTHvH6j8bZhR2I9o1Sa3Qf/kb1i9fYSkwualyiRljpPHapyV5HCdtQk
WYDBqV1vUzvAKCgAaeenYyv6iAM4UH/GAF8+7qnWuh/gnMvoDFtWYpSf4FEtvUZ6
o/z7gGULsk9pClQevqkbi2wfEXke2EW3ArGsuvd3oxY60JVyJsjCHzVb3zv2AqrI
11GxuCIhjv+2eN4GvHmPxI4DCvtZMubzazG5QT0IvsEGUFlnPcJWsbBGgc4RblA4
NMmyC7KqYTOlnL8W3HTWn/w8CXSWKG7JiJVBWNJ0adn8YX98wBGJxUYFoaCWu+L2
fKPv0XDz0x1oyLIf1Wo8Md47X7bqrBE5qghn/8uAeke2AWMxXElskYvyWxZPzHkC
e95aN2S3+qGXGAU580gKGq5WCsXy71PR7b1rUJT7P+u/20okzFad6zHTN9jsDG+e
JmYBwbxi9BV31NFYbJ0XBS0K57iZDRQA6megMfYMlYt8ijQuAtSUCBoZK6nD0dGz
p0vKqpcn5vw6mtmnyTJHeDkAEKuK7l8MQLE1/qcX7f65KLP8yE/MEKiSnuDGZ22c
8z1FeS639diPirXSuFtZOe8sLT2YrfFYaQMBzosjzjLQybl6aCpUteuSawSbPNof
0BnOe7HCUAWmdOOeOpbfnOcAKQTXKEKZJiNNE3JsY9h6urKM94abLqs84PE8ARDJ
QsQs0Owg6/sjyk+JpPwZOnRaU+XqjSPRoLUPdPHgBxErNWmSIkzDp+yQ3C9NhqPw
rYvvzsZgBU+9CnuBBl5/2vHUvsLD4dSecaclGPjSmqqbL2IptdfZ/ooDMdoQkIYQ
kKFxpGnaioxxaUw5QwO6oT//ZczOcZxg/+w1Vq5oCLoNY/4A42nqZHLmHLK5JbmK
OpoUmGPncD3+kY8oO/9O14mcCDzRjLQ9DkWRwLCtwWPUxayZzIwfKkHqd6qP4Smz
KKrCYHEu7gC+EzvlPQrvkKB+Kz00ykjE9feK+kHuUsf22cC1SdsdiayMPblcq77Z
ANQN6ZCPqs/vCxvowTH9rUA3pE7EgnBmzBarieKXe9NzGuFKD3jEG+nHbyPDGoaB
fKXq4UxYaz5lMzwipCrLP5FFAll/F99Oo5GkiDCjpt/e6BqP5t2Ho+6i99qrg22H
XCJKz4zy0H9uuIf8hLfk1SR2hTEysa8jDAGTebTpYLwp+DdonQlDJPJiFQ4spRH5
ncnVCOm5HWeN/QwMwymKonxeFByQMsKxLJiqrNttsDGBkvB5nV51bGyq9bBJAGkE
NpI2ZxQBWdoG8/wy7bnfz21NdyLzSPZIPY11zu9XkivbYFEp2pFIGtSv+Bc12KPf
jfm2zSWl7sXDg61Jo+NcEDJntkXPNwIttdYKxji6qZhtiLUYhjn9yo3YmkOJ3FO4
MGQouuvcO80wx8IRXLMec6AOmJVSUfwkYpvU4nlE/483z+blLzlIPkmvGb/wZLAE
iewxoy3fWPf/QJcQ0y63bX+Wno52W/dnZhCmrx4WdtyNTRwIwe+MnTUlHH2FTYYH
1hsEzDDJeZVF891+y5Jj2ST5pFBphwCf6Mi+ADijc5oSblBi/cdlp+aD8bs3B2DK
xg30VWB4oeIXrexuVCCJxIRcIkPk3art5qP/YL5Byn2/5To+o6OTDV2xvarNCc9j
1OmzteDSdcmrqkxs1wV3qRyDQ9s2bVWfZE27Pj/AIxsSgMfg3mlmQfw4nXKxZ4+7
7uobHENAHQWcSGU2J8MoRX8CNlkSehDHhRhoK2PTKDBXGxQ0t/jaFWCiAX8pf9Ga
GqK1gj1/Ra5fTHVKhTGofRN6l+Ly1F6PQEoGl0nuUrcRPW1eKTkkmA14JwkpFUjE
v2N2wmHYn5I9wRWTXj13TAT+iEfTPKms7aTfbB7Y0/fy62U4h+SJupPoKHoNRShH
mqLGsO+uUHRPHCfY4VTE4ipWmwWCgi0sFDcH+EqjgHdtUH2OPKg8e9EeEQmmTx6z
U/XDNuC4TOliL9T+cc4FZ7uYRa3yChE5xqTzdYK1S5ORNZkYUdbnr3krcx4pl4lY
kdcswLdaehUMsW26eBbKynWjYRkm4qKOcPfnrTZ1svDEzAxEJdIGg7HzdXV5qRfP
af7MR4IaOdAEbafvefxAAW1moKp4nASSpOB8ZLncTeDsNkzxMcenXLS/O7nmoMH7
xEPs1uDSYFj3pdtCXIoEllLLMiyaN0ULgvDZZ2V5l6DDN79aC5OmRTt3qO7VlbWb
FTXf40aJvlMCeGL8puPvVakidm/wzRcHhQjWOzup2E21v9F81t6OL0pH4ceENWjP
JQMyyEOz2bbJlWqC/m0QGQBfVGnCQ9izQKwQXmyuvb7T9KuzGlfUJDlnPEMEVAKs
5Wb5cDSLSY96oeU1+Te1HwzFC0T8aM8xGEmsdA+PAalklqgSquZ2SI6Gb9ZFQ+Ve
VTfbmfVVj3439Ifoj7maPt72G1q+8YmvpAM6IIETxip/f79eJUFZqKRVOcFX6j5K
o1TTv0M8b4z7uMxCQO75ZAeN9g6G2ZMCc3PkuETJ5BAfLgMPMaWCjOSYKCg6NuIC
nPMcrJpyb3jtIqtBH3mHvRS7FDTbG6QGmEgYPL76rKuVtyrJW7EtVP/6Yi194eZD
gAYiBfRMPv88xA+A6Y98YdWA9qjgOoXIQCOEKRaQbSO96IqMNeI+EKjXCot+2VBd
2EJjQ5CUWJTcyLgeHW0VYUcZGdMhP146KBRUeA/w1tNFAEnfqTFs7PewXXRpiFKc
KhaToCcWktK04wPkSi3ja6hhe0TVSbza2Wej4s1gRuP+ZGjdazf3Bo6WKIsGNRsp
X3zUnuyRZux4XKLb8YaePTQUm+KN7YietZN9UMbmVxklx5BCKTf+u1QTXXFJ30T0
ngbHWs+jznRp2u/qKDh7oLSUr+ZOl3gk5KEuZy1XB9naAibyoVIdKkpm7/xygh8t
I6JnsyNFNW2Qny8zUicgH/93MSzLcR/ON7Qt9dLOzvJIS38BxBM4jj5UWqpEsq1k
H+jRD9YcNcvt3FCMf1G/ZcEAvxaD/fdxcblZgu+RCoYBGyHUIEqTpu5sOTIb4Ut8
aJ5Di8TY1fRnxMo8lrKGfmKA6Q4spltYgpnNPbbwyU3m0PFkD6zvr53at1mPnWTO
oemjdsz9iZ2kGHRZyfvoZ6DJhN01VYBJpB67OLcF4HOichgw7vm6dNZyfMv6Fn/0
Qj2Dl0dug9V8G1Yy6JF7QmMw5awSY11Neg0nryEer2QWwqpyJlvmY8Z/wK2WtKg7
vWH1X/XnHSP2BjQtVUJZBa6F2VL+9Q9bQErfCLWg4kQIhHNioGNmSXuND0xCBnft
u2iovBN0WnvhKM+BuEAuUjb1mLlyGVT+KJScEk+HfCxW7qc02UjT8OrjXH7E3abx
qqHrbYrkeKUhDuhgkIjWUerionmWWIhygN2cqgTB4NHy4Q//kbVcIRr7M3C+dcAV
DZTrRClWczUrUGBIMbge6VN0nB1TBYNjMeWwki+NkJjlfEDwRr0IBYjreWGaf4m0
2Ax2yLRIUV+OmtJRrv0K8Yr6SZUEdEvHreFqljO+Wj5s3MBa0C+FNHBNksIfxxJM
yUl3/ohLRuALYOBghl3q69iEH+Sd69SOF9K/PCKfToyWK7Gt5bwOdOU1bxbQtWeM
BE0BqRJ+3iQCRGoCnaeUezDzuFUSJPowugzq/lKiUiAmQzB7Hh2LUbuCIL8bWkHH
jpXkoV2f7VBtKSYkmW0jRoZiRH7s8tJpD5bnZBnYie1oavWgnvLNhBmUPChg/+jj
2ca0VMpo5TLgzERyyf9sIhmjXDpVdlV4RhWa20sBr98uKMF3cLZB2qKBIF5UmGLe
bXRPsSHPBK4WkGsW7vj38e4LBIX9lbwRA9WwT6bfVY4Tg5tObxdSk5pv2fSn415d
L/zmUcSDqcEpsQDDMMjc1ximyE4dyIWl/e9BTn/KLUyeSmssKwNPTZTQxaJGiTuZ
AKpGTBS6P66ATEVL7U4IEYFiWsAWQ537Uz8OTecV6vWqclhuVC19xXQtDmEuQkoh
xhFE/Dx50Mf/DvRRsk4OUk1ZUGfQRBp8LdJlxPRdmaI0XnfzhTbOvpMj9PgG+9gB
Exsoa7OiYns+F5SllKlOGx5F91FzdMgT8EMOwD72j0U0s+xojiiHnJbi/mBFgCqb
At6Ab+3hMu32tIuF9fwneq6atYQiLLQxvKYAYbcWCARXROkZUK7bGxo5X3v5EgOe
sNXDDiBbmMIQhuGMCqEGKAsks60aZW6drbfWkFGaS0fXfVvoeVLm99Yebiado2vV
g36YNhtj8Ih1GRbpS1ZXlkpNtO2AbQpWU3p3jBIz5CdN3dydZzJiUiohSJVJhe7B
LbDeY9rW3tLuTy0qEP5+0BdXuHaamG0KS3ei+dqvSEnBw67mRHSqvgRUApdVoPfA
Eg/LniySWP/Hun2Ud73qcHjcCgVQM/JPQCp/m9OzH5HlFn8X1izSgXoRFW4T5S8w
c05Dymcv48+Wu8g064LK76INGpAbUCKkrey83OAeB9aEk9NF4GG5zOq8C75/EF7i
hwEvGAnjA0SNHIfEtqm599UmYHze883HKJwTTISj7DwezaLZZDuwSsTm8tNQRxG/
wYmyYtPcsYmuprKfVCfruT8Q5pDgk3E2pC2ytVEwx6q16msr1wRG6VqBGoZaV8ti
AAFRHTLPKUC8g99h/kgY70wZrVkGLf9YVhmxyJS81d+OlsG/gerZa1U9+EKRDaZs
imLzg7SekDXGnXx0/5ZltpSqKI8/31J9KjMXPzsNZuKlk0ayw9InV8RzTWPtwtLg
tspRk52sCz76PPjFBtO7aHTYH6Wy+XuLat9FJ108LRulrY8+mRZPgrgxEe+CfKQ6
3+S0iS+h0v8dBDJkG/jrHkPcHyYvA6l08dR4yAaMLa+XjSRjX7QLDiMimGcMb6uj
OpydHC6nsIEUXqRjjgxVKndUz41K/f9075UjRMEYGikg/pnzzePZ9OXEYkc66+x2
aA5/MXxaicxSJPQxmaathNRAKyz6t67ZGvjbW2NKG5U4XkNIdtqQ2bVRwyj8Uj9N
rCGJSPfbhlVJ2/+P5VwlUiNBM4o7y+dRma40bGByiDn+9HXIho4UkAwFFubRLasj
rvIJihQllUwm3Tz7BRu+y8DTn5v58L7dbXOClrskPygzn6gIJMJy+vhA0/sDOKkV
F0hGPdafyhMJeu/VEHQlq5SDM6MuLq/0zExLBQmLINM5bi94fY80/7VhK1mVKSTc
7QIeGwsyRhiwLBWIgsuWnLyUI6C18Q+H4KCZkAOrLDGUXAHv28UBymqrO6kwLyLl
kf7RwX4415lTLv7h1ziVikXuzfGwCu6zlpOc7F41Jb43oDGRZVoNWnwO7XiWxDHz
7iO14rkGaEQc+IHoKYqzScNxO9vRNuiwcon+cMK7neSrzNlWhehLiW8PrdUJU9Bo
lFI31SWVRZciKoqe2ego4stcQANzppSy8AIYzIk0DSp3tiJvwtjDm9QrG94XOhz2
vjkbOWSnqmgoDNbs1QQei8vl//Fb1LKq6eGSYKKExR/07KDZD21wVJHZ0JllTaDz
MI3sl0aGOCmIvIV2IYXvMkl5XHCIR3hy29mXDKUeXdKuRZzK5jJrGlGzVITMpzCZ
vHrEfBLtLDQs1qtTq/fCJRWlIagD8WcTPKtq4RmxY4o5LflezY/WUJY4QucD7H6s
Z83Qqubr5578LQVOeJ0jggmKdBtPqMs4jvFAdcr5gQWzInwD3lKf/fvutN6CGDFn
0eDopj0Tp3sjGR8B660+2yNYeE8SfgPzUxm77q3pbh4gyonkCDgjGdEtlDd4Uh8l
6GAFUQV76WWweXCT6lF2X59wbjM1E3zCzri5/Cuqu3AxgehzTZiokpdgaUEEvKOj
Fylw8JpOcdYmzLP+OUuEutN721j+6Jrj50qWjS7ozAO5sNNiEQmTDsPi1aSXRU4W
enQvOG0WHgRY2lD02KW+pgvtgWtICgR4sSot+ohMHa9b0UAnfbCdequk3T5YoaVq
4GCnZuSk1yiWDCWlxI+xBiXLP/u++7nFx4z18M3+zDQJbqIsA5Cgnp3YV8PkJJsY
b4P0cUQ6gx7mo7yPIghgW1SpDeTUyr/dE2sSPlRRKuUR0XOW9Y5htwoKkzr9RCyN
uwnfAqjeq/cNAZ8BpyUF0B+TPDxe43GKC4QrtGi8lZVhQ+vE5takpD10m75xPKri
9sUi7QDWO0ji1EYghjtSN39whxuV8679fIvuW4p2Csm/NIPWPTDOz652sHBk1GZ2
0capcostvhnrvEORdswIMmyhZsZWIIoum+xqVk2zR+VYH/D//oIBsYUfwsZnrLmh
2/Bs1Tof3dJbrjNyAq2tONSv5JO+jlO5nloMkc8rXzGtgp3QeZo9Ap2LImeFg1kM
pb6vFelJtfH2UZfesJfOSLBw5syizR6ob0mmEJlB6Cp9m4Vph3xz2/6hqcAigKDL
RvCjgy+pSWyDiYRdSb0poS9oydb2UIK+9e8acDdyQKvd9zK6mfH1NmCNTd7f/Fwk
F4qQj+zBtHKOYrDZPXuIOylJBhKVmbETmIzTHHXObiVZJnavKSpjafZjxuH3jX2J
aRUSjqyjf8GTRUIun0L3C646bDMXvMwCMcP+adDaMrhj+WSSPsv+sCdKW6Jd/l7f
BMnQAwHJ6OPmtvmGl6sDHAQOQ8ZDgLD2UgsKVJlRmrFPnz8cY7kQoqlUcKb5yw2Q
PhiiqBvrNlZ7eS7kbTPp8jnn5Pciwiw/m8IhiPH0Lo6KhL6Fcxg+etlEeLHrmuo1
PlrtFYLxAeU7sjoy+LYyT0DfU6oBZuUJyFbBkzPd6l8ss7feWcxsu9wVLGwNLqSp
CI72rPX8dgPAIlmaU+F2SUwOcsGSXW+KtBCUDgewb7anqifsKCsHOM+mwZDRPYqG
gNXsIRLhHuIU/50uoVjBxcT+FCtFoVm3Pkc14+ngWhRmkC0RqzI03vZVMtq30tS8
XEGjjku2NdHfj5OpG32lNEozt5peQJllPhTFQqemnt4YIXRD8SHymKo7tchrchZX
spqDldqwNojS0N05l+n9bXK0upkgDUYaBIVEbZQo4uOYRl/l6Dwhqg22pLMs54fU
QxwTOor6sg6GlXXG8Ky1GNkXwDqJ2Ncsf05K0aRC8Fal06AEVmMXn0sk285unVrS
FB220tUzPlWtM/2QUARQMZeum4+Q93d551AgBMxgyyxFb5HhF4BhKY5zZqqHXhv0
41rAWxIuxiLqCqY6FsAF1nSMUQbg5D/niwfp9iv5W2AwiatAQ2gL+MSkcPbcXtIL
+uLE+DjJFcF80p0PdKCUv6i7VMycBbA9v9b+wVYuyLRw5DI0VORiAJzWAFIaUC31
pKx3H4mxo0agydJHb7XLcSMe4r/G60j0bxlDMSrMwxv1psdtt6wX/jtgDhckPRh1
GIEXMt7ktctZFUWcqN7JdVu2WsJXiHR2uB2bT4lfZq9W0cBozfzuEACglC/gsEJn
TwEfh7krTg5GOw5LXUlKH/qG4EjVSLDYB0urDxeiMomoG8uXEdT0+B/NoR6Q+oK+
jc79qRcbifE/X2RP/8fbKHsusoC8/L/w8s5Lwla+zJaUnnKqTH95n07OXLzJCoks
xPI52Akri2l5WGRvKA1KokVcZKKcqMTVo7y36nFUKai5y+udn54eCI07JKuBW8ZF
OpO7HnCfF8LUUXB/mYBb1lfLgQFBzujdkG1Y0Id5HLq2Gq/fxCtOykI+4sgT6q6s
mCF0QB2VKF0neoRCILp3qHTtm6ebcz8Vc6/crIoVaVG1JRtDbO0dP/9vaq4XfGyr
nOI6TIxeRaBWU39tPnZV2rxuAiBZjNnpwAXrLvd+xZYKq50EnYTfS11S3zLTz3va
zxV4KuyvB/WdDDsePkEJc6lLaUyxpuV0hTvJRyXaUMLvRhiibqwx/87aShjbLqHp
/V5W7JngNif3oeOJt1ldrcmYJly3HFDLXBRYiATsEwbgH/LwkM+oXxsmXuSqn/BM
dYFb4h0QiTW2dS8EgGzqJQDr7iUUXGnYoDiTo3XBeJ82Mpb2Yv02Tmzrnnzcq62n
/3efJUPfq0/jBTkxvPzTuWLeRo5YGxS7A7OEx5+Wm9qdTBihT/gkN7xEnjGPJsOT
pj2cdGRfL3WT0psCRjsheJerUTLxDv9p0WV3u5+CNzG2L2zhPXXhApob5kWEWyVo
B2vqNihyOiEVlEU4aoOLYyLIbcsaHPNXp6tt1jyxIV7CdTLgRtrcu2/tOorhcbKq
Oh/Ar7UTmuH6X183xhoEuxZZ+wff9MLOKFcRr+QtgQAFgTXxu7D+fxopX6Hj23hT
XG8XxhScFGKxu3Z9rwKyaxO9UGzZjji8cT4vC9P+8RXzTtotIAPUXlQHwFgw7pe7
O2UZS5Iexe8OXLXjKi4xnTA8dd3kDXtC6FrlFy7/h3g5RoyctW1VQzJu8a/Ze2ci
ZHinUaWnHuP0L7PRliFGzeurtPyHGiO6mDg39sCKpfnP1ptkgXHR7t2XZmwRU1Kp
f16LL5tN6KvXsdoNi4mtpeNamxx4U2kuy+MfI8lAr7S7hLyoHYtbEVVuqOHsH/Cu
/F1MswqsQH5kgrh6QF8K1+Z87PrH4V/Q+HWgXQSt7I9/TvioeBJGknk9av1+Blsg
/Y9d62rKBBBZFoglTkqHyC2vWkGd/Ha3NuS547SQiGOtnvDM0Tq15xxTFMlp+8zM
BC+0B4WZLuUDufH+gQ38Hes4QS5xGc5Mou9WIxksYgh7FQNaA34Qv5HPE2I7sTVt
sif7Wkrp4fPAsT9PRQcLHqdmnHumpGV3dEoGLcNYWm+S+U7aZ0dD0GGHBTg6wZal
Ip3gM1RqX/RhCONqgnLeeZPnzBcD5HgBBTmZHCJsbiBbGN3wrKEKFSXe87Pcnwfx
LN7BAfij8YF7O1RDf48LUupOIpM3Cv6ZrX71pzbDeikx41u7lmv9yJonF24vQgGW
9NMoMCS4JspcrFATwSC3n0U2/qkI+GbY8Qv85CJHyfnGDmy/2panKL5Hh+78d1P1
BqRHkHRgsjKcKYyH0HLlY+Gazp/GUcnBRbiroRID7hfOss9oKQU9ZEf0L93pHfnl
Zy0Zy35j2NVpsW3TtLHZBGb/nrbP7H2TpvISg5BrnM8U6zMbtKAGquebGxfv5I2j
tds+n9H7cV4KeHq7q2gWqDf3oyoqw0QE0tri7Sm84CYBrtIexXRoGfuQ1vHxIHFt
xl6YQnSy/YBBZgsaVjUs17QE8nfSD3Z+wqyABOPbl1beM+6R7aJbM9Z8/1W9gGTZ
N+PiUZf57GQvd0LBLy3yaMLRRSlj7OOTPLwP8ibAyaziBMwhVG309zsAYJRiDbbW
+sqUfQdKEPi13wI/FpYzjdrXzQwNXuz95IhFHuIn32GwBAfAT0st8airMyZBancP
jl/X+ZUoQsnoBXqIqymAEB7iwxt0Pexejpg5uenG5b9+hHCTDB81OVF2igsbSBV4
9NjaLg6jyZF2NcWZczd/wVle+ALaIuth46J714MF1hIW5fIPmZosPDbTpK1F5Uyw
uFUTThkYKmZnCDpT/zLJ9tlKyLfR8B3+NMeYtYTEhJWEmtvZou7ZaYKgvgiq9CSY
7O//RQdxd7IOc9NdleKueNDigQUMNivANhgEDuqd1PlUUZaUSW98GBoZSau2T4+v
oNBt6Fy2SyxbpaHDdQeeVWl37n5EePfBEikWgPXDJ97J375/EmRcQzcOIpu71pEY
JLNIEaOxFuPD3qMgDRsG2MtFF25ACBTyIChIrG0dYnx6JFcssO4kclZ4hWeZiVcG
487/UsijYXYaZ2ybRDAghV7bXQHnMxRz+fMrT647FDxSgDrXhAoSowuQgUbTGKiy
9EJzog7Xdw6mF2LiViJebGs1otTtmnekYoIxQkRm/xTSNz+d4/d0gJYM8Eskj32y
XdR9rdtQE5X9UyoLRXWnMuIx2kC1lcQN1LhmuO8s5jZTpTYvUAAmMbEGePe/L8oJ
o+tALz0Pb1LD3gMScV+EdAW3lFQeDpNTFi2v8l2kL5zXgMjO1vxILwsrF2NZyGkT
hV5IBDuUwpfOYW9Y35x/Ye8kqNgbkyKMOnvmZaQXhNxFkkk3+1ePhUiglh+VLtRR
gBnhon/y0mXuBFm3v2h24IU3kvmtq3Q6q6HzSda5cSLjddTz/yj22oCpjNMs373k
NmXwjqgtFzZyOl7Xk2AjruGJ5Mj3vuG4tp/HISt5OntRCx9Hff+VhU4KAr2GzL4I
K/Oa/RHmafGtqCNV4indRjhdq2ZQzR6rVXimK8X2czzmhj7Cv6EBg6Yr/vdU9+sU
rMIYN+kxjjC9MIWu4/2CS2qG4QIYNtTkmvcZj9fm7SfvV5G9v/zZJZWo2Y7bp/Vt
Q0jra/gt+bYzNWlSUGG48RpwFU3TqdT27m39HhMCo/zXDyWdPfHtVMuX4seXDP92
YupARcPyOCVujEnU4mkVfTOUtZF+PeMdIHEv2Aq2hPM4vrb4nt11yD18dfxpdORA
6tNfTmbqI+1bbwe9Z9UiFEP0JzTC1oAsOtZ7rVWb5DjSr1In2s+8qbSPI89+z1Cn
/p3VF2idczFfCHJIRVh/WbckXSYZx6g9uwxdMwuiK6tjvIZNaYeT6gS1LVw9jyVf
5IOdqqIUbFqXNTcnMeON4Aw23OkONOrH6d25tYL/uWxjYMVyGWkBpaRUhJFQqfmH
BQL8c8BWq4BwRnzxaQRrCESnQnzeWmXDkOqQ2uivdfrs0hy1guN71R69NUKdrQo3
VVdQfyc9QU2VXuifu1mEydnjyBZBueJMBsX0Cqs8rEfVvSEfYliy12M5HiBiNDTL
IYoeumHZRnL5nNP9Mnypb4Qnwc4i2PiQJSWwjSOfcFAEePghOBXhCMFJKG9Kel+B
6M7izO1UYIfgqxXbWZFqlqlwhRkZx4CFKKsp5PGu74szJmp1YwaGV0hniUeiIINs
T8U2Q9ct3MCpmXXQua+QQ+gFUCONZ2CROAyFpjp64J48vGEuVOQagi1CO4NIINf4
E/6TRRBjDW1aYAPiyEtlDhxgh5BrqhWMA7yQk96AFyWUoN3ZQfq1ck+2TuOgT36z
g7Gv8ZFToUZraF5VQYa95jM7NZj3kXIc+RTL4Vci1B3Sjd5/TVoQNLMgWEgUpAvW
ax5LdbNgvxqc5R0XZNxq7kBgl1HlLIe+EPFrar9JlcaHZ2Z4k0tIItlZo9B89l/M
zQgl43/QXPTo/2HV65RuU/s6FJGpS11FQj0K+NzWiCs4knSOKqNvKsTpXiPCBvdH
bEddIel9d0uMGVQ4CY6mcb+vknYchicCVahsINQ2IGz0Cj2He+16u8XfkP7+vTVK
0mhQ9ZoGcT6cqWOl0dcRgAEsdVmcJQ0eMy61fOtelkTCNkUNBuz23skKWdrDeo9e
EnBwsG/K+i5lw3+ohLjoL09YZLu90AcnrZ8YktPd2gQU1ZgtcvFxlkQ06HowVjwF
bIPJZEzAed9PsuxZ4HqKsPWZnxkHW7h43KSVD7QjSyX9tiHnLDN+uL2prj/U9+nK
vSeSt/dlr8LV2q77HWZqfM0DZgWjASj5LjbV44tq2AvYEGIz/9lLITOVP/9aJEQr
TMXr/vjWlC3b92usAsLkpzGZ90TLyg00LVTqM5wOQzGBZV/tuQdP1plhNkpYyF4Z
BK0iTFBKaG9EAVsh0PhBlknrkkYNVJA4Zh0pfxgnZVjC1cFsxGwb8zH7MzcA/2wF
VFW5j3sKtwy18ms0j2SSXqO7Wvbe7Hop2XXm7ZjHuDNKk/Y9JcUbBmXXOAEiC4Jt
/eDwDUh7j0a245hRocS7N5oKeLSMXwOkSri+ruqJs/3InuUHCLr3mddBC6ENLhHD
KvjeBIRNxI9VeXWcQehqqqG+RZB5WaEBptzOc9nqObqmvU2E5ruHFdhvRCd0Nqpl
gpI94HzOpjaCTK6Q8mH8+SKU4//bdQegMZY//ZeFAOrBYq9AKTc/SrRzfaeGmxND
B4ozu2ZIUeDNC5QAY2v1rGSjWpXH3GWc8BTZgk3Y24yCLVGvikmbXe2VHldj3zxn
zYn7yB2B8Zf6oL7g/k5y/cbb2zsJJzb2Y7EmMtDCEDpb42hdZnm1k4BRlvgRwb/Y
V/kuyrvNFqvAZ3uOz94BY4DAg6sgfl/1P5I6NkK39Az6GgTgt+4hR2PUxBuOLQbS
sb3HUOeMLA6PHIp9onhaa1D/6ynqRiz9Mu73MsBYQZTsBuLoL+tw1xUeCWQ8jm/G
1J/ni9w1LR/hCfDpll4kJySMiEpTSHGdRotEQWc2knPozOiV61TzgDVUe15VJeGT
WDBsu7VNpO1Bhe7J1mwBrDUMK9JMa8lNmIbiCvl0X10XNj38ReI8nzzUWxX34kx1
8VcDtQa5xPolQNhyaa/K1LmigrGZwjFy3SPU8eNdDiijo5qO3C0rgs4D1pDnX/am
t0yBO6zdyrsZu91SAVn0kd/dql5aNt/7jWgDfRFKe2bnAk+fUhh7PV+fvRFhVIfV
5iLYUx0/d9gIUdc7B6ek6OKdRYvWZKjqg8ApEhUyEqcq70Fj0fJ/aVTMVwD71ZOT
v7imrPAAJsreN6A66vD+QfM6Y+Hsb2/jprgAL9U9v6HmXpWPNrdX9AePmbZg9V+2
lRerO9TZ1gt1NIUmosKAuR04OmezMZSk3t1MO7zvdv8kvQ92iE6LBgGLpoIYtevM
XjvjkaaLcyrMQ4COVFWJwlJ829n1CbqrpTjtS4HbYFxOW4hDllJ/mydGy+Fk7aBY
pCvZ5M9lDH6ySRZT5yO7F8E76k2P4StQ134pV+PoKDEzO7kPd3bJnzHmM3+cGgCB
ID2EATsaZU2EGq6R2r1AytgzBwb8Ou18VkEXwuoZLcytI1BCNlEArioWFX6j/r0W
Ie/aTB4pgoogd3qX+pe7CjHiJyK01K0YyZGjojPOeLQKeBgoWTRyOQYXnDvS2vC2
uR90aDQW6qyRsotNl1wto1zb2rsoEQcOhd1bg24W58oq9scSsb5HiFYZqSNkOhry
qvotK+yg7CIHZu6tvfkca8wMpuPhF405vxfP0vmEA9HQiR8Iv/nuHuLPKEBflTe9
N3ln8JhhkPsE4m/QuEA5mvyLbmsC/sCAHlLUdYP7efJ0w029jExrehTmZVr2hZyw
ZIn1/JTut4QkVWSP6cCIr94kQ3fQn9u/WzOJ+an8zh20ah5x+VCKiod0h5tAM2rV
749RGYzz0z/PZhyvy/OQXTsvX4rt4wJwP1yQ+ZxN1Pf/PFjnGu+atacF45qZFbPW
92pLlfzOzw36GHrgq6Aerd6ha7NrbMFBKeC1GQ0qMccYn2wmotR1C3OO5rDorx4N
mLeIeCFBBPfq+XprVzVU5I0USWJbfXf2ZPpKtj7VWtgc/nlOxZEWQv7UmJ9aj3Wn
CEKyMi+NsPYXh4HbPB0FUEo2dhn/vIZmRvA7p/0xjh7AbdMGG5tdIEMG5vFHoC5V
nKtHSiL0IGggmyNLcBlFL3+Ia/AzYNqilWdXa8z7AZmQHWTZVthrrik0TolqhmhT
GdC+oD6aMRHsRH58jrDnmtrsmVh+GpnFj0A57x1yhbt9lYcPhNrtq8LzlIcnQY53
yCs/LYfbLG6PhHOpXlVu69vHkxV+zfEDClZFTM50eZAeH/vnkbyP/Q9ueudxxypE
cbVODiv0AEaqFpezfLBz3F3zNQPUCE6tAWwR1/nl2JKQcM/6y6cXXFCjWkkDTRrA
i9+GgES4J3Wc0BKFl4m1Rv7s5qGec235Xqcmn+A0tX5V5rFeakRkVvsYKtAEEZxg
KpuP8Mv9tSepxsNH+qInRWR4/lb3l6ZDCrpZsY3d9lKpNT19v09Y4M/37kRZUB37
WPvpgHtX2+L8Vo97J4ocnyNxKbxMMTs8DA7uY+i70fd/sovCJrKsFOomuOHJ/4np
K9CBUQBMTLb5vLj0EEhHDF9u8xqGNz9qtxQkgyZKLzv+W67C+hxby6w1ezTwriCX
bqY5H6Y1l/NjBWh+bJPvPQRw3Cb8oBHrRxIoTTkliDtSMnkNVg18wv27d0ijLZWN
7S95GKXuvKWkvmAcS8i1xjEBLUOwomVQ3bXUaFYlGZCSmeIvrPZVlvee8k8r5GFd
wKkyZZ5v2urIXmFSYmkxTc3eAFe/YSgLHZWYnfHBmVsF30H7309C5YhWZNDsu3rM
JwvFJRKPKBavlDp5pdRaqtj78/1NVrQXrwI5Hj/D/OzpPV3c1IX2vr7N5BZAXyKE
cmJ6rBYa/iX6ykftGWrurq7FB09OXScJzt74r2ghB1lqcvQV39QMeDGkNWXfnzrE
F3KYWSfayM6tyhbRWITpvbvM8H5xoXYZvyrwInJcC5bzRJq2apTLiB47WEs1RCNG
kibFby+UIyZeLhzWNiYMX7tfEMCzIzBjQeLtXtfCGyGTDewmHZhkODAecWMs64nm
g5QYnzhFdFfJCRrHsBDySr5vEB5TuWDPpz4PTENthiYQ+KBKzslpl1FetJIthERc
Wu8IWpJXODPDK/8dazjlZkJ7BA6xHIa9cK0xeavoGZKMF6JomzaLFb7JN+dG9tZm
Q5qn62yFOUd02HWAzx8AQONpElb3va9zs/5e9/iafYkaIItwkrV6DrZyDYIj2yPQ
TDJ11J4GMhDnQvBRWj6TRdWQ+zLbJLlwXTePma0SZXGH8VQeaNxDBadUd5saHFIz
/1n60qE4riOkGDzRkknCb77FeGEFHwcFq5v4ZS3nXlP8viUXlJOAi5rKw+OaIQau
orC5a8eTJu+sDii4skHfnSr2Xr3wG/YUbJIcUzsx+z/gPREfc+fOZUYTf5Mi4oLh
VhVXCltUd6yQcRaWP2glSisc+PV9OUHZzb1o+eO8BP5Iise6nOvwLlQ3G2QUFxpA
mjs2D0UFfuCRdadzXr9t1zUp+/w36lkin3AaFQ2xGCsh8Kx2DAzhjVWF48qHB1fc
LDruWjGQsby04C7cDqvDpXF7IIGhFpOWsdT2XLXy5XTgdZcKbgHRwrTKRXi14Kqh
wY0kEywnRxDxAM+t4L0iwldLZYfJiNG8K4awX877cQeGDNdE8tcjcKwwQ0qmA7Uw
3otnXbZ7cXSMwt96BsfntjrMlq3/qEqIIfVEjPbfVQ/pmPO75zWCD3UE+GLvQPgd
B7R2egOzGbw7jiEbZcEn1AzaPOhv6DCfwFnbpgfhnJ8BRA6N03R2HSjaWGdEC/KO
gsIMdkBenGL/Dfl/P2kNQYKjmNMFRbXkfg3exZ9O8DfRWZZYBqRAIFNj4vI95rM6
CJFej4fr097llbrDMPk27pzFsuAQcdVIdJgZJOZ8i5D+fkg8uLAtvHYDlHo5LBlj
CyVrJ27ZksPN90ItUbyR8CyvTH06FvHKvj4dwXUo20Qog2TTwvGsbwWP/CM3Vpg1
syjGiMv8k3Yp6mCnhGNswTtiF3j2hcDhDF+leIzHW8YJ9zqO0q4YkHeP9alYCT63
zNZuWCZ3lp5GJbR85ADH1l/Hy2f/0m7GU7PfpbsPUr2ZFZkf2luywisXpGhS6rXc
ixfLwH51S9R9oYwFDFlpaIJ6iwSptdB7gMFdahvclbP/li+0QrT+uVeMICahAZcW
yOesMVCiyUI+vwGkl0kNuU/v6EcP8tJFDVZe2ghHzGySCc1AumBhqDJdhXeJvBCU
jUa2iV9tdz6dJdUr0FTqIxKXtI5zbomHhvKDwpzzrw7PrvM3AZQXXgivABtry1E4
xIh6eNJguOkI6aEsIGBnvZBipxXgX7+P61S3I4kFMCV819aMZYZRuSmBLRRPCFVk
JPSKEiwnTOVBptmtLEtF1KRWTbvjr/Ys19xp0QStCiGuJb44CF1oAz9UZ7L008Ii
WCHPUz2ow4quKYsuO+YpFMJTXirs+Iil+loCO/kQtElQSl6n2upM2o4Gv7kzx9kI
qwifenSD1RVClXSpWKhO+Ir+dFBTdQLRQrI/9z/x0c1DaaMrOp7PcsWtKpcvEpzz
VnxPxCZDRxCySJe8Sf2sKyhcI40WzyzFY6E+x/y/FE984nSPDOCy/J+5+HkmrNud
dnc/rkW/yx7e/q9Ia+EOa8It+a5UsnMvCjKznqmYWbot7PDZgiYl5DhSxMUthyhM
nr9e8NItYtLClHkVOQ7P86nJInpucXD9Jgq9MPmIdPuTVtc2swCpMatFcFQKgbHL
X0sHC4XzAnTDT7unBJ/lLGcMLMAooCSmIa3eVu0t3yfdiXUwkUKTZRIByqYkYcZz
buXpwOjL/BmRIs0Tb3zWEledT1mM5sTDgBr2qtugGmpPXLHICtMHxRXTBWzKdITG
l8BlWBXPHlqaxiwmC2BjDeOTkladIR9qaSLWFvVQ6ah2uoEj4BZj5IjFvtv2oEVF
HF42NWOv1KangqPyWaS9L1ve8Pn1M6TaZBQGACxCKvVNlNMdHsL3vYpt/C2cI4Qi
GTT4k3MCRJJ9QaP8KMVgLgQAIsNjREPbjEqXZuIavoHGk7YA/bu71ohtYh7PCCDm
twyQGnD5ImlQiGXrJto4My8pTik065AyfOH2kKWIYjRyYvzsdfFnC8siGK/R4CvG
jthahCMno6lv6wmESSQk/F4wsXNdaWtoLs7gWYa3f4+LUGGvZQw6ev6OEfvAtwv8
MYliOhTQgj/2os+agI0SIZbrCNHKhfHLpAK0nOyvDc8199DI9K3pYdldGkTLLzk4
5T4PsInczlyLKw7AxFEs8KwEod3qiOXvBx+vp0rJFkih9hwJDTTRHxRMXDpUnHAf
Vch8e7pMYbcqXWjRsGE150QYzfijQwdymV6BrU8Ui3yD1aACNnSVZs8hvwN7blsG
fjP7iSry4xbPawa1ve6861999IV+7bJfR8YEXRoN5bsXgfHuZyVWFV15RZ+uxtXC
6OlhpIKA0CV1MNKW4hNFU2gWiwFPlg/BEVW+RllHbjWiuzwRyldmU/fseRpZEdv2
du6ZqE0HDh8rTwRHxcNmMZaolPyl9GJyl41aETEflxcJUi4xxnR92ROGrBHDLLHH
lcgHkOh3Gu6rzaeWAKbbZD2bfkpspTLrb9ow5gXgKzHPAoV0K1MijEji1lldR5wH
BXDBni0SwbmOQ1n8U+M11IrhZ214fBTtcat+HiTQ5zrms9FWXueA+X2ZVTprykiB
U2e42bRypDL0XnRMwKozbMDwNbNbPcpDyWNoMpj0SwYdJLl+dcqE4RYzVfS2XBmP
70Q2TXDF5VXfijbfyyI3aDFu2yET8v/QXY9jcUnK4R+jlDcSrJRhGD2HUDkfQA70
VeUtdbKkD4wiLQmp9cn/+caF0wiKmQhFu9+mYJA4lL6xRZpq2wkL3OSJV95SrtjB
NBTmxU5txUUvSN17kBODK2qRI1q8wVqbgj+cSjX0etTrX7+JHOx8akG5YEMJl1ue
7V+BTJ+tE8jdgNDRPSosKvGkTET98ZZ5JuGll5HR7Htb8Iaj/l8Cw5HcrtxCgTIC
F+o9QjBnCfnRY4qP+iTz5bZWfSpiKT1AXsWnXbtoXW78OTtk85mKQXEoDBruXLPb
HnJLApolccjmJcpELwqIRAXSsQG60cYaRUkHFfISgSGCaEYGe9OLZdvrZst8hpKX
sek0FeTF46gQZp9msWhyscxOoaPfBptUudg7GuKfZQYPfbYMBsmB3nMTmsnmrPK+
r820XuhzFOI7cbI05SChih9/IhhmQVPJ0XW+XRAe6MQAZQ+xWE8v/kDNpG5baHpl
YS4+bMVfrxzRGrAg9BIHiLFU84v/iBB4t6T9Jc/OJ/MBjOs/JEKtzb1dcekk2CYf
eS0yFQIqe7MhgZrONputb14VPC/faK4dMxWqT8mgHFDTG0fPIQw1xBuhdhknPGdK
Onq4klg0kqEfttw1gn9e8H9EaSSna4fjYU9AxeYywLqJ7n76EC0ELVZ+m/1Nv/hd
c2Oog+ofhu0AzorXYJDUUm39wAcoC5HvuBILpnCXUh0X0Ck8JstNAkTMexAtxEHc
FqWDfOBkGLlS4Zv+dDVTT0K1w98AciumHJocnM/GPov82U6orDvFBbiuTs7BWY9n
RO2+4W8BsObjcaMI52Cd8BSKptwkl4s4TxM11F4kEYmvUnF+y977Jqx2AP1LLiMh
bp2PDrWchBMT4T6S2clRdvGuVVYmh1TTdPpdUoarZESl+ghjvSdaAuBff3TfJBow
BvgEYwCD/bvcA8sbCeof9RikpYCpjOjxl10lleYdFjSD6RRe17u4l1r1/JsfvdC2
LuCBSENKrOEzWhlXFSHkM1NSWk8pVlyYmPcxEycshuntiFX3k/EPdRDrxSnZ5B6V
K7xdZRHs+w4fbKb+Xsntg7XWyKHZ4Xb3K84E94kk34k/eKcb37wMLdVm4wOmkMaa
P5WOxKrUM7jHNm7bq2x8Lrdoc8vAHL/vx+YakPvtml18iVJ0WO41xyiMrAfu8KyC
o0BtwyOQCxKQviyhvBgEtWdFgpNHmiMVLJmr0FFw5YWvoedkIasjqL4kauOwCITC
foxh3gO8UJce9Ez40GDmqeoQ1ErilBVf/sATchjQ8U1cCgtlQ/tIEorGmQUVYW71
wnd0X8doaZfI+H66s/Mqol49gqh1dJSHwMxXBNlYo/usB3zGR7hdpyNGARF2YatT
s9JX7IELnXrbc8WFqT7bVlvavnwQyYkOrEe1c+JM3cTJuTOSBfnkdMyyOMR1G6Vw
gprr47ACm5HZxwy7t4WHXRIs6a+C3Tc0Zr6+paqGu5ULziFxCy/HIlMm58qehCNt
pv5Y/J4WPozTHnJyOJNYmpobTpbg6Jotq9DtGi/Q7uy5PNV1RhOf16l6jMvvgFKa
GaqEDXDCBSvxvaNuC2eyvmE/YUwf6Pwi++osHle7N8qszbwWYKxT187Em+JfMxcx
P6hcei2DJPsKCmy1w5AJbckBJ8YjntlGUjQShgYWgji3fKCIfhyWrLyc3zCDQCev
d/S1F/UpB4H3yBDUATjZ1mbe7avIoeoC3YIZmBfsAlMQnNpWRFQ81xw/txWYU+m+
zMHe0t+6ENK6AjjFbPxdq7RcQ7eCm0XJTziAxfiJey8R0M32dvGeYf2WBNdHfOX0
3U+efSV348Eg4ylWQn2qkAAeJRU217+ZGP0nU+pq4HaZ+yPRdIrzGMNgqt+KE5zl
/hbqF32oQ4gHmJBHxStaJ+KA//RL79uaVhEJ3VIN2PCRtf8TvZ1jx1diSdB+G/3h
8Dcokuh6AfsQCS+4BUsFnA7wmGWx8BPqiVMeWeRvW0o1d4p3St8kH/0pEgWiB6sH
IlV+RBluOtUxraR/LoYfnV4nYSp2SrPTNEJ8UwjUOgxr0uEtabJIqzXETEmExMJ1
zugF4JR5khhvEVNHP9FhptGmSY/T2uE7BzRdiBVr+ihQgAMtSP2zERjkFjUo8I3w
IyC78H1lfbn/diviryAlsKtqNcS84XGA5BC7X5f6yLMcu0KqFsv3nEiE5TJ+lgq1
zCii7eOWUCofTQDzk6BOJ+yQ+Ttq1PZhRToTd3EWt6Ru8iG4HxyRYy5GMsd7B8hM
+dSErsq2iQ5TJx61A4OVskSv5crXgrZ7uKac5csCAlJRtqlbSzA5qYX6TwGitUox
CfiWARmhZ9xhZq2o0wsmrIj/vfn9V0fmJLsXz44OVx7xmz2CrzeHE4xDLPDe8fHa
rrqj4bk6OwZPV6TSqv4opPERYbpzJEnSF+DoU29YYXimTzgIuVYWXLs2pCqEGWiH
67lyrpww08LEAtOkpYO4XaG4pBKlMyZ4+5eup+TddLEgg585PIq0hwzZexm2tqLE
+zvmFlQ2T+kiersTwJkCNsAMuTiPDS20ZqeZCEMaZlY8bL59i+nTms9X7PSa5Hc8
dYrKi2PzBiM8CEGHVPZjSKQr1Jo91IDFxjRGvop+t+y9uxpx4EAoi6sWrB4T+ieU
ZUR119C99HZToLji5w6dKrCHaU5Tws4hCeFCYOqO5GjO022hfj/FAiqrnhtkmyUk
G7UcDttx0y/dp7SXmbV3GtBS8tHsNrDdMSCoV3DtL17gLNrFEk5Q+VTZkyci7CXX
TstBbWELyyjIOqD3MePzWxfpta4sapN1zkKjb0Ji4kUYtKbyz7coRuD8UNpwLTc6
dOVAh2BdzcxCzc4+c0T7YbuoejbXjPTgfLnvAkxXO+SFlC34SR3R0Ksiu3t6xsOV
ulJVnLz2cDm+wl8erqzIQ4sCDgNLShGwNOGhAGhWty4Tz71ouEIECtUaOCV7iVR5
SqrVBOKn2EuRT82FZ7ZD01VsaCz+hUXAlCPyvMDMnhGsqyTzUwoLbqFBn1nVPfvn
V1MYxplVZpmqcUojM3dIyRADarUPCJIGA5JAYlsWGYz6VSRRxB8wwv/debXqHtIQ
Q4FxaKeahxc5N5m6dvjwT0mKarvZPeMI9qVnxaoJnxEBKkfgu39H2u2rjjrujxsa
gBcZsHL2Hk1C3x9vkzgJ+eyBMkPVLodcoP+5sH93jmzDCUXprQJCD1H2egptnmOY
Dva5p5qC9TTl3SB+5W81bZc4yPXmsUz166PmdPpOnR8tQbpwQVbGbZPC1JakPi9T
H/wxlVihIsMDsYpfGlfkJ9cFTJSGYyBSkg/HIsvuWOp9yHL3wQ6rmFuCJUgWZmYZ
u+03xhHmwKhtgsE/yjmPTwAHdax3bU5G21ONgzqnv9j+4XYGF4LA7dVmDKlHDI8u
4WzP/TA/tb1PQ2LvBPXIcyPKIwwbajnXRWa5BVBKhXv317nY6RgIjaKyd/v+EzNy
MTsyHC4rMdCIKm4agONFZlHWAxLm+cIaOBKHbJ8cHTsR0LrTCHqSE34EPK/UIjiw
lCeo4wvr6NLnt8OJH8FgCNYcPlxw7P5ubdzKog/z5CoQSX4ZON2OXngtKf7+XPCj
8krTxqUDgIzNDWKQIc+fyaPy9qzccUM7qbA4kNQZjaSKW8m/NZJETVQ4JbyH91J8
t3ehi5vHzSRBleTeFjWKwRrGNOLmMvj9XzjU9MwzpzOPq2I6pjGAhSoo1sEgX2kK
G7utUZ01vR6FLh0N4WX9G4lKL9pYxTmaPnc50pJPDluEZ6SUUZxZAv/lw4X0Blax
4BFH7SrkqgrSL0x1aimP0alppcgI3cOfTdaYjzRigMU2d49Pn+za9RUPgMso8xy0
lrVhw5Jp7L1nTBMrL6PNzGTlkWw56kANo5aKNqTFbQN0fflaEiXNgIHMcbDtbssX
Rd3IAEp5WrvDkriAM9WQOpS6n5FQi8YCLxs/HRea4092xMTCEqdYBgaAjkL7qK9h
ARkk7NtFNgSPgBz7PoI/E98dUwBbUdYULgDdGIzJqS3dw4x79fDQpwO72JSfL5lz
5tl0p5n3gyYltqWhz9glteUQb7xs+zR18eA0m6XnXI8ab9icfi3X9dk+Ax+07Xcp
nqVwmEWspjMyCk3EYE7Ox9LidG5xdpZR5mqQXtYRa6RkhjGzU8PJnpRPJ2YBv+s3
Dfvq2SFxM17pb6a7j3wN9AItvh12HUsnRi+i6HAExc+mmx9guSo/TRPf8R9vh3H5
agAp+KIv3YdboQl8GIU3LgASdfmtYSZriGbNd5TTqSKeq4kqvqyYQ+ljXhE8jfp4
Ecu7LH1Rhsj6QFszuiCBmFyaBvyWqYJSiyB6iNDexx07JAKP1ZUbIi1MgSf9CajY
UfOn6HMmHiLDDYuDGd+4exozJmmFhc9JMmYqb5seYFS218P7ZBxckARw4s6gbs0k
2HsxeKekuo3JfZZ1XsbJJznLP0CnwQQi1WMdPPMubXng8aLQVSZZMFVbLMFW4f5/
VGXSuRSevNmy5tN0kiRaBUll34E/EKZOjsb/JxMhQX57hFbaciSltaJ2xxheq7DA
VJWj6s6zgcNC6sZ8ZtgGCME6AT5IlWLRNuulEPOX8qV1QevH/pRZh6EUJCdWPcJi
BA49YkjdyOKznj627vqsFQtSuaVAMl4qIS7jz4qon0sKw6p12Rb1oPkRbLFnaAzo
YYTF/N8ZTe3IaCxIZUwJOvEuwOgEXcgMJjCboZKRaVeL4tuRcnHxzjDIAq2uW6o7
1zFu4OBJ8Nwnvx8z3B2g1cohveFs8o/f7Sv980z35TRwmpNtjcyrGmDPtfleU3Xm
cj9YQzUapQldr/lb+Wq/mEh3ahb3oEhQDH320tqxgRpAbtzxUWdxxk8ZpGGjNSKc
c7FvOV+3BJQTtxmim7n8ZeAiy9+sHmjBK68/CFxe5L3YhhXW6Vcn2exu0CmJSpqy
odEjtmmCKE6dda58w7Y2IYTcJ+tbMNtE+8/kX5+HhEGPosPUgQKTdI7EwuADSlqm
0kHBxIN2rw1/28oUgiByRx1bnWRjWDcw04dOpn7bYKvWUcGFxjwY1GSRA7nlsmhw
H+PGRqyHCh39pKV2EmGA/CUTuY+SxrnSyOsGTnW//1QP0v7Dcku6mAMMCzk3fKZM
gUBb5mQi7nJ3MjKdcwHQKASnvmaVlM3HkMJB0QzVqZab/d4v6bQSG8jHqT/urlQu
P/ZuCYrdbjzffYrhjmdBPOP+jekkz5MixOPi+zZYT/8Chwz8dKl1LH5Z3sGydOUV
w9ZlBdqj3seYGWtbWL9BTHXrrjOAfYcHZIWsX9/Kb9xhPjUSGchtYaumlFV/0fSa
T8x5AWQ5L/xztBE5LBvpOy4HkGPouLkqpH5p3JE2hDSkHxgnWpqRsHvHfSEXMbLd
Rnh7MXgFDF+affMpy36qXGKB5ssdabhSb/rZs9cvytpIuaT/wiTpaWygFffG9GWr
bi9E8orkkjZZmKOH10MAu5LumkREC069warw9DrkKc/TR65sZdeJCL04AdMMqbRd
5uKpQe08RRs3eBS3wapfQKUgTVla+SIOq6KUAUgPwp9J3myVknPbB+aTFG2B3KCB
iUS/AsyCUoi0ZOMqKIv6cPGwqCzhX/ZyVKaA9MyepcEYnTk/GHONzIwkT8w65Cry
nGyNxHQc5A3KRyCzcg7WLj3iJatIHs6FY9u177Hm/xyPZAiOmrXjvH3KC9DO0evM
xd2i+C9/OLPtwUMTH5Nu91OkzH4ozehjEOU5jydWlQmMZVUM+itxfnm/mMUlK5jA
MBhBKw3Ob3U3IbWasAZdYh+7alJvKWTEC+RhNzOqYi78Kxop4aZ8Mqjx/Cx1M5IS
ZXGc5NACExGu+6aoafeG9NON9X/QJBmlvjpiNoPatoUwoFmbIjR9t8ji43UCOq+X
telJFTCqzfLR84d3sI6MDTfDu3KNy7/wS0WSgqjFWR7lTJr+FXEJElXQQ1rIhFqw
nuAC4MCj9hBuU6KrbjQucxEbV21u2zsRKB+0PQl3xD8lzR4vtCHJZ/Yj/IrENek2
oDeMm7Hc7p5zXsdT0g/yFtHLlZSLsXsZF0kdQBPXP+rMMZBH4L7t4/wNgfWIsbSm
bH3sASP4ETF0lp30BxcZkmuvSCAwzyaJ5iRynFF/oLAtzwycQSLOevho5v4AzV5i
x0O/7Kge7nj+fNWXMB1Q6odeAYEERbFWjffUWornRwo6vwE7/+CzELdi63K0JBKM
n4Q4RGHO6Z7k60Idck8xaQKFjJIeiP1OmYQG7Fc1hippgc8XLnbaXBAnS8cRLU6a
zqZDgnHeEKVf3bSjJTN6soaeacov25DYH+5b11QPpbSY2wjFpqC1V6f0D+4p6MCp
sFGpn2jaE6SLSy3cQA+eThh8D0rnHyvRk9XmnTrhv7F8YFMS6cnAPB14dad400bB
vvjgsWTq5L7dVAK05mRBU+RPSe7/rfOOacw7A6oBGkYn/5TCyeYdGYjQPSLGtcbo
LklEoiWzzlQ6DdrJI7/Rsi8SMtuXil5VnYJMqUQ3anJZH4RlpfLtaDuYnV/TLVvi
z1gwHXVFvKUgkffOfb2C6JMtqGn/s5kj5RF5GXr06ubzY6xmvBGV2A79MqKJZ2P1
nDVCy7pX+jIFljOAHV/TFekDVJ0fzvm5lo+5UC/rEyct50Xq0xmZew42o6u9Svqz
8did1qjg8fqwYMRyWU0UxpsPtjfLKM3IqFKiu0Tu6Cd6AjxB3KOm5Nx+xODPxDpN
LZFwViEhFvYRO8dEkroh+MC05AIpufzNrBPyvzl/bKhjVEAXC4c3mSd8HI9mTcNP
0tfOTeZzXAtnXoeB5ciJGhWUx9o4LNTPXqkZB+uKPoNB7kMquttEI25nfj7G3AQD
KbKp4Nj8M87JwhdhAiQ1JWK6FMEYRAgvf0Jl9wmklBRJKKkAVS8TGz6zbTNutUgI
5XnXasZvAnGcNgVpEGWiCod5tMtCus27XZsESnXb3YjDBlfs5rD1ej5ZyaYmRKsj
FJn+p6RfZBZZAKjDIPBxyP8rUhAJpv8R68kDlGMA2ALwwuZ4x+0JM4F798K3ncgI
wW27wviXEopKCUdBB85xtnDq0dhidpz055TWQ/iol0N6hyTUM1SwFBnRCGNt/+6H
yeRfLcZr/bayQURvT1QLZkyWYhzAEbgxrmkdSgx1lZciKQTzS8oQG9v9vcrT1Uus
lhx8DAPjj/7LY4EMLNhht2CCIBSundhuTEncMAR5S0Pmfab61RsxAXNXmjHMu/0c
Vha5w1izMqpI3aDAq6RuUpne2EV+ummGAfYAcl/DaaidKnYpyF9C1wvNJNfvM5Y5
OL+9mZ6el60XdRBWWE/OtDaWIlHdlM9jo0D/AmZ2iGJ94Y/sKPjyVt2syzltzVAb
3tLadH/dTdpmhj3YSwEQ2DfqwxUSB5/H37DQiCbaNg3xz3J4DQqcsxnT+wnMX6y1
uFAlgE4yHpX1qaedLnqxohr3VLCTIlluFjLsF/W6y/qmPUp96jRgh84/o2lIMeZT
At3Ez6k8FrgIbBQK0RR99YEOjKz/pbCahIOv1ZxCQr8TjCzztLZ8WWd9IIRjsCUL
NjBSfwnIsAOl22+vsKfOvttLP3ENZN4a4lkV/ymR78iJt7tCebhYGIj/tS1HCsNV
dOgGXn0BWTpgUovgDbWBRfz3RHwzuWMXN3dwUpjnw4p/jmc56yDQ+V5hLY4OKTDR
Ch9HddsYn+lTh9hEsyE/lwHGXimdPbOJIwRfJM1yiUnr+Rzj7p5uO0TG0pQS1cMt
mad6/PgwACJuS5pMI/fqNK0coMTkjB18QHjMDWmkO6GRss+045LtOtnbuTaaTsjs
mJESZd5lmGftxWlgdqQ5W5t1RZDxMBku3FofFtlqzBrPUZULrXu06b2pQ84Gu9wR
5aq3wHTD95dtm/k2xcu4LVUfO4TZqKceChNiLgYee1jhfLJ+6lV+peew09lbL33B
9bdlhbtQ4uuNY37LoY40FIz/eKqGT0vviOV4+JFm/3SFK6p7ym3eIw+FWI3h4d7C
L7bcLZZtNU0d8RAHf0KbQ/ms+WaERiVSZ/5KkQenaqWp9jmwliqhf+5cjZvln9dn
5d05+kZeA6TAjqtgfYTP+lJL0JweU8iGc/sZfuF3CkwNrF7QkUuCXBdc9N8dD1xX
N44Rfzuw/K6LmZe5yhzK7qjC2r4k6t8zuAaK38iXx5+9yWY/GaSMGQxADhR4QVeV
mL0RlEsFWlphL1lG99SYCJlrhzyD4mQTl/ff/QlaPzXaCe1d7exTlvt90mYvyl7C
XFq4xQSfitkVzWq+ZS1Oy8k+lvdRd4VJskSPby6w7laP39ODlc0SLXmBNXnt8F5W
Wu0A3tJ2VoZ3FJcIozuZVSnaUdood9TlW0Da1epf0fPkL9fdyoxrUzqgIP3CbhyF
zzqfQyy2DZAjUkkkO/BxxfR6AinpBf1uwxhH7gZAO6kK1aOk9w7BPaqUJ4hRkdfU
BVN6EIqPrQ3pQQ2rMclkkf1iqkz0qJLO8LSA045G6KDDBtiSmfbmSTwMFS4Lekke
FwW8Cs/0CDwuTU5xHPUQNg28l6N32cro4wNL+PDOAFKGESbrqBq/6OnGuxIazYAp
mBBrb/9u8ogYaZkONba7U4WcN99QtFsjumwBiV4X/gLgKendR8o0cCj2bHd5wKBB
ZX2AYopAKD7ZLQgvACn16ReINC3QlXu/bYLe0xEk69C+5Fat8g4dRe2iYDLa3yIv
yhESWEC/U3M4O7Y2MLNvHm0+Bztdy+pYmo+ncSrKa0RnJVsQ8WUFN1cDeyLsKl3Q
mDYuh7FrQAcq9bdj0v6FgdBFwaB4lIcmsu3sKMeltoxWhxwhLLCOFdK50mpuYqgR
6WeUgh3jbUsS9nbqjrjuLUhB5Qc5S0v4VP2z8Iqub4iyy+bdiIxg/0NzEY1G8Gzt
ABVQVTSFgzN7i47PD7RQ10cqvYIWlz2cJ2U32koFaDYAgrjhD0CrYKBa7hCt5UXH
bmLwF7L7lfHoRaal1ZvetVYPCBf23Okd98hlqcwe1dUVFz6nikATu9EoKbdq5owm
3u1sdczE0zGAx+aJ3qZV6SdekvaJdynDLywkeycm8Y9SKE1OKZOV01gDGkN8TkS7
a7AhadCG8lAaMEDSxln6sFAt6mbAzczH6H61D6+FxyZHCSIrrZTDDiWLr+cZdC7e
Qks4sruQ9ZMoriaj/rO2jY6M1XhOVvX46J8Poc2vJBty4HaYFHIESyg4pSOIknCN
yySP+7aAhjnhwpMTQJo52vw3Bv5m1t0Z8fg+s6CxsqrdE4g4SJbf9w9iwirwfY1v
gCijbaVXzSfhydS5h9MseDCaC1V1GGmaxQBNL3PL9Hm8Ird3By06HxNdu6ms00sN
JTIdBPgoDd+/ApfvxqGiK32YAekZe68gQFX1dB06csiupdR7bDr5HCeRx+6OYM/U
A5KxEs/jcZsGcjOul6vJz/uXBdWRZukYakVYFKjo2xjTTvw1jbxGHx8ErkL4LIMG
lVW9PpGZiAqlZ9KYMQ0enn8qGLpMYFGbUiyVTQsskssDeB8lqgnlAx3j5VXSrYFn
t6iEoP1pD0YkR8rB/41nL65KTZGoDC9ahWp1wg1+7LZdChDixDAa6Cmw/xDBZIWH
3ZgD5trt5JM/aDdMep3aLZtvT48vKIg6p+NnW8RuWTZ5AM0JRRahiJnkJY/efFyE
6RZjGhMJsGBpex8vVFOZP7HaSqRGN1myv/MUGsuWqNB8RC9yk+utvuPQ0OycyfVZ
vU4knGbKEtxi5Lk9Aw5/jsoqVwV5dJjkF38JZFFbxb5cPn3zdl1d9NGOxwoT4aLS
GhdgI/V3om1bL6mpdeWwuFvjuIBTozAgvA3WVX0ERkGxhL9nhLttT7EJhb4UIGI4
5/Ix2rQlvZuBqxiWC3r8kqNPEOrJXkgNMRHphxGvEfZuZMUL2/uYRg+GiE/4IX4v
oFPYMuwoGiK4Q/r3my5JGnm1t+T3iRHvJm+ww1lsZgYzWgc5Lm+H3W1z4B+crRkV
RQAiH1qkFPlXpBwMFwbYjD/oGpKzpKyaLZ3AQ2lm2+MUI2PlAmsZHZkxImWUar2F
l1h7VvUIr5mbBmj0OObbyd636oVEYT5O6frVFr5QutRMa8hX8rr0CUANCRyIboEk
7hVbS2dWoSMtZEdr0ZWOfvliIM5FpVXezHllziDfCAsPkacJrqw7kD7MQ3/+Qfcq
eslOiZ6aokjZ+A47j4k4A/q63cwWCvgL1XpRTnjiFBafnzrpZoEuPGEA+71k+DFj
pYv/PuX8+5dM9QDIjoMX7mJWnKMZK8Sokey22QDX2tWf4nd6Z5FLVBKixmMqkrF2
5ui/TuxQsLs3JJhKkmbGsQt/J9UfyDLG8wvgdZXTb+ExrTZfwkkDQWe/uYmqRkte
ks0+VVRCZF/bTz3v9wpuNck5qEaylktrodrmX8i13Ln0NzL3975paG+e7HBLB2C0
Inew8Tc0P7Oroq48ZT3ox8zJLiZeA/DQlMKpMWErscjqeCfz3OrwPe1bWNXlO55b
9q5JggbVYHbMtvfk+G8M0vrgHuH4+qoPcRPRW+4Izut3LiBUjDrdZ++6A0E9t+Ws
S7TWw53gwbUeGyYSLhc61Cx7wWIO7G7tGtS/ePhEjTux0au7QVLGaSLZ3Z9AJDDs
SMvCFAaVq59YprLwgR+EU8tc7LaFqBgbaXqbD+U20MYrxArTtl55p1tId4aof6vk
ePfs4bEnp3eIzX+uE6hD36J9zrfgZkyTs1YLF0VSzTsEY1WOwkYTwACmx9UVoRR8
L70RjIw2lGEHfLRcrPlgPSF+pd0nKCutEAu3errCjHFWjoy6mDUXwddcfqsPEbI9
TCHGgYZo98ocW44Z/oS3qWLgZ9f8d8xOngqxzCZ8pHO3W0IhW3lr/c1Cse5cAb9A
hy8dwPb78or7wHTH09YZ32XhmZ/7rYo+gasounsBMVoydH9ZijsjI1lgaNmBiVA5
Az48jDGu0Oxq9TTuzsbwAa3ApESRnyPk1iKukZls0Huv700Gj8cG6wE5vuvCWzwk
1RKlUGE/lD6cf5RHLOSxRnRep4XoUwUgwUgZOBC/x9Rele14Y7v2YqkoFhEpFsLf
KGaU9CIx67/j8NDPtx63mCkI7i7cqXsQWDcZ7lkQzuRnP1tc1TzBjs7nQAlIzoqD
wbD4SzXNneDkJWATyvSZbkEyFDBJRW1cAJDvPHwx/fxDbwKSZKJiLmdD/40s1Ymb
PvTDvSAibLo53XwAXFYFBj/zwOoqjkid5pxNqvSyPRf7F9bSAbnMSy2+/SsJZTFy
s1SiRaSYSfD5g7gtBgb2KuxJQPUD7I2gECASbNd2xwrwASo+l/ZRqlnSn6OKSYej
pJ8dEOnMCw0jUR+XIb2T4aUJU8yUDtB6whMvb9RUTqGFYiMJdOUWXP9oemmEdxXm
jL/IsfSmSzqgJ9hYlmB3biq4yI/2rfRC6fG27tibaCrkWfDAln7RReL2NfAf4o6U
eLqD8Uw3yETA/DqRTM5bzlHrhSSCO0yH9E3SQdOLDtWzYgt7Uk8JyHht+cG2azZm
cMsqGSvbx8oP6RpojD37M8fwMFezdSBHkmiaZDxhYAYJKu19tbm42T636GSbfaN8
OEHCvej508bx788nuGvLHX+bceaPcojsCehj7T/jgsWMg9w9ktoDtMw4Y0wqTrL8
2Gxh/pQXp8DWHkRfZ0ImytN4yFCM3MHh3g5MLI5mjnMAY28c7rFvfGZAZPiWIA4K
Cwj/mc3rTCaCJLzxGVFk/k64qbMx6nZ5T1AO2AJ01+8cMMr8ZwcFAk+V9jLI7r0F
+nIazEtv4KH6FfOV9yf8jOD6AcQZzeCQ7IwRuxcEwemoHa48LleNvsWr5FXASbu6
uQveetvotSp5CPbuBIunmKKvYeyZ/onw6fAGm4NYu6ad84GWhyd5E4h4+W76AAVp
hHRLyUja3xxEZS5pFNw7jmnERnJoKva1yFRFTy8KCrTcIKeQRUIFVe6XaaZsaH/v
PtqvX11KW3f8LXNgTCmlOy2Es+ETQw18DBo4gp/ltHzJ1sKrvutJUTOf7LQAml5m
UXBL2F7DgTC0NaUToGhhDyjwua7GJ9J2dYl1DxI8ZJvSEHyZZXivUbiRhui/gTH1
wUz3Uqt2pVWDohOaqQnuS5ET7/k+Jh57b07kQRIGqj/vWhkD7IR+e6Ig2kNo6aHL
uRaufb5cIerk6rWD0w+p2VUHCoOoc3+9WPkDyeLMhnzOVYxvQTgaT6a4e42fWVRG
zTK8VjONfvR5hjUwkhFwpRKnykKCTT8rIzuViCxZfNvlH+IndNiAiiJy2M6IMKRS
FcYoZp3PE5md5dwKObH9bGCt1sN39nJjDWVlPDLmB96VhtENDY9s2xbpaKlWJg8L
PuZ2wWrjyIaXzI8RNPuE1fp5R9IXSTEQgc7nw9hxnTUA78MMslzE3dCDTKoumA65
S/X6kn0MFCJO3IoyYwzFNBiFO4hZZnwiFzF5wXZkhp1yBssCLNpEM6kZryQEMi/C
KRVhSK23KQBLrhcYtDghVh53dvGchJcAebeBxgyH5BpEpzgBtjIvAhlxiVcPLi+e
bU4Ef9CmHARK2W7DRohV27BFrHKPvqM4kt9mFcmRkrAR0DPloUsg+/wwDUVAxkrz
hEM28+LNnm3i28GDh2u4TUIM1IRAZUXDMV4SARoX5W4Lgc4VO11AQKpYzB+Hly+p
I2LXGZ6CnnTgJzufNqTXvywn/eCS35H/AIBV9InjTRGp036Wu0wLZ9nQe5iRkQZP
SYe+Znmiv281mzmmZwobKhJ/PUTOzl+OLI0xkPyYyyKopi1OuLWbSpKjb4RDXA+h
tLBZTgVa93N9GFRVoeo2Uu1mNbGG9XaOhxDaDI+ITEpGwGOlPQ18SyOkh8NUeHkU
E53i75jb1GxvumhPbiME93SEsec6pHTtvFR1ujqAazPBTbdnXIwZdZOz6y4hrv8n
TL7mK9As+F7m4akemKCY6VcsFWr+ToPqE59SY+hogNFyD/LKHz9wpbyY0AcaoUkV
DfxJOf25rqLJSmrpQDaGE/Gbk2UF88gLJl3IDMHpCEJVSgPjnb2yltjR+LgxALTz
YMOpDXgRmR2Tw27TRcZuiCSzQr6gbH8ebDVMaC9tZu4sHkaMlrDbLeix/1OvXhCV
NxoYDXLGNtG4t3UvPE1i6JrxDu5uAO3D1hKqtbJnvtJRuPkM5T/VTxZWk3Bb34tf
ZWb8rF9lPvK93T5DcYlN5xdnJ9n1HVFamaA76LT4TI4AV/BQRiyUD6N24/G1YQ5T
h1Pov28dC5xLmuiQp0xQT7FV93kwEgxNJ+o8tbkmH0qdFPEvxIx/xKmulnOUxTJq
3OW7OG6ub1vhLAZHceSSiPJliSKBB5rHfCjwm3eeSzpY2Xu1/oGVFjNfDMloal/Y
bZuqfF8DsK6loy3ff/LRKewv7FPux6q9qOJm08I3foYVpfbZQuytDOa6dt6Ylrul
iy/z8b288bOXY2k9DEYyv32SFof0JpXKxzWoRt5bpxdEusgTl9JfMgUsaKid1IDV
9V17XAWCdb2G9Orkr+dpMS0zhxKpu8E+qHf4HMJEFOTSV0brvtW9MkEo1M4xfck5
IcDgILJngSmWqMljVpKtA0kg9nKg6RdhPXEcSJls3OcD+5uD+YAjjneGDVz2R3ub
JoE+VaSfmKYRjcCfcLOJfm8bOsgEHkNX8sbCJCq4RLlFTaTvsqXNGzaMogNXJB9s
XQz1R2PerXiHNcPXHWK5v5PKYsp0wJ6cX9hRoATlAwatLdqctUA31DISuSlM0Ids
2ozx2/s0rrAYeZKBHcg2ZPyo5gu4XSaQjm4h8U7t8RCbwOmIV/dsUtaC0CLv7xRW
PFT6F2soE2OOWVJARn844TtidaeLVBKk8iY9Wr3E2aRyqFptE3oHuq//weBXbdAC
Vt6ruDEIMnzo8mcCOkolFUzJSJY2/5+sJI6CZv2JgjYFa4M7BBQ0Z0DIOdRdokzR
lNxXaOOxB7JNJLvFnfq/L+/izZsEGZOcBsLXL5dni+s58QgDiU6/bRFRkM3jsrqn
aZUV/MFBEw7UbJoQr/P+/FYq9hPKuwIct819OXmmMssdNbN7OG9+8azL8ae86nM0
2DH2fXTTN5rj+kZCUVf/wib6/xqEnzWxxSuQTCItu9AjUvWeCN8StztKYZCaS5dX
zlII1hEgq1mjtINFulKgefce1Y9JxjL4uCspIl9B0JVrO2IA24+ygUx/blNeHO6t
bmPGNA0UVh9AjB/PG/ub/X/WsI2K+DBLtzkFDaNGa+za/F65T6CAfbgUCZPoaFI1
Yk1zi82Uwqu47Kozd9RqflVR6HfPNAGTq2eV18UtvTWjSsI+dGqzzscn+9tjaTI5
E1Aa37EtUDwf+X5kaeWTX63YE4dcHaJhLbn5Th3TUxKxdN/8EssAMLUkePQzJTy1
ULJI0mZ6kfgESY7yCGdJR4lxPW6I0ecqTkHAEeip7xhVHi7Sp6YDTNeiNtl1KONc
Kyt0PuBP2FsQtxHp0UmwGw96LU2bpOUYPKGBbEjIHmjyBqvq6bUj35e/DdOtZ/jp
8wgZw3h3badP+273YMMMs/6t5H/SMLF6J+NnEkp1cOTtZsVsFxbZV0iw1NrxasJ6
phi4e3vxQ1S4hrslN5zqg7HWS6lybjOjv/+xalOLULFKDHJnM8uGjsgwhw9A6qwO
huayjHAPgXH3H+rGwtg6J43ZP5izOXzcuKUyqxjL05wowJ4YeU4pMkOhigIQMe6u
hFPbVP7dOvPHTQR2hrgdUQ887G0dBvtuGKQ3XhQL/rBX5gbADECyVQnGoRZ3OvH2
zF0eXp/5x8LokBVjeKj8xijDykR+ms43WDx03jI8uYJiNVQ0qVzR4yDupuwrXp71
RHj8EeXMZ6zTD35sRe4FQdkcgK78QOTKe/8qjxMeJxGTE6SBgN3P60oN8qycWCEs
U/vaNFxOSAHAqE6TwXP4/CuyQ2HVkZhDf/+o63ozWRTWRBvJV41hIVISxiGRY5GS
55PzG6a3VzJBmT6u6cQmYRjF9JnSqp6PKRv/HUIsKlOHx4o7jm6RJWhkvwuPt7Aq
J7i1eaRWziTXSTkW2fH/vYkZ9o/pxsL6/FF2f1lAU6qabNzzZq/cNnD0/Aorg1Sf
lJGu8S1aVtemNeJ/aH26EtsPV62+5CMaLh/988ihDUea48pBud2NXMgoK9q823/M
EeAJzjjbrdJWiq7umw8biLy3C9e11aWrlzUm+zHIyfDKRvZLnJad30Nfq1rbJm/W
FmoBnNodRw7H3tZ2+qoFwOEw8ZtaJtyRpBR+MHaJ+z1KaI7p34+P7y3sABYK5v1n
fXeGn+o2C/arXv8+jKXF0t16as84TsrniFssNdn2UK967ysc8HZWHPxEhk+AiF8l
vTmdBt12fx1YLYn4AJ4n/g1H9KOmGSVcN1Z46ce9LW3N2+HFxIpsktrLpo0ox4g8
hNvVl4JuJTHXy8JzDe7fbqM1BeZY02oenHV36Hiayni96iicafTqPAqXO1WM5D2z
9APgsPTfYojJyFFbMg/NmvHjFdfX9IL4q0+fBsrkXgMih5BVsapqzCxmPKCyZ5Pf
St3kvtHWyCDWeiLkpCRLmZYm/cTyh36N+6J3C4wtv5xr2pdUQwy7OmJsKgSYB9ci
LSmIbcGY6UnWIYl1OuR06iMS2vofAwufcPYxQVXWLH9cPiToiYQ5lEiV6f2WYZ4I
+XHJ5AIajTHOBVcYE6ywawROg/NfAAz+SR/ZBCHEm97z9XNlvKCeaDOLSsRX1GxZ
EDLRwzFtywEQVUe3Vj2P2wgkziliC8snKZanoDzy5IZoqxUhZwyeCoDsfldzJMGm
osDVevVjksZTiwktR1ehRrNzcJrPDZvH82UrpGIu6eLSUFgSi6nAJTriEsOVNjMm
PQRjvQuXMkBAVsV6mq1z3XlfSgon6/R6o0Gb5bBcjFSwBoxYlfd1oPVi+whazEfu
6HrWD9RxAfeMycn9HT4kOzxQrI6vv/8H5WY3sLTamqesDipsjNz/xbjZaTB7o8yj
retIvYhctkZ5lphe3okNdnyFYSPU+erXeP/NXerzeQJnZUWwMKh9IzurEY337CnX
FDEoqLTP1w4ESp9p0ARloV8+s9rt9s/WMt3J0TKXBatvmrQ7xKo/RpTVq/kmycv/
myDRNk++q1YRqyVjcwJ4TQ+G7BajGk7WVLS7opxfelPiB/K8VwEslVfBjtTu9VGU
7RH5ILOySRd9QiAcKO5kFpkSQ8tu2W0hdmfd4bYIqzU0aiz+c6fRabjVblO/Aq6N
DGflDiqq/2gNSvU8V16XCUr0pUo+VzNjwuDmk+xO2smi0cRSZFHHxrfr80j4Nm0C
Uy5ZeEkvBJEh1GY+R+YiDSTzrZA3q0+gHxs0K1bOcw+poMhQ6IGoHrBP1QbTeFd5
k5FSlZgzZorJMhu4cFKxOtiY3SvApHbYDbyo9X+rl3Gl0XfN6yPw6UklEI4TGRn0
nokxGiXmcBw4DC9mj2rORRyx+2c1rm2EW+isKNJH3AWctZUZumyaEgLVJPDI0LDJ
KQKyYWoAcw6b6UbzJpMpFzzl1E99DpXkoOUQBrIaL9jQg2Vc9tmeicWicP4K8Lo/
mwPeNPqiE4bqJyErgMeNlRdej6ryUr7T7PRHTamBf+1b2eH0zABC/ISdJxVSXziO
0fet8L9qQ4BdnxQULczXhT/wzKioCTl7OAUaIkeFZ5Ub3Y6W/re+b6rgE+05QO0q
1W8xGk03eiPjZKM9N3VAO+y/MGXate4ndDW9GFng4xky6wETMKbyzYws1YOccLDL
H4eJSO/6uKe4F2rwcNWcfsbOsRb5V9DmfNBGIUvMrRG0mnp9gAOFg/qnSetwqo7m
ywMVNstC4GbcIaYkJHh4JSHH7qb8vF/cR0Ik50OzijEAaUIOAJg5kJ3cLODxrtwj
CV5te88ZnRFUL1yuw1shXp5e9B/TA94Dps112vQJGZZ9MrNKLOWTilLqCtFgNjGD
VHPfy2TALc3bpZhyVSnr3QgrLTahIqYttSq0g3Tsf4Y2Berc6ipzBICSuDp1uRS2
WVUBFkBx0+nw2Cxd63zSWvfbwC8bqsuFojavJuzlOtREMEYTQclCLv0J95yEVdbo
FzTXu9LcU/k/mfG60s+H3N7v2cEyIk/6iiQrI/w7HFQtdMb0CflMKcwo+xApGyfp
lRBqafqRrn90aFUVeGcQ/N1p5vtse+cpaUQHQHLUwjoPMdRc8k7KhI1/0sEysATB
goIbwQJzcdi1AICpNsb5M8IuemW3thL9/OlURN/vfXq+GPTQpzxWSo8nhOeZO9fG
Nq2onYxhatkGFKfmcP++zMDSS9RpQ4PQheuV++uTlHkE9F+Q3qNlSRbu3+Qvr+KN
08ZM7zsDg6j84jVsL89s44u46mCXG0zxmzuYt68WbF6CeV2jw/EJQpHlZiQqEFoi
aR+2hhpfCR8PJy2ZQ98ywOYhYHTkLvPSxQE2KdlvJu/N0heHKoiiEOJIwKhkBHIt
rpzDu+31n3KDeLqIUm26db6MCerHLGck2SiGyxzW1PY/7kfx4C+Vg6zu1Lprj2Yz
pjd5Pz6I7biBtNEy+Xb3tsK1bS+ym/cyVcHIQvXRvaCwLKGqTJGkUV3CB2Zlprpd
j+wMvh9LPjKeDVubQV8BzgMY94Mhngy/af/o/pVyETcnRq86uhbuBZCyOXpm0dq3
HBzPe2AADj2Y/TxRd/aPWz9YPboEZjY4KOxwjTEvNorh/7kIilTwAU22SwUtwSJQ
Z7+V+1eB7OwCMMlTNwNVY1AY3+J8Z6kDV+NXWtIehCbj5Cs1fJKSnGxu1mdLmUe1
1Kk0kStGEwc39mAEtpzV3/sW/4vYMnA5r6Hy1Nmb3ZeK8Zix4iB6l53tpzUz8xJz
tH5gZfgpJeSrcMXU9P9zD4BN2i7Qn23eHgibb2WxMrK8kubKKgeEY+jB2XbB9cyL
rWGXCH7AL0ECUDneL4uVXC+uTTC+YNm2r0lOsOoYjKJqB39w6VDNWkYQBkgF/Awc
/MZngp0AvmTaCRF18iyieDQkh992Anv319cLPviqNjNKDTOGDHY/dPUowY7ZbL3L
p4ZZu79N4akw5IarxfZiT7LDl3vUd/RrjqSEzh7hRw+1s9d91gsop9WW34gcNSTc
AKXmGJd4Ukan1l3GQKnBYV+bR3W0WIx0CIURbglsBhEC+GWtRlOTgpsfKmYzeBl0
6HAXmupdPkGrneCYNsgPdp8AOcceDvKNKr2MIQsaRZx09S6InkrmqBWD2drOwZK1
Omw3bye9AaLROMr/RrO1cqrLv6K5CEzkyvJ5/LaSOG7f76Koh+zFPDj99gj3/rVU
+ptIbT0j6NmTbsQP54bGLgwnh/+rmjfJGBXVfGonKBGGnjWmMhy+OKcDSSZ51QEX
6bUeAzo7HTSBiUE4BdIFBGU0YIt3lDrmpfCXAmiIh0w3lo8zQt22nFjwyzPu1zgn
1WSFOAomJRR96vjqyYAGAx6tM8jp5tgME3V43jumpZWQlZlAwM7imLz1hTabxlji
w5f/loZoYfe5hDTEug49RPE1jBOKyvO1JXHAJ/7p2mKvhk9GsCFDFlcnr2kpnQYs
zVZ7nxkFpTvEbXXkDyLi0lzu/qp5Nwakj8QCbCdmhC/P2mRO+YfhOHHqwIPQO8Hd
wjUMeWxIS5nyGVp+ikpizuZfNVH/3mjZtO9/aXHdTqC4A5Bn5bpd27z5eUcn+2Ee
GnE4n9MlGrfbhCCnTBcn5kExPSZRqwRmwDOq+57GLUVO7vM1g9UzfUHDnbtaZyN4
dXJfyHGVveXhAF19w1dTA3a+2+vjIo3F5gM7C/peaD0LTSG0FOpinpb9N2skGXaC
rlpd0T59kGCcaploPdurtMi60jmpb3WSOA+oJ0hsceC6/Q3EPkLziW2FbNQE4lHa
HXc0SdAzx6rv08dAsvt/3PvGWzQVoAg3C6MsBmso3CgUGkcku22LDMus/UTE3cK2
cx9vOUt8sotJCBOszqYHbGc4Q3P2Iz85nMKwL1l4D1xo7OPz/eR0zOZ187D+yfyI
S/V2+/2Un6aaN8zLgIQxQ761UOb/3801Hi1Utj33Ma4qf7QFUNdqe0x5g+BJGXeS
s646p/g9wVjnUVRn7syG5TYeuy2+FxGaH69lmiUs96lVKsDcVjwzfrYXYyaD0JWR
9sD0VAtaMOa/M3kQl1dvyFFESnedSYstzKM2T032iSl67YqxdaAsbYMDO9DP+W+g
/nCg0sbrbCFPEzci6YxTnb7BzOgLOLIEW368dp2X8d5bgddMZJdf4TC9kjEJbNtW
kg3pEGcQQkIsbQJSjx5kCOPy2qLe4H+bTpoEUtDAlncj3XdeJ0muQCPVmaLMn2gv
+uRMrwq+YYAvt2nr5bix+8+Xx8GJs+fGEg3OV8vwVWNhCu45TP7uvxEywz8NrVH9
2WvhGsByh+VoIm6VcJyeTvscANvB6n7MNsHmRS3x89om4S0kxzIUB1v20EtM5DQV
pwjMJMenWEsZfn7vyxala21ccGAyuwgawO4UgeMAyyNB9fakXtnb19vfZuyThJhd
/1KlIzZra0qR+KhkTaGxing63WL+vt43+HWLeP1Ry0MXzTAB8U9xpMajWbu/n2ac
WJjjo2ifwNmJyZ3VOsRIuWDE4G9Jrz5DSaA3bNCR4N6Orc27D4z7OMOTeg0973wa
YGmlCGx95SJypXxLEwU9tROOU/YMMmBkrYdy5Wtg70mNBnaBmFF39TeC18UeGNzY
YhdXUAeZyxN6mx3RLw4fIhqUi5YSp1D0SAfZVSeVJt926Lm+m5IL4S77B/DccVZ/
fgxsJ1PezMTvRq2p7pTFEoz37VTE5nnT47aA6xEc2g6F5Q4e6UOaW8VJuZ4nKwUq
v5QotAkmBSQTy9VtoEml+oYlk3uB2a9sOY1dsASkAnudlZiHLUMGdl+mkfb9Tj20
1v+QHLEo8sOvubhVIOeEyqKSUjnQkudQJoNhrF1b7pJywbg6V/HDERXq3GJgp6Ep
g2EZz8rANbGyLGncBDYD6VwlRpGiuuaA/ygt+5zUhuvdRdDzr4hKB3QGNjJIrXs+
FVZOXs41LCVAvZAHxbFo6tSHnq6CAmZBFYAl+SFF5C6yBUf8u9vFghEabQBzNhem
3HYVCLZr9Yk7PywjjDB4jybMIPpF9A/9TcdbnY2q0zAC5WyAQsMBtJEvvhHpT9C/
LDnv4U9T3JYNzTaXX+6B/pjV0ZKzjjWczTJEnpzLlj/EGF+ypH2/6hghkBUvbzCG
Ksz3HG9JkFkM07vaysLSvSoNhsSPj1rtG5G+/oG33L2jwKTOnVg1Ie8ytzrw+CjL
Jgn71ss5kTSxT8zcHFJKb8gzeD9nEvzBMNZHL9YrX8M5SAlVqbTH/j0r0LJvQOau
h26PzfoHSKO+xwdIOM8KrASAImNcd4G9CyqDShxhUQFOqtE1Rx8Sb3YZ3nnYFyDu
yaFMQWVWBYqJNgilL7lk+8/UsnCUt5H1HDBtgIGV6jDxBkuNEZoYzBhW46QGlnt7
Tq+9b0B1nl8FnbZpDsxVvZ2+kMQ8fa+hj5efWOQkHBOmdh/2tDTVuL3xUFaKy+1C
FjqcOuVQ6rDd89k8Ju0aiF+L3GSGY5TtD0rGo5IA+DUKycfboLnW5qPaCjShCPdN
Yv0wANtWD41vgAVrAoMDTMejp4ty3wS5Ewz8LduwwHgq86DahIKhv+Cu88cecB+j
5BuuOW5W0Hyw8j/IQO8+TbsoUM0bwMgC85lU8PrxPpknHfeEJEOZcC/6oCG/xl4h
T1lVARZt0D7dRRvTCmAOjecjkP9PCp9yGROo1ThscSxBGEh6NggXu0VhXWp5nQR0
M9jgGfAJiDcg7C5AtSvI6iJwlvBB/T9NpQZP1DaQZKRR8BT/5CDVeywXiqx+Jn5J
QOrPn+LuPKnJh2M0LwOk03gwxlxt+TpMJDGHn0chABMl53r52kOD7cAhhE8GCyzy
dGKYgInxxcUXvAcD48VwltnYiHgRCvCxPbTw8AAYkSwq0HGf43lH6kRWEv9Ojvul
RV2bwH3WqXJfZnKWMm4//QBFf/4YqO7EZUuKOouhSqgDxP+ZZKcaXXJ26KwaTqEZ
sOR9JkpAhS1m/y9iaDeazqhemkxPSckmnZpiWR3ugIhDYdUfALXvO0l7JCqX/9/B
Fy5Q/6IYhh+fvEAUJCVeAUz5SXF+qfjHNZqPYFmhKoCEemOLrlcKQtQMG/a/pOH9
yejOWKz+dt6RuljYdjjbcK7+6MRTkcvu5hDO3jguDUJOh6bmy+BiTr6oWAlZ7S2S
Ozs2/qjfnkJaerzt3512QMuY4R1QnhyGgtg0y0X1/dstigjSOY9/+ArVIX7zX7W9
TTM1hjPxe7R9O3CZFO9K5nBDp5IyktKHD+XvJXnbdappPaaF3LizK2QLqtQkONeR
OQWyJQ4ByJwOpKeQ1nKQpnfWH8R13VkU4eV3PWxWnxJB18xSLQVrWIkXqsEmhVbw
QHg19QE+FEseDqrwrsLdYM8IO9j405V1TIAqQBwj6QwbZ7PiOJikqk6GUh+t5yUd
ocB/8LNT5cbBVPXIWgNnXnkdGbJBfCNEx04G/2l71+EkeBv23WjiNVp7B93JCKAz
TRBV3/FDZ3Uf0jFVaL8E4Df/ZEhd7cT8+3SHthYRjK+MAH4KaQ2RmneoT+LRNG3s
sQzbeDwFL585Oob9YDsDJuPp327b8PLq0BWmwPVgnJodTRyjDicN2GCc/WmKCEh1
5ymAmFLMWshmtVZIR/xdVt9qasU9al0GIjqItyZfKjel8DldoXjdyWvx4CjamSuc
WcyNRYJGmJpWQ41akq0Aey8qdRnDTXDb/wLzmP2wmCJ9unU2YislVa2FGJVqi74X
Jmxh+itJEGVOxiEd+eM6F8KN37cnW9Go8CPSN9Wq32wkT47tt5/3d8av9vgap5bB
gF52zGbe2X9lu3AVGiYvyVGjQZDUOR+HAxFrLsBo+yNBdyOG1Z/LowesDP/R1vmG
xryH+jIxuSDxndy2q3/UdWLnYo+F6/12YlssoxXSgY0CvOLz1lmdldrE4fr2zbj9
O82IYd3bZ0XDJYe2+QGtiTRuBud5lRymALp11XaCnXaIDCSVSSPiqPyQWyLUIQaK
kkmFuBg0r1QLxE1sKB7J+I1izgmt1mNIEbX+a5Mayd23DzDV7uHIPEc4ww2WatRk
1wB+CYaAxygy/QuQMjqgDHqCv+DTK/0mnjYJ9EforEOPTZmxzfu2IzfCfiAG64aZ
fGB46FVnqEe0tAtKiYpQAvWWy9qDKQKJP10PFXrrelPMGlbuokonOsWvZhmUJ5Am
lRES+KYrFqIZO1nLs0x85xvIVRmf03TaNo2PYJgJ/PcQKARczSVCZrwAnpaXedwO
5ho5OxgQ1QPkG/C5ND2QbwGmA6SYmxWT1RliAqLmA6eGrvuY5LeCWIFfC30eNxsn
Kld7bq1RSjfPOYgYmlW9WrYE1qeF6SrrvCHrSD/BA4tk8cimEPmaxRXTIgl488BG
munnRTLzzMRhS3xvHK5xAvvP2+pQGDWnU6EiyaoR2h58su0f95kCxenI0vtcviq2
pvqbDQaoerzWTxp2qGVdpoHGQSOQ7vvVUviME5+Iry/qWjpcbqlZHe9gY8IrAjmN
gmOYBkrQboyQ31DkTIeREWz2nj0WfezqPK1bkqRcAAPX8YQR+7RhS7QZzb+t/XpV
WdU+QJuayvqacz8iP5qEIlCv9aNSEyTyw4Ndz5IX7lYYTrkPDO6MIANEkQkPTTQX
u0ykhqXar1MyQExW3lsPtSDE4kstgM16X28XNQRfzx7BP09qNgZyULFs9Hmmv8LD
4taqjpppoNcMAxtMfW/jdL9r3joiJHty/xGzpXsxJkWR+/UeeHvaLZxV5BmBLIQU
V9qI2pHOYZb8zFyS2VBEJW1nHww8pUtrtLHEKb5Vwbb8HYNdyl8lOAf+n9aIvSF7
bySBBDt8oQRtEwdOdp2v5c0hzZViF60oS/fjDG0eyODrylYtYI/+nn4w7jvc0P6s
5GqCtZrubUCqNN0/buofI2Hdo9YUauxk5ggVYHFKh2yZKSUPKeOA/HE+OrtP45pb
1d9oy4zKfA1coIKK3TkxEZr3BQ2LGg6NVb1SRX9LxGW05oQwoJyg7HQU7TbX/i1p
qYToePpxIhO25Lym2e40Y6PA/hi+4wrSsTJqhIdfmjFi8d95/g19dwB7Y8fovf7q
9pzzAF/5JDBoyy4dS1Ic3J8SdsJ9OfuQ1yriytYJEg+sZAQsbJ1CE/DBlzjBXNDb
J4L+PFbbA390+FMdzHmgZk741mIi4Wgy7QqF9SCY3oRakphc4Kz/ITMX7xPbSu05
aiRqcl6P0nGJ8LYiMengtJgWpmrAmhefvQmdY+/erTiFlAAXPyl2l44UtYLw0wzp
guBBtu9SCL57hSjIM2kiaQ775XrK/c258t88WhPf7gcr5uIXi2OhE9Po+xc8QjgT
LboAYKRMhZ0EaCSofOHnBf6vJC/rv5QWabslNS7YpSPdlLAmZHzbREu7BkANcPkI
+VUaLtCylN6dV57RI/qhcHdPs9cRm41GfG7LYoanfB9fKv4dqP9EtwMyTWdgJite
GcHaXjE9JCUCRUSPgmTqWBpMDx5QAE9fA2giMs0xOLZjxBQDdc8WzqiE3lMfu557
4pO5W3IJruKJ9HFEVS+dfGrl4idlioUa+UKBwlw/+PWUjkRn7cNQUT3lGp8R3/+z
NzeOw3UJnQ9lzIwDKVU8F/+nIaiRgLdqdLIAFN65aCoymnyKi2dRbCd/nEGl5PVM
h77LO7NzuWEIWhb1KSBKHV+RXONxvdb19VDA+3HDRf27QADf7qj6sh8sfCu0BTr2
6quL9uKpyy0+tx+M7IHDuxmkPoIBEbdGnrU7Atq03APP5l9ZiuY1dp5vAtDmuUQM
tmkUCWQZ8zzxo/ee8R1AwVBmFuvEJsyQtmYAXAt6KmV5crY7kROXQvBwfp+x9m1k
jIffSWq0mYTkqIbAdYalci3RcKEZTMKIzQZdjz7ZRyc4R62SRx5VlFIbT5yh2o/p
bX/OBDgphJmO/l7KRjkh0rjiiyP81+wpARqt/0bWHnHaJuLb4wmCbQXcFsobHEx+
lcDfFDmRIKMB5VSkBjo+XU/rN9a+FywDngJlW/mdnuH0gny4PJvo2cN/LQfSJb0J
+HtzVvSM5ynTgITnOni2Dr+eXCEiw3yV9h0rI4d47P2x2ShkJ9ZrU7sXlD/muQLW
/OU+eeIGHKCb1HF2mSUL/k1wkOn0L4QBnI7/Qgfp0hRPdDT1UWJp5SShk6o2yoo+
E0XR6LmPzoTAwzyKrzFTs+w1fR+MK5N5LT0vwosxyDAbRteMk1p7qlU7pbDXWApK
cAPPM4+lrfrkv6DpU1bDT558hjIwI3LOVaqibvShoIRAP4cl/VHbeQDHJHairJM0
Fh3bO8OSxHhm2XCh0JzdZqTvQriiHH72JghOmaoVWjRniCFXFSrwR7IJS2ATn89Y
vHoagXervklCJBcyYfVbzn0fQhAlpufTqryQKApPpVCmlVJH7kKtUSjmK8wiRXSK
bIyTzhyV4BJRmGgsIaM4tW9GXVlbMBn7r03O21duo9dtIwHQDs/iRRzatb0LOuiB
cOmYEnMEoF6Yu9Dpgf2UhJ6EmoZMurTOJTRT3hJYQQso+FW+gx8fKoJV5Sc3NzdP
MMbdk/g9uZ5VUs9yZirCBhPUCqGsZTbigBIC6/ZO7QBmZWEICUCoKiZjLl29zZXB
LVK4w7E6cBie+bXmKmQWH2H0kPsCKpIRV/mX8TrgoxndX//WBf3JAuwgyZ21MCo1
Ssp9Mpx01e/bax00c4NJo4y3qPy0bX/zTidP8dAeQfG269hEnz7TKHWmCSL2NuI0
bNezdIT/DG7JV06aWTX1OcodEed42Z/Zol52o7VjoubbdtwGJaYdJkYRTsGlUF9n
WtGpCGWkSwuNvs5xlqH1pws1qoptlTjQR+dS7FeWXd6Aw7oopghm0I9dMKoeA090
kOXEw49qnuBNLoDvCz2Rbd1LrgEaIH1TRPehusbeaYu7iscJjzTVdpH/H7yOpj04
ucu//OuAPYJeIOdpg8L1uFP5j43x+BuW1EmKasDlBlU358gb5KVadY6kq3wBUH9H
P5rKwxtvetHd5kLoAbeN3PA+nd8awh3x9neHCvVixAWlZ/zr0UMxyXB/O9LKwW3J
TdG7A7UDAuGzdt+PWBbKEVD37DjgXg6yjmuQA/HCb4rUfdE1TXnYu1lMkB2qDl41
qsbsxXvQ1n8PvTz8W3goYzlBFwRbDz0UTmuO+nH2M/Whv9O1N6UrkgQMnu6qX6wV
LyZiU8aaM40t9ql6hEIt5zelzvpV6DjZO5jRLlNv4/5x7OofR2Q5t3iliX7wbCm6
Fk4yDAW4Yr4FkLqiJp9mp6W3rPx8CI+ZwrBj+Zdn2dwzUapJMsU+qlynRbuGVxMW
nXLvxNRbAjIztdk1lOvciTvjfwg2Zx0pa9En0yg2+OJAb3BTgtCNppG7bgu329Lg
dkxgXcaPF16elEGmVKb4kEwY+jXoOpW4DbbSpdgUH96yBW9K6R8xuji1cRZqJxP9
i9z1tZ4CsdpKu9pB2eu7E07BPtwo2z/Hnt+60TZRWPJhg0MFpEtd33NHrtLbaw46
3kVtXiEAdgAG5OkWijcwqz7mwFDUF0pwt6FErkvSRBjY7cYWXmCMbPcCQ/7imO0f
8iKMz/Nc6SHahghG2iLMzobSX5jVtC365BhOTM0kNlG3ZXv36ss3Uom+pKYjPHdm
3rW9Ac3g9F7giXUcxyRUypfjMs7YgJ3AMuaD1sc+vEuWGgCTtJRgxmqCBX104Uyj
d61A/48fhx4duYFD2McAGbuHfGEmrBdtlejUUb9broepKVpVBCawLv1wTaZF5C7x
ohkMZeCgtCCNya52yW37os6IYipdDBBJyZLku0c15doYB9mdyoN7ms+N/TDIXbTP
232BlAim3XCOFmagvP5sD/QQLg1ZclRUhCwwWnJgPqJuXt4LFqyik3j2zpltgFFZ
hzoDSq6wPSDnDDx7oKB2cuMc4+acipLSM5ruGwcFCD5Qj39kfbk0gvJKoV8MZQaZ
dOqhPmDNHNOJYQ0LnbTuXMt6ABI63AL6YxgfbsCuyu6a4w9kkQc4QPHo9asx8K2D
/hrJwyflEIokYk48cG5YiF3dheRBwPQzG0G3hxrtvZ4tphp3XDSxzh/B1VDfEh0W
H4SkgBReYNZbVjJFq+9CrQAQCiND4xA1IsI3AJmBVnxgCtcCXr2tNKLV4B0v2d+t
8Dgf8pcihL9IwrP18fnHoLPV4LqOSd8FXPwRqZQZsyI9mrKTbdsRqTxBNSp3cRf1
CXUZ1zgng7dHZdqxa5J7GGROiKW6xc6UmxKdDPN+cjtcFgcsd1mbUKpAbl6uSEC1
2TlO/qL4hHhkO/mZ7u3+8qT5jDqSgEufJsyvc4+6pZcO3cv/5+1mH9iLzVuVjrig
ipzdfUeNj9NjtY5xMEiHMsnHogD1f/4j6wBM72+zA3MYXXTi+MPPctBgYLROJuUX
N/KslDG1KeJnmDE4tJk9lVnwOk/fMmdl2ZcV0/6R+qYJ1TbFzK/Eubuk/9OZ27yL
/JH7BY6tz9hJ4kP/SZUpbfp9nydgehSw1YEdco04mZUkTD9ZYkwZXq/xnBlZC8Bk
aI4QGO1jYiumnQc98odsOho088GM8C9PjkdLAipXv/xbtWyijq6ldVUduV1ysxzs
+7sM3qEZMpRx20YrZfc/JUWZ1/jvrn/pvRifXkv+vnO7+BgS+6/TnVhZmkzA18jF
tApmZEdFoAlw1M4YNgncrGOTJoGy76n9UKxn+729tk2b0T/LhYgQdoT3lHf18bBS
5aa80bwDPJSnKkmpHF7vBFxjNFxgNQt+lMiIdxCXpoYdIGFin+kci3m+vvPcF86f
jpcpu7S8l6JAC8TyRBAT0/AmIwFJ2Y4LJ408JAIGLcn9u1CKaZ5BKGzLF/5X+W5/
lo6Lyiqy96MBO72vebBn5qhdLnY+yXAADYMUBoLEB7/z+MxtiY9U4kdYlK/nWhMZ
2ZSF1ZJXIn/IePhAYTysHfFYFTEJ1Io3Ft4853IcFegqgJ3qiRIodUksoBJT63J6
6haH+dg/wjPFH1C4gdTLG9eEKAJz8IwPH2MC+kI6SV+41mN43XPRJNhUWU538zdz
/8jodw1qGTbnMN2av+P38ISbo4VEeuebBzia5nQ+6xlAgyGY6cu8+pVkwiGK27eR
CCVxhw3Vg1EwmdaUa9X0dr6/7UmbLCFw+EzxJzLKHQYh5Ke+QXkigLVXxfHFfdza
4geULLP5Lkx+pKjo90sbfafz2CpqJWhzmUBO2Z+XoaLUKlgaC/KrbU+0S/UMu0Vl
IVrLv+U7XgpGJyhIezSNAFEu8SvCsyexJEz/YtM+MGHS19xbb5ipvTxLYgsSKScY
ka3r/8a2foVZD1L91J3p7QbzgylvGN4X7hUkaWERldsypm7dkRdJ+eF2RU6dhF9m
ZTjL939hAVsQVQmD/KEVNjJhHwwY2Kqa6YTkVW2zQJGSP1QjPvrBQarieXb5N5sq
SPlJmKKyJP+l7LCsf16MG+CvaSVd+1jOsr5/btraS0Mb5kGSwVSKOiv8m0viSqBN
eRmbBJ/SCoZrXJ44Q9RJR4yPPBNYorYl1SgjQCL24hLosJqI8cxVZPgRfKnCm9H2
l7U6p/J3LLMv0lC4ogyvu3xeXeBUt63mtziR2OpruSoEvTmrWoxOy8fg7K7HCq2d
DyChXy7ssaPb9HFSi10a2eKsgKXYW5K7eVPiGPMkn8O064ZNqJMIncvh6mBH2dU2
NrvQTCISTpCgar77rg1Czj+TXPld1xCFlOvOnx7IECVfkGWSzNX18nrHoYTzAAry
7nGkakaJWjEOunxDqSOYgi5EWZBEnceYpTQ/q2603qVqRnNZqxlg46Cb/Af+GmZy
FIzAs6WGNDmkm0CNahDoiD/Dm4wc1xbQl4HH1SN7TxlS1H0kpv01fc8+2uuJKqBV
SDLexZnrEZ4phlP3UPovxywi1KymtdVmPIpcoLQON5UNavoVKSxUlgU5v6Q0h0PL
L2qYvUjusZfCrjuDd5FLSW0BKLg+yK4XEqWLCiKuDMKDVC1zrIjCQNziAvsn3yb+
MS9bxw5WDNRqVv0jEe83y29hgX0M8xNpFLXm5wkj6HeKpHvijyjGQUAzrRb04wjV
h7o/hmTjy6af84ik5ytEvX+G3oZJ6axyG+NJJtf7d8NKNIQMpvFvLTRxWMXh2Pbg
bH6I/+PGWWTfc3dH6GL376r4XdGZvY5NoFs6rwTT55zjesrUgHE1eoNTlqyXF62H
VDA5Umz/z2XSUfbIwFM+SMv0jq3tkfyhLHwUt0ILsUxrGChp6tqZQuLyb3oK/+5Q
3495E6wbi8tX1R9GfB5i84RQT1M87zxWFShu6y2r++y7v3/wgYHoVQzWCT/Rv6Gm
fMhEm7Ge2hf9/mM8GTqr8qQw5WTKhrvJbzCp+itN4vqXSrEG0tKQnAjMmNY6Znx2
IWcpsgEvFOhLh64JSNBnZp/kckFjJA7GbXHiZwIBu2ReZArXU/YqFmWgMSL18Qhx
b59qOFCj0yQg6RDgAd2zeOxYCg6xw6a7fVoULu6ex7gU157CrglQhpX91/klAVfY
xUnXMjMspeip3NKCuWATpfpwcyggNV1uJLTEw/AixUOD5zUnu5G0dJITJFMKmuUo
PR0zpcBRyuU7ru6sEU0qfX/V+StsVx6dI0GEOC+48WKzBDI3sQb4qvanbig6EfWp
Wqtqna6Fc5Fc0J5m9bHUry3cOUqBZDI9f8x9aPbrQUHPAe8pRD+vEyxj2XjRTXIY
BteTuMtRm3JtaI8dapHQHcIVYeTfVi+QJyk+amyaOjZrbQ8S20c931mswH5hU2xA
/GfGUf+6++fVcv6hjyh5XxCE2r9Ivvk/kLDFlTK4V4ipcm6p44FeQ/DNERWYS4yr
nlp7YhRu9+2CbFiZnkk81+eN0/bW/nyN7vnwHI7qBHXpS6RKZsFNpL0186jB201D
0HrPzHTS/uHCiSytI7vuswe8Fi6rZYpyJv+P+FelJRcYgIkzih6Sh9DPX0Vh39uq
FsVE1JBx1ZBLFCNtjjzxU2GUTMyKtZ/gVIBHFPh63ITeBi/OYNQ11nrHTV6y7xGw
mUhghzxGkE+QIoFhlQrbqxzOap4f6xqkqhgKs56CC2NRQbiTzQOg0ktABTrWkImY
V8EIZUWB6nOyDTeLDobn3AYX4h8uOo5XrwLATsnfDLK7K0ZSUdMC/mVeN4o62pdg
uQliElek1dGuFt3QjHTxih4qxewsCAaeo37XjfU9rsE0TkWCnmC/THOqhChgOayD
ywAX4eLUabg+RJFUgT9BA+TSRYVCDzJ92fPqlH4eVszba0SBMHIWuEgQ5Ytf9ni4
9tZXXnDPyiV/s1Paszo6roy8WrL4k3YhzCogiD8jTWbjy/zn7L7POILLKcHKoPM4
ki/eO5zli08Aq1LDdomdq3oqpBu56yN1GbMa177dUNZbIAYMepVkjsZO5cRblIjD
OTBJovAqER8eSGnvHP6bfotiXnpknV23arWkk3J/GA+xy+G0MnsCrxI7ISMqZcFq
nNWbeN0cwEsaSzG0+lM6t8B/oB5wZ5ndwBidsfJr9fdr95IIswyrFrCMUsNCiTcM
VS40h/xUywXABhmIdSRhKEnoBKGkW120OdcBIjH0P8tNzJBmvfoSX/xEqS5E+PHk
it5QlmSx+BmA+6CapTtEedASfeq2qYkbtafZXF6aMX9R3dG5o6o6s7waiZ75ujbm
p+6+1As3NvgMB7B1aeFlq5E1+K98YBGRC8ZRRX5YR/3UR+Jt9af1/1MPyN/ZCb6a
VogIJJUT2ayCpaRUnGOUvSHZ7d35oZjPFnZLxZTZAXoBaypDyY1VD018mElOcxw+
rljASb0Bm36DpnPo1AOEJUsiswIAa8LEglAXaMn7raQ9SXK76KV3YFlJpUgT1oVD
YMndnZnZhZHL2TO3fO65UgXkQ6yvby6hSn4jaxOU+MWB1QxAN7XDA/QxpJyDVK2Y
3hFw8yBG8YNNbo/rSmWcGE4NHxzmzma0UWKyMtUqzkzHLvREv0WPoOhqYZ8FHNAS
B2VoTBnNDb4kPSuqUElZG0ZkOHiSdCI7PyHWWk3k8rLJHDAcK3FVHIUYy0xPmVnK
N/quAcXMXmoo09pnVWorcQ/cdFTzzBBtsCFswoZiC6uiOB5NiWxvlGCXuMaeFoNP
yE2SCDk/U4KMi1kP2bU6RdWSyPepKfzGPvdvuR/oPVDjmGU2jaBjDk9oLdlYgqlM
NqwQzVcfvCnS6tff4rlzV8rnBg6Ba3Iv/UrvbxOTVOlxj7xDDEfm6tjg4Mn41b0H
ZiCNSwvVsQjmhfnl3EhKx/Ts87vOlFN/n8tchae+42RXxGV5JINlfDP7S6aGNN7S
kcDAlJ/fbnee5VXj8BGADeJRkXwL6BPcRfa2qz1k/IKfi91EPjFF1wkMQvJbSr0Q
fJ/AiuhqOnojsvB7tYUx7ItmxONtLcz9zlREH09yeRWcADT4Hlu8Tt2qowcK/QP6
htzN82tuQMIcEZv2B+1p/y516QmDlDElF0swPFy7Nq/ltP6gDMz6MlbvhDcF6YK/
wTSgfP+fZFo6wYxEqvPpayO27psu9P8aIZnpVAzDN1VzGT/faasT9i0eZQIQtNt1
kN3l+y+zywiAMPwcDtBpFcEJZCHfKDHwPw9rpqpziH9Cgb57fB1otD6mgfHYWUmE
vkd9UbMhiZvfpIPgi2XJodQTCYVN6sv3ZMf7FCsd8Yfs0KwZt2H1AmUmDZfrG2Si
CMqSCD69hH4XGRv7Ckqr9f64Q3M9Biwk0ZqHS8meu+Cm47OyL4OUhJZjY3Ai7wuc
wMGB3TOzukKIbDERI5UAFmkiloAWuYl264lSNJEFzhYdn0vjzMiX8cqJii+GUyvc
Cdnv5c9JO97WYeNMxb8XX1CfQeMWL/LbXyVKQNRiHAFBoVMHwuvs+WNloXTYUtyY
Ier05/SZmzU8Bss+PQ1sHtCay61xiwwETraD2gTxVmPnQ7InRXAEsfEAxbc+JWQC
oousiY16uQwbGrkOdzetbC8hApBZoOf6fdKEmmsMeMlRxEY1IVI2d9Z9IXDIxk0w
9xu4SRrEh9RaisElgmZkXFu2kzc03MMmbIQPXHpoqP8xGEekyvYaHbM8OgHNCF+d
ySTSJiaa25MN+waARpT9txeQGVZ7KuF1cR+vDwkCqljLbLHFbHyPS9BbH+jM+P6D
Oynfrhk59GbjZl1r8ZPDHodYsuhmsYM74ODUwMqNCRAPXwCLJgSWi3P74r3OfxA9
66IY9u8+hjvx+8Axz/AszB2NoCbzZsTNIZ92Y4lWEYd54U4EdohSCMcGekt9iOf7
TsJZwBa9/y2x4wVGmSdgnfUoX8EzNpKgSKf5yzEIOHcDN7atJR3AiabffEmXi3/1
ssKGxroJAEoDt8Y7j9/q7iJPKt+fw5B8/f3LYyRhpkEHs9QLosZ6nP74m4xgPvb3
z7+YxXYtXu09RMUAHkVPENlc3Yhgil1d1oUrHUphuBsrRw5kQmfCYkj96/zYWt13
ulLZykfjpKeMgUZWczlr8KHRFWyXnjmX7hs2Lh/7EHCWE8K4jRQ/frUUopYgk/ce
2sBODahPoEcOkqD8hohF1f23xDIlN9IA8srWIdpRqiXB6kbP9fKGZ8TSlotU719N
QxYHdwqXPyLqsxldrM3jo7k3qy3xo/6owRZDjkXSSSqW2E1jaTgFA7v1/0u/xG2q
59vRAvZIbQd4w+dzQeXMA+i4c8smIEA9RjKBdYWzjlboavsmI+jH1L8zsv6S536y
Wpk5yh3Cc9JaFHDaG/pXVpL6QUbd3PMvtZ2YP0JT4/bnjjPY1AiYP6uiPioJ/NJK
LJyTqAXk1WRg/n37oyaaqyVjvEQWhNEY/mr7cfpFxef9B3Q7vLbGF4eAXOGgqrUF
4K7LekjL17JskU2rwaSYp4mWUWC8c5iGgxbCxgq6wKwXXI5CXQUZAOYiqaLyBksk
EGQiai5e/WKVWA5fk295dqFjF9MPyPtroFR8l44xCIcVVSKTZmar9r6Pl7yAEw7R
g4/DLnht6GKvSNWF/HjpTgpC+dQK/JqOQ6mer33e9ZyOmI0BNypciCEsOLmNM1EI
ABbCQTxeyISuH2go3Etn0cSUfc3qTdWDEniVPVyHes9xM/MA/iZpTNmsv1Ck/ioR
3NlgIGAwaltaNHKurVS7SlULAYjO8RRe4LjIf1BQOEZXD64woeeoaB1CPktUFoKr
3Ai6ekQJHKJr+miiapzNCy4uvpHI3XCgY6FK8UEh+oC7a846YK+2UFQVMu2LRzrd
AWEPDS/CgTzmDssrTMNOus9JuZhbZffSm6C2slSG97X0bhq4tqAH/QnAcUFhHpkA
yY/nrcm5hYH3Dy7qavIETg92AzWhsM6tOJG7297miy9ehlrsgR+hkcnW04DiXjAt
JD6fxlXhuOpHiyLV22M5yKZsZ+/a7VJv9m5LiXf8IF1efAdRRpE52OXy9Wk+wz/2
2nm9fQoWGcYgqyVacZkhBlDDwDuymAzg89Unvz+Z27ruSIWattvP65FeFg9k+4ws
bTSTZH/CJsJdZIjdIXJ7lbuQssRagcxnMR3MERtWWtg8nT2zRpoSc7qsBGgvxTiO
gzihvYnZPcCpzuYAIxccYvYyZtglzp+3OOuZUBDlD+Vi7p9lcxA18sDLLftFGWMO
V0f56m3NTlNXE+eNXtjAAHWVdWi1y/Hj22iSObZqGVSkcWvw2GnqLmV4v7vGol3l
YsoNcQY9oTHprDlvzmcwnIPwF2U3aKMg4qvlbSgSaregu+fBf7E3WezFfWohFToc
KRcE86z6IdrcfuH3BtiywLbRoctyJYzSxVrGKcbMJHYSna5/omYMk3L84ZBYt0gR
x3bYWXW75BVJgSomSPmp7IKo6iIwzTJUEoJXla3BP4rw4/DEpN7AeTRgCqYRfUL+
nowm4z2dN0uP0SsBpae/xCnJuJtwfj7tb/ofbjjGmT4lYDbvPEOwyRpwHjA0tptu
TELjHb3xFIxXKYhSa3aDd2pSPq348jK6ZGmKRx1zHyE4IHJDK1ZY0Ej9xIc3/yt4
fmWaUYQFoKpZSQeFDYFOQX8WcefMVkp4eZPrWVVmmPsZM2covZNNWsE1kxOmp9pA
bigH1FwpprJvsM0nZwxJmJUKtomS4vwQZnzrkZ8qr59Xe6pQ8BIgoanSk7gOJqPb
Tdl93Z2tAbAuWU9reGUagvvvs7CAwx3r6L2/MQUsYWlul9QOeqaqtm+hUjSw3Bvd
1RedV53NPehyJxtcvC5n2qMczH7y/u/T28wNdqYvzkcDGOXNa3X0zEbFCWZQ/Sao
BqzOyKsA1baR4fMlfmEiEV1ZuBjwUqy5bGqV6FiCnTN7kJGw9b6k4Mp1PxIcZYLi
2GmPfmEb+PGArVQ76azY290AjhHgc8+BMANIaz7gX9QWuQnS8JPlAEyZhPaAsSl7
8GnERVoBnZVlsiJcsEl7S0PeOQioz6iLf75XwonbZ8GFjdvD6jYQVNseqOxv0vpk
90X3sll2G3xXGCCHQm1Z9Bt5CqXKhc4jNxKw+RWdsq59/HXE2zblwS5SlEfgJGSt
AOi0ewqbljPMCiVQY9LTu4xTzQ7EH2CXmEj79pn+jVOeYGMwWMQ7jzP0IMKLKC9v
5qv/+Nu5+NI0MF5WbF8nr3faqIlkMse/96OjuoLUC4KXd3S68451l2nHhY0Ai3Yg
GK+O+vMqEklgsxLrmdb+sBdwlFtZcSoMOgW5MH2uhv+JyrB/fRt42qGckJiJPOlO
jABia4NhumEtfNcEWv6Z2z3bKQqY5wn8lDhXv+UziNfYfJgCn5+CF1l6fPV1YLlR
IKD2q903MJvhXC00E85fGHlP39oeGWCo0Fr7A4euDpOVzRI4+ISjNSN+MO56Q8dH
GVyj9QCcdUcSmDP9d0mra0QZ2cEm0KGijhtgrv9OcNjhbMIYKcBVtKWt+2EqSqYH
lPQ81B5H5UOo//VsZbza3SNYufifYq0JyuZz16BUwrI9kFkcWjqSrPU3pbgVO9O/
QYtbMrhzU6DHAgUtlNqmzsvPsUZUYwfkrXCAaYMM5S0AZAt5VX3MM1kWiccQCjs7
T2uvcoLVxrNQtBttyzJnChnUWq+FzjaynQaeZRNanI5SPZyF5rMM06j3WQrbhvRl
fRxNzr60GGJFp1txfBLwnB9O0WcYUTBnnVUjCXHyV2epXiwshcHmiu2eZXiHK3IA
2CFVWVmFEL7gYmiGfrbpZO/jXKeVBtgK+kTGISZ3eusgDyaNXhsBiUybR+4Ap//V
Pt6I/IdXPpvwAmFispRGnwIP5kvAFqTgK3mobgBVWps5+O+ABmhOJhL9NVDIg0fO
mD9PaXNK0ROhyIrOnvCHUDGYUSBeJg4K94eS/hNr8Xs8+5npF2rEatPzfB418DT9
2wyj74meJ0KqEyRXE92a1xeDmEBQVtylbzwohnHb6aliG+n+tuBJzz2YW5YFlRtZ
qiqSTvC1teXRkW39ZIOMQ9FaMOHQcMwBb2RRV95vXdEK6xjamzOSawM2eRQXATAc
o1Xs1+X9tMxSpmGzoDMlN6At2XWFgLYMXgHhkYLHyC5VW3H2Tz7xBd+Yu3vBwxJd
CUnItNRRX2m2E8hHYONjesqc7SKnC/LHD1j93fVEMttF4prSK8t9FZqJdQqLCmW3
lLOx73R9GnepSCSnAoHEVvfDGMxaCCmJ7mi6F+wclcSm65z2a3A9l1VqDL4c1M8j
9lvx4GsmWVet3ajLQVSeMvsEyfpqGDoaaF+XKZ4kY/Qh2KWm498WGDvI0kcjU8qR
r2ECjXD/x4pYvXtFkZozlhbFlKBjCIgi/KXkzJCglcg/C4WyR8IrOCsBjYT770o7
aWlX8LMb2J7zuAKBqzEX4AGDfoNFki1kDTc/NuEn/5PWuVN8UnX6c99POpkkRWJv
Q106I5LhvupKLaLb8V2lUtkEvTuq9ldWGKEA6BYI/Ncjsy+JZ/j4NKycgBuIVDP6
f1qSyevWGzYzU0wgJKFWYuknGyO3XfbB8V7HLR2ovCWJAbc/N8gTk0dgmkzpH62H
f7CBONgYI3WzH2OpKmYsxyw2CWSXXsUY0ogGNRcIiv1f90Zd0DRi/kfoXmy9JSZo
hIxwy1MqocNV8YRron51xH12vDEcim+spiADyWriA4n5kEYNpT+jZe0XYUFCY6wI
QTGamVXAj29rHjhT3S8NT44aORK2LCSK2/fF6gLJP9Mr/JTQsAXDuqJ+6HZj+mv/
+c38uZPvU0LoO+05gvlfniHzI4LQJys0jztH948JBrDvf4zwa337CNgXn9kkZNBY
Ey69N2lxmOu1BgbmPAwJXQoMIiWc+iF0Piz2lR0acwjePSqlmIauomHgkLuAsg31
AKSbzLA3O1B1w4QOIrid5fQR79SCJMKmUiZ7tIzZjnGsPFNtXGLyk/cw2EYmYpxj
1EAB25kLTEy8Lq/OD059mnND4UaUCZzw69+PTfsGHfk2F909yILsBnlU2tPWY8Ug
/21ZLUzFe6vxgPtxMp6pEHNQ2z4+iTZvqVoLU2x0IW9vzfG6QnfrndYQuUJwPvEl
6AIJ0wNloTwmPq4Lbgpmuj6N1gYwiLhlF3edDjzcDJyX6FSXRYl5V3HKQ2QKxeGw
clz7V17Y5JdCYp3VXp9NYadSkST8Ap0T2rYDAYQz9dL5rOg6LQPuehyuv65ZrieY
EEtr1bnBU0hwefOg8s1KFgWAJ1rVi9bcYvMs1EM1Nt2MEBZu+02k6FW2yWQBdZlp
5jNzdrnmGcUV1HeDCFI+JOtPMTI/b5vfqidGdMC8V7HxttliLFGWl0JdAdbr02Cd
uDpYF4lKSnayCOIM1l7mTYTK0RLQu9VqFbTPkWDM9byIokgR7ps3LZKX57nF0IpH
HisbNYLUqCm0tGgd8H95H60VefLM4+OcPvCyuQ23xZ/q67Vw345+hX/6J9i8sdeh
W9k7mHSqgV50ROFmNCYu4jt1k1tWve+pPp0KaBv5KaYXGcrMjjEGDrM1snKDIjOG
iqsXReWPquiaA3RIDJdEPcAgpQeAmMqWjJsPA99AMzRMidJsMlcSMRaGAiIKcqSH
o1RIHMqKuHrTJsndRyToA2b0eVqdTZsreQ7XW9CQQSLBvI0S/X1XOn2aVhyQK+bA
oZDXjVPJoFVhH8yf5dT3VmC7CxP4PxXlkRj8WOqtWac5kTV71pz1wZ4SBIktnFHJ
yUSAQkSibTGn27wrd53dYmkq8hyI8QZ2UVC9ATrhupHMLZmViq0c9lTlWOYLd9Ee
4jRkqORnASLGKq8gB8d0nwSUlIG621WOC9cRmC06GH4mIS6+whJJr9bHowAOA1WM
iEVNXw++ztdKUl9MTFQHGR5RLtoY4lN5HVut3TN1r7xnS1K0gB3CxB7Pwbd170cu
wV3LEkZrsz6ZsvC0UmZjMh6SBoDmwj2WeNqDcXU1NdaKsfBU347XwUFiJa4TPEus
X/7w+TR/vtViB6P2o530Zvk1ro1z6UVzNG8RCH2IMnuJnFwLmtV/8hoCG0Riu5ae
Qn2UYB5bPYPnJRBNXW6tHtAnwxwJe4gNxLD002bSN1f6XkrmHj2JLe+KyXYNxUxR
NZAb8x5VkbNESyRqqzUjrmD29PamaaJ1Q24kUGWEJ4zdTfLt1OqjjMX7M9Ntj/N5
tuvHxkCXzw/dXO/da6Wf/pPwQykctG6f/Hpb2zPy9MJ1ffwaM0lU6UoMe3btCx+Y
WWPOeitiKYhWZLlQ+SAR9RaSSdzO/n22TNim8G46SygN0ucBrLJPvSsjT9bY+x2H
OuijfBPf9iPJAki7JrIOZRjVxBVEcOny/ftP5j9xCM59Z/YokN7OPnBlPeaj4Lvf
nOVEy+NZKg38BGJK1PddfDhog01Y4UMLxYsl+F/rzu8XnzDZlpnpZ0b2ZiZLZ90f
GONF4MdlcxD0T8bwwZcyv/Dd9nEDK9OOWlYastOGncYOR4HGea4keQ2bYZhxSyQ3
alhj9mjC0WS5APg4HeSkHEOeJ/BAFf3gX+g6xbc44k71d2wHTHo4cK6wyGXyCqg0
lJj3Wh+XrJXuZVMdLxj1jR9nYnRTs/9ry6cmbEZFvdhgvP/06hLMvxybyJuPrOiQ
ts0hh+3CPnMbg3RHEkjSuonigc7n+Jhids8UHns7iDflE2beEaTnouO17Phhmox3
U+FN5IAw2fX5JO0mnyGLd+MxIuL986yXvCbJiWcR/3Af8utaMuzqCGj5Fs9XzOl6
LyjFZ3dL+YHzh2bEqvEzSP4LfAc0OEWCsPtVD72BOqIY9l8QbPoxzWWZQBt7Fheh
J2wEQMvbcG03vfLAq3xGrndBkJs/OsonFWm0iihI3HnrtU29RdjpjJcuy3aEZjqS
d4lmnyY9myQTl0Jzg8J/DZrCRDKSrJoLQOfWQxggBUjTFAPspTt7tBvooOFozzwx
YdSxLjwgp1+xVc28Zh9NrnY+xEMDHXT+v1vadiUFw2pnUIGKQ0V4c/k433T7vDVB
4mzBPJaQjV45TDZ4RQRmRl9xJIC7HqG6lONJci4vSOsTrOy60wTyDcBDoVKO2cv5
nKDoEHIYZ1B0BGoVhiasZBnIHV6WcEWKiSa4O0LlPxmkI0UfVTy9Kn7QbJ0twp+l
KIzjaFvGapUgA8A0wdiGhE4IsXJMGURUtnCGyXNZaiZUPS0TRq1g1kvsjfBE3N7m
bDktOlapwsscDsokac8xxlyyLcMFYVcLljqbiGTo/xV0BJtINzciW8FAc7nsh6ec
PVP2T3Ede4nX4ihozaW8MMAaFMY7jAuML2fIlZCGC5STchfTi1tANzHCui61Pp47
YlMf8ZPTBB1e+6AxcoIlgVr43Ilvk9PVjB8amONPdf42QaCZB0rZudHDmjGkzJFw
VcWr2O9W9jdec1o51s3zzlLXHGBO42Nu9Ju/6g1bS8yJJS4kghxmoloasZE3kh1F
7h8DfWnLbO9ZKP5ozIld8buGTgEf9T+QyVwImphrMu0DcV32nZqsiQERw/23REZD
oFmF7Ao33z0Jx1/YDPBWIrJdzhc9z6FZJ4hvQaueCq5Cs5n7QIhngDPjOZil9PWq
fhx7Ym+cGzrbnwiGdqacR1Kn31RWCuPOZHheHYKpfV+w21ujDZFBgtDZ5gPKO8Zf
vXp6HQ2qCneA44L31jhszBpUYm+tzrpjeOSSkIhqdRi7Ev1aqbWI7VdsLO7sn+ys
aIRM5xGrQMpzJz6QYaKiRc+vA+qOv9dUEatXWd8tR1/mJt95xIG0kQ4aRr+joF8o
sO6Di+8OUaIvgPi092xGdqVRsrDda6y8ULs2ySl/Dd1JczzqZLezJnzrXSmYertN
g+gnTIyNABc5hyxthpjCqw8439xoQeSc8zoomwkenUYeMSuCOC+gItf3v0kHjfuI
99EQMRsZ/TUJ9kaUCjvmtd/U5DoSoGa/ST/QLDozaN4rP+uYEI2EjOte+J6Shz76
CoXgDGXIwcQpLT1vCN3xqsasKrTeCxpn9eDb6eZY0fo+XQY84CLWxfAz575hus/b
T0FLFQTMdVPOFymc7RwYTY1Cx6fRfXXTDgEebBTLWxURmNKFDqjwmJ8MJJP8dcY7
e6t+qMLUHB6MP2f4Ze0TsH67RqkKyVZYOJKzy67Wi2o+mancfp0et20RF6d02t1P
vvLUkUDGqUYf65loR3aD4ogIQ30+45RPxnRFQVpdku7W8qvpsUYBiSdt22d9HplR
ptb6SIqMsNaPLg5tBk92psQfj0pwrzUOjVwzcPc3R8xRL1sboVVyKfsMGa5p3L7e
nizC8scgxihl16jyDx1TE0dGel3W740wAbO2/HJ6bL8G/y0SDFv1iXWMYGKqifsW
ygqofsdcxqixkkQsbytsiC6F7FyrZN80QtYjvNNaX5wrVuKHglHoafEnVARafpvk
DOd03luF2b0iTVDPiTOoS+YN0QalP+7JtuDoIl0pqnqvRNtBph2Bof9OiLQkjAmT
i/3eA6++lOyAVzzLzUMn84upjNEB2AVT6Pc/4Sg3R69V9coZXmcjTcXHIEfRYsZo
Qn7gUKijFBNArba8vnoc2bxTELUO2mOo8AIClfbRFqStxZf1givZEnjWu7eduBXS
nu6XWuKrpZs+Z34rGQROnIkLYZcpsxKA0VwI0lunrd1YCLuH/1yliS7VZ9/SE5NE
541C0dBZ4K7CsTRSn954dVJ+KHKpQ9A2Wix/JJgqUsrNhp1/va3+K+NstxWiT5tU
LZCK8wVVUYY/9klVLWCgv2Fiojglfabr4hrbEVMc2PQlmIdFNRQKK7u76IVrSi0A
FOf90G17TsfqPvPSnV1K3twjHkWKA9uDriFfZwwZuXLp1lit+kfIlQispmDeSYyB
p3pPV489aDPvYJfb73dZTL7gMf2MX0mTIXkScc+xvUdIeAH4fYs3LS9gxC/vt6YC
BhA5zOaKeyCV7IrQj6tejG4U/rKhIoEPrba7XUVdqJzFbtYZc/GEysdx7Yau0fFQ
0zKzqQDwx6xBwy0jhZFGva2HKw2sTJYdoOW3StAaDnEP2Yh/FNNP3c3/ul1P6Air
vE+wL/Ko8rbEYdzaUWOLVbSPq4qqMHu3xqchc0x+WkJr+Xald8nYE6uBZCKYQYvG
whk4MUDPf+yf+gAHZuvYD+/sUpgvitkxp6b3ouM9KxVK2a5BD1T2FSL/PppL6MWM
3fHU2G2Om8OKZWhS+z1h0AoUNlNl4OFGesH2jJTlss25iRT7LalJgxb9qOZgDBes
j4BoXaRmk3Fl6Xgf5qOTDynAUS1UeP2wtpYjq/dpFY0lSXkfHMf0SKeWGwcv6cu7
dvUHXaM6qXmiJZn/VhieH/r9PKCxjM+JIuTGn7m8+o1geBFJAHPoDfPtnRI6Ll7A
+BujUcvPwV7/eETC3TMaS4ArUvTdsBUf/76lmCNn7qkvVGnq5uUcVReFEsjIiwOR
UVYWd3qOO68fMv/rH/v3qrBKvth2DZbaQ0pbjOHVqMbgwf0hTpRXdW3lUR48aCAA
Gr7OeN8Qh4OETdozBbuHTo6LDfHOr2Ru4vsTOmjas4N4lNFIpRp0xkaWeP5AF0xE
6sbAFZtxwI2zxzreFkrCgJM0lojnm2g1YCPzEnMxVVH7QKpNoKmIg1TwC8mYar5s
CMsaRh/Mpc9B+aAs2CXZTCJa9iXQNPEvxeZmlSyBX42RnQL/XJu3ZIg4gtPB3iWH
UDLP/Wxvnaj09m2zhet2EuSHL0IP5rue2DgMyyjUIBLeBcoRdN6FVE3txM486/x/
EOt8nwNGgFoevmm/aY5HP46SurPXl3VJ2Qp7+vfKKXDTfRPIJtsCfPmVLHg0KRzk
UHaHuxO+S8OegwstIQvDeSn9gscfHqfrmizPkk2dkbwdYoU0GJ7zdJhra41/2xDA
gfbNSCUK7xDZr138mxlL2j81q5gRr1qUbnqonYfuVjXpkvX/TrQuioyB5cE+a2Uf
x7G0f12e9Vho4KRDnko3HdfUsqfgYjK2TmgBIHJjh6iWU7yhCoKGaYaOl66X1RBO
3cxltYP2FTT38Xee6JrA8RCG8NsSLjbZ+BqfkBa+YMUs80feSnROQsZ5vEfXjtUB
JyPXhADtSF+/wykTqXSFQtZcMEZNlEAOxNwkFqQZxMiBuPnlTeTE66JBG22gMB7U
uOjfEfs3ZsiYdlSiEzwBVb4VM3OgH0s3uqrVVm+BpCEPqC/teE2r1ueBwqHxg8+4
7Lev1uusct8tDDOw0fjNIJgHzTmSjpi2FoZI6oLt4kbs8lz7M5VCjTmJb/5WgWh9
SDJ5Sun2Sp8gy+ZgmqqB1BfsecJZDuNqpjGRV+TwBekJqQuliyFvE9BKgvk7DblW
FkhaP4o1eigg3u7JlgJn3TZnPXbN4jpw6IA6BJQqJOXVk1TJZe33t4QqvFMSATUl
tnjw9e2LVyJY/7FIFZBNbWG2hjwQ1ObHUB6DVKZr0Jzu+MxcnONiVvFLkPmwpCKq
2G+C4ApT/CgdKsDIrz35O0JDa3/qxIJ/3yk3mBgJJlHHxa6R1KLeeN/5I0hrMYmw
5QQ9gJTFxT3P7XmHIuyafDKSfWV/hb2LbOPk4bCfLrMJm9MIWA98gCtg+nAwnUXx
Nc+p959m1ZWMJ051s7iyVEKUwe/kYc0qWPDhe/7nKZd8CNNP8vBHaTjRbfN4NQQj
dlnl1I25lJSkc6f0r/u6C85DzLOu1pGaNhr/bekyU/Lq3WxYXD4Uc83HC7H079gy
PxGbn5Hg8HtpIE3As9q/h6RC4aWzhv372zxS9CrD8YJACiPF960dUtDrVbgKA7yo
3lRPpS8ntExZPcmfmV6G9oe1mlSrzJpYCMJoEXF1a9Wbwqdh4iQyWTaWGnZPkD+K
tcNp8tatoxGiyf7ej9uYUuNV6MPQ1pvJSuLYcbKqwVfpvjrj+waF8d7nOvtBDhgm
OZI3W/y5HKvp6AcPEZ29MLxE2mV8o2MTsp0NbTTX7Fk3rBYZH1txogFxIjpXu6yD
8vaWt10RB22YuEgbFgJSFDvSq3xgK+g6S/I6NGwda4JrZz2avRq54wa573rtvkHY
l0kbdoemrjByPXrr+GBQ2Pf8ZDpC5v599JILdCEE1SPRwrk/m1DcEPfhRRSb1a6n
7MCUX76HDw2tYtTcap/jnJf2XzFW/EWUJaPsgfqN1MdL//XMuIhVIWxe9QgkLYZ/
XMmFQAYX68wOjUJ8hj0nMmr91QbQjzT0qA7WBGtEAfF8s0WupLnhq0Gg4yHLcrKZ
NllnqFgikTLwg04nCHRudLNeTBOERnxepzCkQB03AtYuAlGNchiy9NqS2fH49kJ5
7XHSn9QvXmaLXP93cmNp1GZrfpbVT3w6oKQzMb2r/WAVE630a0raa9cUmCbDtXZS
VrgkzAThab/6eIzOGJ7cz3RNWx+4Gux7WtHmwLeC9yUetJjjX3kf3yF+3Me9DQeA
g9X/tD62IEiku30I9bLqFV0MbSUJErhLuVkKjPgLvSf5l9IpG0btWIKm8OK/g7yY
NUZHEWxboICOcpJoAFWpYK4k/nlAlPFrMwfsuITQHSrLT/Kl1OVAsGry5ejsB3TT
eR4MeOGRKAep863doKO1Ic5dlaevlLkA+tqUKowVOYSJCbQmrywYQleveGUVxkxz
8OjK9gGPghyH8TrCDEeXq2sTrPRDwSGHVxCHPsUaCeGJBDEiczIZUEni6ctVjkN7
oSD31IBFtm+IFKMALE2qLT6A90dAXlQ08zz1SNDha0Q5LnnI2if+K1584NY3fTTK
dNy6mAr0C6jz4fF6cpRd+UIyYgagUIrDhUkQf0V5w+FhR4hvlTpJvT7MwX5IL1jw
BLA+wxPXaFEDe/GL0tlM7Pj334MbqO5vX9+vv3yhRfmK6ngUMVmmo25bTpDrInNb
sYl1WLPUB32+4IiI2QFhQv6zkYXc10YfS5QIpZRdcheJW5HhDQm95lzgUptE/Db5
e9GgrTK8w55nv+4t2nAZqO1RUCY0krzKrj7EFQGKG0ii3bX8LncZhgAX0vj68SKN
99jr7M49ZPPEyopvBhq5+n61ojARoyN0ToyVgI//4Ai1gijKva8bv+NRBlyTwNGt
KkDK95AVP2yW7b+gTyVB3bDdq1f7t4MD5MZH6ftGbsJKax0FYK+xWOx7bD1xDgBy
+MXFJEQrBxZVsicbcHlPn3oaFP2luzWEW34rdeYkKTCXHDGGtEG1RmXuLpaAy7lN
yAhd89kLgmLZ5zhpgSjriHeX59hiHYpCdkNHND4HbRQpBe0WQ8cSZG1TsZB4QRwG
alQtHyH62HmM69S2M135YFZJ6AfPv4Qnfq4d4yWoVcJKPVNGW6467PLt2oLWLAhk
q1ScDY/TO/ulV2pYzO0GyshbNH70gNGJDpXPl4z1G62MQ6wz9ArBIuywlK5nyZCC
ia7LNl1jauaOEkDiC8h4U6ByM1wVWkUktIPjWvNmGNKmB2jPZx5+mQilbDbm9HZo
keC5MaVly4CzUJs58GM+rWllrC+5EfS9XPE5g6xfGK34GZYJ4wZZ3jomjCVWqV8S
BRpSJcslvYsgCyzyZouXoYtPm0Bjd4BwRqj4mqF2Ry8Mmf/ESrnplwHozBLhaYaX
p+JGHnxsMxYlEETLV7ZZhBZLbzDemzPILPCL9Nx3GY5KClkJSR1jpFKrd3mGN+x5
crs1rZ0Q6OZAsMbFrALKzWDTIV6v3wrsHSG/iYbqNi6EH0J2o+74r88GH/iEAOYc
JZY/ChEJDmUk0fQFf25c/yEu94pNRsvedqzfkSZrMX0P493BtYta9trI90tzwTPo
Pk+D8/eRiF4nfKpVY6ofG2SN/0heceMSj15mS88cPenNvV0xgXeZKkE+brx4ZWGW
/4dsJ3RBp9oLxGWJlXQicEbRIZ/bhK4e5QFPB7bhxLKl2X11a68PvDgT4jdiJHXx
6KVkK8jHm0jMCZY/NZbogigQoEHrUTb1foNlyH3H4p1Ud86EpMuLyOAbkXcIkDo4
VIh88YWCQ+DR1jHxhZgWyWxPOaZkWDHxbMotcCm1mooqtXUMD+t+ZKjImxTBD+1R
bB6E0W1dKVvL3q8dQjHDW0WtS+/v5bOzX5PogVigmMMP3WWGLEqzkZAv7SJX7Jyk
tlg7JdQAhABeWIr2GJbKqIBfAaLRj0JouNunCNZHPrWJ3hYwxV65Kug3N3IqRpTw
OqoFgYKZSh75dgomXLl7gP2d85WvqqV/+075Mk/mzRHrpAamH3jbdI3Wf3cOCbwl
GBXy/tfRZrDsx9f7/B2Zju7ASDIuGv2RtiIyvF6dmXyRovyhDwRbKRJgBunW6anE
E4mkKdZlHLZyLimUwz01w+xQon/HinSQFqfCtesxB4uVKPcqWBOsLrGVPa4r1wW4
Axcj2pW2Q+roNhBA9RuYV1/bg8wBhe1a3L2XaQtEYAKziE++/c3m5058Rdt3iLMP
GEKAAi77IGk9bFORMUoFBcUXbwA3erFTw2MnM4ujAEHSq4VaQU0WCAdsPwNAXbpe
J39DAEnMJaihqQCKkexAo/AYvwMUTKcMM8oCbw8ixz9OH9WocHhfeQPAol0ngfXH
p4siMOuUBb25qi8NEgxvjYTb0j2liqfEEiyE/p4q8UacHz48vdbNTfqJAHd0CEJa
wIq9dhMmDJqxVzcx0d2RVD8f3PeOp1HzUxdkQwLlZ2Z5vobRU8mwzjx6un4iOUDO
ihOnHybPuKk1phuPkYHi6ErpvXxJ9S0HSodR5325Mb+4numFBo5ZqpQxeN11hEGq
zfehIxN1HylbgQelDuIm6mNSSjuBs0aBEImTU5Nlsr2Br5tkAsyNbWR9mMoEK0bc
BspzbXRrtoJOez3e8nST43dZdEcB9jbZLbFG8aZwwl4e6cyp/tu96BiYHaxq+nAA
6xN+PXvWwRdpXHp2bwNrMTFmkzb3gSP4h3CoMQOfnzv/gI/fAZBC5YbFD1bcGaPn
KekCvIjgk4X2c2ABMgSEPqUP3WArEvbGEOwJQrs+Ea+kVdVY/qqBRicI6MqLWpNq
ok2vFHLIijpFSEFsqnzpFikfxom18YyX1tbmBkzXSZN6WMhrJ/2p6OmPYQvSyZ04
KiMKpeXAJalLqjdw1NJ3PgclsXPwMWl0NAMAPcG8HmzOyWEbHF+AkueAW2Sxg5ZI
DnAGuToZS4NrPWRAmH65H9sGSwZArKB7J7f5F1acXnNAuJwwpd+xxsa4dFv8wBqZ
Hc19sI33zAxP7if3Q+Zhc8XA/Q9/s54twe0HAi2aQ9X26UZsbBkCIgbMPqE2a0uh
QTngujdDxFs9vcbTKQWKnWRSSMd5FEa8UdhZqlVxBXzxZmzsgDkD7IbsSkS5j+bl
7beavgX5Z7wlyf6h1Fv0w5AbEs1pJqfBFSlNWzRmo2btsh6RLMTLhCwjX5Bww946
Pu3G6JHiaM0P6CUnWkzc+qPMia93r90J8r7tfG5Ybrj12PhQRIOV9Zr9mzON/6Hk
S0hPBx9D1Tnnypbl/Gqz6Y9NRpbzPhIA6F/z7tGr2lofF/KNiZwVTTAifDDxGl46
47KAIg4zrfzGt5uLK9D1QggoUo9M3o97oHQVkRwMtaZplOKabIj/tA96Q0V3JpFc
ADUQGbIpI9XY3XmxtX7Rsg/Sq7HBOqbkOxC8PPVz7/LypUbCZeH+ZF69Pq6q4VFY
ZpbBMraP4fmv6tHzDnpVZIaGPffz2yonEnq0KEaeKhxo3l5/6y4pEvxiNekUpPAC
pc4XUae/qbvAOJcR8hS8O5IAmu1gDozxIZIW60v7kE77/n6IBNB5EW4SV+lBVHwm
YlRqZLnpCpMg7g04ZaTPemYeDEFVf0c83qF/LUoY7fuZv9lqYnAGulNUlrMdYbj7
Y0B+iKVjJQyLXdG45FZdCIa9o8qONPf6kpumY3OChat9VGKiwXDkDqmnGvGGx4Zp
9aUBvFcT3L7LZUBCGp+vHPq1maoGhMPXKUkmlsb6EeUlyS4tW7QEaJhcaHOTOeCc
iHNIpMwAPL5T3BYfuMruSHM7eQJfkBRnVWMpJqnYn71l7BSSxWz4WjHHXAgZ/zqX
x6763QnRLhOMxPwxvwKKkvllEHINcXTjghtAQKCKkvnmDJW1/OG6R3MuQbMDcGZa
YISNQsRItRmia0MZ5hUqAeKABsXXILTTwg7swoyNMJyzl6C+XMjGExXy/FQoha4F
PYQCT++RBlcZlMmQwkaqL96BQ8TgHYOVlSPknUuBQNG6SigqftXbP1ha2pUCJs76
g3cjrKgFub3JCRyDXtvRCV/99DvMmffdpmxyveA/zpd5e1XnSbOB9/IPF3/Sx2K4
RT2kEbXpgOtrlLGQraXTR59DFPiX8Pr0WtLzeVlPW37ivnIvj99htTI45WxneRY2
NPUlnctT2SQTy12zsaUPeS8XqMx92q9Xyi7l6jy2nZNTE3XVUVk2W5WwY4OAOg1U
fjmb/VSh47YGyvCVOKsBCKZbmCJ6JvQV677UJmmP51V8y1CdH7VkvOZ5dqkjqwVo
bAUqd/XUH5zDXNYTY5yanY4VE0nZ+tMtfUAZn711qTG8RECaybTwKSwhTTPfQ0Tl
Ysxb1IW70fQDgqDQPao9lQTSxXv4YNtuyEHeVb19UzRexB8cLHdKWiAc/Gfseiop
cB3lQdwHr+s1iSbEsjmF4dlPjwnhZloP76FeJuhXF9/uKQuwtI8tOHcj6l1b5ie9
AdZjT3nHkKoh9cNoQO5AWR6K4QMzxr6t9GBGTDUXmXluySksIGLHgE2O6hmUuJxA
1VC1O9pHwLMaKl8swQC56XZeMhtQEQg69XRifWt0ZsR6fk2VEaQqyDDPXDGbMCe3
M5TlcQ8MlLruiaPAqaGcRMjWO685z/b0cEARu6jo7s9rulUmnkZ0r+Q9dYYdpONg
TiC+K3KaJE4nHdcfZGCePN7zu5+RccjF2RNEuSjCi8pFN5wk3bz0bIRw7eJlGj4c
y+iwNy9ktuepDFYdS6N4WgmoJ66BSDPTLH11B6B6AGrl1Cg6eV/0vUSxhTOsaD3+
5OdtV8HlrOkm9hug4FQ12jq13raVpkHRvFybmN949qsPqq8xbF6GsRazIrFLSk8D
2Afymg3gUBkgJrMYTOHuarr/G4g3F6T7rR1GF63rmJm1nZsACyazEhJQX9JyZbFS
qSiC6nZ/MbdrUIOpW89kJHQCJKZ5QiqJeWIUXqdOgmRdDktrZARf9L6KJ4Hz6lH5
aisnpjEHInTcM+FIEPJuY0/5U/IBp0pB9HBoxtXJWXCGU4TSU4EKitlJfn9aoEm7
IGPH+FyskYtz2OH6AHpU32WtQwVcUFX+EFckdfLxyXjgpFz0r2jOcdRAZ/pX/FiQ
o9V4z9jX/HfFGTOV4PUB3vak4tn+8DyOfja4HEvqtYcNIQPFDhJPz04gFOXhkkOu
AR+ARdfIAGkbx0SyniDJPJjG4ngMhccSL6z5g7vfnqGNb+GHosEUEIEyImbA5kcV
j5gdXgdmSwVFWwmJlY0q155Iv3x+DldDociCN09yPFf6JG6XrFZ+7wkvrkRlTX0Y
Tk0ZU/fli8uazZUqODXY10tP0ckLUXsu9DsEiDTWGQ0sLrZkP9CY49Kr4qlbxcCQ
TqFWFcfr1Axyuec/n9R6KQDlWgBeuAPIgHScGyOBdXuIQRv8a4xRphQZJZ40IPky
4EbS7xTveXFCFZQfNViOGctNM+XhoH17wfBDqWrPbw915aAngJ/MJdU3ovd35P0F
aK+uAG2TDQFxA9/rudBEnutFm5m9XFAkspBJRmeHvdcn9Bptw/8keLJUfpMXHqpX
ZA0MZh/T76GryvUYB7R3vhEVdgUwQsexdSTMZcyGRnmTCse/AESbQVTTwEPeusGE
0pA+TsZJdg4PQizlXucKVSjmT+XIIZZAhl612d981ZpVK65LBJUbtGQspWOZ0Zrp
jY6QsT4qIEH7CJmLPYYL7MrjD1LsgAohMvqXrfFhEArFpUnSC6mucWiNYhO7CkaY
bxqogGK+TwuuUBKbtHNmIDyAytPXVjS1sYIXSgUGL/bfnz0a7cy0TinzWz/1SGJz
MvDO1evO13d72OJ1PQJl0y3drL6vnlMPEDon/HA/3MuZp4vG5KBA06TzxwSkhmew
aCurpEpHdD5yh4J/06qlRFsBCqaZSgO8AL0KZcdSSq9scbps8FiRYsRQYsH7yT+c
CAv6beDHDo41tUzf3c7lXI10FUu9mFKKh9PzzzLkylamoYxJCShUABpbojfdoNZI
zOYVcRX0mlNUMkM0wUeo3oN4dNHHrF8pCcoswwajWEW3T0o0pYxNQ4G3LdmimyUQ
qBIUtyr3e+QKcnV5Gc4oa0KBNkzIDWH6mzLzJbhZYMKaN/hL6WiJbSIerxIEFlOe
bCU4n0nPHFWYpR8UAf/HzhP8KBU6kWzftdU2AnPr1MpAHeHsO6FvevIsEQE5HrEv
ENNM08hiCjwzy98hVfM9LGKSlCEy0S2LLHmrIGsNpSBitd3bME54JuIHAT0o+M8a
AJu9Hz40wWP6UsGWRdPw9sAgwjeJLvo7P8KmriYCposUGyeAfBDPKG6qFmXdQOJY
YUASgP17cl+GRre8JFj6nHiU5Yemv6eg+OgOelAPxI0bpDPQICmm7i6OFzAjn9RO
yfpdEol/nB4TwFyhscjHCfwN8uNxbWVv168zlL/wbKqPdtdxhI+UOpCEWqXEbnrb
QsLCzzdTKCxntYF810UB4xkwZQnDN5+8S0FUAtgnFT5HwqtmmcrBEAhNdAdegFM3
KRPwhypYy/LMhM6eCjjHfLBb3298sKEJTiHD5nNk8cMF8GidI7VNSSF5DOPph8Sx
aTWD0eogqULzQ67eSaSnXMkphagC6ytAsuqPI0fYRCgrdjsDPifJ8OeaP3glMK6m
4wpLrz1HPQ2kY41NQIxeJDQU8o6a0kswMSGj1FCf1OICxdDiTgsFp/ox1sfTdYBm
GShgo+zgroHaE7eSqb7OvbRjWSmKFV5odf9iAfetjnTS1Ei55Or+yaeB3ABvombj
emMHlZsPMQyOaepKofmjUyK14QxW/UOJPWLt4NfT8vM621M2B3b9WIqzM/y2e6c1
2355LSXGTG9JakO9Y9xa2NEuzta+bZhzPBp3YFsO/TsNyPYYzb/WHvl3VHUWb6YX
kwIWM1vSs2gKJfm0i3CQE5K61QSSux6fC/QiBH/iYZRzYP//WdjwH3lnfy06ht9l
S6WTLJX7n72rjKLSpKYzwgV6J6RYw4QZd5M57x+5doyZsmYxIc1ugS/NpguaJLkN
+kk4L8QJRCAzwyFBO3jNdutiyb371IolF5maQr0JvfrL8rXdapdIg3rgWB5arPOm
HP2n4mfpaVp/IVQyrjvZPDe2AaucQ+0IvGA2w5YuxnBDMyTXnwP3noUfpAD1Gkt9
gPdwCpE7sg9iWeAj1QEA78QYuGl1OnA/81xDyLN7UKHl3Fhk0SGvQmI35u7tAaV9
ko7V8b2qJUz+Fq0sph05pk6pkRMZts8t44B91e3AjuSekYPGiZnAJKS8AR+Qg8V8
S1EBdjKkA43I0UTjz6QXsjxUEAbp6MMhfVjHuBpKp8X5+g3Pi2VPkGBLKfZrt7Gl
G+S6b2krUnb3/+5mYSbTtyn6XH4BO5P0HczLtxiYwaZ3L9D5GHeHKX15IQYQ/Gri
chd6b10DytFex1E3S0s3UbstcYXPoIpRDc73jq1CR9K5slmh6L3eNZ8B5kky1oNo
QA7RnqAoGtm8ji4CkVhaZT80EOSIYX5WYvksgnfayUD8mHcvi38OxF1kZvFyQoAY
U51Ots48rFlfP/x5C1GrGH0P9XbPMDbkOVJJNgz0mBceiaz0Xp7dqz2z+lU2z5A4
SM66ksMUvDZiY402paJ8LsJjlycEPt6N6GSlhuXb7FBxKq5jV0XaGEV1pxQrClO5
kB7C56MobzsgqLitzv84a/LaPwGxJ64G1uwYSGh2Q+0SrtJAtdlznb6lZg9uALNN
MffWPs/vkSqL+HaS72NRYKMf4BWBtmaPsjRk1XIKAKtVUuBv2BRBElq+C2pgKT4T
eqr28Rji6pazjViE3SMhNzM45nEtjqCJTxtSuhNPucZ9i7n91KYtoJpTqSUMbABt
sPmNdMWm1xAhuLzH6NWpZ4zOTTxni5EZScAlR9/+av3zJHfeqKSF2qoQcfrNxNz0
lVzO3bAOTTSOJeJaKHlchj2ElzA996411SXyLwGy9cEheMLT5Ju+CnhYGnzg370g
/l3QWYAe8V6tbW4MkrX07zH+57iY3F4Bz1XJSRJw07y1ehL2gChKmQCavol5Zy5g
5QOzDweRCELhEVHiIm0ngg9J093nNFPu6QNv1FP2xmoqgVKS6gUSzNMUBBe82n1P
tCR8Ia1dmIJ7MdA57Rf1IAOkV6LVdihrwcQvtDW7B2ymht51DSFTD3ifdIjIdPN8
w+JCtq8ABldGX3Mk0+heB+vLNlrabPuwnEeANT7DnVfwV/3zKv5/wFA/6JlX9Mk5
5M0sxlflCDklKhyBag717EFKjYJk+GvIkxWIbY68+y+viXgNeyOstvC8qJnVx0KZ
p5dE/zfPFiadyUzI0e/1Wtp1bfY5tZQcEx51O5z938g39+GMo9k7t5J8d6FdNZp0
OCph/LbNFAxVNtpDiRpSo4tat9L5sBmgM8K4XeWOMjBXacFOU0R0+X2sfhvi3o1A
48aXzEMqSgaw2iVTYvFoWqcR1Bl98R7NLCsZr5WQcsS1Yadh1TkARRZQYmwZ5s8T
lpLUqA5+eK5iOMsMiTGUUr/MnmpwtIhoxE1kHghsj1NorWGAF1wuUQl83uJPNgrD
X+YrdJNY24GICcl+iEFEyaB1iLQRshEFGIsOrXSaj1fVHfWKf0vJKoyDwnNybE9i
R229G4macBc0LwQtGD2Fc8TO/tb52vi0LZlsuSjnrPCXbO5DN4cVnE40WXsBc9FU
KAs2btAxxNFMN1TUYYcHUxhu0CsXg9aLVzVKPQJgsVYip6M0CfWPc1Vvc525ojek
i6ZREDEV+U9GF/5yBycIyc8bq1jdXv2klGNDidy8I+RFTfvXEKeAC43dhMBdFvFS
jNJLJAnuPbnmtrdCPBOoMFC7/pxvpzu5n+9rYxryyyTByrqPBwq/aNPzaMZSW7IU
3RYeZnUFkPnDyr16hNdEUqQKbumFuRVQJqpVjLTmexQgGmDv4sv7km3dLZbh84tw
aK91nlaBb+LWayRDs74JbUQgnPzShWjpdv2nNqOcXmeepBaxaFZLszid4OvBxPao
FVdJmApYeAEj6rWo9N0t+V438MI6qYEwEASVxL03Sz0UV7JzjNj9pjFR7tIye6EW
rSbvbocY2Ggt/dWD4iJb0vxjsnhjtil0wJELofd07XkrX/xF/YAQU7PRfHOlhMmL
os+cD6Z591/RFe3jgnph/IufSh5kSOElVe1TcLHiEaOX134fuzTfgSR/x1Z2yMEl
Ly4NGU4kiX3izeChUsg1qIpr8mnNQbJt48hbatbsPDMsMBGaSdTBh+lXoufg8UhX
3x/Sm/8Ed24i7gCECAfQ6sHznG6W09v0HyLNiOzpsoscBjIkQmRcxI8WHO/HiwOu
82CyNCWJoEcmQ6dZIxYPRXt5oexfDf2kepz5AJ1lMYHimVJKx1ExwUyVJnSuB1I+
9WULJ0lqLQfUfCFpExIJ0fHbZiQU6sIva2iijB9XsmSmSFhwJj5k8czDyBTGg9ec
ZJIsTajWqEx0HmUWS01C5TmUbZteiJomz6TG9gRppoH7vvZRXni0UUpwcpAnXbiI
Bzb7VydK+CQdhXjDlKfSYYi6DVcoK/VwkKRJyjdOs8A0HL5zRx8u+lKPPeDDJpmo
HS5dMl7sMVTlMke3ZGS0kfs6LvWG8kDQVaqzZAuySjP3dZPBWorUGmBmITccJh6e
fS4Zsd4zlQ8z9B7M2hBfusVId/NvCMsOd8CwpAgwg+s7Gc+HQWvcXVuyt4FFDELm
JDScdSif3l84tJCJCZM5BlbflJ6G9OvX1fs1oOEEMHr09kdMqCLQ1inKeMun0IRA
gdw8RDvABCCJB9VMq94/l/Q2NGvw7HQWBmYNYlfCEFnbf8/TxOh3wL7pE5sBLB4H
8pptiwIpbxd/BJ6BCoITr+OgRcVP4yZ+Mmd7GqFfnWKXq2mJQ/8La0Vz5AAcTYYa
XPuC0nSaJ9nMHnwVUyIMLZXdNcIfezoEwM98FI+IypRGmPIYmhk8ONCd0nSmjTve
pIurl/566vz8BZAta7o/XDT4AX9pzAGAhRwBENYOh7VToNna9HaPLcN0jctx7J+4
uimR92wYQv+M5OMhi94ag47KkP2lUQVdNjQf0SD4tz32dT/7al5R3+Uxi/g0EO5P
zFB5Nd2INickeYi34dzyr8K5JMjK71/bSkdFjslsOGpv/ybSGVHFMeaFRTlVnUHF
iRGT/KFlUsAMozqZ8JcHXbym0QAalcgFIqT20rX1NxysAWP4/3cTwE0o6Mui7wHo
BkQErEOuPrljYQsLuQnGdkvSR/g6P6j5w+tu88lI1qwSLWX+jQ8179i/axE/53Z6
4fyWBPHs9psXZMWKYb2altdTYzdSqn7zTseJWdCJQqmgjPw2BM9zMN5fO/cq5+pH
ZWfk0RoLHmBns4DVzo5ya0uD8shfnuVoU4P6l85M1YdzDom5GXKsXkVKEENGbNvd
GiWHvgG/9itnYVJFFjczzw7b9TQAfSuWl2K94nRSbQgw6S+HqiGvHlZDToxmYh8S
dnekzFomInuu2wl1fAUwuqB6Em5+gkNiLHK3ie3HBrjpypvfRVJnMyxdx1lk7+Iq
nbu/UIo8IhgVkCjwzAw0fIC1vETSNHRYuKjBl0myNhWf8Koq07LqT5XKyOnO4OqY
RUJ2dQRjE9T6xKzilxeuJ0JNgJ22/cHSWk+YgOHjiP1O0EMCTX5zovldu7EXQpKF
1PNQIWI6Z2k97GgmcefYNmzSA9mGQZShtAfGyQNgn5dLOMc/Ga+RS35dPE90ps0v
MIAII4j5X7katoY/AIUaLDXzVTFpvBg3RXPJ79pyUjEWecZIHVx3YREg8IFZWFTt
nB4d5ksPUKVdeL97Y4Y9ff1H7gXGNA4bYoMRJ3GC9i5W1T7L2bjBsgRIhOiDaIT+
X2KwxICSKJu0/XxYFdXg8VUyWG77/mFTSrqBMuybsL8RvH5hGFju1AfcWMN+MUYt
Hl+AXcdbb6rdaT+4/qGr7XndBrhNfVs9fyzoOQdLo8J4QgtmRzFTWw8qkDzDmUCq
NRnQz3ObfoSvscA1RZOwuc4L9q4gpEqSBx1YUeDGg/N9GrzZl4sjR/IJUVJ/ArQ4
iBEfwG1w83gXu2CcDgMXZKwPw84ppQQNJjGENOIuq/Xqk3BqS43P0X91HKfOmvyt
929Df2O9GRGMAGvIWHnW8tzwzrOYoYo1Cr+CXAl9+lmq6DUdZpeN9K1AZ37prz+w
rhqbRiAx7yctPeN5soxNGKj9u2bv+Iq2afiGpuGcBShjeIZVZhu6dx8+W7yLfeKE
7sG4dwM1Ld9cTTgWSBWh8Hopt5IKhq/i/AwQCtu9uyna2/ymIJA5ZEElWkHyxmZ8
E31Brj4f1RMF60bS+zijdrwgK2TiNLzokKkBpDx8gpccKRo2RGnd4HcFsMMFVfVF
hq5CtCuw7SKrGZFG9FtY6yO9+2z7tBKNU1uTBsek0osgMVSY5iF/l8isWWrl7UuE
t3OqFM1jWdK6GPqcZrGwbSNbfi8VZOWSZFadathvFIgegVXiOjllFNyrIdp8pdIb
qTQ++DiyAk2lk1hlqEMo8qqMbfrautcO4nmCap7KxhLeJl2cD11S/ggZRvg09B+d
YLndZAvC4boJZA2GG7Tuc3W9+5sItuU9+ICnd444wv0sYa50+/LS5OiG5VA/6Nd0
VGlvm+FenUErDhdAPx5ktuq1MmO4/OlY/gYoqMVZt1gEDnMlut63o5YKwgxdSxGn
6KnevQ5Jbw1bCWfIbBFGtBvh/RM2QW60QZMvQqRTowx3JwFi0UKo5/FexYarZuyN
Q3gDGIWEofOEqg2o/aeQlSG4Zns/PZaT597uUEbr06ybEuY3MLE8Q83vx7WKloAd
OpFZ8rINJF9QyhJUqjPnNgNJSpKUg1nB+BYMFUXmpqLWiFsHOrHLcXRgAPghrVtB
tT8zXtD9/HpPtIvQ0IRRhrPRt83QAqawvdvIDsJDcMRMxc6/N/XOzSykWFLWr7oe
g5ufrsU8H5uNkJwngjhvSOsV/Im0VFPEbRSMWkcUZylqXuvPAADcEmQbuBAT33BW
HhI0viySj69nSzeG3wg2v940C9rzt4Yo8GAG/AvxhCnlwjAjgc+bCHiY9lQYaonW
xS6aNkCTl8HQ+0qJp6h+7xBQcBuJ3rmnsjpcLNmrXwM3gyO2mW4iloWaiPrlW+Nl
b/32zfhkOsf3dYVEswfpQI3flUmCW038G6eU8LGWqE1XMuiGEfKZwonoRuOFQC7X
n6V+4xs9l9UmKapyZ2rxvK9pSRTfvpBQpYV5xc1QABZxMawSBB1hC0ucUuR8Fzdv
5sfEPTpf9rpSk1YnuVxwHVFyGSVz/mtDymfWr6rInIyhy6IwBOZn1e3KOh4XughU
p8hKsJpOiko+uNil0XxMV+dJyrEH8B3CDrVFlTroRx2cQiTedb5tUVUAshnCECtp
u9tr4ntCZFF70zOFnJL5fcMYPvo2KxiLJS+VeyuCV5JdZGiBuIoGmYrcWiTJvel8
XUhxb6ehsZ/Z2UcI+EwHEvzusMTkUxe+jlzzJEB+ahOiT+zCnV0rmefd0G5gpY8M
XVk6zzyAu41jgUn5BfW6U32v7fUHXGR9sX+3BAJILwLqWs1dyD/kqCn1jXC/Hzcz
H05xU0eB3jVOzEJfBCXgjNf3OBkejiN7vlMdhAZTjLvC8yGBn1aVU5mL2IR8DjEH
QYNuC1ckb1cXThJ77BHvmg3A46Ux3g8gtieAb7nhZ1YIO/jkmvKJu1WgfRhxMqi/
f1MF1g1NOIAWEp8HTqXxX3EixcZutcPxtDx0sRSPnqJM5E3VOjxn3FYeRqur2YPr
JOowzUT3Bq4GVKDysM0WUikyfqHIhb6m9o5S+S6vug1qRNsIBt13i70et7tsBkCN
eElJV9uUhCBm2xEgSFpul9dM+mWxBsYITfdvExBLGQa4WV2QQTVcBRycHObWQ61S
9cF5G9/vyqwKgcg3eAEOEjflAzNTqow+v0+sISpqEOiobbZLtjcYuSRat1DSA3ku
cNKyhtTrMVOaZmT4NNjqAmF9+k1HbDphvgG+265f44XLpzoCNY+BkqVu+Tui3Aog
3OzetKQ5o8XQ6JGPbyTZAbC44yatIKd809L9/1hckrJLytFwYIC1Ibgt4l2xvmVM
Oq+rbBU4sFPDev6lNRB/Xnr1uT/qoPvOnURO/cF5AJYanVmcCcv0NhuKZbwglGor
7orBIqryfX3I9U5pES/dlTMO8488zV+JI8we6Adu93fMlzCgvnyI2uF8qq/Dks7S
Jfa5K8Tv8VeqmDPQvvL6St7IcDO4NLG7O0YRhloTRDpCO0SFf0YglKakSuq4GW3d
Z8d/jd8mhq/a33VJcRqPcYAbUQPYCpwCjOyo3Y/DHqg8RQdlbei8eEhFfZzU7piY
rgn6vJvTNz01FuxwW+w05hjmImTYADqJV817jRo+KeLY8v2PCYrKxq9Nzglb3Sx6
hTpxDJZgHDVqARhPa1jjxPBtsTszjk9oV0N/cR+hKE4wn/IiZYQ7FlexKyj/7Sce
xxwjZWm1HW3p4H1ukst8v+OvmriweVIvYPqz8w3PCC4zOmjy9z2GhkBojVJuiLFx
X7injQ7QB+ORUUaXoZUXmsXFeLUO/qELgXGtXEqF+BBydEZ9SWdrVkq+jygEmYWM
6GPusp2WX7prYQ+io+7rM4UXiSdVkdJ43nMhPHgBpbtL6bCWQBYeGRu9m5xx+HUj
7c4kzD0mpcZVxx23kwWELmuXz9Bv7nW7al2GND6GtZ7SjQJgR68aEd0JMKjcPtRO
KZL+jwqQ+rO57ormPJqa8WL7RQWvltgysbvYw3X4volrLfiAjZP53+xLzKYnGUNj
FkWFxI87SYcPaN87MnSNOyApv+xSZtY8pKawBF76OTAKhkR1NCY0HHSaXA9xtPj1
t1YYxm1nCaelf7XOuDsZo25RKczzPza0NVcw5aAQvRfL2uG3DAcWoITtszlGEJXW
DZSzVkL9SdNoQYGB2X7MfajDEqtQkVGBDjbvhOV3h9NbpzyH1FcsjXUlsT9/e2AE
/T7FxmkztwJfSUCrnQspbt8B1JZRH7j5VETll7M0TNCoFGpGCcXL1sCHkt6FBzyr
AzpyD49Mf/aaVjXHpD5g7kVw8OZ5cxohhzPmeykG2wB2uKaP5TcpjgsBuWqEMP0i
avQSX3ELgrfpvgJ/zGuXSajuzw8PQ3QgCrQXTwia0y8jGOqlawR+wO1oSjLVAfgn
Goql3U29tCWQqufrfeLs9Uz6WNin15vKLdxtoA3hpM0VQatkKfA1XOrgwVNYlJVs
+HbBQelTW9PiujnCSDAs8qMWzaXbhKJlM+h7ByeytVqwJZ5YmH3TDDrh6NKOuRqs
Xvx6JD/9vylQfiaFI8IQAaUnlk+gGm0Rx5s1W6vDmq4GB1tEM00C54qxjIuWNvwt
kO3I4pk32sj4M70MwexK5FPpCtXle97GP4bijTnC9lwbZITa2CTE+hqi2HKtMLtU
F/I8+CQBGzJDhIGqQt4Iqf0qhxgW8nIBdbUKl3fBUMVsF/nQvM1kU4UERp5KTOOf
BbH3pY7vgHnaKmW0drg1sKin0WUPn/G+pUDc/DjsM4P4Y9FtrVhNMFBQ/ZlC7Qsu
gKyRhzE4yZ+e/680kM/IJbR41a1pqGlx0r+VicPUHpJKsevNAB3iTSPbgCuKQmdu
n1yOhZuEAY3cxojaLBQWElVnv4AS3fWeKQWR7c8Wuxwd/STCtYxgQkNqWL2O8g+c
DsLxnmvMeOXhc2a1O5+NG4J3UzGVMAglRYOQfhgcmIQvlX0i+Nu1OSmVkVGcJKQ0
ltwBc+TSyuRbwN7giRz4sslMPtqnKa4MyFJy/at+hr0l5ZjhyL3OPjXQd1uq2qNk
ROpCO6e+5s2FW+SyT0PyTPJwDT03Zg1fJGRBsqGeVEsYg8SS0+k4UcWa8ow7Q7fY
TpE6ksdAKxdRDx3OOZfDr9Tka0N0RieN+82Y6bu4H2689d2jNz3MT2debXHHUF16
EKRvYnWPwZ54cbiJhhbDYY9sWgIVXxGRKhJkO3ZG8Ctt9xsKjrCBIglHZN6XzH3l
usvQqFoehx7h3EtnjeJC6FsUgx+RdQg7FAHj+hYvcr001ZQt24Fx/8f53Zf6+Fsh
Q+1DJ16tTk/btZVE+bu50qkDVK5beLt8N6xYdfSsjwDRIfYCZhVnXRBEo3CQDn1y
YbnJRIWDiIuaGrUM/MGnwO9XAyDRiX3jDoE6aw5sAJmqsBNWEjKDO7Cnw/QnAEGb
2YGMgTpaztCNQV+GuTqCTho5hGHby07D0A7QC+9agaqQIkZLTPamULxs9sB3F4ii
sXb5McIA/KPH8GW+5LgJf0jTAgwbvHOncRNX7sLpIN2dFZwNNpUP4wQH8zSFfT4Q
14P3uWLo93z3OfifRCZhbQPKcvVZ2+NjxMTYWww1X+6NKDZUBHztVPpC6tw6GQ1i
m2/MitBvmzR11rI36LnWM0K1yB6Vp9dz1myeeVIUyZ45ZbYI6TKC2r3IjrETZZ07
522+PEK5p44awB0R/+fFtzSOVg6PIXD+kkUslsjJNbHKbw0SjfsJ4o+i3xPneKYE
SIxJhZxF8E34aflSe4UT3p6qdLLLJIV/B5lUfBEN97vXOgdDqGh9/csk1ZTbXxe4
L+BP3I91c1YROV294NQ54IGZh3QjK3eC7+XO+NbehRrBkZuYu5sK1SEZk+bA73J4
WbgOikDRCFM1xI9jYdl34b+xWGkWPWmUJKNHaJPB2iyR3mklWauJjYZDQtobVH7w
UI2Hxd5GNNEGO6JVv8Fbw9Q8qffnVo2TVzH7IHbURh0BE5F1WU5/A7Iuc8u75Ahg
/kEYUFflOKglCeTTo3YNrr2hNyZ202hXcFYOnF+BCu4wHMfh/SaCtEcw/3NsgxBH
SgpxK0bZrYbOYay+/KLv6ols0WkcU6KWGLqrz1YJpMuMkDnlnM1axM/DXuOOYnuj
wZ5m0O0ng1IQrvZemrN546jywJUckYsD4hI2+QTMesUUa0GKRLaz7LJi7DnidDiW
eAbGQPvMLkxlfi3Ex6czTfNUWlLlXKAsneQRTV6e3EGo4XBQhN9R5HLS2E8lfxL6
d0/C5YwnzHVZiiO3wDoE7p2sgAZ32EizNT8ipSrZEYtqv8TE5AZlGFTrtxRUshP3
WCpmHu0jNkBUoqUvseZI6G1pJ5lQd914aMiQZCBiO7tCEN2BFn1B3HX35OTmzCC8
w2Tg0dKuVtTujmyByU9UhfF6UI3Nz/oy3r/Vsg1/t5ITFEDl9J/PqsXY910usuJ9
9qnux+KlclRSfV/F7T68ZizBhepkYnl7TaWeOO/iKhhJi2Xr4T2Ae9T3476ObPMJ
12KjDlD3lk1Vjusb7yxkeZoBX99oYjJZgM99rTKGmcWK8+zW99Ym8simk2FO04mu
mrf/o4T4JhykVJZHaODxnz4+AaORfDgVx9VAtP5AhNk8R+lerClEsdQPvD5ANxuK
GeWOHf2DMmhTAzQAxu4szHiPCitpiI0jjMUvDXxpxxusIbEca8MJwlKQlPtkyhRJ
7n1xtAAE6ANwRwwdT12Ab2VLd3fPwxSfLn4QczLvwQFfM31YngvsroOLq8EJ4Dmr
N0Uvj6Py62WdoV3h/0y7lc7O9uqjZIKgYM81Xz5RRZtJWMzL3d361Sl+5zIRpwC7
ckeKo2E/8Js4+kXt/kYo4VM0QSEWjq7lNgDNeptOUT4BSbkUQHegbE9WV1U+KU7p
zBOZmS4XQyPcpzQxG5qmQtwi3Vso5Y2j7O6RDum8kgLSDVWIQQv5Ut2DU+rQScPF
QqRwwkzW+AK5jvPq9Fb/bg6WVtxXrOPTxrd3a9m3iBmBGwO7NR8KRHroTex+psVV
4X8+cNjV0PdYuF99S/e22qUJhasWKYFNdXNEniZYU24bOk/T/F2G39qgG4blmjQo
s3syWvKv0U0lN8cgPUo5oAOLauFpIgOmTQeKht6CVz8TVqP7k+2W+gzzq2mgCPRO
sRddtsZCOGz+SdBTLmIXjWW1IukAHG8qx7AVfAfIF8XkERpj0h8n5/Bbmu1BNg+c
9DVNPmDAlW3Ve00Mt4wDrikE7hN6BIgto4qQ1O22+T9fekd1E2cBfZ4A4s9WEAuD
eW6I8wp1HbXIi7pXh2KISbDDxJi+8kAY3MwzZK5dwfPfzwkgTRZ7e+rIa7kjonCL
m6UKBit736NCbExxHX2FUT4yZrNq91XhYDPKiRoEv1w/PHPn+iVlOtIYN1r0ZE5c
mnacR0vtPFS9e+YkMiVBV2kxMm7xTNxHJuNBVdKZlcxRPPyUQETd65H/y5pu1Ht6
tpY2EBCCc3HmmGNbp35yuuPDYkO3hRJJ5mpRkwYcxxfU79avvk793xTvSnozgSY6
6dyny6kxKDNYZt2nMqHRX7NYdibwXhFN9BlJwnrd6a8/Rluy6dOZ9wMDb4sTtsei
iYEwph3k/7sCFScunzAK/Eqx0PXobSEnKHM2b+07DwlNms1rarGOC1lKTxK+3D5C
zTQdYZHga5M95iZlfTYGXG+E6MxAi8w+y4B57tO42FFbmNnXcSqxHIH7r7gTvtZp
xsggVT8tfwrMJGfhRvgcsrVF9rsQy7TjRjyTboj70KgfTccwH6WsRvFp730kCowD
CBf7Cu63Skl0bXwGsil6AoKyKZpZOBT3vlHdB3VGiTzSbxeSqcErgG48BP0644VS
bm5mzUb9DXfwTiDAOsD0PwhhnjnNkJM6GLxjcfD3brFZFHaAcEXq+ZfA3Zclo9HP
vNfhrcMTFEWWWdHA+RORpz5oKaWbaDPrbFrExJM7AXy2d0yy2GJpWLUQQ0csNO2T
IwlY51awE/4RsmFGDy0umQH0UngnChwwVaXRKZPc2d0nqI2Be0maxA+MP/lwXft3
XzZo7B3bXm+9hjJWln9/K1ruybf2GxPWuI56m6HYufpCp1gc1CD7bn49EKIWVDQ3
9JroYuUgV+v/0ZZiQABcMitrf5AMokCPgq2Y80Id8RLLRRG5zGUvzA+JANGNpEq6
tbCt7WtL2jc5IO4VUZzwD0cmz+nFuKLTGlkIGupcOD0kzdxqcQW7IWJvIbcJH8N7
MnigSZCv9Vdjq89xHFkL6D9fnBAW2m53FOmjc2fdOEoHCL2L+zc9Aum9bbrvsTzv
pQTjlZNV/Cg+y4drFGTreKFYomOdbwIWtFL6rnTHRbbkTJSOHbC883FhLVmVo2tG
mm5stp/jYwjMSgejK86gt+K9tBEcKkmNniNbC0B9nydpYwmRJOCm41rpi0Wrjkmf
YLDYCP9wxA7G3uUPJ5feiapYUCp29GWRJyFfKq84te9FG37Vp1k2gdyImIzfO5Ww
vaD37V0NQ6VFDMMgbxzFjY8y+CnxkIYxTpISWKgE/MRun6pTUwa2HeTbGtfq8+/P
vAPP4ISky9evvWHjmOSzxrktJMwchWaehDvw+F9fEzbqBOHNNRExlIhAfjLIHTO3
+d0eGJSiHCXDXEphTEOacN+Qg/4Byl/4p3DtbDhmYw93Ld+7nDNsHPM4f10/lxg1
xc/7Z9H2/qXjQDPgV6kh9/rkiS2X9uBQCvRSWy4VAjwBnaVfAQuv7iwKzq2FfJf8
36yHHJTRwzam9BoOU05DdLvcagcxjXF5I79i8B/dJTZbCRcFpddG4cE91+9smDNa
bsfuaxCLUInTeXWlNdLS6Qw4QWjvRbSB0ntgkU8QX5/ywEVwywNMH+7KPMQoKrcY
kOQmWHUKgxvlohK7J33vnmDS4z4ruFTqXegMBNHCVfMrCY/GClCE4hwXUJ4VXewX
LhxgLtaW7N8WY+9F2UKIwjui/wT56n0Z0RPKYzNs3FCnCfxVljZVqA6BnqcIPPAU
k8Ijl5zU+s6XdvpX8sPngWqI1MFYWK/+WT/587K+SlxNN5IUcf0QC3za/+0qIJw1
a+X0+ndFVTf4oP2o6Q9kQlxgtxXEL2zQGEod7X32DSac2uMO7ey0zUNHXu5han4r
GxkoET3D645ilcGsbIyF/QPZp3unP8rLgRn43VyvFNhP2do+ApO9nlt97KKwaI6o
vUhXX+jY3ovK1lAayis8/zxf414CGu63K7x1dA8vpLJmWPr3LcI/hZ4wCcy9gEBZ
claByDm+C1iyKgSG2TYd7oj6g1hWdktfhbN0584Granahwjo+ShMPkL5umk5jqIN
KbCl8kWmiNyxf/eSMnBRe31QmSf1fKzLppTsQtfR3b0QKPe8+RLcessGa5Q4i2q4
C9dzgiJtiZ/7W8+2swfCvMTfI0HnNrtUz61GFyr6MOtUVqrlnxbejtexvN4Uh+R4
3cvnx2Afmk4TtE5X6BALjRKz+ypysGE+QdCBEvWOjOhrsqFOfVpHb5hdvY8RHxhO
li1Nf4Qsb5TuB3PNdo2Tz79If90OciArqHLqihPBg4Djid8AOyIUFllZMb/iP48w
XLX8j2T07hWXlMvT5fx6IQrADNjqQVP15ysw7hW6TNxsWlx7jvuAcs+nFe6ciXlS
r8eryTnK98LPUteWIt50NxGL+JecGOUWMK3G2HlWQ5M+bzvuDP2kTZPW8GOj4Yyo
/5mIF58NMtqX2USyyVR5ccXerHi1pOZiCitIHj8dWMdezz1+QVadMCH2RwGtOqK1
s6PwTT0aaY8VGY35Ke11Cax3NSDlLD4W3UqZqA55euoWh17mZe0xVi3Yy5p6BTfk
cunXWfoqLgtW9nv7oKbyr3FIMS/UNn7SE+YlzCnjsQmDQeghyJQwB9RykNo27tA2
BWDz3VvWR5DsmrZXO4tuSk1O3IKct1ChLfIguTvKrcK+uuPLCy4WvvDLX7hKlUfL
ELU4mkfHn3d9aI1xW6hMnsIA2Zn7gMPT1imQEzGwu5iMchMCcCxdvTqIyU/xR8nX
08ZRL2hchFdJcyhA7cydYhtfvAjdTIY2m/k5IRC6Su8dZU3WDAQnsNB2Lmu8CV3Q
ooSgiTz/ek8VBvlySqlPSVaxyol29/6uFqGJooVB33u2hYcM2bdj05dxDrc1Bhn+
hwFwzOq1mCQBB/ldRCMQWCQ+cd5nDnRAS5QFVNhobBKmifdLMNs0kiI3o3QM+KMI
i+RDH0WpUtAnPEqJKft8Nc3LPWi0xVZMPLp4vZhUMyhCsueaSLts/R36NJyDD/Lk
I+XNS1Dmk1Kl/XEQKsiQUPWmYASjX7kNz6oEGVuCE/8fz5ZsjHiZakTgfikBOJpx
Ktq0X3jNSzid55OSPZN0S5xpL3O4E98kIj2N7pHUVJFctfOnpQmbA8KfCV8OGl5c
P+O6NsWe4NghvK70jnK1b1r1N6XCDhYq8gXNk9qfnAyZu3e5bWv6W1dDljP1VsFx
6O3413KH83OW38W6nERe4sc2IFR62jry5ZOrufnUmuIiI18wpwj5xPzpL0547O8y
Y+FAewfUONAgVIwT2f+uv//snAe87wm8JB1SjqhfFa6pbKaNFyCnnvQ2aKoJoxBy
1jl8eX4cISzuq/vTH8G/NnQQX+hinBM7eRFUhnnGU9XtXQ5sTeG4D7dQR+0AHpOe
iDttTFHIQSw2f4zyH7tISHnxv7zyyHU+XdeBufeISgxCHDfFMJ4HWWdVAfq65KYc
8zmv+avTWPyLQfh/BT6IgVmM6vNhoqeAaJslPN4eQ1wA2mu4fn1RBKEJEdBlg9A3
8J9Z4i4Su9REA4elMBjojASV02Z5yH3yGnBDVErWs8jOBNOMCJnXAQwCv3W1bR68
l6cHIAahU+MxKhOrZZk4/M8UZ3/hts3oGNexvabAUTqO+FYimXFE40PmQ8u9FYaK
ylr4RBhX3KdHMjwIB8vu+IMRMpk+DP6x0+oWHbQ1ZPVOVnveIEQqFduQW3uFI/hB
qsD4yOJh3OmUXNAlwQZunblb7w0LA4wq9XrBBv+cWznh0tK4DY6jjyHerotMVLxH
T3wJA4qAZAqsxylJbTNjfzBQVPEEhNBPZ0VQdoStlnGz69PlOKGOvj7NGvYCxzoW
Cxf+vnmCE1uQjVQEIjA/U9F+mrKGTKCODl+CXk32bNPYBwRa736jd1dGhiryZoDb
T+jKSGEFtEtvg+Kz7gGPPwBwT85oeUJl7LrVyZy23UoKntuVef9CjdoP8+VXyUzC
JB3MyKBbqqdfTOxfa8Y4GXI+7SoCmJ/J8R2bvz6ZotRQChNE7zptlcYMZNy3vip6
Uy4OWMHbqvUuEG9SWfq5jhzs2RBPzl1Vd043MxluQSQR66msy/JA7JaZOcgHhba9
26t2kAak6pFIHNqFWVx16h/q6ww7M0yv/qdn3SomXw4BiXlljyFTpWpHzlqzEVOV
F70I8bAoaY/E0MY7BOdrQfhBss2V96TrrSaBoJeVCNKWPS5MJFoGtUu655eoduEC
MOZI+I+kD1WtXlG8yD0S3G3zj69M6xP9bjruwK1HUc33/L/nyjByX6+CCK5BYSaN
oWB9o1SQCiXsp0R1ShsC4CO3im3TM0MuWrRnepT/8SyaFnyngQGoeNuWAWYAoLI7
owZ/UtKNY/vJ3xld1M4G1GnBQUuTHUKrvf/6byPvp3Jzd6rNnY85OTMOVHxOeA4O
3a9C+I00s8J3WV4s0v0ajAR9xOxW6XKwbTGcw28ZrKpQjVSyIIDZlJMl21QzkHOL
gc5ireSQdpEAR4r4LtybP4oCMYFN4rRRCT/Zujo3KfDq4NMSH80vcRtBOEmW90gz
kWD9pNMgP8cRX8p4nppCPhw73wa7v48djyMBFa5NHxSEzUebI2VDbj6as1yjZb8e
vns2BMpPrl5Z/WDgtgSHAHCv0ulq8sujfDjbf+tWDbnR9+Sr7g+4E9S7MkZyZ8cV
ro/NpYHWWIT32T90IZgHm86k24GQD7fsIEKqRfkdYxMTjzcdJ5KFQUV1TMNnft2A
qhEEG6AKfBCt58ICRASKv8KMLsoCEmfZ/bIsY+3PdqS0hQP9LtbYBWjvtPtTf/gj
2/1QgPIQUDTuEyJXLzfcm8J8VAktos86jDkIDJCkJjmFP4+cZSOoL3Y2WmdjWcNs
syEFL4QpHHJ5raZ6nEhm0XqpbEe2QNIXJW2tezsX8vLUZBQxuMAK6X6rt8du/DVx
Pr4lEWJ+e41etCZh4Q6tBsLQCPw4Nqp0j4KoCp4vGcDoeBTgKF0cX7HGBYinkSmC
9rjXKBCjKRZLbPYMQZLMVe2y+A+5Q1hr/NKivr6ItPbD6tn9wHCMLk5q7Qe0N+gE
YeVgCfFyg2mhvTNphOWjbncwYMy0YdDZIykaisT059D3jrV1J0ChVPup2Sq+q1aQ
2aSsGquHMs3oalz7h4tF4svkm0+8O0veUbtHb6jiGhQjHuZKIZNh4ljCZHzaAdLh
Lc/hV+cFaon72DIoEgscuyHPVQba7H0kLwMkEm5OOfWQNQQaBv9e7Bfwa73eaiEZ
JAg2xBXNsn7paFfpqn/oHOzjUrKDwgHU4vSlw5LrNR7PAbMXyK3nK9P7dQu9jTv0
5g0WmfoCtwbI7L7FkDagssXLzsQ0KgXReTVXGMcBkBBJCANmGPTRQpnYKL2xtW/q
9HDLU9CEmBmP2lVG5n3ybeLYk0b7hxomGYNpLXv2uhg9sIRLpdJAkwX3PHSH6j6g
KIGr4VrYvP5+moI7rWprnf7Ybh6EgmPyqt/nL4G9QpGvnexA9McvW1W/nLJjpz1U
Nh2pI8qkiTiukYeKYdPXZmf5h9Mp8UNecyyVHPBU1XmJdFqCaIlMWPUfzGnHDMFz
3V3G0+EFw1ckkJj1pohWxYkJodh+LTZKyHGgCgraUGNAX4mrneQfjqlzKD9ZijBn
nnpltlpoqqOumWjjU7MJCQhXyG5axCk7OY5edXzcwD5oDi/zhIry2U5uvyEM2+SB
IFtLIo3Z0D7aaUlIjzdq2GuFUaAWM6ZWXrP9FY2nua10EirQ/lywji8irGXGGPeV
0r+Rsx3HDgipNCaFrNEc0lev1s40N9Q60ROmkOxBof0m5E1TpdLj9vONe+jbeS7y
yWMfPbSG4+OuukZP1/bSHzEE8RK4PHvdQe/Onmqf1OuWcltqhR+DoHRpVK98M3Y2
N912coC9NxJRKUwIU9cq15OXmzGuBNEHxSgZOp8MykXargIfNKfjFAPS6wO4iOVi
kNdbtwFkVasWdDZgm4SjiBA58P5DUOp58/3GLJvV8PPPvmk/RmIvYLbl7TGEVu/q
lVrMn72LzmyT0G1TzZ4PN534ZGO9e/KraAqrekMOiLxkkT9ptJgvXpARR/aL/Hjl
G1LyUa5g7COMlwsF297pdEDSOAtlC/Kpc3TshgtDrENO35VVciZHd2T3UF6YKVgr
fWXDbhjpvOPRTw/zxh5Jr4PoULFqobeXQTRC6+c/6QIiFDkjgWHt6BkjlyHooTMS
Mxw4rxcy1m1zxRPYyJR+TY+QZLld1WOyiGQ9q+8sshjWcy1P12YvNG2ooH98FZRk
OmONln2Zxc/Iu4xmTnWKFnlXjZKSPYyWnhD2i45OXrL/0+ByeIWnD9EshAQXpZ78
UodQ9QKKjtqZnX3Qs+AFVAxwaALG1DScVOoOJ/CaFfLRpwNCJ/hS23MstSsR2T9l
0atNRxvDjDw0i8SuzRZ70hDQe/8ZSW6o2UO2GAWKicgJwwVJN7zbwdYAUzGlkvhd
YSxlwP1dSmQRha1y6TpJIceUk9H2bvnDST5HlIUIGjT3qQUIXUBH8OZP7u7EQvgL
Oo1AUSy6tTYpGaFQgGbtT5HQiRqh5S2zkI8zUtkF0XCZZbgvIhKpmMaE2+kCYLCz
CwHp0vmfzsYIocKwEJvU3CuFBtjXdM73BZEhlezInPa6DRK9FdJ7X0xAK27ynRqg
iKannnDXmgkMSqqAnuutOSlrxh6f4FT9QERzr9UVfEpmLOZ/7rUZ7uHoHy2ESSul
XiQ8UyBTNpGYyRcHrSpqt7nuEY6RjadUJUlzoBc9KmjV/SiDy7xZ9x/9jEsUmYmY
siDI3aFmv4PrkRVyCw9/wL9xYXczS4T5VNx+gj69uxXJXgbQCrVjo5YxdTkwQsr+
zAAB2aucVbTuLm/GSidCgHa5hDNcH4mtGvBt/LFJvy1YRzhii/vNUjUy/SS9cGxn
AyubV3rn27oCFIodyDxfQen6O5zwhE3Vj20DWOnECN4SyBbsacDet3q6kWz+ambY
vxyGZWgnG9UOaq4XAhduqC+jW8IRQWfEfdz6uo4sc+wNX2p0RxiO+1qryMz96beY
YipWJQ/echAZHodPGozppmIUY3Jo+ep4DyethrJw7z+Lpz/ybM18xUT1+mGrMzC+
Aoi1zT3DtzhF4gA8OtiYq7cctn5rJvThHJJw1YgL06zhofcOCssp7NsN8Go26cyt
QqiXHfij9o/TvC81ap7tVEhScBJKMR6kDshZdn+VSO/8k9qSwJSlSgMFstK2e2n/
7wPglONSfskXOGkpmNh/sKX9iSjK5r78EVhnW3lH0O0UAB54+A14/pSf0i6BxlJW
jGr0nERUG97jmVZyZUyCbyaSQROKXVMUgtqRVucwAD3Ato21z9gibU9PHUmGK9C+
+2qeYzklfZO++ISmWySf5grrmWL8ZIyH6KdCyDvzfVZQJaj1T7IAobFFZyykRxAi
RlxvCTNprsJ0CRZprX6X/rmlgFYys0EZ86LVmBi0At6eredABXDJD/eVv/ZMDjUk
ulE0JeCW4j26bA/6HOAyPeKsIlW4OKNIhJzKK/nuCbcGQKeMtwZu/K1AxxVUbY6E
MvS3xytGCaBmWPQVUmqLyrrIMMaRf4x2yp0cFAQudbumcmLAIj1OYFvvHkx+s3h6
DikeEO0Y/3K504d/wpo0z74J0wIkIfjzrDNXWeUJdi5KBWeoEUd4qiR991ttZ/6l
vee8J7QAM0HZ9bXLx8lpOvSPRYu3Rl16tv6P6AyxPbcfpoWaxKx/nmuGTfIdpsVE
kQ6IqXaah3uT+dV2ojHaGVE0Z94Lcs8Z6z5iR/lKiLtbHLcrowLjjP13MQEsz85P
LuyK71BynMbzUgn5hdPWxbvly94RsykizqQGKiMwNwlwxXyjE39yeeVT1Nd2mKAT
IDROIrYfpvpg6bhYZMjAHJNwHGesfcyMSwcog9jhF5M5K6W+6kfg08MFIRm41CV1
eRPBwtd0bHYxc8QPNHu9zbkykIb/ubiXuQlLMSgfNxmcwgZFRZlhog8XxTheFANt
KfSWvfms5vPDdT83hEZym6y15qbY2dMQUdy+9F/Krfb1pxb2JUfh+LrGPcK75z7u
rmIROBhVaZ+4ewVBhxlVssG/w8Gg0RACU0RFNBaGDxQ3iDmLFBH24Ky61dEsAll+
JPjtA8zw+KyYO5k0yYn+sYK7BZA0c3gqPWTHowmWHBaWM/1vXc+giSr34goMayWE
EM4CtRkIG2AHdyM2gSm3pXqDeyYRwwUNLoIMjIL40NXY+xgW5diH2PyEaxMDJctW
KOS399JRejRFZq9C7jVFlcIbGrBDzWoK/ZeZNdItLsne/q7wWR0xOZisJjJUq/yi
aXEFdplHGE6JMQ2eSnkbI0syPSTsBJC1TN1wWCphPLRCmwpL4eEg1gwNVOzbCmfK
MCt4lrXO+ZhP5+C2kOA2YzMJcoyd5nrGfl2Bm/m41aCMB9ftXpSwtDV0+6uFVbA2
409bm+FqD6qQcR2b3eJscr7PSwhWcKM0Ack4OOqoRnzP7/+m14sYWmfNtkg9WPzq
0Hb7s/rJFKtrACZwQ3pnD2ztsvyk0HpwQAYYv++JI3M1LP4ZgJyNnkJZLzf/opyg
Ub9oRKkTPXJffMKzdZr1NFdBzzkuE+XQdHenbTVSyKd3U1n7naUbzbTEIIPF6b9S
Z6Ag9OFaSJtmB32Jj3vYQEDI1WJp+X/Y7bcJ+DGTQSncfHp5np1MKk/iQfIsgfKW
1uqwb4sNeWTK/gwh/zZEnC6uWSxZLatcTNZcrIrHib8dFjyPZXYCAiv2l85QuQ8E
cfHgcwz6XfdxKh7txTrPD0/kT7NfEdPQFhci0u8Za3inl5tSSLqMCxYZFUmVlCkM
LTvb3UX73h4Jh1GZfO5GRIc2nuLWo0GBjI9wKkIM3UuCVsmkrjUeCKdEt+7zVArj
kxrZ0gvW4j4yGCyMt4MG1BgX2aM2BYoXFEgOrnR9ZzOOSXnfY8Ip5+3icgMMhBBg
IKBgLI/IMelwFrPKlhD1DQUFQXPYCbwybVnsju/+0ucgEqm9s3tF4Wfv5oVUMCve
n48Q144Bk3SmKrrmP6tDHJNoexq8gJStPaSGpIYElPwpS9Ahbpb0HmOFdeyeuFZy
9tQ0MkVpIUH5MA3+h8qNYyl3hoH881DkbQtlRJlTCvmDdeQPDIgTd9mNhOqQTWDw
+vyiQ+6ukz3AFv0MdpjoORaLLxTKuZcHwqjy9ocFSfQSYPLiNN6GAL1IvVtS9uj3
CEaf1Nfm0f5R3aaxqeQzWBYHTgUapVAd8gj3cW7JtxIBkm/OdKN7thG6R5FmW3uX
M/oWM4KmqwvkBIK0aSQ8EL1YjRmyWN3ltSdttktllgBI5xEUnioWdREu6N864M2T
TF2SkXxDJWUrtov6TqDkCKSxZSX+7JQVpQU9q9ZWoP5gNdQ85Gp9vIi2SdKiDRuK
ZUXwHyvoiIEMx1MrYRs6gVTzwoJ97Y2xiYsvIBZf/QBfebl1CcJvc73NVQRWYIJv
ANbZIjj0XhSh8oe3aLmgOG7g2oZSa4lEnspza3qHGht2cONJrX3/lAm97LnCvIL4
ShpYeuJWd4FP5vwfDS7iIvaTdTXLiUlNeyoK+Frr9Emo6JG5up2cRdBkU9+DPHIO
aRMo7MqaIjy9q09bm3vDMSEeBCWDikcFYOViXdPzKmk4OJeCNZG54kVnJBfzxyKp
t0V9r7jAf6lFbg88QzxejlznHsB0INrGZG0AHILbCr8IrmFRX/ohfVnVdvBFo1Px
A2QAE9f3cp/a2hDA5EiYeFD2cY3WjylLnVXYB1rAuuIwaN5Mb7z8jPev3DXit1s0
6ZLJ2KhS7H3CbznQQCq0vOXXRTlcq9+MqFQeHyVWmxHNyWPjhXEqKNEPmmQVhBDV
IP5wGXHL2IWzj4HEHzrKGLvI8hqds3muXHd+FoTaSMc7Rs6pbZ5zRBgxDkmDDCqv
DIesErQfwgNkWAOQo+VxBPmVTJCEKHeepOjJcygaSFtdTAoByTxL7DL+fy8EyR4D
YeXOKqxB/LyftmjMysJhOf4Yuo3A37r7Oo2KytYMe38GHjzsFNRMNdSsfF7K6dBR
zm+ybs4Sz3cMOd16t0sWssHwQQgyui7rjRtEXnMYERa4Vhy+b66lIrhEV7MYj7cT
uBtAXFP1kSpiBnBMOolOBFktFbE9pfCXG8boH6kGp0CMbXv0I9i8X/Cd0gcBMOI2
bW0djn3YNxpzID0XaBFi7XRQJST+Yf9wDzhGU5er4qUy/V/X1qAJzvhRrGqgDNUH
tTgJ/YF18dQdBXmULVSeL3ChnJCY7dBaKMuQf9Aav4TUW9wZObYFv5slhOeREgqE
jWAI0cbaECg8tNGm+tTT6TqziZkmdS0xz1qQO5in+ug5ExE1fMhxd3NzfXOVL3e2
Ig+zoKJbHv7AbYegTAs1oFY+T4FhpNXVQY0TbsESGdnu038xhJxQ82EWWKfuhWce
ZR8CTUiKrTqCzMDcveEKMcxT4AlHSpp/YhNtElme1OYi+n1lTnDrsg9c61Ciz0CR
zgQIbVbNFmfWYkHhPiWKsATh9eFnt0Edal1dfjkGuMlR6+MYvRHR0ANoqFrVMEos
T7Ki7gvlF8VgNDOEw7M4lPO1xDZoPT13VuqT/yFupKGiGngMSx167YHuHbmrVqi1
vWhowMJWIxCbhANIf7+WQ2caQwE2QcgCAq580klaxfl2e29cxnYXwUR/lTWmAVx6
mdnkMummQr5WaWPbprTKmDQ97subqJeGbNH4lB1ejCOyAZyMYaTzg5dHL9RQwl6E
uylCZ/hjfkxdDX9jcsLbQCMzXeg20v1qWUsQtk5O9f2sw/0QMrGYX2OTRzI2y68q
8UiD+Zn3MdcwsIOp318YP3cF+aHSo+7I817hD+puzK1NCDTNSWybv+A9BIYRE33S
4JRwt1Sll7ro1ajZ2l2VfRSSPGFFNVMp7yYwBPntL/j/Zkc+PEaJhGCulc5meT1Y
O2ifSoKD8SSWR8/KQ/cvfH1Y/r43oZUEaUOevmTo/QB4ia2cSC1ychlW5IbIr+Z+
F042LrW664ML8cGiPzJmq1oYlSR3TLXiLVSoFTDcEIL5nAzKWEEkWLbAtxG4tC0o
zYAZ/9SSQ+2NGBJK+QWPE4uw/JQ+0WIY3NJ+anXlGEs5h9TLC4gg6+vTPLqARdRN
1WPv2g//ZKea7drbX7l0aJcAbvoQp3y67wx7a12CPntDtQ1YHnmFL0b6mNVlm/IF
bVnRZYju9zlihvwZrR42eIxVRWeW843AXgXLZzoj3gMgNqQ6wwhujTD0ixLyrJFe
WGu2SlUp7iFWXcaDTj89U3NjxlOxhvsD0UiFyAYw0yZkIgxixQiy6N3/HiBEUzh9
dcW2LEaUzOBOFt7pBWspwnW9OAS6AZC1qilclojzczJfUqbfbkE1vFs3ppnCS9PN
qoLZQ8krbVlbcMZ3gcTLwuK4U3TlEBLxZaCgmbkDZMijOTwHlvVXfnBMEEK21Oia
C77BakKGytRoUoD4vxLXfa0szSY/8hc3IJUi0IV7Fz4gniuv9hRpnBJXiPeksnZ/
pvUIx8VniSq7UZGkIOi6BNmoWGTbf8f5GCfyzO0TBgPA4xru7VPn1DIrf4Zp15Xn
jUq6wO2c+NvBKp/w732RHTzKGRy8uledLoY4qAx6bWtvZ4NLc4fD3gVp4dHPENoC
/CaDlVGu0nbfI5Irq43ndhz0WnzmqM2H3RI3b3CxU+HvNtRHVj1szv/0wXvSR+ic
O95moA8hXsyXA8DSFrMn1UM9l+zvC3QkuqnG0ichon0iTYzcywygjeRaHj45Tki4
PWlJiL1JAT8B5I5J63D/Z+qxl3OmtqYM88u3cZu1l5SRj0YNfaC79DxsYw3I4H+J
egUQMLIqZHIgA3vFmTuthLykOwZHK7ktH+j/Uk5TM6+Zw+4sjtrLVjy9gLZHvfSm
repEAryjZ91rNomFEK/lGt90nfI83A1Q0kW5eTfkmG5p7jwIEQ5nM1Pdi0rJDabh
X6VjWyuQefIJmCbynogUyBIWxDsGG2VVsmwsnXIUGXRrxgfWUHAhs5CbWAEkEGEh
mrV0ZtLslsK66wohV2UgD3ncSl4vATgWtBmFfYvDzHB76x49SHq2+CtVrrD/PZI/
6A5Od92R6r8f9wxBBJZ0n8azXcS4BL+9P7yel+KyekE3i7Q+DUzXv1Eiw6/KMv1z
d3+6q2ufc8jmO6h+TE1wpsTIdFMzv++cfzKUBjbP9adozIkzUCgnKIYSckjHpuyj
PS+91bfNuSBbugcF6RvQtZHvbLj4h4f0Cu4YZ4uKn/wlnw13eDJvbCa+L9nuBuD2
QgGRcATvJLzjUaVXujz9REyX3s0zv/HeblDl73hk5aGjacxtn14G1yO1aVHKRLKE
izlaTGxurX7+3CMxaJ1q25YVO+vu/02vgwmD8ctNpeGcaRCI7bY7MvkDpnjexUlR
lDL4atmsb/CTznA7ileRmPcJtBi5pJpyzTRXlmsQv1yro2cnlYh6vkF20NCRbA2d
J6/23ZbYVZ0OiyJ6XcM6VTpHgyY+2bsV0/n1/1QTUMVQr8nE6A6LYNXRV7I/qVdc
tYk0NLLX4CUg+7451wFcFwzV00VEW168SxebCXybDZGNuLWAiZDcfymJtDEAF2LJ
n14pq5tLDeug6V77dgIP2Ioe6IxrB42VOe6A66Juce/2SqQgdCGGNfvfGjoBhz+7
V7otDtqR0531pDgqdveMu/X2vYJ+Bs9SpDlEXlvqxQxRPapvZ8tBlKkstJLV7xoT
xyoSHzymZ9kfvJFJFf5iifxgq8VvmfYVQIMeilDdS9mLcPPhHKhx3TK6hPNh8rp6
3R1B2pmovkuGBDsuw6VZuhHaU0CE1gdbQWqfGopgeKbFPDDxWZeGiwtpp4YmK+b0
8Qo1IVZ0KZgV6NQj4EM/k5xGjbU0Ftm6Hs1zPssPCWvGHeRsVOhui8IiA8Onzc47
U4QDXPtgN8SORQsnp4oavSoBSnjbH6f3nricpL3ZUls3ydUZhlkX5OkedZltgTF2
NlWJuv7kiSlwNeiAgM59tL+3GZPRZ4E4EOtzcdLkQQ0ol+OTlk3/0FlK24E9VLWE
jjOnsD5BEK8MAg9si5RnS6o1j1YjPd1dQ0JVBOpBF4JAYnIpH7aRSu3hea+bWRZ7
uOpggs7dTUoSrzTeZP4H7APg2u7mONEXSe0vRMIbo4AE6P3yAV4Va2NIFy3VDiRi
rWgGWIsJaV26DZxEeDOpi169BC3G7gFOgC7VKAc+Q4agxqazct6T5Zb1ww5G2lRU
wNxMJazwXvgHVlLVzOxCRy0UO+foKUifnJnLPKLggy8VQBKECGETP4mG6LU1nDyq
9Q7F8Q1GuYsRFK/wA9gd8kDmB2xPIhfRgsttfllrku1vuBqcg9Zp8DtsuqzlraFe
xE+D0VCtrbgnZ1wiBUvwBh+XcAprIWb2d/0tybx+wDIz+bTqoTOlRZNcQN/1nwkU
JLA38FP7cEuOnFgd0aYRa+l1n1wTD2Q1gXLDcnwnbydN9KWpXgJ2WVlD6yoYUrKz
gWGVgb3ISb6Axa0bcu7qI3zmiuAqe7LhnXK7NgkbLLVKL+JvDky3niG97FTf4OGH
/E7RslB8GgH8Fhu+Si0S8MsUJ1H8jmkcsg5kTM0ZHGbWWEmazAB6p3QUdoeyo2Yh
lxW6Zvv0LXLw/w7XnfwIuoMPeVqYAKzyRwXhakQN96upVYGxQqKeSsxJyZPF24QM
yc79IaEIQUAAGsqamt4/ZkzQzOvfEtO+pEI12TxcaYAY6LIXIuBy7uIa5GuT1Crv
eX6DYqSXzz/G740oB7owdJyQDxKvLQFnDZj4mx+z0VkjV+OwqCitMKPg/LWqbTax
LCKOKVwBUNwc9KggAPoxOC6kVfulx69OSi2DgwzC973ATqKBibXr/8grCKGtesIQ
xrc0huGjz7UtaUIaNaBXbj/OKp7bjr17GV9Z6xgrvwXi+Sy8UqcvNgQtM0SwcyGk
cY/5tbTitFag65Dz0Rlre+sQMe0EJWNdgiqFRxK5Q5GhxjTFiDP0fV3Q1qyoITXY
Y/iHY46rMAcAOIEeYznmkMsd4+uR5/aNCKc0pj1fFdDSLOnnvVmyePHCdyqsF18Z
il6vLGmU2N0uEvwm3ZAzwf52ij5ObjJriKRV+fRrcDHiXiIyDG6jkjpQgxyTH4wx
Y6j63bfQUPxtA/6hZ8spvYIlGVx80Z/sfODoD2Cdk399NZZTuThvzqcadzMoeyhc
PMDNIM1qlzUD9TNg/nC3/VApfxvA10qvMiQbTY7iSWnq/+KLtmMCTm5ZFs2jnYsR
IzYxMNhuR9MtBhBFEY9PxFnvpXtRq6t4I4TEeA7En62CJvm4G1gyqVxKl6W8uDtM
3yasNBKS2p2J/j/hJjZdLI/vLxTskRFaihCAop5ZaFMyY+IwgWjLYPN9GjsUtz5H
O3d4seOBnj5Ovoq3+YI/WzUxhGRtZWwXZePJC2cQNQQtvNwZyC6+1mXh7WUqG5oj
68yz3N3IiEF/ZSIzpuDhGCqJFVbl4ET8jJQOBQrEkScW8o1er+IjnleiPFOQqMXt
Y32Upqu8UgF6FuBn9JnCtS1XsYr2nHD2abnGTjvGDHMbgO325WfEOAwN5Rz8i/wX
ZM9qmlCSbIb4tOZOgt5KD/zs7tBTZGQSlPhwMHWks0fWeE2LXTdhN8Jy45QP+2nD
d2h+UeaVfv42tp7evaZzJ8fxwpXdV7EklHepndfJB/MPIfGvmWoRaxcweDznDYgL
9yiQVrNnyuKZDiRKQFcU/03uivl976mJ4qCw9qkTKD/oJIb3sjVkM5Fm/XMMBFfi
Jpo5CAFTDo+uKM/h8ABZSwr5ZtpoitucFP6DlRWYaiXoqwvZFiiGiCM8dL3KlWRL
D6QAHmfTQU45+hrHkRajeWw1wTkP/L0384QZs4GmZS15r+02H88sJCFd04VQ3Qv5
Q5amQGTFJIjgL/hlGPGBfaGs/HZJG/gPeW06athh8OnF5ow2xjYiN55enJ3A3Mcd
NbYKQcnwMOHOtqsFzULcc9OLp0zsTGzG1x5Pl7/tT8qMHElGA+y2I2xJwM7tPWAe
I4Nr2vOSO2Nkui3HqJLjnsLEKipKPfPpzS2g/Xb5/qBPYGFqVTtHoJEdSmg9T+Cq
BuTQHNlGR/oAYJSN33PmplxSe57UaHACygmmFN19gNxgh7dytqCXGy0+ITr53J/B
UdCRG+ETpEGaF4RoX8Xj7e1X48mdruntiLFr/UZROo/2YqUdDFs0Q0THsDWtOeTw
DDbBEy/mn0lRcVAQsWcyyDXKzFprNzToTNtABSxJDUuzv/L2UIET/LeH5+CObeH9
mY8g0Ej7Iy3geEK6vu8dmwpi/WFm8QRj2NAHd2Jk+EJN5odp1B21ikkX591nx/Ff
MvNhLUnf8SewTRUq9KkChEPSs10AJzNS7xjgZdikdCAdjIR1y6iPOeH3rIYBvm8A
ikyIE4G9qg5EAGbBa6x3VbWy+AgOtG/zbdp/ftZl0NfRTVxkUBHFR808PukXqBET
3OS5xNzD6CIS/1lF1udSByYXMmY5S8I06yVLWTh76fdjdZMKjsjDf/Np9WqtGEaY
K4xoEJ8daQlLgxVQnVY7EAokiMPtbL2HN/64f/LKdY7sxFyqEW3w76OijgxbMTVy
fcTWMV2NubKEIQiwbSdtsWHuzOfZGFlvGjwt66dQ31yKGYiNES7Ohlc5/AzmvFgU
ifXognCAMXqpuIhs+uFyQR8JE2KhpglNU3Zi7KqCFGvqu/y+OWxi8K9ar3nL56f7
Ml9snBtq30u3YrdVFcwQEGLMK0qukzldq13wGNYVucTBFGjEig1H6cD/EGlfg8pp
VU2mcgwMi9KYHUAsOdogLzVUWffVmo1lU1gZl+vpB+5v6IrOUgbJruwbVIcgNB5V
2dcbgSgCcVmBGxukQ2EViTdIAnILae6R8HYo5rv2UD/v/fGp9UhaqwejG41a6yHx
k4Oq6qkRH5OWch7S8hLG176Zr6PLglF4ama5Pmu7CCXjwgm0qp9Z2BNyzIXb3sEI
psFDsr94gXD17CG1hmTw0HdtuvLByZI7AB16kPQa0bfKE1ZlRKH4qlUgw1CkDjtV
edb7riSyqo93Ix/5GDcuyEBK6UI6HTnquHofLNdiiK3O3ei8OeD8f/He3YntQL9i
TXwvOAQsLrW+L74gdQpcYGHEiEhJrJF160dsGjRStjOwZJXuLhnlv5cau5YXN5yS
IuY0thmq6jIxt3K3QWi3l8qI5nBxLbTj4k7iO7MoIrMru341Bd3COa5fYID0MkfV
+IonnxZeR9P/6yhfJEyFPVIPcHYy1+mb3sFOsi+mT46TJgargqoCQDHMrcJmQgzr
ln2toF3Yvbxe/Jyw+9TXYxQDWh/nGjH90xiZoVzdotcwsx/ShwzEtJzlUtktdmQm
f64s+e1lf0ZzPcKJhwGa8b+i+mt1p4w7bAyXcyjIC9ED/E0YPHvaPsnbcWQ6seE2
2/zuAyTRpK3KzJFvDI+YyhwsDuyaeKXUKiQmDhLA2DRY6hY3W33OEvJYU4sekYQg
TUNdmuogdRnt1YkPxOyHFQt89UW6aVWE/PApwnOf83FM/geFn5WB126DIyjA/zP3
TBysGI6fbVf7wiOU26IiY+N+O0BcxmtcR3ArA6dZZU1PN8BlNe5jLDTbEVmopX1K
bPY7GUNuW+fW0Txt2eIucTL9EnU0zpKQlKFmHCK5SQqZJpPWneV6EJxGJmZrEKWD
NYT3hlKImTqeEcwP29occ20hDiNjF4X/oG7ba7X43UsUylQTBx1g/E8NuFV06Tzf
2ltsDoaKYI6OqPU8J1KHS/wFJQmj3lhQlRP9eRHcUuWfSGKTPRSkGT/Z0Ke7DtHn
fbvM32c+sSeEeDb4OcbIw4r1uG5PjCYz5Ru58hI4EiPyby7nT0dDoeKB9eQ5huZq
JRdAhg0wRwvathTy6MmUMiurw6HV5FSRb/Ulnrtz19Jy2Rdg1mdKt19r5YjVFxdr
SYXgKNyO4n4ia5w3K+tpEygIukgDQG1Upho79fHjqynTinWhQcfi0Y3L5xYICk0H
JKbzNmdv8WhN4HCAIZxhdBB3sllTuadL2GOorPeenVvZ5uIG5LQgPgsrhvRXO9IS
aXzyWHlvVHK65+nESWr17e7wmQ/Kjm0UtPlHTNP+rQcOTR9qn0214uTgEIVnbiOm
mgZTRO4FYEinqevEbioKordPEiUb+2ML943pVWQcGanYOmd7r6ZfoUw99VKlGbgm
VoH+22Both6f+YjBO/feXIkPSwF3/EgqJYOIGSIF9km16Cff5jxTmhXavbf17Nsj
e3gKihJ6oJzE+LJjsa01GKdMPBn08i+i1rPgS/4w1YbLp4Q8YjeiIlXVy6wGgznI
sbYH89mIQF7ocCm05/gnyCrB+VGMdUhYT/bxih/Fum220f314oyJIFpCvTgOkTyZ
Pzml1q/BXu9xF2gPBPyel6zvSxm9ToJ9aVTbibavQGNZelGixNO1MIqW3heHZzId
MXSKg6kSL1p6hHWEL7IDp7856HM3pzQFSbJZcKejAbM0W4zYFpG6jiqT32qAqL7Y
qh6YvGjWpY5XVcnLPzkoWwJ1RYD7xry/0OYTRzv4Dlxt0XhOloI2q7/xj8PRVZx0
mteyJZ8MAREZN4sRbrZGYa5hl38BMlxv3XCsu0TuDoDq5RKK5O20CY6HOdn4+b2f
z4BGps76Vq6AfnqjS10LWylzH1042/apDv7GKfBDQZg+KQSUXXCwrgbJbzB6AtDO
EfL97iwXgvRT5CPJ+zgqcZEOFqy2vO1T1BDDYl0qS6eak3iPjxOOIwGg0LaEyPxH
dRoyl+b4QurkivdB3WQPQ46EieD5RYfKkIiRTcz/mk/+jFfAVuXd78oen6Dae08t
VoKxlihQ9J/wEYZJzv7V4zflqf0MKxNhr3wdCsd1AbD1aU+w8OtJxS034F/vhWW9
LfnUWoTiYyu2LQbb4/xTc+LW9gqNqW3qI3XtEm7eb/ckX/6HsNnIyr+b19ZDIqon
ndOYQLNcQcY6Ixox0X+AzKC/ZmYOPSsBpXQiRYmPu6YgVdUKCDuwLgqbNBMtZw1q
TVhrbWBtSJxoc6dkcZPTvOkoCGKdBZEL1nDWZrClkaTZkDQ9mX98vIiBrxxcAcd6
iD9H4WGaWze/I6Svj3uEna7dj0rEAFsvhMlEss/ukzdlOOV4u70o9r+oTQ5CPqo0
jZvRloVP/5sJW37h3FyeHJM+xiOA0OapqWtrFnmQmxzYKDt7ZKzq0eykpRkqNq4u
sMTKEs65227ofQeRDgwX4e6hDTe1YSWSd/hS1qqrBVu08iCZt0goVXdNmfKNlZ6c
YRguGVetKAKcaoNuHxUMKabwTdPQ+9l67bgY8/MW/DQQ9rdLVNRpJnwA7YMaAgL7
PStdOG1dU5iFoCgVtncueMtsq382fC2YqSs0dxlzH/LeZcJDYmWsEVBz4feWE7/l
6BiP+ttpWiGMrJ6kWtRr5MOqFmznwB4yMFB06iCinlToKi0whq4Yd7F86vgUEeqS
Jbiwqpkhc3ooZ0yEM7tgmKZi9pzSiNenn81tLg6WBbCaLI6vBZ2TVbSaQkC1Il72
+CtqRdXLSOuFDHIsUisdHzkWomDsveozgMHPsEhvN37GyUBWS9p9z49bt8IQT45t
7vbCgOjv/ICxmmTrdBodnQOWqzmco18M1EZZfWBFrKd79QZ6tr37hx/ZOHiyHy4n
doBs9OFKvxbNDTuYutURx/bfWsRoSpeJJ79MuEFqvkVcuRrfwFwWnNqDnHz5uw8M
sXeEvoECQN3udo8Mns9lJ2v2LkyMtP3F0qnt4h76g4uFlxEFC9shg9exoISsL5xX
6iAanE8lK9K+8lUeNna3dX0vNvDsPxdceRfkmBJW4c3mLQi1R94IIb8RIkswp+L/
qAFXERDtU/o6v4wyEFmPEn76ijRZReMMykNbH/IFfCvDTcOv2RsyLIeXZvFgwgxp
KWz/Gi4xsK2YRDs79xu9nYanV17kKIueurk8PbnnneVVz+P6x9E7UcroWR1mpsq4
bleO+gnLFaxUXjx6GxW8UNW5LC95jaZmp1G7qP1atQIhmWR1LnlHh2IG4h/MhqtU
eA8Gujw9ODIW4GexAZe+e1Xg8JlTAHQOjdqeKW4Ab0Uix0bafMXJbyjAsFGWk0ho
84MFHUIxT6PBnQnXY/fpB1WU7L7z/sfcc+2abK3oqSefcoXUlEdvnHPMcUk/frNm
IazcSD73ajkci6MYHQRUMQDD5cGpzmkAQiPKqOBCZFIjeruhp/HhuAHBRSy4Adux
cBTMrlCXiRzj4jSWhPfm+zKI+sZLd0h8HbsZjS4Rq8F91TVpyTG4J6igrzcwWvVN
pViqS98xCSSxtLIRzwsMVzx3akazARo9lvsgL9e6LW2f4iVb7q2mFdcjtdshkHdM
VvZZeSzXiuIHuKtQkG3SkICwf2QepPvzBPzVnAil+/qQ+17Y/W0RXzeisK2j5TB1
N5oePce2VEz/IZWG/ybA20Yv1lpoKMEp8KrkID1994qMiQsGIlj+gr0SWEY9LiS0
auV0CxI5JGZYfHbhjhmk7KLdmgMQ4fkoZ51e/Qk4OmjjV1I2xAr4001Muxc+iLxR
2TmLM4Y43r7yV05AgD4yx2Sl2En8QsRMOWaL+80rlSp6otvAxEueEUimRnbbP9m8
wYdhsZmH9GNmPRSg+csM23Erab4vC+PqJJbyMYvzsQgmboaItvEGtNGFCYbPjJVX
zkRlkeebzOEUnFR1nc3LaxUZ3m+AMWdvSxI8MuHbYadft5AbuB4F49hRDO4Uv8Ot
TuSXPKMTdLpf92tLmfjgnKBeOqz8pExadZKd0jIzjv0R5RPqJSeS30ZFXSAnbuuT
2/WP/OuR3UXglhmll0h1KoFQHVxNu9/3PiGCRwx7cEr3bZmuwNvuEDNjhVmw1blX
Z+I1MO8Q929UTTBVu9ur/R6NKwc0sNvn0s9xHCPbBQxpWI0uJLoDcUXT4e02CpA6
f9QYlLsijbPQ/QSeVBOKZGPbtOYsxplXNSBzJ5ZgjO3MBR+Br65Il0XLmNdRDARS
ppdA8aanOJk2hLM6BGNUELPBD8A1buxq8qu6KUHRLJdFipr7X09O9+FXpX6hl3M/
tq3rXJeJo8yIPCVmABrbZcfi9uAenULlYNbzxl+AWVtddBjIa45yYrFtDFZFugp4
etSiBmgEDxKQpc7aSplGb+kwDfDOlIULPDzuy9s/j4vExx6rc5v42DIP+DmE80/4
dvAWc3CTYE6ZBKlXD1uhslMQ+MR6YW36jZYJf023b8ysG4O3e4zCggOty+oXAHNY
m5We54CQvnG7FoqRE0JN+FIOBn/B5PaPY70wwqapyBTXMS7/NQoa7cc9prL2K79Q
9PcER3nYOZGVmm2Bg/1IYI1wpVYnFbGWC3Zgz1AIuW81cel5H3JGFrbf1rBGHc5Z
MM7JT71bBZb3SyjCLCIkbBKGuQpziC81w+5oA+zPMtkmiJgho3fy+Trn7e6s5Q4L
QHR1pVaa3wKWPclh7dE693m62RWdnxzFthoHAGMkAKQM0zu05QdzJDIUFCcUjy10
nWsqe6wdJmexBHXwHoA3OopLJhNw6ffbX6p042314FiGfSm8oJ1wtptHAg2MEFnm
P63HQrerHENZdjCz3CfBsQ4GAPvKYb8DbdP61LfHaBVhjM6ZaEaRv59gvk1AgT6+
3TPHnW7aeo3HMEBrJ3fcYNnlnoTYIljw/oYfk3rAOXqkYE5tO+HOwAG9jgZCw8nP
LDj26rVX6M0Vrwlxd840bjtNlMSp0uJfo518sgr70ADQuRCefMHcPvj7WOehtiOA
AKmJUmgMvalgzEDe9rg7aTl9JlIAAcb1tWiNOv0Q0HdZzJmO2ZgIwCcbAiuXCIUI
g5Zu9zREC15aZxnjWZZpWgBup1+UFWWl5hjLg1ujKsOVbMFmxV6TGpuD1HJy5sQr
3pl+Kkf+NJzGVAafZ+d/jAKKBPAB4UcwH8dUKmxW9M5RhstCENm1W/e59ChJzb+P
tIf+9RHq4FVqEcN2u4+qOfdW/CQCvKDDa7rw4tT3VEyaIPmDdMg4SngOUG193i3R
IXAwnrnyEi0ZlT9mubtIcAI1x3auCzwwHi5wl8aIMb/TpYLM2FOwMpWFh4es9RC2
ahGpMuzByezrF6C1qPNcaM1ME4NsuYS8Ra68Nepw7v6bU5/Y5vqe0ctYG6fHmuOJ
3+gd8MA2zxm8hUar796tV51x0M1S3sriPhrkIg99WSPJImqAA5X7pPbxTdKG68ZB
5JzZAUIHCRkM0Q7vMFsk8khPFmwtTmZ9JkGjJJjycuLFMlb4GQZiNH+/Y4iZYAbh
gmDB+5VtQD+JmhCbWVYxTUgjSDFid9UvMDI7c2QeoayGpy8XNDETt7ecSV2Fxljo
UJQswNAMkh1jihXMSKeuueNbf20xjRwcfpm4aGMp2+UIP/14wFgeH94Y3wFdyrGe
7NzBHEgclLJYn1cNx/PQnQ5T9jldMSamW0fuxD/UGhlHp3IRWzjtfSRQLTpxb4X6
7AL5SiWlJsTmldeMvbyfn/uF9+l5sAo9HxOEEpln8O63WFVqvG5p/BvZcRLkJMeE
9wvbSeYx56gGbSKPIC6cGBXZb6I2vWsW4irBM9NxmXG4Mfb3cuzZSrXdKPMAJMNi
zoRcyXPHoPLtgBsQQlInydioDKe96yQePC06z0I+qlG/kGjQ0KsZOwZjPxJaNGWh
8FI5j4pS6WK58lmCIILDdFLcyge5stpWKa0b+uV89/v3gxn8+DjuDmt5+Y7lm/ta
yZJ9eofcvvhka0muxKmVlHsJn2cKSMBeKJ1mmpYD1+Y5QHMnpPtHG8t01iK1E7rJ
4D/1RUuCwp0CBUTod+cmQLoBYkr69Eapss2B4ntHd+/lCwngEL34LKKTr4/0ZKAG
JOTiQhSkvWUlNEeLSQlAxaDmCmXWDOmbkRPDdEh/K5pe0xaSf38oo8mON+qPZqA2
H7IsgXLfMpBwriUjY3BHEBIUujng5QLbVqkKyh3QI+NClz7oojCSTYxFJNaef7DH
yLewqhaaQB8QzAiyiu5Gw8+81p7/7JqGSaLCvp5ghS1P/inLr+/3/vwLuw9eWGUM
gR23tF8V9Ij8KpX3blzXFju84LjT3F6ad938dHFjeeJVKfRzejhDqbaniRBUqzO9
CcOMA1GdEIFiW5tB7b2jV8OQmF+zibPQxeC9uRCf/xxFBTvtSWgZfyzHSvhDJusI
dKu6RBTXXhKgQoZZcI3hA6gMq0LHPqQwESN4X5CEO+Fr6+HJKSINtdjNoBLXINZe
6Esn9BMlf/Nk+dBiVKd/AKlZD8n12vTx9G4a09HfMVX5jY3t7QPk/GquzTPaGiMV
eLFVVJT7E+19bCSWddxxw529xdpUsIK6LblDrdJQUUkiPq8zrkAjpJjs1MH4H8ru
y9yqpQZH3wtH/iVH1I4r4iHV2B+Q6PCbM7Y4edMNHcMw/kXfCeJbxsg8olm1IP8T
4W8+h5wPHavGWyY89Ty8EA1mQl2YA4ryj9EUPC0J00DWrAPGo5qUdGJcnEUEgpG6
18HIRcUmZh0IFm5QsHFTeTGbonHQ04KVezlsSRIDgwy6zUg/ApUvuQuG4xjyzO1R
0TJl+pAca342XZ/hqxg73Py1MSWlY1DFzOCFVUqOTSL4bq44YLg6lPpDhoIeOZY+
IZh9b057FNEukR0BVwoxal/jywQystA3yD3ndY4zDbLgTVG46md6ZU7dGUGUaxuC
Gx7y+9ptiOaov43z7M+GfCIw5+vwYApizQH7lBrSZ/p3pdUsQflZbY5/MW2cr+iK
NCMjDhegny6zdBlw+/FusA7dN5fIGMykrtnyKBbX2sGlw+URFUAomnUZD6mZ6CLG
qKQDb5yfadUO+Ssd7amrhgBntmm8HWvWWL5ndijFwOuItnihWyvohdOdoCDN9NcK
vE4CvTCCeQho/nT9FXF2Tw1YgpL3TLXRBlsEz2BToGsFxdnwm0KNpdwKnqx20lS/
pqsHPD//eBGeMN/62H7dhVRwIgwNTkdtbF7sYpYlbPPdztd4r2m5YoCtnEQnSgaF
yboTNzBByJ3vIWm3HaoDCyljVsx0ajBltWx6rQC828IWNcQ9N5QNTvwTdVIG1HNv
OTK41UawhtwvZ8g2Jd8KQKqZtpYbSwqMWXtUqGWqeo+/pcjszknL1LmkJDWZ3wIG
kDzUWg3E49ymMgCs+HgQo6gHALsPyqHoLRNka8hss5ik4drg16dEq0BXbiClQoVy
4ckFZ5T1Estz1IuDON02LVAdEybEFb3LaxxRmSkBSaH7w7ZUodzd4PkijTivRaPk
16nWnz4AofhcxHQiVlKQg7igkH8Ly8YQx8gNUIhPfm5vS0lVJCszm/036+BwhMQQ
gAE0tVBsEVRwdvWp5IhZGdcMhGxP9nfJJEF/Qt5MILrfgMPU3WLodCTGPVJxoa1E
FDlXQYruwzukPNRyTLQli8B9NSKG7KqsVf8LquhHXJASxz4vlgabd3vbMimI/zRW
PrTtoCuNJcr0LUAV+YG9lLABENj2clrYYx2KAkFkrlEVT/pDvwvcxt8cMPQn1mYk
F/oMbaE725x9xdDJCEO6MW0TC1HIdKseTjfjRjJzIWAklORqJYiHx6eCmcuaolrk
1NtxRrxMWqxn/WpxCprZh4JweXcL3uLW8oJIvSnSWLiy91k+Y5fYK4NeuaTTWow6
rIE+E+NXlBh9mDrHejK+OaXHuRGJ/ocvklg4Q7uM3sEOEO2O/uPi6jGOLvg249x2
k+B1mZhplkZXPGxt5Plx5qX3vBCYBUqDwI0uzpbB+AMZK4437TS2WU6aKPhOkNVp
hyL8AQs4YKwPrvPYOeDAqpXGBAN2+HuZKyXEOe7qFK6Uw4H4JEhoIUUqVAfRlOaA
tfSD0WhXWicr/Nw4H3Hxv3U5/0JQufr1UnmdAVFMQtxcNgPYGy11O3TOz3bSJTm7
GRD2ThOr8tTXe9oBVrg81JRJvbX25CIBVfDvxcbmuocqNqWXZCmecLpvGCt5GmSs
R1CB/4t2YeQDCeiGfyrHMwJu1AP61Jzk0X/atOcyw0x5i0WFkBXMxXfaluLjnWQw
RenGRnlgau+X6Ps46KRWsT2Jf8S//Tu1cKd4xMF8kaYgGNk/skZprE8/r0UcO3Qa
Z1sy5ssZb3dy6f8ByuCofqJNHMhibqBF4Afg+7sq3l+U2qlxkTu3R8Gtg+bo8GSj
WusI43EvXm3Lt+bpT0GUxso6VcwovbqxDFy5j1JivdxWNfbvuX+2YP2hYPcRafmK
9u9MBGPgu6uRAjdgzqI93RD93/bYKopXJH+w7fFHI2YMfjEZ0yIzdL1PlnNP/XGk
uMH9SWVO7kSho0YAj1AbxjTIKw2WedTKux/ibC8QB2VYEd9jbUASTBg2B8+swppJ
dbzopygJ4uN0CiTW9FqEYZo7rRRuv8GFhUzgLrT1kUNqf3fgOXTkVImXzUTqsYEk
c7NE6yGjTiNIX7l56x8MJIeK3d8Z7JgszM+D7PIl6dm76dG50VPU5uvncPE9gtPV
BffeBvjdCiIxBIXBdnzYFbVpRhLa199+6aRbu24Pts0TEjwJxV3NjIQs9e0elq2+
815PvAvdxbedsgtI9TXzrZvGMGSsHoipUF6wg/0c3FTQScVzgkubUaqXIAWyWlF4
q3HCZrbXdcqTeuleCOnSLnBd0GXkm2KKxGSdBXuLJgROVLqPGUlvfamef/H28Ol3
qxn4aO+B93kKnotbUqA6rRtDpoKzb+PinFE76oKoHsvZbLgdAg5mIwMbJeNr+0rK
OwXEVCr6Djgkh4tJqTjTLbhDFhV9fdvz7UYF8IqJxhFSqLG939eGt8M1j3LgOPxD
tKW3588KSYABz0vHpyWrbBOF09Mhox0FwwfUYrcrJpaLDBk6Nhoy7url99UEe24T
Dk/VmYdZUCqEgqk1P7Mk751UZ8eeVkmQUmU3kXjn6F553Yh99Ev9+nkQT/UyzOqd
C8WboWjMEqP00msuNYyHVXKlTd9yDlsUeuv4GVTZj41+LdqmS31xAoNuaZ9xqvJc
TgGCJl8m4sbI2BRcZtRRCmiPOe1QIIsHDe/My+d4Hd7oZR6TRvmrkB1zypB9AR5p
k7G0oPAVyVZMU35ojCULEBhHbv44kJHY34cGn1zodrRQylb7DLAxI00C5298fqfY
ZjJMA5HeqL7b7yzQGWd/yeJgpL2+mOWTtUzYXAAg9lMW4x5uygsK7G67fKB8Ag8u
LqlXY7KaoJ1vgZxd7jQbIbzUGFkwKD1iYfKyD8okfjNxxmewlAAnaFUWZHdRDD8b
GAUVNxHmSa8f/d5zt+EQiDmLxHwg/084nWX9Y2dVXyLJ31QdcHuN1i5RagdcGc/H
yruboqR6glSuLbHL+PcUytxpwA/256rQX0qsSG/LhL5A9Ee94N53Zv9Udv3Xrwm1
oAXn8b1SFUosNPBz9ZDvwzY7y0ZeYRXz74NUpXf/6ApF76XtuPcxATJlpwUSRz5k
z1FK4jcaz+t3swYpVa5xp7lWlAytzmXtKBCTj+JkVI53sMqAqyXAw0dCvqxs03Ox
lhMjTcECTrTG9mgLAtX9VbnfvG6mcaZhhSVNU8M1OfjHpde+yz0NXc6Vwc35Wstd
igy6+siBEgRgSYiY6/a2E/9kOLZ+r2QtCDd4ntZ+BCkXAWLHUXW6ogfs1tGPUBBr
bD90+bpj39M7SDxzECrysIz6TFIaZ7k1ZxqIIjs2Dd2JRCDc7xjwIUeSiAOG6mY2
7B/jLzZOTl6O9wmuFtcmEE610ksc/pKYNqwcoSaiK3QX1RhQI6cOIecJRo5hPV6P
BsR3HAjK4UtoLEFmdi66fQQ/WvDNG4DYHmyCJjouGxbLqvUdUcJRQdSC7c79fnCU
FheFboDrg+LyarywsA70dE9mTDZwKjX8oJbwCiR95gUMPjvWCD3u7LUiLQszsQwf
Sbnemirhr4YjplG0CYYo4b/nb5TiDqok/iduJi5ToGAQUVUKcwbRN6iJZm1l/Df7
bvaFn1+wSXA+OF31kuCAagZERt0c7KEeK9DY3ef/yTJBWh7aBKZ78nIqmCLL3mmx
yxzdUr9kMHzA9v/mPyLt2I0d0UiJyh2JXMkjMxB+dxmR+QrHTVbqZclWDMUapDCd
veG2q7dtSJyYFNVYLFmPw9GRXllY/ldjBa7B4cnItBRRb7WHYcAkisyQOO6AHWvQ
EQ3eDRDLPDx4Ew2gHtXyZaj4XVliFr8LwBVvlABiOVVQ7/vWi8LoSHjd9XJLRWM8
KHD57/hh9LhngwbWzk4ufrZapuTSG07xkdHM4+jCujcga9oPiXvKGkcRsoEdwOag
oobGyVQv0d471bL+eactTod+SIjSaF9n4zzm9/rsq9fK7J+2ix7veKA/7rxfhvqD
OpfBkKpaauKX9pnqrNzFzlaxoyH9Mw16xTyOdmg8evQbcSVLmqsXN8AHJBjp+Q0k
hiq2fho9VFtZteXBonRjzcYfFf8Wq0LXs9+G/Mn6wVL5SXd4/jStrlf6gwmrCbHY
cRieQvkhzfnq2ENf5n+Q6KM7fB1TgqL4w6jyAr+7x+Iw31d/IvTqsoct6AbJKqLq
TmEqBgRWknOoLVMn7RZQ1JsVs9gif2Pm0efA0ZAXOMcvRbm33DT7ovCIAGyyuFQX
ckFh+vbgg1HfhsyU49b8fToU5g1gakYAgp3PcQHLb+FCLeqYy3HmfG4U1QR+7BL9
5zniWmXBR5FnyMO0N3NdHa8Ynysd9a5MPyPWVzGWfiv9OwXuH3WSiNu+celTl7Mm
I7OEBhX7Cqi61cvmKmExvDmqnWMtM59dM34Loh2aRw5Mv5WqVrSfA5fGAnRSOURH
B2lYfa3o09EFXrBUyYXZh9mx1TRk6ZOhT8EZw0LEzRlqbV6m6tJuBKReZQNiBHyF
rGkqJf1WpCWOyLZMb/J/y/n4fRJoBTvoKnzMlOUSA2vvQjck+Tju/aCB7qHbmB65
UdiUAF6hxROeDYYSrSeZk8dfgk/h3z9fSG36f9CxQUgnq1dzHvTwnqZMfD+dWobO
HQmu6hjFLqYdg54w6DVVsfWlmQWxFJtO3UVpbzBhg65ggTn9ayFOVFlDEbYaFuVh
6WDIT1M/im3jzswvZSSHUtOi+/1kX4d9ZIS51kLb02qcZhIDiDtzFGiIY/Gh2FjP
11I8Jx4j9rhmPTi8vC1EidlqvXrIRIoJoKhkmKpHAkpnEPsX2xhszox4prR3uafF
307kDx0BtRzqOclT04MxYRRddug/jAcWZ6lfp/orbiQIpQzvmHB2Ox2Ttv8wvzo7
JdgpXmAylK7pcXEhxXaZUV2yBhB5Bx+dfkDpb1WUlEeIUMQ2SssAkdmw3A5h//mj
0gpfvkuODq/xBaNE2OqKONH58qnYe//BkZswdavEEUN2+joTwJWRgnSHLxJbiPPf
/SGfo97bSgW1j6R7mU/6d5l6cbt1tJ/qN3VFG9ZoPE8iLXSiqQu1w54WUIXK6EJ6
Hd5EWi33l6uaQ14MXN3JrbWmM2zljB0W3hj89lan3zO7dyRgpFek3xCkKPZhmss3
tBGScEwa6a8r2XQNauMt7/u5TBVYCwzcC3XuycMMf/xR2ncamz2AchX6XjUAMUAI
h3nifoOJdMcaMBSp0CaClfJ/k/yKDaJMH1vSOPrxP9WOxxww5vC/71YIR3N7TFnI
G7nrIEXZzJaQYDdZp0NIL0RchyUMQlp0woezUst80UGkAf5IcbJ9EAzUEIK2Y7/w
wDxpfPoOcTpVWYN9n+UU7ktEo03ygX4cDvge1ZAjAzo1els8XFOQ/3Es031H3RxN
VtX/ysEejkKzmDTqv71MxW2icFkvbKZfU1LQLjqXvBefPebITJwrTEpASXFitKe4
0MdocrWvtLhzp8gCVE+p4Y8x2Oni8kaOMTPFgkG1F6mq8Dw6vQJ+6dcnA1DFP2Xc
OhQRKUQX/sTYcwuC++nVBZz8GXHiArRkRXbNvefe1pbmdlLLLIRvkwcpspd2Qij6
K6aJ7gVycOHaYR2pYYaZVhxLTfhiHEUf3Gzn2C2VkBXc1DSvBI8UX31+s8CFNkoE
G8sF9haMYqvJX0Vzqgv8vhGI0E7tVtUOwSL4PjDug3y16UwrnOYy9ytDM5pKPj3X
VIvxm/O0t7M8zqJ4O5duVCmR2RyBPnRp6bMxp9ChNvleNtbl43l2u/TsIJm42RpI
D0u6ExG02TpqK73NHRv/i0Ox6+s6dbT6Ds9hNWLLHC8YLUg4lb+fNamH3rXu0SPB
g3qWMvlGFtsA0JiCLbPWQIxoegfYOixUCy3oKqTeC9folnRxxjYcAytVF7fpNYFq
lAkkMmlGjg+1bx8VpRVvVFgu53bsSe3cxEGixZyE+0VbCW1oZUM4V7j5dSkoAXoy
N/K/KjqVCITW8L5K13uZGyOo3+GtPET/j/UEdyHpNq9ovsr8Pnsi1Pt2+tAUh0qJ
Yy+ImbQRMc7CNd74GQCLHgGOHuq0usqROe+ego3siWcJ2QExZ1VHKv8HN/54aBlq
slW8UHn4Wt8HswUoum37Hyxi4hwReS5kXPDddkCiAafyqimkutjPeCE9nlmq/zq7
tkTUM1nzq0OlGJp2Ct4dCtKLbp702St0DtxwXWeQFDJh7H67OudUcKUE++z0Mr30
bRWUzWBthALzYPSI8QAloQb8cCO5RdY+qOYw1xjHsBeuMKKu9eXU/2xBql2/merf
zrEwOSvWTb5VqLbRNdcgeqenIS/aeDkKspcg442LPDC9n6B1Vcd/ht+Hy/ZAu3xg
Y7t3O+KQ8TFfjKJabVQhc1kZiNrFfj2tpZde+9Mm21y+Yv/3GctHqvuKMiVH45lb
QFPkKhIWrRHkG13Pq1iVGsYXbPqkHDTInZiiqrbAsRXCZiqmJXuXzacohQwINBAY
cOgAUv5I7Sa43qczzrP7Wsus1+CO+564fe7kxyibOKVSqMNXSMV0+jKaSzdPgN+g
mDY8+yQ5ae9ZujXYyrOPIaAnMtiRWzLx8u1mXkzvSsdzIfG9+MAJHhqRuzb+P4kU
PMNJ54dHjW+/yMTmWokZ0nN1fPWP3nuvZdJIMsvoYPjXLZYGariP0fbBCimgexdI
nOhGQSiPHk558t+evCDUdD9g/exkc60sWTGCbkN82K8PQdkulzW5EL3BfwfiSQDx
VTTcENTaPt0futAUj97gq3zA6xaWTgjW6dugQ0wduklghI5yhzRC7+I2cZQvwqtG
9suAJ1IZs1zmmgHW/ZnPBuBZje96JDx5ebJSrWPryDa8V2RCZ75A/Ns5ON3JJuyU
McSjupWn0IeSIuLyl0TSA8Xd8k5btPiAEDCf/Ln2Bk9lXU3qtvzAA7xRUaEC8jYd
P8WdH1/h2qaXNECtpWzcBnMQmnG1Jtxy3g0Tga5j57xbf2A1Zy2zLpRIHKX5IdBi
qcQXdxo/pDgCVv5NVoFHuGuGDPaFhUF0ZHvfJNdxYeL3oVUdkR/yjQ1I5HXJk3Ho
F/yrs5IrH5c9f7xAc+h1L0UD5m89pTw08jtXoZGhnTLESd3crSrWhLRJE/SqqNtj
L/e+E1v3z2iXQTbG99W2dctArElzoudD8Zjcz6f23DXScxBaJp+B2kn8xUK3yCYr
hRzm7mkfnu5a/xYeRvM/bu4jBz9rkwMS4eSz0WFZfkKG7jX9rJt+AtL85ecqcYYf
s0/MHiFW+P6WfTyPjzj046sdvXL2SftJX9sXDtTWbwP9oPXWWoDSuhMhkLwVtSo/
zDy7r3/gGyQCchtFupO4yHuIc1RYh5s5djKCxPqqIGeWP8jHBj28Ti8i0ubPIIy6
P4haRu+kHjZ0C6LiyJuI2mAKBbJrIsPwKZCvZCpe24LsOkczhAEgf2Xzo+p69Rmo
cX2rozhbHFEwslbR1YzEIdEpo21yCSCaYBY2xpjb1ycCpI1InGne25JzBeCmf3RQ
brapXkVualEAU12SGWzGFprzLLUjInGT0L4s8knDz9ZM+r8LDi8FmNZV93uDWFgT
NsindImPTTK/+h1780b0SfxGCWowmiW0VshqQ4fTFvprNiSYy6Rt8UF6O6PTSurT
2IOUO/FoQw3RRL1as5MCoqyy385Ie2DydXYWVX2rkyKHD7VqDeY6/auiMnMaoLwR
w8MU30uRJR4mjIp0xZmqjotNtD1YN+qkDt/R/OiEAo2b/GkfLg2i3DWtAJfeCnHk
6eanDFYauDpdPzkipeF+6cLL0ZVZkkdw7WczKIztIlqNfRp/Sl4cGxlUjTqlbPhw
ivx2LGM7EfSqIvyOEU6YtWsAWltTT9GUaz4d9T7C+MPZQyr99cDP5CPqEU5WNBO5
g+seYg+OPlOETkPT7JEgR8M8U//O30n1Lncwm9OnWgS85SFKoiJj/iXYZ8oTcd0z
s/aFRIGneJmlBEqIcI+o9w29W3EvqUKfJZUPQ6hSIzwzaR5bRp+etLS5CYlsEgGi
e7JkXs6DRvAVoCkfKcYwCZOEsBG8zR4fKsI30PRMFB09Fu9Veh/h2sdtutSBAZAt
+6+RNzdHGjhHqzFHL0dks8d4mkBJQaWHmVE7g4a5dHMbOBlk/7yo9NbivvKrx9Zx
rFCsMfIxW01TE6LxL6PJgeePXxBjZJAEZBskp6JOJautMfid2SlaXM9/4xKg8OM4
ajnwOy0ZeSsrTch/svrVb/BYseCKRN14wBlw3Yl0nE3yhZic+P37WgBPUqr1PKCG
Hvqus57u6QcuR7BKPem8wyg4/eOo1eEEu+BhSVA99/WyJHPUSmNVW82vOjm5ORkh
+h/MXI00N/D9ZILj2M0ziel7a8GnQPFGTTbU7RD2GZ/AHcCe50nwKK9TielBtpiY
25p/lFogRvG6lNIVJ5M9gTjhBi0YclMwPgtCFS4GD6Z27BcEg1oSC8xiaFhNpUHy
PFFmzYk8RiA3BKWY/XdQVZIdmyzPZAvpxbf0ToED6bkPAB7Xc4Ola1oJ1CUmpmAa
V7gFxEp/3tLw1s8mA2FGlEubx41LmIdz14zj2JwX0UEZEQUEkJCjfRKNeFrXgmr8
P4Z+32KOUkFaO0HdHoWM+SUleHFe2C9CT/FboVttga0WFLiuPVFH5QM1zxcgD24x
qXdE4e74GZoweJnaqaeZh6FYKggUA9zW9CiLDul32AlaQZPHOREumapBEZIYEFmk
IgXffE7GcaH4rgRan5k4KvlvZS0BqgiS7WzF2MtkLXcW5iPAWKX5KwhSSLwR2b6L
mQySrqcQkJccnG0MW/eqQ3eJyr0DZe0tlXFv9VmfcOVf9zFhNvzsmamCIY/BM5sY
2+haYx36e2cYi0+C9SLn1dZev2VUx3C0ZcP40/5tkwfodovj5KBk8u5/a+l8gE1Q
2hnqsP1njayaCe7qJquIZSC5LoZIykUJjorsey3R3xPodzF9d/e5L8RfXW/KbXTm
uR4/J8rjwZ5uUsbUPrSTsiLfrqe5NOvGXAerK7mw8UjiswLbbLj/bGbx1OZ1t7Vk
EOYN5c74sPcljcRuR19eDGg4apzJK1pzMUrYRrazIqFgfwdgYyF9TgX+W78StLPs
DI76VaRHU8VD2EkIfuVAVzYzmfXmQbzSU1x4cCGHWD+NgHMKUm6edXBjrIdpjKCQ
Y/elNZYHFbO0prYw3o+2z5DZ89xaaXy9/VZJfk8VFEeJakRvWyFu7VI+/8vJTqgn
V/8KwKvwHRfaASMc5wV6GLXWVQ5yendFdVLCHI1WXs4br0aZSU+xyMITL/UM8tc/
kiV+1RtIZrp32L062LcLTNFA7QvPifvrvY+8GewlhV7KfYu9cmT0lRLB7hLSyAFH
h25PreabqzxzMq6UNkO/s2WPMXVnyrQn5VhdM4Gce7MJbxtl5ulvAhUhvkUsm9GU
vnUtxbXGF9ReqEin6uZ2Kern1Ts4BOlez8bLhpynYeuwIIAr3LQiHRWqWcnnI3r/
gZnd26znU86jMcN62KyGrMHi8eYrU6CHTXmThS/eyuXnuK0Lp+jTVgdsqr5quhZy
/Gyh0BsiyMpUm0MIC/ZfkjdsgLS/2WCcA1mExafr4jzk/xZrMv7/E9ODBpn7TXOr
OpUmp1cbAjyC9eLHHgh8NVbmHTgy2NIkRA/LgrhDLBO/2uPqJ5YKNhUqjoaE+wCw
OjEIc7hcOYIlXIhoeRR/cdPyo+46cOEkQ4GD9wuGUShfTwdKcTkPM7+4Dc9u9+Oo
pYJtpj4Gjfuok9S/YafQMRm2QV6re9f1GjqoBfdQuQ0MU8lkYEdYF0dlkP5OQ1TP
uWnmsVqwK5h7ZgEtFGsy+ntDPQpLAzOPBTXinfynxERobY3eyaXgGIEzBEj+iUFu
u4nMRf9uyTvAZIqO8fU5cynhmOsvU3U2LKZl7Z/xb6DU7WmIRahgpGGFGVoBxs8T
FOEmusPT09YqSyxH+Q5/jzhb0GxE3UgGGpqFpAcQvPFdRilqc6bULKqAyu0wGF/a
POHu/yEPGirr3lQLvYflk3kvvrY/ciWJHOprTZUwl1ibMxwHMADIaMbZtZeG5DZo
zuIN2cvbwCNLgUYstxzLkBs+gMC50m41jwgUhfBOneypXpHF4J9jZeC3LEcWmdqY
CwNbp67MQcbqvE3wQX5/l49QrlsLPIj4cuV41JCRecQ+pnFvObhW+9CSyvhJN2UU
qR2XJheBi3yebPDDvJesKFYh+Rvs/KC7NYXXj47r/05iscJMrAp3z1pF7MhrijNh
KIy6RSoVm0Z1+huUkNfsxRb/xsGIa9hC4dBkrmgWY0fEE+w6EFrPa+3sklPlrGmt
Ld+LbUAHIdQeqaOdSIoEyHorXPoB/3nU8Mfb3CJgw/MTpNpYb2E7trGgKbtWdK3w
wMSabIKOx8FLboYVks4i1DmTfsmgeVdtFQsw0+tL9yi+J4o+nIqef4zVWb2Gw0hr
NyP/Zaf4zlGhu+y+ZAEh/30NTg6oxR7Z3OOMoOQb2x833DCC1F+Ws0w0OpmBb5Cs
9Vyzjneyf+gvi6PaZj5AGwrZ2tFaqDwh36ZCS7pzzYSCDYIh9S09k7DP9Zj2T6i+
B7m4Q+Xe3CjZVm1kW1qQ8o4kTok2ni8zE4edujBetQkNcYOmBFqhKoqrVZQUGD15
bOzX8Vl3n1vanoc5OQZ48HlV6PYMItRj6jOnpez9gD5ZFXPUJZCTo61Iyf2LsQUh
ut77th6gChLB6nw+XONz72Q2Pze3XluYFr2Hoel1IpwijqyEXOgsQgy7rMHC+WN/
ypZ6/QWZskZ6XT1vzAu/eLYiwoRhP6X/YAtFPSESHDo5/wygQy84fQzOZxMAwjoF
60CxcD7QDNK+fVCV6968uuczC76lw8T+4PL4oLJFcbEHkkQUoPW2UIIiw9VpKju8
RGYI2biAS2b6ZStiMK873XipVwtXzKA+uQXp2/c1wdw6UJg4GsvjM8WqF8zLawL6
ilzy+kApVrYnfybRESJKXSKCVCbDKoCiFnY6N1GX+KpQGA9hZpz7uAvkA7IG3L1Q
m6e1EolJ/xnBAwwLqLuno7r2jwgLpfhivrhXcGak6LirtVZB0yx9PIu4YDS9OZAY
9W80A1Pmr6B7QIjlM24PlGzqrd24W12Y7lMB2+8kTuisdFJ1s2QVru04MsBhpfay
IoT2BUpNzA0ow373hCFMOrDLZ8cunHv2l7ANzgl0Nwp3iYaWJuoc3y+z/+YVcBSQ
oC+IF8fdZ1ZscGqLnrR9+9CTR8axxoUGYkDkuGPAkoI9HloeVx866j1ZOVVAk8fR
5Z8CNlMDKDZhuH9k2mATMlklwhDWiOJLzSeoklAeL7ebR2ts/13vcEl9oOpENijO
Prb13/F+MMY0Rxck2xd1ipMfG4eRmvJK+d1ZaTmpKJJWRIoJ3pvazBRN6AG4QmkS
bxZvijUAvHzQYTs2aFSamn+ScANWyzdWyIpx1revqk3RbHg1Xm96TecqKyXx3vDp
MT/er7PGMT+fIuD3BjZ3PMeKTSoj4Vwid+AV+7dS6fd7moo8Ua7zmd9cCh/pHPNZ
CHNzt5s2i3ljnNdLqv2JnRDC791R74IUOF7PAa7XleoV1h3euJawI1BlEIaCgT/A
MnJZY0a/dB0vKjgT1pq0XvNDdlDEJpQj0VX/8SVy6BC1b3uJWTlDvJ5SZc62f/Oi
u6+lg03AYxSRuElWY42LcV/XbvpXtcDuPpfEhpMcNbpYEYraLxJ9JfAnE8MvCSUX
uxpXEJSogn2PRkkq3AbmKZiwD9VbJeVOUmTJQPJ35ceKGL9MoKmEBaTewu4zTi8X
65AC4WeM7Qpl34LujdM9jWbm5POAgUstLxxSW02ahijTrmlN7ZIdsq/rLXtghxf3
zDIQdCwIY4ghAR1WEnHoNhJvZq3WXTimhbgIJC+ViJNc4NXVhcKYpgwaZaAvY1SW
NUjx9gmrmP8H6WdOHPWX/OfY9+DzO6rBaNRkVk2eaPua5MNBZwrKeNDxOvXBGfQ+
V2JEKhCQKi20Fi84A9jAuZAks+EWz8HlvbrHkAM9vHRVloWltBocS/YHeB5K9X/x
2zLYcpe18wPT0dhAhYkbi5U3IqeKULrh42YlFZDwXfhXlBDeyUcdjTbnxIiUc/sr
gsWFccJqFDzwAPYzHmDjOpKw4tLsHoYxEFdeD22pkJ1zbXoGReXrzXznrAayAtmw
Oc9cbZwsQcPS0iNK+ES72Ki11sfYFGR9YbDRu2b0biokU21nEXyd7E0fTXSULQJn
mOD3jl9Nl7AsuOiO0dVaiTnzJ1FbCU19634pLztcPuJWnewYBirz5JLRmI0waEkg
1yCIM25VgSftAgjTsWFfohXOxLNH8pkyBgxAQvkbb80UNDVWN716UdJ+0YSMgPxU
+bCIY+iZ8ydrOPBRTOQS1kCunjQgS4cZPqLKg6djVdfS22xSj9igpgCN3ukG9jfk
biQZYnAnGofiriXn/MgNSSdTvngOI/iI4DCiEvAGX2GPQ9L/h0eJBGmWaccLHNMm
nw+kj9ColYsYayzwpjECgiApsrPZnQpF2gWwljlbTkrefb7v1XskdpNjamFGET5s
hPQqX9n+CE7mf8eRQcgKjhKsxjLLMhH0XfCgFxO8RvsQsNrl3jZwVfPZWMxsRBCL
2NVm+UBgQjGei//6EaruPJFlTT1CPThELsygMRYf+MuyCwvjwSrfm7HgOtyLqKf8
oWwuLXm0rGIR7MEivKUI0JqaWS3qVsV2gxWZElykACwDGVGxK4KqrxCW9n2A7y+t
KmtY62eqxD9X46poQRfKOGfdJs7Q6CfAulXu7P/+xWHhLSE12YSk7dmYfzHKyoAA
OBb01/MSY+nrPvvbt8bPmKlkD/nkeNqi+sKrvVQkzYDp3eE8O6iDlZBAxPMNJp3c
Mu0bCOycoQsZenkxtkcO1v6SkpFRyZaKMTyYmULhpLsFVrBYsrf1BFFcW7/36fEz
y/xkbw9Lu4Rb5eV36o0LrHRdZbcspykaIw45BbQ8cN7/GxL0kE2e03O296DXi+h2
SGx0zkeVWSFA8/wpc1HcDkCgJLdcfHO3ItBgv4ygH3UxSZiEv3J/TfuoJE1y7yAR
i0VI3lxb0Wo0Pme9uwgPBjLkiGAm5QG78B4uhRzHOpiTEPYxy+iFicRSA69UGT2G
+QGaZa1owjlZ7mwsqNebKux9sEqcljVwXrDnZFwCOShnVYd1IU77fue+QAcKC5RI
mdt0HSzhZ63CPf3XJ00MX4/6mWYxmxrLDvk+H03Q61CoFkuQJK+RwrTZSCUA6wmT
wq3Gm6XlCgraqtivgqKVDDmypzl+Z9tYjgo7pCi3Qbs/2yvqAaSZ8QZrSWK/HmrA
NvFuQne/tIQghcw5U2ckxAXAR5GBovH5e4YYvvuONg08oFhwyIryKqdMWVhJbj11
ThTGVjGEj7Lptzw/wD99vaOHAM0h0WQ9/Tq4oNLS578C94Ddy+C/+RmLbNPRNXyD
3r2pzXtE0DI/MSEazM9WH77Fq4DzArsfEOPFTgcR5Wl1C6zI10Iz6ryV8LlJv8VY
GG1QMAoAP/fa9SJVGB4IAd4Rf1x9jUDf8hQc5ad6rzxKo3wPIGFMWCme9/3QIBUM
D8c6WXcydIzUT6Sxyy4yLfDOK4KzLMvfZwjaO8+OZzR4Do2QvxvWrTBoMgzULIoP
WGGEREn+U+Dt2/VB1fYGVA+RUN2xJEhHgLb5YeuzmQ8tetjIsmSDdbpk99V6CZgi
cRV0TOJH9B8vgNTe4LAsColIIOd88AdpLISi8T0nWSKsdSKyVQGIqbZ/1MIAetWO
m3SidjweGZbQLeR4u6kUy4vkcACXm+SW0qu3yrZEK+8kx9KgDOUi5URbrSBA2yK4
KZTgDLzWGgt4rM5UpXlS6Tzs6elA+sxs88hD05ojMEFTARbXnd7TbC3zEa0RFwjU
1em4TpJ21qFLWDNh3um6/fVEjX+3byBmOsoF8OGu/11lk7OMa8mCl/SPHV07zaNa
Kk+cO9IlcUWuu4U+XZr2K+ZVMUuqlBVEKQICJTOZMoREQGTdgw96Hqqqjv+O4up2
3EvzxW7i7oGs8gSGwi03XcjxfGEIWlVBc2cGdrjmsdrG/K4aj1GZekvG6IctTcw2
UFuH9RpNtfWoc4HxZDnwQSAgjKkuzY6I3S3XqruO3PYYMOLC6v3NfZLfX3eCZBSJ
hFc2ws0LSTPmTawY0HFbR5NTLs5ZZ2kLKvEvPojpWG3QGDLhsDSzSIwbFjLbKTil
pW670xaZrlSE7ReQPlFMi3vc7moI5FsCtlZEPY1NXDMhdXaFZSdfaTP6K80E7Mm8
th4rVY7DotiyaYVCNWFFKlNxIRBK6PPOiL41YwRt56FPsTC35XNWtYOu66Pxh9l+
Y4cRXmyEJwLCKPxgdXYOPdAxVAFs2LpYnfrYaTmVH9DAF33ABnBytwAzVMjqjLpb
70hoSKgmpvT41gOeYsDmPX5dfBJFVUnTlWE4jlqm82x+Gb5IRIVwTWu3WEA1l2Pq
om4KVw3T7XNMtmrGh7X60/TW+2oshudYU5C1JsIes8kth3/3cX/nxGYFV3kldYml
pZBNJRfmk9CfwvngrFDnX6EnrqGIXlqsg/YCHgcpQ7e67wJ360zNbgUBWd7gyQiq
+gRdo92/DxSjMtbEkq6XSvnR7umZ1S0qz3WmzgqGVWJB+CwVph9ZSwxB2/7AHRZ8
YV/UmPnim7pXBdG4AG60BCmSNJDL29t4wtx1hiHQKFCLsoqanHCNHJnVqnZ5SaO2
KdmCbwnfeZOc+JjAhtwnU1fCfXMpftpG0ZKtYTy+ZrpEqXcWkLaSVU5omKowolre
1QboxfL+RJmR4cOsLIudRkMvxPSMwGYRv3xvpcMFvbNlwaDE/E9SXmQmytQLvT4k
lJhpSSXc60qXVe/Oj8TQm2vtoq2vOX+EfW2yAhjB5qeenPUzT17dfB2MuQkidf3a
7rPZRIabgECehcvvDjPXPaPHpj3XMRJXVfkIshW+5X44KSF9DbUm611dNtNiJLLq
tvyoAgTGzThdiOdwd+Dj4i2X9OLOlatWd+iUedCFq1U13+63Pl37mFgbknaPGkxx
fjIN94e30i1AqTzCXBvqJ3E1YbPjpWZO2E6BrVp/pvymUMdLKkh5cotxiNGgAeTS
4u5zUh15XzCHhUFsfDOQY+SXVpT+dKwxPum+xqyZUed8AOjd+3kRFDTnwv6j8m1+
KafLH4rGa03oJal9I8va04MdVM2ET0TG6kAALFh9LdHAffWVTIkz7m7rXb180xTd
MqOoPEE9omAFsrg+ORsasbbI5Njk5sDIDjBdf7DkPhgtfR7i8vZnmiOJZC85mZrP
zfqgwEzI0JdN6Qk9VvuLSYM0k9kY33SIDhgtZeIj510ROjday+k0w5pr95+pM1VB
nWcGKAKpxhVK98wuhADIiUC4670TD8KAw+h0T7wHuZQlYRhH8P4GKHyn/oBJ4GVY
zfcxZpnKE0mnnFELq+XJUeHChr3VIp5s9lmkKXEIY4JC2i//oiIKS/RY8GEaBE7g
QiFzCCtrG2LEn63Hf7eEqXh3O7owF5ohlvS7769K3Sd0Es7FcVOVUeLFKHLvodlS
MApW3R+T/DdxCFHgwKx0DOS92buo1lHuYCZCXq1aqjQI/lL3rZqZddShgXGBHJTz
iqCZmlhDo6nRTMzIVajHhmEtoti5RrS9CElpasgnTRvYyjue+mQSrS/Od0XJbx+3
xmTt5HGJLERBjIsmHjXAUnLbWk7h0GOaQSD7zQrdWlqAQe8Sc8iszsi+e93L8x4F
+5POmrTJSS5/qo9GHnaimiH7UU2ogLdT+NCQifhPYHyAAY0rIsCQnqFlz1UCDNUf
nbdKlTaMRW38Dh6UCw0BpDoPCQlC0NwfMUWQ/O1cFbXacwDfhynYFB3KblssUJW5
gI2wPLr2jZwiQ1rjisPbYPgIAkB4HSNZzPWttmKPx1iubRQ5nqcnwsCOIUtQ6UB6
Rp/8gqNqr0WnoZZ8NIn0E9fCalvkkzeH7pwyHZf5ev1Qsuqy/uVifF7yraVN0TfX
ulFNtjA0L0za4ULQVGY2MAvVxGl/L+YpO3wgp9o6/JkInlUp1sNAPZLu9Nx9CmXT
4SpPrMmKPMmbFy3JNGJEl3OMrMJ9mKifAG+/kR30YJLQVcv9bcFA16a9U1qs+ujU
uFyLwwh0P/1FMROMdr9us3XBE1kvjo95VIPtQ+f619T61Ds0t4UASLmjQWIadXIQ
exgSE6VMgQ+ZpHaKgBwiqlfhulP41P9zvyaK+veH+U6NK2+irdk16oP1AHLkcF/g
ik5915C4pyaK7MV3HxHqlu2dkuuSGS4KPj7RD1CtVG4t4/HGK4U1nHb06ZVNgjk0
bz3EPP0EoYmVvZWiiY5Zlu8Jl0YYYN+LMtbBSTdyXTVRuxCS5PK7I0fbeAK2o4Do
ukDgUZlcfzcpQOHm8JaLWqFPsegoGarjyRAdKeP+tniL8P3WBZ7TgvsQX8J/ktH2
plS55hH23Bfjh2D90xurRE8OCyujOVsT9iH1/x0GWLIHCGydyyJw5OA4+Ho84Z9L
x36Ma6cX6WFrkFIVtIf9mI2EMuxy7LE0yzj7RUwrYThr0ho9Pw7j7TYXYq9ZoDhu
zrHUn7Oma82N0mkPpD7WR/nnlm6CzyCmPHN0IUrBrMlcqkYUgwRB8WHJT/qFmi/G
SuwX8Riqwu/KXfZ0Ymta87wOaMkOaOaoNTnU/UI8Qbs/hWEWi6JFaq1+8bftody5
s8JFDeh03zwLev7gzPYgvfaFxSI9mpNjWbmbQra8dXKCBL+UAczV6pj9uCHSp9Ii
L23H6irm5MoU8/EoRhGQGIz2GIihtlifuunKgdCzZTl0tGnIg0iXJxWJXeCy15dE
lwfmlNeQDven/yo+9egtIwBJp001DQe5Vnb2dkp8T2um4XdS+auydNnIZ/ICtQiI
UmpEfAUe/YT5NSfKgIdOpKWfjFOLyYc/1JI94c0v8+dkoigrS02mpuZ2H33DKL62
bCZhcIA5N/4y017jisxCwpe0Xhk/b3VAnPRnx9DtLN8EK73i0jODqiUqinTPngEN
RaNYwQ/3axmfZ0CCB2YoIL3vHfjwBerMsQ8IHl3jVDhkdTd5SyXjS4kZJDJxaJIf
P3pfypn5xexPOImiIjb41AxNXRH5tl4pmLkImu6KJc4mHCCzLQSrd1WxyfQbSWOS
leRgotxELekpfgfCVSKU3NF+QSF5vD+qxPjhAcRdPr8EF/p+3DXJTOwPsNiqJ7fz
Q6Op2NnnhSdg67qqT899a/bnCUorkNw4g1qRXQh+FMVgQTuktnQljKniw5FbylPu
vvfTpC8EXhRwhd4fSMbRH8HOO/MBHFupOfT/O8gF9nJLMy97qsyc1BvW4VENkKjq
AQ5+44lRnoUf1Z1s3PfOxVP2Eurs1XtUXROCNY9kl8XMr3N9tLY4LOAsgg8wzsDO
s6k6Gstw3oieRZn0XN4dRzrnolLtDeoVgn6zewI2sroE2uxI19mzMPG93129ahsB
018nhfqWOzaQSSNQnG3cGK0Bvy9or6hMLF5nqo977tIntU3DewWcTR8vxbECgwT3
5jkqI648l34tYvLRVvi5j5eKuHaPy5+vPwO0vOu8V52fR51d1WCID8vgWGiaUsJp
2UtFdFz6k9Tt/eiOz15HgeQJHxEBZaVjZi6VofOAULuZ3iaRORgOqRuAJX0xKcpO
DcBbbknZIorwHs5ZuVXo1OXcfpot+ts4l2sj6oKDfAmjmH/tywkFW18XrOKQK/9Y
/TCc3q28UNBcV1BjGHtf2IqITLjnXGv1E2DRjnvZXGgWCzkb3EQXeyels4dz4H0M
owILq0XKS2ci7fU/6F/EDsLXlV+9/j9Uh5yVHV4YeyJmYn9iIJXy9ExmtRMsiwm2
FRqd8TASNBWFwxcVhj4ALJEBZpf/61qS2F4UkbpvrsKcieWvLWb7ysyvDd4uUBRt
+ccYLsWCecLChy+7b2Bdqo4cTjCie4RAqlMBma91fZCpWmmCwuGgDMmGDot1rLvq
qPC2dNJJCku7pgh8JG58PMFKH1dD524102E7p49GpmCV2PIzpKhlP/b5lBr+8kO5
emhaKI0jRdSfW1O8KLiUGCPyQngoLAgIWVn3g6wZT+RBvs7yrWY88zbAR8GbR7iY
c1bdTe3XhAYnomWjIp0PdpR4woVWyvHwvfREh4m1JQ+m9t5Pzop05AzQNrv71xPX
8zmXMRz5/BvYV0d7wyc56Xn3kNdrI3AlfAGK08dOpsm+2hC1LfmdqkuZq2BVqVdD
DmoBa97FLA0avpyLbcPeAy6Ck8uefDXjCyqJDSVw8tPIl/XoYriPMBj3LqE67srv
dqKQefr17ELYj84PPiLG5t2NjSk1RgHmn3mKCk5CFtgYp23Die0DvHxu9la1ZB6B
hCJC46BVRtIxmtSG9v1S2KR0TG88LY425bj/1+r3Or58yDYhwc771f8D963ar5N2
Zo8PpKIvShU70HJ2yErukBc3BxUkV42B4qaiy3pJIM4Mg+TyPlLGeLFxAkVPRFGz
wjn06OHN64k2RMzZlEi1Gy0W/0jhbylFBxzCRas6+Enbu3FDWaOTOKPn4QTpLkJ9
zsRaV0FXSb0yqM1MfvTWj1IDllc5WzIntnH+aBRBUnSPGnOcbEnKYbHxztkMeb/S
HGtiy1aoiJCTTrFUk1yWRuX2aX3eQ/CNSQJlsF+1jCETMmisB9/qXxEe8bQyhqlH
F3+oJS8qob7/hCxmTB8GBJ0DghkNa7sHA13FtyEn+RpQHHk0NoDUes6IDPFFXAcW
voFQjn/cq1rgC13UKGjRaWWFFloXsS+9BMXS4q8BhS9qzEKxqdzVbTUE9R/p2wL6
FboZvr6HTU+RswRNyHvq8g9UvzKTtuCHwczB/tG76ZFpbEcGgbauLBwf0Pz8TsSf
Rd8nMavL9jbrPe5s+vQmG5XEZ6xcTForeFrsD6ynU4sc9RWDbcvoAB2KS+edWLnW
ccJWFBH/v+JhnGFZxCfQ2vUZ3Nm7fFQ+SzwsG0YsatJbhyLNfcaZYuZdH6owx7QF
GSsjxAcqCllA5PoQKrCKVAAey89n2wXGIwpXWBQ7vgykGO/3Z6t+UHl6zJhCNfmi
xX4QTDEzE9QAcEC6+66Kg3Zy11olBFSAHTXokPJ4G7sDIB5dIACDBcAeGfCNJyhA
SesQJTajSG/DKOP5pY9NaioHze4RwoI/NhLyFTMINS/pUHhB8dDdoKl2ppigp1/P
mv2Z0f54ou3KRlVxw61OOHyJa4jeX/HAku5fR9KFkt1MGRp2Kpxu1Zb8n1CP9i+u
L//T2F8vLJv1CH1WZ/FX79KOHSl2RFlvXY/Q0/Y321V3ndK3VLpRe4bqNZhloY2k
oMPVfTlWmjVlKSE8r6AHeax1YE7dcJyg8fvU5RGIrd4aVlNzpWWUw/cWTNSYsgOm
21H8yxVMG/2TcdqWQOA5XeJ3elxLDO/gyEdh6n5gSLX8jxLVI4+ja7pAoN/lrsSj
LYZykQDXZOZih9SCh0Fqe2ZW8apN4KSXOcP/1BtocXZDUaFESfzAGJfOzj3iNgOl
aVG4M/Cci/Ykoa5iL6g//BP898jqHeN8zD24mlWdfPAecSxKfMaMRrlgucdlZTb3
dMvpmiK68/PWi486KmtGzXERPTh59e14Pcvk0kEvKM8CFrp8RIGV4J0Zq3ELI8HA
I0u5OaLnIH6odd/h01fGpVBHeVU4o+amNIHpvtxOVHACnFDx2UKrIXQEkM/ZPvIH
uHQvwLvQimbZM7lAEWqNsB5venEVsAvIpBcVcRxkQ2PWOuzopaBvYxNgS5SN7LII
lQ68bISk2Y/a9Hn94fvcYR5Satffq8nDnfFX+b3Jn9Ze1MIii66uARQIMbTf6pN0
LKwy2n9LOWlf00D1R4WgGPnVasBs60goemXg9mDam7BWaeAnmFIzTGOR/lRIU42a
I/k8pK5YB3Rbk2F0ZJn/ZR9Oa0ap2AtF1lUScJ10AsB+UOOvD5KlUnrHhTYWYYAO
9YE98vzg9AQkckGqrcc81wTMxNjfNtT/xmNMLPmGtKCwBIb9h4rezeQPgQVrugqF
GvN9NSaYmagOPHibB1tboNjpz5jIL/KqWxMikQXXaqYm0INkUHTHIRwN7zKguTwZ
cCCPGsqAA72/H8tvz9bqVv5kebWAVzPAwCkHphwcJS/mEdZcg57aLKWH79a2CCq4
1Vg+BwKYv5Q3QcFl32dJEjGK4XS1ZFGb0m80+T4nnlrGX8qRY6ne8Dk2/FV3XDdp
JAwFQJA3c8Ite9BpwH0iG+WkMY5rniSI49KvndF8/shUNbOrD9jgcOEHqPWBK7qb
BopmHSHvpVEVfit24sRuafpl0lg2+kAF3DTdVaFfpmcr1/61dZ7pKWZryhkW5jRD
YH4ZOxVNDWmBnjflBmFM/yfUeKMismF22KQ4O69oBrelNJbZulsPMEh6nu4tSTFr
4bChJVaX7etVBTpKGIUdvFKuUNa/LosCOlmP+UCVr9BVXql7ljP33vnVLbm3+R7k
gCiXMyfJA9WYjKc+Hk7xj60u8GEy5+Br6fKMj/c/OzBeJOr6zGx3ktX3LZWc63qB
Ox6dNFW8+wbsZCsii6BWtUNZMHMk6OGfnI8MMB7W8vzWHqbiLTXyc9tKFrQUt7ZE
cqy/XSYzrjhhW55sYfQb9ZetCFG6rDr+H6jd9msgPVJJW3m/TgXbroIE1ZPdniaN
VuGDas25pUYUZHaYlVMMUSAKPTTba+DaHarDmLGp3rM4y6WyqnXD32gAYFZhN3uN
h/GXD8/GL0iEx40RH8c5DjGxJpAVIPu/ym4CbqdBCUCpsMQPXVmZnyxsY3nCM2UF
CwynFGcqzzal21mjWucXDcJl5OlCJzrMDyK/qfe/tMwVraCTtFP5ZgGBw0HeRMiD
d0AHI1ohSE+I4WNIYhIOpbs9RPAgX6zwF5IxtKxSl8FnkjAeqNRfOnIU7czm52Np
VhJQkD1hw9IbK+z7j5xEYy9+81VEeol1pNp65hUPxPfEOkrL4dD8DRBVgoVfaUC2
sG2+EVq8n6phVKBbnEmzuywI5+tXcKJnF/J5zMWaQf5T+A0An5ux25YYXFcm9O7v
a16m0LelXQSEoLnfL8Syc+FqOjxtdTpX7oQ86A2doc7Wp4I4nL1ToNJSZrEhutTd
mUO5JHv+RbRktWsA7LqVuDiVw1gFMQHOVPV00PlF5hyVFTOIAxD2hCCWZBNTn/5h
jbST34oZ+//xZ0gIgc3kX1jaRmyR+iVlr8Ys1PR2Umr2jlyBn1NlcpUQns0ry1h/
z55190NYVfoFdV5Awbz/a7+czFyX7HVcdcIB0mgdgLdezdLi8v6ag18b+vI8lj2R
O+Jjk+utK23YWYXvy4kTIKHbCCuvyZkuKjU+pmC57qwMoeTlvnL7AvYLTyEyzO71
nYHkGDEZE+UMRcFSAqZSxm+pHYm1axhqE53g0N2MKsdxkflPhIqbfYsirqby3kJM
38qSx4bisdKZyL325jv1hip38Z2lSDxJ/2T1XG2+JQn5pNNQ3YCtPo5S0ci//GZH
1mBelDT92X0lglHfmMqfkwTTMF/odpxYc5m3/fwVqgdtdV/e0OtjE7SnvG96ueCM
Fj1hIZx6nWrhQupehxQLO2Np4v4il3srmtKfG4P0oIPjCDA6Acq6Thl8lshpV6LL
5CNGQfcqFGR+XNvuXLuoCtIrusF3E/SwkZDHJN+JMxoppMoyGDk/5bSFXt4zJqK2
rLjDM+GqjU8J0a97EjBDZcFF6tvgHN7E5cm0UG/d1wCRFGXdOocrb4uQ23xnom4y
U/t7zinMtUsSQoj1WIjLSYwgJfg24N6/OH7baoxJpt3TfbeNmItDeiS9orZsRw3y
arfHWTtf95RbuZ/XNfdEBDf70YbpGnalHplnLhdUBsy9TJhC3YRtpOnDc3AdJn+m
ErdjFMN1j+6VTqkds9FIDJ6gZK3rEhazxLRwcPoI1E75Ff2RLvnwfmloArrA+pWG
zj684LWP184WDuKsaTML8LgOYI5iVj8RcDqXZK6XG/7yh4UrsjEATi5RtyeXWEfe
WljaGxgTGvG2fZsdydz+hbxt8ghjdkCQF0pXl44LTNv7ljmVVqVFsuiIusKU8tHr
yB1kk7i3rOAtwy65CUtz0GJ1DXd5CO+VX2pw92ybkNycHCS/f3PAbSWYprjQ8LSY
6vkCcHp1ZyBjAtK1rZ48SAIk3nZMKBPK9BtlVtBvP6nQFEZiTI8LrDo+db6CIsGZ
+XFCQVLSVXv1d5LtRch64R7vPItRl7LErcUDxfF/MOZnLKSFk2oxYIIF5xbRcvE+
I3deFt4CMWzRiCk4CIeclr7kK7Pp24yIL/gr4/Yi1RnCGwsQePNe4Vi4asXlS1DG
G9Z+iVBZ9djfursj6QYSlz+9SckTFj2sU/SzrPiCFIAYzwzjYde06fdvBFTyi1Z+
L42gqNAHcN0HbxvvNlATZVkX/wPSUjUrN/t8gajW66CnIRg/xDmvY4TbGdsckZlA
Zqpp6Pu8/lx1OqA5K4LB6XpxM6WLyyzH/+pZL08QfecgpCliH/o9qQSblNrWQ4Mn
fkWJRcXKV2AITCTZ1D73lYMSCsiwNiVuIExg8RrFZVr+Pq5GaNyVwSc+tIOYVJ4x
OOCLbOaqojr8KmJ9A9qxgKg/mTHQJT98x0NHQ1RUCW0qV8lB2HI3K8K2ja9A6yeM
5VC0bHpNRBOYyHbaHIr18NsbZDcdZJplgumjqHTCP3rosZR3sJVGYD9wHJTsewBY
8gNTnPTPKQXi/xOzj/u0Ws8QE76o1PA33dBepHSy/940hNS92i/a5N5a37aFgXi/
8DYQJnJfD9zwS0Czic3UzkAIKuNngyjpIP6X3qc0B2BxH7gdAFi1MnvnSQkxc/dj
BwC3vDNuOkNUZNRSa2L728KwfBNY890Fm2Ft47Lz5BOgEtdlRO/WQnZxYjGCgDYf
iM4sn8t/+Av/SfKNXUWytenM27Ou0KQJE8uOrBmNOXMNlQlIhT9DfZNgb4RBloEv
pLIyTcvvKORqHhmNfxLx6zG0SMViyKP34KGJWWcWfzoEUsQmEFQn1yz7s3hwjQTt
mDRoRlfdzWVBu1PClH3ij6DDuHs9FJhi5IHEhEu31OKUrwZJtsLtRUbUFAqjq8FL
U+OmOFbDf1vvt7kL9y/noJUb1JXAHIV70q1nEdezBCrqmNWs5cGKrQApZ7hAFUKO
1O5h7deVrW3GvIb/8z3OvOtEPg0o5Fs6aiaqC5dJPXUnFmnZIjylbKFJw0p3wNPL
AP6f5oC0jTGBO4vyT2UL3m2uV7pqWw4vK30X+PkY/EOFgss4FnrXmEAy9KUD7Dbg
mbSnnqMbnWfI1dtYHkt4zkYVthIt0UqxO9WALEI5iRjDHHO5BVrlY29dEwu1bPIp
j4agWn+8yxN4XXfzBic5ypafV/CXgRvny0bBDrT9N01Tmv4f/BmHdGE1gqnZfU33
dEV/DjS7DAc/RaXaGHU8B2QIY04LyZsiFFMTeBZWAboobuhRO/2Rcl7iZzCywADs
FAOd1uAjViJSKNDjHAIk9V2SmehTmR1awMSfRpig3q8Gaq4MUJlMF6WZcGqeylkV
TdzHaV27YxUgAlnk4g7FsEjDmpnbjH11SGiWDEHrwF9ZOhB3cnf3OrtXSERJ6Wwh
KrXdUDlpLI0y/MDipwZVUxo7e+veX/dg5LRfA+H87i3iGfOnsY1WnVebwpRQqbL0
1Dv3rcMzKjAMMUFW50SXAR4s8KFl38AXi7PvuIXW6TOyUSsSHRjqmMow0eFX7tYQ
n+2686ec2uorqBVWigezou2UsejAriRXprg3LOex6Lw5+HaZ/eybdgA6SeH0o5UL
1xZNlt+hZVx7+tk7JwvdNBW5UzaQ1eOZETjhoStKma3WTUUEo6xIDL3SbZivTWQM
sY3SvniytWI8QLeJtX/LJmYT4IboqBB+Pn8zx4G3uZTz4j8JUubu0h+2VwWfz/at
7FgHfRen8uUMAQVv9YeIlC51Lav1jZFsvD8sl2Tdqs4d9VwEYmhO3tFtrVgnatVL
Oxv+51lIrGtkp850EoZvqogrduMX9ltcd3KIXRXrnKkaxj8DkDb/UTxN4ZA3ZllL
rqMFoQPAig4J4WOZpqj+Zhboel/RKTP3bDb+NvPX9VmCQhvrd2sBOtOXoZJqBMiK
orlvj3C0xNzmNVQRvucFowDRq06gUxkLi1cnUjRkiNdcS0mfvJja5xEidKpcIzaD
rb4DOWEOGaTVCgaAZi7UefDmnngwwdJr/sOcJuKf1Yb4oLtzo7L/xm8IITOExrqF
iNvwq6bsryyuwMSGlOSgrnze7scfkK5gaqKJ36bhYf2lG27K3QyQXYZ8FEVHK7o1
clm6yZMXLUPv1sCdpwcA/IOknInr7047dS+2nPQrJd6ql1fKSslZrSe6m5Johx5C
t7BpYnuseI5n2V4oIb0+tHRmIZ22dKUST0gVOAvO5ym8SoQNvGjIAOGxQ2mEalhD
rdp9AVeSjRqy07s7F4NIevmbbU4tc/dmbPWMAwKYqbN6Y5UOn7naVsVftilgTgdg
tBgljDDdrxAHREcAleVZtTaTYjYEbub7qbRKx7tEnNdKIA/bMNdLXWJ8AmTTwhWi
TiKJdpD9GBybXH+Voslo22h0RJ4bng3bVvcYyZCx59AAHIeWsE34Pe2xeOuo42kg
Kru+7/12IS3ssRFy8sH40NQB1vJswvEwYktI6Lnyw3w7gkyKqajZM0+yS9V+xZmu
4FxduTzUkYj4Ruq4PebY1WpH25LnXEKBUZ08RsYjHS61hDTgrbGH5v/8N+1rofSH
FSlWQtDmqSHlxCUH+v/RXvEHwV22CVbj2avds5DkqUyKin2gE7s/oWhdyOJN471H
DM/U1V0BxVCWE8FyNQBzEVyp6nt7klxoi12zpsAstGxjTs/PxP+oo1hK+uEjyUeK
S2GPR21kKpC4cDhSH5/D3MVYIjIirorSPglt8+6eN1tngEwViA+aUEZ/+qqT/0NH
joEAgeN9TGzHlY0aZT4rJSumdQ7VoEH9cgjRPWtmiE8VFjsTJRmUtJcN6RTeNJLf
NO3bjVv63R+OG7c9j79jtaRmqOw0AkMb+jZMGEcyv4FL8lvXdMvH5XEH+isk6Qto
7sv4X5GA36kIq0uFkE4q2AyztqKbPjzrgQu/NsRDF9ea9LFqWO4aDCVdr1pDbVNg
O39wvJ1WU0ZLCQLkpui5hh14wtIh89QK7Igz6kYGvGWWH3XAUFgUxpBAMOHhEbtj
QgiBIBJvuMKfoLjEvtcYg9FKlWDZ2Yf3/BZwMuCQNyoqwItSap8UCvI7JyOscpzl
fnFbdaD9rEYIBJv6VrSQB9x8zLMSe2Obd6ZXBmIpb20kB2YL2rZJ/EUBOtjm7B5+
5Bl+ng8KLItTcM2WoteAaM77iG3ZMPXbWHZkx5dxpBVXd+zzmAh7uvldhdy4P+3H
qYH7iau/VoV5vbAwCoM8GgVjHTbrWE7KKxHP6yeauUjFW504JrJpF/2N4esHqBuz
4HhYLZxnIUMvtfpfOLD/CN6ATVHah61VROyM22gRUwjKpxX9XTlqUntUSInQ4KZx
fbVShPxfQ7idfdAcE4QhKkhRIMPb41P08312irZy59YJ1s2vNXWQgzyOyg3YhyNM
OWMthaxKW/N2s1jmlF2+pQK0FiZ8LAcNWOXc+h5ulo6Z/3iYmp6hg2Y7Ah62Gi/c
Vtdl1AarM9ZyPWOZXtXSZA/ornecrFXBdqFWUf/+Gurll/8g/y0Mexm3ui9s6d39
QWTbrRxy+ToB2iRSgy3vdJ4vDBiCrkpt5M0HNVUV/Tku+AUBDoYiHhLSRBpFbAqL
AiJUz2Q9e+pG03+A/iQCeKcQuVqIyqep8csLmnzTNwtwRwhHoNgtuWE39KzsVzRe
Z7WikU6wciKKkit1LMzn77rqjs84yGxM7XaegU+uzPiP3P+jneNj5IhUynztrGoO
dChDJswbMDdfCwHvnucPHt0OrFIZWpv2HUqpbeYPe5kYXFxek7M0Dyu0anf0eb0f
8XVdW8lfwevoGDJpRsT3FmZ9l5GcjO+mGdgkOwmJEbAFwFWkZVvFu7Dm4RvWxVHs
W8/i0HmcSyCwDzNF/365qD9idm/lEER7P5p5Hr35lrJIPmdken0Gq9j82S4O9jMZ
LrDeehwfGkFJxHZP0AdU14GRPiggWuwvCbnR1k3T1fAD460Dh63JZZJb070QEY3+
DRXhO5nS2GjL2TrrROBtALwwRb9khGmLZ0qLuU5PPxQ0ftlvY42T+pCFopHpu1tK
M6R02OFVf2iPatl+gbIpd32A/6qbllAa6OrCqZAq94GHuupuE1Vi/Un2LZ8lC2cA
an8h74ohKZ8Bm9QLJ15JLUQe3ov6W0Tdpj4GW0nFK4OhaR9bMclYrx1mljsYri7r
umAR9mrbUuetAHBg3KhafzXTwl3YbOLJkccufl2TZz1lgTE41lCMesvesLLbNiWk
yqe/U2jXsv+csIjW6DxP/Cbci9b8HKCYahRjjH6LsRTvTYfywRcO9FHAiDZ5oVH6
DIGXERwlSBFAgUPSm/WuFDia0hzt7ab5t8Q9cbwsKqUx+yatnhuvNXDUH84nkMdD
S7MnBNv3FZJWnNiHRo4mIbe/d5AdrL4KKfKgidZygXGxa2Uglh7uTu/ffk7jIPpZ
0uUkHKu9SGRlqmAvNlrRsAJnPzR6pXBRsOe5FwhYBPxoduAi/c3XF4VLj7GlXsd7
iBkEwlUKTJ8rnVvMwZnj7CqYEMkYEv3rJ3J/UHoIOVmCPejCHczpKJdyq0/Z9GoK
WSCibTKHUhhMygp0n2TVJCuFymse+kc2JXxkIoYnM1jNK3csZ/H3H/sZZorCKaK5
I2CUELJYF6rxTv3o1JDLGW+lHcFbfsh0xrVOBRO4PQnr/sagVxwmTczr2MpJb6PF
P9ZOueBke2VHGq8yxO5X+cv55epDqywzB9TDYvYx0StBAP9tkv1YzviIh4+eynUa
7vu9jnuMOygoNpcEuEshhrsvUWIOG8OOh0wa8yjSk85iQU0eszGCnkL9jmgvcceu
i2DgmWR/FkQ411i7/w/HO834ateBR+k0Hxiv8yg1CdA6e+wfTVuH1mOsL9Eo4JWM
RYZ0ZYE3v0A0l/ekqPzSFEqAyZNJjEkCGOVumlV0/tG3Rle+oaeD9gyrsK8HJE9p
W2S8YMEVRRCGT2cZ6ahWTLrk5COWO55BMDOMf1qiyIYfZ7/GADzT+G+AZ/AMwiDI
TFJhT8Ze6QDXCaSV22Ody8z4/U1qVAcxLgaalwy+gb0fHHuiQm0Sx6bMMWl7c4VU
tw/6VwlPh9HqIlr5nWhqcfsdYK8FX30oxLa2DABFo0vAdCXO36MPWM1qHU7HTyti
nt6FoiQ8oh/JUu5RJJh95Ub8X8c5nKxQjc1LnFoe9Xe+WksAD5WGGhucLv13wCUS
53Jgez6PYQuO0DV07GYvB8b8fCAXQ6SMBmgdXHOFjuTI3gH86eayOiiswGme+pv1
19uQrOKOkQFtRB8McBhwWD/LcNOO1ylTLCNkaMCklQnc8dos/98F/INNgbgHhwdh
iQYN4JS3bMRLjEWJcXpLGpn3fYrpbu6MiaP1JH1FAZxZ/T3wmO2/eXsfNLAaQf9d
sOM/tYv2H5z7KJ5No+CXtxub389DINYbZVvDSdFRPGzq5CBK8sHlTeg+kGyWA+SS
F16pQgVMoMUh6rijYLQbn7NKSj15Wdu2fnX0tEGFv1Rlqlw6SrO1haeltGv9dcsI
9RtIRLRNuDl2m7XiywcX1qc0tT5ISOz17MTHUCbVbQ6xVBs7QxgrHP0QBABsL9TP
rQAm3nA+CqUHyRp89g+i3t+WnG26BD3E56H8j6CJdZ/QOHmqQgYR0soZ/14zuOHP
pMIKjSkyHpT9ftUZFKecav1JAT8pXN9TEjO0uIxuj1EccIrtpYKszmEUvGuOcsOu
MHgYcr6B83j3JZKCDNtb8StJbaiXpb+9DNfL3V8MDYgiT9+psB9aGtFYJcU0PM8m
yq0ta+v+mIX0ybQszhlnRenSWPez39GhtVR0BQhpPOMixWKXD2TOQ3xi2X7cTWLj
IGwWzVHtoK6v2y5f42/w+sp+H34j7L5KKTBho05f7JQJvaq2DQoIHEEdKrCsyVFK
5B1YjgFB+p8jtLmRbbJ83qkQQTvLgQ/1XhwU2nWf9rs8xCSFAmnbOX9gn/2/YChx
LAYDh8MM72pQ5Z13sOtO6VrqWhn+o0m2UgbBGtJaUxEzXoTQChnPE6H67gHi5JLy
UkJmQJSrkpSx7lhILywVbq0ZYkd2/hxIGEsiaDA4OLLVVdRpyJ94HF2J+rm1ELVM
BfA/2f+XFNMECz//kuL7ZVz/xoCTGBVY5JnYyNqZerdBVlZBmMVAGBbDVnvi4Rb+
2arHqOhaC7SiGNKgHomLDBcILT0O21KQ4WP9efqooTkOQEd/pqya+KRRrfKFq9Q+
enasmlFqsrViq/zzaGaiX3cPirlF+CadTo/ScpWK1LNpRzSjzTJdVvZij9MiQMxi
SbIm0G+t6m1J5RCazDy47GvTquNKBOf8++x0aCLzstf8VsiMimq47j6v1FSXahnj
zaDPLGnhqh+9qa4Gcj1nRisfgrbQskuMu1WIYNf5cvipbovvvrfJR/6ZkAqtzmO8
EJi1BqrDjJkY8t+Rr7VsqZmLOqJ7UJE08IqD4uxPz18Colc5xoO/BILt/DT/Nu3g
vWZ8/tOl1ZfgNeVIlo4xJ9CjBEX8QU9qff8RXYLgweOmYqERhm5QQq0yzG2NIcHS
lXCo8bnB25iyANJlwFhLpWbTWfwtXqdqTmo3UVoxe7KczyD5GWal3fw9TZ16HYXK
mwmuIF4m0I4U5WwIoi2J4huYa6+FrnNEArOIaWKo0OcNTbronv/oO1Eek2rusku+
NeKLsIOZy+SfgrnltVFThDBPluxhA2H2QEpL+gAyLy6jHLyuf/OWfUna7CSboXdO
a5dhRmf8ohwpu1XwtxalsA8puH7DHZ3ajGjxJV8z5OwRdQrftMqmLNW56guIjb4A
9tQEHWbBc//RczdM7HopQwLbyAiMnsTDlcyQIbq+uoFyatWb8sbuf6VRVEk6YW5L
0J9Pt3lHZQKWsrjo6DdL2eLGabWE3UeUL4Zwl4DRdl+JAuTPyKiGELKRD+rOXMcZ
VibIsJmY6l8qJLUWXQMG4g0sMQTeVVexqTi2BDKv0OrlKx7lufoaotqNGXMhjSmE
B/F0jiwfftZyUHz6l05xvIdffBIzdu/Ro1oC03hwMngz1HAZQKtd5Yf/cvJd5Ul1
yKxVfGW4TTuf4SWENTMTjCX8vvNCnwUaL3drJ0h16nRxfUAJIhsHhGa50jIFTizD
kg/e55C32LJgzG23EaLz+KQHnEm8NyOuHwPAvcmfIFzJWYVdh8vnf3ScjHwqngsL
Hnvw5DchAczPQqrM6ZMlpB+eD/YfwboJ69dEfb6o5fZQ4VGFlnFrUOEpVTJatF0o
JTOJLjttszuTNlGTifEmR6U4z/rsCQurO2rmoX4a/IOHp3b6nf1HdJCjAMwz974l
trwecXlkAajP6X9fBdDiWpHBSheFfC9jSuSWJorzwMa8983aTZCf8CaYKDpcCeMw
2vumW2mOSIpZRVCqFNlPbPDj0YzteHKhZbpdq/7NZgLN31auPHJuNkVjg19PRqF+
Wp2vfTmQYdLTUTlRgJJeYTidHZntUiakxLHEm5xr6Fh7mors8UIrM1QP8zFSsW5v
XBcc0NNuaurZpW61ifSaPIxk/t7nAU29pLF/+o+Z8MvagmYyEBHBNQTJtYHV9jaB
ujwxDdfkerzCiaYzyX/v9D9Od9CtQKcLVI9x3UOOjroQgawKM9c7F1oVYawRDgid
GZZqmC2gMF785QeAnWDJaq09xsx+vYPbmDS68MQUlnSpRGk8kDUqBUW31HpwZZAY
pFENljiHpVDp4Ky/vS8ghOMoboiTtKt4yUzdRCGmsZKvK9EFwY2BHqKZIGSA4NL7
s8mzNVWb4S+3KD01x3maUDnGGMrc99jM3o0NeNeweQeyENf7kOdlJIpKJ+J9vDCc
TOrps5LjpYWfRoa4fAU7O54WMaiywH0vDX1Hg8TfH0ETnW7c5loVNou83KpZl80i
Tbi6JjqXGffT7M7bU35xZyBr96GPZS1gkQpj7TlYe0QmIT0gcDSOZkeivaO13OlG
ytLTDVjzeA/rmRJNpofnRDujJkNoatdO6vFZyyajBcFI/T2aKcVWPnrkdBpnVSJl
9CT/AJMZaLskwTdVBC2EyaFzRRK+N99x1NOWny8dn9kAcNqq0EQgEL9f9PxY6vdD
kJch2iW6HfWGNltFjd6PDFjDY+xuyENR/jOvVGZZ2mMZY1XJauH43rYNqheIUojJ
sUffe50OmVaMIzISnbY2esQALrj+dhjnRjz1nxBTIHyCxu0x0juhkvUV/Kja46sp
qloMuDHgvOe7cSTBpucFDQwIk9y9QIG7ckv+QNTfJshKWKcYy9dB4x/u3YhSCpY0
hixrJ4c1LcsgPFtzTSDbzXQuLdYIhKG+UPftmiO3nMhwDIUqC9BCfBw9jjbDwE6M
NbJFMS222RQ0dfY+DajPhcCSa7jmXbjZ6AtBKt9oq9mJJgfJzZ8aOHTzX7lmxckR
niEDKXL+r4CSbThYQ33jmxs/gfJR3/C1IEo3FiW9kfqW6I0fCAxzpOPhOtY3jLh2
0t6bdBBYWGuAoFbe7xO3DXgNffjz0nRN45xzMlc2cIKAXKIo+XM5eAvSfnJM+3xE
nGxuOyXS9vsjBaDtxWB0AfTYlICYuOQAi/nL8MlzPOZTUaoLRE9iXJBQbIgyCa60
M8bYKOnixwLg/aRVyISVSM6aQrVC2ufjg3q0DBZDuAL/mazcCTKmjGg9UT3Xl9Nt
h55VD9Uahz16NYD1EL6mqc/fVPA3BU1WqNt7RXIuiJdRwynstp1sNfJQ0hSM5ZtG
kX34zMcchpN4Zx46ek8zDDOY0VwkCGyfgLpCygti0HgPno+VVBxz4W+56vZ/Ezhf
yDa/QtBeHdzUs6/bgK3R3/rHwayJ8i7L4J4MvrvM8oz31g8IZZBpM1wvVkxQOYUf
nuvyp9mL1fVXhaTfefpiAmW79rdMxQmHLfMqbIBc1pQ3S1NN/s8Krsg72Mx+/WzJ
JxXZ7eoVYOJyDOJzRyXAod5WbdNI2LSyNe5UCWH9tDAlBtM5PhD+z+QZLSTl1nMg
YH1E75iqfZPTBD4opNMcMtNV78wD7QHASupigpUMlE7bRzHvvp4R9MTDhdf9lPl5
x4T0b/MfMKrbSmMLQxNelWxqvYC9rYd6C+dLJgus6+k7ZQF9BgNMwLgO5KhLs/3C
/JZMFrmYOlHwPG2bvaxOXm00Nf6se+TuR5Hf3UMZNsGd2zgz09l42B3fnaelqRXB
oyW6+rjnctCTdFzuw8ev1t2npjvbQb9WVAJIzJP3kfb0SYcK5lSl9bDOs6q3qAiF
PckgxmM5s8GbaGCqG9/tT0qSASzWbOWcryFyW1lywtv6raFmJTV84D5mCnZ5xORL
mp+5clKiYNMQZomW+GWs/nKmj7/fSX0vKV1QuPrf3RQDtdLZbc5mZKh+FAI5/myz
rje/Vpc4Qc98OqQt363YwsGgLvOPyWZxOh+95sbXuCnWlx6ycDwAf4k5r4MKbOMx
ECeIx8jm6H9T3gm1wsE/LJ4U9wdRB/BgTqMeJw8pTP194q28g6Itv1kw3PnMcmo0
D8BPreIAEQDABQ2c+VDx3LJOMkiHDbArzaIdePVTCLGmmY3oX3f7draPT8z8IP0i
wJhVLsy94T5R36zceHz1CSI3jfKJ/twDqou9UAGa0IjhiYYP+htBi93rn5ept3Jf
pqzEUWCV7DegkYHUBHTWUMbFkVTuIvhcVTJwnVBS53A6jpXnUqkQl4HcIm5QWSVN
M8UT8xVvB6NHEaf/8RDZrrT8QLZY5u8/loz73W9aN9Jtyy/Kt/HymqRX3OFscXjv
qPN6RR0hRi49zyDOQkx8NYIoeDUB86EnJrpn+S03y4v/F3F1VOEewxSebTUVRPvZ
6GOLjfD3xwwdAQUqZ56EIi7rVOVWLOk1vllH7ehNx03NSQCPGKAoD9d2mtiJi8xc
dX/7RDqx4XFDELcgdtJaPtlcM4DbTooUql4FJfFRjPUcmFl9k+E95JwShHMIQUNp
t8GTIKF3BaoWiEI47myGWs6LSKKlm0/hyYBA0+XPoRi44SemA00abYLERQLQp2md
XDahmJTmskizTvWUnMSWnZDKK2zMvQtZkKx3v3mXruzvQGefP76PiuPuxk0iB/R4
nXpLhFU/CFgMqDrSrlAR4SKRqaars/OXiSYuSkPjH3zq8dIfkh/bKFAjReHeKDSV
E4skKbYGZXxiimR7gv7ArZ80NR7QQ0pWqzWnCTaEtq/F52nlLJ38X1JQ1j5Re9/9
rPYrh7nazC8+b14NW9PRpcLs+rbM7B9SlLZddPmTZnZlPFEcTsHW+XFuL2qwnesC
5FgtKrrFGBRvC+ZqIQ6n50k4lHG9SZ/yH3C43LSHm5ZWTcokhcAYkysUnj9cbPIZ
fdjQyqQBoO2sYDVxpEIxmmt0gyVXdc6br2cevMrCk4a+Ub03iVRKPHzjnK5BoSES
5e2Bf5L/A/yqxFdONr8QsWLz2T7sE3nCEvrzzsEbsIK5P2NW6vi1ADNCXzCCHWVc
6IweMHSZASrYoKUCafBC7ak0aJOE53xEk+CLQiTiW05K/e09O/CKaBzHjK6BqeL+
Y4K4OGUlNezLyfgOg2mXEhdAJxSQqzi/UUVlcwGh0NsByPa0s1uOWdYfOatEVEf0
fke564I3HpEAuEWe73BNVGskjXpBrxCJ4/so9nalPKapZl5hp/p94sQBMOLqKnHB
3qq31CvCUIvkUs2GzR22kxN0I2wfA2+FeoyTNC8nJP6dGfdpQXGgpLrWbvI75Cfs
Alb7WSgBjHeKtbfUFkJ2wwnwqn1B5CcpUl/Yz9VxhSr14Wkc8OvRbX2tFdDlnBRt
Pbzmb5Zv7wA8GY37qx82xZpSXDjjXtdwXAYtbr0nIO2iLchzNLP6PJ36o71bqshx
yRv0FIfWxjBMcfRfQLPJp6IO11X6ypi3EfSsyWEpQv8a7Sd2Bfyn5Pjv4B4PyeGl
+fvHVE9/bPV2A6APNz7+xIHGOi49Iy0j9UaUwC8pd+l9kkuveYxccpNusQl4Wosy
tgtb0EUD/RPNbKA8WiNP1IDcLPiR5bkJI/7jkARV2tp6Iip1ngC56ADIl2t9HtJt
5KHqYgSAjwyUkyED6tV80VYNxByefHV4gYWZmh0eiVeJZT//FrV/yp7FppPTV2XC
/44vze4PTngppim0yD3dGTCEITL78PF1N95jsvCd5jVZjL8mBGuJmhX2tI4Oeaa4
YGarplleu7UG/tT1jDeR8krSKwmtoMhs95iPvAc7L65xHSXWP/z0K7Hn1rsdBS+n
pj/wG8fxS0jhmTUSKhDovAtdzaOFLBnS2m0HCCIosqRX7AamO+CETUJmq/GgbIFT
40uAlT0ExA/zkAhyKzp1YD5yvxSAT0dVTNkHk0hNUGXWRsLN5Co3idEZXKx7QNSq
e9ugxiNihVT559UitTw+mbgpfjrFcslgxHXyYyog/mqUnzXG6UWZWjugNgTY72U5
gN6dZkpmfafgTDg5aQIqVuD5V8IzpDYyj5sEjcNM31Ges0jWnBn2GYBTxv7PQAiQ
aRlpAA+XYfjSbYwt99xFUrIZllnE+oGQY6WR/zdTAtQsw59Pak7ip2uKxpijgOte
NWNGBNBVv5YB2aY74M8cTPCBqD7oZhw24SzYGKDJBaYHUcv56uQCQ1XWbWksnWol
Fc7MTmDbaf6h8SMnL+vS0zS5S1bByKW9FaJ6PaeqvHfvQFfuSW6mOQ7T6FRknBEJ
4o6e9e46ZChdZ8BQ+eIQOISa5IOE+VMEDpf+Q12lL1wAxSf5Kbmp6x8eFVhB8R4w
i9Ys8sBOnPCbGn7+ysM/4BadZE33TD8WXsTJp+IdQIxbBXy2pNhLL8JlRRizN7Al
2+ifJZq7W0ufw6jylxH/kNLn4qdIvV0MoYzqGzTDvMkbuFIyOER+oOYIGyxoK7p6
mQp8+DwUbQgR6YWSGKR6+eNiVy1UmaTy0OFp02IztGkmyZlinyXxwELPN6eUgQR2
GMtpM5kYYbsB3FbtesBxSDwJJ8ZWnICxmSre5wHYHNUP9Wo1HOFH8/rQuJOVARXp
R3eVGl2PVD/kpHQaLL/VK5kF4FUjvWFxRps+2PM7HZ7JZi/ekOTO9YK8Pk8UFyWy
Lvt3BntIQINEYJPOaLfNucs4lpIu4QYgwNbktWIEV92XP9FoWjU3bfyuNTzNQg7H
ufrj0T2Mb8WoISXErLWkJl2s1A1/ywLBM3tp7pubWjsfShiUtqO2SAVzTusj3AK3
YcmqLxaUnKcjYIDn0QqPzLYrgl1v070F6ueM4340fRl2TyZncanPDwHq26euqml8
IHFX/SOj9lt10A6I6KIvZhBzeQ8ZdBDa64ba9VKLtaDIGLvCML+FGCPQ265xVsHO
6f9nOD/1NYvZHxeu00Y33H7OxwiXF/zsp8tjThG8akzm7r4aHndh8nYzua8dkbDc
YyBk4Oeynd+F5fCYLDoIOMj/0pAg5DUL4tB1OP86V/vl0cIWUVYMIAainN8VXg1a
KgLHlWJ9Yg7zEk0Q68TDGHq3pVJiUJvfSqH5p/2ixRnzgxIfxWZxK5zkuztqTjXg
kbPK5c5GBRvfh6DZS9S+5o06kCmXhjpBXsU6detr+lRrNyHUg+FOK2aivHAlyJgX
+zyE11izAu54YiMtOZhmP0UtSrnvZ/3bn+PQLNzmxtOCwG2dlTMNTcu+7ANRf1Ud
6J33sr9UEox6dk2PagrykhE6xQMbjEi6bpWBxa9uFiPD5mhyJkj5MdxlwP5RcS87
vkz5VfKDD00uAytpunelxQckzZZ7twl9dcfLGATQfjeRxSNX0uA8Ofkh1OAo9D0j
NqRLloO7c+sDwssU4XazfeG60nM2qyfgxkjYg2CdWsaqYGgXV2t93Nm8p6cfENah
z1L4VVjr0NHpTFtZCSFUPLvRQbRtAzuCOVWLH6H9jAtSfPjL+BNUNo4iFGYf3WiJ
CbJCB/GIZxmCKp7J+YJs33uDHY8QltUSayVYVVlPbX5oEwgCFqTiY48tFmcUwblo
U5MGexIvSXGOjdKRrwNF28Wc/hFNsz9KT2bxE2HO5CRkAcpbj0VyQvrgx63mlcAS
EWQ73TYbg+WV1iiA9+5Ji87fG0NNyj0mAfml45ggEsznJTHkuctCPGnzVdHyXOJ2
Sw1Gu+tKn6A1eVpso1rGLemD2XYTG5zS891X60teoRAaor4+Le3GLFlsBDy55f5Q
vlQCXWus/ZezmrV0YT8znAesK4ZACbvsLBf+2mc82LF17ltr1Vl+c9OMchJztxvh
cnTwEvaMcm7rP4ECEwMvI2BDgdZdm58hQcO5n0ACHukQusJzyX/pYWpIJeLyDpvB
2LnFNuMYA8S1GVwPnizB74WyRZToVJJ1O866sgZioS4ysNlp1b2EUgNfRrrZ2A2O
qWttA9xRR3lbKaLdIayZCimJBOCe73kF0XJu4gvFbs25MFLtC3oozLQMNOOjbBWX
8sEYbnOTpRKT+qouWyBP6dZ0l9Cyvav/OEuw0JxgPaS/6NmY3ex0nBPSrQU+YjlH
XqI4aFh5A/uTpBZfO+Yng6CNVB2zi++yfEbfnOi3gL0ZbwFd1FZFbW3PQsJlJkp3
glVcjRDEpBRq9EVl1Xz7LhKT3WLf/K9QjqHU6o7/pZfyAmAD96HhnFZjkr4TLVpm
BURa0KWgZO24zSQwiRRFMYnAshw+Zy+A+SWPSIPROkfedbEcAfyH/vQizYM66bhg
mIPaJpdBeGni5Pcs47xlynD8B4zhGtyTk5qcUhAjvOpFNLCIHdHhpVxxSmhVtwlm
2G4b9SvuLjkqwPJtC8fiKsBP5WiS5lS7oJ+PaTeWI9mM3JZeStazUxJAK8CuALvk
EK3pn9A0jKijD01gLDET6o1djsjnRIQTtp2kxMaQHCQyjrCreExz/aXTFCqqiLTY
eq10P2rNQVrK0iKWObildlm4Fy69TQ/wEOsaCZpz8A2ilg80cMkxkUnr/fE9HzM3
zPcCY7hYrW6zT2QfFzB1ncSTzOUmECkAxtEkxX38B5Q7vhsgOCmV9ivWKz17fJIi
vASzxbrkPHKLoTWQLSFFG/JOL9iovRx8FHjDDmfGr9waEuNOt8AZqeV016a0Cytv
c0Dun1Ri5YnyXHIVSL4QgHtFCQKW4+nXfiDtY4jxU1nQeg8GhIlEtCyDlwR1veOr
EkJffVvA9bKbehc3amkcLjV+VRHE40U098GQfOhnHF0Bmwx6NWJbSSO+tHpnVtzu
HXSry6NwNaE7unpMFn8G4yExM1oA7hIX1y5p3ev9ReqFGJux/l6pAIY/pKDnEqLf
Uijg8hf0D3F7qcdGwUQJ6XzkTRQrBVV/dxT8kOvqW9eA5hOPago0jy8/kc1SBU5l
CEZGQDbleSDX2FwZwv4aEvE7rpP3cJMkQVzOKneJad3P/MPWntlUoBsHwqfdcrkf
B/n43phZVySgldQpEcgDPYnQoU0jXt8toy7+BEIPXh6YH+uQnDYxbSKBZyV45NWn
DE/tl2kL8hKW++t7rSIL4/ocw6x7Ft2pvEPnVVLNyzIECVLn+5HFi1shgQ8ke+sm
jAUv/4MoqZGzQGrweDzrmPOErhSo+tWAnfjJ8pyBKjGrnPZbPCTZSv6Nssn7KKqQ
Kp2wcB7rXBqxpVMUZpLxWzmQ9XacCPWjI8KLmvSbZCnVgSyPLi8A79jpyL+vA2Sk
lNpHbSHQAVHY6+F6Itbctb/u1wRZuwIs+GEUpOrKF262XlW4LzzstLiqqIHB3gQS
KEFq5dEcVmKNUhKpLdDR2wmkYIhe2jv0KChiNMnmR2oacFSJFOQz6M29Y3qlayX0
H341aOXFj9jYzfu6pGvXvK8UuFgp0R5iMBPDe+WfFyScKinR4kyZPsmSUWbTzINc
nBDiyGqQ2jKa3mx0MDldhsAQOJb4/PMs1bu6eTR3MVnUEHbMKSKDszx7BOYc534g
TuSPtLt5Lskz0/mf3GRMvNhw5v+a6RKT2KsYrrcajB1aOgd6fXvceUbGt9vW83XM
p4Z4yoWbaawnqm/r/DHkPDiGc5npDHdHkU8+Xa1T6ykQt5BJ2RL4/1xueOF4avPV
572P5MDRjnDSycT01AdANsIfao+yFLv6PTIHP/X7wnPNepCPf/y55VJyp+P2uSlZ
Cbvmq7aXVTU4euTTERy3OsYrnggKuZZ4ecby6vzSEf+zNdcpdJmpCJQsMJg1NGhb
kaPCraWW7bkrSRubPWej5JNYXOWs2xYlVrGYlRoz9ESKk1H+o3LcW6B5tRTE5vzr
EJM7k+PbZcTyta8l8cZRwOchEmcqOnUEdb4NeNlYf8dl8rS2wxCBMLp9pW3Cc2Sg
HDx18ciMrinDxf50Dl+GPnwkHb3JR8pSoWKaKfnAK+Jr0x69VlY6ZXAWNSQ84AiX
d2XU8m/ybwjZFUisFFqiV+lHacfJBIs3Z50C+qaY3mg7vF0pmMzcX1wH0FOCa2Sm
NWt737oaCDwMWWjzuFaMXQMD7RpyK9ONpFvPZTvh3TbmcDBgenLIN08V6XRnymDA
lIOmVt6UnOM9/9Fvf9gUbW4AqKxV68gaJIvdM7W9+fTQCjhMNdsYbzMiC2Bg3m1i
vwbD04QWAzgx8bpfvIgFI7Qw6MKvJHMLLzmR2oM5Ci7cjq2XU3m1LwBQ694z/udB
DZojdZblffzrNbHwZiRUb4HHWEhj2RQxBZADmyqiwnpNPGkHzmE7eIRi4smYRll9
vxTitQcUV3tyNgQ7Plel7BBCY/nbmrsjlCJ/LsmXi5IM9KeOFD33bXuGtqmNwroF
HRihKjtsY1Z+UuQ9QaWZGUP0koZx6I/C8xeEajAl411icIpVZEuN3xR0kVW0Qscw
hIT0C4dhaI7N1T9+VrIi0mLokG8M+Hqh0SK1LBaN7/8r5NOP7BzBcP7BvKT63gdz
YBsd1tvDlvNUsi+qZfjMMAqvZSWhagCoSbYZ2lwxIfSsIIi/YXOJ6JqlRVDFmins
uVZLXMt+piqEbJJm+HQNrMy1/TMPgzljaQev+3e3/Ju1xaG7GwgfqqMzRFeQDTsX
T7J1dL+6VGTaO9GXnvBx2Ybj5WkzMmYw5jn0ea6O6Hcw7xIwr5xSbew4xiRfzp7R
By+HIO0yxIBDBdnv1n8mkUDTZzUkGk7UGPjNy7EfnZgO44urhLirBZXeo+xWp7DO
G5MyTkusmFNJMkLO506J8MBM06HluSJWslfwIurGYxXGI8MORxekGqiaXrHalM+D
httd4on9p1PWwAYxXlg33bMRETB9Z30ZVXMzb/WMWSK6HofHuoZBEgFJ1BipX/s8
qe1QhB48Z5POxG8xxOPWdfM0IQzt5fZsOT38rq4LeFWGnsDYxmdxMIjx55dW4c5V
L3doUzMBI2Wl7+YfCU7dyd4hv54X8uhcHbyYZHCjdoEJAPr/QcZ2qreTj5PRfIga
z8CJHqlwR/6B8pQGwlqclqxl9l+Na1rZLvVZmCW+oDeq0E4T4Z2V8lQz7gtaXTxM
2db4U34rUpi3RbNgHhDNfzXWoDg0V35hIiiprurCLJ7LAeqkdZ6LoVhZ1WgrXgqZ
rVfSf0yO45ANQTHKsnfgIwniw/9vCEPGjToQs0hdxDoJQrHA+8FnNN5a3lxVN9XI
xqIeeoOcFUZ6PWx13w61eD372HrZzWVJfHgmJ/owLREB9ulwp0ev+CMsLdb6M9u3
8kz2zRemncTJxytTZYgJ6YYYNp1DWO3SvhAKLIz5KUfuZgqSegUuZSl0qMKBlQrx
mP2C2GfmOzfm/yaz1B/hcnqwA1hvvKPYR/gH6eK3HUXuXbGwO7R9s9lq0xKgfIh7
k5euJqAK9CXuVlUI+OKvPInqBez3qAPvVFTJ5x/A9FlcqpPgzCEXVuwTPVUFZKlp
ZdohJAcv6/RM0W9n7t1xU4fcH3RKOodaSzW8Fzg9cTRDXR8rI870sSDC/M6W00Us
lZhTJ8Yfp2BmOGhS72V/DzealqDeVH0fLqC7h84wOEdM3u5ZzSsU3nVOhbLwSDOx
AdUyK7bP4aghKIg7y3tDRfdnbDSUlfxD9d1zqvn9YaNnoQYGa35pgUISNvBY4f5n
hyFi3vOK+2JtC6+r7vb/wEJecv/YFrlcGIoJts2X0+hQtUhWabrCUyZR5baa4Z35
Q8zAfpS0Rh7YBv3vP22S3cmBv6eVak1x6ktQwU6FBhVarc4gdkN9VJC7lcqDLU4I
+MFvfzlFi0o3WuWUOtCFcZCsn5GUQqQ/P3qUwPecbVKz8HT0QtPkixyUSDdv2YCl
aUlfob/NTCsoVL7WTQ1ENgdFiyxOjjWGFx/lv2L0etvqTKjnP0F4iqBoAy6iQhWe
rVwBkkbcmkYWN4m9qmnrMHP1IEqHrzvB7NjTKVobyk/Ue9Tln463HVIcI/Ob4nNz
ijyIlqPG/Lg8cHH4FsCMRNR76fRhGi8bwevwbC9c06WYUr2DlWOln1DjdXQCyVmo
u0cXLQx/rIfWp+kNTSiSsu+FlDvy2NkSPc2d0OQ9yb9SpT7+ATPEHpRl1ul85z1m
p91KySaaI0q8vy4BDUb2wPP06nn5gtT59Dlf6LK7ewhrdioEORpj+hzB9jNz2Gzz
P5M3eZFecR4y1cJu4tZLSDKy8dwvutLUwEk0jyS279kF2JTD3v/6Vk9bJRAzJYUQ
7FXqLzyoqfDwPFw0NhQEE0yMpOejL7LZqp/IDgTbZ2tnUiVkiDMlK5QRceBQ5Go6
PuHJDzcr4OMwXSzddgQJNAzM6w24Y7lHdUpjy98bk7lDeNoTVvX5yKelvsb35UUZ
F6LtmGMX+UcCnOLgwxcrpch5sk96PpRy+dkUzkiQ0+ZNtpnEv7qfID/oylSCRl76
49ykV0z5j+rejO2enavo9hNEq1Uai++6ebqXkIr5yLEhHyw2jLr+kGzD1jdDfbL5
pRteFW/7c6IWuwnPTnqaJKTCuLtQOO2POy5QGO5E7OnH5IHxqeIO9PTSOJ41kvm/
WhXdlGhptYru+oA9ZZ4IHoxfcS48ROBVs1sXDNexcX94uowg3F7TFEF3REmFyY3K
5ioHtlfYoVzbFtfesX4bbxeYNeiDrnD74xF8t1gyd7mTsQgNsGrLEJ0yCNTu7/9Z
zSG1fJCLB35QO/DSBTWpwQ3HumOuEW3WUCK+0sYO/Zd31caXKXFrTnpHBZuZue7A
utC2HrJa65Zo6tx6lJ4AA5iEzeCFg2oAhnYwlrEmg5WittUHrtwHVTE8oMugxt6s
NtdtqgY3kFHyuLi+M2Lwp9CD/ijqHebUcVwAK4l4Cm3NWdTrQECnxsfNGjDYOF8V
zGKdyzjDPucnYHnPNhpwWblKbrV+x16wdX/+jzXWdQWQdigjEyHEz/nwaf7X34F7
ghZiFFlyAiRfyqex4LBj4gz3gKDpYTsZbcIJH5T50bsTY3LF5j5o3sbXp9H8y6MW
ZAb1iWeUofU5QLl4LSKbdPgKGvhbOnwPPtxpzlV1AhKocZRXLuuWJ/xg1VBym29Q
DPzih/9HlwVRczil/xXkoiJGqr6R6bDuOVT/zZ62FX2fzgQaJ6qM7HUyIpHqXaWt
gHKRpaJEvENlUUPDPrtdpxQaitfsy5TcAOs3tFrPxw4BMAPkSm5pepspj7bfGDXf
5VvYNjGywCaWfk3XunbxJfvUWhGD8vxHHA8nV9S420AttF+JDqysxLloEiygkFpY
lqAbzDCP5pFhBIrsue5KVI5axWN4IJDJx/nwJ1PI1/LPa/RZUOF8Apq7iBgFVwtb
IgtW5o0gD6WsmUltY2o2LBQh45a3xgr1ZVOA8fACcPZSV4UlQacMpwx/nwQP6sP/
hNb/iB8ydecQYGOW494IWkSs5E7abqY0N3inJRHIXzwjKO6fXTeyzsZ15Y80M0Uj
v3U9fgfIrkwtmjJLTwn6V72Mawybpp+++cxbnQqaNiI580LFFV9HrYGjW/iTLWu7
B67FECkI8dpsGkhZ6be2siaYjcQz2yJZwY5VtA4SF9sY0L6d6ratiEzwgyHGCxqW
ks5WI2sYGdkX89lhzjZoLfvZW1U0Kt1JRWBN2+ONzJ/wPBvy09whUV+j3g5hW+u8
CByEWkybAH5viHZS7w25E5YUO1zJPTB16t3llV6g0TZsg6hc4B6zARYFSJsKxtQY
H/N1SHRq7+VtvQMoDM05e0ckIv1bG5O1UgPe7ePa9hF6ml17sHh8uYWYfkPfT/7E
JDOrhFQwstvr/3qLb4Ag6qDt7JDu/45o1jkVoPytJkN5XX6IXnVvNu3k52tfx1XG
04oXzdSgIYcutZQ3360Mrd00LgUtSXrZs4UCwsikjKU6WF5K3EMZOOENFTsl0w3F
/qwhj1wwilCudH8/4v6PjGuawFny3iCGg4g+AyZmG1AXySPDJL7wAVtQXVcpQbmG
4gfbI1kSNxy7v2lEfxhStKG40cNqpyjwVLmzMMs25mmYauxEh96DFU+GcNuw5hot
H2qwZX6Ju13Pq10vvNEfbfcuEP4W5OSC3d/OFRdZVjn6uZ/satF7VSsmfot7feyZ
IBXPbejmZ/x6dhbRDkj5YKsRp4HCFfgnbOMcoWrmCyB0aXZHAXOyq733ZHSqIqrV
/bpAUFQ/nRhxhWFWDGW/GlVq1pL63ncrxB+Gko9gNADF0SWL8rtmo023WapMSVQE
tS3Aq3G81Xfo5Rv5m9yhaFccsNo/M34B/NdBGrg4ZzZMHEOYNofnXwcIDNiE/Xwl
JjlQvQyChjKu4k85vO+J0ZWokqfzgtwGCYSdCpB+EC7/Vdp4ZeyeNWn3ZCZice25
0COaom+Il3KGdLd4ifiduFQyCrzZiBFSh9m2vdjfrpx3jJj1I2K94DjaOVzr+3wi
vnpMCkxAbe2TYHHks5RMO6pN0GP/Edzfbkh66ItjjyQqD6BPSt7C9kpUOk3SFDg6
+w+31R06zQMMgbqA1hdT3N55bUFjGZ2cF9dHNmfQBfL9v1rTM1k6+dnQXH73usXL
NDTffVwfsgQX6wJUDgZaCUKQhAcf1l4CWlVZJmh6bd91tAqvkDgujKVxdKaiSvd1
/+6Yxf8W2yL7tFpZm5e/2zunDkcXTy54jp2OL8GlMJ/hTBzoRBrXsNfBQM0SZ2FM
NRnY4luHtCWX/kXnp5pHPXXY7BLCms2h7wsmmmISjygK/ZOD+hKoBKYNjX5bpSFu
qRrBR2E/HEG3u8ZNikn31SgTiTxwd4hkSh+6y/CcTXKf+cR3I9opsms8lBM7DJWm
as+5szm2txm/EUOX5DkwN5eDyWKvzcFxNAdnc36WzEx+gpfVAXbM2dWS9SkuqevU
mgtNo7AnboEyF1m5PHnL6BiOTYQ8o92bsWISyEqyCdz+G0ZwwBVtE6yPKOTf5OgW
JdGwTg2T82NmNN6hENRXtuYDjj8vSw1d+zAk4ThNbXR6GgTmQ1me1lH7Q6gXTMD8
6x03Ideyyv4YAbZBTb29CpwH+rSnOqIX/u4CVltyVX5dYo+Jm0iISGc8sI3V9RjG
YPYsNI24WDfC7i+VLPf9cq7TwwJ1qPpm4FnTK7h196IAvihP7dO5ryV4rRFMKI75
e8hG/SmeizaecjPeCg83C112BMfFIjXWbZmXe0IvvQjo7GReYewhjAN6pWtUCMCk
SWKkCIKz4gMQVfHqvcRfYL9KFUZg0yoVPXpmBD9ydilhT/LXGzRJhBorkDCQAkbj
IfD7YWINWg41HMtyZ9sslDSOcNhuEtKo/zNNPI30XG7tTWyAyWipCnKvNGhI/UJU
WGgk2w3uIjczguNtOVdJZ0sWO1UClm/UWNK9OD81ZxLiE61R7jX55YoMxdp966V+
UdyxVHrDaouvvm0b8Kzp9J0SZ/wIQOGAbZuupCH4S7af4CrKP5A57exc0cto+SrI
mI69D9QZWLpj0vZdfzliz+uO23rVas2cYsiFLoj4rW24cbIt9gQcHoFePhTSzd7R
c17Tc1lVeQaVY7EU93vfeTzDcSKTBOIwXJ+uDwNVdyMjUfbHYQk5t2FGROpBBf+O
ZGMFlWP6+Wqm1CbrRQ499k8h0vJmse/Q+ldeX+Hl6gsf6ZWBe03AHdUyo4jWz8+D
HXAvIvzsDDjrMpo3xLV33jm4u4n9ngFBJuB56QS3NEkQHjE/WcuvnCtmNwG1QDWg
zdrIzVxwQuqE85fKlYQ/SySYvk9rftM+rDrDJzSfXyXHv9D/iH70mu9lcAZmhqow
IaSjsjm6azGprusLCJOO+c0kCfZNIPI1oxnsQBQyquv5mVzjv3RDA32nkAXy+WUO
1zHZSGaNvxynjT1XHVG30eswEHMjEWkuyyYzypLG5XFI0BjOXXw1IfK0nArc1qiP
+TqfOpY4Z+W/ITyWgdfc6OSW5ePTvvXrdlbBy2I8UC2jvOHxxz/9Rz8mAPP04ADF
UPRf4+Yl1+xQ3fDHHakMw+XRnzVAGz40Gc1HlK36ntxz/ui/GpCLg6+7BI4UWelI
E9QqO8dT7jZ+kcQT95GjwzLETx3vz8j0SoVO4iayhLFbPCuFjqAKhBbQ91LXP2D6
4MTi3tzirq44NFeL7WPfgVOqaBuDHJTTrfbZjIeXq01pPf5bXb1sVaSCGLT/gkNG
sZ5XXIy8MkKE2wItnkWO9O9RWrndO/xVHq556Dq8jVXSC685D9y3aDXCnZQFEmU0
rW43TRFwY7Rm6mv1Cix01KD4LwhTHKuVUy/Q87ld0k64VZsMCgdbJnsthElx6t9m
fZhb9waOPg/41Fac9DHwPcjf71pJx8nW8P/zfZFGFGnK3kKigs2aiCJiaHLa2YF9
Ynh1sxhAATEp4S3jHdhP183lar6BKSsuPsk53GJScp9kPRNvvnV8fGp6Ng0ZMWsI
f84lyT9ekb2ena627G/dUULqJe2rgjMmUwniMWbor3pFxFivyoLcKi9i53j46wSm
wZhGj+7n9Igt9tQ2f6gYV7t3U1kU5FowEA0IOVcuKem2krGgBYCoVdyjDxVJr9rZ
gl6aPYJI7y7PaX4fKuP62G1s0cg/p9Ff+0ih+utpoNHN4JpM7Ob0Egl/zLAIIy1a
nKbOz3QNwXFh2sRpJv+Hy6s5qAIJs0LkBZnFIOgzZAxGOxWrn0B3ATKmUn4Kccpq
yPbBM/8BdcLKg7FUcZvK0OrmdGSyd5GdvxA+R3k6g1bs0u07XZY8sAJf3tQHOBfk
+iA1lhR64d8p1lDNS/lXzZXcHsxAMMGjICw6vpVnyevYwRev4OlnUhOyL/4ePki/
gXThBAGREvEE/VdSyaR2ZXj9c0TAKwEhToTWDtKik3BN5+O2RVagp671ypiVNDiz
LvgPwT8ASQRxjfp1Ro7c45dBFNoicYCDuVr/VKuoib1YnA8sUEuct2I3ImG1gx3T
9S/n3BnpAMNAo2T1oISggnHESzV2Pslng/slnSYgh0rNKHdprCjZe0dGhs13xqV+
3lrVCp14QLmKjRaCfnUuG9cvMmCFBKRglNdAMP+AU+uER4HRtPLqw39NAjVmDvCt
6sROgH3g6/mzZxXDt28CNHxWlJvJlBgPxAbX7j2DCnTD/Fz8oYuqgMxjWmQWDghJ
9XJS0FoqHf/txTjBUC92LZNGdqNns/NNTpnVz3UsZ/SfZCbGGW5zBOQb0rpXbn1h
5DB1DolLeyHK3G9taXJRNKEM9q5pISQ22K5N1QDui3ozFXFVMOoyln1nVerLlDfX
Lm/r2eHFps83eflRqkT/zOegRV4HMMOPa7aJ/73GynmpA0MMOmMCfC5oJjCG7tyw
3g2K7WR314C+425+f3Mmw5E6ngMKKyPus0ydr1L2onoS93ejDWMFNoFJAP3/Md1S
dmWSd3VSjHb50QM1O2/8ihjebkTo/35y8umQFrPgGJTdSO0tb6E3nYgNWOabXQEE
gHodw9dWVoZk+QEgt901XMlc3gVoI+i8/c+u5dJJZU/yj258A7jZqMFT1ytY2bCv
OEssqlR3J/ftqQhrkGZQaoy7Y48T31ywKf81tgUCvQz81nkNbq4YGZ8x31eN4/jp
4777iU5ziNAwDeal5nqCkx9jqnAklKhoGKsbcfmPSu6iMofiZ6f02b4643IGGDAX
APcdIBngPrmYBIsOTae5m4eS9rCeaWhLHluTAMg33TZ/iE9qdjThZxHpIBfwggHc
wNa5uFGBjePAerLehbclBW8q8N8P2s80JShu+LTwqQ+KNeEazd+zPEVKr2dXi00Z
ZeZUl+vTp9PI+LdAgSERz6aiXaQbCp517p1MgxRJAM+KQWS+GEAWdHQLdVho7XmF
S9ymI72sxHHqrk4GeJX3XNLFKkVxEmD8YiKmX1d9BHphKW1+t6aWEVUYyZXsKkVt
45txbD1Q/d0guflwm4udhz919QY4okdWEFeJnCDdPoPCr7p+6fgzu3VZbbS/lKoN
DLaCONA/UfuxuoomrDDlN/b7XFaTQ1+AiCmNMPmXAjHkma82GEF8Y5L1XM4T/BTh
uk5bbihSHfDxMFqMfO9/QmWLqVkqb0QhgFca+XWir+fcKCJ3alqQRumX6acQAW07
bRGzFI2i5xAHUPOav8HmENRLdBz9oBEuPwtwREcsBieFFtwgmkQtrznkTPtW/Y3M
VuUBP+D4c85YW6we920Js+Vvibzn3YLQ9m4VJi89yBgkjcT+DhyT42Zx/R/x+u6i
rkDDuDpzr7Jcn7J9vQwgcFkIiQg6KMgEX4B0K9nduFwfGSSj2jq0DpAQYB3kdX4t
y9ecbuMPlrIWKxutAU/G0hJIja/d90RQBMIQwYYbkxwgUSMZMn9te50fXfd1vond
233DWjwTcllKsQC7XLlGAR3zj/iH+2HFODiVrdQOrnWb/xIVQ+Q/0gxGnDQZgQr2
kIoQbtOZshg9r2dM/kzLz9d3rly4021ax900kjSxl938emRKN7kwDu6KtlxnkYBj
nymLME2fcxu9a6lTfULNn5KvA0+8ftt5kljnxInsE8QOb4hJ9Yu9Bfxq+wD61QHR
TTH1HSMWPd5e4r4irX6e989FwltqN5oyvmRyEkcLAS5ESPN5o9vp37H1eNs2H8oT
rsTgb9lUMeefKB/6G5d1nKxEGgHY81FzVllT/vMh1GQrqEpanBzUcCSocTSJZxoi
INLsNE/K5Ekbmeyo0Jf4AtOcxerkZmd5tE1niACuBPaZhTV6/0KjxD9K2dWgTc+m
V+ZfdB54cQ8P8kR/mqnAJWVF6x/CqcIjVa6TWhwUZNaetecurkd0VYVUiPx9VWp0
2yFKGmyen/H7VuE+1L7vIOcNYX9pxQ8xSDW+j9yaSBHhAK3AVUSgWqlny9FQ6TQO
CA+E8A9dFDXj3rtQd+sW8RybjVGtaTI8ocWEnD0FHevekDAy12Vs/Z4ceXLD3A05
evkkukfhkWXWFQLPPzndTmn/EZUoqdhkTGQCXxQ6rNHnBI3bUMbAnjImanU7aqgo
9h5hJuEDi/+fyEjEpqH+xdwTlRWXY/dVi/qvJUApKiziceZYPi8TbXsqO1Et44v4
fHoam6Hc2YNFXLkfcEL1O9n4qGH2G01C2z38odJmc5aqb3zuY35P9Lo2DMvzTmim
2UcVlDGB2vbgFUnRpv/K0/GlxSQJVCrr9dY5BrF9dTDnQGNqxJs/F9nmAEQopNZQ
+UuyvJHzbHiwguYxM5jlSa6aXaChR2z6CSUjj9aQhKxHW6jzYH6zGmej+6MUofdm
2CNhXx8ZegER9Larxpv+Ni6ZIojkCtcJBelg5EH8WR8dow8nVyFecw9DbwMMUmvR
kzRLVoxruQjCMtEozphUbd8El7Rwq6mn7dY4j3y2iDgbM6FtpUzuKeRG30cWgvK4
3RMVGYuupckQ2cH3utX7eNfOfGj4He7EKdSCi2XCsOoLcWiiOnI1N0PYyZ5+oqNK
FPa1AoChZR4VCTM6xZBj7viKD0UycTPUPMHx0qxXUX1I4t0iJqI7sgmG8IBsy/f0
6DzhCfef5FliYEBOKwqqQNJLLDksvqXWIEKIoaZgshYnp2ryTXul3RD5zgiyQSP7
w/cjsN5uxQaiogc00pmX/F6Ga5UFZYZUkaccLMCancnxpGs/9Ifa939fN00JGVVi
hVK/tIQPqO8S8P5225piJqTmFRyiUWo84kiMjPUDw9uSKN3Mje6SCHgsISLhl6ji
0ULpo9XGUNA/6ksjKCBO3WZJV2pRSmH62FvtqUhnzwsqrLpeWK3Nd2oy6MMo2cAz
+enKIDHYm/kH077XGIUxsBrwycf1FwzAt2DzqhdiIfoqhbuxmvUHcB9zAAUbodGz
RiI5QLpWlOLQFKY2IUbSbels68u2MIzHknRX4QKiI12AStmS4Ft5wyslqdPxaeOr
xZ6p9atjo0TNHMPkWPRu5qUnjqETmvHQYHejk52NdacT5U4UZgDsXnQlxgd28DMT
6/DzXexxxwwlbh1N4KoVdcSpaHx2OaFqSzgwZudpEhiFp0PS0kIgzeOLElPRCdhF
9FfenmNpmZ3MesjoBpvGJcXquh6T2g2l9z3uNal3QH6mTCYoLKcFFjrDnfGYkJx4
mWnu6o9Mw7XZ2tCirBMYk31m0hxGuzmh4oF5KeKlzLWCqgXI+atYSwEkbvJSPtQc
l3mcfkyb+P7gbee9723n4CufHll3ZzAY6IEnt32Nc6kE8zXKl7d+H0UurataYGre
NeSZPYS/QwPHA7No8tmwQJ2shyZkwJYjjDF4hA5/CegqO/1Wws9x6M1OmT7FEasl
RVBIWxZY4Y/mIp2M4SnyJVQ3BYDjJd9ecIabPC1YGSM/wyCGwAQ/UqwYprClVumE
Pd4asZsWAIlzgSTOXAA0fwR3rrGry4LDOTyAMHzoPNmi0QnWkYwMDFGCkYQH7Y+/
vKjJ8a8+BjQ1j1eg21MAjxuyAHiCA+W6/Czri3j4fk5Pn7XUrMkeoN/NGq5VAQ3z
FabiPxqqNoqGF67gWoDz3coqsCgAIJ2eAm/WHtbxM/wfwLlvnbYwb60lPUUvw9AR
4uGrSwtqS8T7gA8bUXxqKe/fOSV1tfgATuK0WPESshlNtpiH0k13mpqwFZaqejPr
8hpa7ympA1mSGdbtn6W5dKCahIsbiE794oKg3FsIxB51Yq0248zFK/XSm0/cBaQU
USEntEInHl4xxIbIjdGiKSqe9mUlfEn9bB4nCSotWLw9SU1gRS0TLJTs4eorUWE1
3ZLihGVnhmdd3UP156L5UJPsd8mltQ/BxCmectpYGRfCcDXm+wOMWWJU7WYbOH8r
KlJYt9i6bpbVep3qG0/GpiTtuTRzD0Lh+jZtt2wCTEZi/kAKILUxRAIYYH41ktg5
iQgdX3PH1DWFgcw1u50LdVxs7RXaZiFIuEuB4xBvlayX6Gwx2JNu92RHjXtd2HjX
ifzX44BhnaFmqJM19Svh70ZvflN9qQHxdO30xg7JWNWkWLq0LTTtGJISZcO/xBpJ
3pg7lCutvgBzFppP4HtG+lgMWoZV9Ff2KAYuU0Rn+M3A/sQ6F6PI+lqIZNnHBoEg
kNxuWVQ8Dy08Awfjip5msYi1O2iJzdJCXGQXMzACyFR93UcgNQKqKQmZmw5ZAZqc
CVZdZKRQT1iQ0uEssXAXIWnoTSnkPzP/xwX89dVgB9MlNzjLXH/B9nr1skALnqAn
lTO3UomXklHh53z28Z6FDShGSUvWZzJMtSMl1wJptIyJPAGgleJQrZHKNfG98B8Y
5bnw2bM7m4eyBugRC+5je8hP822M0+lfnlQ5D2j3QkEXKd1RCKZL//wA5jaBXJI2
xykdG6C6drLK5lrs+ZzkKsrR9Gs0nz1HABWQeyeFqXu5Sq7wNGyB1+rIOg4nOvnu
dSBAwWpBANS0cQCzoxq+R6qUKn2wo1a2Q2MYDKilzPA35KM+cstzKDktXAzQi2xZ
ZyUtoJbu8gBMifmZEjEUDlVJY06W5eRAQ5bFBek3zrYBRbKGgX0THU0rKjJOzxIB
jc0h3iQn/i4q4Or63iaFDoz+sezmraJAT0gFBTwkbnZRlGI/Qj3vw6xLWrtd7Mmx
pl1ICnT1Idxb7M6xIfe+jukGatOeE1TnwgVpOQI8c1NNEYfl/w1zCeuzEUOfVrfs
wD66fah5E9IPN9ZfIeTgCNyTIHFByv7Lzdg7u033uuqn+Gmfx01JN638Ptj6iz1h
ozK03RNptUuJAA/iIe+WAuFdqJKbGFYKouqYTVeF2fM17sTkxoi7WoKGsDCkXhBF
HXmLDLgWmj7scBVeoaYG+KY7YcUPYZIHVVZ34fx3N5NmUKcSZzu1KZoQacmKckaC
afTsBJ2PcDLmCZi+HlSPekzRB8P10SfHJDHt9EmecdgmlAwQZh7w7QLWeFJVBuWK
bvNBa8bCeNalZWyT+NV+lQYAn5Q2aeocB+vhKppjWs4yfAoHm61cRdCBDMskXL7F
wMPi5kk6xD9lBhkaWiy/Xa8nA5bK86Fte5eWg/l4d19Jo/RvwGmSeF6BywfHfyYu
MPcp0VXEIArF4tPa197PhWZFXotEyDSeFlmvq2qzmgp+iA6ky9s5JTyWLuk8rjY+
MrbHl6jNzIcjW9pm+96AK6hFj9muaXH9pZ6selvXiULTXZu6+KN2VhALv/SXmPmU
X0W24iq7bG/xdU5Tp9cjD/m3mXe70cSOcJhP/HTzA6DoMHGnn/ddLXfXsMJXd6ik
EjjAPOZ9AIaVxxMvdNxkrX8i7Bdl2sXyRaAErSXRaWzzRsi/7xoL2mho8+9iHEWp
ijk/1W02iqZGEsC8QFdx+aQ8U8z9IM3ro/CoOFeCXOzi5OkaqOVz03o9t8fk/tBi
iALnRgxDJ/7IV6xHHDzhqMC7lt1F/QfMKuazDFzfyb01kVAs6f+SMppnBMQ94QPt
eLHhR2fqYSrEh28T9HVHW3kzGMIDsPZH09dLHt9HOkkkWaW7U7VDhxxatLoDDTI7
gBm7I5/xynW3M8upGRcsNGI7hNwdw0QwD2u7bDMCr5hGOBh+5M/zeBrJhtnGZUiV
0B6o32fkRcMcwc4h7Yf79bhA938rU4AwRXHjDze0eBXUCcAIVwYeT8MH75eB4zP5
TmsY6qhk1UAcPQ4dg60OuXnJvAcvX9IqtnxWMaqCe/Rstx1rwO1BE4Z3Ql1GYVc9
4CbhlWIduHNcGr2BqDDVC+roh4doOgwV3okTRBc+VrTlyMyyocAjByp8c5r4mb+g
SFSJInJuJlzDMnCD84QrCp6sQPYSzDj8LXWZ36laC2wyhSkHxxtQ0MWe1jCxh1lt
0lBtsVt46YNB6Uwt6Md5a2r3EPl+CIfJtnB1FogjNG4TnciIsC8IfcnWatirUpK1
UWflAEwHwj2dyr0s4iZnPhAZ3cE0eGCkchAmUc7pXCflVmSWYfwh9aonn/iWqw8c
RAeFG2zXs+rbJ8zx8DpVMAY1seCx8Npj3qcJvToCYLn0r6Nim7HUAWcGYj4SPHN2
hKMl59lkOh4y85ahiSw1NAHT2Ow25DL9L46jdseI+hXQdMne+MWEM5d6v6w4Ry2V
SnVXSIOOdMBcgoduhNeKg0+d/4T1OBWVglF0r7cFbtKyi/NtmoNY/GdjzajuLD75
s7dajyVKG5XG0Zh4RKtJ957f04SZWv8rUcTqHQt5FyjTSp0hGaLhJr1ujaoQu09A
gnmhSoDbVBUjHxxdKM8YmTQ1ad05D6r2UVzpVPZr95GJPC0rm0PblCVU9E50FmHl
Es60TtKyfq4oCEquFQ9f1Ri/zi5Rh7Ob65SD7PiO9NwzUfvzXLgGFXuZRMG5Q4cl
tosUOfNyhIZEqx91BrOBzB8mcU5Ac3cQf3pqFX89f5Mq2Shh0qv8sBOPFE+NtDFI
Zf4jykU0i3FLzbDweNVDXtAnk2EbYc0IX9ZlBvcYsuUC76M41hWfuPd6o5oFKswa
KSo9GyFZyJ1xSU/QBm/HKpApMqFOxMDXfZZvLg1ogyDK6Pjed3ceCrJvXrmHX07f
anfNS/xgw8Gp9Aans0m3T7kr/bijf6xMo7GCTHPt/XeKi34WNs4zyTGILoglDfJ0
LyebotlWMcuLYU94HWmxDA5WhWiEQbEQCgkT4FRAH+yiAHvf5PgZaiw4JWc2aTHQ
9E95PZl1qA2Dny5/WkAQ+uqfLHZ3ya19knC1aHjXrfjmcNTlP5Sq2hIWlcTl49la
tvSa0CTgJcQ4UviDcQncHxXWfLA5sNVjtmwpic2GRgaqTHMMnYWbGElHMFsBj5og
bSUp1uBrNC1AxN0ZIQVea6yB9UXH04g/NdXmYL+i/jhx/Kuf2lSUkA1Amx3e067s
zY3Ey6byY5IHN7KKzSUkiPqgFGEUGGhx5wdjVHI5LHbBkDdsSJvSJl54P2KvYuXI
juhQKWwTXG8TC4kGLr957syZKlJ5dw6g73NgeenmpZGyMvyB28Q9x9lJY5iej8+Y
gZD11iuNlLSHEcVaQ877ug7eiBUODa1ng+BWMZ530BZTkQxisqfc7wK/2bdAnI49
X9mvGuJ1QUdl3O4TmKyyiqJW0lauZaA+EkDy3ebFP1tw165nJqc0aBFaX+Y4a5zW
qBgojnpizN7UxLI/8mDZao2kkiAp7xU8IFlduSuL+gIZF7zx4NBqHCOOmxY4H7ii
RIpecCOyLjgfL//KGBjW73CvmsUzFOCA09sb9Hxf4e85HxIOUUlXh3ybcv7H+RGa
I4I3GF/P/yuQAK9fO8t+zRtQLMBxFZlAkmg2HhFiBN03eS+Mr/t/u3fvn0zGw69x
7IRf5wxUh1SXdAPLneNNhYU1Xoj22Q0iQY+C6u7p+VJI0NExWiDTGSNmsZMhlL1W
xzRVWnXRZmvYxayyd5rJdw3jpEmIxHsYEmw1cYF3BLMK0h2w52nvlWbJg7uFpVRp
dNRXB5WcZHRbaatj/qMGbGiFsitZoD8RCUo6WuQjA2jj33M/0445KikNv93aQcuq
p1cBvoHrMjEswGDkRj0bNqwnRh3Iy/YDapNi9vx7Gazoe0fjnuEnxMymTDheAJ0z
WsklyfOzOHKvg6A0lTsFYAZ9Qhjd8p8SG/GLtjxi9UOzAqXAPuUkayD1+TRFHbSr
dN2rdQubweceNshBLFhSxQcgjMHwqO58b1gP9sDs5k4RrUPUu0Lea+6Rq2CteLLQ
W2U+0QyieYmu1zrwaWVm4CdLT12O6w4u41rFFFyGeJNQAnLUsivFLn43Krt4zMIi
RnMIaOUIxhYG0ZjynWbfC3wwPojS06tgBt3uZHWqCfItpQ/NrrXo7O9iOG6+wrxl
KMzr4hwVkhWTHUCrDS2gSCteZ2NHSrWuaHoPFzOvHVGiWTNqYvxgyuvHLThi8mls
X0YTHs1jWMIkEr0364vmEfwNizNsqLWPchRAGrCUMS3u83G672C986flzJmysVlA
z+yMGSO5PVr3nPJUPmYgvn9JGAjxADQnfUblmlpZ7UthNdrqT5D8/NpVP4YjDPku
IuZV8QdZymET8T3Aj+pn/fcIzR1ORw9mn7GfgNCnXTIcX7ZBnbCtNjrehBYSAUT9
0GK2Plaslh/nVSXgMtg0Rg6b7B68xhfAudttarKxyLBc1qzCLJZ56ORViimz/0be
N/XQ/wV3Lp7nLTXjzbZUMxCoxOAqFDwvoVOMibhqcE94m7MsLGEZB7VeZYBpOYhh
i7UWoIbjZmrm0ByzkmvK1+TnL57ebgvp0T1FaJWYvKgkNDzQj+AxeFM+lAbBFuXv
tWMhRXvbVzvjz66xWXMhKn33D6SPDzMVoNM4mmoguZTuqfWQhd1nDyKy3psjTzMo
WzUswI6+yei5rLlbRzJJRepsnmNu1Z/u1vUAd2eoEgWMIE/3++w7EzhMqlAEoJC5
c6VEGNYt74e5QF1ZotmyfGZOVIIOf/ZLZC4mGc7a/aKpLoWz51GvbgNeXLl7DEVT
vT/9xwVNonPG3WX7gj1TKCEkJTkEECYy9ftCcgPffUSLFpnnkmeg6lfjRDj9cWoB
7WtVMi47Awj+NjnChNwH03XiRFes3BW6EQ7FObkH/FlF/V8FZ0bgmZA0PgPOXjCc
YFrt2Riwh6jlH7sJhdhpKtD33yPUHoSv9g5FzfORSOr79mNjVjlVOFGZr9cBjAuU
ycEIP6joz5rWlky0MZbNYEFZaOOVVTnRQ8WpGKWDWQF4l8daiQDNfnU23bKJTdS1
jB4XHBJ/2MSYKaF2ylpnPV48tL8z4CboXtsLgioX06dadn7JP23oYvV78F8sEF81
NAEG7J1AJ/rt2LilBIqDAJyYTUHxtj0+b6jUdlJv0SASEVFb0gsspX5b5wZTlnyD
M3fRxYR6DPDxNudontBvRERJZIUu/RV1yFoVfkkUhpX95weHxu99SXt22MnHq1wU
Aat2kB0WG6MAVeMbhBtCnTu7v0nUJaYHc8rf8n7fGWkTp9XIVP09jZfadM1VCEAC
GSb1i146ti2vqZHSqLQOZbMzqUW1B73EbMMZewxXOCzITofO8kPv87w/tvcYjFDF
Q8vilL5xHLsrmmMXFrnsRor4p/9N3+xkPLgP9ehlsIDuR6fIaJu1jo0asd6KA2Dm
vV1ZgOx+avJkZF1yxweKMK3WI0XMfRnl/11zQdkBmFVxrIXjLfqdj26E+Z/L1JeL
BX8zEokRoRKxF+T4rYzVCjzsk+I/visfFSnC6HorhNeh3w4c8mJDSrvL2JTbM5Ms
UkRpgdi5n+GFSyX35bmV82UTTJZPenlrha4UEqgEnVUsrjSZUcwgdq1OOxNiuY7N
vpDcAJTsSA3XcD5fYjjEmHST2gePNWcw7YyOHSpBjgjqkFrOQPMkVZzzIwaSMpdD
vi9wSsB/6KahdIip4NkHeLnWPys+hRYCQRGTtVnvaCGFSFBHsIWhkFNL8Zu0gHnS
+nIgEHPf/N+Nywb47LH8JOXshwwiik/dM5t+fHQisV2QxPFHx6OxjQYak7HYSbhl
eQC6UJlxLy9Kw9ISWLvOF+Qf4ZOTMfrqABXt0qQaWuIp/uY1wSr7v+1cpW97drMM
XuXi5MSygpEAqHgL2ANLacZ3rIvdiEPVq+z1vDm/FPmQ01Led/xHcBYhPfMWzN+3
nfGTT4uNpyXRNqm6dKQxQP5rPEP1EOWH3dVgNXECp3D6YSUIUEXXBSdp3iXSW0WA
qTPffJgjRape/OqD+tM0NHGyx1hM/t6Nf1PvmY7Zl9gpIUY/1gyaz45Duy1OJVzr
H1x6jqdqQE/tyqdeikHrsgnpcf2vfBRhFmpnFE0PPF0s2/xLKW9EEJhgAvV5BhuV
s2eMmXWeXDpX02LOnfPl7RrL9T53GkTd8BkUgcbat6WgmWU13ils0KnOsKHJ4TOz
2QXdpxMV1ylEXQeF7Lzyo2psR55dkMjnDGbyFAvyLYTg1QtLtmkoWEiGcLDkA/yJ
zjfVEJe3rf7EtYWHANbckIFJitufr/O1Go/5Nxpox/fJRG8tb+3f4gAjTqKG3hny
gX5K557mzXwllv8lyd1XDw0Y6SpAP5t/3Z8YzZunnSzxgRioW5dVL+Kr3mzJlE7V
pj6PAwlGmdtvoXbcS7VXyYiDcmNAkCsI922S+gH1P4IlCqRzsf4OknDQ7P1SNYoQ
QP55IbuhYkC3HQsSnr2KRf/iXz4Cd3qk2u0ZpXA2NinIpLTBjLktBk7PTE2DawtF
eP9c/jFmG31DcleZiXX7uloKhmIquZOF2FjD7lUkJEI2PQGzXHSMN9NdAfVpJpHs
GC71isszW3pZHabYP07Ae4NtEJfEXUb3IBc82LuAE05r4gRGqcUGsqKL+p8fhl3u
E5iOeYv9N2MHFAco4C47p0hQ6QypXZkR8Nbujc8fEaPW5DN6DIil5BvOn/t15GPB
NRFuATLQJvJfapuP7FE91bRkKF3/0qkbqmPsDZfAWk8kqvLZv6KFAKgRV83eSwYj
//jIiMudgjxblnGbMFY3Bu1vmALbvnk078YgLBQEqv3w4nzQT95t8+rSMNLC55n/
VEwo60sgYmlN0+RC+PlhE9mRipnYfh4sjQha1LfcbAX84aVaOfUZOxqxECEVL4pT
cB4Cu7dV3LN7ngEPCYPRTao9RHc+qm8CP5oTF4UWx7K/UrpK19UHHFmDyVvM+kep
4nCbK8ulGwc7CgszsmUtQcdKTchf3bdX7irfy3G17t3mLDWKythPgRbe9COwr+qA
lvk+bXooaXlUXoAcKONmj5WC2rWTVmXoqGCvbZQCqKWTIr3fvkW4FUOk8BFLrpyL
f9cyaFjd/KI6T2Q3lHEyAQ1b0ySMDqQ86jsB4TNCkye4mLc7YNiYdA+bJ6xOFxKS
2Vx+RT7ymYacQh080BkeSB8GrlYQDoB5k0NJO451UXgPH9NHmHHchJkDIlpD3j+K
HI9wVTG6z6Nih+qLnQb4LRyyf7XrskQKzO33zZF+eV4hHX0SD70NbBRDjMNbUtsN
6ksX7XOdVH4UK1LoIEsnRJlJ8aZ8zI7nSY+nM/7IrRsiCJBQQupVPKWDzw+eB7M2
Lp04EDP+fiMiHlMQjmP0bSkqSWpH5oc4V53CftkGE2WhisXfETXI7oyuBTKcMzeA
K4QtDytP0PDEJi1N/HQoKXjr+v4rLPEFkJvws0YHLI76pgAUP6qo6flLi/qhoIQJ
NtTn7MBO+mwDHaqschStzN32OQrl8OvU/MDuKZDh8sKsuPPuq82Wx7k200e0zQyA
P+IjCxWT/BloEJXVzCMy9jYwNsTnyXo/Dk/JerNDh5CFiF4GFaEYQHYZTlDmglH+
yGnoP7PbJT0w50R/v9QkGOKTB1JwCfGeEWt6hOu1eORylpsZtwrTfT7zjjC9UeP/
FBuNnZkKWxJiRD/ZvBBoIweP3+FJXin1bgX0uG5y4kZtC5/JZCjNmo4DX/8KFz/c
c1P54Wl5zKFdJD3tDqTiBfGbHyNFELay18vVd6CwGbQHa2ol8z4DjoiEVKnNElzc
BwmNbOInJoIlLPND5Uipv2b9wmstTW5nDsMDJ+9cgI5C4fOov0wMxOtQquRqXFm6
12bNe5LStA+u2AdxiHSsD8uPQtfIK0JGxu5t17nK22qws78m8W5ziWRFHexu5+8s
FrePKHlkOG97MgiswzAxEsYC6v1kLLdZjKW41V22kEbKBkmrsYq2qRmm16NG819x
xwrC9U0rmsGNzyanx723GkZrs5znD7qX9O1mOIMZkfayafb9mW54Y3ZB5+SHlm2T
00/WdoGLAp+aX2FbicoX6IfE4reDGhLDE3QL88mZlvc7FnmKx+bfc/quLHplW/uk
AUENAxHcav+tDOjA+QcN4Y3CnNGtwv5PvZLie3fKHsFJ9TOyvzPr8XKVJFm1FUbV
YpPAryXV9bznB9XIHMPNmW9r1/WLQtEhYbKocPiQKrbDwi9ceqhQQuS6SKe/QqOl
1tICHYSLqLsXgCndgc1kdtlCG9zpVxrgQM3Q8E0ZqMG1icpeX42sUAifVg2ySaoU
zlZO6Sc89OPLgk/WnW97WKfRTeAaQDF+k/D9eJ/fA6fksKkjFPw/WjPEXUPgm4P1
YNeBxtyNm1QAX3WKfLxxfotZc8/hk4iBDe5GHcNw8In3PK5FMYe9/YOGNwNM91ac
OWfXijMK0pdsDikJdkv+8ww5N6/RZaO9FDvll8B8BrejffL2pCePnga7EPKjfmT5
ew2+Par+FcUc3qhcvUmhl9CELWGaodERikVWm2EppMn5OcOvS7kl6eoN24wcPEjm
DiCGJBYJblFggs5rkvYp/jWtODZgLXrGeKfeZMJK5u0wWg2bqUatyOY5DJ4JL7N8
SfyomU/BFGl0piVPOw+S2a8n+99EOA2koS6aQoD9sHM7amtjiQfp7Ad5SYH0wAEl
q2AjN/1iicdcYpKNpkkxNBgu6yPKXLUkQh5apRKCHaZ3czNYO6CLrlxnbwc8R8U3
r4ygSqj+GdFnBzkU+qGHpzWuYAskkIIE/JE+NAonbikHZVKB3Std7N0kykSqaK/t
QvMbi7Qa2KiJnpayIaDEc/L3BPHXBj9E3kGJLkg0c5JK8x0hX4cqNd6y3qZgTkMN
X44XYGlmajLQCTunXW6/2CCLY7CKI7fvTgWU2BF14QiCFZxgEmcKx/MAbplyfMQH
q9Y9lDkkz1ws45zCX2cGJNkvdp+HdhQ5u6hLPq+z4fMcs51LEnSDq3sJc0FMQXSS
GbuMW55W0DzQSTR4ZrP+smsELHTvie0UaEaexiiRuFUaTouDKq5OJ8GbFA8o5oSz
LDl7t6C+yu6fOmAKLBn+kmSDOAGvGSIqPKm1KSbYUeD5o1QxKN6IZg4oWHER+/LT
OXuw58LePLgtlR0ruLXMoqnP14rgoGOtB+jm1GZcmLcM5FzxkjoN8Wdbsv7bsJfp
lycOs0duxcvVznFDzPo4v2UNRLxo5I5u5WrTQEax8cgqzZeERuI4k2xLlzW2y8Jg
V0ZhsmHeojRQmwbtuzM4ug0cG01STBorIZXouYArOLzFIX4/IZZziIcSzGpyohaU
hmmpgBbtl7FmOrJfdkFkV4TiNBK1tF6X1w/1b6TkzSycbp6gykEMj52Uti69/HR1
phBmPDCAfBhVDw+BrdCh7mt66kwVmmZlISClZB48mdHiAlXYFtRjKxRBdzxBZThY
vFdIKMjpznUBcGd48rXVMKUaU4TSi0Y28Q53uBplJdCcwR72/1qV9+BMhft/Ux0z
uZzkqFLe4qcBSg+/too956FoiiYlZkfkx8kbeiRWlTmG+u6K53L1N1oIGFbR/POY
Vc1QFHYRQUQPonccj0WXOcYfC97kfuVBglpH4M3BzR4P5eqr6gAxOt/ygyyOArM1
puGyp+nntORvC++zEWirbb1hAwyzY8jp7/gdsfxxMReWAmrmzQxWXbh5Q/kTlL1k
m8HGB/gdqqHZF2n0Z8qa8iTQLZBQvw4DvtVMn7LzME25NZhz4IpLPHK6QXbM8cTz
g6V1LK3r3HSoeUx8aHIMf9Ol4LvM2mrDaLvTzknffziAuTCaEoZLXva9HF8J6EGl
PTIQEmMVHNYZFnGIjYg6HCvF78ShWUTH2gBpGR+EV8BMVYSu1C/wYQ4wid8WnThl
qu9bmVkX8MsPYryaaTiZXO2leuG7iyPHkmi9GkRNJ7ej7LNzCc6V/axOdI3xb7X7
qjOnSmXVJXQ5RQS5pI4g5QHfMRePSEb0sPdjSL+8ZV0/ybfrNwIpyEL8aytVCoM6
pgAP4FKnWhfXso1Qyq89TFZN6rbSBJqHs5pCOpcwbcSn97du4LMgJ8rFyzVvXEGs
wXf9g2w4YdCv4Vg0Y1Axah46Ohx8WIGmpHOP9Ux0xVJ6tccX+Kkx1tHDgBiSWFGA
Z8fs+B0lW569MY3pFEuMqkg2BAs2WLIF/Ip0Vcd9WMOm4ITmN3qxSIEI/4GDFhlX
QZhX/QT8pWRcpkRsVw0hUVHU8HYWBhtTUsd5rv1XfWHaeqIM6XiFuoDQf/clJP6J
Vfm6C0LkraSbYckNDYjpcaOpOPBz8/iJ6CIaH51INuIg6OrBk0JlxLa/w31biZnp
49IDiYuts+mFspM/HIW5wXW+0OwZuUrLV+IivG4MbpVww/ykpP+YinaKAqmLp5ll
EOtpOkdDzjzlIPBDtVbzEchk3+3xe8rEC3ThwOtk+dRdYPd2YXvIn+bTjcTl2yV/
HaaqG9Ci9MD1DkhxXRdWYXYv1+xjMlxt5LuatVHvfToIg+97y4+gVIZCDIevLdrX
hoWloK82uL/TFhD/kUMZ7SpuvqqUrp9/kLiPD4u9S4xCKFeQGBtovdw10/yhjR4u
UFkysvmL3zs/5kb6IPDJmD6+0TfbKWfhwwx9eRR5Nf9Lkdvbp26gaM+SEIzlpxYV
iZXETy7uqqX82p/RoVUoCoN4IkEexNboEbDCi+fIBwQ24ww5P7gqZP41kfuv5M4v
RR4QHFAegDWyut4AZuHvPzkGgfalyYPsybmeFngQ4zthB5P6d2UCZ7YT3O4glTx1
6o1Yj5NOyyj53+x2NDjrWSXh7mkfLMX8kLz1CaJ8yqeNHzNRMv7uhTGWnx3xM/Mi
SkiBNrhnJrFNskbL1/HS39sA39te9ZlYV1Pr0ckhlgQ35txyMMpw7g5jMu6bcG03
PCkFEuvYoLhfn94snlix9ddEtjALuztBLPpCnwZEW2jO4QsRN0saIzC8Qj6UvnAA
Fw/dIoij8Iw0iGyKbFh5cdD8DVKt/ZiR6hfYHLuPz5z0FgPsqGNI5SotNDOtWKkk
ZMZ7oDz+cY44uFb67tTZChlVLDD7P32Z/1rd4Gs34ve+IUKsy6VOiRwHHJOvmF+g
j9yQIrCc4C0zjfRZ9aLjIh67q2PssLwXU0nLNIUGLSrRKguAiVsTjMQOgzNZOiBx
uOfVuw7yHxJqrvsrbCmX85YzlX2+it3oV9JkY1WZH1WL06mwGXdsH0QD4euYBQVc
0Afkkq1SRlYcMrs7fpWrv6GIf1BKaJWlW3Q2VvgO2lJkCLoLNi+qnTEwKKTpVuCg
U2xS9SxGvJz8tfQ7KGbxzhgc2+wcRQh6ItfB1nWtWn18yTV6VMCqzhNeWhQmPpMA
oyDFpvPjHv9Hx14/epoRRS32sgp9I/JZukXpgqlNNOZ6XnuQS74G2CSubymYWshH
1eiJKLquKmkxuXk9BbFFMVq97Q7OZzZzQvBXyuGh7kWB3Gj0vz+s0FtaPZQWDfXr
pc6EVEFUOJYWydx7hSb7KLHmz7KK/OKyMUKdo2rpECXaxPqjdcyeZOJ7OjGiszlp
uhWRk4vuFd/eRW/mc+4BrQWXfwV00vBvQvH2qJeW7bWzNCoUeK6wWgo6GeEIz63A
NqwePIRCWYmp2h2w9SvTPzunPyDkXcOWVE5u3Ol9SwkyFkjNZzSRCCGdLBL6TyYE
sGWCGtrH0Akok6BpCUzXa911mGVmZZD/PSO2v9MwXmb8siEbGKLxcD1/6HV/x7+R
00xZnC7tbKWeJ3hWDmecbJnWmorKeOYNnZJ4dtiqNy9ptEcFKxvRM6V6+Cwp/Ol5
NurdyXEdU78sv155a+GDF30Ee0H8VpLSX+yJmmvNXUZY8AM71QFVS18Kfo6ol9pW
24M574ZsZ+vKubnxui9xtJagGmFqtrShmujJ7glTaojYzO5bft4B06mB0lDroYKw
53YQs9NeTeYGbRPpRdzo/TL0TAgNa5sEvVL3/ZzKP7pTkyKFkGU6zHy+v0pHrmBy
v1a+dPYb/MztoQ4zZpnB1H6v4Su2HWfUcvuT4zgi/iji3gFe6oI8NK7ltsJnCVLV
qvgn37vj2PYaNLqRknOFsO8byF0Y+pDFk1w+wD8wN0FRQ01ZYJGmvLJrwucKnHGu
zaqZPhglYLn3Hu1zD7qnq58y3OxD/PtNYJgsNP5/bz+Ud/WA7otV06W1Jxfw08BS
D0dnMFz2upStWQR79EWuHruVHPO3sv6Qkf9Mj27d8shh4qTUYwosA4Mu7DkA9S73
xQiTaFA43q9NL8gC5ITOzUzlktirteSxBoWypdrZZfC3QRr7TYRKthtKEDge7rol
Xlyb3kEx4pc2PCe/LmHWPP1t3ebIUwxKCTPmhBVPKjKtLj3C4w0prEkQLS2BHi2g
cvT2YKEBCC+HeelQ6pzIZK2BlCpKSP7H0RVcjuq4IXk4SbUDb+NsLS6pm7uqh4lE
/DYGijYSaQB1hi3Gy5hWk01j4t0fOrSbJHFZVQLKl7LnhHAy/TEQhs2OQkv6dgfj
3grOQP7ZjbdDUP7cEfuC4BN2YbT3INDiS8coKU/znAKV2Lw1UPW/bt0HfwUyAhWd
Zohl2aoRe9PAiBxafwobqCkYDMbFHOJUJeZANKZZeU2cBUt0bbhyWG45czFnX8zb
KEIFioUzwJ4qg1YYkGmR/91wz3lYNIzQ+t2Z9YYjFfvYcVMf3ACuPHPggBLIwHK5
EkBOGv2umoLRv8yc0qlSFGByxv5A0U1o+EtxbeesiGgxeezwnRmsqm6cm9cNk6bG
MCeMe36h6xLkVRQUO2m+c43v+uwuSU76wzrpeu8oW+/j91U5ufPw6wGCbHRhW4I7
xXUyE7kynN0vSQmYE6gfgwNVDrTNr9omYw4YJ0GZ4fcV1Tm3fLm9ttEvGdASrldI
+CsprK01hWvATq4dbJxjB7P0hVS7BXflyB/8kP872lwsNyYwJWPNMZwOwHDMRM6E
JK2St3XKicAZZwpoZwbj+I3TK33/SEoMiy2D7ctZdGUhHtVaKc9zTF+9XuS/t3aM
FL/izJUY2GxLIs5arcOS4zW3PENY04rHcW/albiOH5CWwEs+nsxt6/8jCDXBK7hS
GDytj1sIDu3DLTH20Kv9pjyEQ2mjK94LWcUvdoQh/ZCl6s+UPi2wio53odf6JGYo
78PyHAr2COa06AusUmdGOqjBFHGMkUDpY2DdpKQmSXWHtVtI346VWuhA/kn93uz2
0dNt0jrRji6icE9g0uDh+Lm1qeyKvXJiTpMY+XNJTHM2mYoT4rKifE9OmozVcdB2
+pM6Dn2CFXx/sepXkgVLOizfQkmTJ+vghjfIRqopL63JJtuaI/nC5o3JeUTGkTkj
JjQCPaEwsUA8jjJQo9okvqFWIdkgdBmPOaGF1x1lcSp4phkj35C5vRoAVw6hvvuN
Z12fP5D5qP7lRbJJrr1SSfB1X4BJmaL4eOirO0jfFW+53XeDobgTUDH93ecXc0pg
sA0LCkxY096xJC9KD3D0qn5z+0U4XYfW6OHijAO3vEj0RJqjePqqnOQolf1gU2TD
SOCOxWuoUGrypTtGWPxmIh1AseYo+ON+Ta9ZREMrQiDXT17GAamjQlnddtyn++Rv
BUx5dWg9uZclLIr1qm6kxqQ7cNTV6f/VV1Og6GHCVdr9sB2sR0eBDE9Qoe+O6LXq
9CogjjMtGkbNMLOqtj3mZ4QLswUrYPLqY/teGeZ02wtOuHUHINfUmpOottdM9WPg
uKUHIHUmBH7diFGnmRfRE71XuzBG0WSiKhIosKj1w8qoPFV2g4xTF1s1whvDYby+
X280XNdvuXIr/QepHTU4LOCaDUWXvotTLvPzX5Pyd6P1TvDYTd51dmoZ977s5j17
NBjsd6BZo4wpvWjav7E8YJlCAHnt0Qm2ZGGloHBD7fQt3J4P/BaEtuPKRslTVmsu
c+vbNj/88jUZ5xD0IkHkXdDFjY5yY6EFqrIq6/iu5AIGdmaNo3FduPrsQczoTdI/
noexolK5Puf6BA7ZlmzsutHMXMnEMD4VzEshdUohpfH8u7R37lBZpjDFqbSitVEE
m6a8+hE0KS1hHcOhKLKJDeyADpcSjBqH69Yjp3Jod+mpxjsICMLSV0gaPqWqM3pE
eVMRzx3rdz29AWE4dLBNHiGML8BQZvf5ay0INx1VQmNGgZLtKjNwyLA1GRPs3RL9
MH+s7TasyNEmnJCORsfPX3ntCfHRYu+GsLOIOOH5J7TidOzxDRQ+Kx6UZ5bPUh7Y
MBleNjxYz7ZKV/V/qWVf8sb1oj8EAtjKeBRFJ+6PA2kN1x9JWZ+FudvqhM/TpEki
LKR1WDrM4Xz8sdHn7Nt1DFRusGYudfp+3WXlcVdSPowaG19hbemaGGXirv7D4ZI4
X8LkmQtZG9fNyGXaQpC5T29LCckSF2D6haxoWOuZqtBFE+Uncfo0/uGVJu3/k5jg
cMYzXPAttL1ab6ZfA43YjhXu/YNb5PKdTbmrEgM3BJsReqZQFv6bF10HHuGVpTx4
oS97/pp00CDiG5RHNB5wUfSUn8+yowh3w5nFNI7ChdynK9qVkpP5W7rmYU4IVSXa
+Y1iUIE2VJOC3yearMGWHT2gacIxl4UZYdihFW4jOaWKpURmYqzNu9ZY7pEABQnF
gDZk60v+BN8lprPNbKCLIp1SWMZjqKXLK6AVNgyLH/lTd5pswzOHoQO/+3I+Fmh4
53X/eguU+Qmbn1btLZSIViQ29Mw6LILXUnfY+S/e/F93LQLG9DoDy+omPtKQasg1
CkGzL5GQn067GKCQ4pUvEMjk9uv7ScLKgtfEkCslV6Qqqtb67DwmvGbGbWisM2LD
7eUlk8XH6YQyWjjp811UoIpgDYXvFp+MdcQYtsoBD8EcQNFasOJLPNhYOWbr+Hv6
2CT6LH4BuRav1Ok2hK7WDhpABtgXwtvmyhaLkg5YHJ5CtzrjV5WfJ8enhYCm/1y9
ts8uoHkd3Q67055wIJJX+wWW8Ezyf4JF5slGStiQV3LN5AWcn0xiCbYNv1FnfoLt
KVjPViGXSjl+eR184T2iO5hoLLcI10x1sHJzJoRlugnqX2IJEnc/rO8zs2a4QcOk
TkEUkr6uwjTaRe1897Ksp18zJZt5phrVY9bA/vpgkLROXa3r9dUUJC4IjMndUCim
/KapslYzjTDswQM0td2q4PThrPyWXo8BdBvohy5N7+FgLqjrBQLfkLv8jRI4ClMw
HxAwOBqjeXezlzhdHb7lsXsvVn8i22UrxGwvblrzk4pQJz6Rv53v3843q2rMMFAP
6hly+uB0dhzkw9P09yHWN7ZGaoKWgAVhL8GGNkOhgzdiVA3Zd/8ENSuBxKaAs63L
apQZy56Ewzjas2yU52qY45wq2xTFNUMs5Ju3nZ262+nszjBfQVTXMbKQ5zkd6ADY
OeamWQKj0tDzPIrsW2ggZiOepaP9VmCQqaIfJd8IV5WtRr62baeRBHqpPTba6jys
8mlencckBkfVVgQL7ZODIVbhhiWs6OgLYIaV3IzvsGUsW/3AbB7d5u89+YhUj4Hw
9ZYSzEuEvUjvUGtu6f8hQSahrY2C0Htr3ln5IMg0xCrBhyugD7tpFwqib1YnF3Rj
fCpNCEx9Ba203jp5JgxPay0k6vAFSCUfMRWbPUxKkXN4JqTzn2VS83HhMYkjZn2F
S9IithPDENYgqubvAayL6xiv0YdBMGjDQHmDDhOdem4jQAEFlot1CxgT8wIoq/V7
WlXbfOUWqX7erSpJ6uZ4XSKM6cun34vSLW2Q+GwB9RD1EE9d3Dx+//WgLbaSI7DH
7ldQ8N2WExgwm2vL4BIV+IkdwNOlIStM+GJlfTYDq/pkd6d3GIRoYYrPuE+VMuWO
aurxx7ZGenaFoR+VouiBPAapGXVC5NQC9KiASLpl64XI6r/DskBsQ8tIsH9NezGV
WsPjWnsU6AJAHbOBdzRFldd0CIv2mZdKtr+Sba24qq8p8Twj8SY4zw1Dbd2gspFH
AlTobshoXiUMU70zl1FYznseA6slKaJYIeO4jclORo4ndGo3sMJQ7r31aHg5hpOK
yhy0ytrN/ReKQZSrRp01YN1DNWkKSaH6lxN0HC4v9bGOppYFldCJGHPS+wskb0hP
/uRbmXsjDQ/enq8+01mg4Yp0rhV/ACzT3a7r2rTTq+SnzXuHu+44l388ECYr4lf6
HOXPLYchgx0aapqmjURb8M4U2YRkmFTTWWUeGC7f6BQ436s1CS38KAcQDnpRGwYl
luAFJZmEnvI0yDXV2JPIRpfg8vrg7w4SXwLTzkTfs24p3mH8ThXy/ajY9FIYcroS
19e4PyRw6Wf4dTAhOZuqzHhWa1DqcfR1f4WcMq61L4UO5bS38ydGd0LoELvPb/72
6Kbhtqz/C/GqR8/QawsDjzYZdI5FJsTc7Q+2j50eZ7Ea88ndkulKSh1tAo0gf7nJ
ShWymmmcVzz3kwa+JCUxktbU6Yt+cOq8BKU+dmIC+pDZtnB0IKxdo0TZONu4YH9W
ToEmR75pgKevzGhhf83DI80uT2QJMk6p6ZFUqbr0cQAqCDtfBOIT2c6ZXxl3Z0iY
X9eXhqUYtL5xQXRsgqmzBO1X7d0v123QBdvw6/c/G8Y0bQ4w3nZNhg5lVhbArwtm
+cEk+qRAObipP/bJSnA6CquAchwEt6pB2wBKY4goaki61D01vCLNGADzV6JqvRp+
+ufKTJQiaupX95k5Wri08D1MS8XqtG4jO13soc+MvNn/4S9A8u+njEroJjFWqbBV
sR/ZmkCH+ykyz2cx6sWh5gifHN9blslJtISnZuJNrDwgT5RHg2iiSrvSNOHJRll6
mGCsl/prKkmzl/Q+rXnSbh6SNsReco/UvZt2stqGHn+ElVJD4XD/CzCVLlBidfkr
yDjTBZb7p1vEjNTYI0pj1kTXD+jEEvD/+UdBRk+LbxCY45DIE7L/ayPyFbpoEh8e
Uu/dtvcZqwh66TJtjgBC2sOFTuBOIqwuuki6D371/7yaVxLwlVqfjec9U6Mstb/w
k5HPuaImONsnyhba87CIdFroHFLsoCjSw7ZDBq3ofiRYZ7/0RG2STLqIITL+0H89
EDt9WglaqNIxJaHNueUMqIuw+0X77bscDDD8YVean/pRiRytI1ryH3oO+QKcAyTc
NK8+ts/62RsaBkJfrV46K3nIybanp4Qg1QQwFrdC6rjaFggLnWBiTaQC3i8EKq95
Wu0ijSU/9x4Lwtty7Bnqx8LZTrqZ9PImfS+QP06dKLBhRSVSy9iFKtNu/mgsqmJJ
ueV4kHHMsCpcL0JGDkm0XTBowbqIR48jBlf9HoNG3p9PYe7KVQTMGfxgn3B5TaFc
ND83khmKvP8s0n8YFamPO5tU3u4TG3e80fHXpcHenarrN6oZpWZ/4OS4PDORK7e4
ePvhX5yHYfgIfzdaa8txaISu7G/aTMQITp9kV9Ra7wD/0Zp5ZagFdauCI/LB9zUk
FZAFs/dQ2AVu/9GAZC8not+RGeOFxsJO3pDWLcimSmCtpMfaW6HmqX8+Lgm1Z6Y0
7nKC96Kvsv/V4YRGu1FdgTl2Jf3/zcLJD57Pv7i1R8Hf5x/Rf9CPkmVCNLgUYF/8
i6cBdomnaLf6Gk0lg54ZtMd5V59o1EgJ7MrgY594G4ngHmbAdeKsJUGglildTgmk
WuGwf/cZJZgRLLr7jf7eWCHFjyDXLz01giuj7khc30yzOuFWts1H9UaMI9TKu8K4
K5gA8z/tMl7zRxWON+jxHbLQBDygXBPExA5GqE3M0EIK4IHNOVQNsdsT25Ar4a+B
KfxHSahnX70aPkMmF0XQITbk2IOzdbTkhzxFIaGgtfKmjHfa4DHbjKA22Chq4rFW
dY/JojiaSOVzwAfDY6c1mKxVbfpQWE+qUC8j+DgaxknWC4ZeY/rmSV/MxRwGXsVs
bR+YUxYi3Wd26sRvjuWIobdT595gjVntmZk9cZe5MDDWgc9PPpdWTs76NOFP5VJo
y4V2EeLGyWCqcyVjqTbGPsQ6XXwgXwNUnwWuGuR3o5nSSlOvPGFZWtVYPNRWNirb
LVbA+z8DGqXEdV1qYcS9RlgIYjalij4hcIewGdVtr/TBCWjnUyQg7E7nVwXYvEvb
P6nQOsf/Gc9shGHfkiWVA97A6y1Eo/zjoSXNk0/rrzUIVlUz0VhIvrocFgjh2e1O
wx5b42LUTbNK1J08MhR55YTSDkl3a17WSHLHDSfQGfaxWxemriQ42UwbXiljLn5I
gtf50woX8vVDC/LLRB80gkl3FmrabnHe3q4jgig3FzJYmi3pSjJaI79UWVgUBqqr
8rZ6ZpmArY7E+XcYttmRuPiW1IkWK2aNThAzw73uR7n/GO0jTpI68cSDSI7KE1k+
5G/jqP2uSt+CzQ5giugeWx1OkoLwCNqaAk2w5bkogvpEd2NI1Fu54KAaS2V8c6mD
nZBLreSvQ5eFpGcs8k+mzS7FZnSckVPp6qnxZibXcTqYApjaklEQM2/y99nSDwmk
39a3rRJ4W2TT7Pm1Teur92LHnSsxXDZoDHccd619xyIC2yxY5HT5FuILFIQ48iq3
a4payaPVQKnqmrmFzTmUa+R9A1USXE8siCRCzgc78WTne0aPN3fm88SJObfyA6cu
eaQ02LQJ4FsV0shpBJO+Ff1Fy7Uvqm3NnPZt9LLfFMlm+9yv2SyVFHDlkbf62cSJ
f1gga3Hoc3O8sBEG8H8MfbunWsJtOsBQ3xqX3QgE3BaPd4RIdIu5UsshR6vSVefl
2jRthtNCS7qBeL/7bAHwi5R60KDonvDKXBTssa7drKw442sWaMmNM239tFI9113o
pzVXhJvVsMCqnoROCBMIvfhPndkfGLYYPQsPShyp5wMJ7sWzuN7fGfiFYni76wEn
zoK0LLJFTz5jCpZ4hge5GYKXKXHnK1+o3oQlP168FmxNgRFwOSVUK4AZcwSMx7zP
F0Ts8aP8Chhmwz6DZ77eRxcxgUxXpREKaM+Q+9FrHj2pKDXY2lIDUc6RAoXkwWxy
k6KZ1/CfI7++vtZr81J/z2H4Ex4cETbArSXtWzVYOwZE1ip5ieVQFgFPwRSc5gDB
4rkZyBG3uJbxvuxaY47PEuyGDhgGB/xyESpF+yP3S2xAdIGODfJW6+75/XMtp+Dp
2sBfxYCd46ck4tZWJnXGkZRxuHfPkhbnDFoMFdA850Ext6AecQoGac4K66I036sm
kvDTMEuRzpNCH89PUFbsbhrr/5f8yP6fAljWdHoH0zncpjxGwdsHg7YTfDF9aq7P
aqhwBGB1u0odxiRWSelZ9kAG4AukePCshTniHIZ1bEey0AlaHn6gzi5BjQp5ZOUk
C30okP0hfId33Xb/tqYvq/NRVR17JJEaNRtoZZCTEJX6q3GQjHanSCQ64DUK/fK2
FbJ90VNOn6r0Zdmrd7LfxudqnJ/AyyvZZZ1C+XGasTAxwRCNPAnwUW2eP30Zrlzq
y6ouxskSdzGmN6OHf0ZTgEIs+bBwusm20JTUqOyEEDC+AAec3m8tN00Fxr72ACLH
oimjW2Njl4FGZ/gecNaq1TFuTA2SbCAINrW0oUXotRgqGmo0qMGaNFWewGJfM7PS
1nfzC0L0RHsHNgKGRYITv+1u5EOEMU1PFMBQOApSW3pzU+K2TjWdt/v9vleJgA9k
9XRXbghdOUQJo2VSECyyhWSJBMiMfynwbQWLoHorHEjPbS3sKG0Ikpac6+VzC+ev
Y5jYQPcEB2SK/TdqEnoH3ex1r3kLKJoDaqaqNKz3PQnoQIHh8ktTnBCWBALy9Ajr
sLuO27tVaoPVnghEI9Vm93qGRUravIAbp+O0Q9VyRUMeUXwT/P8q9uRux0LfG6k0
psvwLYZQpAp5wKWXTsZY8gXcUnqBllPVzNqLwERK/caetbUXpFav7gcZhz2pcZ8B
RTW2OTrQlLNHJB/yIQ6cpmNDa1ubnsmz3v/h4WVBNqAZPYSpuNo5QApAhbdjrfWv
3imF5PgpmvkliTP3VEuNoN6iUXi05aJAjJx0sK1gZV3bQUTIOYsYnAsSqknBbla5
0/4X6R3DiTn5k2aHVk9YnTcca7tbkDgYgxEjtuOlMkGn3k9F+TjpMUcTpNcNZEmF
Kg1LRlHpYK3TmIUqlfOAGhIZnX+pB68MYahHAv3s0XpDcjz5KW05CEV6783bORRH
MhJwe1VSBHTbV/JZIknMMO3ck5iOoQvNXLfKCCN+5IQQ2+29pPqLTCnSEL6V9f8V
ucT3VgN0NXyhSCCWAwx5h0URuWNKsrD5Kpsgjnpqr0wTCXB7Lfn5fJ60l0KYadRq
OonYhsPaZmQL4x2QVxM36IyqS5WBrN68cSWaqtmxUFPQ1DH3lDG6uC6cqJgmmOX8
0JIoQTzKnu/e3ImLigNyN/Gl2rvL9F7+oPPDOh3waxnASDAiC6SwMu/EiUj+3X8a
v4QCyDceect6p9Drhn5YaOETL0noXT2fyx35yCCYq+ZIKACZ6vRvKk/qQHj49b5T
01AiNpSkK8C73Rln5x7j4piS0IYSFnD1df9rpxmTihcWEkwHSnwfOMKSzHehoq9+
axG5Vt99BMgrjKe7qIVJUBuJL/DYD4DvKM/d049OcugmPLxxnEzZlCVhVJiLknET
oRp7QBBl4jTZ4+/kv3Ysu+r4hL3h2toITHT77fd9dpoh9kSPRZTbLCozRH4MUuSz
Tv5Q3Zqfe6YUEJb9LJGUx1iTE322mi/J1izzeulQuuo5GZJBJCyeNA2aGufyle7n
WVfB1zKXWDX8DTJmevp2gitYjDFfsafmUWraCfertQbf+AhxcfHfztgWkTRl6ZIA
SsjnNJZ6ZVlQkhgh6E/hTyx1WdGo436ymyqkw35264PvG5OyvU+cvOeptKJ4hpNm
Q8UXXFXUM30UiiCtOFm4La5BSBGhtXqvnZ+58JSYOaoKAn98lG/1cYdNj4mUbkEX
xyDxGQzTZdeP79lH3qU/gd80P8BCVjdVz563FleMIHaCl5lOV/rELDHIYGQOkMFC
kd58eQb874UEmICp6oownI3kIMxIex8GJk/qI3y0lUW9dsRlO2kATFrhk7rGBqsr
mj6uTosAUR/+jt+j9/wiPUanIs0LiWJ6oGsneOhBruE0LJ3UtIVyn9oKg6cq3B4C
bWYJ0PneR/y/9ZElHnWmeW5QkhaJb2hYxSd7MStwXzIHaHlONg/sl/9jl4CqcXI5
MwS8THmDR9gyxoZzFWYkAMVwg/zuQzToent/THP1icZPlwefXzE/7Jvhd1GEvpK2
kMTygSYIm/OeXqmcCdcWgnYAwHw0EPhKk6WKx5HUflIz/Cj9Dd6quyOKYyhRaQpp
6iKqvlSO7+yUJqjToGMKoYQq/yuywEi0JkT6xW7ZpCfkGc4x5rRH94z8it8ysraW
8h955Ct10KEvqM7/UPJkCRDNiRUvBdFbE7iKSBl2WyKp+lrrlN4i1v/XV+imqyUw
5GBGt7bw1xX1XBKGQbZBeKUB0LGr/3A3fWu/S/sWWm1lXq1CPN4o0IDPgpawUM4z
sRLUx6m1GIT2CMvrVGyHb2reF7mu8oAbtBY8mkJJOC2Nv7ovS3pjI24jrHp8Ch+H
hXHets9G9tMYRdgc9hkbHGiLfhATshYafs0skgQtQqwX0luRCTH5cEUCISFYdT57
JRViWiVRLUvkNmxCz1ulzaaXwiYAtLKVYy+PBPQO0d/rpmmmc0T7QN0YHwon9tA3
ooBpYzVpuwpM55Hr1P4vzPg9rL7MepAzjWNidj7RcNblt9Cn1Ecfjwfcu24epp6u
cdT4vmwhK9TMJjTzR1F3+bl+7TxmKavwk9keLTASa8UbAk8AooO/1fwGM3QlpT77
ySj/FC4TFFOlZ6NY7wtmZqDBGn8m+aiuk5TpwYKAn7Ez0UARy1ZaCSH5OQAPJ8lg
ziCF1EEtH+IaljXyw4yTUvltkFKql5+KsbChwI2LqY1BKhDXr4bmuMFZkU7NZQfq
Z7Z7hxCduGAijCVawRLswut0VdhOJnuoHc/ZsOh+Kftv9lGYdldp+SEgpUS/erpS
XSZMXh5oN4Jj+s5VSd4obFWbxF727DQelZo5NXqycFAP5Emobc16HqucEkU12zbW
aqeEYPmWShHtzIR/cj53C+DFNMmn4E3xTdtbk1Fr3aBYznnVd5uYlFZAgRKpNdF7
5BiNtCMKsG//SaeXDMxhB2jNeRlky2VcPp/jJt7WOfRAcUR7X9/ydiA7Kmrd8eiu
o8e3WGBk/EHEc6GO3yF27W1HaR7Id/Bl8lZulkSjfTU7MrgBsLFygslTMC57pWHe
9SMqO6biwXpMBZtgFgZEpg8kk1c3DfQL4BZICOvWQZ7lUV42876+h9v+5neeQwPo
l6StAVu5o/vriyFVMT3qh1OH6SRvKL395SzftLLeOrmT9UKl0tGumLFCEmDbFEAF
ixDhVve9mE69hYhBNcdyTiUQb80kABnjzdSxyu9TKezmB2weOzJd6jKnF5E44ZaN
DNF4xzOm54qGOUTgWAd2syDDzDelQBhgIdEgTi8K7EUymbGHgBMXbiVKo5dGYVaK
Dy3anGVrvhA7g7b9arLR4LCjWtPQDNeXrqlH8F1nCLpj+ATcA9T71JUhzCr04pvU
d/duAQKawjPDCgSUZOHSGVfl8loG6LcV2zRQQCQFejxxRm9HRJKQ2HK6xgtp4lnn
NC9Os0SayPhzkcgETNwuTBuyUTpyUQu4LyL/1BRfgWOq45k7pEFxpIQ2gJ0ibGTb
ZAeyUg7eynpKy4NIgXKx6jFxXh6prCkIf7foYExrzsfpDeBV1+CJAfbJpVhT9A+t
thX8PAuOC3+Foz+2C0ErpkfEQvH7BsrVJecZcONPV6vqUHTDV/+i55y5LQF7nCzT
UrgFgR3/X18AmG6MzJy9dP5EGjEWt7H+pSK+5CO6AQjWnnxARYVVViTMnntKpPVJ
NLxLiLSee7eORZ5B5Q7LLSH5vEN86gYjxRoR7exbwzdtThnIE0QnV0p9avKv3RY/
NlSBkIiKdW1EfxCj8z5F0y2pBtsJMnWfLKjZxToOaB0L5mZcxcIsq1wZRd8KQPWa
UMX1jSPeWRD4Cyr6gU0MW6id8Y3xRZ3DnAxRN1MvgSFYrDpPgTWrvTQuwVeUtGIa
SSclSdVIsVElVmDQ0ILC9zcH+JBfuRS4NJrKcn9D4rz1FQ5W5yzh6p8tP0/s5f8J
3yqGqNuRGYNHt/bPf4y2w5fYYKImJqZqTA8IdE8nebt4eAgYopqgQ+5KEWkjyzOu
qG7qUOKeAWHHK/iTv1Cd9u058555vYIJSBK80k4NzcBzNQPiDgt/IghKyFtNDPgp
q5CTblEyHNkxDletJ3uY9bW/+iMREY3p0lZWFUJp/vu5GeUGLMaalDRJbVMSODbD
E6SQiI+AlbSDDOWjz84EXqbuGTwRdo82Q7imQP+CGR14U98LsVNW/+SMEB501GSi
UfREar2qQM4qL5PVpd5XzgMMJGOC9nuZhb4g+rXaOAZlM8UZwBBa3yT+4tDrF3lU
L8Kxr+yUnqdMppoGc0fBFFZxspXw8YHdu/lCfEbHTYhrZq6LkWPVHiLoKiOjWSH/
Y6tzc8uITgPBZwtHh+GDPYweSb9RSOvJQG1WI8wz6UfcEo4RQhdqi2NPwBiYDcA0
VUbl7FwZCG6Gjd2lFUVn1Z2wYtJY0bcSOrDeLrzMIf0r0HaKqof/vy2FuX2o40Hf
4NcFedwCIrdd+EWRgyH84u5UC4UwwOAWR0dG5JPKAZi4Wignr56NwRoq/6+8DxgM
waMmXBorxaFLZzp19um1Rt+TJwsrTRfGnPUxdUHyUxQ3Xxt8ZF54JA+eUJLOhCn5
t+wMKI0wNtUSY/Jdu7DzM7dh7p16fATrU2cfnBKewapR+EymnWa5eWsJyAuYDTXt
jDsnDHkw3FxmuwaewmwXDkz8s+s4uUKEZ+yQmFo3DBhvIasTqEkHmEU1IXtJStmM
8pbbVITMC1K5IuJK7qcO1KelAfWKQIwj8PyADUpqhraq7gfnuEwJz1WU+KUo16P3
eFS2OQJx/4wZrppz9cyYDLyLcew1OtWgIFuEcjXYeDz3r8gqTUAb026Xo6Ff5eb4
Vxv/nrrx9jRu1D6cAV/a4ZgDAQtlJv/Pli20mjztRz40qi8fRTkq2Buiy34ejs2Q
TdkNNNcPoL71eNC6HOeG5YKMw6LPxt6HNHnYiNmYM5p9TIWuLUoh8QRZIhHp+dEh
laVMdPeJ0tM4ni4tUafRjOvI3TKO5SOuEgIKMpex06+2JkYev6oUN2n3iQT0a8g6
rCYxT8pkN7XBsuTkDkg/q/C6jXWmzXp7j5BhHTWLyGJNDOGuwyqR32nxA9ad0h0y
6Nre0Arev2q7+UfVjE8P9cQpqENUexfJjMKCuTyMFajbj+td2L8cKE0cSJqSUPu9
l9Z3YmnA6nbFByo98cs4hFR4Sb0j2m9Q0TSfxPLTru/HGgPC/UG85R+m/aaM6y/8
+egFv7/gk9M3dHYKD/6X3orgOOmp3wGOZyZ4fSLOXjB4c0k5hyXtdaP20P9zWQK5
0QJA+49NSdAAevDveXBIDJM6SKo+o/EF6TE/gSjKG9X9QF+15dV641NuN0T3Indq
VHyz49DcnrTkwgLSzrzmqI7uOG7X9d+pzsOBNhdLYlZ7YyrfRerDNUp7CjEXnAK0
43gxeyIhOUVRsikZPR1fSdu9EECW1IEqxL1qhFKa6rMGpZkoQdr0KVhVeJb+iyhG
icuGmrNKKwAUASoVhS5tgoKjU2NpAJaYtV0no2o/uoTh+0hGk54UtpC9X+/JDNfd
HNheufuKOK1hC3iNyQcQ2HVr4jec9IJG+m8K+YBuyR9ZvUKm84Yc6EYwh8SGjTdO
zK6X/g9Mw1nlNOqKnpI+KHwkk9Ft2UB+7ikhJ51gLryhRZdq+sP5U/qbLnRFYtQw
5IuSSVkjKJ8ML7hmHhq81W9knliEZ8XcedvhISkwkILz4C/DX+zOGJKp8R5pkx7T
AZ+giSNChziIpPo4rHT6UjCUJRECrq9QbWhfBoAgMP8W25UdyVdor1OEyImxonqQ
o4xD57DnGSiHQ4dVdhY7f2BKBcsAevuCuRdDOGU1BrEjPFPeX4Dt0YrO13PxIDg/
NOYUOkHM+tWYbMFZTV8p7SH6r3NnXnnfZVHN8T1IbfE5+/NYQ/5zQdO/CF0UIfx3
1WgMo6ig7hMbm61RZg4oQkZDyH6dQ+1M2KP1gn2mCXh0SWCAYfXbta822L/ULmio
iaj4st4fFDV/yvClgMfY/YeG/3oC3mM/zrwMxbf71BOadP3BiUHyi9xlWflP+6er
ZwBH0JnEwRRYrKw3YkdXlZWQNEbPusy4/YPwhXnoeLZw+sTvePVnR2bAzWaqeXrH
BbLFN5185fPPA5X6JCj1F5UwoTx2XX3NAN8Gbza5akG0zCgdV/2cDVKjylTKsxpg
iDTaVP2b5dLZNcxIY5uZ7bPAPbYnRZM+tLk7QniCNWlXUpu430GlGtLYsQ3X8rNb
5uk+/2MLocBeLu6hSM3+OWqJZg+h+Y3mB4Ur1nR71qgZW3B4QFCKkvsNbxH0jnc3
jx7+f7DruyzZfgCGAd9hzia/fMbDSSAmAaYHqXuUaxSZkQYpR04bP9rX/8WK/DAl
Ho6r845lhAOdogfnMzKn3Wn/1mOZxIp6AyCE3xPVSTLbD8IMpI8QKQsn6z3ZvP8f
lQXQ5Rs0ZtUe6PJNbYm7kDmrtnSeO4XWsESge60Fp7u5WJMttpbrVPtYKl6+t/Qe
6pCFRNmRDRmvgLIFiw1k+6vcY96Ye8lfhcEiQr7aVDguxD2Sr5E/TaT8BPpiMgoI
MX386u4b+amPeyDuWWTlFBILw3SN6UrGMQoFyUmN62Bnpa450H0i9965+cngqm3S
ESzWfggFPGOlhGp5UR42zkaVDbXKSfaWK6USJ8lBCmQGDMlETOJFvuvtz7QfU/yu
DZat9eEgIiT8zSfgO7G1LV5MXVAqGDgvOUWt4mdJlY9z0gCMHVoEj2uZrcu1pn3s
qy4RfufKdrspRD9ESUHD3f5iC0EmyUNYnLHwpIGX+gfEABewzFqrQ+ddIR7sC4zC
fLqTwGrXiec5wRlOoa9/scyqCXYg4C7+Jbtcxkpr3vgeRhzyu8jWUeF54tSKL9ID
riLMu01FWWGGeCnLg4QgVle+9wp0HuY5GA3gySMfdwUJGjGZzLsqwEHhQtfeit09
8HS+uj8bxHnA1FA8Kps2a1agIMAsdzNB1CjtzPu0lhU9fyME2bFlqnyOp5XZZE87
YDVj9FNWeF1jeKVe7uD0/97Rj2Msm9TJKt6yE35Ccqaj4UpX195pyNMyFWFpoDu+
kklfkc+zu7zRFikPXLGFywbat355xuS/cirL7nYuTG+q7aeMoJL51H6g7VlMAUo5
8bKRFbGM0DGBb94nm7o7R0uP+3oGwuLRJf1zsstORDOQXM2wdB5ZuJ1XmGdS1/fh
6cx6p0bR/yo2dvP7CEWuGVqZjDiGT/eejisFmQ9l0oJ2IffEsbEEdgio2UohpFty
dwImb1CWcCdoNxl+nSIFDP+PnKD8KEUYtmajIn38orrd14jifw40kwXS2jUFY1on
Y6PP9+tIQm4Q8qDHSTid/KBRfjHgs15/V6dMX8jQ/Ci92T0VKxae3w2jc18L/7U9
6b8Erh0HsAnDbB+5TgXS1yHMtoMVanXKj0t6Xx07fw9krH7M6d8y4eflcfHo9I5K
PyRQCnxCnYIyVLwHaCEZNq/9xqGGPGrL+IRrjLE8K/850IHF+1tUzhNMYMun9VsF
cfhgA2r6PiW+sstXbXa88WKmJmkNNj2R5RbEpjPSpUEl8j9WhZvpNzFWwEenEr3p
KW+YX18RMQtGiXB8POlTOWYrzmxsYY65O7g6mkHo68wSCYOV/VvunXu5KZ+oem0S
zh4d8+hNQmERiG2WcAMVf/l2fnLMXwsRmOBmVtZMPsNSQffpNmwblOJDQPTbZ6zJ
E7JFKHKB0CPQSCYz7tGjMDaWXlrOjPfGOEMT0bZipMfboP0M7s55Uq79gV21YKZ0
9aWbA0yktU9ztlyzcuJAmUw3TDqCNlk4RxKL3ou2ondeniUmBMITigxz2erhBUh6
MrwcIYsgrUAcFuW1aPqsTvjv6bYckEQ1iuDyfDyM9RY5iseI1XACHekSdyULa1YK
0diX4C8l/Y4KnIEPSTEY5ywCam5FQ2rN6/Qo1jgEFD5IXIjmOqjXdqTB7CU8VakC
2egKS7XKQKlfTtG461ss8Sa3BRX8VdozMrIOGn4oonsiHDxKA7OapJLfBiw00PzR
z9IDCt2RTvAwLyoqyHowE/rZ8R2BeiRMhQbqIYUEm3fJg0gRVzBQRGojcxofJDWa
Dj30yTTDu0HN3E2fgVjhu7g36kmazwspnsT3nAX7fyB67kr7TSsnACbkjAk+RrJL
AX9WaF5v2O0chBZ0OyOnJphxT418Qo0r1t+3zA+LfkUjQdZeQuzskqbyMWfvZKV8
zo8FfFcrOFSICkQtOq/Z9Z+xXMPOkxpzpBEiEm4Np0+ns+A4U7bjawpt2HUTC8i7
Fk2uYDkcLnKM036LJ7rRzKnC/CexKAf46nWDGGC6+hDFchuZ5maWIiwrDRj+vCxP
O5nrjUPEyF2W3bnjMVgYiBB8PJuEdFl0LXDzTz+GjcjKL+OqjvinKEEBcOgT4GSa
Rqz2CR1YIKrnvkAXgxukSeyl+hMsXxLoBmVjsJPj1pvtthKKqCFoTGh+9ehBJyOj
2zA4z5UNsEtpwWZCpTQFkFWNLyk6SIWGvsxsz39fHGUo4XcGYO87UZlGsjzUkabN
1bfVojhnoBtm27BVL4gvMWGQwP9wnc8tux/AANhesLQ8SP3Id4UhKQbRD7lnERJK
o3wYdNR7wIi3l0fhDCVFl2Og73peKSQr0apw4WFHiACmVsFfFJb4tiNDtJ0Qs+D2
oRX41qA4amSdQBANn7nrjqONrTBRw+NwZgCRdsP/jHb7w69f3op/SQ1Kg+0+IIQX
/ShdeG61wFnv5oLAY+I72voOwujUdUtQw1a4KTIGoipSkhwF9qvt/JwaVMDnj6Rm
YJpEErK/+GL33oz4CLjMnZnGDpn1BKjEQG79Veqy3P7n4vrn7viLrYMTmGDodDJ9
dWGG+zVFnkXw70NnC1KzKAsyku1RVfmSot0fCdiiUgYrZiGJ0T/T+Oo6ZEDemrF4
+3HSVZrZsv0ru+yWbxLHoAzEcsF6jN7SrxiHz+yWchVCyuoLQqyO0GcbJrvChpo1
7wnspCH21aqZiuP/Pozl2ya8MraQwmP+4gLi5MxJnlu9GFHd9DZJyEtNvx6g2bec
iTvFga0kolAUZBX4ugR4Pf0A2J+1ZOeJXJuHE9M9PSPYlQLT0O1WMXhxlUjJj8vL
ygZAarondmHFo90aA/2zJaCmSsFqZqIjLnqa8hM6USTiM8G0xxKWJF+kDcaSicUt
0lspHAHWTfwi2p5PCnyUYpXkRqOAHWNg5jO4NoGhRodABLIsdhgOTx78zGjnSx2j
iOgy8rjmAN8c4dnE4T0twFDj9Shljka0kz/LOknxCySCpVVtlEvAfzzXZMhW6xBp
MCz6CY4DnResQRsTH/UaM4wyUdn1orzW5Pkgp7czfgLDmsDr8HH2vzUFjcO98Q/f
uArujsN7CaIhC9JUlOkKHPLEb2XM8rpHvsPVOPBDi04CNIb5wgRziPhX12Rnmdmn
OrghIlPCx4Y+rEe9/EhIlDGU2+3BWt7bzYNWeZ56T8wOMPxGQwD5LBDF5N4ILkvj
dRhAWNigI6jLm4RWUSSIK11u7liQ/eTCM5mtURZrc4zNsR5AbRVeNL1kPxU0nW+y
zQ71bLBwkBDLFAU8cm4IQAduvfJX3iPgyRBF9sJlBxdSYJX4vG5zePhjqtVJlYZJ
llLoCIvfQBpblyGIvkPmKIHZx0VVty1RIyi4Osy/BRFiJl3hZdaxDCnt99NYL7XK
tEdVZp6SedA5OMhk4VeiUyXCmUxD7r5cN1CN1mJcqj8b2AAeu4lb4H6IlNAxjUHO
qGtGl2eRx6J3e1uPwGGpX0ycXEQCRB/4+XD6lqaQ+fnQSgzim31mokTrKXAJKeKm
wnVw1Cox6o+BdikN6GfvH6RR2IIjQnz5VlmLe672i/FUdUu3xYZjxY9u/TlVBNNc
XnL0eAYc/lzP0ffxZD9Q0prV8ujCLBBQp+2jq9iDIwz2QkBtMUiMvwf/Be3CtSN9
zmi6PHjSu+CYkZ6OmBNXfkSwEqV+235TtMS5G/Cp3Lz+hCtP1d866bT6/tHGDXgB
NvZyBevjAfoXapNoHkMBIil4yDSRZ309gWcFSmIztz49/nkpvx7yGk8uIhsLG0ny
+ZbZ0EY/1MVuo4CF1tYhZw9X6oiL/zCdHLeybkt/Vmjbn7LpUMXSMzUjXo14aGP/
iDYMy7Q7rw2OuBixlNUG3ABjzPR7qiutT3nx3qFm9swOPR0SGQJGClKpabVbD4qA
PaMVzp859n+L0eYr5YqJhHPJSpbtLqKFp8Dwjl2RftCt4QNg3B8Me2tH81Dw9/V0
TY+SnKAXSTO6G3bLn4R1uy8772gdCxIjyaP54m+ofoydR9hYx5vehwAagwk93rk5
NNTR1SQXQpIv6jKTtS6OxZ6YtE3wvzHKhW3ygDcTo6CC+0C4brPEpMvx4SWioitw
gdYbvWRbfCJCbWBME9SrsxPOLQnOqsKLf/zuBx2WblGlaT8Xicw7uIwrNoWKdYd2
xD1+2oAwd2eDAP+0vEfnTfWpRC0w3IZb+EPPx7V4yBgRtQM8gFdUyGiagE7GsSQx
yjT7SluOR+s3V+lbxN3vb3ibOEKpXaeSKYdqAHUR1EzJ6Pxy/OCJngyAyXN691ax
TROT5q8/lVpCaTgYGYJxbi9Ve9zIe8hvnInk/KluZ1X3f8yyp9vFIT5Ram9RBKe+
10EH3NLbgkJDzjeCl5c8b+iKlwiCdY5PMMcOukl5rb+OAGiVmJ3MWEqbzdA/zCrR
YqK/C3aWiA0Fh3TgIy5bBWFqQCotOkA6tRn0HSvcApzMh5hIQvOuWzX/jznWiEbo
+LPXnXanGvqqsnzEJ0qvobG1ptbdYP5AX6sFFjkN8Ss1x8URlCOG2jw+odTE4VrU
JCn8jwREIHvVU21F1RQMk6z/hZp9zUBJrxsBKEyzJvkWUU4iwMQ/09shf08WmdMD
6iiFKq25GDiVGcK7hGEnC/rQhUDtaM8SdHOSGvsqk9amrsC+lPlY5T1FTE0bJHfD
/tD+7pemDCLLDKbfy0sKILjLrvmsclncBKMCnJHF3NiyzcwtkwMv62Be9xEWhS9l
BI0/Bti6BtKEpD9b+wPWk6tjDvLpedfLML/bGCTef5/oEW9ssRK2flhXFVQhFTE8
j5vEYWG+l+o1nWF0kkEXqJVKzgpE0lAORdDrWiqEH4R5JjxqnYEX8kByHc7x/xmF
MM554uvN94oOq6ppmi6CIjBkx8Tm1LCRX9uAuTOO3FbQAhtfT4UycYpH6ymAP5YL
U1xLz0uQAW3mrwnPnOMCAQnU8DvCbe4/Bo+1n+8oaVPdMKWx3BPCs+BQdKktoTXx
HZZYJKJ3JlwtLkEY8BwusEgNmyaCeDN2GxBDw5rgmYDMuVBAVtXo8eAt/D/bKYRo
/34+HAggoPMdQiQbNrEPv8f4oTohpNFLsYUGlriBV81AZXziPcXfClQVshWFt5YC
NbuMU37HDh1DUPdrpfBkfn/my/HZJk4yoWlwdE+SfAXNQ9Q1FXQE2zk48OstoizQ
f3W1+3sWzzy/ChYdyZQRM4T8uV74peWnM3sHZluA0NLoXvmOXwUUmBn1j8g/ybtj
vXLGM3AUDuihqJAPSXrpGLoNwlfSXOOijV4fd1nDcsDkGerr2++wRVc1RSLt+YyV
vkD0LGsV3jxazIXTkALEP89MWeuAIWkOh2fW7iSyCplsWeqtHKTwSWsN1z+D06tG
zkWnCqfpdORBBhQaZRHZMzE79uyVHaaMf8dtLeQcv4DXo2ShKkDRlO42afdYoogJ
Oua9SgfJS+47P1nuiD1jDmEG4YIcE+Zh8wWi/C+uISWVnAjdbo3tRoel6LgdZlFg
yag79bowGKvFiwnRpNvIXYis0gL6oOGTO5vvTt1vazy5n3HGKYuBTUC3jPtO4Su1
DO1WB+rRsqmkVfDfpnu1oNlwgNdx+Wkv63NOYMJJIrnTbamSGGdmyO4HHMZQP3BS
EMjlvthqto1/5vIlfLEBGuxUNsgsFKgdS/f+Pn7IyMU8e9kdcPPfc3Tk8W8OCeKv
WpGn0n35oZModWdGVHO795wGwMAak5i/8AxqPWMlrfEjRoHCLsNbR+bhRI61u891
BnyYnXw6tYgC0+jKvnsZQiDffI3Aix67VTwpuYG8uxeMqnwuj5MyZgjNTHPLAp/M
42wxPK/RoTUF+r6xAH7eHo3MADs89sukwbg3BqspaOjd9uZN1lEgdHXHH0J3e08W
+lQ6/QGye65Ua/9OXw8JmXN7L0x/f3IRbmisTSTvzhtVYG69A0A7KH+g2cQsls3h
jESVJL892k0fQWZhzgLdSTquGfw4KTFAsXfMQejcQb1DYU1fKi6zrcXL7FSBwxIC
Lor/tQwaJXWZNSabtLzZ4A5RVYK/79dvmcYn6mH6JIYdW6CNKaz3xrWUAni+/PsR
wbSJj3hYFnoQvMXW1m9NO04QBHcRHyJtJvFq25EFQ/FLgy47bsJ9B+JoOoFfTGgB
XVvwbfzQUBbxBM2cOJwH6I9ZPM3uBDSz8cb7bo3fa/pCe/V13w0UIx7miUOvklEu
R2c2R2cdETF2HsUeq0Ku1Jczf8uTAvKCcwbHYTjvSyZe0IrjEKaeGfvMy4VjFQtV
Q6hdrFFQjHeuPdICHbgbe5SiSTQ+EkfPuo3jjVqylwckXPac83YfieWgGRfyBXAy
yjPQKWtDdnTZ14zQgzpmt+wdpmvrIvfVFvm85v4RiMQk/DUyXuxJY3ub6o2rReoA
xvEJT4UcnE+aNaeRXcoi+fr2D4T+9/S80zbXhuNU6VObCpeaiVWXSwO2420bQCf9
aVcO68Fp+AUnNMTHpcO5ATQhNZNaRmRB3KHa9L/sSXr90kaQDZooCaVXzno0Vh+K
2oSgmXUtnSeAEe3qg4AcKWZsPC8DDdoOXbPJL1ZTTa22wBnMh9JDLgMmYaZg5J+o
eXGOk8naNgkpIx2mz2j6c6qDq6TaawWyeKxrGjc0u3C6ZWekmX1jlWYJj0FwIbOg
36P/v0wO61cUFAGfDx207ILxpW6bN5ha/FT1kzUdyCXYQY7mHTzl0Npov8hlwigu
DduOvI3k1MKG0/3d7qiTrjO8VRejpFyJpaTRWaxv9Dc+JksIPLOPx8x55ZspyXkw
1fY4q12QN6tiTf+j86RNd5NIEx+6ntEXldgUF7z+FdN957r2Ht7s5j2et7zzDIku
nriYq2MKZv9z/eq839q7As5c8ezHlBEfJB+j6HJpILJPe3uti8hbbatkOK9me9Bi
v7WmWL45v5+IL3OTMIB/bZa+uW+uQvznZf8jyFZQBMSiS0FkHnpDP7ZIZcSZlC7h
fjbg1VvHn8b+gcpSmc0+G0VaPQcvpQIl4qTHDd2KM6xxZhu0wdZ+dOfGZK+FPAYh
dInrJPPgdSuAXvGhyYI/aEzyv5uhOeU2BxZ3Z54n/eg/tmz8n8yWEWPo614NP2yR
5/3JUANsYjQYuVY8We8+UtRXG7QOUhqDA83AurbB4giZswTd/3d9Qmy4YGvUKwTW
lV3xmKlV1foZ6zoGXgg7cm8jnuzT552HiCj2VLEZOq87FBAikLS1qAwYRpNhXZK2
twMNpLVr7U2qFP8LQTYx8FLlQ0pUiVGkA8GGH/K1W7Fj7bbQlP5m5W4SXWeRLXxz
uI0m+MF2pmhO2hmc6bRumY0NkKddAELGpGI1HJi32of7DQ1sB0K2qYFUr4WV0clG
f6QowH6D5nbbnXGmFCz6JgoX20d3V5VSzWvt45U3tDAqwaBBZe43ZwRm5CxzIaCj
FAFjoVmxwf8xgkKU3o+Yw7iIrukAPitnSJTcJ7NTQRlcEBpQ3lPyWL/i1tLha5z4
fVRuN4rgmtlh3Dkrpn7i21+rMdI6ul66jqNfamKCjF+DIaEfn0BfQsgAkEY+asdY
zyS1BHAN9+Up0XsE7RkWusZk3mMNK6DxTjRiC2TUOddc03RpghdYJFmX+745XSML
HVGwbfUb//THh5bZuJOhV6KJ0BtokHcqz7Tsmx0D92mzfDg4JMc3kOVq4ojgJtPT
dtSPQXKfNdGvrF2+NJiJFvD8cpZdzs4i01wu9yN8CCFnogQGrGQ9R7WB6BohRdZv
6Q98B+jhpxpuybKY1dGOFsBl68v+Hg6ki1p2CE1XjNm/zH7TOp1lIpAGXG4DvWya
3fgeqWik6k46SsSnoKcjRMV8jBQ/ca6ZKuwTxZXJOEIjK/7RZZS95QgrmFm5OG+J
dWl3KpMFjmEikK0FuM3vIZ0ulrlhI96pqeX3CXfWmv80gVaqkwDNCM7BUFkEl4wy
BukcjNsrn76URXkqYPghX6hBvpZGy9G/cM47rnfIMiStivUGqv8vrl5tQgv7Ve1T
Xwc+2njRCopEkQzT0x5lfkgsWHmu1x2j2SfNucAnfydXJuHqsv+/0nFBruNuGNEw
jYbApYkgD45f7h+L9ngkBmnb9ymt5E+DrzVAZq+LyEOKCMSQ46yK4wwBcj2fiNit
RGNfZhHZXidRkhKFIrH8JI4rAucSn9In3GcK8mo+2SBKF3YRRPvFRxrSnmLz8MKj
SJs5KmryXx9ZjU+jpbvQSvvK6Pk9gh4V8VQlPbsb0ssBQts3z65eMXrcS+bRjnfF
ipkrySZ9ODhvUnfEqSCd6qpaLq2oYQpoJCa/h+yGpBzpXPZoUIBEoat2BoxQyv+1
ZwZ6M+KzYafX5URVNA8Ki5TibSXv1Pd9NpNtDZAJz/9yppc3ym2JXqYzusUVAKBn
V5+b9qKrIRabj8pz2KxMESSaS8YBlonMygOsyPuGQQ/QU78EzvlgmIKNQkzziJHt
gQw8Q3os8Y4C4SEZmd0rhQ+k6WFk9LWKuNUtX9zIRpODDL2n9qnuoi8/ZoRAYj9L
DHNsMsbm3qGPEfr1ACa2CyBmqxyjECDFziBAOJ3SKNVn4e5FeoJx1B4qsvxfqpUc
rfKaADpmkV8dnmAqfDyd0JBofiqPGzOEWpD5PhfTlfAyGBxQoy73Lv1+cwWlaRtt
75KduqAmMhxpZ4SuVMoHubPI99Ff6hWiTC4zniD0RYTtlT6WAU1DZWko+nzxhoPw
SbwdFTDDcM2cvLW1FNbwIBLHpu6jLPv31PaFsuV+rdGHGUDebnDTHWl/xVgEO6Dl
8Gr/XZ7fRPMpK4+dtoX33ftZIatn69XtuORAU/KRwZY3866zMyU00hKo4RzFFunG
FY5khFJdLx0AUN1MzL2eXcYtgRa9ZzYTHB/oGNkrVWQ0PEQR6bwl2oP4D3I6PUJn
GAP+byeLLFb5UPCZ7IQHzhN1fuVqAePr7AsnfIlGkG2wgsx35ggo2CYM9W233t5R
Dnj+n5aQzRzY1n1DewC/5dfxPOx4nGjoW9T+H8H2ygw/z4Kt2B9KP55gbvCESp0H
3kqK+ls7KJb8EXbSeY83QsnxkFPgYrneb7jG8uS2nHVLYbylhHO1IkcKRgse1a3h
ID2uBzRgbYroha3OGmZyC+DZ39fQKYGDKIFRbNo2sTPRm5y80MTPN7mGX8wFOUo/
tW1GzTtAEjOSzOIVSMaMVfsx7L0FhgO3CrXrFossagRKOo8dW37qpqr69Ajlm6p+
R4055mezFMWUDn3qeH52BaAU9zglCpfuDiF7NOtdZ8dHudgYDJrwzi6fsHxd2wCi
Hzt3VjDCR2qeTxBSkaWSj4uuiPkKq6kqlqbkFaUmMkm4Zuj/4Gts9aYAFTHmcK0q
5Gh/lADDl2SVVQogHx8CKF5kiEVkks3Xjv7wCZtTX6pwGxjEdf8kX5e2hRVzNPT3
Mw5sp2jJP8SaVkn6L6H5XACI/oWXo9Adg9avqhAyMkP8M5J37ZRUq3UPpxLUrb2y
i04oWqp0vQSUevlNaJ9Pl9pwGdsX9Vdig3wG3mEM1VyReHveSDZ0YGxNYOaKjfX2
D73Ofue6ZgZMCoOB/aXFAWhKZ7SMZX1xx3ybpAxgGBxgTJUIifch3efuIx9J9kSA
jj2jJ0wOTFosaZnnnwDv6wBMNfPBBTxVI0wNuq3fZik0dTpi5B+umT9eGzagOC53
RbUoFZ9sHg7fhnNbB9avXDniCG3RTZKtMBUI29Q/xBsgpV6gtRH9bSM1FpiIHtaG
ZuMXPj5nB+OOaLHgg8PfvzHLKBx3hjjHM7ekaqAchx7+/eyLuhO5vTygFnjBX2AZ
sL9z7moUmvBteeYIkuTGNKn4V4xcTxlS4Qikdu/kd84yHAd1GhUOgppDR0RkY4UG
8PimHMxq6GJkMSlPc0T9jeq+sIOf7WM26SIULLZapXGP3jknEUjb1JSXCkqUxojg
UbHXB0Huf9kAf48hSU4/L2m1JB9rOtHV8YjfHV0W3CP3OWgiPo9K3bxpYKknghFR
4PHHMbvoEpwJnTC1nng7Mz/opmnrU2xBxqrUiIe22Bd/f4FX6cwaXzFIX9xdclNJ
Hp8O4so5y5/NA9kABLePJ6L+rZyjyY3rYvbVO0UyHSxYDqsvzqo4Hhl3nlkdhWXB
Np+OsqGIByLf5H9HhMvnHPAXi+Rsife6SKHgeX8vK06QJsaVA1a+tJniybk7gyDb
7beeRLBYBPbGUb3k1auvnA0d4npQaTNniKG40oJDzcsj4n9VhIgsKg/2UO3k6h/p
8x+m6o0TBcAjEoM7DkHBocOL/jXvnlusCCf1FIUJjaJagYht9jDEgP/bYEeIoUTc
99LTvvq90jKnOtxlgxITQa5RqdF1awaj4IspxishSFYDTgw4GaN+Jaii2yfv99Wf
ff2az3WpDPDmJb9CsTSsXIrsI87inlihhsMrh5YhJGE1uyXMwj08dVlUvXAlffH3
xuZW432Pm7taldYVXDsUkvyh8f1Nyq6UNkbvPaPCxn849lplhGRS/yMA1A27B3jh
06O3dXz0/SJz7pKJ6H/fXtxoHtue+vRMagMXuzl5ir9DaXtJc6H3lRwz7dAWoBOd
A3/Uh4SNyxMx5yQUHxcDmvKkJpZ89m787hDLW/VtEKhtywxV8vhkQt1SHv9Kldiw
i7w4Z2qzWAfRiUJ9SMhI/Zzf4EDiMI8E7F3Kjdew5eAiNB+p8iQPx/scL0oUuh53
OHRWwn+FMeSsbtMu9oEFMgCf3XkNvE3ntfztv0sN11ptN9NxJsrlUFSD/+zzkvsr
uM7Xyxp6itVw6LCYSh0U/dVmQcMj5Arn5t7DXJZcJMupcuTgmYWxFVJZSTCAfuSJ
XdAzXSxLTS0eMJmXmBBL13rS/qMjg6rJ/Ihtk38nFxlaI9sBYqYrLFM4Bez/V8K3
Xlo3LvenmzmKNoVaqTFWQtltUgLbF/10km7mYCtr2423BqMNFTGLcG7ow1BRoyr5
HvJ7vPcPjHg6T3AKofaTOYJrMJ/rKumu5SlpeHPj12Jo7sNtptx8PW5MJjV6mfFR
RAfJn7bUJV3iICuzlOt3dlOi6NgiuCbuvJVtnoM9AGU3npn1yNXjQczXnFw7I283
QsJM6jW8Xo0bVckOh9FYVXi6L7uRAHNcXaCLfcDoe6TSwNjzQxX0yDM+gvsheBzE
zC+/jj0NMRgao2URmiOF7FRA6BpFlMjrPofWGgmesK2IgcLy4vuYAKD0A419UNL8
0IO5WfS/NGOd4FCPW0CtBJ27naUR+Z/Fe2lpRtuL424kNDgb1doz3/Zhn8KrmiBM
wmOTMSw4VV0QJTlUfQHzpyR79eORtYXS+oa0j60CY3G4/zSuTk+duK0nlV1aS3nh
xmR7rydC2vuABMECWWqSVJmKUthD4dki1/KMK5NeqdI464ati/pcSBHky4kAKQIK
FwY/Yd9nC5iKf0wPT8x+rzon//69HxHH0jkGZglOjUH2Nb39/Qw2w7x5YjRBac8G
Xlg9z574P8Zn3MsykJSQPcNPAl/JnB78Q/+ZN1YFJazNr9XwIihvs6Un7yh6Fvsx
J3nu2gQ/aoksN7XbmOTf6YGVSmcZEnr9+a+LiY8tP+cnVYkbgrPQUJzC4k/iHX6N
ybUxdFLzDNyo3VSyvjKgb2Yv3CazyI9G4ugMODiemn93BnFf6YOEsIFbjfF/gGYs
44A1gY4PBLZh4WftPBPjOXNpRjFRPdtwg9GbO9LAZOWPYq1P2OQgrmktAr2Mhpun
wphqFBTuc1YoYB55A9J0TixQRiUFSB5MDedd2M8j4hcfHr42aHjDrjuyr1T9N1jF
v7Mr2WbMEm5iHgdNs67LyV7GfCNvCvuaqyjm9j8NP+CxQo+U/NEDFLW/O2f7rS8F
ry8U6HR+N086wZbTF+9UjGK4vpBn50h6AWrkGW+3H+XF7iPlcwOScfeGjFnCoDTY
oKwv3d4QrUiAk8JdyHIhaGcFBM9i7NqhWTSqtDnx0AvW92oKrN/kuKqFTyTDzd0Q
66E5f/4KBihBnUZN1VCvoaRkuWOV89pD11EahCbrbUsBnUKJgQnzNdDDHum5lb25
imZ3Dn9dnG6LOpY5APzss4klAg9CBkD7l4fHdU85QHVzfqyHHqTmnwRRpVB91uZB
1Zb6NnHGAyAchSTOD2A5N7m4jnpjKkgxRc1vR5blBRA9wJSYp2KbExtHoN995iIg
LsbSpPYgS5dg9qdlxyF6shdfeB1ArjFNGbxdix0oKYL+PqPv1C0iOYuoMtEaMJWA
YREch5oVdcuEngOHhwivwNZshyvX7GxsCWutHMaFF6tIu959PyjksL75cBzXGs4t
fVnvgnSKbPADBcto21JyXYkXtTLnHVAXq27fZy2YU1jU4dVajvb7yfbx9HbrfCFV
lCEaBx1g1zuUe7ml1Jr/FeW5zzc5Z4Y/Y/PW46hDrvjmDQBtczSrRf17S9oyS0r9
0kuYXSPxncQqVvBV4myveL+pj9oJ9K2ofEx3MwZX4dcVm7TKXlykJ2yZGClqRQZL
t/7MBfuXcIkusn10KgcMlyMrn9e+/3N68bvzinXOoBMa9aPO52FQhTOiN019oXov
bLtR2/zhZKXCuDnhotQXIbX2gKu4tKyEoPMrdcWQRtqxXvxQhC14T7aQAJmqbFwr
OV00pXyIXNHczYtBdwbiZM1kUG9w1g8WgP77+LfmQka/VJ5bXl5Z4oA67JoenOUD
HUPHVaSJdq+DjUfiqQ3kkfFOtiXDNeuuokVb5Oi5JmeSy+W1zJJjcCtryeQKuuWA
49KpcABQ4pJVHRw+LIXWgiHYond4XtMwIqaRt/NyEyM8u4w1G6bMLI9nTB5ZALgS
mLkTNS22JAcD9Q8RpMMx3K//EWtS1xaTbIH7mK56ei7ttmeyqecVD896YBFknkef
HpYGGpzQSLNSXDfTgKKG/MbGsH59dFJQJ8H4u9ZsCwUAkf57+madcydK0DAEMJgG
rCEDomKGpZT+RfLx0sBxVsFhwJT//wLKmRnJdJW7uAD0kRnESxoUDERuc+xWmowm
FbsSr7LvqRzWwpc0dzyz6Fp2uQuf0DrP5TjxzI2XZiv8DphysPlOtYhxtj9yvf6P
IAsp3bNBlF1RANZX4L3YHa6IkKwW2q5pSD1n6YotykdGUZtCKqhvaDxjzLK18baX
JG7ZUUIyxgV6AAlD/LDmFWn1SiVfD7cXX0gj9d7sjFYuJhYO1l3xqWEHSjOA9SC+
C3RSZraNxoAAgYo3/q4xm9eMAGKYmH5nQ77V8SQLEnBNNyUsUj1jRzCoBwWv57Zh
f30neZdkjVqLBlhKPpMfSJUnaJj7aGtjxICo9mZ2L+4xkgSpC7trIzw7UpEBeY2u
zyIFHpQdtUgynvw+48Dazty0L8CjSyLoE5U0ME8/4iZ0P1iHN7Ex+CwBHq0KVdCz
QqVyTsG8PTKrR806X1JEfMWnxbxLkl2/JBtUiZlU+XcCYAdCSGJUIDkj3VXBcoXs
5kRDYipAy2NxV84BP9dl1BOftHIYb8Y7FPGWEL8vSYjX+Y+oy9zj1lFPLdmgDxGf
pdAm8q9NtWTI016inGg+wIsh3m3+KZDYWmAXsEt8c4xY8lHYTrTGx7Ypbk2vyMx6
Nc8s9MkhyeMqn88nJZVoLufjd6dl3+KySElRl/E/X+m7pUvS8Foz6PmZyetN4juW
K1BWyjVldrkW6TLjjcjTB0QxuQ2vFG94ck2MASmwwSTD4T/imrZyxNe+IxPUMZFR
DM7JG0AlEY0LSmFayv1/Jp4RsnuDzXmXgXgiMGGVylYPH3L84v6klTT4DEjkRqVH
peG7qNVOU+4hQISalKXRN5chKH41HRf7rgcWBTUUpLndcIWgdtMBWXHcxz5g+6Ej
EwkV2WNm6XCiDfnFk8s7chPjSxjjElgqwY7iv7/6Rl9nH2mlOkDQ2nXtm+MHFWbD
GvO17vadk2EHLgFMNvKoUfVoBBIwIqPtP1R3Fid+8zYpYXMDzYZkjyH27MA8t92y
rWnrkmsZikrjlW6CjeerpnFfSFuA5/bmT5iuF3KREgDdCc1hCllSxc5aOTKB1DCK
q1vjG04AhDT6Bz9xJ2/cfwm2Bwfgd9kq0Qi8jtEbwVlGamMjRFs7pwJWbKsVuZuU
VNFO5W9l+GS6cJdpsDBGLQyDqq4DXFOoqOysrmQoO/pbaZOU6377knrgWE4NLWPo
NbaeRVEbaXT4qzOLs5UjrDaeZzfukqcIFwly1+NN/SFXw2A4aajG1uh7m4q8gyk0
21Afzc1l/hWRKBSvg9qFQYheM6uKLTSa87sAnxInUYc7oBje8o/veX5exr2RYJwb
gxGlO9/tlKWnExVIvL6I0yhMSPBybI/Jh2FCQtoD6V5HgPM8Qdq/+Ukcn4ZR4aTY
F2CCokbNC2VPMMNPb9VB5InXRfDqOOUw2gHf9Brveb2XfasiwiUwN80wLqQJkR1G
FDiYa11JB9PQ8OdxdAxQxz6busL8Ph3cPtEi8ChcZkvGhSyxOW+lNq8vAcKkkSDU
DMJKY+q16N8PAVNPGMjev26kctRU46SegHPrVB7Eh43NwNFvOKX7Jynyiz02SjrD
9l0k3xAvN655lIY4lBm9RqZ5z9tXCGOfu3lovhL9MyszjJ7kC5T/OrnUog3cBOL4
IlqImuTQM02yX9Jl/sovVclFkldB4PZrY4ccDHDSoyBZdXO79dWyHy3e9a7OB9HJ
5jJriu3i2xzMAMQeFddpxB6vM03AIgAwKubD9JcD0lzZywgYX9cttFgOj9DtnMht
nJjOy/wPMc6gmABekLHp01VmH+xxyIz1amLqumrTIIpP+uY8oNdvsBOyy+pZuEpJ
oFJMHeQlIco4JYYgJELnPut1jGDYPhHnQUDjq3AK8kc2gO1IyVyR1BTzvv2Ow9yh
mvogetzSHI+n5qzlX8cxzUf56UHHX6Z/DB6vR9bnyNYpY1pCVrT/sRfOVxu+lWPn
GHcRnq0/Ix7UqjD9J6K0lhmzyo2x2gLpXMKOYNmbyJIL5hqWo9aymOPxE+9Ezjvm
elRNVOEOsVZ8N+SGHLJ0AGKYeBQhp61NgGqo8AluRU/MTn3gvyViMk0Ogg/96E2u
elgp706DZ3JZWYh41meTBOEofj8r0kx9HQemjXdeJ//z98xgMS/ZdLxE/wMzcaMW
yBvQ/a9h5yROvkRR3zQ/dEs6SSTurc9ViRhABrsL1EU0mV0QDteEqNyh26K+kWub
ei0sOsjMU3/nm7e3LYINzs9nVAbtfJ1TC0p79CLzeYEtwnhT39WUqgN/52PbX9Tz
Ut7ePqjaBA/STqqSFCVT5WwcUJVsZa9nH5VDTx/wSPrQarhW+ftHdKNFew/STPap
aCRzQgQQAGynSQhc5xMG29/7rdrZiQoCqNbs2bpjqYEB2yZRTanISa0lT427IPQs
JpJoILzpRLB87b+c0IHriFAbEWAdw4QgUz/nzEnAdFdXjFeQbc7qKs6fXzS1+iew
0Jf4oXC4hqt7NJh1vEr/9pjFQAAZ/uCtoyNwfwh3v1jR9hT3B3eTfiIGJcpBiyV3
W7aHMQBhvpqUl/MVoGD9PPbVvID+mKDNS4RhSi3P5Aru36eTflIxP+/akWNZIFm0
0l7R+mdPMukufF7ES0rcr/C9+CJfwwojsFDgeXy6qKxgefqshZugvzXNgOdu05lX
3J52BLDO5bWQXAQ415aojf3+asQAvxCNCZ8CoR5sgSOwUgomQd76JcpfftqZKeQm
m60A217IfiwnBt4vuVTb1Enlc4SEMBbVSspY1QOZ2lZrM5/YrTYEinwyw7jvRsn8
e7dljcrotDYJcp4QREZO+bLAdTj3U8qLBu/56cYMpGQglVIAd5j4z8fNZOARVI5e
oWZScn4IYVj278EfZWZhZQdd4ovAcE4pP7+tgiefU4XckZQPRBC4/yCCg0EO6bGJ
OmXEDZZ/LYsjPy+yMOH+syy+cDHlp7g6lQxVZYYEViN2Zd1PPOACWYZ1+DklVuNq
y1SJ89M1unAjow82sZ36KKZWOwzXRjTJ96rd83NlELghCU6/anAgSEJAnacKRJCI
hYBlEtk8uIDBb4DhkSBBUXPPtVSqI4LlJbqgcYXv+Sce3EhQx1aozKQy1yU/5jgz
W79u0C2WfDX1iXXrymdZd1L3UNUDRWFAKtO8bn7/CSEQxiR7Mw2/pLAc9vtsG7j+
yE+xCBbeVSFDCs0sMGNAhOka1ptG1TgDNLmBsDeQXeN5G5ZYivBnJz9ycSuxGSEv
Z/8QkWrL8UF1ZAif5AGRax7/MunLJoOmGbYMh5RrmGiZQ05/hhFGO/Ma869wP4Zk
iUOLfarxNDaD1+cBE+A3z9yq/2KArpxfQ2hLZFnOIZWHjrWJlvWevtKgvbCWMoXr
qlAjrXGCRY6gLvrwoYhF++psCEMDrso4lKYW01FLV8OtvHTCCEz2Dr3EQxJymwhg
GUHt02Nx0r1ooIUb8UimJIe++y0gPdw7Yyd9O2U8xO6F9uJXy5G1UQOP+49q+EbC
RSYcG5VQGrR9TQmA8Wm5Iz6E6S3QihgM5x3M8EwWavyFFBbCoQR7KPQyu7t2Dfqi
SWSBEuVoPazOs87GbW+TjH/dacuZKPhTB0e265ZfWYPZTaVzz+ffOdYnaL5CDfdN
jUYwlD/TU/lgmByAxNNukjKB0/cQKSsMn5DUSyozTiZZizOXB2zjUln6LwiqhtWs
UMpHqwXvhltNHTpic+7uewcdNYJGIQPWYbUMbSgX9nVYwpYb0HUAqmmQyydHtY81
RkDqBHinwCm2coonaRzzeKBt7DWD7GhjfWu51d9uEDCCt+p9zk/ObxvRefBAtcFN
754gnu8gp/N5HMzdGJg+7oS7DL7cbpmu83UUqOiQxQT8C1vV9MK9DF031AKEhh0K
zXlyr+oyQW2ayUyh+fWdRBXBvHhqQvlkkpKZcSX1MJl8F21hvSztMgJC5i0GCj5p
MP8U0OlyA4qc0vkhGkUJk1rcOqJrwgNqzxhbWn0a2T3T2uPW1KJiVd7+hNcRzWLY
1XZGpyh80Dc3n3zOjY6jHWXD8WnHdNELfcW9yAn+KFh8C1DMh4/BpHj6rYiNgg+I
7g+oJbzrZLo5tX3A6azXU23K6wApkBuI3/CK8DAx25mdHygMCsj9SorZk39Yadlv
DYN3eMChRLlU8eXccI8zQbpurMOuL0lN7m51fL3O4m6QYkRzbLUOS5q1Ofva1NBO
qj4Mhc64NIa8tLhV/Q0FRuIlpbibYe/dxjDoVNGkxuiyHPW7dNzM7tdhKCtzfNQh
h2QArep2xZanuEyhVHoclkGsWyUdXuJYPk08BDDPoBW03Cna29y+Q6IHaTj/50wg
8jk9dM3PKiJH6ALoeTZP9gofns3zsGtdcejAxrPLi+OOoEKG4hV46SZZ5p19oTyV
bg9RkWWo4ZYoh3PUlTY4mF6f6X0JXHIPEmlv+RMwUadYDf5c3MUblc55z5sGj+G1
fsLLkeGpm2xYoUd4OLMJo0kF7C7TJUNHCSvrtLdkpvPjrc8LZOxttHY43RSTvYUs
btzheIkYXTRbxYyGO1hpm9HpQhaKL2spZ6qTDy6jzjwHSw8Zd4p0GjPwmSzyu5MS
WFuIrw5W2rf6VKTquaUgnd2Bg8zJcyMg2S3AzF36zEkZojuHjNmUf0x++VaPZXOS
aKqaYoxHVEdZJcUnjtF9abcB49dsgA/hYtlJEchkCxuEgP3dr/4YS5D8DC/7DFXU
yYqnO9k5ViXRWL3Pjr9kTCUE5iyGIrdlGge7P9OSPzEBZV0J/ww7SJtskr/KdDgH
/ENwZRnSAWWSiP7y+I8QQIS3Bg82CRMRAKUmOZ45EHP3RuR/fWALJMtJBtWZMxeu
pXWIDDo4qrvZfa7Tyd11kIzxanKUaDji9FK6z9dOUDeUSMeNm4eCT0aBYdQFlpqp
YRwWVxnh6ma2G/Lpun4raUwfc+IV5wvhekP8zmkGzA+uKV/0ndCnMDIL6PZJ+k6H
mDKKlIqc+stt0x7x7tydcn1ISAqxcPZuB1df27pUWU+8tX8Wj6DAizvZdvUi7/l7
n9C4DVLlnn+yTGs70Hp5Xsz2PbZBgxp6Cza7NIIuCgRttzXea9ZC6/OZxpOvLbmJ
cJ+kWrqhW9y4U6YxFUmgQJYgu5lJ5yICnsHtftIJGfJ8lJs7oX54PjGNEGlHM30b
uyR9CyHx6uK1S7Vxldno8mSfQoKUT2/ZuzBGD+QZNRtCThlY+raWpt7KZZoLXdx9
knIMaMotd4wBJ+HLkhZ9buhrZmkiurhU6FNR5f8qAKpos/Ro/HVlBqogCOxU2dgN
KuMAzXjiPXAxlpyksEmPzSlZETjGvYEuLELYxbuQfjvOUOajE1rbTM//nCPOzypL
xIXusQyzklNVqTaX2nfzn4zO2FvyWDLZNzixsMDfHzA5yic3ccSbiICJZx8NH4FJ
SQjxaTqOfcRxe/84OuJNwWKn4YNay1YVpjYhmaN2ZOJz2T2pUMPmgG+TnQcl/YRB
/KqPfHD1ImcI5OdbvdhJuM5tQ5j+RzdRUmu0agN+L3NaU6Mg5WkdyxseIOBRleQL
FgwjSzOfulD3aTJxDY486G/GOnfnrigYLtDogcviDNubmiQ/1TeV/njLpytIJCJE
m2PjYPvgCxWCk9oNYFxEdfvHN5nzke5ZF051d0Yd+Ep+2tBCUli7IpNuWVfJG2B+
DnolCXN+5QVLjdG0/3wKZLa7yIfQ7KZ51bt3w2comYn7iwLSjsrXuTD+UUhA/u74
hdO5VWbMpDsCNMoQlg1oXjsIkzj2NYai/4ytQBmp8iyh7dG2Et3hPyMAfh6W5S48
AH9DLSWOF9THnrq+DoSdwjy1DqLnl53KFSLrEZ1clyIoIjqN/x579bP8Kc+AnRz/
Ccq/arh9JjK3y33lou5Gt7FV7SxomC21+PW95JxMeukZTm3Nwv+9+XWvhyhkBCfB
yvK3ny9j0sWxPkTKiec9j61BMkh5iw3xNsqkTYP1pesELLV1pJ7ujY8PCbj6TA2G
FdqTgdi2aTP4+aB84HD/n4+LK1jf2y2/MbxcsL1o+uKkkN3pIa3kF4NAgmtK/w4D
OFOs5NeS34k1OoDS24jCcR2DV3SjPD6oLfmHPDlIuFMAcmjwKJJOG2+hVxLLn2av
LF5vfEGyOKzdTZjeP8m1ipOaJSQ7u4MuBqZP1C/iqquxxXcpGzzdpNz8eNRAxBUH
N//saYmd/j68y/ACJ9oVTzSnse3yfcj0umwutIRMjTTlgssiE7TIOYciOWYZSHvn
Ln++daCGmeIxrRcF6lPkO8mN6jD+Dc9xImBzblqv0lttmeLic+usr4F/pJEnMxtl
ktScSrb71dIJamirRF6SsNwLHJ2Fq43rxDu8QxSmIMkCkc1XQBVKVxn8LgkFQNFi
K/tY7zMd/0bPThScUnA5NxuHwI8ieZG6sNz/XzIuVEoZC4UVAzU3Sr7Rkp1qH2au
83oG1wcr2b0mY8KPv7t12GdEG34SpnB7pWUyA8FIR3pRo1ZqYAwL5ssN4cD7sI7E
7Fk127q9sLUHy0FOgqJegFRfIKQBYlxDJy7ls0s8iglQVU/wz+nbPcuLflyppgHn
QwAUvp7JMsSrEtuxMJ0g8RAvBp9b9gLix/tts63VaFv08Whz7FVZ3knbwI6TfnMz
jMttBqiItYix2CVF2xmjvLvir3U6maTSub1T2X+vCib35NZzX142jvylIjMQ6qam
LivVhlg2u4stdjGdzWnwYc4O3RGumf04ZUrUUoCsF/gJfHtqHLTCxTyTZWGNfq/h
hEq824rPhPC8VD6nfkVHwSO9qwRhz01t8gos8Yy4j+OH8jcf/Ps7joj2R3G+wQ5i
UFJkXXixrmqJ23orlC7VVigbbGcgtf97U8s1Mdc+Rv1VsgRefbyR4SSL37pbryIl
JIVva5j13rNQGkh+cMMpMGSps2QalUnJugGBW9/Bd8/mLqDfctNGY8PpiFgApqaP
/gRj42QMbnezlGDDnWTGdnTjCBouNGAw4HJJKZMcs8Ppgn3lPhPwG8z9K5Er7QhZ
Qs982tiMGO91nkFX7dyIDTz/o2qLoq848NB9HgCgsMlla9//c3NqDOxRe3nbY2L9
yx6TA7K4A3V3R0OXSzkvtuesXC1GMUYhMen1+R5NYrBnImz6+TmTC/kNvSUa9vxr
skcp1oYtqiqf+REYBtndjnOkyggxE28HEmTtUKfZwWSjUv8U7qbiFN0CEGrFhIca
bwu7S9TAWdARVMUKJS4WgQFlcwm96PVXHoe3f8Rk9uOdNBdXU0xg03A5GUYvV4gm
5dAmsdlL5mvPNTkoB+ybrtexjrJjR+HzPyGs8ke2h+h/EIvqzeM73VvRk5P8MnK6
jFubK4/aA7sWke6I2gc/v4E2DUnD79vpOJmML8LofP/cWv4xsv06N/cYm8YmNNiz
k8MsMOtoXuBFKyIenpDqv5n4TIB+5j5PzgQIhVVZ7YIXZACvkYK3ddtF+Ginxthh
bjX944q5D77klzSoVRGNUL4v4uFDfm1u2kA6El+ECIUl907xz/VxAejrWY1NOhvm
Y9kSoQQo4zYSM9fuNPGDfBlgM08J4Dvrx21Y8ZT28EziaaJxOv0t2DYO1bl0Ohrl
XR7N+XzKJzpUgqSBfh45qTZmnVl30UCw7gdjKRyNKhgR9QjJ/6K6gw10e+gqlb/o
sbsy9FwRvs/sNZ4qHnRp0ooQ4cSHL+29ovqgmewRe13DP3U6sDtiCJAjED6Cv3Hu
AstDCmFgP7HD17CRnZGU014tleUU2QBEjw5RNiYrU3+92SwNGMiaGMf6thNjxVx4
x9VahBmp3y0khlgdYGk3ngeTm04GCttKLhJN+Oh4w5chvsg65OJAcf5QFxdLat83
KEY83/QhE1BWzyyj8gQQo4xb4z2RHLvVBL1WBv4umUMenc/a0/qd4ukKgPxH8cI3
q2O/N5DaOpmznZkeuSMBANcnIGCw/x9V5b2MMLf6HjTAtanoi+XHAJFOwawMaelq
W9NwJq2EyS6Hvinx5/4m8g4IJspzUvx3HYYJfB/jvOMz2vp5icaUmR5EUfvnzHaC
pXK49wT9Jv8CPoEYkfxWOd3uOZYwyH6P3EhgL/P/8+hGZj3iN9mcEm/rWulBkuUT
nlb7bZPkzZT6JZqf7SHwud+lQOweAruY4nDvl1fU5NinT3KDXN8hWbgHXyYTMCIo
Y4ymPgxWsCSLn0TJBQDmJrfsyd0kOBySKZRogB46BnqL3oAPFieD2k+mVwsp0jAP
Hio0VzmxfdZvi2QbdsCYVY+NJJjbknOr4qMULeQLtQQlJQ/u0BkADZl/2kPeXknD
k01NYgwSbWO5Lzw7yiyMw+/UzrSQvNv1RstrL+OeMVRT3pd2xY5KCV4f/nY9xAoD
kFYG9yxKYIwkgj/BUhziP3mK50HWa/ooA8QEPun8DXpAfgYOGY7oiQl5QSNLxalP
Bx7tqqv4Cjor5CW3peqkcI4z4YqhILq/WTlJfmGnFrfRFIYXbIA/tbP4YSz7TUZ7
DNlEmD4dmqKhmFASrnqAow/yq5bWaj4ZMSuaqza8mwORGTuzSyoEKo11umjUbm6L
FBEyvGrNLALedKjc0GdpY6XIoPQMc/ggJnsrahjp9rwcIFFwsfgRu0Y2GRb0wuE9
Y1xoWyaXwAO1//wNCmEaWsrwAjER0kabl1CdilKgn8obyhhB8b3bClFr4GQ2EZ9z
c1DhN5Tima7w/ECpwSEc2zLu9qJce+BmeIgJjXlpJ+jflGgqn3bvk2lf0s0qnR/2
hnSC52pEwDfgVfie99zXedkCe5AWpJHyji/C5TPNWF9CVF4Kp1Qr57yPA8Fq165z
/kwcWih75FE6Pw0z8EGC6277gdHVSBlNYzaJ4DwFmkwzg+8ATC/iDlhjNCYwBdjA
zdDE07Ivg5mIxxI1UVmv1lGXMgArFF/t+JK3CZdxXAMrXz8fMfa4hRhTxVMRHSh2
pnmBytF8WpR4p6ReRTIZXKEN31pGtLbQXTPHPSmq4xtVI0aNUTH4Xl6kTIIRXNF3
8s6VV8lk2TbQB90BGpNA53qhUF2EuEFcHQ0O1nUCjeaiEA5lFCHyiMKhGEDJR4Hn
5Yk+H3Dmz6XlLNQL1mMaTkzKoTjO1BWr/fYvvuI+6bbScsKLTskI7vZjWD6eyhe9
2sQVobnp1ApmMsAW5+DhwBnuYrxlJKPn+Yzh7iUmQzqbxRCUi2s2dpMM8CUA5IuF
uUeKb87mk1BZRN7mk55C0X0gvQKleJsjsyjV7KZ8wZtGJboAe1OWAeWqV+Y8FpGb
6LVwAXKUj11SZjGLcocC4fYGlGtCw9fgK22u8vGzsJI/XSlLTHlooQXiPskPQ2TW
GwTx8fygcM8abglyJhEdSD98AR2svmcs7mwK8IzbNhDnB2RvvKF7TU/MvSQdCjjv
9qaFyDsnVxgbAHhr43ly/VsG03sPIoGshoQfpWq2jl5z4XPgaembHxhEpXYYMu8k
AJwry+v8f/J/XnnLUaCzFQ/2eU50mQeh3AmbZa1XzYtYUWSq3KiO1hmnAOhH5RMq
Yv2jLCmWJ7NSTvAGVteHu2w9KAtlKTOaKkfCyTy3C0PhFsXjRZjlHBV7RgsvN4gB
ItrUOTd13m4KfkBoZZFYyIctmQ0Blko89bdF+EFv3ckrHNNydn24i6+Zq9zhe+Kz
YumHsOY+7Q/GjATMZvfwafgRzUWOa6mDAJpeEq/iZS3SC+m5IAG5Nj7VgQ9TDsFC
dlEKRxRCJ08dVs9ZRN8piLsnSFCW/HEkjP2ZzO4U+F50Yx70qBCndP2oaFZVRz2T
krEgprAsAX8pwmew4Wvc8kVtR4xRhrpVpFvIpzaMSSHNDpwvPaJAIrbU6dQ3dSVy
IZG5oOZMBT/MXIXL/R7GWCU5XVecVUe+jgkyiKjWnZJ2p2aHdq2pEcjnoGwvYTYO
i9MgObatQblIpgc75C0Fdz/fFMWnRzqr00Lu+J5D/JqVeGpZq5H2RWBVlk9NLm/2
d1tWEJXKPrDuOL5MGMy54H1BGwb2aNj2clvRxvbHiue8XdhVrKokCHeano6ACHoz
zL5DFEX6oYt9sn5mxq5d4y4vG0wDYGGRoqw8hmSgn5P9I+5lolpnaN+o51xbAq/k
MIHESmqT7STubl7j6c9YgPPyvPpPb+XDEC2+7fs6lMpVX7he7hcmM0zX3Zy3+tas
53VINUBvgnF15l+a2Y6ThKptlICzQI7uB0ij2SXtDJxdCj9UaumBJUSkyuYW5fnK
K34x+ZRn1x+7TlNefXwFf7RhzSeum2Gd7TSwLKvki3ZNHqyUblb+kIIvKdH1uWlW
rsAe/nLC1dLlfbd1PjUjTRNuIwAtPmTW+jVYkOnuydHujJp5KIGZYLI+F3QzSMtL
6CHuFLkN97AWB39T6b4ZU8Uhw6x0CH26+kDaqV5/ZqNbLeFq5iFb7gSbGMBddhA1
hEd7VrJKG3nRYAvLExNFnL443Xu9e31QkeOU2efODojldvqoa260FMkZX1o620f8
y8vl30u0Kk2HKQeADPX++F7WothMeGiBeIKgSbNbf/7nx7twwUN7Rx0gHhydvavT
xAEm+AjAbmtDAZ/2+/GyU74KZrc1TBIgidtEY4ZESlrbkfbk0H8vBe/nFAIS6jft
n/mD0oDVjgsMQ4/BxzQsnCR5hY7UsYZx3JAFrlkjao1IOaDQlFbIm5hPwZL43SQD
FjxHrM42mDjb/ujGjCirUe51lgseNtT1F/wz2fWLgqo2fcyWqxWiF1s+j8HBnx8Q
EqJhQc/xzAEAUt3I1ml+9zzs6EqRVUQNM5YQowmqddnHAQyj55jZwkY2PgBdbjOE
WlO5oGxo57BuqqRx6zXbZ7bxmWYId7Iugnb0ii4UqZKBc/juBBcmTg5MBPnN+4U9
+rRhWfNsFfjYAZID/GJWUV33U2LuFeVkmaFI7F5iRgL3JmxHRiTUWzxjKoJR33HJ
29V1Osf2nVDQ7dykRdj3bpDg9UrsePcTUnm3EvVLDIBamTvUuWWy/tvnp19TCeoS
aVIqdVyIr7vIo2zh615ZYCjXwIu/loFaGs6khrDyfugCrZEjVmWExsfwKpjUdQWF
LHN0l30BBrXUxYtfHMgvMzMiTU0HNmy5wWSB5ztFMAsjMbgYg2lqvDgFgcsYgosK
5EH96d5F6xO0sm6DgE+IAfVjOvTiDy17Z2Hn5zpRBGKnLnjxrrf1qcEafK+/eYz1
PkkQvLRoB91w7GEQVmMu+IMIlPDQ9xcUhslhsOhbwPH7UXpKtVC9S9KTMtLuh4IM
sSbKz6/0YX7tv3H/V6EcUCvqtM1ENu6Mge6sa8g5jihAh+HrnoAC1wJBEZy5xAHw
tiDGKrHvBPAMfvr8oKOALt/TY+2OC4VCwCyzCO9erHvulpJ78BFVrKzCC8gmBL6B
qraLf5u5Fau3KhTlWPJTz8+IBulqtwc8tHmQXqPYDVYdx7+xFJtpQ/TamWDtij+/
RUKOpEKskfYwfODYj15BvZMwAChY/E+8aST065C8bDx4EQlqLbm4bONc0cbzKAyO
QObIyc2+EaXKc3NnPEIyBM94aNdenLXbi/KapnmUbYP12ifPEDjSUQt6P34tdkwN
eHjPyqXemmvL+F9jj1okPrRSnF064VwZta1uRqRdbPXBy076Mtb39DkX2xGOueaT
HDvXXzHgC80tFiy8B+91AgHK3v2SDeta9jMw10LUxxqKgTBVfPvEm1uSFgjZ40uC
N3f70cU/banAIw068M7lxeP0cNAHrTF7a6RZSnwavOEcuQ/H7KWQMETvdHC4lQDp
5MQhjr9S2pFRx9Tvwe8Y5VNi+c+3YJ81MME9c0ryKFJHUQyDWGzvWYEZJPk7kMbe
5sJwSmc81bKkByTD1wepUB+/DlykKvrwC0a6tSCkTRr8kJ2Uzzrb0149OstAEMOm
tgKunJkqIUaXozReqMxzV7cgoac9ALgBzG5tiDdWh5F6tLfJgFcf9/N8pWB7mb3O
senwnUu0/7XwIJXoxZYrUWrKdb4heXzUlzVaE07ZDJOB2LMPDJ0fTmZ/NREn3wMx
m89lssG2Vm2PHoJ54PYoS7MsvC6RX9/8TTCRIHN1+xWkdoRyvOgNuO9lEjl7edz9
BdhoxxsrmUPHQ2F047FqluI4D53CmoCxpQor79CTprbxI+9MpA2oTAR431SlaBBd
KbB6jbTNpVfsdr4GueuTEbnYTUVoxSyYM0shpppToqKEGA6/0WgkbzIS2cwfwcDU
HCh22FZ8/bV06ZASJ3Z1zsG0Ho1/CMdQd9j9q+47EXvl1S2bzx1yp/rOUKdRLCMJ
DK+8ItXCGTxjxTpMY2cN7Zh/hfPF7PGf5txDP3k36tyHg6z+TtXIG05S2ys85IFo
CgzKYddxzON3az+IjPr5bSkT1rkbF7s1dQUArOw0YWDodiUDYCWIXwHgknzxLWLm
N3rnLsh9fmJOLIGQN3/JtwwjQO/uYTU1yIKSzIMya/wlQrYalUwd1IGv4yjHhQEq
zAZw41jQWgOQHBXzgK2QTPpvJe7JAB7hj2vXZALrpjxNxd/oYP6OVSM6jKbILsx0
MakRRZ7V4okgG5oijbACgwWX+t3iY+XyNp2XENXEMOpBISCtb84hDFh4vfzmb+se
/lKHBXHpxMmeTk5tEFdIxbCHlXINSKW4uEvih0rMTXeRJo2faiAyOR6tKWNP1Hqg
srA/KOdKwPtNQGwK9XA+DKP93kNOeI5cTC/wEHd8A8R2t1AU9uhljOIym9pIjMWv
+pPuHnbUesj+RaKv4LoRB38qM7DQjkVnt0umcWLrPNitDIul56nUR80wzhBjLJcC
/BLazyEQh2gXfkfcBLLE0lM17iM1ruJe7gY5rS2fBD0jBoFFBvmIKM4yxYxl1DCG
Cx+3PvhpBUXofbKWbPWJauR7SAMtXO6ciW1hgazOq5Ie+J65eAYks1TEthgeUpR8
dNWkrnSn6pYjTKURLDTXMI9L/e1EJQ546I5e91MEl1UKCLcxWJSUMQIgteh/IdCE
2Mxfjxyd0UrQHEOKSdULPbW5d/GfxAE+scrpKpg0OaMn72Pjhy3oAls4ynabOcWW
hTYAINc1ycARv2OBRBY86cgNoss9nZdSslW8VGo20cIeU3+rs4l2/gh+bzZl5Vam
GZHWrVStuLOx05HcBJrb0hL/EgJDZeMDsr5UtYTv3n5WtEqm8NnI3WqaILzBXRKZ
jI6IZbM3n5ZR8zKQTqEcRx0C8tiaxE5kmDvdCpXGqtOK9N47fzZKOWfkLD6gHnOq
15lfsyO57GXg1hPL4CTD41KmZ9ZD+mCO813AJ6y/k9o1KyiBh8ocxXVeJGueus97
vxh1qbg/8cypyJ7xmUuuWL+17OzATr55dPDGvvDvxzG4Om4As5tblHbSeExPJcYl
/2UReS9sGLmUhYXn58rMaZLiqmIII9V2gjk0z4U1Nwak6iNcEMaJhykdC5yUvSMS
wg9ml8drHzLyrJYb7wvLSyVeNTFaTb9NozgTvJWRki2yaPMunCbzbQcs4O+llPp5
mrsZVZpxsoQYqw2x7AwQFQjoAzkmPlXbjJKKJ4VXcty7yaFXXazTlHoLz7u9dQs7
dDQKU1jCvLForVGGBE+/06HULPeg5lYNoRI1HfL9ZMrurfEXymXV1BiaJFgSIh0n
r6+DDgBS33pYb3UFrcv2cc3hYSh3yKrLZ8MWFK5tlGwZn8QBagD+MA/ams2QPxVk
P4fT20j4SYujV9wP8iETSN4mMiucvUt+NBnYgyEVR0u1JY+LLAAmWxCEhveCL6QR
JsZK0mWuLHsyR2j3Kn4LTtFPsS5CX9FS7zhV/67ktqcV81zKaHM+eIgnHLIhl7y1
vwkw2hoHDNRcRc43T1GbBV387cl6LWdkFxX8n0KsPWwP3LF3lETFLFd0zYJsnTN/
qyyCy4u3+uqL4cDCx4IVv6cbWu9jheKRL7/p6tlFZOmx40pt38fkCLtX3aRc1uDq
3tcJlVlA+hRpF/WcLkfV8AFy9xHJiS4Rm7Q65sswE1rfAMT83e5f2LUBbn2Lt/zk
jP/DIB+BJd9/zDlRgT/4U3bXrjNLgr8yayBSAYFkVeac80aPE20sdpbFN4mf6+kr
m4ve0h41/bUmxOngrJo/DollE7d5k2COoUeDlIT931gR/QOFTqq+vecEJh179I6Q
S3t3yhOsl8Q5w2jwKrguKvg0fqrGGrLiR1aZAssYU//KvnPDQMEANA3nCdSSC3q2
33mzT3gGhbzCK2XcEYbAJtUichgD8UsfkBZFrxFl0SpVY0LzgdSieV/1M+KHRF7L
C6osyIf2EKBAEBbSqc5Hjrwzn3ITE7UmV/bBtkUDn2mb9YT9DdE3kxLINoaNG57o
OFDTjInKF1myRtYwVBcAujW4DeSwUe+EeeU0yA1mnGXUCkAKp9q/KuwM2vctBnft
sPHkZYNHHzmZBv5H535VkllDJSP+Pt+ZpbKiYzxBgVxeMmd/XBX/GLMlHFQ2dP94
GUrI1rkTuIu0hZ1hLcrpcWbboWVZPz0mJhl9mO3swlWmSuV4Yadz9Jib1Zf9s51y
59P/kvvK82f6kOgkG+DukT5S+mzQvRXoO75EtFVoFFdj+t/fZXSBh1Ca6wqpj7MP
oMzum8wBCIYdPuLbxuwu92EC/pQ3Of6z4SltoFkgs8vr9B1tqqhmnaOGm9pm0nm3
r3kOWxUmL/dWEbqAGtV4fT6xmFynoVjIcUilM1tzJ4eFm/xYNTw86jG/QvGuNG7j
tOjTOvs+MGC6ovT5EwEGvAV1Zx1Mpw1MXK8HnCHCQvf+1ri8MhQZtzgm2YquqIRl
gu10B0G2XYkmRY7Za141A3rrZkftxPeM6ktRVIABSxBvK0W5c/3xafU89l9/Fxi7
XTm4zlRxkQQxRNsi9elRp+GD90+jlhllogw80OaFP/kISy+CRyyeBvrYE0b/KqhA
ZvEdSP9zoZBHTdsgxj2+S+DOi4UrkdfhFNkZdQQ0N99EHedCmFFzmIzZajgrOZ2V
EEGCtlYX8pi6y3wEmyaNQ8Zh4AbTkLsl1nidh8/9eEibXow2SgXjXQGUnNDAPjuB
siyNoJ2DzvQqaFy7NSIW4BVuHZuWELl43WInflH7fR8wRiTkkYC9RrU06Y+qPqEl
WP6csYxUmVkepRwbydOJNN/jH2XsIclaz/QDiW+4wvV9RFKe2KwpacZS2LXBCGtC
I5eHApnA2LGW6AjDz3+uinf+bdj2Rgeqx86NbMh4MEsi+lGL6B1FTUuDKS3PR3pt
CE53b/3Y8EQs2HgHDeDAPUXOEiO56pYZQgsJlMiC9tFLYQC0Of1fVq0Ejjr4zAbN
rVQxIWfWZ2eVZVtQWJvbgpkx4QUdzwW38sn5VNEF9F6vA7CvBD63/G2cwpadxOFZ
0qG+5XIKXfiYTaE8h6vbPOHpVJXBviNkiAjon+cUcwUbGUkNiURN6KjIsx5EOSoq
72zh/G0imE0VW741kQfo3tCvfvppKhHHe8CLH8ufrttwAZA9R7nNrk0GBodAnRnL
TQ96L19LzuasYiPGUnllkY/F1+HJmXvcXeRAOOdxPRPMCcmA7mUgKMn6zt+mYoei
UlhoeXypuWOfwPA0XPw25uuBkr+4K0ojHWuYSUVLCJVeCCFXBvUsSTuC/jlJDgpB
D51jp/St08br4zxirb+GHgJyBw5W4JkSzvWCeHs66lhW0YGGDX663CdozMMvMLYt
0eqH7HxgXGzGPIbhmCIU6QrQDFUrb/f8NO9w9RFnO1V98HfJQ8UXTtocnKQH05ez
jGI3jAoWJWCh9y2DbLywXxAAqayX7iGklLFEmhDKl3cHXaL22my9qGqugvcMlfgI
QJ0TcF8dBUPCNPpEeXK3karh7dMavqbv5vkWI5S/M63NlH24z95GZz8scpw60kR1
XYapTAV5WHFVapagleFa21cG8Rh2Xhgyjxqa8TjjJzPiREM3CuR8nKw52QWmVBBR
XJu2KWZrKVPCB0EiC/dBKzYAe3QxE2+FftL7xQvHBClJ9nkc6uHs8GeMUeavyLm7
WL8m+UzVVhidWE7c+rbwTzM2uJ+uznSDGCu5w5VyV+Eq5yEfsZDObVJV3RoF7R7y
SSeC7RhT/FDSFVDZLOP80xtSbDTpZLPmo5HDYGruqAvHzFsOx85IYZmmCL94eD+d
2qms3KYxJ19sSRUTIl0dYnIOLsQK7idXz/65QqFf1XrHSkVgLjcHbkrOj72Wg4bF
v6Q98KFuoxMhc2WDiopf4UaNASf3uILCrG44r/Gk1NerhfAvexWxNurlKsRW8oeG
puIDMguESbqlaedb37XJYgA2qvnhAf87eflrnKKHVi3UK937s5OyBeIbw/7jeUwU
hgs2HepJuXvOWVKy+Uoc3VUOufMGin6+pN6ESKlSnV3eeyYU8NzXUQZSf0lM69Ea
v5BWba5DtHytdl57o8hC7ctwpG+qcm7QZuyQ5+1eH9zTdx1aXDsnyLaa94BZNJpq
zwMtdKWhq4bRguyJxsIHnsVq+Wbz4OTRDjCVueXWT5Gwf/0EjGjJm+NC6H/0RW6D
mcziXOJqKiJTTJuaEMKg6ZCyYWCQbswESMnMAQNuPEktPxYZ4yIZY8R4FWe5f+hz
+OT9pB9EXXWh76i8DjzkdZLSz3bJeK4yc58JWuBiyIuFtr+L3BXL4Ov01C4aBuvP
/WAT1Uv+cKERZ1dpWNuDJ7r6SUbaJiSoP/fCEHYRiTHg19FLCFJFeZYzvFrZXli0
7I7TqRtCw3WdLM555abMTeYhHlTLU3aIZUmemHLKkquyE1b1IiRMJuoOVfsPhGYB
yd3Y0sVyElB2vpYxkdORsFToNB8eJaf+SC+PX3nMpyAULKEc5agTaxCdbAvIg3RK
53pVigx/P0xwZP9qVZ7lKS5j4epj4t479HgkLs+OMPEzcySurYztBkHTbNvnP+92
4mypUn64gqknRfi8CsRdRO65EDBVMUdA4Aeyg0aB71aTbGUzyyx+265yK+Tglvat
RkUgHvawxkUFjZyGzFANrwKahQd1H8g5f9cJjXg9RI5JqqPLMiRp4giv8bk02hhf
D6mPSvS0G8JL3wW6K/yt3XSelOhQnIKTrtQaavEikv6uL1J0hTWg356qUaJeKKs/
HyQ1kDhlxdgEJx3yQfzxckePAyuWkYQM2Q8Opl82cf9TqDXRY0/i8n/X1Zo9danT
bwiUkevkSlMoHV6FoCQpZeedsDa7IVrSXE96LBT5gcsz2KMs5qX2r7HrIApL43o+
0qtD1VRtCFT91aIHoaHxlnOVSDjQoOnKnih7TF9HjIP7jz9SWMIoFf0buX7WA81B
fy8QSyxYsXYQDziaWb1Vd1TdtADLftWq17MFBAw9U3yzTcCTpKe45tos8OdvAr9L
MIxg6XACa6CcOk2xtJIg+wQBVl2vxbFIZhp716dbUhuSqpEPWecmi475DNQRjI9B
jjt2b0ScXkxkNGLoGKZaMOYWQ/AJpIcDQOswdWJWgsN/jlggUws4Fm1MQIu4xfGQ
i8n1GQIDbz3t/ifsScap4SfbcebNS/UEy1pYzGLRQUBDlNd2YmMw0xDP/SJRStx/
jqaPbdcBWNVQ55pGtZw4d2XueOwl6BUZB48APJyNlKt2yWLkFP1vsCNwojE9B7il
pVp+vwoptGhAdlfSdcfqSkvtUDbuzM9WTX83TNd0qvo8LV6TQ35Mg3clWpF6eYDt
5apM8QadBaGNcuWau+Arm9DMPvcrVdTU3/7k5U0qTpc6KNGX0klZ+HBnN1IXZykT
fJROoIs07GsrkFcr3631kcwCxTvZB5u5bqixYOHB7nFGXg8z8HwFZdxVafcfTHcI
LZeiPeEBN3u+b0m1AYJ+aZ0MLh3IQUkjeJA0vMFkMFAKeLoUD89WJMqU5SkqqsUB
MHp04d0aqpNBw8ZcgT9+ZHhs3npzQq/W4qaRmp0mEMsIDoTcnyBhNSOAKy/7sGnM
AiG37Ddczt4KerLX9K0usuv3NsV+yTPxNqeVUciVTcT2NuOtX23dg0nrbZbiVmAn
/P5BKODs6QZdk0WN7D/TwdVRpRS557/gOyqbU26pSQNZCxmSAVBaRTH+nAoYg2KO
ZW9V/54pi7mHajfMl6AsXVlP52FyqG+elDszG6GsDg+uQuAa67r7KXlFNQ58KHoZ
nIm8NfPzWoH1imTRLcexoYYDuNQo2j5A8cqmXOSCoAgNl3W02B5skJLpwoC3rgC7
utbvtgAYc1v9EjKvpt6fTqtj83m2CV+DCxCqVHEgd+km2gp78iZNNZwT7tq4j2BN
h5BdOUJIBOjCBwFuOrBeUigaci12fachrz8egd7WARBvvQcR733qhbVUGKbEqc+3
Znc5Z014lKmak9Q2/dXJPo7e3dRZ6VdzXMHWD3EHiFOyytZAfEGet7E+1eU/AiTt
8Jw7NMxnDkXyvIhRTv6Qgkw6Y9cx9W+NuCKpVKGtfbc7HowfXOo9TdEPr81bjCaF
mlPNqkHUl7/pcFf+BTow6G8pi0vzKZn3qvHvbk7mCbdL64YQ8CTlla1OYUDN3iEq
XPPiw/Y7AN10sU/vvJzfyN6ebTbqw6Gd5UGvznSYPQ4nikngzZs1RJj3dBXu53w3
zkouOszlC3uOD26B1erj5MI0ZgJMRSEGnW4Y1g3tYliRdYNQzaciqpE+ov2cO9A4
ESqxZZgG7mZOxdlUdSGPYagN7RGCuCK47aXQJkCUEMFAzsArgUH3i8oGh3kRhTUI
LUUkTSYk5xZRU3jLnDwn0oE8HEtPKBRa1pfZ9S70jgNiLpcayoGExnk6QHdaxLpk
ap6C7PaJMlev+1SUQQuUktqCnneHXvfulKW+0H+uU2y6dnZ+dD181nGfVj0AVlmN
NcHmXV727P9v37J7vJrMHr3UeSZA2I7oXhnKx6Ur49k5rE6MyJsNh/q9PacQH0wf
JxO9GZpQvdTBODG9U5RTOjnPNnahcIQf01JxZ78dnpb2JGe4LzU4yICjEVhi7cTu
N7CTght5L3l52771BL9e6gviUlJs9jvu0FgtxabZOv3EJci6G+DpfEhdzCEUZXe8
zL9RfjmO+VbNdcOovsk5roDht3cPn16HdLO/MzeG3jkaHPO6y6oY8klnAqUu5MAr
PWhpbDhi4YEiHCaCuf2QhPX4LTWkZrVb7Dfw+D2zNAYapjv8SWO6JBRT4t1LHbC4
LYf6A81ZOjD7jsdT4lZx31LaGMwUDZq658ncpDWFoCs+QbBjDTh+UmyGqEjHpCsp
8tZzKbjJY1n1jsj1+MQLl/MOqtKJ/H+IzaDJ2XfnwtxUvefw1Kob/42bgoEJvN8z
aM7/fmu9eofoU2iOIs/dOPzqokvJw8pvTxfh7bO4PKxmEiy4AOCZNYgo1YdHhydj
tLBXrui0C/3LDj66D9XJHhPuaI0ndBSVO74NpRr1YXIUIlPsg5DvXg5IfkZxuA7l
gkNZhVMQ0xxWXy7OtilRxuGHj1gAhJ6/WDIwcdxJCfIpS83BeQQ/3TppTVLvQK6l
TFJDZJZK4yBcIF4Z4smBBB/kRuGdNjqtdq5dTWHzQ2ib0oF7FneGIh1Mz4Kju0QD
OVWkQlRdtrOmBdZNfeSpvC2lZofRe/S0WhSn801oB3C9wIk8GqJFkmzP/G6Baf8E
Tkf/q25xMaRlwIhb/Jt1Kf2qAqi48Ypz4FLci/qFGbm9WsUq8Bi5swZ6By2caz5R
FQHgty4gL5Ym4CRpJRbdLOmZ9OR93mqJ2DlgI/mMjdmvHrqyC/YZShxQYBwRpj6n
jz9tCP+QR1N5NDAQnNYn6rtInFKL/4h3t45WKZUMVFliZG02ohXEa7SoUMiA1uLm
GGMQ6iflg0+gJtuYHQZeq+Hbz6rxRgO2FKe45wz2cjBZ5PnaVPVMLKIn3EdHr4NN
IzZlMUE0Itjrmn7MgN0ecuXC/ZI4quZA+Y72i+2x0iovYn0boHm0ztN1OTQZ69hB
htZM76O8PYNVBZv00ped7FH74KT8W8qu1ghgfrhFVQmlJQ7c66TNlQkthm6Np+XW
3m7PhiiuUOaltXHCa21nXSI6IlD0+myeU+1b3jjtpNElFVk1w5SyNWpr66+QG8NN
vJJwO/H3XXMfSB0E9eh2UjoNvrY1TDDQ55p2/qAgC1p2ra/yUour1TS58oSr3DA6
zssxXWOLM9sxI+gXFOpufbc5khlcw4V0BdqA48rwuBRapL9JhcfnV5FmAmbDoDxX
3sillK1fk5bVLPIT1w/o2tD3XEomhHyZXM1+rfljYW/DAq9mO39mZHuaT5FjJE52
TSKnw9sl0o9SeJ2lQrC3LJlbox3y4sag9GOAkl59goJpan1x1rFV0EnP6R9bDVIC
qsLuAOIKw5Il3XqBnaox1mVmNkAjVbAXlz83mpajMJNoLvKaTd+w9b46apUyTm8f
jTSHwyY8kiW/52hbMBv4xy0W7kaFaZgccdlvVGYNWcTdJBYoW4akcuW0cdeNwqC5
1w3+1rGdiPyumyUBo7rq87xhpmQElt63L3Km1oxT6gFOYwq7uDGc1KBw/rXQpN9W
18G7ZEULm/032lkKDypvztkYVqe6NNPj0q715OWNvGeNuyPa04mSMRi8SSjqqZQW
+aqzM7MesRnXDoEM/7uqEKedRNRid/y0TlKYZTXQrdO9YurNGQpnOKUZGV1PVNI+
ocvUVefa4fAjDVQkYw3jNm0740h3AnkVVGKhlLBfpux12uV+fN8XDNbilRHVNnRz
cLW8Bzv7gE3Qna3J8tSx2eZWWkXUHD4BdgZyMix1Nt9OcEM2qUYwwuaeFCgN3EgN
bWS4AC9dJe5cT5UlTIS1a7J5YZJV7ldI3+DwYJsMcfX8bDrwVvTENisnVeWOmCWt
vPa868p3u5AkGzRyRWK6qpcv+IlMkdohQY2jgyJM4TLYCPs+ne3OWL72NLW0RKLa
BK5H2wQI80qFXpiZn7pn3M4/FZyvL6NPaLaOUquQF5zYKDxksy5yvXIsDoFAZeQi
EDoe6keq6kpIyPzkxqy42uymOag0pJOeXVAB6odzGQtiWuBzpM3bPWLr9eI9u2Y7
ud/F39MyIgwweV+K2L7kjWKJ6GeDn1AdppKNVN7EICEvgXc9bJoGE2sYnmiWs+FF
ZPGrF2BVM36Wojd/4Y4vlXvTsfii7yWmjqF1uM26zvxc9RuAsFjEBnSOMQyfYl9f
AlKAoziFXao7CuFX1uv4SxVDdACci4b0CUISk7aknLhoT2BzE/AtCle0NhRGiw9J
5dvGOCrY6hm+Gy6zWm9yG2h2+ixJ0IlmaXMJMOEUXjhA9VF6fd4Xqq1FN4hQUAO4
MoQBOh6xKkh1kjur2EjlzICRBpV50CNaBfSFmW/leLW1ZCqB3uUuRnpJw8vvCIuh
wRw2nvZ1iVcvXkWlwSZwfrPe9iHJzSFleHRentj+m6wscIRwF3osYfvm8GOw6sdO
y98j2CxQq3eYmfgTa1Eq+KHcFEARgjN1BLxWI2SXoJUjGR3at/F+oKd4Blz3fKfG
xue4R0/PFNM+DGECcZoZuCOrVeRVf03Y0s3FNRpzJH0Jycbun3V47TbrZQq/O/fd
mhex6r1ub39oKeGGsCD7jr0Es0KDDd4GUKnRU4wAc/0EH9mVX+O7eMlSpTwaRwi6
wsjfjLaNDKiIPX9ZufF5ho489DEVUPD8lNJwmxIPlYxwk4ixAArpEfy3FzsSrBjS
7grE+ISSz8nFFo4IB6snXnwzZfIli8E4LxCktM9a/UWfb4Kp1sKM1BrL2TSIa6Fi
OY+m9xZbS6MImJaeFaeea85reT1vEP4jry7g7PV+L4tGie7bvS80Q1AqdGD1mTh4
S69X5ojj0onq30jaB61rZSJarg5SOfaH3uQwitFuf8uKFioRNWIg5BuuONwp4fvp
Af/H0U4/M5MNLPOjIB/TObBkVhmvimOzePa84PuCbQwcmyomEhWEXVNwv8w0xDwf
6ZXn38PWm29zTlFc12grdZ7UcmkBIWfGJLpN6c9pqNjZOP3GJ6+Fh8l69yv7WdHY
FSXQ4FUgwvJKd900IkcHJ+X2bCsWCwvWq5rC0HOY/YSLc+m1yLmiGj3hvitnfoj3
N7FlXpCPI3VW8717LfhV+cL2gerLT35DR0e+Pq5nHGM5vzO+eKG3xEETLVoYTGLk
CN9a8Pe7hUZ1Q5LBQfFX2W+T5+oI9fJ7BRmTA60DzZyAV6Whfuiezxk/JqOrNLeI
oR0Urtrm8Dje96PeVbLGYGEgQ+btSCPBX2b1YL1cc8loswmm1QF5UdVH34GHunfn
t8UjvyEjg8XA/PvPJgiTpuYSuFrGIsAWFgweqnywe7FmLKcwtCwiB5WWwtMKNyyZ
4o9g5VSBmQJW0bkoMPw8+JEAt/tUL6BcDuYCSCIRZ1mOJpsn+PrfZw0DCAEEkcpz
9mKXkpml5MvNIBXyzah0JrbfLPmKxUtXzXjdd98nfoTNI5RWd6flfXDOAQ1sKZqM
XGtrWDMEcZq4HTl0IKlho7fRKmow1jEK/bzIGr9/zTxd0u3AL6EwO3vCmTITCz9M
QgJpniSgEH4X1nAs4JI7xIP9lbuqY7l5V7KGAAsBsJIlpNC84f/6llb/jiBg1H58
MoSZ1T8WnQWXYbHWuMNOFcJe3OTZ/GjRvmnBIamOz9W3OJBobxPCUq4mWrKyUkH9
bFZJ9MhzwWBUCbazgLe74SipLWdvmiWKo4llKVOWvnOKQZvIzGNGfzOZc+uuYPEG
blY+mG56Tgg42KhCdrYigfnL0R0fcVbSw7iyPbWsySr8WDxpdF35R+7aCkH+JJS4
GKOFIVr8loGCWPdNC1uPbmx+jI9dSLrzHtHAun7SZVPOfsUssuWFEKHDcBKL6N0J
/SOvSL7SCYD8j2u72EkoIbDKug5aJoAA6EoBorDINQVmMtWInXMJn7Cu5ltbp1jm
CUTIAyk9C3QyoxgFsLVu+pvW00NDTk0cZ7I2YK8JtwfDSGBVnPBk5j4sgt/vt72/
K9LPNtiy10FRQBJSMHOMev08JI3aS/hpO9AV54Sd5uk6i+0KdMfmPRJRl2wXiQPg
5wcNoBh3PhQ3Vt8f7TYoNUuvV4OfWWMHUoV2rFo7hdyUb+4m4iqYqYsL52+2FOWO
9MLAehUvLMfloIrbhOFRw/dMHqkbcCWSdAzOUsluEYMTKt+F3IbkR8vuFRe8YihV
LOp547f7KUWPMu2zYT1ukcDeb5tey4oeElBzBia6SjU8GWQn3fltD0OWgzChwLgB
b1wPTzn+CgbQUVjd7E8j9XtLW8JolE964VAq6FOluM7REcBnSxsO66CYyayj+yhf
u275ScBzxZp8sYClZ9ysL6Ij3OoH1qme0gAWzGMXlfxAlAvdQ7aesBGMjiNJLaq7
GFyckUe2DkdnsxYWIW5CRB2A8hczxbrL3G4f0YHP86fz73jLCGPqS2YlUcoLNzXl
439bRKhMgGVG0KQ5ZjBpEylBnN1o4uIIHJwsTth7vBa9vMX+e3sfrSuI07sx4qkt
bTaWNvxXDfu1JfQa60zez9UkbBIyUb7SRFwpx2aH7DPxxeahp0dsF37ncKd/q7Kc
B2eCFVQ51+qaGJ38EJLrjscvT++FgWibfo84M8+KmuXA26a3ZU4/PXwBvfDH2jDs
7KWWx/NRTQ0tMKRTF+9mlCeZjGRQVtNl03wbeGJnQrb7H+dhZjT0Ua2WIUNOhAPM
M7CoO9fsKkiRQD74NM2Va/ibgaKjsA7rJUV23X56rFWLZDOY4llGCgAQITPV7Ilj
+X0MJqQ0LU4hHUSsqIGVnPDc8ILYkQFi+U26y0Ozo6jqc38zzbhy0yA/xihxS9K3
+5519IDQb7ZVKBL0w+UpwtUPGXQIW5rl8FJsmaY/kxwxVfGEIKKNuGjV1diOL3mO
dsHyjosETuPJ7GZU5x6CXQ4yqPjw1Sx27K941u/VPCKbpdQFASG7d4QcQ4y9E4UY
Y+5ZeLLUHG1I0c4UACuuJ15oSa+C4As6qfwPc3Idz4angekDQfI0nLe8LsBO1KcK
mBe32TIHkcqp9mYA2HzXVRj60ufoB1dJX1BMyDBEeFWnpp23Jtzd880M84cy2dli
QWA12BciKNaVYvFpuXyg4Wq+AvnHVBodhwGcPS7CXimWMMfCCkOy+Pju+1MDzCGm
M5Cv3w1xZeRQbabjXkxMoTtjnZeG0bqKR5/zw03U9HoHjTPLmnoPHmfo43i3/IEn
g1FRgIOYrpfK2SwngxexejDcV6eqPxFN39gEzLGzQOTn/43bagtTVHkmIRyKKm25
n7g2lRunVUTUT/khUhToLCRADA8ypZaL6lw3JdWa+c21cOObGnjDnrCbdSCK6Ysw
Q0aYchd2zmbsLCY3/AFz989/QGVHMW3SPYvxdD6w3DORdcKTOrIE2WCV0bnLeawm
UvEpexCdyqrhjoXm8p/yt9LfeRgDhVEkYY0MleXyCeAGWKsiPMJdfqqMXEs9Op9X
DWH0i9mMzLa09JD2BD/NGuMKTiw4uRdYLGNxWarh4Adq1z6bEfgG9MOUPRGzziAi
fjIZiwkMlb84Bn2h0dCTF93meSSDKM43f5Hcbmqz9kb6I9XC5X9FiDGLov8LCHVA
56is2TzxLH7e/iVV+CgTdLmIk3rtRrniMBpWmT9p92+SooAkfkLi5hlVa3EFuXsR
O/mADaGKnm4xViuoviH7NVNgQ2Ni6SnBHBedTExCz2BYrz5xRleEizlECzN1sPNM
Oi2HxOyvUfnTerDXOPK2JV+KDxhM7yWym8FYACbjFvt1BGnrvhQAzzsGa3wt7iCj
dyUPV/qSr4UtsGJfbClyAkLtgftFTvDOTvp8oO1NjChnt47kpJuKgGEv3SUI3Q3M
HIuJsHplSWrtfQK+g+i25fhcp3JLsF9zrc5GnutYY8zOdwrDixOICB+9j49UCZZ7
caBlel2gatk61oYax6BUxJvDmoN/eErJje+G8VCzRjZvj94efVj02Hnk7mAXrcXl
axGnO8RHGAjA7HttW6pKgjUMSfctu/uz7p2GKOSkyMDMJjLO+JmQ10LV/1ef6b7i
p+A3s686gsxs0qK/xvE2uUDFsg4l5+O1ZvfG58AWQ0nQoBbfOPo0EY0fBQQTGa/e
xFnSsXRCa6nALbxuHR42M1S1lrfxn2vQX4BIjZsqAds2PqGkOJODgfQ54lDjbWZL
Qw/M4EMH5UQdWPqE7I2BaXbfRf74q4tQ9XjhW/XcLZfaPwjNAtse874pWtSX2Eah
5r03rQWf2cpEyAzyFqVsSvivcPrPcufammctbqlcpcSmTXcZ7sOZ84GGtjBMxcfI
YbDs+3yB4e/5V7UizLwAoduoLF50Lr9mPBJzXe7/dpjt/ExJJ+9r7Fb8eAzvHExZ
XQRB5CZKhyUaeipdEWv4OprAX00VEkrXb9p+NqkVLJ5wANcSwqSb4MwbzZ+8rX1W
UNsjyQPg1EnqW2Lltk/vQJeQA1SP8CcggSnn3Ft0AvI2AErLmzDiQ6B38D+w1LuU
pJewGM89jI7lkkQ3jWHmN8K/A/C4SX/Jj2/E1Kwp1E/EbXi6YYruZ+CUZZLXwA+a
86d/T6N0w9zethZ5Q4HnQz2rNgDvL66UTmcyShDC+JM2Iunra6d2eyDVf+r0CVpS
UUMY6uKBtgOaC5rG+4IN0QUT7RTZYpGMAA8AxSqu9c8VUDp6nf770sNZ5xbNfGFt
XJYptLlTENaflFJtQB7vudtooe6Z+6WOQFN0qrOlff9I8cIj7FtT0peBplb/Q19U
MAq7CK10g2FDKjKNaQQSaaNitp0DIAvaealRLqJ3s4J7LWSUbzMS41gIfX01KwB4
Al6y1K66MG4rrUrIxTdWkvNKGyePhCjXOPOaPogWYWqm0iVEbFNpX+yzDMyk/cbN
tWO/UggX0YfUeSkyrBh9j4lM/iN/8qaYw7idrI6Nrhw1jAjZsYg8d322Um3Vxm1/
knGLKWOpm+G5b8XWQ4CPn/oEtw/W7zq3ReBOfI55zDtnSpCaDbA5nbxza9SkyRw7
MvOgRHoOxoPz4mlFkzOuqqpVqMbdoW0hzWQx4CntRcNNSSbErrK+7/od6Fyzhrlt
UlUFXITp0ffU9v+mXj8sNb3qaCdLEXH3uja/Cn8QyBgCNowfJ/eyGcYzI2O56Oed
2nIUUuNCxJA9z0f23ZQg4WHpxRuwbIb9Ty+6p3UjLRNdW7Jk4t2yjAikU/2Kjdwt
PgV8fYcu12G2d2S2mx6E+NK5p7fUrORXHsA+gsOp1J1znD7XWTyWGwVKuJ+O6PC+
FIZF5EOHfVIXFKQ6N8k7WY5YyuBmjqz3+RCuZA80WL8e1YkdGrK58+KhkOoqE0uu
KZMHae01Tu793y9sXgqvyAeQxe1JEQIl3CQWDvZn8ni99/3xcnOC5H3wJLqKVN+m
QCjvE2EwOBvA5sr1cApxyHc56gqOzs0HCNs/Rc6py5o36qmiMlL7TW+PsrGycx1v
eTKIYhYQC1126YZIQvVQPOZkl0kfc+R+smSxKLbyRNATDMuTL++BAL11cyE3m2y+
chcG3VqDmPH3GrSJU11rgjtqypibNK95I5jMzVheRGBPwXwJBng034B/chlzWwue
o46NJBvpkGJOvubg++kQTahKRC+upIJr0NTY4SOVV6qJHVyn3K464RxabGKS9wZW
/HB6NUzwYsy2Xhh+nqCxQ11+DChzcgk63yt+mzlKj0XAJ2rm2IJ07MRKJEYKxv11
UKES/xXJE/S6i2QamRVzFYOPDmBlgoVcXnwplh8G13oEHWkVnUMn1Qg1OYwh8k4x
87bB4Dvyc12wNOdYEaVBkKoVYd3AJDwJuHnf/zOQT4/gL+1mD46XXBKwNVnkMVn9
SmieVBbd7xsNx/s2faRnRwveclidBJYn0h3AfLqiVf+0N1DZED07AcZzj3fyc5KP
6te+QQEIrSMf9tVeOAt91gmsJuyc4Tw7Ah1fTTEWGA3Ndqo48U5336txM1bihjRU
sBAw8pk4gmbHG5txOoZ0YXKjx5yyCpRY9iyuEK/c9OYbunClzMMdfVa4yUz8uz9I
8jW/cVLuzd8vTgINtWwcL/FoL4apVDoXbHhN3Y2P+kLNTwhXkkIOKtGhWJC9aiOg
/sPeO5cUVVPd2Q5kDxn58/wgc1t2lrd52wodIi3wwX6uKdNIMh+tAhE5kOESGKpq
EAtivTOva2KvhsXx+fkiwlKKRF5sG9lehqyXVISlCNPcpm4/MP9OYrk9Dcpgj3G/
+A/Dhdxm2uJuEpSSN93InMHYssTuc8M3WxmM8e3UezD1Gm6crQl4jgG9+gl8U0Yd
4aa4Uicj1HrLyDV2QrozysOAVdDa5Dlj11iFnkFBftBIeWUeHAZVXt7/EwN6qdbA
zgj2qhvRZ99t3PLBqGc4RdTw5+Fga3tnsTJtmRAhC8FoG9GTpUHIFggEvjQLw4Sn
WzXOXxm4rTw1QLjE4jiuTCQe20nVbLEG9QRh+c9lgOCD0Ljytezb98nASLR6Vs1d
upYK5X9LTn/HobCEpTb0GcayAblsbmO/MK+9r53cztIAEPjQFr/ONnc+3u/KbPsZ
c8hbzhLSvSXpwKMaw9rmkxFftrYkI3TtlZBrXMCS37N04t7EgIp+HfQayb8fFiE6
RsN8OVyuE+mU9kcyXN21M6Q0uIDn4kGWVSI50wkgxakIslsxWcSDYwcaLycqCRiC
sMUCpZI1qS1Osv6Ved3Txggmkh1Nshfu4KiPjJiG40PjzO4ryWhixC53DFgY9/wl
Ds+gnh/o1ozCSk5OqRbnQeFSJI8UIO5Akp1GJYqdvKGPesc4tjICBaRzTbRma+IH
2hneh5R3xAoykJWWNXgUQFQGg5GHPDjJnb95XT0zVcg7EqRDkhURhu1wFTNn16cx
Hzm2I5E49xhLKNDCpWHxNul7YcxtlnaqxJsexgxQdUcEjICqG9rGUoot28x5ZW7o
MTEnAC+3GXEOkJutM4FudgTugC6EmIqh26YbCPbEGJmK0KPCMmCkWpuCtX6aoFuI
qLSZHEKddOI8P6DgbQd1X1PoEkouJgnnIxAzIoeipyS4sJHi4WusoebRmBauH6WM
zX2NbolZVwJblBWC03xbMRg2ttzT0D+u+y/p1Zsl4BqwOz8bw3xA1x1Tk0+y7vV1
Ostm898LctQLfbQkst/aaOHAp+qFDGuS6OrboOm37FZtFOgvmO/KTI4GM/Vzb+j1
gWKguaYBvC2ed4H2gApJZKsZuXaXqPc5OLLNERL6pdU4ZOlxzIBznZOv4pGim1oV
ZH6NRu+9C7CgHyKZR2qq8L2hoQZMy1Speui/vftNXRqITvVX645Vd8UtUOMtohJY
OXBeT0lwMj3gG+HCjJcuJLKq3A+sJ0yBnucpEH4G/A5nMfaUNgpyrGD/iCwehnGo
lvxUVMDJcidi3IEoWHnYiTD3LBd1b5tCvXL+hXZziVIamLBYJHv7WeiWIyCVruHB
37tFKdF6LJw2Uvq0J09GiiU3Gl/zGzV+ZQcCsVqPnsmTTjoiwKBlES2KZ7OiyPq6
xOpD373aPChJCwzQcdCfixqBUbo+h7YROm9ctPR4cL3tsJd028rh8uYxsB3eYMct
kK1O3LM8J7AgkgQ0dPUMCEJCxD3FTcHUBOaAzVyK5nKRGNuvx9BvzMvX6/3VHJpD
+OYLJtMKv/PpsqL2xWga57vdONJU5nKmmT52ap8F4KdhJZPDLaURTW8o7hXAWd7l
K5XQO5bukW+dzqOiEr+OIJqDlDRL1sSx80CdB4HVdM7SkIwAQcu+2jlQ3R+V/cCY
x/P/BkvLjZWlrDHz2Wz7ziXO66uhvgH5ukQ3sE506TPMRxtp8UoH5QzDge/PtHJk
zwwT8GRlsn/8KkE5uB4Y1HUlRUoiaDug7Ve8T9jybyZNjthuJDIE2z1u21Tb7g0M
uRkFkTF/xXBrQX5ML+j703EumtrNSdDMoAcIzUINhUQ6lN0/dmjI8mWFJuX5N2lG
4zn4OpWEKVzDA1G7woySBQtdbAtK1MSm2P28HuGhJhzBjbw0HCtV1Lc8RK5oyIvt
vTgOdeMAVAlcBjxULxnbnpPKX3dCKdEjuMSRjiiWlsKtByIVpNzj8+12HeaprvrM
nLeQuCJ12UOw9x7FxBMMstpaCGfKUa2M/EREeSidJ8VzFIXZin3VwcCpVCyZ8+Y4
v/C0ope1Ofjf7FrloYwjrEfEtxEzqwgxf5Mu3gQc/+usdoFXZ3nzR9GYhoNLzm8l
DR1SUujr5JFyg8a9ZjGxHLuHbAFGIU8XhhnvZNxntDAGrOCdtEJrBWZh+T+iWSp0
Hmqaa5NwkIEf6qLdcl/Zv4xnlXfzBVXroOZ0+m5aFCslU4uekJa4QY7xNgXgmBrL
FdUYwxSifcCIa0mfiEfDAMzmTuKh3ejwqzQ7oN9S8z6kSEbEHlhXVK3AnMtCUKpe
w0oSDRDc5nQn4pReZW8m/btlp6jvodL+Hp7XCVmVavnYYmgq8PIDfmqOpo0bridG
Sc6zW+fYaLuWJ960WXP/kzRsnJ7j4HcVdQaWTZ2SUN8vXTsv4klkyhlJbzijjMBA
1961J3EnVPnQvjxdteZUmdiKfvrztNY4JNnwi5MpR4mJz9PCx80VpOzra/U33PaA
ipzA5qK+fNIZmN7iEzsB/pjv1SC4N2oeNu6xte9fwM3z5hpJSU4/7zFqngPadu0E
uPaOORgJdj+Zi7+o9tiwhteOTIvn3GVog0Az5sRgdOzcsfn3Kby4L5gcgikge7aF
8rc59eGVPENPYT4aUDp+pDwd+QJU1hOuizJ+OQNSU+HLNigq0/qIeMP7rdplycWz
J7XAfl6QK72EZmpxsvJChpauAV6sFP9ObpuCNCaRUke5KD/xcpzXprTrVyxiusAt
VGwy+0MNq7NAXX1rlPvYuTJxDgWobDUVirid3j8bezrcYBeBo2EN3LRSW5Agfiel
cr5mTE/qXmUF2+oLj9eVI8cPiYLyYQYOTcbE3sAonsmfnkE5k93hUg5anH0p2GYo
kI64P9PDUxhfwGmWs5JwMxNFah/VszQMEJKJgvzaS+KM4GpML8dwWGHq6OGDPf9M
kca63HXXNR0s/C0KOCZNM19dJR3wE2F5urMSHomOcuG23aAQCZ7FziEvKk24NbgZ
1lHQXvqXLQxkLDqRyRMhT2/gRl+jbV0sqkUVxV1LYtkberWz0YTdy9w3ST6zi+sE
jOADcQgIKzevYGK+4DmNuHqHTAn3T1nTc3ceMlDVPY2nqinxPHLcnAfLJbOcsmzs
hvwk2ljWltIZiXaECEHFlz1k+A+Utky5ePKIgD2ow1ujPImA7a8O5S9e+adLOhr0
I36Iw6XbZMCdMQutzoaES8XBBxRjPFN50sdC1ntNhVVkmKOOOJ1J8G8LMWGdSOch
o6t0dPZrZJ+rXlZJma/NNbzeAv4evPfGIjNS7e4AzzscbqyX32L3oPP85u7SaCSU
jTyxjbdXxEnL+kB/I5NIETM8g5fCkEy1XO/mJz8BrsEU5BrlGSfMtS0stFe2bsKL
twb93dUfhqkAQScF646OrNSCxzRyl8wgFUSL84yzlglGQlG5dVXhnIknd82JYvR7
e25nZvt07Lxx5pkw7ywj80Y0/c5szWs6lZ3nvceJLB4UAuWafoGEUzomiqoYYkb6
9fAICWVPJJuJWboLR0KOrn0v96UXiQflDgsuZRxyZcef8C1sLBT5hgJU386ZDttj
6PD2nvTvmJ1SPkpNnhZ9pQv06e+K4Bg4o3/7Uh+GFFhQt7TmargiSr7dQQssUXgm
Li2vTslzWcj2zksJOsUOUT9mUXqIV4GyAEOrxTVV23K5TS+1PWuH2RM5hxSii2o6
hepxs/I/pgGKa3VQ0X+VHuG/+UcoKhEJeCwMZ4lgfL9hmWNqS9ywyf4Sxb5OTRCQ
uDdVVTbtC2abCb04B84tCLA1obecwuPzVYTYZqtftK2VJnPjb5+RkJcTM7EzP3LX
mlQktnxvTXeq8OJXkfey+Zco5QHnXzNh7/lIS4eqBH778DQgkpBh+qSvbKHaJcGq
B0FNQ+5qiW5txWXJWYClWo3/DrsUBra6h+5WxEwvquT7atWDpALZ8CKHjVsjqJ/J
gW/d9xTJHsu4pjPDhXfOeTF8U+TU+ZbXnVR35yvqdZejjH4LV5ykVFof+ADC2agU
lqdUkrUT++GZvMFtR0+uvYitwA4nsJJyVFvXLmHFSoJwbEpfVk0lQJ1pughqWu+3
iRjOLWDuiqnskT7pp9qdaN0OqyhreT46S/fBFPrjiGCXSM8sjEyPb9iKI3zkHCpd
7JqHweQw0tnO/ihg7l1m9A1VelPUemquWSR+ev2K0cYckMV9o8PUUkBDnZOdNtGF
3E073Ud2j4LVWKPK0a2H75yvCriBEyjJqx7Y9WgthWSwS3z0SIS3TN43EVtrMzvY
CjwUQgVV/2lUIdQ0H2xZ/dwdI5jzsnhzOTKfdOe28FpcePMss+AMbUWF8XdgQoW5
utY7nwkCL7115ostOk1lCs1geRf6HxIssEQ/x+tQSLBB0iUnUidwhWBAqqjVPTva
ZXN3Prb86KzEzNpUuYXvJJSKHF+l2PovT0sbu1xR/LAQYSf0v0LTTlKrlcT7aYvI
463t8zew4jNNWtKKV8miUEf7STmEhDTrfiKQ81hNvpx/ZPeFauTDykhhPwfWRY02
ucsXyWTRb5Xj2hjbSJTUqU4knQzJKhPUYkKjoH2OsKaqX6UBU8OsI+4ZkKH6/+el
zajommhjY1gMnsCWvBa/qDTo0Ukjs2/J6OYtigsImW9gQxC/e05vG5FA0WbxSoOK
cPtGhKIgfVK37uk7vE7oxrJYohDSZKaXr1S7nQE2MiOIPem7YRaovLGtONMdBcpb
zg4g6yzJ3/VhW1CGTHYG3YUVIAZXRYiYajzo4Ln5Z9CtI81EcYHjlpjh09a0DlkK
u2fsA7dJDXyRGAhm72ytN2Sr24Ui8PxN++UlqKRCmCyNkHWhAzi0sAirGBrMKevS
WiWgcrn2GpG1UqFulFsRn0AYT8CV7zVzaLASDEggHTyZmLnDwwGE22dVJ7g9SR2p
pBx/MJ/OIcy1S4hQ372rFhhfmjbAiFK//V/Z7nzgTmLz2VqrV8GAYo/Orkdt5IcK
U07fVvOnNAv9wBNtItJs4a992xR6lpFG3+o8zAAdcNWLgAyCKkQ0p/7X5TmIda6I
smVUsbG7v1Wc5p2aUj3MCrAycoAeCtRjWerp+r5C0/UqpHWi+A+zDpgUPVWEs+CK
4S45Ljj6sTtsT7hmGPxHVBjU5I45Q6OBrinMFdOY8hDnOrlc+KMLhD5eiaCx18aX
iOoNnJwyIyaaYBuUIxmsaero/QTfFpcH3P4Kd9cCQGBY3sNUhjDaGDW2lQumTS5j
259Y6wUkVoHy+gCpOjVAkL6hcEvhN7U7keyjp5dJQ+w/dMmR2Sekz/PcGSozjly/
fNkRMKj1OzFw2rKYwatnlLMD5RAXK+Kqx3s8h4tbPoDcTZ6UwDhTGV2hfGc0DWZK
OKi8STfcZ/XOc2WTeRPktLYHf310j+/En5mlXKLaxSoSsUfrNiglEJRvGGkD0QR/
x/zYV9HcGF3osACp9pNNkY7wC1Gi1iJD2Kqjh7HHAlXnCXaU6Yi9cI8AoIImysKg
P9IkRjC0bEQBOq0mb6Ah0pKEjtXj0YWv+Ri3/ZMe5OsnnH9Sw8SFX/8x03APvGaJ
3PFrTlDrh/Pi9KuAMrYTmuuDXZZaper75s74nmDcIq+kd0RcUX0Rhjr5nbKHukJh
HgjaVGP0pFAPHOy1nqtiVvn6NjjUu8a4SNrVw02sazhgjs6k9LQZtEjtTBM6m+m9
AvD3NN+XNeknkNs1JdK719IVeDZgAwqHM+J/2lt12uGrEv1qJzrzzDZzVYsVQCFb
h2l+EhoCO/UEgU785UdVTEMN+7gJX63PsUIRsjge/bYyv7qe0wu693Deramux/rW
un3U41ZHYE/mN/pIX/sYWKausDOdJ42qBiehLohwEwqe17wVCUo3YF+HV6xSGqSr
1ZNrOGxkF2itI+rhJaMvoLKtM6xUC3qSi35v/HiRsceXQqGDqME1Sx6bssTNDd+f
gcOoHJvijSs21IcgwFIctAWlkBJLY8IhyxBLF8sttrOtwWSvsCDjNo24E8IvGnCM
cGh7ttYjO1CRedxfcuy1D8llJlirEc6VjJaih6Lfzb/VkS20MDQ8ZfoQLLAMnpCw
28FgZmtZ7y4Bh8jLyUi7KoAa/UwWxUgjUJ23AGWyLbETxUH3qM3+jGfxdalm7xNr
3A9wTVkf50Xi/p2B7MxgasquW6jDir5csk+Wxr5RwbvbrMAQ4n/jBpELilneIH/p
NbZDpvoTaP485Q2TcxMvl+V8xdLqyJZImNOscN6VVSnfjm59d87a2kH3dCRVwv9b
RtZ4V68F+uufItwHrOr6rdkzmxe1iCH/0orl4361IQ38VY9zTyFmVNJai4/4E2qf
1kgwf/3w7rthpqeDh+sBkNwxlT0x7nGD8RJ6NJnowQ4be5NHXZ9J7MVtRPZOD7ka
c7828g9celWfJziPLcRt807ckdUNx5Rbsrpw+Vpkk+us/XY5XtOdbiDBrxI3BkI/
vF+G2N+Q5ZE/5rW+GlimNiHJGZ/VcBd8INfbEIkk1rL15AvAM1uugKsr0S7O2Qzo
dYMvheZrHkYmfu3rt0j1C+jHkCzrLzebYr7XXgqLOBiASlaZEQNTMOuGRduj8UBi
MFzWh4pU/2fBm8jswbdT6LCKiyrCKnImcJnNL4R99Z2rj1ns11mpP4JpuV9cd4A7
Of2ZWZGxvtx8XBkAvmftPe5Ng8EzDYzoNe2jjgIHVpujB8BQJaW2A61Qknu4zAB9
N38uIyT8ydqNF1dcLBKKPSx9khgHWLTav+gy1VKEcqSLF6gez5a1N7J+PDADb8eg
jAQDCsDPnJZElsvkKAIHoB4+h85tsqjEumu6PAaJREiPFK9qasKJbxp+lvN70lDo
spm3kBgL/9BYXoBAUY/7FlV1HZ1y9xmYOdtBRKnu/RbHGTtcclf92pvabfGXHUPJ
bmmOMj/llK6CAxPQi4nuyce2YPvDUliEN9WTCaL7vXIJrW/nKr5Q6AEjnE0F41+N
dKE9g38TCbkNwH/RwjwzNK/FjD6j6e6eK9Wc8O5LtP7sCoRmw9QqGhR31GoaD3GO
lIpHIBmWv56rkdwNnpG4NWWG1kJMy4J9WtoHB/BfDlIIOGxC3SZKL1YCQOZN+vIb
DHt0FwNVm1E9ByvvKMRUOMustqiZiUxoj1d/bvf6umMRn7Rw9za4rUwnYGaWqLpy
io5ygwTT87xQhs7MVB5nFY2mA0Nq7RvuJAYO6ajJvH8cd0loPK+O+413GYvC6SWy
BFClG93Eb/paclKqDs1jycTDJ04IX0wf85DVFSzJSz5cGJppq/v/tzfgA3QCv0YH
U7ZwRg1ei9EmC0w3wHAk8O9jq78Lo1JOgBrGJLR702BhaTTZrURvD39LAqna8HOi
wsYaXoczWP+uxoAlX4I3pZvA4puY0heg/3JK08trgq2UC7yvj/L4yIKxkcQFJy5n
QtFDoo6wbXzUFZhSlXg+8y6pFBkOf1by4RASH4F99ANanR4RocW2o8qLDn60GzKR
DCKr+Ea5O/e9cd/G/6ss3b41ZhMn1u3I7DFHkkHm2IBjhfjOgh7CpEf2ycyLlOxR
3aQcqE+j3ku+So10PnrV0qAVHxF6KTVpqkMiZv3Z1CO+ksHLGD6wFMsJYLZxhnLy
U6qwheo08mXNZlX9GUscis5qfMkc8x/I8/nu6TJydaAzRcPr5yQ/uLo0ehIV+IL5
FfWJ9fy8E3nSjfiA71Wg5hTAAa9OYagTYIvj29c9VzOum5igDwXCr1Ri2k4M70Ea
6TezMPA+27nrUq/kMsCDvzf+GQK2ta3/fcMJMrYjSX9oGoTYxA2ABzcJnzECZhuE
KouOwDN1F/bY+Zk/IoHR5Qt3gZOc2C1hGG2uzCzxBxSrrEdEMC5srb/Jzt2NOovS
IIULFZbPUIWpeB59FyjT6QbP/vngFkze3lV00eHqjr+nzKbbhujomYwMiE8dgKDH
/0lMXTPgcEq+WmoxVaWAB+lRq1NWE/X5QLWuOnn/g3o6yjh5y1GpZv9UfXIZM/YI
BtTfTqqbm/4O9ZdDozrqKjYH5fv+CR//pSR3K8VBVpPmv5ZtYqPrf8gojAM7OHJT
mG99oGUhPX2PcPHSCY/zPPewApovl/zdJy0VDi9u5GxZBZrMooHvuiQpk35bzgeS
ELflo5WyM1sE3Qzx+PuQhO7hnGLMVjqdIqOC0D3WW9jLdWO5mhM12yWj3FxMq1JO
c8NK1VaPvGBdEfAjJppDQgtVT5FEFcEGqA+/JR5zMjzCr2bXG2u89yX8dXbC1mj0
Pi/pLOqdn1eHCcvY181oOy64h7rt/0vQJyBCg6r58K/B5hFqAEuhs5Tje6sdvemA
xwmw1C3cDRMOHn95OehCQO3L68B980+IsuRhviZlp+Mi5EtZOfSOz1vw5NzgoeQv
GzdzKGm8PUP86ZED3ewvV7iFlsvo2AB+Or8QpSwHVf3WJo3QaKgsMFayxDxA4gkb
Iy/Hoh1nlV/h8+9nmef+VtQbsPeD5r9sTlDnWWay2gMkktD8REN+plck6uRwdIsB
PRFPVWO5us9psndy3Rk56hhtNvOshNtk4inCrY+bWg102GaNT7La8PQYEo/M7Bp+
fo3IehjLoEqZ0HzB0fMyORob1ksMPyP5SD2TPVfXCYEA6ufG8edaNmlpZDnw3aOu
N+0MYbOKhtlA4bFT9maykKGdUYzXgG1ab1B/xpj4wa1bZjL1oAzw5gm073/DtSRR
VovPnRjfFSR+FtiXdJkoycjLrfO6rd+RP+gwBK4fgjtPdxVsBQBWhoV4IZG+NpUj
QklhIvMRQ84JVnxhC4E4g4u8HwnaAqQzrm0fo1sTAazDnHveqF9hfonu7KJsy4ZM
CWK7LOXp1krS7hVr9D/DhW9NkbCb0v+odeIAJlhxUkLZjtMNf1UkK+/t2Ysb11Qa
7Cl+MqD4T3CBEhFerGHkTwd/z8K8hQP/DubAOtZoFBc2m5kH3/QIH7lsZGeMMAv0
t0hAHtqj2y7fPkfZO+c2hEuuqWQ78SBceyO480N3/69TnjuX8U8WR0CdZvS8EI9q
m+PBMhoAuzQWbiYZfvl+Hh5Z6qjJ4RKgatZuDjKgB2Kij+iDVMCfEl7Wa9A6khUW
se6fWELBA40TM1tYUlWuU+PkLZADsDE0031kg2vfNDXDD7aeuYuMhuIGLFV1A2pZ
Dj8OQhS3wL9kcJ/XyQ6sxme5cw2vHHOBLeGrjZne4WT2jDr5y/aVYgFLr7nnGh0d
wEF1qVOCecFoN8zSrPliLJyi5C4vl6IeXU9OHpaJhuN/dGnte4I1jdxgUfBu0O6B
y6Zif490NqAU7r2IwvzCZVVWC9gHZ2vqhvF4TNfjpNvJ8JKxoJnqXA24NRbGswjO
M4Cic9TUBtOjvBgZU6sXK/Yit5CCYnLJWXE8bOPyJBPJFar0Fj+iyrqGJLERFPFX
4hYgul75186auljL93uOvo+IpBBPMYmuMoAptpnl9ZCJi3S3hceyc2U0riF6jRrB
cnBu3ZI3ogTUD5quhLGSCcZ7czfwKF7WQhcfuWrfc/4VMP0obNs1TImCtL3F9W5C
qRQwUPVD6HB3OZ0vUbvWH2RR9+ntVyxxkj7EGW56nb7zGXHwkOX1mGsiWGxxSecj
wYHKwNf1y+dNslpNNz41pv/GkRGTLIjDC6J+e7StVjFXi/FsToySWl/HUlgkX9M4
CGDxdGm0HOEupTdpRBAKUj3xoHeMqKe7EMvVvRJf/hLvN7NQn5rdrngWPhhn4EUW
eNsnjyWRLiheBq6917Bz5vuDGZtoKPTKWDlz87Ywya6UJ3ucRZC7BiOV4A9qfGv0
4CyVxlFdKnGnCIvMJ3xaTa8/qrgnABx90Exjy90CWFR/X9Tco14qrCW0I333UVHd
Y3pRrGkYlYc3+QAd3Mb+D0vbNEH/9BmlLbDKOLR6sgb5ThGnXrYvL9yYJhTu238t
6HmdavVq0HvW+qRNf4JR+vmTTHVwSpSDXAaK14Rs9RJU2fCiJx46KRgQUMVFn99N
ENGpFgkd5ncekI/okvxiRaxj7Ps932t8ZxN5sHWQ5pSDkOFJPQ5IDHDopSx6JBC/
GLJpyKIE7i1EVuPbXWZl0/C1Vt5BAVDz1RH2ki2iITARtSxsHgqvk0ubPEPqsyEe
T9ZF/GS+quaUiaZfrWnDpufwycMEgdgo9mTxDHJmIEpKrtVs/dCVsNKqGHJNJSOb
j8y7dmavbKqaUTaQmDyIVtE/HFK363nOtJjpuzYDxot5uYBYfQ76JUTL3daQ4uQk
Koa1TxDgK7Sy48qT1BK1yGMC9z5OXI6rcmS/dFIfgEDUjEqFZ0AnoLy6AyqAyCQH
Z414WHYvQ5amNP4uSYosKLAZVvMQIWKIwuixf4jPE9+kA6bk1Qr8mR65t2iT8MWg
3DUVZowLvCLmMCTzDNdXueSMMkVsifSTJW07a0lsxe8SgoqfApWJZ9QFmR9yOnNe
U/t0kfX60b+EfQIwuPZLlCpBFAlUkpjvefbDSBmkiE1M3U39oD636gMH3MjGJFzP
fDkZX1kJ9e+ZrGRiLgjqGPWhhD07WL9TJ9Y+VffKJRjDolVcDHX+UhV+D5j7FiVC
CChxfskkTFgumnIOGFvC3gZbnIpldCyezcc1fotUFtvt5kV7M3xJw+//4pjjs8zp
SM7A0sv1DBxoxEbeN8jB98i5MB9EnPzcbzjGZ/+pAmxbJiiXLC6TkAtXgKBO/GDt
qSnNEtRLJNbEp7i+TWeg/cJMdjUXB++B+smnVfoml40JOVO8xRUAXcsfr89w+xrr
896BxiAW9QQb2JqEMx2uHLbX7V9aZKEIqXPhfWxMe6Swq72tdifMVG7lgBRulrDY
zvFbAzkntzYHtfI7ec6HKFqLLQqzEnNYhudVaZKi48Zu51FRttRNYJ27ccjTP0pt
GefyYscDP3T7Jb8AcoVSkwpxzF47Txxr7fpc67NQNDSQmyA5peIp0jy7X7G8KJip
W+2hxoHavHsQI1/Z9n3b2dH9J3XAxIXc27whL/S8QH1arAwgdHewulgbSYBdVZe+
x/zRo4kj3gT4DZhZWd50flZeVQr2XS7nuyXmkynDczIvI1EWyzdnbRNMSiUOoFXi
HoNOvE3QMKQOyBlwFHFwDGqMUtV4GqoHTVyGJLFCG8zxWYfzecJxC96XBOtGqSAO
vAB1pX6B2RQi33k4T2uGvw9vDpNbE5OFiezFGlzc5i+MNbq1wLBpXZ4u4iEXwvqp
JK8TchRFwx1vCxkqWWEyR2RDCkiBHyIXAlg6I+8j+5WJWlfGw4Cu7MwDjCkR3Rp+
gE62vShdDTPUkFsFhpSHjfsaKj6esUIKEqrlgk8HbxJV7KwEwNIqTAM6yaiw0WM+
58bIqT/r26RbIcapkQmhpiFGn2LcwkApGa4lCEhmzBb4OH07Kf/RKXuZp38J0ads
2a08Lf9njfsjcD+Z9RW9QuD+WYJHMVUj5zBpfYaz12z3/7nBeySOnMxdqpczKwSS
LWlbUtf9uqw4rC22Y/6lCLvklZToMbjAtKx4y3Vy2xo0/V0ufxN580Al7Rh2F6s5
J7CoWLJHOjhAwISvPLlFopsGjVVrN6c+hRTRGpQpca9FAbohYsWKK+KRE9ryQUD/
3GvKKWr1bKJhBfMAhI7lfri20712BadF417N8er3NYLpnDX1KooUcoPnMN91svm6
pUjiRxMPsUYaYYGXKJA80YLeCRPrWF1wiMWQRZGTZG6IJdjUWT5nyI2doNExHtPh
ijOBAESPDym/wptCnVz0+hU4UJ5bRcxE9NDnjRxwDGmNe01VbrRSZ2AOKVmyeqWg
hiAmhN9HjsCmA2FGw3HDIzg4qeduIczkSUMuglZuTvl5qpjBbl4mVPf/ro7WP7DJ
//kT5PSijW6N9xjdS/yg8mqYeg7C358ABxnux6n6iU+t3HhEbUPu1u+ICZ3oJHJq
i9ZEQv5UxQPUf9yKLKOsveddNqT+9l1R45HseqLIYlC+ezFplAITwHVzXIMFIKbO
Ye7hOM9x8lcCCdB1ojbZlGR2JAglmbKx37bg/06o0lNx0R/PCrJNkzVa8KcWDtKW
15FQSmqZSXdBQRy2Vpa/7dwiZAYLISjOWFH7zfA/LlYXGHSLJU0G3tzATq8NVFsf
4ebveHcejlOxvaaHeUID5+GNFyKxoTMa+pYX6q8d/0UDaAv664YvbpHPIU8pZ5Kb
lOyv3PU5mk6KRlZ6CgZLPQV3EsZnxIzUCRqp4nT1CIIz1st9RBtUZj+ePQw04C8h
PEWRZq63d0PVweM+0wXMxzD+O01va+N2lpIOSgXIQjBSuPYzCw3flA+Iud+L9PKA
tlBHxmtew5xJtq/OouKC0Em1/t6XefOgpHq0QX0rczQtLejyouG4GtjNyfCf/srl
jdLZCF5q3DJQXJD9L0gO6abnoO+GEH7oUIactfA5o4n7RyBogiG1L4smhhzgJG9E
AN1Cunz0Mr9QRoINs0c2yIGptDoXeoHJv/m0ImzcMYf3wUzLSRQx6CR/XHFOBcrr
z9Vcivuf4Zr3fIKg+eRoWFgqlQuNKWGogIbyUOZFHO67WiBKzWUCH+64IivyXhA0
3HguBuXZAgQuEwvU1rR0s3JGW3xkGAUsukaa1vABr1kToyU91ppOqZZaDm2+FFEV
9RZsASyyCz4ECWgZvFieyOXTYa/Y3f580dedJumS6XxfFIdZFi3fX2u+O929FcIZ
Db8MsViYyud2cZCihbX9N8tHa3D8tNpthDlWKR34SFo0danLrC34m+hiSNlDu78v
LDXSSePumgg2Sjm1/YTvbt6pooQ/k8Vz0jvUzHDRyLz03qXzPibgWzxoQ4OuNNbu
HvXOM12qJ2imHZJycifA/IJhGmyw7GP9p2sOTwFojPb1NmGxYQFomOjtjaifo4i2
a8PTm9GwLKOy6XwlQMt2jNEHqF2CVK2prosbVuXqSAFjgSyOGS1H6OVses4Dx14D
f/u9LWxzTJcmDIcIs6/rsuFzpiA+aASvkIXyb22pXVn6xMmCo6GwTwh1N0wFYdl8
3Wf1i3HSmYYKn0V8oEwiEkdek++/sNrcr2SwVT1JjQM+Zuq2Qir0swxX/CPWXDyK
WbLzWYG1MVlR/COPrxDjS2fpOOreesXiEFevcFZHzTO0mT6NwcTxLlTZTPgtx9dc
muekbaloIgI8+vbPPFA7xp9p9395DKKAbEnbjGuG0v0tfkOsfT4mCpiqZvAPFKeL
6p7cnKPPfCD0TI24LHs8E1PyTWLlUcFTvWlrFHT3QqCh6RGvUmbmc5srMdq9WSV/
a5TVOUqG7J7lKqeq8azd6OBe5WOt5qL/7qpoSY3wnQ+PESTbtP7kDbkRIeqSVKcq
+k4XghFbNhdaXpBcFIU4IpwVADo8OD0tNQYh5G9w41txnb9oqyM/wVIUwo/qG9Ri
YQRgzcwKIYvPoNa5b6vpQR9hkYEVreyxRRcDFylVDe3XUckVUg3f8L17jf5vmAnC
9ULqz6wj7VXfSKkMd+1I0V7EEBgaEXXr+8GY5tnlWfFHIFXnefJ53mAHwL3jr/ol
hUUH8/+v0t915Sr7dhjVX0ut5xz6dhdRBE2vJ9xHi5wAHhNiUIBiHrwQOoOsOUHi
bxgLvPV0Q9M5i9KhYEFA95sG8qzDhsp/OXdAh+ROHkav8f7dtlFjDhWwkwYZiPEU
HZ7ilXhKwwSDA76+VVbEYtIWZLlJnlijJS6e09bkl7b9WL0CMVql3XKdpZbB1c4n
vSylVleu1OdF1qEES0jiiPAztskG2mHGWJRlWfQifRfCS4Ku7PyWx4PYyMaC5oBo
CuuizZcAdWizOC/Qv2XqZwHar0klSVGoRJUSnsESsSNcwUWQBmYh33xqopI8FRL0
Q2TuqpgqS8vcjHmkZ0L6yHNZU4xwF8m6+FMAIUy7kK0QoCoCxYxV5rKXrEZzmZTm
djY3eIpvhu0elOEoY8a6E5LAYsknIZxPngAXD4cqIbj9tYtmEMapTuvI+7vadty0
7w/HNM3cNtrFHOg13FAdqVNu1oQTXBJ3PD9+07/umR13gJ7RlExqlsx69TYeeyyS
6PmLxZRX6uk/u2TZ1TyRQrNZSEcumzcLlmAlV8sOyDL81gpvh2MtLTvHzwSHR4iG
MFbpPaF+pIbkcQqeUhY0hFoD38KXpFyC+SWAPLOPfWKsjQHoeXSahPLBE72CMc3e
NElfm8uRZVarVPiWOkzmyntjPgThy1Ab9iWKR2armquWIIphT4UQfshvziexLSOT
mmlWyo3iSV+aH+6Blt5SHUC8ompgd1z3f7yGY/yhSGlB2Fv85Yrn534ludrZlo3h
86cJ+TVC2m3i3KPP/+Be5FgnxoCN3PDv/7k6mRnZD+wIfgsrlNZGExvyRc8PYimc
U4A1Sl+HgKrEUK8b9q54ueCir5Vsa/pxwrhQd+Z8LGIW8ETL4g5Mfu0ty7T6rz9O
1ovWg9rx1xUvZF5avZ0yP7mhlk290BRVfspdNpyhEfjkEaruj4PrjRLpCCPe9rYX
p6OJ19XiFALqP7MssdZl2wYSr1GTvWASBLUSrocqLSEAdl4uwItFKe+rnxdX8NN1
5bKtWaBg2BeCc7au9qQnsGkYF3n2ABoZNIYbpAyFnNkgHx/De036iSQWRVXz3b1L
kG83mHPcCY3X6nQ3PiNoycKHFdN/ktLOWV1KDUXZwTo8e/JEH9Qdr8WYdXk2d+PK
U1L5BGQxQzUGQbPr0mU0SvROOOlVxCSzZDCZP2SrPkXx7eHa40T8FRSCwbARuhxV
emAOmXc1iiwDC41T5SonSFfxZ6M1RPuHGLxpQm9k89uTFFqjbvT4VsS4+qWkdxp7
nCBt3xBjeSVI24zOLf0D/d+sxAj+n21QGaO5PDJYArANFSxTVmkp3YlVClfTMftb
uvWTn0VYBqe6oeNRuRKpMcnWs/mSSXMvDjxeSsMftUNvNp0x2ifFwY5tXFAw3Quy
xkfuN20g/XxGRSYLjQDlmC/OuQ4KY1IpIHDjc3/32wctw1AfrBOlm2BJ1KS/4wwr
T14wXQLw5x9eW16A3i4y4lmXBbFWO19BWFurmFjtPvuw1Gp39uMWV/SG4MCv8N93
5doZcTrHnEq8KnyTu4EBEXYW9Om4lC1yAdx3MCkMKS51p6kGhaiZBSYXNlA8MkhH
03MQxT+L//oeYpx8HDd3a5erfGDinktkvR55OYhd97FnjaDyXyck/k8+6Ybzxs3q
DiBz+w6sUAVMDV0Ca8iqWlXGI0onIFJBJS+t3esY03Qm2RtDqCorEkHM8PK601y5
B3hnBtrxaMB4vDRjHlso7zKeQXjvnkGTJOxm6MI2herKuD+e8lBavAM5e7rtd79+
t7iWXujM3IDdReU/Ze9cC7iAno8h37+39/Gv/woAE8pDVH3hS8AE/09lzLfmFTQr
LWffoLyOO8b3yXMTeLBzNo3UIhwcOKh3cDV9PLq2hjuxPyhbi/XthencuTJfbWIk
gw3p2j7BIsk40mXhSTxKvhPQ7RGOjlYohtQlvUPjDwaKjZplS9OSDcViy2I1/KF2
Kru4FbBWaasTr1F7jZR3OJtdRqkXEReRdDQVrvV39BxGPEOwLMgew15wNGRpgUK8
srCG7LrAyZJVhfiKenP/CdcEAaqBRloeWTtk/h3nt+txuFH303VXS3bhn4/EUrKv
yZIWaftURwwzegz/3cwxWDGhWmTCr1acAcakEHmwJ3qZtBBhbqB+nTYDiK2/1nqc
OZm1UjvIdFBLvnmTyHBdtMo1yAHu2NiaN4h2ScBecWw2vCU9ZrYR/bJmVGCLLS0v
o3QGQGb65zHs+LVP02VDMDK14dSmgF+mtwHQOq9cTHz0CWCsAJDscqJUsKCGoAOq
/7G4PFipswhuHZ12ZehZ6XtWlfAAF9GfG34W8ZeWAEgNXIwIeu9sHNuI07jZY4n+
mHzVDSP8D4F7It3dJZQq2Kc4kPGTaxleFxHGVsTtqCkcgiv0VxXALsoCWzFuY+6v
Q/nfPZRizMbGZQIYpVFisorKsRtkPy0epj3QGOR1x1ly20ZuDZ11SotwssCuLkvV
npD0luVYMwwfsyFqCv+G73G8Z/0N2ND+mAHGSaIDNkrJHSdHjMgroZWt3kOeSHy1
D0U/1EtVLq84jufiaWhPCEDdgI5nvJ71r1EW/A9rrq34TpFlQmzcrNqGae4UucG1
zw6VckWt5+FFqn4x1Obw4Sey2DMBm31HRLPn0YvvN7+KZh3htRMKCdOMw2/0u3Eq
5tKBnQ1nkWPNp7C53HX5K+j/02HH2C0uxjmV73qJBGBM72i/E93Ny19h8G/reuMu
JrHrBzTwDbjSAnVg2vbnCLklZjySSF2vyIDVe6Vy9FQhRLATG2jhpWE+fUGVdf/p
62WzVnL8/gbhN2tmG3VcEUzbRvApZKVm3E+IjEB0BGe+OTxUYS5sI+tduhiSEIfr
ggoSJoxbkrctpHLnP0ce6zYshOnhwqkefWsdzYWGxNBG3ZEpUC4OzbG/QHAz34Q5
JYHHiUmk0CrMV829Q/d9ktFhOtyWOnVysTfUPweni+isD2WyEiV+i/R3CD12Cc/o
Wk12iDf1f6LU9bcqBsjVWboOBiDzwmFORAXoyfUmUAtEQaKicPCXhJx0Ggf4iEus
NE3Rq4gYbNwKluego1o/uImVlpXaoBEJqzSmPB8iCJXMKEeVwnrIja1wvq1ggQ3K
2LE4BNh/WuL5L4YsQhyFNliUJyRKWH6C5ThBmgwi+JWvyGDKj2hfoNzzoRm5SKZl
DgiJ0aH+tyluEgWjvQAbMhtiuCstWVARxSmHNNaOCyUjkOSHMvHXKs4/C9eoT+mi
qXcVpMP2cJgd6vc2FU0vfs7b31BLYnTmmpFtVXjXJA/WI9Qa98JXOoA+R+EU5XuK
kBj+JBBxLt0Xj0opotN+HQQFQDvTDWoCp3rxFWJAv3ylI1UwBGWSXvXWHqzbas7Z
n/ipPkHaSGy2Q+fd84Yyt3Y/pIsN+PkTkEsTde2GmCVvah+KuT0Htmmu8o6gQN8H
ma7eZGV3wbVT0JivMZQzW8S57D7wWyWOOexeQUFlGIboHDpdQu/NxPZWevX3h/ZG
89gPFD2F6Zif6VWZ3Wm5iYye2ysWmrODgQ00hTeKbnUH+12kS8Ulv90ZUFEC/5WO
pWesJVkQNEozdBgcpqqk3O6RlPvjpA02HXfiTYwI3DJvSFt67rPajkisrT1DvaBS
Um9AoiITn0mLgVavsTak+Dex6TvfMeetLjvVONafD9orNl+V+QjGcF6Sag6MAbjn
+u1eYj44sqz+ONH8/bHPXJmJTYTcPSsIewJcK6Maz0lfVZY3A21b6IprAIhLLrwv
pA7LX81mAo0kTeTEi/LenR6eKZoeI4B+wHJoHceXKfqqWXkH8/xnaGlKQTaXmGsk
Klbb3t7w6j8SZ7E8WlYp0Zpy4wKUJcPk+E4W3lntQ0O8m3Ga1REo14QfVF4jqJ0S
terqWefrC/fxpiFvotn5miiSuToEJf4OlJJqH8h9FHld/Yj3zP2MWgt2vkcqa5Xt
bsss9YZ+bswr8zYaOMNZcKvUfNUey1qOCsZippFdUK1MMKG1Mq1PKZ65B4IuIGuk
+CInNz9Mv7LwFUFNkGHj0X68soKlr+8fMjSj10OeLrr+Ybp8admUOqmrO9Rh2hcO
RlPoGQ7KGrfqSTSDsSsM4HorJT4H80cK3G1b4XK7w1YHiGyVfK6p66uB2rjmef/F
VDlQ0JB6NTzcfO/QPeh1n8W10VFDz8g2alhhpsiItpok17UQHv3GFOkvqMUQ/ok/
jzy4fr51o5fzG8F76tD/OLGtXyfjm71xiC1OSP6kYEpa+w9UXudGAmzCALVQ087p
ltatoIhDFOvWNTwi0f09kjMkj53F+OzO7+TYYQnSDugG5btGlrYGppQN93Xgf44h
+XyEsG6mAODFzj5fvXkF3FLh46i9XGOnZyklTYQ7f8p/68AmWTLH4u26oI/bubfB
Ck3JuHrdWpEeMILhRaKI551uO5nAL93amVMIaFcE4hsk7kWgcv28LQRRLqPfCERP
xIAXilSebm+e+SfMwAxNgOz+xLpMlYc6SF/nPYiSHHdmtAhFuVVbO2hmT5KxcbzO
2GV5J99Cnb9vXbXMxxVN4B2oGNVAZHk+XVzdV7D316btou3wb0XtZx28rY5cKOMY
4Jy6a/KdZsAdj+ijsnktunpCkRe/X7rngxZ+2lgKxJ0k2I+Mu8winoWuMPya11JP
W5EFWOFykeu7cf0VnMlluBa7joh0d6jrWzs+MYNSNP6fq64wq+hpiRgrpE1Sacxe
amPv5E1n3nShxCunMp8JfKIBOOTturhh3hJF1jRdv6lMAUrevLqF3fPVIDxEaAzR
FxQk75XSten/iZJKIACxd2osh9b9PgMpCog0tr9nsioIqq0oj4SPWYAGYIoGKv3n
yxxW3AAQQQ8k+7j9qCWXGiSvTjvrzoy+4r0wL90V2AqxLq23mPB7f4srzkx2L2C+
ITNVnw3M17p6xgbhololVZ/3baUZSiyl4mBv5QsSOzR4Q32aPvDae7XzoUN5ynaD
iIIR0hprP6ErfFRtS7t5p+DXyPqGOqdqBG5Are3aEcuV4+vJVDTG87LTnRKMPilG
M931BfYLl62jZ/EQqezHe7tht5AhRCa1uzznOjddeb1IVAI/fj28yfkv481yK67f
IDi1rDtdiPopF0wgYyhQAvTiwXAfYVTnpWvZO9hWUUFnNyhGOPelOX6bQ2okv+IF
brIeKeSuOpUiAwRcVNjgj3qf4NDT9cxLrHc5rh90ZNzjvL8BWbWLwIy0zwofjXPq
1Md9+LLmMVx2rgLdTjA0/GRSq06SY6OqTAKR+m6CXkxaxU2yrMCd84l5t7kILzZr
nS4voqo5/p21kxcFVIyJGriWobhD31DfIZ5uclzK/h21ezFdF1snNq7r/PE+6fGw
y5GjFc+86itLTzPpGH2hi/pBjmzee5g4hPYpSmhWh6Unp0fG84WrzxRY3U7H+V8Z
NNVxJeX5jUc2crCK+u8mT3L3CaCCfpky7Mp+DCvjiJJ5xRWUNeyPwBk2T6wnTVmL
VPTOmfsCZWQ6UUoYZifzLTaNby/iBDI9PRXFFzdZA4jFEP48qIBTVARSrunmPZOg
UbzSSHjVOT5Sj67plcQALlEiXSv1ngt4Cy5n9NCp2hOdxblinyw7Evf+u8xVNoh+
3Ti/+4ffuHRsNgc/cziWRRm40MGu7xq0dx9IiU4EcG1js5+ktgdVw2j3igfIZMK2
OT0fyioLYYDBk7kEcZ4B4rB7iUMhkcU0RYpBo/CxpvHGhQTsJEYhGbElAOI981GO
Tqdy+fo95AzdbK4p08L63o/bDJwcCOw3aNheoQ0FYfAci1pkoyud0ux08hM9JWOa
VlddexRI+fqVPx5zJNHPLPplz4nV8ld7j5vK2nTrmpJdsGNvsnGBcpACtJO7Y9sL
8+hfekXcoM/KZ2lrngqhEtEIT16ItzjlwSJA2unq0jwg5GGPuyF5tUsEF2NrI0uV
3j4szf/1kN/Jiod4itNACuDkuN74dZ2ZMa/Xv+WUBkMk3/WzICFVYImfk9wLIIuQ
XKQDKwML9OId/3fPf4xHRB0n+K/0a6evwz5P7MoWra1cZes2b5Nhk0FAAt0b4ThW
LcczUOCcCBVtCfp9A26/iabQeb6+Kb064sIy5BIPJHwTunVo2I1yj6XyMwTY/hOo
sPp1J9gQ2HdweYLI/e5jSPp3pI9XHaGgOErmOzm/RTiY+oqQrWwrmb2JweH9QpLm
SKQebt7uAz+M54U2auyomjoQwTMGCdKX5JOfKD/SJCC3jiqJITv9ew861gd8wkdO
oKQxyCAR3DBMm9m1yLOHAKKs8Iu5qxo6hdYpWiKeW9LNg+8oKeXGed4KMYUKeFxP
MLK6RBDC8asrdwa70PHobSShvfMMOMVcNQBfmTcLcl/jm1mUEY5+IGjtE/i/UiSs
jyyFg+cIChdRYzSUl3HTGweAEM6itzI3DYYVrjMSWedi+YIaQWvGzIgiYWN180jr
UUsLk9CxJqRl9tJwxkN+bm0YuM2CwDdAOSTOB5mGX7UvUcqkq+th6Hvn2OAPrtpl
S+k4PBHL350kHSWzxajQsi2+fYN+ULHonhm7ejGQeVph5vLW/b0E8y8luOBjG5ME
cyls758B8+dtYZ5lGuyUyFbvGZv2GXTEhQPFtIoDunkQj1WKXPSpE8YTKPnC+5dR
J7Q0f1kf++CKY8PSzcqCs9q3lDLbkvFEjoPMz00FwqIwIDg6KHpYwPRQTnJz+jxb
ZRdoeNdJIe7mN1NmkGhPzap+LFfHXk+AY7spozlYsnf4CGoLg43EYUvbS5gkl5yk
MakeY5kPVtsGCM3OsSMQyOe40rFbxCodRu24fiOPrceTJQVY8TziLFKF/2F7tJdZ
8nbMUL2dB5r+J2Lt0FqzeTJMxEzVE/hKMja/Peao8Q7SF6VdGvWmPOPqLeTD5fGq
lhqTERrVubGTYc8t0eB24AGUNUFgUk0iloSQhWNiH1jqo+NkMZO4VGq/gUci3N+0
zMqv+FAVScdzC/N/bJf1aSOM3nMhXU6l4dqK27DrryGLCnXIFFp1WoDTCMt3tW+j
ABNQlpjwXhVd8KKX/xulMQ1qPYgrboWdoafH7ragf3ih9LajtxpWyNEKrSIDs94H
XzqVPDwpQwfYiaRp4Q2Ievq2bgitWUMDQxf3A3HSCeo8uos5xbYgm50GSwF/oc4L
Rg07nLhucmZHBp46zZeIYTT/EChqkl9iP2LmmKcXNh6P4OfJDwhHcdOoU3gKrmRv
aciyjWGiYzGwOdmwuTzvaKEcz3wRbZD0ZFjD4eFtcD5R2rQ2bWAPcnGEwmP8NqOg
8zajUbvcnY2NR2x9EoEpPqfv3Z1X6N0Yb6DnUW26M7CUA1SE0JekeKQ1pQAUP73+
ltRmy9hQE9mkLF6eHPpe3plZuimrK7wfucsE/pnZ9ZdrV0s//lxugFXZJ+BF5eyF
j9OMk2eFwXV5vSMLVQoJTAC7dT9ISPhwvDrGm6JFtqQqKeH6ACHltn2dNFK65GG/
zp2bJ/BFpZ6zrNciZnpdRgGrg7LkLKGm+ntaSoLGl4drbNix02aT/sX1yS6vyDeq
gTGTjBHkREWEN1d2EQO6aK04s6jgUeqFhFOYcd56OrlIMZBdSANC9WBJLkGBs2uT
VFcanWx+QQpVwoa7J2XsZtqICoydLowy3kM4VFGh9Fm9PxDMr5ltPFfVLsh1HpwB
YghD8KnJ0Ut6h80+UDZBPF+1mr5NkAv3H7J4J+mbO5crRabzPBDZiGYRhFBgSUKr
ugz2hGRTDlT+zzPWyqvI03UBim7S6xTELzXvnFHEUT3/l9FegCAr9mEZlqB8iy4f
WOKfNLZumqY31B0FyOkYX6KDjzxbC42SzTjo0dkwD8UuJkMuJo5DFvIyZW/7r8GP
128mC+WLf9jFhGRdd4fIUCCR/Ec3jXAUDfUlKYOYQxIflcT5b11/v5/LctFnR0mB
j1f6rJm1QJUdv0FzX5ykzdDjUNnfZ0j4WUB5tPv7F7ZhFoQAFuaQTeM9+vHQ+2Wh
LtFd2SrbAmt5j2eRM6eZWfXz8EhzIMxtBjkvX8k8qc26+eSeq9YmRIqrdLgNUs2Z
5o0bOv1psRKLVOeNwrBoXXMs3Jrz5WM3RVNIzluz+NE+qoxoDoCnaLbmL76ghY+P
8Zso5cyWyPqm0NAjidwKseTP7ru5m2z3afGhFMosc4dM8oiqoU4G5Jf7CuJ2FfR9
Pw+i3u69QdKLxxz3bMXwjeOowGAShJYlKiS610JDUGjjX8hsGOZdYi6Ey5Sw4Rhu
J5rcjCkBLR/CsbG5c6JOQ+EteVEIr5hBrbG0vkV2Uw++0zm2I1iK749WTc/7yltW
U7ShjPk3jWyQQBuIdbNIa2vlix8ZExzmuC9ffPpKsyBRvivANS7D6kp5aSOMu8IT
GEOb9gWgaVYuRTIvn5ghVOrAqFE71DdoSuhFB0X4w5wOKcfoTr/JmUMGDm1mcH79
tm005kJXprpzsenzH32zXe1f3bhpJCiZ7zKJd0r05aK1KHplJudutlt5RmjfbKR6
lBnuDIy960KXLQtDeLveXu/K0aO3pOGocelTIrPMKBa/zF0pTcUk/5Pgmr3Qn5bU
e62XhxcTY2cXXE0lnZDLQ5YSQ5kQfVoEzJiHLmA10MJGYCh+7NKaQI0HQ2OH3aB7
JR/n6pdccXPkJjkewVEoOpVL17xe+fatoPVsFMHtvn16PRQYN7ayyXLKFaA44QDN
fU3VFOjzEKXghMdjxe2fO5r+tyHwgweDHgtcVMULChxBFgT7LR9QQa4aN/ae3NR2
dcrMjojVbTQwDg41JRe+sgshWuN9vr3rHL8Bm4+ixwsQTg4yXfPbPkvDLRhROJe5
KTGXJG7RwkGlDfUzJoYwjB68HoskVv+iArLsDWFRbcbySxz2W8EvAgpSaGSifot6
01z+5FMydxlUfbytdtsBKhNcx0nlrhK+f1FVz55Mx4XUOncWm6wRANaNByHPQrrj
ZEfztHT+6Fnhfhbt8JWRIGOk1QVse9tVy2SAZLQfXT/LtGbfQ8cJEhR0RXfszBQ7
nxvK63gSjhFt/IK8XBHVltnvKW4Ic7xZLzHdzREC1wJMUKBu3HPCmYxfmx4W6Sck
d+0wZ5B1iWwYUNJY5EXbcWoLUXz8q/Nu6XmSYST2AAIScdUVaxX9Nf6L20wB57N+
P6XFrT5r1Qt1i4xY1G7ZSK36OuBuwudUXJsUf2IjbCibSfpXdhRvzeY3HpEhnDLb
aC5mkdsWO/HM1hAB5XtYg4lSmFal2tMGCAiL8uUJ2mjtKNIPoHV7JMQsup2dSWOn
S9Dw3AdQ+X7rJsCIfYJ4UmRWzMfBXXu4v8gdzUtX/3Gi1a8BO7JF0Q1bKwaUMeG3
NrMJGtafRHSxaUvMkWc7LfAYSrSVAK9UWS51mk8eIFUOhJS9j4ZwY8FdZbioqdvG
eEvZuOR/S6hXqv8uFSHHLFXq3j39DiICWLeYvHV2Mq51SoZyjf84FRDeYCPGFnJ3
bWuZ0S9+qmDCSorcsdUPIILPrJj9l7RoWhIKqNUs6Pra06NO8TYv/Ep5PPV0PcV1
IH4h0Xu/8vwqHRsiejHQYIsiQ1peET5k12VGtZdT8E4ahgcqNfcSX5dbyLdP1xJZ
WsbBJT8vENUA2ud4p7FfitjcljPgxa9NbjHLvjlhez+QieLo4KM1NWEAmxyQedwa
bhQPhi0dX4i07OzVuu1KXFABHgFOdJ0NqHo4xKGYpFrgUDtxFWs1INr5SmKnFxGa
hEfHge/6eMeJ6vj7vaAwmTVpchBdwkjF9tTNYnXvVTBn2VHPMpYWkXj6t8RmEUL2
6AAwbgJA1ag+ovgSBxx+ms5/Bm3WREku/GNQ1oY4Yqzn/L6iXGBpwT7vmTh4+YOy
/N/N1i13m6Y+LIyVSKWJKBMZtlartC2KLG1JR5pRKshsFET2ufaLVTcVI81o/lEQ
VP2toM+5UKi8XuqssDYgJfjHBwzP1QMGwaHl0OekrMAAoh1wEuylepFoL2Gh4Pll
ZtQqk+ie9269eTWKYpZ1vB4QGrUbo8fOiVc1fe3WGoUJ4hOzQ/C0SRNANBtVHWf1
qzUzLKyQI65XLlveR/kEwcw0mVreIubO2RsRIEJrbwnTGYi2U3FZnRNA4YoSrC++
oI2SaY+VHDL2u7Z3ZS+DnGOxaI6ipKTUu9YioMvAFspepEWOXZePNPArpMTtjKvM
WakYiu2Q3ko0vf8Ku5B6/UFOcY9SYXjLfuP9ake1kNoU574O6pWGBBSK52yEeHjE
ySu9TZ+DH6yjutHFZMTUgrPntMOpQ08lvW0lf4d+AOxhL37AGzKokfuKuybo4VpG
/V7lniQ5PCSPFtYICmUav1j/7TfNTzqkUfbP89B2KrnpttV++ZYa+6sTMqpapGpq
o9oaqCh+QSqGfmGXus73HvIJT6w9h/I20K4sVg1TaRikSUtH0G8BvONEUfZjo/8v
UQBAcgntZwZ5AYQW5mIXHDrhcec1epWtpb5HSiWFGskD3x4sXm07oRGs/wADpAMR
EiIDDiRR/qtldi0pAOctLhmmtivbrQLlX90gZV0UwXajU6vq/gVbvRZzcIWUq6P2
gtYjQnXf4Zo4XpJNgX7LFcxx4rJaaVPG3NQraSAMGoyPq2e8UTB/eurJPVFoaj15
qWVIOQlTKQlj+RQ5T99J+l2kaexx0Equfm8UHcMvqf178clsvxJuJxIanh9cE6UG
0hq3SKPVBe+lcwduRgNWn5WNQRi3daJBfZDY1V4LLwvWlqNp/wc5ToBCD6XCjuwz
iL1m5MqJ2MrrUWxS+iAZnbMtO6TpdKIDzIJL3tL3ttclQVsjx33rnLbmBW6W/nym
JyrZluOe20vAmke1R3ymvOUT/RMy5oq2dxSc2np9e9IbzBXUsG91Ad5RvbvkY5sR
zdh/mODQLJZ+5c0F7Q/rZgPx0hSry+eC8WRIWB9E65AUGf30ojypOnY+yckuZkFB
aL1IsE4EQDaM5XQrG8SKEmMWVEg4I+Qz+cDOfwQ+zxnSPWIEmR5xHW0WKCeG5oSK
wDleWIaNjv5puDLetd+3ySCRm37ipoZFV5LAGmvXG46SWv0Evc9dVwrIJnyZEYCx
X2PjvtNrNEd1eS49/siHbVj0cviqYOtHvP5zsnnajNYH79i0+nW6bXLm4ZrME99g
xMKL/eVOIieH7ZdV2J4Zx2oEoz2nGdfF1VXk4VKyxaYSus2NIZXrztCjGbltklzW
IGe0o7ESgrcG4j2B1ao5sKPS/7a9kv1GjuFDJ2hFnPdjT+WXKK1HDMVj0XHV5Sxx
9kUVlVDugSfbU+auRW78ZjW4b2OH4wjrOSNMeWdzpsUZTHndfMAWVv/gOuTFLpmO
K92MKx7h6tpYjVRAWn6e/IiL7gy0iNlTSD1wa7iNYw4gQELuP5mVLsIitNZYrSlD
Q+dz7iWKzVdQlXHqwfM+g3FUwA1VR0BxtNijtSjPRW4jyMbR+pqmBeMz7cUaS7ou
kNw7n1HZbtBWU7MqP18mhJjUtg5kLD+/lIF3+KpN1KKVVD19vYcxk+QO3tW2/rnm
ocQOFCJslMTbsqaynM9B0/adPHsUQ4bQyUh+JL1c3IlC4oiSxFR40Kvw/efAHE7j
wLDSCPz+eoQTIIrQkXKP2JYkbHpblzaKyMt4impQ7pp2umDTWmPIMWhJDkhhpbd/
Edt1dfkEJgAFX0vlm/suYrhjQZAAd5NDQy3kjzxPTZyuAsloVhk/3vR5uhgjDFYu
QSqLVr4X6vFKBJHcxWWRbBQEhGROUNTkUaKtEQFz4j3WMTbTnQ6qLqbIFfmgK2tO
LQ13yAqnSt0KMLKDEYv4VybcuC25/7qLNRn9vBaERFhMxyV62poQJ5z+a4kNfDVb
z52SHRwVPBxIUv496IK+ur2OUFcf5ZHMf4A8vpxNgwG337XJbToqtQvim3K8qrXb
RybDWBKhUUxUGAO9Lr6gmTuwApVHzS4ELU9uwdUwnBWuuTBhIubLMPHf9oYC+6v2
BBplKXnek0gh+RyBl6YDPG/PC7mJmsJf6EQ2neKVPhRzkZ/xDCLPLKaZRdQEVUov
pDKHLvDu57iip0SDnwjnY4AleN3Rdnphbm4SnHSzC+QKF4yP7gZ+b8bc7h8zxCJe
u8DDNInElqnqMpsKsIODW9gAvfw34GCCsi7OkBkTJucy6dBGY3MsoodnKh0lTwD9
7f9JnfKE0LjMzmtuEmz4At9BxDP4eo8HnfYwv6TKZI3i5OhUX8I7zbfVagSRAK+G
rcY1Ul6Oe9pMF2Ay8f6NrAdlTkxZmjhHDdntqaIaMyN+VZj8732VhdC69JU0eKbg
A7XZGwvnyNRmyNYge5tftn1xQGwNSDi+wD/byKIbIe5FsVvgiZmBtn/F9L9FqitU
GVx3FDv9QpgYkhHskF+g0C1/NfDDDxedtSv4h2TIMvVU7YmSDMOZ56DVPaHtgioZ
UzF1AiCP7cHOejDMby69UH7tVdwDy3UezW8gjdyXKsg64f/6XQmai6pOeEkICi9E
UXH2tvoMmpbySB2C2lVMkAo41i4UXYi1iQDjoNLYE6IPQ93wGEJOP7sPajciU4Vn
uwB+d4tqXyUvsa0WnF+Fa5rdYi0rOBMyaHJpn3ZXqcEh11pUq9L5EVuvsAFP+5xw
QIU4ENcBwmBt221ARcBwQC8oQiyri8k2DEhTWjfF37nkGeFsUbNDQUXwYkPFgjZN
OreXysbyl5xIML7zcuCE5/YiK2j2JMWNM6XfWUeNLiaQVGz/QgUXT3bdHPxXMjP+
M81/Szn3plkARW5EmjtNvr/KTunKW/fuiOqt2a0V/rriMzGoL+Dv/AB2cPThnTGx
ronnuWSU8jRcVbC24GJupzuJ/nGGn/+wx9Rhhqdj4zr+uWGivR9STak0muz3u1wR
+1sD42mIy1reIEIM/A0dt7QiSKyZwZCGXmz4wbFAJvuICIzDYuSJnzG6sdVAm1Gb
8gE585txQfAeIjlymgPTaq9kfnXBtJiQ53274+ewXpIaLWdmBs9ZCwKeePGRzRuQ
Ai4EVSV7V1iO2Vv1Ik74Vu5aqPIREdpo8CNjja5ZMhXNjEMFDLkQZa3se/ElCjws
mtxNz+GZ9q1Y1hEG6BJv+2jnVjcAjyQbfpt3CTRgK1esZSZRpHXdQGIQ7ltOZctY
iP2Vjfq8ruFSMYKIm7iIeuUhPhEw7/mBI1bDEHSj12JwWUP5r49+LMtroVPCrvLa
zQZE16zYFwJNQccu9gXBsvuXWL6o6tzgAEcwlaCnwNKKbR9ikUiDsupnn1/B96Du
0L/uRxkbYUBdB9Ul6/8g8rGtVAe454PnoYGEuapg0WykV4zt/NEcHNs0aD5gW4P+
UKZTDzGwR7J1Hj9eLGn4ujeEMPcXKdaG4ZBI2KC6RdSA7xuKlK6agVFhMmRCYhkA
CSdaajAHOmab+tzmjgoUaps5u6xaH6rAhsyXGvz0icumM7iLSowC+eStreWJcyQm
q1VnP5KL4aj2xLQNsMgtyGsyZHjTcdAbONiL9Gj1midmsQ9BS2atrOzNMmBvXlaG
S6078FugnauzHDeJNwxpHsRXPslNKcIIhsCTBtbL/O/MOb0oDba56b7VDBUJQYl5
7WRyj9Q+PDcPW25d18S9OELGBEzJY979mmI3VggSqQvEyTMNHr40+/WeLE3r5lDi
EVRMLKHAXivpMc1yKu6stz+WR645D77bWzXLnfVXYLlI2DpLef5ruUom4H5yv0ch
46/3ao7fN6fZI0Te6/rHQVYeGn6bsqfoxbCS2o7LEzVqvH0X/FDuDgI2alrZ87qh
ZqSl0YnJiRKVU8z9d13gykga69jewRkFv6znVsRN+fDCyx7yd6CZTn4ZEyrDxSat
FTUOG+QJwdGxJRpZ72T3GmYNwjlrJtX5lFiCBGgMVYhoBhUbLJTslVJuq8ESkaYg
AW/dy+VYHfdxUP963k1kq31zaDIvJUUfRa0eMJvfDfMcFPF4flcnS5cbNZ2BWr1y
CaUvD+xT+JbOIx5onP+vVCRXzD4J1q6jeyTHB0dAwEGRcsSxhRP6P2cGtQ/zXuUX
g5Xi24zxlqi4NxXJT+3FskyYYSCJ45VDtYYhlOCMAvHLtITnVvfgYik0kk3kT8+p
iMvEgj9JH1XrrNERaVw/l6dPv6hcqIb3/ggsR+lM1H6fAscZ9FUuhOvnOxVqEOFv
TXkRn+TAGH2o685svaE/jYz+zX8fNx0NvcW+3aK0GyWSEs6DFt6h9PHal7NVaY8n
VAovpp+MzwuH2umy2Kl0GmxKjZSwzaGrxIRr4bJy7hS+QSDX5tKyb3J0s/3N3NKe
pipQFk48hcHam7EfxLxAC8vknUhBFtT7/vALglsErkGFjzbXCfciiSTVB4XjRKgU
GMUgAejFKL1vppwXs4c4FZSx1hhN1e3AHGwdIv2I52tSJMfcsuN9tfbz70gQGYxO
oFGGpjMm7/jgC8SUxXrPdoMb7jJvzM60BtUT1YzpLcPRXyDRAAZUOuHQEXrEMwmy
BdygM4e24EoxvZbRqGiLuHy8COsO+EPcOXZ8Zpru0W8WpQP4pgCpNy6PPuydhS0o
7KuAo8HJSxpXVBrbpXh3efvQQhVAse1EEW8OGPpI+v1l/ZPv2MeOQmRAUITMM+TF
JHuWun3X3ocpHrWkEtZwbLHZAS570CZEf6l1x25BrWhj9e4W7KCX0YTp/y+gYbAx
uG3Mv5blaewZ+PtAEszVJ74XOsKt/9SVYX6w7a0nee05hlE47HN53dQYBNeUyL4l
q9feL3NFJ1At9ylo4lbNT8BSSOOsbglM/AFRHbjf72BV7yjfWhrtJBGO4hyGsIRs
N7vljGhAgWShTnN5e4M19ykKrNkQJw/vBaI/O/ZBPjNo9yG1Mk4Sxh8xaOyi7HaW
B8V5MXpI4MnfaAbn0LxKvOeVb7/xVsPs6AQLXq6Kg4LpOz/gRv1SjI7QRS7B75gM
SYD1kpXk/vKzPQ7czosgcOlGLNn3EQslIFvX40MWwKIczVMoDLxVqkWKAJb0PsU4
mV6MKJnDqPIodIeiKugJFvlMMbUyf+3nwrApKfcl+2PDNiwBbi1AkC2hKFh7WMOv
B2bM/yookW9xo3/FfSVGzbt0evTDZkZkkdXu+Kf04fHVqmy+WaOjanVfghAy/pJe
NuzwmdVgNf4GhMW8ELGg6aTfvES8npiJ1jJUENLFHQz/k+b9FlBMej34CVLp3hjI
Pte2JVBsiJACYY6+MBIMUUvPA6qp2/qJvqZam/BR6CatfSXNVirywOx4z82NLgnm
YdiqM5WunbRhDKibF25ylHVp7wXlSyudPkBwP0oAqFHV07P1aez0cgKi3Jhm6oln
i0cVwrjhpQD33StID4rMXnroVpPx3kl58/1TehwbNwNWuU2vq4sM26PZ0l6cQp/O
olmYwEYwlqOMkJe5hwXxYBti4GHyGk/egOLt2zUC7NqjGVn5d2/3fQp/Q4jZwuvZ
q9XQHBMI6TmklpLkZ1JOeVp6TlkhhzQo/bc7TA5WJVSBealz01HS+ucH1Bm4EUal
34Gt1nFRNkXQOX7KYP38KcU2MIUkDiyPkNiFutR3bSlZ69ODhVDd2XMck624/yx6
ApDDfbQkFJnzEvDa/ZTCYMSiiq6CvZzc3jlVW9eDXraolTfkl1Iw/ICag6bJ8+6b
j77I4TeOCJFCkQ6D54zDr1RVc8uSwRuK+hcaF00H2L2uiV3pxnELcF8fJ99C2QbE
jVk9jhK38UZ2Jntxi1XA8lN4nHzu8MxcCSwMRgfCzRVZGW9MuNst5o1CeRUKgb8v
ne5BERL+m4D7BH1ooZOXosGrB+rYYpcUGmzwf6DwFAFIN89PFxvmZ+lyqJylT7VU
7Z2QoK0SJT+ZafanPDKSSVbVPtfK3gqBibykVIyZr6ME4WZVKbtkmyevnAAIsvOI
uWYlyg8OZhs4mNG+p9gkl/nArLP4NB2hMTZ/kKJXFfjyBaB1VWEWbL3FKdXTa+ab
Kmp2isVW/oV/P909rLEc2WBfpWKN2mD8HGrDaZBo3v1AsU834xjtB6lbEjfqRPY4
D/ypPNhYyyiCK6glfNVERarXhKn+5QmbEwXt90Dqn+sd4S34J+HwvDj3vYOo694w
DVg7Qeq74QgP6TvhFZ7+SoRHVyuJtgQPQSrKI9K/CYe8Vr31NjD0ji/8HSH9cufL
qfqEWtXCk4Jbr/N1YtEyTStLCER/wH63EMO6dnY6q2vYMirJnc3SY3Jp5P+cjjO3
KqRJOyuw54gz6PQ+emXNVkRv2GdESGT1HEKdS3hOPydyh/LlvSeWfFQxwk/A6BoX
euBx8hjaesMvO69hLoJnwEOnnA8ov1vRBBNmjduSaUZzenoSRfv9w2Ve5JJGPkCg
aQvboBKN+cWpA3sh06Rm5yMOgr9ARunYiEf6JdofkF4EHGiUyJQFOH5MxE6VGOXm
T3iO6ox/0FNJIFkr7gedE2CIsKqRDZ+ayCyplrQ4S7euoh078gXK47Tt7XcO+Y/s
fZNZgTQyp9nDZyDkkmo+46aMPtGermerlrvAdVly1eLa+td9OlzKrl1vZdft3xkb
NqUEoQqp7POQRlOXXDyAzFaJhsnNwr/ZBOR0Ks5wrldddJAUDK/Fa3f7xQtk04x7
u/jb3VKWGDiuXXbl71sqe+SOEE3WCN3d9t+C5sAKvm/B39hAPXdjpaogGyKMs20h
Jg9dPRIu4i/obNkl8khHl4KNCip5xqFuBlEXXQ1AQXQrerRrhFX1WYn+vGFwUBj+
mgJut/hUsypIT7Ys7+GW0YaSG/eWioVt5O1UOihcQkhmgfFTXukyNWb9vsThysbY
kSbHv6+DbRqPAnMQW2UhjX/SkdQH1qYew6zfzqj0QwYwQ9FdmeIUp6O4VpWz+hdx
/WiB+O47xXxQhhXw38ZNLqJWrJ/F8sR7fmYBx4WY2it0efZLZXYz4yuxYbfIM3oK
ZI5aohyx4jjj4o12ekZ33UClWM3RGlKFqaNkFKs8TiJI2Lh6YyfPNdLLETYatXTQ
g/g5sF8EbcSP9gKq+C4BAa5+VCpcciPSBhKci3trm5440uQpB1BlV7RBkHiW7Abb
kMfCNKkGXJ7KBwItixJlqjb8T6a4vT9BN5FYBzltv63SmlRRnx8w1bPaqGhpa8UF
QEY+viT5FzXseaACiteEs4iZDHJvnmyZ75GwnIr/yW3S8Vj7dc1ZNMtgoQCJx5RI
yVGz+I99kjlSruqT2Vdecy8zGb+q3n9mqBzXrcamaWBa/ypAc1pUgE919Oh8fTOB
kZs2LFSGtIEJdPJwgYodpO7PvW/F9/EL8WFfw0WssSke2pUHAM18QPZb8qQmgJAC
pKaZ5EdhquGDamMVwog/kAoFnXgmE2M0WzmNz5FYmzR+Eq6UNnDecMcEaSzDvkca
WdV4RyklbIHLL/3w9KMuYjrTKqMcb6aZVTD2YVZQIHElJhbeiToHLNB3WRdAg0JF
d2enIa+BGa0r50lsWpROSEZ4726/qbtN02ioSHoqlszjZHfphn90NzBuMRKOa9fO
WYFvShnHzy7qz17+WTqwkYtCUimfEntdnaqPDbrKss3y+6Ix3qzKJT4Z/xOyejFH
IHT2sUUGMkRnTrVhM1gPgbRn45Pn+N9qNFyCf4oOp19o7iOVhHl5Mnv5cVf6Yqsx
fDG2npNsBhIQscgEZwTgB/JoeJDNfjsLrHMeck+dydtobqrziuFHDfJB+FowrSI6
7xze9+rCsVCor7R/l/W1i0dZgTJGjyZdRdAsIDBkMKQcHISjXCg+koAOz8Q+g4AL
yc7Sn7ZhdUcUEB8BYjkAaNbWjM60k0tgxySWmy+GHYhuRT8IQQIiVspHnjdv+6XN
fk82mG5bJlMzUVLCjkBGjKKm75p+wf5X0fhS3ClTfqtUzR5nZgLX7dNw5orE5QJq
F4/46Dz/Kz3Bldp8NRAdjqR9WeaOIuzl77dfN2FNVywZfXGhcAblnf22SVSzGT5/
jb5h15pSGDG2HUsBxVpxFQVhPDhGW1wrD+Y8NyE1eMVSaSl98EiMlrBwMgrsyjM7
HSRmicUQp29tFUYs61zQkwhMnnzOg0UHExEaqdiP1ZC8HA9HoDxdVAuaRNwaMwj+
qkjO/wLbSpszlvRTPSJ4Bvj4zXTblJ68693IFMPY6bgAFBpFSRgSWrOpQku7196u
vRj5sDWVRILryOnNk3UCR6H2bGjxEr/LNiQ0NKXzU7ME+SByjnWH4398VCyIM6ha
pe4MSr9KKOhdeV5yjtmpIZdqFXdDBP9GWmjAUwg1kZPCZjhUhXrwfypiImXM0Yf4
D9LJAD3cwXPDfH/WjANNjf+ER9mMaetPlV6BQqC6/nY3szM2Fs1PQEBuliev2J7j
n3rt6kDZXNLqC7UxavfrfYOsHdqulZ+TegAbdaoSVjzCdurCjWV1o/ieXnuYizUd
/mBRFj0JP2PDCQHXo4ui7uKR3yyg2LVSZDZDnCwqYphFdrX9eX0LLYUoAgYKA1q1
j/QJ9UZq6HL01WSxC3F6g9H3A0eSMrdA2eOrMjTKbuJ47lveDI97Pb9y7Yc5K1yI
soY7mu7VT1ULAE7AfnSrCqys2UTojrHJt/n7mwcKHhZzvP35WkVmq50016r1QcP0
LJkz7rGDF7NL1gGiEpRwQsW92pi2llKFv6UkGnNHkJKX/K3t2ze2OCWEDMqyh01K
V3wd4R+sJLhrHx7X+DdyBJpZ9cpY6BecYA1hECslyGirxNdXkV8nEzWZa+RUel8u
6JLIge7WMWylPdVekJsSydo6MfVrES6DkN3UxYeY9m8int0T4xA6zFChQ5DwlJmO
IDw8pR6COCd3VCWuFusrzUSnQg1CwUVofC0BZ9psV1G16IiLglZnkRPKMYrRXVFb
C1z4zBn1wIZslLmp0mu1WWbrg69akzSZInsPauH2o52t1BmktS7BokXrm1xcM7JZ
PYKA9G5mTi+clyb8aftl2HGSsJcUkzz8jXun7ujH0x3mWRnirC3FzBGSQt9ID8uY
xh7kXGGwsOITGE7EIwoRN/5LaZDm1z1wJ5XW/ruih5JU9ysPM0Uvi4Y1o1rTH827
i42HilA/g80fwGpIe+dZyTSiXm3Ga5tRqSCrfoEsHecu8eYNUXYRZKJCWlonrUbO
hukKXOeia9dGk64Wc0Xg2vXO00McVNbueNhbYK0ah8mOCu70VqD6C2mB10FwGW2Z
vAyZeGHUqIFWFnseJ0ITTz0R+BCEBs0ihP3MBYp/R6DALHaPYrr02VSyXURk/6/w
7s+parQrGbTk8XGDW/oumEX/zbWdl8ZVvsybsEM1EbfkIR06BVQO5M4G+jv3bG6k
etSWU9hVoMBX+z15usknrE5pktJWIGZPz4YiGe3nj9kjC2t5Y+msx9bda57cqiA9
n1waFBmUzMX6QvUFRKP8/u0WOfAz6kTQqO4aPL2vTwBDJ5sOoGQwjlcLkfSQSeNi
jWPyNJ11u5JMCCl1vH1ufTdPYjO38W4e6MpHDT2ty3agB2KU/04wwV/Qznlkhivg
p3YNt99tRBx6SbZQ+MyoSMzeeZEapK9dzik4Drrxuw3e3Y7Lk+Y09M6Y8lgY54RQ
VYLnALTjWHYa9jPh07eNzqDshb+FW/9mErZn2IAlKVqDm1OZvSC9/fkynqGm0fvI
DanOYlgaUXvU9yUIJju/qqlBwjNv/IonzowHxYqsSHtZsPC9R9S9GtxKq4aKoAQn
HEInvhsRTBTwZq1sDSKYQHHGAzbqEMdAiAd3/ejTgMwVbBYVgZP/eAU7NwARNvee
lMSIQWFs2zLASQyZrVJ6BZOtZwSqRwULF3BRFAx+OKBslqcuu5OfT0zeVHsI2CVX
rLQaEb+yIEdMXEj6XqiuZbntpwowgM4KE5Xz4tk4F8VwNvFg6aRhcGirZaZP/Ygx
UUpE+sszbz6Tfzgndq//360xMr/G+u9/xGc1N183As+1ruErQ0PofB0ZeHh1HfQp
dBhxRiwzLurhP3KhJFg9Nx97WVPV1LN301nWSsUkBjxXtGbEhTkJEd6RB1M5bxYY
MA+HjdwQDUMyc4v0Xpe+FToiRxBz7AhxRpwVuoO/BUGag/TONZQLF2zhEAXHS9MW
HmkKkQtLKEHpOfz9R3H1UVcyep+l7yRj25OftB0cIgK3a29UmV5jX2+g6FQ95siJ
uZiYUuszHpew7z4m7nsLifzO51KzYNL7mhEsKpYRXbSVhKoxrazcLA8eIVvfByfU
6yLqqZdnZG0O8s6zIAWmFDGxHfObnDroZHvSN8qU5Q8OQgZ1UzTQC58zWgLuQqoU
fRULbEoQcPotTQ5fQZAtnGRgeK3qp/97zeZlwo3TYlokglEscKHiSvQHhNakfjga
uqLFdiUtTVoNMcsjW5lrRzUu1lHldd2g7HGfzAnlYqrXlhuv4TStx8g7sZXZPt9g
iTj/nSSC5G0vNiywJIugRAzg2NWgewDvSDL73nfmV77WnUO3+nV01aAbZ0Dl4NhM
3IrGJftV3wII1witWq9oH6TT71dgf6v6qrjGIn9DrDceXw4Y667AU8k6rp66KDkd
kIw1DFUB6Bu7BlKzNG3NE9k8wzBUtzbi+v87kaODGBnsje5Nl0S0Mu784SbtuYrv
nhr9Tmaf8/qoHE6SrxK5W3SkuKDNSmhgjZqYTKSf5jNjVqfiFuJ2hV2iftnvkOsn
S+uZ0BkDTszxbHyiaijPuPCJixqlxdR1RVIJwdtIj9/NWjgcCwPcakNzXWYtSryv
0tmWH34qTLgsLK/h2npCdPJHwkiirMut1/7JODWkR7XcZRN3LLFXHH19C1iwMYeq
s33pF+TP8LVWfUscMqXHDHd6Ai0exZCRs7925mkZh/0ANrh9dYwixp9YtKY9XBjW
VI7TZxO4nfWbgyNBljO6cOBzFKe9LoUPBWLh21bdxK6/qlSPkwzf/PBDYk4m9l/i
lt7GuAFneVsaDum3XmAMwNZlmUR0z16STOmH23IIAb6ZOZ3K5GTBEPgK/lIvLhCp
G/vWNBqzqvhfwyyS0ybYl+KLZnz0lhw5ad930Vuco+LBX7bGqYJh9bg0tDmSA2d4
vo+9TUOiPPKScK2DyPUcr4nc0LNdSjkgCP4wX0NzzJXMlwZZfJLgF3kejArXx3na
RkJREJsMzCDe/f3HZQzJWluhVftlXlWqIJI6A7lhVHpl/jubmsa+H4FeqOr/C9g5
r7xcoGnG/+cvZtlgSceK5Pb9fRXymeKnlwJBtknkLQEXq4rHdndupxI9SAEAKUWR
05FB2e0IS7rOO9G1rTvfLFjOx7m4carNqHSZpHzBQ4qsdBXBqVi9KTSedmxQLRSR
ZmctVlMzevj1qhC/iLO4Yt6sAhPlwh6IUhrCKKZiPJuzc9iVSsRWWFe69pCw0YPc
65nuYjLoKjXH/skVD2sVYsps8lKC9NUOYtQzwS6GiCewC2Ec02Ji4E+S2CuHXiBS
8nF9nrflCscB2G5lmLbNUkJGWx81ilyFFAG3BNQlui0kG0p4OnwS5+Icf+xeQyuh
a7RyAtRhed0Fom/dYWRTnEcErIm0UKU1H0byXs6ORxB1Plyb5DZMwulYi38HDkub
K82HJL1HCm8A7q1D0fWnicNKbRwhOQgXQjI/sVNsFEFB1DMslQhU0f0Lpt9PzWM7
eMtQfKxZ/PMo8S3o3NNztYqQYRQdDTxzU/SXCVraBr9I5XhAxvIcqqZPXtYTAsE2
Grr4+y9YDIlVtUutIlx0OUs2oEp+zIQLfi1sS1wpr1TvxnXsN13kt/qqE7iMyOHW
fJ6BxwhX7AN23AkY3noR0GENZC48/f2WgeB/M9FsOqJeVYe3RnLD44nRxWCRZZP+
u8U52DIgAmgv7I6xCHudGykJYkP0X7pxGYNWeMK8t2BQBlnInegI1XGXg2eosRml
KAhMRruZQgf2EAvJSg4BLRDNaZsAgd8kB+TNEXFXzmsgMWveNeRfk3SYObgund16
aM/KfrFQwZv5rtOJ1aRtLECWjjDubJ8YxhocAQcVvTZyPiKCW/HTdZCmljKBhav9
tui2gomYvBINY54XSQZRi/zBCKMOVzbgfIP0r1P/71bmmkgqlrKhuF6NzLem6Zfi
RaBA5jy/rYZfhHYdIEPF93/ZzkwkXn0Pe3/wi9bIhcSjHlgXcc16padAz8L2GkYn
hHdYVGJ9xeZ30Q15XdhhM/vt/6wVgX0I98Bf03y/dtwmkzyWUzkqvRNxjzmXKepY
+vHMtF6T+H2RMvAFJXvzQlSeBz/Zkxhz50CptYK2kWMXeGh2WJ7cwwdOCSIYuwK9
kUlBpm3NMDJ5jmgkz4xBpnP2CrLc9Dk+GCyfwFk8mLvjBTpbJTTjcrGK+TJzDGjT
u58FFzTCRQQChyRj5WF0RNTHCGUFlddXfgyzob13ND5mOXbz9FotsacduS6HqJbC
QmKXroOEyuzjpoiMYWSAxYsxViqag7JmKBjZ07tL3qdJNFQkcF/UJXi2PsmGbeRx
eJij9F+XBiuYZi8QW88ySgm1IBdjMXRcKRxvPeSb3s2xx1HSmJ9Cxf5ST8jNEwkj
V3NwYn49MEZqgs2AdeiyRJ2QA4ljeFV0DnHKsWORPWTEXEZmFxdnryBx9Wlr/Fw7
mmeAoyUcPxQUzcCqUbKX+PafPUIaIzSw/8pcRYChitIWSYKslhxmO89pFNN8qdms
Svhftetl+lfCFYgI/9IYOemMoZUOmmg4SEN5ymFFc3srDrpemVEaMAoH75fS/8SX
pUWBJ78TJ15rhvNvq4wwH2FfMCcu5vCR87UgDvcBpVKfPM4uMUkHP/2FylCDTJF3
gjaPo1wupwWy49+nQMRNmIeRMFolUrVqTzZis0PhP1xTbG8MvRqk06TqOhrIk2YJ
T0EPf3DAzETJ6bZjiDjZWJOiYGNaurEpA/PVWzbB+29H6I3rL+BtPm1bdZUgRVI3
CEFDs60b54Tv6P7pIGQrlMdqWUThB0nioKEiHPB509LR8GZqdTLNWbkXkJ8YAsxd
4sVX7fSNyTPRD/T59wTjALF4M1gFWdL1AGqvPpbGBMrfrPY3z2YzXQPXnSOUYBai
1KKWBXzeKiCOgcsfURPuoodA078qUZylBEFdIKHT0PyGz3QOhhIe7dQO4R1vTwxi
Ry8hGPvOqr+rpHUOqCAvCEZ4TuGA0aTQzn7rq2Kc96b403OemcneEehq9myfiZp4
Yefi4FUBc2s8wK20d0TeDhttVu0vtlOTC8FvRff9cmiaLw5YTibQ624ztXU3NGWI
wnwdlwb52wfwPEQT2sa1c0HOqnK5RW/EissyhOCjNMjeFoRgjhulwn50o+LZRhpu
pznt5VtNYrRM60wdYm4p3bNTDp/fdJ0bL+FEKuHSj2btPwRx+fU4CtQF9fZiiCIn
SCkPw2Zpmm2yShexR+AOAjbSa2R/+AuROItKN9r0xq8muPVCFW7O2TZJ0pUHEZc1
jTEZs5jc+PGjyMMA5drhPACszNnv2BECERLixn3GOUb/Q+0V1m5Fjp8VLkhcTga8
7bmG4/e+BTF43JWPNeOzY9lbvNbLhiNSXkVCppJBZbkVAaOSv+zqzk2XgaPoqhoS
AwS1fLkOQJwwZUOU/ufh8Jt7bMXWUYwvurwKRkS6j4Dsc9nyTEVUJajf9v+VBx4D
7VGp5WNQXRSgc9JrPTLkP2B6Nv2fiJgoEFAR7LqWHyXV/o0PT3oeZt+D/tBDMZJA
Zv1UYcyIu0RhkLaz+Wkn7le2SqazAcNyqYzNNGBvtBp5DuZ5gNEMXCv02k8VnTGi
oXfIrOT4fklzw820JIXEQFqYnb4G/Xr37t0pMpoezkIFKIirCgrIvheoHhaaeVJI
DOwY7BgJ9oq5WjA6iu2V2vrKcrbwMl8d3vcoeMXazTuB+PXarSylvG3DLhFmqW+8
hzd2AoY/kfHSwp3sM3KqNnQL5Sm7a8GBAHPCIimlIhgIPJV2K7cMzmJYhELmYxVv
P6SrLcXhp3vXwfl8oqisgB8wylEpDGiXnzWG7t9iwwZ0LSV5/243h8Q36lg01Dyi
h2S4ZKKEgezQJLFl+VYgWPXyU1kS3keTJ6LH32KTWNhp8ZLvF4foeTrMIFqA9YCM
cNgh1KDGxTuQB4cbOnMEs9bHSLnZYRoIlj6/xhIpoJFRHP6d5mRQ4E1BhEZbl9PY
ZqvvBy0fnDijxMr8jPekxFR578MxO3+CejxNoSSqG+bEPNqHR4hJG78BDxMzs8iD
BRYkl7ud/n2mZTKJgahOooMfQMhpVdRy+VirlqxoGr4OoY0UY77PzwiskG+NHqcN
rQ3Awma3RFbilfP7bp9s6pggqy9B6Auti5Q/RfxoeEK0G8s2ZsbhqBgU3a6jHrjt
z3Mqu3OEBV6+AQcciTQhTjZPOONLSA/RZPlRrykPCDq6XmAQn3M+XkCePgKclteT
SCbQs+od85wvvZEsVd2IedX6zNWvmmKV95woWqoHMEpXwHgFuAhQ+fsmioPdyK5c
0mc6RmyGqkGbT2rkEq90YnYEcxzvHqWLRHtkGtj5KHJvbBm/9W+/aqjcyV5nRk2w
n6wGXX2Udgb844tvjPSV9EutCHXss3Sip8xRLEA5LsoivKF5XPs8hPiXHDuBgZFB
bME1TgRlmLPT53oWOyoXZo93wAsBTfMj0RzcU25wNw7XYYx0BChDyWd/O6dg31Y9
i53ATPhVwNJG5ZDNwMJtM1vZ4zrqpctHSc9bPWfyZ/DeuLSC3Sk+MkNPJsiHhIbW
dbJmxGm8rECXyoL0n+CpAD0NN9m855QZMAiE9UG9Q4Eh+1+rRZAL5xD6fkcJSZE8
z9M9hkYf44Fzp7lm9C6T4iPG5h2OJuTJg6L8h1zX81+h33C5oRYsIbCNFhvsYwF5
3fh0eDZp+LkwpF3euLt+Hvbo53dJIeTbpqSqHw2Kt/rt3A7KDkiGBeeE19Ws6vYN
d4fsBiKj9wAO4itvBp1gIEl0MzHgnlpKckNGqt4Ti7tWeIH/40F75LxUJOmfBSJ5
4CUk0+N3IFzT4oWIS3Qc3OLL0UdNpxJ53tJ1j2dMWJgSyUkynb4NJevnNgwfwKpx
4yIAfeI7MjHyJOsD8Bncoz7/f0v67vCD1y9j50ElobnvnzIvwcRt6uPc3hoe/io2
2dHsF6naUwA27ZfJDaf/TctLldVrmW0BJtbhX7A6Ho7VPKQzNk/c+mIjVA+cLTid
oUeGfXD8NyNDsMRUzi4BzFsElp9RYRvWcCWkdCxIklkvBluntjdGZyeCVe7RaGUK
bm36RkZrSDzn0FjSjtSUTXfgkHZBq/RkXRQcb/YGLcRA7GgfRp48G3n+WtRRPgmi
Dc1MkWJ/QYvuUb5GzVHDnmUNJx5CVCMaTPIfw1rCGVQEDAz71EhiX0a6ubXbecN5
GAQdLDyvVM+ZHpMNWvhgNimyyXlb6fx0Lric/6Cq7yww8bkcj8UszYlpVFCKoYOJ
7IM+gcTBfHdpEv9/5DkaGWMh8/T4zS4ocTFK6Bmw+8OeO7t05qHRcKPMiYPGEVAL
uco4feZYLoZkKN56WFQ1rUcRujU8U0E+AY4GgdeI2itRhO5OHZwHI0w6UiDUZSJb
znPV0gElfC28F0UjRbE+bMW6p8t9Eq9pqOX/JYaiMzYopi2/g7vnH2HbZp8JrPqS
2cR/zpIl9LuTtLZOWomOs58+Hh1tisJqnOlpuM4/2V499n7CaaUrp1LJQsWMMxMR
TA1NB/mGPJ1gBEBz7qNvQHGFl29neBFUD+zMw0q/FF+Q097a2YAcB/HgvlaMIdwZ
4eTRXd4cJvrdYTfqzmtvHwWEnvQt2vH6g4zniE9L0O/6upUJSGoOZR3e95zm9b+i
tDcPtdimJbs4uRcGafJ21W14OW4I+kaU2YIN0Q9yjY/jec0y/srneB+h17F6eHLn
2m7Ui7obGLBvS3LPNjQsiFfwOogtN8k6YHZwYvnTQjYNq3Zm26cA2srxJKz5dfdj
iQbFAFVJFNmyQMfuverJ8dumhUbqPafvxjy2I1J5F8nYX5vmaLDE2jFlSlyEwZ0v
9fglTZPyQJoxvWvprqaLVwkHefrof/RAqrG0y15K1cGbheTUIyQi18l5iF0Y1UF1
Zed/fpNB/rAQucTOq9oYxTNUaYf7J60HP9FvIrrCt+OmvTSN0KoStL1Rd4y6KWgs
vIeSMCKP1f5yEkkpOFbRAys8T3688bMUCefk0qMeXkrznjCPFE4oe9yDa89tdh8W
gknmEH9vaUoEHvZnECnpssgASig+6X6X9TbuTqe0qcYRhiq7vp0T9L7sM5xJYt59
b9ZPpnDekLLx1zaPQPhq83Kmg4UVsczoXgD/+xewrpV/eAz1pRUefDyfLzrAZaJ/
hJvSBVB3R0r4xelxE4llhVUeWDCm9O/F3UcOSLZP4P4Kf57pKzdQhNidKSXU+6F9
q3q5Av26ekAOvGgJ7JMxQSO34gLQNubOO7RMF7kW1L2Q4P/B0MB5aOeBvkuBc/AP
EepjpFgqtusVMutNdwySA66CQMXJ4a1KkR4KNa/4DOjF+B5u0/NV+FJUOV0owu7N
3HMPBw1r36qA62bSjDMeDC29qM1K/GT9F/Sv+I+Au2jgjSSgzomHFbxfXQ3adtHl
4TqJfTrwVo7HugyDS2Je70djLJxR4lUpfHLJ6/5sy/MwIGsc0fAa/0Q8Dp/sy7HT
xWULM/gyTParfz8YjWeQnEvlmSj0SSZFd4Rk/Pq8wVJRgmQ7qAr6XxLonBOqbtlQ
oa+AyInvE9x1Jbnca//WvjsMTAE78/Jt55YbisMWYy4hzmXQ0Jcj07g1CpWN3Gyr
MzXZxWu+kvhLQl/mxIm4vdm3uZ+PlDBRJMbt18Kie7fOoobhVyRS4BiIdsS9Ou3M
Qw0KeAtkSGtOQFNBjDSDgLctn5E6JnUUX5MGtiE+/JUA/fy7Nf55kL1vSX5BhH35
j+pcKoJN6s7qz7Gaw93Fk8bBG+l/dvv+w+U14VkDJjOJ74St73QYBSIC8DwSKC5K
+2ttumiAj3P9P+aZ/rHEYY9NctOWc6RfEA5Ab5k48UyaOOtkT2mBS82GCmfC2t6U
7NRI4guuzSwuw41znfYpsEoSAtlP0B3y/0vJJ5MrYFZ2I880feszn7snOtja88DS
vxZqLJ9lVQ4vICradFriQ4zE+5TV/SkcAkaUzIh9fVpHI6VUZ+zxgw5q+7Jfh2XM
4+E6Fj7mf7qocPIIPW4ux7CTpPftM1q6jQcCNFBcj5KSkUIbzfF6mdilLuhs1O9J
owqRCWnSfXwJZSWEuYDIHGP7xySd/pPNeo81Qw2pqyH9m/3CtUH48fvVUJohZXGP
F87HOdJ+KYbc2pkw4dR4LM4p/B9lYeSQTefmvhcrOMvZxBmuTMNO74DRe7eKlcRZ
ztUPkW0DclNq3yNDZBqNUTf2+YroUTvlUEWNbLd6KfvbasYlRZoQlHWxR2beNDFh
T8VNbkFnBhcfQ7BYTzHkcMzJ9fsUs3Qt9YOBSSgbnzttCBLucT+UgvFQL+yZlaDD
iiFJh3kn+uefCQnTB2gNMdcZcZAChjyx0UoBakiazzvsREWhe3XjCJI9ic0twPkT
NHfFpRa0SCX1Zd0yPI181mTizdrvLgOgTsDKqqRBEla4s7VljC5UOnuoobxD/I2g
wQEH97FbE45NX5y3WaapZYk7d+VldzZvwNZcw06VAhr5eWmIP2kGWgLerPL13X//
AH4mIoO0KUFG+4i+sxTAPtPsENbcpkkw7EPviJYfrB23Wy09i36e+Qb6bFMO4R2C
Szk3OVOk0oWJMiUePdEcZNM/jAe959Vt9rPMTZFLVmTqkCIOkLHxZe9fAUO/svwY
v1RPkN7QxDgTgdivSCrxAfvnQ8G5Z6qIwZsfresfeAJ2ddZGnL+T1YWWx8kcHfl+
quXx4Bz+6ujHo/vAMfAYR28vBhk+7MUojb0Fb9tV6OJrOX1ieXjVB8Ty43h5FK5J
JtulzUSr6rcEi+FT7D9hRzttm+gdhRs7t3WsXSVcJG4NwmuOgH5HTiDv2GSyprnH
7owITmw4I4qjbj/pkgoiwdk1+UPw6IcpynEzk21rsHogZ2LHKAGgcmwjTXHIzrgf
3ri/bUghg+3DHSMGTqvdsrqJl5PhB1KiHgLELyJVDhzKtkrpsbm0YuhE+7BbkNUW
yZqxdEClLXqwFqeCz/rKUOKLSwXjpThjRTpp0/HgsG8KDtwmkIlS9xPO1UFLzkEG
2riNI1hwm4DELS3YfgZ3n6N0GuIPPYHQmz50bfSayOsnqxYwIyhU8mc68pWMr9iL
JpoorRH85C26oeYT95fLR8M0N1KccH2onJqDKfAZ70/kFSiXL2cJZc6xOElgwpDK
l5OB+TbmKUXdWwfVPDcFaFdzXIL6A9Bf5/Q0h5mEkV6gyHrOyhxflp/Zx2kgu50X
Ydr0lbxwTrfONx+JnOqlaQQb8EZ5anAN1A72tJ9w4KIuq2ySpmn1YCLdDOvHBuCe
lXvpqX2qiQaz/t8QAA4hYbC/XgoyH4XJ2wxaf0nIOyojs+FyPrp7h9759GhongTq
I+ixy5Uxaj0qNrJw//AXqZj0WzaMrWln1yuln2SN5wycggxIEOt/LXMDMrGHp45m
yqmuECc2Jr+2mx9yJ6ZJdYx0lg+4Pv6vgPSjmEpZiXlfU7TSPE8c9AZfVs+oCZE9
6oQq6JnxZ2nW1TLafUsDN8MS+DRFUl1XTziHWh/mbuvQmSMv49NSPzyVMF6NBah1
YxhUHSEP/J1hNnNmAKs09cl8KEmSNDhvuj3zJPJ4+J44MWfoVJ6HnlAKJv0g/wqH
E4E+l9mJPYElAZH6F6dWncBJQt+DT8fynuvYeHAz+kP3CDswNZrWhywZLtPAd2Ee
ga7xGEtyhoY5cxHOBtl0NR2brt73/483l8vW7wsplLXp8o7CL9NrlCEW25qiUCDs
RSZ0o6NHWwOCBSUfhOe1bYMImgIuA4I+KD1lxMWjsyUzpe7qk8KgGgNpJRQaRxlW
iF8POkqYTDK/Z3Lj7SGrSGjzX2s6ev6dd07bs75oP7CJSTcSpgspKmcYUL6DJQiP
vsHwiIo0TPMeJwsk5BZW+cTKRLNYVmQhkgztWnzp42R78inQzEes9GsNBqt3Yktw
pV8DqNgzDWv81tEuBSPhGZFVSwdqWQ2hzDi6HkAXHaCLbXq5dqqMAmGVKwz8j7An
kjc4+Y5017wCi0wFas7UXDIU9Y/FaY1gcMVPdmtUXuq025r9lUMgEnuZvtkMTr1q
2peMsqe72lseiL6Ao+odaxMEI/KkKQxLKt4cG16QL3EnyEScZyO/AIVgddwM4fwj
AyoU7FWt9MuKL46BwGHfxlDeSybRm7d5MlBlwspOzfElJy/YXCsclUiVhAKpVvAE
ThT040lGdwMa2rE1jr/JwaTa+xxVTzWxbpxMWu3YIcPbDc86tCa1c4a1SF9bRCs1
2fSNJ9DyDSCdph1dKDQZtMVuUlGZTK/ykALNapHM9jBTRdeOBgfS8Pay/3DvHnpv
33ZOZMkRzzvjvuGtS1tcYQTf1johQU15CI1mKtMMaUulTgbUU8eso+yMpZN+KUbj
ievuEeggYl9KkoBAnNQjJSSmAZXVIyZ7YydCKy5WSCLMgnYmtwFTLlwslExQSqbV
Fwh8LhJtG7AmKh0qlmgp5BRBp55zEq3ycu7OhbhAs17EvrXpZf7UsCGFqqHS8OcU
gNtivg8l+9kHBDQeJlmqxL4nutidrbc5gCvMIYTgvVTTUWq8mZd1F2MHCabiw4Pu
sj/xN/S2+uDnz6puNflyPW3Nu00z7m2tmWOXpVImJ3UaXW/Zej2apcX38rQa88wM
Bew0TKSZogn8gq0jknIjAoOC4C3AQasjnWSzh2uGV5U9toWWo6Ze3QnJWM6H3WgN
y2UVM0c8WHCBbEHVNvjJSaCP6iCy+cp5HTLwh9YXWI0v+vsRWBJR3DMgmbUsmpvM
BuPnnmvQoaxqPbIQDJcAM6W4E1FL/yVjw7wpiI0njYQD4+MNzdkns0Go2eIHDcO2
zIsWWNI3R57N45BbsOJaqa2N8nb7Rz6hnCCvs4q2WGyYulx9HyIcaqfw/2Y48Ka7
wrfqihX39f82D90ZKM808CwZ2uy2bW+vlqRHKprS7TohIr4+dT9CzCL1lHPu8C0h
hlc9VBMBVudZ1CyXJnsonQLxZJsbr55Q2fkzSqIPd4gxchJbcQ/QAPJduCC3lKY6
/8pnj7EFyovyKvSjia/AuKiE1z4WG7PBKyLMPA2giYtvAxhE3d1G2rx3xnbXVXHW
8qxPAXtMWjXLPQDjcr6F+scXZhSuhHg5NNlW7PFyGxIIX4atCc8aRgaBfe5rV4/H
b9oFazlzXshLoWmEH197pxKVDC4Qt/fmIF9ulTuosfZmG356qctBZUjPKTzStPKj
Wj4VrPKSYfC0yYDzmKGBPzXLsJScKl0UOsHRRTVHnNA62PTDxvhjgAIEZuRQ5ChX
maT8wV4yzy+DIAH0ga1oUTsbYzXbfRWR4ax5HuwQXImG3gtWvObZRM+jftFWLASP
RJoBxho2DAyLbdXXV1Gu+0OiWKaCq3js3cmG+xRVZxMSxuQlRueDP0x+JKzlxxi/
gXVf+qhB9iPA6Grs7BERyokQnOvg34Do/9UMHDwQ3LkhMGz0aKWhbbdNnfNBURzG
kgar4W9osLpd4XWEkSVaDwetc1vmewOCV3gegds20ctRsXGEpFlOQLjS1qvV6BCP
sHXpm6gelu+C6Sk+1AFbQthd2Z8d8KLkufLWh4M+8pemVVTI1gO4T7J1MGvJK7aj
qiThZZskFfAVBD/6MP3doI7CMaoDsERxiBXTHycV+C4kouf+lb9bZGfo1yMUkC//
JmRnPG+aEiGKr+FmEMJlDbAhlbrzqGuyCmjWWz2MMRAL0FAtw6/Wls/9hjHf2b3m
+jXGw81L9YJZv85wk4ex+dSDgc4mFXEqYUsu/BRoBN0qlcn6/K5Cy0sOwWZjkmQY
O10prLohr3T7BbUTQf7BCbINTfzUMLh5Yot1d+eESzBtnzQCJfAeQOBJ5Xcg5iMc
jq4plKpY8P+pa5WR4xgyMv7tOrHgJbZeyGDbeJwmxIWSrsARbqg0KJcmPbnbF3t+
gKlSPv6kBcwL3yPkVQKo4oBdax31k6pEcmyJCLpH75xmAlHhXwZ6eV3PS9HWF5MI
GRGMfUZsQPspo/gLGDOOkjjxi+m6nqhk7Co3sGfbLOcz32gcJl1oZiFbOpofKSRB
/x8v48zexKg8Thqa4Y7iFpy11DipT2eX7Be3PTCDSAc4wgIDTbb7qumPE27ecHT3
dfhjTaJ/vP/smZURpU8t6itMWofi/X0x7gKKa3nLIAn8c6ekyo3J6wj0X4sf6c0J
m+8FiEjIEmLKjclXj/d8cuFR0Sk9hcCx4MnO9rEz58olqM4paAdbSSaNEGWq/bJF
SYh4ir61I6VGhMbV9y0ZaFbciWj3w85BgAIjLHCWxsn/Bx66k91pQW5qQB+0/EzY
EDSeXZzk4R8kBQ9zDpdIKfpP1GJ0HYCxSiSL/ZMV2HA6gihvSHRvxzqs4i5DxncD
oV5rgkzSkXpCebvwAQvWnRzdJGqmcmDr6W2unuhr2JeAzzlIml1aCYJQP4/QcZD3
924h2GncNkbKtmtKC7o72mLGqwPsfCFX/EIehUWLSKbhVvckNTdC56UvvVx3/ACP
DtZ9VekJpkAOTpFOqvgco/b3I//aflgwxFeT3tf0AE2JG5IUyxScaBn1sUDbWqi6
T/UOJChojdVpLcr6mNiDxSQCKvLFgFi6arlturpX0k0ozWHXy5B/qhuy3V83qM8X
fAcwgs/CUVg4mi08ReuDxcVWqroOLjpwW89nP3QRAetehvLVWzUr4UOCy845LwJQ
2/HwVwKnXKrNdIm4DKwDNEUU3i5l2vyeSDhKxjiGv0jcIypjmcDXV+4gpY0RQ0WD
AtMB3TLNQZNsQHIzYHSwh4EQWHWWsf18LE+l0jHvgUCig3qQwfWQyR0K0KGrW89y
X2M+ZEnlkeUOqfGDmOH6AvpQUD4Hl4zLMlVfBS38ZAIbcBMj2koLjJs1YcnJZyAE
Hrd+zH3igzvOt922Bu29RbBoaRIRxnEfGRUIWDN0vrMj0J0k1CZVxUgmma8QxlCe
bi15J5EHcjseW5c2lykqUydhLI379ahddfxxBam6nYph9UosiJgCSpbeUFG3j8WR
OPh7jTfO3nPOlJ/HvnmqAMgFPnsW4f/ekrcN+jfpSCO6OlfNDiKMuAbcPAmMZMVl
1T6TSopnVdneePm2trCZF/WouQra0pmsHgN16dIDvDNHdn2OtDSE9UQ4xHmUILGJ
dlmK0ESugUJ91E3n9/kJgx7IBoqUBxXHl3b0DoalAJwdvd8PJH5Pep241yRe762g
Fe4DAU70CJNulC7SMr00wkjhlqxoYkDd87WTU0047uV52Y7mYwA/qGOmmUtId1uq
9CIfBetOhWnv5y0M3jcdZ5vYkhNaQpk0B0+oLuKDmPpq/2A8yQOLdaZwgRwKuitI
KAAC5POoJg19zHMDN8PR8UxrhBfAH9FlGDBuxk8QDzuVP/eofAEtR68UFmIa9cIE
kG9/xtBkbDmrawBHsdQFn7i/226zvZ8t3eaAgvKRixYZJMZWEPRS51jwUgLnv8xo
4UBN7/f6oALpN0anfmFOw0Ea1hJQSl1Px6bOBb4vioLBgMzXLLmif/8DgQDmZTl2
1PgokIJ/CEHXNpTn6OSJ8Zvs05ka1wtEqGLr26OwG76+QRi4pmQ6IJy/c6J+IHYF
yLfZDgIs2QQr61wJQcsgKUDK9XodE2PVVl3GtAxIAUEu48ayVmufBmgg9sXhR1vc
tyxRwHhPuxMPx674gJ3fpRkpf/BC3PgGo5hGoCkKGpucCnprw7BjBCy2ev8HuN4h
d4cH+LiN+vsVLz21qh/EWmkrqkOJSf9hYrTb9gsYgfKXbe3ZWO85+yhSxwqm4Tuw
fXQpoOoi/Mn9iLuVRwV+GBCgUP9OfvqyiUs1X3mvGPHDhvWJeel5z4ymoH2WIteQ
8uVTQ9Xu2Csoayhpl9MmIPnE4E7/nM1yqbU58hTAljJv6VrgM4M5mesfCarJ01RA
w+tqNpJ/YXtAewc6WBC+udZXLUr+25tn+j0RlV7715v42SHULvz0/00j5ZsUmaca
YsM7wE3xSWdz9YprFSwjjpCmFadz14YAR6kfOvgg4HzMP9NQNz7yLQQaTCkCuZGM
WwTGMcGqDgjEOeObeBidVBelp69xo8PJIOJR5E0sstm/cjr73cuhdEcggeOO6mpf
IUEiMPx/osKyIQbzVdnkvCsVgouC/kE9Fe1U32iSSFeqMvP8VDV4kvxGyxqRQrzB
bUf36DcIq3zhO1b+h0KW8qJ6rzuhIxmA13TOvTihyNN2aNBXyT6CLEWw2Ki9lXUx
JrBPwdcKr5CBrENKKASxX/8aC/gVc9nYHRBTj3MMi5qg2Wl/mLN0+pBig5cvDD0s
zEOsL/yxSLZfDABsPJGdMW6vKMOHaupPsW0Y4Q+wWZwahgtMV3pPCzc4hn2ocFiS
hZl74mgqrzkDY49kTgFoeBmsCehiZW6LXQwGwzFB4Oa10oD2qTHU5JrPt2V93bo/
xNTWXF20X+wHF3kg3s8fr7q863r9dFDCqz+hxpLcMslD7Ov+jeX72v59kFwgwNqg
85lCqCHQa4YdM7U8+ipE2X4RMh9gz1gx++u8Jeggzdf4ouR6hgcqpq2pXPIHBRk4
zdy2xulXBwfjyskdXc91/PV1eIS0QLfCe738eGIhaG235Ktzc7srEOLLRYGyNW9E
KXfuqHevefQuPZDhtn0KLHPgJcEKt21YfySOvJ9GLAG2awIq2ccHYvwte3I/EcM9
b+0MdvA5M1H1X4aNVSMiqbG7BLskCxVWC0gh/yEhPpTGSAuonkNseR5xnpeQCZns
j1ofTFRfngj7EUedreQRpvwvNphz1qa6fAvcs2NwwOD5cm8b5S38tLAW1frUAHbY
hsHHCyYjykPv3kaNEJtD7hZ0phK5ATw1xZvrxm3cDhYquJXBF7ItmC1ruP4oSuBF
3BsJSuwbNuKL5SM7pFIUUyqD7T5XjBbtiZrBwdcHCht80oJ2w083J1UV+7mFsofM
zTkG6bIVUNqDlac8s6wXS+a7Qy3lCfyWNMix/x1TU+USRU6eQk/RsASHtnsxRnQ+
1fs78+KUsH4URpF1QDm8DnF7n6y1QmgXOKhSQNJWNTv+JTMi7Drbj3cSPtNvWt1R
kyjOBS3PuBqrN+Y2g9WXMyOQLE5IF44qyiW2LwcPvavIPFwEZvX4+hnovYIHcSsT
tnKO+9s0IkJyPH3+HMCAxhd1xItH/7ntXS4NBAjVmGQ7aTW1qNG2EjFIlfQZkbLd
nK0qJaZfWu+1FCaofF3jd240uDSIphJEXZ7dt7mJTQNkH7+BZ5z8ig1JOtmllrwY
eOBMRGaXbwpTiFcwNWJuRuLbNkirrroEC+4pHHW9fHFb+VwVlituxo+4L2lb2L5t
WA7HH1Oe5eHz7TEtChtuVq+6n7abyx6vFZQ/1jaztjAskXU82hgbgDRK7v0Wvs5n
nIi8fHtXZl5i188yYsBCZ+XOMRTAlMHYUAmExvJUc1cc0w9NaftSO7/Xc424skAF
948Ly3bWUoBu5HMxK6m978aBx3Bg4rPveHC2MVs9ouUOuJxo08dyOHVSxzU730/E
0ZMaIYX9b9vR5ZuizB24T3kF9zOS5ByeGub7gAf5eKLgkPr9C6NCg2F/M9HaiTTM
kMbq9fSPjxkPzBoEXl/X6QYjyLiE2xfyp9keKBS7aeqcSsoHwDSvRi8HxgRS9N+C
Fj7pSN36SxhSDkeucwxEKD4NLhjfJ1z+AfkDKkQ/5tWgQHtIvWMWPrA2an9NlJHW
86rE340AOzont1RdoULoHxdrvwcC9ozl7u1DpOAuh3NvPYHnQ6htd/Yzg8IYtyEm
QmyhOLKQ/4aZK2ZGMXd8lYD7kZRYNRMev4NvJv6C3LExrBVzA5InrpFO717XuZSW
Qd1jEuW3n40yW7Ln1c6iW777yB31II72f+UTVP5UnCeC6C0LZvCi6OEuHJA7I3jl
7E0faqrlSCXpI7A5tP0zYO87yKQdCMA1P6+k5GVQfzXAxFJQFpRXnnG8FAAZT9ba
gdZbbiROkoHAZ9LottACgwuRlRJ86kbJa/xgPrGwnRvrHF73vQFLS27zHHWcfUmg
XBUhlb65KHEXxQwX2HjquWGgBJXF6Jm+6sIOVMQBrzGqTNVA6C7s4XlHeOmdRoVy
+QB+IBmDpjlqDMuHl/Nu7Mf6bS25cxc3ftxCaHhffSbdFx18/ja/nAziFToq7pGY
jHyLLbOC/VW46QsVYKtRzGxoZxg6XD4NJ90/bZ+IxLdNfNYlVSn/v+nAEAPsowbp
VmfGbC5g4HopU7PcF55PdOXC3KwdarsBiJ/KscqemCybse8+NmtlTpl9nz3POkNg
WoHqPwGoCBEv7g27AgUqHf5sDX3d5UaDhTF/yO8dVkesgyHsXnSo0MxyraGl/mi5
gBCT+2ivAQlOKx3BGJpcBtyOf3j835y1mP6oWDypktzHGCT2lbcJme2yDE19+YG5
s17pq6KhGpalO/wHjMQcStDeXtKQ+3mztiNgM3jpjRlI1Rl6OovVywqH4Hw6QiUU
r7THLZAyQFjKiPBmg7PxFOeW2RJVhM6NmPWSONMaZtl0V9RW/9dsXhN4HdNn8++0
2LSRe/6PVq8MJlwOqeMt2Km2giXwxt06mQOAV1ce32ecj21koXuaA0OzB7UwxyGI
aBCRCFuHL697R3XfgMtCUeVkTgA+3JOjQtTBOWpgQPvFB5G2JDs1HEjnguwmXEEh
hPfy74r3XJJAgz2XfEQy14nA68ZKcv37HiwO4atd024xQqJfypKuLvDPpTzoFqE+
SbcHetAhgGVvx51NDeYs0nb3HjnTpD0CN5kLXEDzpDubAw0l+rnoESGNyYbOr3TO
2lNJw1sVf1FIjwLxf7owpgptl364nxWcwEYiB7ie0YzBAy1MMfjcApQuOKXt6oXc
N0OoonAOVZFBcAoZiNMn7qqSBBmnd14uU0fLuQE9V08F/Ta3ShAghSoBdqOQ6k1k
hxeVAj3Wn+Xojr3wuF6MiL+3G8z5TGWpAbmoftuS6na9Jav2pTxQbJnEKz73CBfS
srUJnqdJ/Y1ndznNPZaEz+fJtHJD7+Rz95EhmN+Gn6jWn+4MXma8NRXSGbaG49ri
e5pLdcX+d9xfSk99sb8fmpDZJ/zxu71IPQAUiHNJ+HpwJ/pLZ55NBBoARX+rURuI
FqnflKFtELw0VWTDyuFRAy9+7StzhMNZJusvYr8suD/94WDvDbFnwF40AnPGuEAZ
PXPSeD6Syo1FFtW8PXskWdFbMsf0sIg9h3LwyKmkpKkXbtB1vTQ2nyGFZnwwgiBe
KjxaBFg4pW7lHw+VWwvHxiL/2AkOQSYFYX+eyVSh2CxSaxJZCXAHsQnzLChMF3gp
++gvjP/uGe4IUQeCn/NJPn9Qv8S2VklGA6bx+PQacI4J1BzwDjEWGn+ixvZHuwe5
0A0IIIpU8108pMqZdEh95ifJ4j+S3HEAZq6k07hVlZh28wo8JwihPppkehIeE8ME
uWpva1fRhH8D0QHh+HeO37OJXrH3Kw2ZKX3hyJwU61yVXVoHfB3NRKGTLmmmx9h8
OB9F2/LnjuLNT3z9F1bEqyMH61OZewwqIoKDes7sooGeh1D0j9I5I4VyB2nskM1z
RA9+6GBE0kiX/sAU2Cx8xhD2ExtJOC01Tj30BATA8csNqTN455qQALAfjVgdSz7E
DOYTAG07OiL+l1Kc9ziqo8Lfse3I9boDZp+i6WtQTpbBoz1jYJVXdp0M9O5mPXmI
gQxAS4ZHPtA+rf+s8w0Tth1GTDTl5b1hmFx7U1dXfWOLeoqAVftowt+8AT3D37HT
PYQSziC+rc5UxvpKyIczUNL6du+auZj6hYu48WzIiRcywmwyVuFaHCyVApUbpZsj
cqbIqRrx1Xic+AOuqC+x4+iv7IFWETqpgCvLFUOyE0IgEQEQ33ml2D2Gc6iLmUjr
kpx5wBp4pdrb0IQtUEGk1FOPzFgtNVV2sENaQxFmN5yYyAxSRjjmQ6I/xxMCxzQu
TPaLILDDEIp2Llm0GHXNx1Xc8JE4MTifA+CxEittb6ZkIqPCoQPJBOC5wwPZBHNB
fqqRaKWilxzDGTFbY+WY876CcLSkQi0L3QhzocAmucgyRQhmB/S49bQcxcqkyXKD
whdeF3TqE0btgfvtKHztc9aC6JosOm+h/+1zqX45Y3OJW7fYLunOAmocNAlXoCrD
7mWUOpQDfqyPF5UyNtW1s/DfpBordePf/nYJV4PO8Sg0aJtDjUtMGS2Lh/bofa71
MRSExe6GE+EaqeWKXdE7i8e2TE6QQCT1fMSyhbvxaJpMgSpcwlMqaQZrQGPn3xFw
h+Rp4ts++pd8LeuQjyR+KMeB2zhAz3449g2Bzy3JWojq6ME+DNYpEHq9AbOWJL4W
uQZgPY7Emg95znqydBfANbMusZ/x6tSYzlMzGwhX6XjvIM0aWOauMp1xlaMSKd04
WvHKgG1Q+R83WrLfLLV6zy/PDpoAub727SJ6tmk0XAoCXpiJj2iHdUjlgPvUqxnk
euQazDNlzVPDTJ/tbq5nSbWq9T7m2SCBb3iVL0+mPEh3h0/73jSSQ57ltqEdiZ9L
WcvkspGiSh6bDfzX9yfAe9+kQFp8SFnpA4WYYygmEZs0X0rRdIFEyL1TtJxyfgXe
/ybH334l72bnoGbpY1/ZcLozgnrrF4x88QVLuRWG2pbLiybWcmB7wkUi1pBEfnF0
U0iRhri0WvWHt0SzOQ7Y5rauz6J5A4IXcr1EByNDC2M8I3xkWRDo+jgQU4xbCq++
Agfuswe1sFQv4BtkjS8FDdwge5OGG6CObFoad4IhdvNwNF40ICfFtX7KfLtFA16Y
fy4QWrl4T87Stww9PKMPqnFHr8jNWKu4mKX4i6GBxRqhYuDgrmTqN0e0SZhedwR9
aYN0n/GadCH+0DkCWa8q9gw5JTFU9Bzkbzg62YNx8OKc5HRdIBTHI+qULtNBwzxe
2a3S+noiQJ6Gr4BYZIo/SpA7QkqSFJXb3G9nWT5fMl+XTjTzvTWIQoJdMohrTsDi
tpjhk7taWSUGppGpIHQ++eCKVqEdjwgPsBM/kkUNrcQRuGRedHxbugY8tPT35AXs
1ASkyA6jwDzgqw4tldmIbvH7ucBK+PmG/9hgOhj88ffTMlnpgFqAA/pnuhzdL7X1
kYOzy3XrqT8Zo/1CZ4+Kv1XK/X3HJFaa0ggotGINMxQgl4IR6zV3u4C0azX+2zFX
lHlTNHezC4eLalfjFQKSNpjtsS+lBrfQFV6p1dL9xcMC+PWRj9mGw5gO4fEUFyl9
Re8ZgDnVqVTAmeqh1Dot2+sHxV+leQItLEYN0YvyQg1Zj5oGolJoVg7JNeW/eeUd
UA1dbWGHDywuL8JF/0E6tBLz9j9yIzKS4kw12zRaRE8y5owIl4/uSCLUxzbzkvUr
5VSUajLWMobE/3aPI+OXoLwFF9U4T0B41J3tQ/1E23+f8nb3T8obixejknRTUKEF
OT41rzQNSoRpKY7Xhp1/R3loj0i6CGVz1oxRmeugVtotEqqnVoQP3D5sB7nvqHRG
fmlaB0W1MvM77Umt/FyQvTAGmUWKqCO6dM9EWR+/Gwumd/4R4GE8T28NVDl0bqym
nAgl5bV1HvYhwZZhADjHGAJHIltWGFvJ7A++0Cg5LZ4sna94GV3nPrK6kwmKMe0p
9NOEzlidltW+FvtXc8UMCL4IoUWZn31MtTTfBLKUIrj+rGKzYH/B9oHFS69G+B5L
Jk/TScfFUXB+jYt4OU5kYcRwSl+HjbU7VGDl3XeJeAjcrkVB8lkFk4V9LYOE25OW
TclRENx9mcIOXAQd7ySX3lT5OgBsTMp9Xv4hcbp0qXLMS14ybZ1Q6YW49D7e86jo
ZM45Li1GNfCCvZYqF/Uzve9g9u5upOp64zH3+jq0LB5wnDpCb2TRyfx87FhgaIt/
Hyxd/owAYdU1hd9pQyifmeeQuRcu2d1ki5928QZahjBvCBVr96QKQfW5TEXSXYV4
lKNv/Py6Citg68HNrANMlg027zG/2p/rbJi6eKWwem8cv6fkcf8UILDwVjc4bBsX
JWLSdIRx9QcK/Fu5IgJZ4HXt3klF6vx9cZONWG73kpRrzzhYBJY4lJd2AiYt6YO3
/cnz/VYvGt0T2QHI3WRmkB40B/6TZKTUpGAkh5mdlhMK6g4s//BilJNJ9MkLni4j
jkPp9KLTfCgy84BKRWAVl7qqsyWkHBD3yIZWIMtPs8ZYwf7MmffPzJXxXNNbByt5
p10+OhFVfm32ar6JHcyjUq1i9FbnF03PFPxTtjlAlc8KnqkHKa2sida+tyZFVuL/
Aq9u8Tjmsldq/xt8nVtddIPNrps6pTT4euERjLTRh6pYqs9eetkzE4b85sadPr7n
eUNMSlWBOvQWCwaoSbNXOw+738+UIH9JDOIyz25MyvN+cfvM11YYTmty+rslCIBE
yxGJ2OwXAK2NbSrVkUf0AS5ZzCtJvhX+b+EY+WF6Xam5Xs3THZ2mk9Sgi4TqOmYc
3c7mk+/VGvAPb4t6XlplZVEzkkHQau/brfSFXQYaM6TIaoWyqmwVdzUhytx3QHqO
QiAh92cDYPg5IctFIZy0dFR+dmCf4KhRsdaJWHdWra9HKc6fbaY7YmHHEWkabOVO
4CBS2swRoxCh8lb8fjIbV3i4ZZBh+CoN1uLeB4Vpzc2ox6i+enLpJ2209CnmIOj8
M3jXaiskEe40N54e+reBeZiJIaig90eOqOUvvtjQSoF5I1PYDvgagKej7fPnQ2Qg
xhD3DgSIVtx2TJ5r5npq1O4cCn6Qhz/P+Af0efbYoyzfbTONdwHHUP96eWLWWn5E
WVLCJMCzjGOmwc/9uMn4dxD7XRhOrRFFP8jHOQXGuOSF8Uu3XY0dfuOTV12V9Lob
xGa/OOjOvdeOoDS4nOsrvrxr4goktna+kyGeQqGQEL1Iuh5U13tF338slyBwRKDg
0f0paSjuhREtKh5P9eEpM19F7YuUNT7033qJ0tjxaKQUaSwDm3pToNHl6QXgNZ4y
ZRQVBBYWGbb8nxclJq1wplXvo0jHnfV64vmSPPL7R2vF7NCH/Rn6mjKIzHOOSY8M
kXz5Ee/S0Nofn9VL/ahRNYeMDX5ijl/F5kjqx+4AmnOYm+ozS70ssYbebAhwZWZl
R6Xex0NrM3X87wQFg+bDruDH8OLOJ3/pSaTm1+2ROME/VCXehbYjM+FBatGQJm4m
KzHza8W0BIWAtuikaow0seXtGAMu7AFi2fx5ZE2maILWWvJds9hC0CuZ7+erl9P5
glaUENJ5EGu8uYjL4bFM08NeNHIyBi7Jnz5tSMwG1VLGrIXv2yMfaeFLVfKLw1au
U3AMmLOhPZqh3wgYJtqegbfs0BXUerSKMAZ6NCIlj+JX86lRGk6iwswvaSC1RMEF
XTf/sRSa+61/xhXgsv3lU6BabKnAFl6FfDkGvXRpF7TXyLXiE1QFSq+JJyr5KSht
USFwmEpikinR2HaLbaXwikwfuDOogOYw+XhaVj2P3WhKv27HGa2JW6ztnWzIuDMk
Ct5Rkr2MhPDVrmcLgvrIPHmit260xqhUg8Ku+gSX9mISrO1Nt1tXRW87efCselA5
A7HV0WAPcpXYdDKuzzZWB86lMIoLSRSLys4YDM3B1TgevgKPuYjLARVYMb4Dfil+
RN2qLlxEwjKLDFQawqS81injxvEiObGYIWuj7xg5GT5WU9xFwo2vjTrkLOU1Iro2
dDfOLgFuHIef8oQyvmsdM5kz5QE1pWfyZCgC2hmAy0YFRsrzozcCabIaL7bP7Nzv
UTl7yQw1YeqR0tNUM9mOZoS/ZyNa7b5vGlBsKgw8T8m0y1bTKd5aZd3IEjlhQXBL
/TwtgQEhp9PYExT2QQkTvkNGmIwuDAlWcgkgwWjQzWBfamW3X7gtKrWZvNwhbnp7
FOByhXBqmDlNUIfp/bQWT8H0izefkbrmXW2ExBaWg8MssvdzlL8IjRgWGDfxZ3ew
2xJLVKugrmvOR9OcdQ2n3iUPJkxPu0uH4CwlLLF/VuRV5ypNWf7KieaQ6XEVXNrb
PvEUfR8zwYU/dHbyVGZB5lv4GcPh8WxbPv3CdE4QZgEsskE8D5BgqntjCuy9XOee
GCrDXYiHXpawzN9Bn6zxgswG1CZcOw15YBd5m4j8NBWW0OHoKTx1KFAAYFt9VKE+
T8WsWBJ13BvGDdHAyyIi9JaMO/WOseTmJoY0Us5J38u1t5+PtGhShzbb5m5JiJx/
36pe0EKjgaaC53k5Kp24K5lD0eS0yNpCk8pyu2byBDPbjf8auQdRGpOtH1icfSBp
aehbudnaT9lWb5WWY/bADiHy/l/qo/lOHBnZJSjdUR2wYqQRI8YG1WviNfC0X5nU
yf3Ma5RZ2gGpZACz6JRWkhL3gF+v0YR3oO12nEMn7Scx55KLGtdvt7GcUr34pb5U
hdGAqlxBLV1YOwJuHfrnfRhKW7c3BqEYQQvMQ6XpiLtIC0AgdFAhaGUuWUgwutpe
Dwr7bwHS8JqUnmXlwrFES31681e7R74wfU3goQsUHXwG22tcUS3m6XtP+Mx/Tm/f
/tcPZlOD+i+//S0wNBob9mmmZ+erBq4HJlej7j47/ziv3Qo4ISYNrqr0kLtEUWuW
GmbswOWjlAg206TWtfp6UOP4oOuh7/JTNgl+SIx0ocNuFjKfZHYFyNRNNegPTZ24
jcURcPRfadFeeYgR3vcdyNlIdNhc/r1gbD6pe9FY6TW7q1Hwkq46npHSd0Pb809p
6PZDoVeM1yWoPqdZ+vUyJMqFs4h4b+vkHOYihbWa0UUtE/oP2FcsuzEdXvRSratj
/fHIk+QHtTA73L1UtlzgpRwLdggZ4GhzLaO6XNpYle27KYBDLFkUTsrHmRTercH5
g8TB6Pr5Yk1E755J8slQPN48k98wz8r+VJtae3KVnfyHSBprl6/CdEZxE4EuhI2/
Qjby9+5K8LLtAT3b3tCimiuxQxvfqThYld6wlLHEDQ3XWdWVbqW687wa3K5tZkYj
p81ZV8eiCUR+ii9L+q3gBoIe8KpYAsTYYlas1vNWyCId+IPD0O3gzaPU5if7peF+
xeoXgOhPFqKePdgIDimWYrUX+mT+omc0t8IwX4V18lZmYwEOYF/VSN6jcbG3D6Bh
JF6uvt9asy2F6l64iwZo9yUT28lH6PZke2JcyDtxY/rxsBpi67VnVMRWVDVKNp30
aXgniHIXKzDDAMPjIO+/E81CI2TktrxUmFhlORkEOqEW1LohfM4wFp5y2tU6HAx+
NXD6zp+JIHhwB5b3YK4Wb936kJ+KU/chX4w6KxIwO7/kHHd1egRX80DW9MWApoJB
aYA33DwJAHQPSHOD0VLYYjmC8qut9dG3zX8WiP394U9Z2xNhIn/U9Gl/gBtTMNcC
CQVatHOG9vQVhgv2pG6gDO7dWwK9zKn5NhgGImxKltCG6oxlhHG6dFE+vcQ0AH1K
yMxAs4ZEDQyFbdrA1+KNj7AH4VEAZMKspReh8z9xgvCMuyQdNyV2YMifKMWJHCq0
3Mk5HDi7DXhpXI6whnVVvtZxaJB4NDaDLuy97urzQEGUZldZEJXnn6GwY8mfivRn
E90U100ybUwn9vbIGqD7lcjbj7bNWQFF231uhzC+Yqp1buOamsd3dJyiWq5cWPFC
s6ufqZBY2rxVQgzmkx0fj3X435+NmhcRir8rc8RN+k9WOpQPb056YzV1+YEhYufI
i4qthBpVk7BbZvUu6WK2vX+pu4wrGmALn3jS6zMqQqR6f061iiXj7nuBkTluqpp+
Ht3nX9uW586hW46dHDZDTqvhq6ncjHg9bEdlSCD6SVTgX1KZMOmGDXnTVFLGE2+d
jegiOOQHO7q5eaLbXXX4zenylnYm1wuBBRmMC7N2xrcZRsymNhwluBYnI/BpFsU0
BDx+P6JEXV3rTnRO4T/09SLuLamfbmotr4z5qocIgk+iX86QJVWsa3QpAT+Tibsm
k2bmcXCPL1oGq7NQ88u7SvYKnZuwKPlr8/gEMzojrVwG5LXlW9nDeYzLMEsRKExN
Ob0XyotXVIq1i1AdfPLYD1+f9UDDs9tzJ/jHuNhytmUdx+YY+vi6W2L7Ts8qGxgI
da4zTu88yJwyiyqhS4FTNJu0bTOalMNyn5pXXVpg2xlw4hl/KQ8G9CmGRlXcKN3H
xOJyhc9yPp52DyEVqoq9IC4hrrhcSvTW9wdcuEPlmhjnInIOtSyODPxDnRDx8/UJ
bFznjy73Jv1/vO3i4+P0Fjw76pt8BFFZnzpK2FniHhOt6Rgf5n0f8GQHbm075iPT
5GxVp0aCzM28CAo5lFRBT4SCDTniZWN/HQ7f3Q4BAP9ikIurVpD9vVPcBPl3LhZR
UIylm2MMK3Pt5OKazhYPJ5p8KssaRZzHKKHApf/gDC6AMxiwZKf32RH6UE2sNzrW
Xwo7s/Jjx6+42TjpRdLX7ZF6MoqMja6TsGDJQr0sou8VbuHWF9mUTmBk55MqvHbO
BB9VkY0G95X2r3gEiBDX1tW0QjOhoY8GS9fHXRnkm87tIHho0WWJNCtJeRad63KL
77dqC6nB3asTuy99eBGMKwausUsCSn/bXFaDpAD4+KroWgH3x4GOr6yZYvWijl3E
bd4DSyqyIcRXelC6QytHLj1wldlfEPZW0tjnoepb2SexewLHk2UkqXAA7CEpwv+R
nZF+w9ssdxMCVJ/CZ9x7kM2js+C3XVv2rXqsjSQYwnSu1gV3pE/H4InU9Y0EK13x
lGgux+8tTbUD5eJKUqFJ1R3Xx2Uv7OLelzNEJU7ty3tqeznO+HHYTeW6CZj/wPLL
rUSBP/BJ+27Q/k21jPiR4pp47IyzwpVXjlnXnUtxJ582ofQ1Lf3CreOicLMacZoE
2LYY6T+MIjDVenRO7EFVxgXrCaEyhs7l94nxcAVBS/rLYJoa0A+aOnLso+Ho5IjC
pINSpKDzozHxNot264tbbjaGrZLRaUjLCnfrwkT03zk7CVMNUR5Xy94gKwsqR8Ds
f1gPmwHeln0+LlbU7AWbRD8/Zd/NnligHRYxthKcuBJu/2pxoehE7lajliqmkfno
msOUH1eS/uvtYAezyUueQrTjy305hCw6Yolzl2A0xp1wHjIgMVaUhD9Y/Ha4y1I9
2SfOeys1Kr0eJyhl5vHLEyZnB/0DX8nBASqHbsQhXGB7uM3QpXP1VLyxA6PbXiPG
OCss9eZOT6KZSt20PVxaV9CJvJAWlo7LuuHNEcNc7JGWprM3AJjWitlFzKFn6E8G
wtWwguvP+QVUjc4412iR7Mpj6OaWkvz0vRe26+JVtObMzbs7NYdDfxE6Epy1PYR0
S5lhBSezgldC0ZwLjOO9mxN+Yq28G9R7+a2Ocn/qBPzToxBc6RevCC46xdMc6YBl
tUiUydEjRGc/pQaZPaV/Ipp8MfSnyl0vo6bJbe+UD4jcjpPhhMWYT0gnLlFQEUAN
1Lm2kaX1HPPCMAqnmjMeysySVx5B1FLZ5PLEFk4ei/e4luqaPBJ7MUHaSDdKsH9b
9AwJA+yL8fjMrN6ewjQ0POTifcw5eyjQQHT+V7SZxjMn/OTVGViLt5/fR0cHWT8x
KsYP5unh0E4EkSkX5oFYjxEJ5Sgz9CbZ/on8+H/r8or36K/5VrcarugbGY5wnkbn
ls3LNGqgVBo5tCakLJAJjD9JlEPduGXA/Q0sM40PvAwweEx+cxBUl3PvfX/Ixqxm
8C9nj7Db+QKX8V2jApx+8a4d+N//vL6byjvFdWNgykvDjsntz4nnpAtctBwtSQMj
Y8sy1WzY+lT4Iz/BFmSeTwbA9ZQX27np0Ty13ZB/8bvbLx2gorw1pNxSUiqOPoF/
4QAbBB6suKF8UuMEz6JIgjbhzxbqL1nOLHmaNo66zgibz3ihU+E3rbjgjEvZJmNr
KJD4Rp3NmH5fIFEbJWXjOqbcKKKND4OWuJLiNJ2lMTAtjQconqOvi6JZZO8qOTDc
zhfQePCpQMI5jgxjKrRUJaZ70sTl4rcdN1NL8BvYwx+uNPJC9V3iJ9LjGKcM7END
/MVZxTXVE+Iww0qWWEQxuIsDqZK1WMbOKuV1IRwkiKkioPUt+PIRZPyXe1kSfLhi
yLDdeEcywLdgN0izsrI01wv4kZB27auMpN2LT+xJ/6yamsUoRktgk0SGMvniWcgR
OeGkDWtU8KNS5fYSp9alxzPct51A9gJHTGDKtigLsECwH1RFznaj8osrAYXG0XnV
5JAsQJMOIsGMn9j/T4mjzLzcs4tws6B3NDXTcAthN9hlZGE7GpPUXyC99x2eqWGN
XhJaiYSYDvDbbAnGJauZSd1gDlopOpMTs+RyaTVxY91Yhq0KOYRvAXy3fyD11Wgv
6+Ld58aVIVcpMjm971qoezpVjuwn0qTjTZOTd2tZdLQJ9m8Akjeawd80VXtGC6ck
VjVJM7u9cjtfXv+LKJFBwXyKjQLLjsAAct7lKAbR0e964UDYPmV0hpBg7J+eicQb
VPKPwVtAH3Qi0TKz5ZrEDOekYtDG013P12FTfbQfb62YK6Wqz/Kb+UIMjNJAC0mc
4gatB9aPriWmKLYwsfSgTUypimJ7ZMpglrc7V2/Z4mLPkUMyqk3RflK9BUGipCEj
spCzgjDlX6WnLIQcn/PRL4eY0o/7MZMkUOIr75+9r0HLT/LaMC2OK9Y2P9twrC96
gEnq7UGphfRIgrT068XMV+Lomq6LmRKsIOUT0PGVgeGaOl3CfQc6yQpbza1P8b6U
v0I3/NCMFDPiRdXosIqD5INtJbzPSJwAvveSrHXf7NL6+YYLEP4E/+/VqXdcZ6u8
9s7y24h899ugpVhGPBFN5oRRNzYQOsx/U4IVCzIv6NcNXu9GS5UV4K4LfjaDwTDV
DlNjDPcDnz01sOols0e0ECf7RNB+rQTTYgmPYIxoHMBp8NIJL31WBVy8jKoboyrt
quJ8NYYucaMtcYzzE3g4WiQhVe93ZV+o5r2tWKWGpmSrsBD8s9E6BaXw7AzyDBQa
1QBlRuuqQupC/2V3T4aE4Dy35J3CCGmwf14kOx8czZNvjdOnfrWaZSdLEIeDttIb
J5yOW3qwYQKDpnDW1mFlw6ColZ7lmHtMDiylgiUo4m0xboxhE2KQCnUiuE0jjxdz
ff+E2hlzg8MUpTDpjmdhJimNacfD4MtZ5IP6vCEjxy4Bb6Pa5k/II+Ub450ZuDlO
irkiS4J1IWiVhKxJqeDp/S0sle9Eu0wMTxMM/9EdSvZB3mR95vFfQPApMf3dA8As
Ft8SljgfGiP7VPs6V1aoKBIDVZ+NO1cZ28h+P1kdc4beE3rM+bCmBDNkAryWX0Ce
yOLEHypH1IxdwWB7kxdyVaLXsrDC5flP+J5HyU91ovnUdIBmDjUcS/hqxtEoalkR
wQeHkcv0lPdThbc30SCyLMV+T8rLd9LX6ix9n8PS3fM8jT/o5nwzWPfAT5RctxhW
oB1DvbLI0x4dhUKndoAPLTDy9CBFz0IMMuwbYLB4KWHeanhqcoDdpe4FRTFq5+rj
mlvH68+5SAMnCpuMdWWypIQCT3GLYcdgunuhyZeTfd49FeAqL1zmDJXEVWVAh8EV
9YbAZT6Z/rFTsmrRrsUvk16MIz0NuWWsay5PEKJBnjIlutyT9vDMQRwkiUJbr0VI
nkvTCUmcORM7P38Fr6zrNd4yYKeBxfupOICKcXXtLWpGLqvfaGlysBxB6AOsHvAs
ilgL1T67P/z1A4x2rh0HpfAYp/ethmEU1fsoWZVcm1qW+BxT8kOLqsSHlZHVkMyb
7htXq6NtB/96pll6gBDLIQY+lVpJeCwjRkVYQavTDOryMGnAH0uQTjfaDwdXnnoL
ZQLp7O3R4FPQMeW0aivOojJ9945yyOttO3jnOopHwlBqHtUNcP6jRrcEJsBHeYtn
MmKhTZm9JzHZ6gt8W1GaF8vrX7m5tWnxrYDFOd4BMkxgWW0RWUB8TDKiSMONXTGd
0IZyugUE8XKRY6QbQYhwf93bTbJdlutcLP2DBzLCjKP1GBMDHrude/bdmeYLVTpG
7FroapLGbo2Si4YQZuwd6n74P8M7vJQx8tU+lOcY3o2fpbfICM4pbZvIaSPeJiUo
tfuUKoTAHQ3kTOI410Tzq5fUSdh0Wfg6VywNTvTuzrWtQnO2UozQtlSwmzSLXugd
GNWiGx6yggsdhcGcC2TEj5N+fJFy/M3244qVWY13pT0+TwqrXDlpoTveVd8ts8/e
YMdJ66bvezNJnAoztMsS4DAJIaujw5S4zssZ9Ui8W+waTgknoZ+7xWjYvjvDnJKH
NnqFgT9wNDueTxY9d87wvcg5jNKsFpRPypDBQm4zdkBW0wTxw1DhX5Tr2VouY9m1
b8pha5hYn198ERknecG9Ok9WXa2VsOKNzfAhxoP+Hz6eQafCnRrYzruemyGBrR1A
yI8UYMAw/6rba+qMt2205PMPA8x+cU5dZE6/mxNf/y4qOkZ2wkyZyf1FFH66leor
tmdafiCZ6g4xpWBAYX7RLS4Xo+8K9CPntSggvoKze6kKIgIS71xlcRf9SLdEsyXg
1BNxP6SyH9m1OvJRpXa4Aw7W3HuQ93g5idIv7ykNrMlj8StenHTdxJUk3rX6ZpBX
uK3IutZZC8zzamEuskdn3fVpk7Lk1+9bgkYIOnRj2KBaSbU/7dSH4lgrZ137Ot0T
yXaIR/2cl9REc5KvOKVrKGfrr3W7ymGuYi2PcASJjrK70FHzMp75ED169p95KJjZ
/1SXlZRA620O7jWSC4+nA5r36YKIXDU5jqSHtviR3HNuFTm8Ejme8MxaNBfxNQ/o
Ff9d0b/i5cAklrgtztUN2sKqaz5FaSFNYjd/6/EmjeW5IMLVKVOtdDp4oIpFPYCK
7ezq3+/5EzuxJmA1JKA/AZ0ugOG7KLRgJIviXKYYdq+WMGDFlVgg6kPpJewMrYlL
Jul6Nyn7KVZMC4dWmBhJ0B4S7kWzPS/cTh9zwhaEbp/GwFAPxixzeJ9d7yj1InLB
iom9HsJXz8cev1pjGf90fdV8zAxCHXATkPaVRG++KC0Q/0m+kMc+zmm/KmDGQszN
YQyzSdH+N5g6N+jX3Cj4AkeTIEErxJ8z4L03oSCOwZUk94i1FWBfyuB3oUuyiX6w
Knhg4xCIu1w/bOV0x85UXIgAqo+4U5yRkA03cfT+XGbU9AuXJl1lq0nSFR+qRe6T
vzxkQsAEX7brxfAYUdA/bKi3o7+/8bCN8wYXxBdm6/Gyt524uiLhIuiBO8jzWLAa
WYziY4QJ7cq2/mi1oQS7zATK/DOUXG1VAn0dXxjHLqGyHJjhUqEyhCMiv9zSIz5I
liszPZDrXajJZ2rUnLBSglJiOaCF9c4jjUbX7dDFZaZeckD/g41LFDBAKMu2bEA2
vNM3JO2gdjq0WDqG04pPM3PGuFeahQm7+oKN4cp/vW4tgN8Ni0earhOV/bc5p8d5
oPQGOlySct9BYwr1cCiJWyAQPrwwH1U4sbaRUsIML9kfJeZIZh9akEs0cLBlKOsq
PAy0cMkKbNADfQx8QFbjibDSj1ANumAiMgW2UEXf+Eh+dzZQCYDsS6wdwhO0xWJV
0cbc/Zeb33N6P+8Gm2TUQXoAfMR40ObCKCEUL5FdUMdElXqcDzMQYnB4tETvoIio
LhljbkmNezDjwHE3RlbuFpEohdpVbyFkUKEWepb+kkoX/RbP7YYiPVGevWJNSfJ4
yci0yXy+y4FDUUBhOgk0QJgr24mZaolBlJUGuEplJq3bAkBwgxaO/ci38cboDHKv
066s3erij6rvPtS4fNhDgCOMU38xFtpKre8i3DdSuc8c2pe+gut42QQl4Xx5/TUe
nChFUv3/mEItUQ6XTe1hJLjNP8IZsb3M73duZBWSL21M4bvE9Eg6gI0MyMSL8n7X
MltTJWNP/NhYIYtuhaX86I7fUVMyxqsXWsTQHCdMkM+Cr5QWjXN0tv8+cGXZMzcF
gxwAiWVlDlkqp66OsSWAs7O3BJW51l1nTjDYo0fLlaD41CxoZ4sridhx9AU16WO/
8u52kSbMg6tp2pzGcHjPxowq4VlHa6zODZpFcqS1Rw46xM0vZijYPo1osSObwaZF
X9IWLaqSJmGfJsfMeg8GNshgcJIIVHH8eh1k8W/j/Ql/mRbzhFzbcnStrhTdpC+9
XO2HijWwDkpio5QRavHLmeAe9ZvirRJvCbZ6FpUlJ36cnymlwStW5dybyo8DcNbW
wB+GSMUQVr3VUFajo5VN+W6TzliTlA3RfaIzqKk9v05fNh3sDPqggOiClWsgdNo6
S15Tv1EkFzRn8I68xdGn+xk2R0svML9qjDd/i9xjoB4+fuw9DHlXod7Yiuxof73Q
k5pQMRBOYl3YLOBSjbGOhw6gE8M8G9xDMa6nhA6rsmFOEgTuZ5aljwmY9Sm2ByrL
SSC+JyciSLMxleOmvwGnKASNdL8iBg7bXL3zCywMyb1OM2JDHxzrhB/k5IB5DDAX
xgScl8eE4mLJ0+i05UpMCzDBt+NFa9r3Ox8UFnYve7/ofmRZJ4+rCFaPbn7v6QPd
suVfm9QHGnuqdQc9QPCsyRqEvnFWKr4uGgguv1Eqh5BO4OtTQJZ8E9E+eZBaadqS
/e36eD7uNizjeFrB0Sjrk/rOy8zeIR7NcmqXIuGy1mnNFssA5Zj3yrFWKBMEHglz
caOgT4qhfKK/Ka+bKWr3q+zoVbWcOhlrDvDKFHv0UZ12xTBdvXxpIfBymF8rH7f+
S6b1oMe75cDt7XmvfIWJzsjfCybjFpsO67hx7BYsNfaTe7NPxbmWGKSeoDQ71EeR
Xif+DJFZ/Ga0+Sr2vPOlLxabDvOTRUE03vQebzFzEas17gQkrHaRxan0wRpzY1Pf
vdPxPpRPrpPlXHp4Lc57/RHbklSD36sIgDLYQxCPJpN2/fG6+y2KeV89V7TajS2m
bMoeqkOvng8lFZu779JJFv1reGUlEiE1cmLsuuzKIUHEEzRnymnsfyfLYjY1tgrS
1Zt1a0+uWYpQaptAoN81i1ej3Zuv5TDLUyi5+XPhqSW75wrvv7LdZmDdBpj4/eCX
tR+dsn9s3NK0ChOg9flT20s2D45jvkNX3xaNPh9rV4pguY3i/BIefhuWUkAp0KET
11tCm48xleDCP2/m0EIYOtgyc2nqRZnEWpH/aZFrygSNCIWfR8+gDCztoLfzeFoj
2C83jc3fwomjq9dVnpYFm1qP9EhWpsuc3h7EShnHgJgaxuH7p95ag8nNDKpjwARz
5Yk8R49o61xhtrW7VKx5S+WxGnDy1xamzS0OgEWrdohxzoR/5eklB5kiZdMQ6F47
wS8jIEilvB6+JSO1vqNjvkTqJXc53aLWmo6PXQpfBDTxM610gj7LSMNsxproXPjL
s7BZk+0xMCXl1ofiq9fw/MUsx9QihXoChBirFgWz98Dxoz+iMvPQx7ZZEtwZZd98
P2zRTDtOCq6Aldt/HxCJqPmtKk4xaB8yTfBOe+BA/TkpJGSKYkr0zeKAtyean4c4
4DAMxswPA0cOrWx6QcBkaHwNkcdGhwlr1f3mtwZodHNr0zYHNb+tIg6gqbug02nz
LiMOh1HE1MIoCnOiq59XJlW4q3STiTY0dxiuN3SHWzVCd4exrmVtvdX0BvmevXXX
zhImceOT/GWiKvuCOuMGtJUyawKsa4M88E2bCtfwOs7X/OPBajcxvh4TQRVttCZZ
6L8z1Lpq+GAv966ka9CaOWJnPG5p21YKZDAYv6pTA8Cgt6xnkRgZc5tgNToOjbWV
5W2qc8yuUYyy5gUvA5ytnADeR82kMB7pexQAgmoHAK1ddw1GbzIwOJVSp7EUPESl
RJBo320fz+8fmVaBEdAZVjs7tTj7fTkKZjzeKThcegE/Xwfy4EzM3S5M6E1C2EKe
9tG0Nn5q0n93AfZvjBvJeYA6jSc0Lywgs5moiVl82Djv2buGHyESCvhhx9JgXlk9
XRk6DzLslQWJWXRq6b3CZEvHHIkC426qikE2IhhZJms8g6GkEintaAvFAt7zHO75
7iA6Zd3JDEAcai6Thc4n7bVul9Y3aAJaFSU7uxTsuqHJ+WOdvcqTR03c1ib43TO8
VNdiNBnqXMqgVt/j1WlDJeNVALr1d6HbKqnpik+8FTLsQ3QnRAzyeKY8lFrDNvRc
wKk/R3hdOqbSAPwMpJLzlepLM7oSJ9sLBHyQ/sTVEt3Yfw1xlGdECsZ7kogYrhEP
qCxf/29mtT+EkIqbDidDTOxGNCjxlehydZd3TiXT3QOeT4vF2M3nevXcRHul9BTe
Bsp8r2GrIBCsIXv8lQXMhupEkBWd/sA9cWPR9nw5GO+o1LI33LVcVPPGbCXWML8o
CaL3Rw3WbSKnkIT8MbSaOWM3e11Vz5d1Q2qiqbWe2ERTp8cwSnvRojzSimK+2/Ko
rnLlTYyLpA5ZPlUjBfU+Y4tMu+D3cZKx8Zm7KDVuOu8An4O4Ukojemt2jezoNDia
kePiEJL0jLqNhubeUQKSIaB3HY/MXPf6XFuNgjC0/Dcrqlr/h7V83GU785cpuFsF
W/Zw0fKZ81EmymlIxJswaR3vmB07c9OydEY3Bs+c2lTjuJ685ybgFcxY8BZ0VSW+
zuZ5Mqx8HxQBR2kQQsp7t5685d7bwMkXBp6lxJpgqQZmE0W4bgEar/zIa8t+Go9F
aD6tuHcI+3By3f+UCZutMPF1IY3+5ux7USThE8ugnjosuuKE6Odepok1/d0k3Doa
+ouADvyY62Uck5K/g6i5HPvw9VjUKzlnU1LcqwbwZv4ds4z1wHsEHWDnLJZU9oG8
lhmiyrwbKzlro9meTkNZF40FO31H10FqlaQ0sEDS5VuVWdUrigSuMRlGkIKTN6ZF
Mhxo3GJlsrjx3PxQlmeORDm4YBh0S+biNQvsTHePXuNEwGq6woWEYdijEn03UKAA
Gve4io/EO2y2db0hD9RwQkfowbrMg9ykdQDwfDj5M8fBlehXZCoIw0oBeu1gfFJ7
F7z9/sZECSNZaXKyaaf/8eM1mI9MtFlv9jw+K6VuM8+apgk4al9F1sLwggAApuV+
+tFSH4qC0Btv8ABkGlbumUisLA9P0N+eA4XToUQIo5OMDQ78UBuYXm+hzdsEFCiS
yQMCBKs3/MhrHQPY2LvkCsfC8Kz5ezCP9EbqTrg7R2mjWmM7gn0T5PILKAFqn7fx
Yn5AjY7JFQl3ObfCjrhpHTnTSxydwnm8+LJear2YtscLwuYTAbXRJpRpJFQ8ps5G
2lR4yczTG67ZjpltpKiOgV/JwtTLc0BvKmxJAhnXpde3KvA3clzwXj3dJVDmz5bB
OoI/MGOxbQJGf0m1g3HHXNvbFQd4m4keyqpSgrpTdiuOLrEP2tcgQRdX13rDmg0P
SCBQHK09cR8qbjBIJHMOMcI9pVxVan/koLhSMr4kkNLErDPkSEPsTdbl1SgQVqid
6qqWNl1JX2Ub/ukRxS6RGsoYBQz6axz+j0jZrTKSfEBKVX+f7YAzdZk6msxjEcpO
DCTqnkrCn2VhnH3wUJUoO7E680HSqgd0vjW7GwWStu/pzWxWOaWdLyukXY6ka4Ml
bqXIt901MGmYQ1nhoE91trYMQOZRfmN1vfRjrNazrdkWutgTnNOT5e1eHjoQ5Y4F
fdY+ZOc/3P1Uz8TTvUTI1FkYvfRvl5kNsoz5h7kB9v+Bn6cv3w90HZcV3f/fs7oU
Z8yUqMGF2XlLjB0zzwk5wxvxt5UQ4N4/VbjV904glEYZoDop2115ZVUL9cWZlmAa
zC+FWkH0KPo8B5U7GOr6Em+e/sNr578Qu0Ebsgi3yo90yYGjJWHG7vDRPjeL5e2v
IH/LbMUUxCBaxpFX746ujcYnvbXYtx16osE5CnoQmsXCc8IMAJq5nh7c5KU2HAJS
cZgIWAAqr6I6umU+j1VV9rtkGgfsUv++jd7naWNgjnwkEqWS5av3iZc/F2KM28sW
i/Zjr5iR2KYlQSiv1oqlu2scz0zVUSqYremNvnLnTa70FLj8PavLFZe7cj3v1ZWM
Tl67Q9/8tLalIZNPyyLWyJsUx51N1RdpLE43rYQqRFQIhXWVbc1WHrI38rvrNvxd
jDEwioiYybFf71z5T/cPgN7IwhdZl9rl3QW/A6odgP2EKm83/41xkBg5f6qLIx2J
TyXdc2qNiluvZT+/FWMQTAGulipRIWisAv6oeJ5pMzGFRYXjU6b2TswJRMKU3/aA
oo5wRQsFVNIzIrRPdE/abVjfKlyI+Z0nmci7/intQrU7gC9eRcWpniS36sFyhkng
UnVad1p1qCe0YBpQrdf7SO18ga7QurxNheSZH+mTmm4wufBrj/Bv3B49IJbAzQDC
Zr/ZO0QK6kfYNPWarFuaikImag+MQlR05aAL44jAvhU8BlohdF7sSqnmGnxhrG+f
BM8w1QVBvPvPZgm3bVEhAY8E+O2N536cTI3EZ28QK9V0tlH+UtEm/UgIKVVBo/Cl
ovFsKbqX8qMGqF4y1FAfl+Mu6leDiQOvuhPpyPG9h6wYDGbbAx2N71rpZgj2zWP/
BdItjMo/B1E2/mTNAkiiqPVuj/lDjZukrwyv+snZbdNAvGUQ8LDc+YC5s/VaS48K
ZSTGQ87Hg97EBLrsHxiZtVRNXFmq+sfJWcoiYKmDfyLcep91ux1U8NIkmvxrFWuQ
TvhYS92O6o4cFYmtMWgPijd1bDzP8dsrKepr2HTg2X7onELoLrc1qRPMlPO8ujO1
Vj4e+KKTLmr6Wk4qTOUIL2phWsJiutDVoIxJi5dLVGCQU95xzdD1ySj7rFwgvmx+
AmYjiYuJ2rlp5pC54OiFpyFqI+Yac8dy9dTy8pOEj+DOebT53WLGtf7nnyJ8J6oc
i/2Njkg8YSsRuCN96zxsC7Na1RuqdAGliy0UxEw3kZbzh5+/N8i4LrRxbKvXeDek
kkgWL0T0PeBImQy2whWhz67xz2bXz01frWTFUv3oU7glV/edTbUkI3TwAf9GsXPq
iq7vqXouipdMvICuuHs9dkeVQ75IM33SHloPozRQm4ENQ/X1u+e49f3fw3P0POHG
4s6z5SZtYqu3QQmgRXyH5+pNvfQPT8/Qzt38gFkQvV47NQp5raanwc0zkhMVylmq
zGoW+ZFkl6m9mGFu9yPuw2p4DoHF9+7HLForq1g/4OIN+L08un6jyMnPQjGqxyb/
fqxSYiHTf9x5GOfsvTOEmb8167WETE5/lvAcsaPZuwSRAc4E7CPe5soit5HuSoL3
HrCZvNx5cAonhEvfscZZs9uutydTh1EX5A113V0dQWWk3kn1WKE9k/boZeciiTzf
BFk0NufC+MFadSvvu5+e7MahNoK67MmTI06BLslKYPeTUFZfs+L2voOUj4yqYQxX
bRGhUhyMwFwKnCe2S3kn+Ps0Mcfz1lKGl92c3Jc0Nb3nna6PclhmNxzilR4zrm0b
2U4Y8MCdnTSZM5/32WAXsmIGgBLDKVOTVJz7mRVu6bRy5tgO3fg2dFyMldCC2oGP
YIQVbBi92MhfsXWm6RetKEmauAs8S3atX98fLzijzkp4Hjt4EROTxcnY5Ba2R083
EOGny6JHb69nRNOnud2GMQLe0CdKxkd3pcq+53vOQRCSB6n2b0RuugeTPIqxzB35
5kICaW1Fz16Yi3SHUx6Y2SWGPZNLlSen4LJFu+X7/qh9wEIbVllA4J4V7hsEzGql
nLSXeUirZrRET3NIzuq2yw3ImCfBoATQcglL/ujsqspeUcuuCN9zUwLcTwN4SZJd
tBVyjmQCIgEr9yAnLQfZssR01o8Mor184bJtF/8ylBorzFxn9v8eqiYcD3RUQXS+
kRgE0YZBl5KMJaZ4YLlcVubppB9smGyJbdMLtp+SfZ9q+b5mmQSKPR8lrZfxYbGN
S837763WiMQ8Mz8/9mauzM/kZ+uC+VjVBVW9HY9lYnbGnqtYYNTwKyQ2RvvuPli5
b/q9LaNSka53u5l4eNu7+jMkBjThm7Xmk1qh/tYoV0fWBg9WoI4BSZoaISx+jOtt
NaiyejfKOjcag1bLVusHE02fxY3riRPVOQ6dvJGlw4Ka+CYauH+BJSfRKNOleLe/
TxxBA65vrJgDvxQPrc1mQZ86c1ptgHiuyepS6dPmamkHK6NGRH0zKlX03pMQIS/d
LCuYyBTFXomXPwShI01lWfkWZ+zEKU9mFsOozmDgGtSOdw91sGsXEiXxATPKlvox
kA/peqEwqvCJbfecFtOP0zgpk4LgM56Lmh13R2VPUMmtR6cX1vXtFDeeRG89UGwZ
y/X6hNcxWOb7Dj14K9BPfugNPJbNKtJEMrT7vGJ7rkWGwpEuKhkQO1HRDrorsZp9
X3EtF+U3GOyCbT7vXt5EEOeYCbE7dRZqH8mWjP0gk22fIYdc9frohytOTuShzv1X
Dc7it27pKOx+eoie36rJn6X9QROeULuQim//dc/QVEK3q7Fo8KTRamABltdC40kW
OcvP2vjJUYbnad4ZvL+AMWW/5rv+rR4T+C7xIRH4cnxbPSg8MAFceIVC50tIktu8
ZbyDYjaRpCjtNF5+itOLaKkXtb93jJtNGWEDvDjP3iSnxjWrEySXWM5RAg2pUeV0
Ryk95HAEwOee2QJUAMyi3XWo6Xbotz7+3i1vNDBfkBE6a3RxqX2mnwv6MkMGpuEV
lQ89DomBAyNBzr+f+fb/3fqIzuDC88dDwToiwZ0KDNl014KQCIOk9XrvdbvwilqK
Xf7G472ODNSwUI3sUsoOi33+tCrwcjtKpsiCMOPb0bql9Kvy7v2rih5l49HfXKBC
oa+zWWdNmeZCZ6QtBGtmKBJcm5g6zX8fjUkbFQecf/pidQGVsGubIucAaP4nnMWt
TUfmuE5+wWoxPm6Q2aml2BkqH1TvpikEP1hg7/8YipjV7mNCi5GWwCGuHH26UKOh
3t7Hn2q1Q/h8p8cJPdfv7FSFq28xLonKLl3/GKI06gQ4PAOHoquE8bFJ5CozEwUP
uGU6+KG2VqAE1YBVQOzgd2R52yd3jn8SEB+eqtfiUhC/J5P7IoFbGGUbA+vhnjnz
RyXpsNZl5pcxMahECwyCogwrBRxNgFNq7crdQCARcxvOX8LW1K7HJYWjlWFz7b4i
1zB5vW3bXkBxEQwC/2xtz84bcf7AAeYX8zEIzK6u7uIsXhAlmWcj9VU2eH69TVAI
B5e8QqgnT+2gsDmkvW2YBJzJgU6hifHCrdx/ALxEimGKahcKgT/pPriYGexrVgDN
212Dz3yMm3mY4Fj6Qma8i7qoEkwuCgfLORBlNAcHyUeYzmcZg7OGjZE4467smFFL
1O4GjDwGz6QyFR4RgrwXw2rP1coAmLauG8dzvGcRrzxSS+lRwySKnVRl9q30g8FW
4tBDEdESxUDmpet4sIM5RpqPJMWa+40Gu8IKmZ+Bo1Ptqf55z64HOPbXI1dfc5oJ
KNylRQvPDaZXf6OU9rbjMOBRCP6o/mqyuC6Be8OfFhx4J25lboUpBNsTJbGy4NLq
il5Gmcss4J1QQxbaX/tn5yhHPVMgeeGfYrzm2PR85nlEli/xQL3Q0wsRy6NXE7rE
VAF2y+O5OjyspAPnVO4DdM+bEuYqGhgXEKrPHU+Xb50PzgEQy1JZS+uVQ+gx2K0E
OtvAnnlb/ZTa2LlH98kHEpIKGXzEL9OkUZ1JmSsj1CCdAgddzBXq2dKdT2bL6FVu
i8FTxuzVmi7/y5QhIy3zzP1FNX9hycd1NgMWMyRYCEtFVqc7D1lwFocJkzHH4gZs
ZScltdRHIP+pLh0B8rsyhErqBcFHrwgfVJAW9EFCkWwzU97OL9w00dVMr1IDP8PK
T2wDpOJlR2A9/XRkqle4xtq+viPG5E+z23RFOXnnDtv/pI9RLkRSx33gKJ+MHljq
CQwPCi4QBW/W4gYxD3vmBiWGnhy3ITIdzL4SkaH3wdLy4C9KyQjbtOs8O+gfGWSN
iS+Lsi/2agxqKTj6lJHQo4QqzLAaj5JrV++voA1o8qpXI49Z0HcPOPvJGIM33BSC
Bp/JqFhmiCOBDKaZ33IGkpEbN1rVqVee26BbyqcEhCtTxBkm147gF21jqC4U9S4Y
r32AhFLwrX6wyfrEOUkjIpRic+LXULDoUytLK9keD85/3Xj5mBSNwyudV53aPxEn
syGOyu1eWIB4TxDUOa9842Mg3T+T/49XuF9g8SB3uNedFd2H7AD4EP9GrT+S9cvG
ic2/0IIJBGep19n/nFMH2VXgyIkKpUAgRs4RSrB4FqqWZmZpUkvxhDeqLJwomNoZ
A+FetIyccLl7ucy1yr/PB20gR3Fn6htdeLiM/kEUFiF2w7fAJtL+WszuGKDZOgL0
da1Ese1Jo9cubJzUH76IBzBDb2sXD2bCrjbZMSWP/GC9Z7VJpEIh93mpz/7Qf7fo
Ui4yXXd0JpvFQ2JpVWPtcdKbQlJZZjqR8OzQPF7fClsoc2MqtzZTPmhZn8JieMfI
pSZhdctkJhzbrbCxMGGcBy5CnxYXHE2Qz7zahbAnscPRv1J8rweb6tJSCZYCdt33
B5AGsvFDpvHHndIume8Mztah/oGjHeOC0bbfta/6qgRJSfcWMy5Iu8kz/tFtkxtm
sDIjeG1ZYQ/NTcuUr62IJG3fok1IQNR/a4LYIUk0jljb1m101ButtpWVuvchQLAE
MZs+7/suZH1ztNGjJjQv3JHBLyHQ3Rfdnmfuca3XMUlh4D03HbARIu0280KDWk+H
U68rniu+tPFnc8IjyO/IiKghWacWVWuNQS0hOLuZrgOShyXMtrdJs+XFYrimHeKx
3/ur4F7UUcisgIHsovdO7BQECQmWTfP4eoMkvDtR+18AKVGrjsZhYj0Eb6r36Z6y
bNsqHv4SLgwRANJzqsaqo2CGvw9CgVFLdQsZLuTipoAjbye4LLHTYlabmxouUOP7
cVu9fTXxFLvS9Aa/tI7hfJHpqqGTqPBhIbs4fX6yXrg7vt+pnvv1wk+eVUhe9bFB
J+sxKTfjnseb4Y1HC9HdopHXeNUYE8kjeBIAsqQvwVdsGI1uFfGBOXQ1Aw3mRZ3I
QiZwgaP7uN+12poRjTNbfSIEGhakOUutKMi8tfC5EtjXbzJRoB5wyiyl/33j3j8L
KAFkpRWTgKWh37EhdQT2LyduJrfr/uROwZS577TwCgyDBcBekkYK6+eCB/KV3yVg
AzpDXKiDWPK8h0i1888QHpWxBFMfWn9Es/EJAiBb+fnIAX+Q+p++Y9ziyYQRgEiO
sgVXiU1F3KlINFJq+Qo6u5H+ehU7KCfO1Xc1mrHXhm/I5zjRQsVMN5a67ZD2WdXS
QGnvjlWlRZK5bL3SFj8er8BXq9rSpBLQPZCpRiTzD2A3ae3+407jA4tfLk19h/+q
B9Z7yb0x1ZkgtxMMEdf5Hc3m63brmmToCTrEZ5jM7H3XtjvAzHNFK2DZUNxi3Kpy
MyJiF343R15OG1WN8kFfRxOVLeTAok7d+fmgTIty8LktCMMYhvJaSqHbnoSr/QpQ
ZuX9+nsJ45xV5q3l0MLA5m66f8Wn4WDgCRZAr6TM1jqZvU8nurN8uws2OebPyaTR
J1GCzKieM6xsv/thNurk6qGUguWXJfMvH1oMmrJIr6PgD+nWCwVICxgw5DBZPzq+
fuGqm4KjUkxX732S0/DJCoABL9rcpEwWFDIu+6XG/fYRgJfjuZNrnpDbZlpOm2Fd
DVkIsWo2cPvVHBraMF69yRRkQrSCb5bw1Z81/Gug1fCjC0vEqO1vl3zhuLZ6JCpt
pjKwDLC1VdQMl/0ZAts1DszMnXRecZsbelA0AkwFPFEANDyXbKo7sRvtL2fUw4sg
fuQI/6GgYA1NARzhOXb5iDbaMKl/6Zvsb3cRSh5AXcivRscreCw4szanAw28hOFB
okEuhLkq5WVPLmuSw2tHT/4kKz7yZsQ3aAoCxCOsWhWALkWlWm46UjezRQZQpBye
xcADketcWm99A4PgHCjFxhRfJjpXGxXKozCu54RzJWuiCfWrjgQNizw2FjfhzUfS
eqTD+JS+q781zuMdacHantmLsZ7e4vLFZaUyjJ37o/s/6/Qp010H8GUzaRoEQBNM
F5i9awzEQLsIOa6ElJZysS/n8jqLmSUJgphphvQbuxrW+XZFYcvN20+f6k5uSaMr
KRLbnPc70kxhnxiUjjofKjOZJyGdYzcfFFRN8+IlSDRK1myPXQK9M3JPncy5dfaR
5TCzge4mzDXBlHKIJVpR2AQh9g46xkKk8p6mu8olSwVz1bgFAlZmC3qqMIClcGbl
WLHPTzFi2/G7jVtES1itzD6f6LND4f1mFS08VxJU01dAmYNzOTXnVyT2kDqXk2Tr
M8Oji9f6Mxn+GkbDVwMnihCw1aT2D/oJ1azvxrieoa9Il7XOvmKDVuvoMMR/+ZOZ
4DAROFSe87zIgl0TUY72oprWoNXBRd9bdi9og202rmIUVt3ZlcUXEo+8wHl+Ufsf
kx+kSXv3cbcbF/VU5jCyJTzPFHeKuSCUyhrgY463Q/2rnBudVEkBeWeN2zTj5ZpE
8h0bFf3tG55f4ca7BcsBfF0h7VpLOAkIOSPMvpwb3kCYdw3+mr/GF+6dNmyc80K3
+IQudFpQZWsq/L2yCUfCNQsl4oYA0Ldn7ZBPYmSb0JJNm6cwj0MW32iPo8T8S1/P
pfh5AEIcPh+TKbRfDjqt2o/JR4zy9nUe3qaPb/eSjXauYlYRy6GuJYOee2Q85/Vj
8aSxKiMoMo+TRfrR3eoiCvrAUn0XreDQMRrJm3G44iycFGy1kQ+ul7K/X2UKT5I+
aBXXWBAm+D81SE8+b5AplDLpjz+WOF/Wq4yTOJHMl5pb1WRCuj/8YKXZwV8YSsEV
oe9ca11FPCl4akPmQ7W7KwsA0ccIwc/aQpAPK9b4Gl3fRA/t8q2+Q5PZueYCgn6T
Vj1mQDbFJKHji/HlndJhLTswJNOvqXF3FwooMfzBLy1nwmhR/7nr1g0C42Lq7I7H
ZjmMm5jsw4nnTcpRinWaUwtdWR5GrFh5WqFMTtam2Dx/+zxzF00qVPrd56iarTEk
tD2uW2jbtBqDr8zbslDH3UhjD1TewJO486pxYlstM8H8vFrL8sd5S1HLW/ES70Zy
u6naQ+eyEE6enKm3uAbLujpt3/3hHTwPp/ccYkSLTTYcvrAYaC0S/ZdMemXjxvgq
0TFFaZ5glLtF7oGPdiD3fmKR1Ke3yqAh3NL8lrBMLQwaVqld4jbQRBi4QzWfKxL5
g4OzNyR1KnPo6kPUkTnljFihft3+VCNSA7eQB3OlgDk4MEOxFHjeLjxo09ClCWUS
LYvYDIcwGp2nppeWf58sny+MuqhvBAH58KOvdCYfrK6vS6YIguxb+tG5wigU+FBw
bUQT5QL1MHK3wXMV5zxhlw/NhVorOPqKhiQ8iRyU83AE4EKcZ2q9yFfR6fKrqxs1
+UjpFhSOPGg37lu8NkvK8kvq5kR/mm5e6osyMnmMdEKJqa0HsImtKLFbNY28TRXS
PgSsfLFe10VO616VFacQAQUiIuuOHmEFkD3LXCaa+dK7f/Urecbl/UFNFBF3Hzrk
Jz/w0sfoeJgGI1zL6yEuz5xs1CNlst7j9EUDOQyD3ju0coUrm/doR3rhSFzfCUY2
rgxzMmadho4ih7weq+TDJJfFmAdJHoKmti9ppGealyot4VsYLzaJyFEif5tyqK9U
HMCR4sbbBt7XaK1YvyFUeLnKKiJEdXOSJltXZh98i9Z9+isrg7OiFy0x8x+1cSij
AEMH77sFR4fyRMdhskLpSCrGGvOTLxTBEDE425VxOASHCtmTeTu+XbK/o1hccO+M
yiT+osU0hmCiv+AOn1BqJ0Fw8AyEGkvYiERiNNuxmktYOAgyYYNeDoouV1SuewLt
XHfiuu1nqPunB2WWu4BchdlKV86hPr+n/eIQ201NcSUG8szdlyHClVZPU+Kjqo6y
cw46D1vQYgRT8VR4nde1QlIXUhn/yh9/JFcnv7fp0dpZM5UTpA15/KBu/6fH0sBj
XYLx6Fq80FnuxWFMSNGWEyzJ3tALH0ONafY3sBAXKvqS8HAINCy3E/ENNta5lX6L
n19eJZGw4h0r5+3k3dVVVCo2xrQzb1ekCdZumEZ8y3sQeMnczxruSBtYbiNsJNiH
zfLqUfrPb/VEs/bkoeloNnwtP8Zqr5UpHKYoFuJ/RCpzmssBj7mrxPDNFtctZpdw
XoXj1ctxjCMl4ZuBgiLuzCwMVIi+hD20WDsQ1hJum2M6TQ5B6QHIXPUWCWROaEnq
6Db5qilDmzxPS+6RLI8TJ3ESoHjAdm1qOkUehNW6PrqOPQ7qH57pG1Hdlu0wVSwa
ozApEyFxmph/F9r12cN6UyfQZJWV4+cdtqMnxH5j6HKg90RvS7WBTliyRyPB0MSU
0V/IUkyfxez3E2rGRICbwe/vak6Usg0AvcD43fPcVY23QbLM6tRBRf18NyoEHcWk
08p5jv4XhkR526Br3w8AJND7QqpljXEHq3xEpMtMAXj0usMG02G5cWyE5vtslu0x
YhsV5vyIuj3GBzh6fx0eRdFF/jrf5S52/6c2TfywbhF6hvesKVxU6eETSiK/+XFK
hWpKnaBl+ZRthRGWdco5+rWiMo39XbC0Tm/yU7aMk0bdsEJ9wP9Omh+h1NjsN9vQ
9letRI7+RSPuS0FpF38lifHfe2A4I0SRdSG2O8+juLt+oFAz1+x2cdX2OLIwiImn
lM6g4zkIdQ5wh2BhYV+RKqCRgiYdG1XaOVrirYq5LRqKqoyjfUlHrmyQQ27c1vie
2bCoZKM2slsV+HuEo3eUAjr1/Z0feI71nMgX4PPwQ/Db0zY6tYJOGsVXesJZLx/+
LpgdwsuzsgABmC542X05QpoGsFesSx1c+T+ou5YyWqAoRFQO4mHn9jyRci19i1Nf
Dw7vr6YWzpOAAfZ/dD9UnQjkaQP59L9LCfaZmxR7XXecVJ7RjzS5zRoW25I/riGe
StrdO3Z87jNJwMTx2nx3GGyP/FEy5vGAXGHpFEAP2IXuQfpsiPbqcrRF7LqmliSZ
q59Y5GbyJDfQyYM6H1Mv+0Azjf3v/ET+OB75ILGEoiAYwwlS2S9ExEPKQ4DMWEDV
fiJJx2uSOaePtihgjaXiQ92xWYpVNkJY0rOA7HzW+tOnFHfdemAPBiRJzGDGyxMd
xrQmoyB6ai/YyIX5iuysEtHiHg4fUviXup2lxca7VnzFFSxGwSGMkkhfCz/lv8+D
vDn4tBu6uw6NVdkXUwtAa/J5ADN+lUKyxC9ykpRnwV+n8YUV6zHgvqCAsrVrRO9y
ytGG5JoIlyMhNiK/UHrGHXNzToxGB9ONdT24ZhLdtf6VvCPF15nvjdbyKJG8lwra
ZeoTS21RRGwtHC6bg8xWXuaZ76IjhROfH0B3mcBBToGJ4xORnzVKIHkfIQmt6IpF
tkQLcLsiQXPlhVf5m5HsGnZyCxpRp3TGGSd7ofZ1IXVXWGvHKftfpIP0UuUxljGr
m0PyRSxpASDGRzBFUfCJwyrtAMY6dlN9u+HZHx1ecdo8o3mpWK6VCBGZ5I+XVoNU
4fJwX5OY6VCQztpAQsCAYV4fn+RUAy2PEU55YN7c8TOCxu0WsVcHFqrLinWxX2pc
RS1/ejtcBcm3FseTP4F4qT+rgKRjX/trNNvnLCiKJy4RnxKdOSRcoZkEFff4V6Rk
/tRDvJkPmeODrDMBObKyrnXvcQRau+nPjikyxP2sCuqi104HU1f4ztmDnMJjohhW
ZX6sEPm77fGh4SStNJlLlHCp8Jysn1JYPeS1J69cET/vKDLSUMkTbzaqZ0o3PWQR
uTAl1mYo8wBisk9E7vrtC+/PjKg5UFr2GYYk2YaxtKG7MIo/fMDmJw+QZSDnb+uS
a9wMEGUbrIyIjMkKsMtEKxmcT7Q1pYSRJDnb1MjcDCRHTshR9u29kN1sSDFnR8mp
gGvECUg/7Nv4/X27IkNcDL59wCYmNvdTUMLiI4YkENZ4vRo4uEnnRg9pL7oUvzlh
pE4OxE8xWimzyUgJlUGcAA04bZbnPdvHHwpVdFCDhkNvI/bmuKfWS0xpEHTs+ZZf
ZlXEznH5TriKPMFW49TzudIqvJwN1RcrFzTqk847XitxDv4PSafvKRLcPDtPlZhN
K5k62MHcU9uu9ea1JJ90LDQh1l0k59MgekAerWyWJr48WXWMGcxsBA0fyMiNZa5W
TjK7m0gmNC4SzGw7MEp1P7fKusubm5ffM1GdS9Z3JcSNMR67+LBGrAsXfDCMYt++
ZwJRSwnkA1ougtOGpsNYpV8xDxA536oxTJOpA2guLS/VrJwwRUHbv1Nu/1LIc75A
UfCNmvQw+P56rxWh8pzyiH4o60bgud/hfqSZa9E5Jqucrxl67w0WhDltK+vCUDf2
NbdSFP44QGaKkysobg0gH2P1P0pKvnVPly9R4vi7WLu9wBdJKh0sXkHDPMHP9t04
YEjclKb7aZWZw2srZMr3dOvFq3uHncikpZPBEg3tp0GJelQo/7fM7qHzPt3DRrgt
4BGYt3VsPf6D18xLP0H1jPbHWr7WfXmNcBdusvAPbf66h1XUh57DlcsDnndz1UP7
60AqYrisdVvOdXasgCSK4s+5eb+B2QvvETakytZgMjzPLC7EJdSY24f0NlcvsqE0
OQW7VRS2EjazB2N+9k23iLhocCutj9IrAkPR4bZGIlBroekjxvn5f7f8jkzkfSrx
4X1kyo7yPT9hrrr5GCjgMdNse54hXbEa7O1bpFpT7ZSBrUmFAKH93eTj19W/YY1c
m0BCpUQ/KOJ3Wumz0WnjLsdD10Z1b+CLsdYeNHeB2/wIwp0+P+MV341jfc8dNEZs
1Ucnh2JWHNWcJOlybbhaJJeRD1lmV86eXQtBdGB5IpNZynASY9EtfrhiYK1c18FO
95JLiifxEo/EVGihPUpD2qsGFgR4LHDZv6WOIBWOGiDKvzw12Fp3X9XuR2T9j2Gj
SLKaZmCmv0nEOk2tV3Y+Pe92sfjApQEGCVpEXvNIKD2mfLDaiZU6iLqIsS+gWWKt
OHZa7Sprn+6doM6CfrmP8Irapr7v+5gtpwBeLC6rJMKiebtFOyhvayZ5hMegELKE
YllJ4qQ+ICQxqqEtxuTaOeNy5K6DHevug6QSrPJAuttPztjfaeCBMGglF1hrY4uK
jTWbLsdxZ9tJ0wWCH1yzjoEhjaAH+GvMloMjDgxNemSyU8WegrQITBINoxlf1t93
kBBkUs3TzsDBihDVtH4S6MG5c96pmJIVxFo/ChlHwYCijW1rFyRy/Q90oB+17PHg
uqngNqMpxAsNdcOl2pJKjJcabuks+SLvKvO7SMuyF1pqSOKnJBSVi+StocHsE7PF
7JKn6kg3Ps5lfMZFYyh8MqWEpiBnMyzwWSe/9t04A32WU4j+VTaMFcAUPi57wcNq
f31gkoXOKtnXek0QDzKtTjcKT7ue0KabEYRN2R122DRP/9O6amsmXAM20lcFXnss
3XYP49+QPxm0t5XVZqMdGpboDHuo57zCOA4HX+KblH/Ot6sEMjFIIDR/EJ0N8tfA
hCi42UW4BjJdQwGITIXQCH8hPlV+UGHYl95a4DiVkF7yhty8ljuuJvhk347qPsxY
ofGcxeGnS4f8jlRyuM8WV6T6iQu5sYMwm/XJ0Oa939n7N3kg5tVAsQA0QDdLnCo5
6ys6tucxG5etpdzxq6W8CVgWVSXaG5AOP34jIc7MR7XK3SDONB9Ea7wVx/l72oBf
z/bsbkg4FZkRqV3kQze0xofidJQ5hf4TkaTwFr5qy0sI/S3V9rBgrjT+tl+OsrB5
/ST/U7d9WQwcx1k1QXX2upqKSoZ/ZcX2lm48r+u0y8cXAfByjl49i/LUjkb3dRk7
fT40R0f8Ipg4HJzd5ZuoRDpgL1ZIx7+HEYr2M4BTeS/8FVusUd+w/l2lNs2nps7N
sXIrbVRk3plej6fzPt9t5/RynlCsGWo9VwKI7kz5nFAdz8Coc+MTajtYxoZAjah0
4W6jzAof3N8VWyh/d83TaPMMdTOULs8MjS0sIgFezSg4aqD+QOiR3XeLAJsYubu0
bSgImHJxFP4cF5E5pffm9DKEK4pTM+eSv+WU1eGbXSXjM3mZeTNz6qVNg2xAJJPY
mV8AvRCuBS/4DWiO7f0Jyr808Z+3wd114FF5qfLfmJ0jPUAx3FlRxI4peSrzbOWr
NyX0qWf/9Si/yWZz32b/YRGC27l4njMhAGtr27Azcuo9WcHZvnPYozlKdO8Os3LR
ojMaz8gPepTIDXQc81QndfkoWAPqGa6ROT/wtiiCKDBSQ3tPiI6DtU8qFAKKS/wl
9OWqM0Tog6DdLOd5SZ3xGD3iBjlXOrlraHhmpJl3Q1DNd4B6hsUA2mjMzZ2cgtn6
rRNEtKBxqX9YcYfbX093psmnYXgqV5Dmls523Jyln5jgUsaTmGn996I+u0FBTxk7
228bUKP7QNiJI2uheg9l9UUmdhYOCog5l7lnZ7LZknvV2DxY70eTEtl8bBRlgiZu
UyEfj2XCLj+W89dj/YPbDMewoR3k+wtaVeSeKhVPJLHBMRS4z5WGTryKUPs3DyNH
rWZeGTP6Fh5RQhPyBuUDJ2wD0iSKODrn3Ogn+f3bJ8flnVzkQhWIVpvnZDfZaKUU
odWymgiVz8s9Wc4g6+OSvHpETghTsCGPFkQAijmimgS/8Q2Nm4UmgV62nyo/qxgt
yLrcsAa9Ow6JxSsnYZYEWLBxSTTF+Bqf4ATdUPjuVY8pwZiG4AENoPVrtQJBygng
EwN2IxbOtURpxhQdXEyiteMj/N++Bd+bvxCwt5JJF0kFWSf0IRKuM5NaJyhu1BWI
sXdibOGgOVXwLRkT1rqDGtrkphbpqTkluPTEoUzTr5CCX3afC7JCGguUJo6p4Xy0
NQDd2/50AYyeJdpe7TFEcm4S1CFh2vplsECdtput45PNfbp6kmTRelZ4ozOEkwhX
6IvLMWlPki4lD/zkfzKThm9DRPpTcDV2K+OGBEztdrMHsbwsT2wALW7H4y25ex/Y
wPttoIxAdU6zjB9TQSjo/nJQlMIyg61H9f/jRHvMiZ7c4tPMyr+xcjFmq0gJKyId
rj0vWDCtzfmAwyaoVSrsKAvMqEAkTaZkXHEyYmMd7NfsjgxzL4S9yOSC+hoThhP1
obet3QHNGCqdwdpN8OKkplSyKjQ5EXGwIWzkZ4C5YeLkr4L0anuybDa6agluou7+
Oxe9vqbGykKw4V9ULIrbnEAjSUIQIlCgAszgPquhcLb6JmaIv0fKFAo1Nb2myfbD
qcM+OS/zSKMolAhi1mI7H+TxxNO8QVJ5XAr7eXmmv/V0+TG2uET+QISKj+qFtk/F
+3K4ALNTXAlRNju0Wdz30wj8HQ5eO8SHxhTkTEVwCvj4Rsam2awyyynGhJKSQAd7
ZKAxsBxwDwAwNEP5b5mLQvsfTPxI3qNGUxL5uNj6Ioe9p62nWmz/HxA54WkJ9V/x
Qu0PgRWKwwswfHp+Lrk8M6W16dXpp/s7skg6p9jC0FQj7GL0sqqk/58ZVLYxlroG
+sGNC2sVySUjuSaVpnmw3WUhBHgah8WlyA55tEtNHQc9Df+eSowXwVyLEgB//KCc
IFf5EBmeN4NRJJ+cz/hhEfUoFLQyOZxqp5CcgltqZjVm+tMyyQDXEVfwI6Bf0H85
H2DiCSuUelntRrECesGaoV6j7TEjVYn1MO7BcSjzA4sy+n5pZn9pnDVIytb3OPk7
Vp5wVmNHG8wW1zLE+VG97idWPzR1mXh/+XpPgYWA3kPLGMV+aCDUhGKJyBLnOR/E
FOOWM9TGjCMbIxoQb4dzUVrGRk8N3I+gQNDNu7o8wdaYZIDTDb8sX7QpTGlPTHzN
V1tujTPI8/sA+fPo5Jmt5DgHOsjVMgMPqVzFdBgHfrVQ6YNae0RNijlRYtmjaNmr
4tW2mws/Ceg0cxkfWfWgD86IrYWOj3YQXDk/dZz7td5dqHcng1G46mHJ9KWfsib1
MhU3HcT35AFLLNYIPmr0xS+F2JPqgPUdYQV96HZlv2N6uxDCX48DnKUX9qw3Pj/N
8HzSxdV0wqjcPk39eNMg6N847OCSzClrVemuL6rTZ43UfMW2bic7pkdStT18NBkX
ff78cL2jM9LOBH9Gs+6V6HfbXXwLNwSTR69wWjqX4c3WufQXcXoLNZVVyJ4DiNfK
254XMifC8zLHs1skK1ZwVDUCrVrjoqMElMytEIWLs1H32e5ElGHy1WDnmgidddHT
Lm3PwbApQnXbCxhJfTrqtgMslqe87imZEyOAL80LcYgFTnn0pYaF5tnTeAyXeJ3T
eDSfrsobrWTQ2w/o/9BdtpJCgEmwfGUJaR4wNVeJOL8IbkCVTVGbd/LDOcguGHAU
0oUo5vQBESco11FEu1uSnBUEfRpf+x25U8cLqaRhorrofChCIz750TVzGP8eyO0Z
Lheb0bAQ/hj6t61ra3TzfwW1e2pS8elzdOxRJefm1DV6dsmX5j+IpB2T5ND6Y6fm
37z1d4DoEcaB7o28MM07J3NEjy8bl5KxkeMXQUMq556o6oUJW++jPGhh0YCj1N2k
vu+Wqf2r/Cy3nKmgHB8cAoH613b9WiVAFKe7XS2qOdDFsFsfYksUoTpjR6Bc0zVm
E5OS7NQrWoEH3muB1viXGUNQ342X8BNbU/xhHhyjwAH4PgrMgNrClvyb0QXUhtMj
9YLxZf/gUW9S69nd6AOkUTGjklZ2O8/8421+59Ju5Nit2ayc7992IqFU9juP8+sl
HF9pQ35sFSgaroxr1M1OREnkJrxYuYKhiD4SmyRODsvvp1FvwsYV7YHG6tvctrqt
4DCNsOdKuU6OOoZF3sNAzQ+JF0C0F9Iwo2HeHL6WO2VLSxW+D/QN+FpcCQlYWObm
tT8AK1DSgaAuvFxgOGKbsY45sbkmb+km2ZgVhncTAQ3pnZLSoujbdYsw6CYat/EH
DTeKmsivD/ScVk2RaCvHlLDRO1FZtrGowQY8oFdrFmlq0Yf2xS3h33/RRhFHSs+W
2IMdbS3y9GGFtDRHGD1NUWT5eUpyMHQRNO+mBdrjee8RHVyLm8kDEJ7uybgB5TB2
H3S7aMaqEJS5E8jF38GiBzhiBhK6Ej7p99fcWNqwESYZCvH3TfyYAwatdcFpRkNj
kFngwmu+TuATtk6fE4GuQr96C+vNpFUtfQNHfQplSdqBR9x+CyEfv49nB5v3VuIo
VgiDLFtRDHXPHijDvTd6Z81CErK/MWOsd2aPVTQPD9XRSZJzwEw9EL+erwAtyOu+
8DSWXtMOOytbIBSE3f2TsGVnCzLcyiHBSn0mfmsaWFapS/aRAyEbpolSjYKUl60x
7SDuegiJ+YTKI04B/yXGbQYBDEqBoSCIMwLvA5rsFGM6zIBpFvCpERmpBejPusFv
zGdrwPtS3iuInX4zQs9yE3XWMmL1t6H/MRH/i11AV5LH7MNwjJf6gbKwbpBj+rxK
L0G87CgAQGzZm+YPb4v2DcNwDVdQ1jvKW0mKA0YkgsK7mGIQ2Y5pQK2LblC4q9kX
7UaCZacbU4q0QvuHxaEiSL/TXEVk87lUc8qfCgQwa8/Q2Vq1u8uwa8o6XxCzmf0C
bDcpE+xeIh0ZDWdBOBX4liGQtQ27crWjCAJ+fduUzsRIoCCrK4EiPirw/wD0v3Pg
IctagJSgoRzfKAPI/fzuUwbKBM1hZMFFRKJ3Araw2KRbFL79wfUbcqoOqLFSss91
Y88fSNuHWvqdFVXZUXczY+7Oa6o/HNzMp/9LGt84dSTQtIolZOwfq6hjTOGO7AP5
+I94yzrTspOZ9k6z6KzYBqyJWnGYkxVqB9iWOTTXS0rP5IOi5BIFJkadrA5uMJrp
ZJiIwbYeDoQI9AnCtLfVUeXYnD2u8XH1pb6SwHNnJ8LwclILXYM7a0TTf6UmD1PO
acTxlMfwiEaF3S97nvQDFLeaghTwwSuaWVu8Ht2D3Xg0oxNybthAuKjECJohYgb4
XqgIWzmmLdjvqAshTswtpTfGGS4tWDcwpz1qK+i9WfZGeiZWSwrqPePvdojanNfp
1EWkH3VPRj5VuyhNd0IwK2AKbmvxAxqCc38FiTj+y5DHUfqORKQhEAlNXIdoIGQr
4O9f/aEUV4LeRu+i3mC9EwVuG71WnGuYxVjMTzNGZQaJhu4XqGKFIrEzh3iI3+2n
t30PQEwfLgOFHk8vXCJSyJcUfUeLBaIvnINtJy2+rBj/3jn/vau0QYll6TCQ1ZwU
k8HwjkqiXetiCDHIhZ71AV5xarVZAx30aftnaZwZz98JkPWxTjWZ416Csa65CYcR
pZtAQMZLECz5o2CdLXOtVMJrNh5JpXO+c0Kfxp0Cd8kEU6IpwD5T4B8NCP1bo8Mj
34ckrx1WgN/Z2XnQ4b+fZkln9VClE0QXe2qj2WTJJNN2gTX2KV737PqK06Hhfndj
GPHGFe4fIlsQICIFUHZUOBZIsanJUT6XOdybRaqBqjyQFEEtqb8YRqbUy5e/mTBf
gyWqkUnH4HVcepxyL/VHXoL22yAjGpFS1SzE1IBmiADWensQbnwyslB4Df46SBLk
VS2jSwgpDnBBFhLOAfeG0YdNHWKGid05z6usQG33t23RGXz0GVGAODLpmPSIig0R
MrRIOzJxLHjO/Hvj9C9lZVzH+VTFIKx6QrlUG7XGWbyX1F/g+POGh1EcTEwq/ArC
10yNVncNCH9bexmhUlGGzSSsYOaJGSO/5x0N/Y6zHqtrnituJ17tcYEEyvZ+wqFg
4virw+tjGhO0eNZ4bDJ33B0zTywQPNq4doQsnkTRK/GfOF4XqDP/WstlLSKLDRe1
2afaynJNWgd/0hACE+JvAJQ53Zu2NyZgAWt3mSXwPh4ZYUHIt00seC3Bga/OahDj
6ah0QdlhIhUMIMmMdtiAYZN6tXuFXGp5mJsM84aJSzt/CHH/lektNiUKWr0ygjbl
LcyJ9f+wEEUyrQOp//2oolqFhXzKOiiVbASpHfGVDVs9BtEz3HcoVFVWrOqjyUBv
whbEc25WFWUAMiwOgXHRpAiUE522ql1gkW7ehIJ1ZSYD+NGtL2NqxDYVyqsmlrq7
N7gf3bt78sB0mgsdr31pP1Q0PkqRKO0wr9XtI3QbG8I2gchErj/YLfj5zv0uWqav
mRJjTZizfEE2ltKTafo0QI2A4j+Ej/DYN1umtNT+KmOs4ZeBJl5lecIS6kzQ6Zyr
0QYqi4pnp4RDZYh6EnLoiCC9OvlqHO3pKSwVj+lMTLT65iMmOeaweTZqTDBR1fm6
ggtJqMxkZD9wUOhUJZbFasa/7rLlJJs9GnPDt08BkRj1eUneUtgxuKNP18466KqM
6OyoGz6HOZgstQwuCN7E8ncHhbnZMqUiUxbRi4hEEaZj/Qem1exgAVWCgqxnGDzg
El9MhKYAIL1YoXzozGW+QPhVj5YKc3ULXibWk+k2UEf0FtgjEYmnuepsdXuKtCam
NPkcIA2VVQFQnAPONu6d/A/ksDVAkDc+5lmKKQ0ibGNEQow7m3/79upACEqoXdv3
hBB7ksLGQ2sifySSvapZfHN0oD19/YmvCQ8nJbLw25a5ucqajETZjKvLCZFwX1v1
624qI2oRao+w0JglpbCUqBHf6/2c3P/HnFBe4j1UL6JuwF8vvNS95V5IrneSLygb
R6N7B+trapILd/W+bkW8uSpZhIIDjNSfzPXKP6Zdbf+g+vvDbYXvTAhsf6jwSMJT
pkL8hVfOGAP4kARnI0drl4yHGxmP6U9LJzTXm8wGN9tMU4g2pYlXKEbu2aW48kgt
rfH5mNX50CLjL4QFACkH8LEuqV/qdqgb6qmOGByM6LCk2zC05IGOl4e3DqyTKhM3
EtA63m7dSjKv4B8YsM+UvEqTD2Hm9MaXvI50r1iW73rB9it1BPMnmyNo9iivzG73
x6j3XD2dAgyguyG0RuAeXUX1EnMYqkcFVhkUeKL4YvqqkefwnHdnGON1P7hqdokn
PsEZqvk8tNwbQ85KmBL/UqjthdgzqZgxWQnjXA694qVOQpxope6+BepGcjdEkXAf
ACRdhVtsQuSX64z3uR6ITx5JpG3Nxs/vAwimZycN/hK+JUobT6VYaedQQyzllTZm
mMzq3MuRh6/eGIFyt1bvicfpzz++1EEawuFMHQQMtHHjStY8IW0UR0GT7qmyHi4O
f/j/jeeG0tm4iMtumF3oY5knjLFuzLMFNsICN1ygZJC3pl5CY+KQ8hiHAYlMSKde
7wo0ZFEws9XY8dQKjgv0cNhYS7vleafG/qIqm7R/qgEHrZVoyE3p6o+q17zHYXPI
HmR+JMaFS6CVHFZOSuRZY/GsjQNkt52+NGMw+r/djGxraYnWsJiqRW9JAT1xqmSy
l/+p3fi9DJpGsKQoGkQOO1eAzjSo70BKHpguLvvwOE4wbdplPABcVwcWvRnCoLBF
EcaxNAsGinE/JnENUr4fYg2nDd5N64aAkHG4PK/yUWLUTxjRgU5HxKWgw3s4eVxb
ejSEb6LTh9Ilj0OwjTXOY/NK3cMVeuaACQgJ1ENk2srkQ8RzteLJ4g4E64AEnhOH
/f1OO28AHnZCb12cYlVBBBz0jgGS0fzIsgooxJGdHSDLFKNrcS6RGpybgLo3cHWO
81nLsaCbHp3/APfDSVQzClUxD3omJvE2Egm/b0z8WN9vdcuRKWdsdOQlnh2LGNMi
o6bvqkT0b3sEyUftYCxrzT2a55e4iQSozCylQsLDcWWRAFGEOqYmbu54E1x6dfQ0
YcyxmaTtxNstEP4G4vxZfPKQoUW3rt5K1kA7/HzH7+caHEkcVuVWTHDKdIV2Wirk
z5NuIVkKBwqyEHyjnwkyNMYJstI/cxFyqnz8tGYJr1x4EXyuFpX+qGRNMmtdiXYH
4rnk2WVX793az97+fa+2COqhohI671IGnrOb85jS6u1y2j0QMMcHZd/77MjAnhNC
kzei28y/6rKxT+F0emT1m3rRApSLKiwvj1C8m7313g7rsIEdbkigstmdpt1b2MpR
5QXrUxZc9gdLnNtX+HuxxS9pOmRzawDWPnwD2J6LPi7TJ5VHZ1TpAxx4yF6VywU2
RftunmjJqjAzJ/6ziMD3i3N82ZhSSNmvN4VMxxqkLHwBxHooaJYVEPBOTgE3MysQ
o1CKUOjhZgrWAPUQ8tMDFmg2c9sMXgxhMIuk+5Ew/4dIwo82k5BPts0srF7v6SdE
dxniWJt/YErhk6z5Qqn8LeEMuOhTTHRlENk+L03CYTes8SmE4NvmXsP8YmyhDll2
j59JhBi9pzAVX7Q+7lyO/CUQxiW2I+ye1Df1hswxB+UQa+AGsjiFMQEz0ral8iLj
XlfbXFiUYxH7GObIr4r9st4vY97W2XxGpok7r1QsBLacfNNbChlUCtfjSpfxhTR0
l8GwCNMwPqd509BPkCmfnzqzSuGj8Tkf45kCyYUNNV7GIn3CWXpUVEpDeEvMgDmb
23eru9BuJWtuczbzRDeXPotN/GQ1Mgd3aPYbd7UBhvMEvMs9TNJyLpp1y40PwV07
aASphId5qKBAMkbEkXVy6TwrqfzsWbN/DNUUFIO46IZjq4G6HvHUnUqCg+in9LSm
TDEwRGR2NRbxSyhdB7LecM7lFYynqy1wksDJ87X27KVxF6lNUYycoRhl2qwd577C
Z0GtSgoO6xHpL8TWESHCPDH4LyfYALK0JC1RKNsRqRpk9+kP7wDEdtI3AEV8DgDU
50ipHJYq9hrHXOCBV7n4S1wzM7QTzQyCK00GLzJgnZYHDBLK4YTB2j6QAmDy8qxx
jq4sZe3IWeTvNot8ioe5HlJJTZl6ESHdxhN76s0aslHMWCJ0IeQDNaAWEn/VsN2e
Iui9WiWmprv17CFgz63f9blscc4HIyWGLsFLyvQf37mucBKdpoAIrGEOuRnNCruu
8lI0vmNjJRiBtltciQgzI/Me36EyETWnOBCuzKdmOCCgOV9V0s+xNBFsbcQTl1Cs
bGbv3M3d/zcXEJmNT4GU9oLzM6skG1XKc5fuCX2KEW60X++HN9ul0B/n3W5x+iZt
KoZoSnB1P7Aw3uK5KilyVnuhMuM3n2vWffSuzn5pX+aDFm/UzRAm541cCLQQTn7T
IUM3eiSUiw3yH3RPHf+y7Iu1ks5hYMAEK7Jc7uEeRtOY4N/+zY47g+6cz5di6Mgp
0EuwlG3E+RM3HXVVNz0FkXAPaf6aB0IMhslc6uKpmSLlyUjard2bZUcUQLfbEkNO
bYaLj4IAj7FYRd9sdc+UpVHXsRizKdExbFW54/5zBSBQYPCXhQOE4ev1EuOQsQIS
XNF0bAATKBWaX2ucxTNK0en/CUT5q3IQs7E0LDiSNo0pHgbqzGpDt3euet6ENChx
Islt/GZGrllchmzY3dRxdq2eI99Gc9cBW1skNJlKQiclcmXXHqSSNAgvIXAsVOA5
VT2590mi0pyjf1SRXhW/Cj+lwhmC6rntOXU5o3Y4dZJuZqzPNtyzYnnfUHkxKEMG
LXuo9MrSerubn+FSOYV5cW+KF/pWmIWq8bMkrLIF0t2E7fkzIG1Bnr5ZHz81X1PM
aob+WRiNZ7DSEGuKV6eQWK3ER0HUN8FBT0g0csOlWKatcq8ZW71mrPTfzWPIs26S
IkjnD/dP7vWQnpgGOqqLpVhqF9wB5zltXK9wxTp5qbZ7G1lTxNzP0LzMWTAD9J2q
U1OI/ajOgEriC9OxohqB4gHT09cqbiRGMHiZ5ank+5sN2m0OR2xDoR6lNP1PS6xc
/ipTSaCr/Bs20DTDQfNupjHBo5AVnLXZRbR7a1STxCdgQWGvhls3GHa6w0H3UajA
Ly79dBsp0yYSdhuGAPnlOpDabHVy8+PGJKcdvwWs53bf5zUAsRoWL7yVNcMIiWrt
9VyOBqEUKdjb4Q+WvJy2DI8pjGNAGEjTRoKBsrUfJybx4z2GpPBnz/ysd2w44cvR
js0ACCDjh9wlboHjEKsn29zwqlqF/zq2i6UuSvN8NvQDNgovjhelm6cStlpgM345
jQfqarQGJZLfFRjVnO9aQtHJFx9aw0aZzpik4hYr8Yn+p+uETFA+3230LXhWWFl+
nQU59Ic/Z1M99JU8qcaYiCnpF7mLjuliFnWa5n03XcFw2nz3r/RIfu/b/UZq25HH
23dxvLAt/xabnt/kYE1jauQl63EOTA6KivcqaqUTvEF++SG7T3Y4eUcCnPEr+lBx
pdQqtUgImWB2iUjn4Sh7E673yLD0t4gqk7cX1rbZZcdiAF4gJNJgV/0H1WZECpxv
w1LdnTB6w52HUNfFqOOodcSIUfqqXmFwGn0xx3iIHIhri+F0F6owww6F8T3Sr2Wr
tt76qm9CNjbMqV4Pz4/stRxIGhZjT2aM8N0ZfPXhXUAuZza4gknmRGyMwnSPIY+B
Bk2SZyCmq1cO/Qm/aAkGCjfASIDYh9n3j29S+XZAxqmcEVJNxAALZOW9DGAPg7DX
FZaEnU3tS4AbXs2dF3NX9bvc6JNSPvclKCn/TCrrNQVzxlHg7WMTGCK7viOHqMpf
kD6Sw4mkl0r9pE2DvCPOHclmpjJk6u47FipIUt6t0R2GnJcbMBxQ/AwJJoWQUy8j
mqs1lMSL/zAHt/M5WLDdJPJGRUOeF2lMS4nRQ+CavOngv95G7Ra3KqaJ/VHkRx1U
cT+pRNx1gWWiMo8WfXQ2Q7L2w8OG9AEiBTt/jWNoeBTGZea9Y42uyCW5M1HkPoWx
EkZnhN05oQ7RO82Q7HiVAhjhyY4Jnzb3l4GhT9DEkNHLNIrgCshkXU12WLOLe88z
C1H/9ACjU9d0sy0WEazod3vp/GQIFBdQfD037R4qCL3qx10x0c+HsmfLPVKvYZd6
Az2SHLV/w5hWEEY+Yu/Hx1T4Bm4ze3he/18guzjP8GVrGCZWcR6+xhjF+7Y+zuqo
D+GoKuLSmGTQHxHcp4jh23CiMT4EeIx0bqhk9KHd8+ysfUTb0XAscQy8OaxdiFM/
BiABKkf29qHPrUytXkbdyeOS8nFU5/YQMIh0pkGzNagz7iNNGRCDWA96izgmk1C2
QQXnYUh7wK0xFPwAgeVTK2dA9VjfS7vZICDRvlllUq7VkSzWzMgqh2La7vpwA9yk
XJyI1MgOYcoTG7/ODjFuHO7Wkm8LvwiY+Vps9ef8NVziAt6VnLsUFGQHZp2THPHt
yUK3+3JT0fLW95/iPbv4xEUpdou+IdxhO7gdKAxy98llBLtq2Q+4iKvAbN8jmCeb
Cx73jESiK+ZtJSUCPREqGmgrcXxj4kpwBnGqoZjbx538o75AGj8ebIpCkBVqFJV3
vRnO4fzG3bbw1Qt3ArbumRcnC9QgEktW4Wu3yNXhhC1NlVKkCkZP4ftWL0xAzolF
LY4CnGb7IyjPrRmvPv5hF0f0n9SDBLDLtx2ZwMGUNw1xecfgmxTbn9Cm4FMFpjE4
aI1U6liCuIQN60QZLiho+Hi/9kLNOHkGEU/qa4IHdaMrIdXKQeaem9QHoQAIxXb+
AS/DsIQSVcNv2pNNRk2vfrytwFOwa32/TDOsi7WeqD/Nab3OytaWhQJq/kA1vZo+
5/2BaHzUA2+BmgpTF/FBVjOKi+jbtFXyR1N8EDX3WR3kYG6beKVoVCuY4kbLohvn
cEGK9YLF+90GzbEvXAZmdPGN+1ADFcXEKbFm5dpOlLooAkR4ZC+7IBHqIJgjrogQ
/i2RfGUPQzD+ulhrLcq+E3IIFmzN0/bubzvRTXu9o6dBfWELMOxeuBhl7HCq+DXc
/Uof8iK1dZNvdpPRdDmSSZFyguD4CW7tAAIRINjGFyOUAFwC1geN7Eqdn+K03ynd
C5dMS6B1x9XHWK8zWikkyV/XPBqUldexeu4EqEELJmjSwVmFdbeq2f70/NzBRyMT
kduO04gHxHC935PsvZ84YQ/v7Elf8Q7TtuRIh1lnAz8HhujpJIj41xkzE+J3jF1W
gDlE6H+DEs/aP3fYqEsu1s2KqLmkduPcr7tFkS/4Zwtx4mTzi21sD51rnPfJGEwj
s9UTIbQPx3uLlObgeRdGGrJy4v0OErC37f/KDbF3Mofs5ubw2JtpGBD7KgbVv98v
RvNSS1WsFn0YuD8qBsoSgKoNHMctTKPo4Bgefuf73qkwXbOqTUwnK9qwdNWFQv5L
rpUeMiSWieQg8ZGfC4ZISbywe1FEImcY2pGxpUcCVM0/0IyfVRb9bJXnW1t3YYmY
iFF/lxME8K0/7GDDRtckPUqghQ+E3tkWIBk4B+5RxCjn04SmPzsofixUoXNVN/9S
GNI4aWzd5sD9HlNVxPMx0opFyoTuGQABUHRERIaitO5WlWPwPA2P4HbQAvGPoHvd
BWIw7+b4i7r/9nea5eN5wyKtUBGRIVUE+lkYWNwVH1reQuYvuGCDAbjY+Wzdmshv
lH8jEJ8Lc32ZiGZiNaL0K8S2hNTQCdACEudM0oTV7BSwfPmrEcm52vSO95pgy3ke
JG7Zzc8W2D9AiGZEKNNKtw4z3CN+Mvvz5QuSr/GDEAIL55zDkpKhBrSvAsexRGBo
aerrqxzQqnkaVhZtH22+DE57b70XcV5p3CMS7u7bcyTRsEox4YM3kAzbL++Fv9WZ
OTKcAvkjU2Coy8tKkdTH2cV8VJPobfzs2XLA1jqYPT2JSqQcOcj25MoDA25YnQrB
H64lZv2hZA+jqn/mR/5kkL7wer0WXKfEUC4SCxIk1tXRHUaMHQ/MjM9OJ7Vrg7fd
Si8fk9P/f1+sIUyryRKQJ4shf2HlkoKvhnVkCmZ+c0JL1cHndvMr2IZdXDTasrwM
D4K1awQzdHL+HJ0cRDozAoG1qjUqEY2swJuPLAI9N/xKCWoT+vGje/NoaGjCAwEh
EpAXbeMzLSF1NsTvyAEngyBTgaQwxGCtCJW2TDcYRELSqvddDwTo2BrHnMvdxgs6
Vlch+jAa5nNuHitpif0KUSFMHPl/jtWPmCgQ5iTXn4iySSxkJc8cm452nXa2E9V8
4oOjZTdSmo9Z7yokEGSuy6OpxsKzRri43wtXFCa/H6nL8iJFbiR3UjFjtCQ9uS13
TmzaC48U7qYwPPI1X5ZGRYFoGoFbV1ixzg+eS9D/M5zltDRhNWQu7Q4U/0xA7moo
Af6uJFq74BN2HQpqKvc8L+qwUuNkphcPDP0z7PXAvtOQQK3QfoD/yCYWtFKNbYLs
wP+bx3ARDQu9eIgKhtLlZfkkSCc9FiqjUnISvZKL6oREHLM3C7I04G+MVojFJWid
Vt9d3y4f8bJxvRmtZVyAlGaWqToziOvVaY4qbYBgmz0UfgfHGdjPYOUczb35hAkK
dfjw7TnbLbzczykagVg3eM0WZv2SDKBnNXKx5RsE/XTgrvZURndVpwo8z9kUpQez
ZgygtFwik06Dwev/iAZw8XEufgmYjU7BtT3zyPKwze/0mtIiYvquFzHbMuHqbw/t
tYGQe+p54sKd/3rNwY9rctDbrTLV/ZSgj6PskAgGJbx/h1HRj1YqDn90N3KICVM7
wi2V0PDEnYwhCK9VXUDAilo5ms6+m+xqRZcbH/saUWh1vuPlqe2rttK33eEytVnL
R0BesfTHxh4dwJfQo92kNygMOM29Nkb7GtloBHJpfPTf4w0fHSOhnMSPq6yRkdSz
XoiGZDUclQOaAVhdzgTApyJKzUCLK6zR3v368oTwu8iG+SKlyqKAZvbfbDB3C3u/
rTeZCwrBL9CRIHR6UBNDgZOHF9Qnthv60j286RtZOjk+tL/8/Vm54osZ1Nqna5ZR
fglxKufZUDgt+rb83i7JnY4x0s7OVo9uDB7oDXgOJfENKcYeMVWs5jMKDyOjTQQi
ohRB/dL8xoLkYx4bt3lMo/qXyZ0e3m+yBAnK6/GyCtZ1d69Yvtpk9OUBSotgkrEJ
Yx83kWVijw8Uht4h/7PhJFzwMUhMwtmGhTTYVJQrQN+doC2m4R2y93VpL9sZQk5A
1W3shAUkbwVAg7x5kH4y7OniushdSc5sAXfrxJDBbtpPbHayCKIvoT3ld2VB+5Dz
+X4NQmzb7jwOiUk7GveIdEE7YcyAML0yHOpAc4ZE5z42buF5zSPP0OiSqFTyP/2R
LFnbjZvRUS4wDjBWb/CFFzbCln7YlBaRQ5gFBCz18U0YAB673VxkqW6PwWGgwIrC
fLcRmvGiaOBgm6+QALiY+CEzwXqp+nmZ4DnI2nRWvKLmPMBSN/jURlfOJgB8Jgjt
JBS0TsX5Fr0Dm/G5WansF8x3ZON7FON7295rNdwKZvyL+3ul9v685bZ7hEmQ7irW
lpm4bdTbS7Mp0k1/6AfxWMJWYHx0DvCuL7wSBPfoiARFYkk5yExlconOV2p/8XnL
iNj2syPKsET8fJg8uBSgfo9gVNXJ978xjPUVlY1FzWV1lmzH3w5PTgej9o88T+3I
n2t6goybHNuX14Wi4Mmm8uC8pFXw2ao1X0n+SBST4CNpHJn3aWffZr9HW7hbrxjE
GaAnRUdFUQPFT/eevAFIKGcXwGzpJMxumyoJo2vN+zvDVz59bTiNJmzonISZr0rx
XNIOjlZTW1Tr7ILc4bqkq/y3kt0okRNIcLGKrirv+RjM/I2iWdfukTKKmlUfMFlW
B6BD19viUngyuzkZ9s2kw46fiAFZk9u+sLRYIpJzIkaAqpTKqnvsEapD/zfnSu8k
WN609kuw+mA7vKqhsD4tiTt1RQ7uYIS41AS6emfuWBo5ZNtCgpB2IVyqm0GSpNjG
V4QQlFVxpFQq1slIdQrcZsFU8H2Brd8Askfjgbfd0pJigKHt9foLF6SxW6EUKfT+
Lb1YRjHtlhzkvs/ghb3qL/GRD5RpnyBDd9tXOqnSFgdQWnO/lE941em0c8RB5SGO
Ixl5hwPNrV3eZGFloeMBn8qQyS3HAQuybBl91qUSUB08rT9Ybbbe3H+FqWBw+i1K
+dtXfOegu+Es66Kexj2nN1lpkiSg6sYqN+Jkwo96ojl5sAqWqalrcRTpOWyi8rkB
ai4ilZUXk3nIbI4FJNQAEVfLZ/vIsowQG775v7Ib1xr4EszOwTyA1iZTabDEnLY1
nm3sBLCC6TYwWO6qv9ESXrt0E+uSNMngxPODeSKNCoZPmG1VfeZo4dKTSq4H7ZcD
R8ZTLILMzw0HffrcUdiCJyVqiLjqcu+6A51WlSd1hZLBu2QsRl+wR7tuFGA9AtH+
r5+iLfHNRwc8W3z0jf3u8RCW2JyzgleBsFs/hZOyUP1pJ6t3dmhXd0nJUe70Slru
6JAgpB+S3nwbd49C3bR+xgWzXAGfi+I/cOv/V4yJpnABI19qWuntiTWntV7rFlV9
TcqtFHuEYU2OsTtfLumOHsZzUSqvz/63r7IOAlnPxgtVDDqFGkZ22Olt1K2qKB93
SzPTLPTrdQVirzTgJ4t8yqimhkxgxTcT4xku2krLokXM70FMkL6WTV3JqsYK8VFP
vN4l6s63kf5I18q1nSoaBewV8HLDwUuYxvNWZuIIpa8sh+QcUu009t0q8vkrqswu
FOqntxoUsrdDrdejeS19QlUCVcdQpbynm8T7h8v2m82SJRlwrPzBPw0CreS161Gv
dRjhbjO5QCjRNXWSXXerRBCrAFVKEKJ1KjHu8dpAMIIUCoB1/mg6Iyz0qvjxlU/Z
pQdHxCPBYAr0f4olCXVIlRUQbIQtPWSudYG/SepdNez/HGgGiICqnqEUVtmiB7ML
fa36gXQrit61OV78jejohZaKlw7KS3XIYZ5qWGCV0vgnzRJ8bnlnAykRngClX1MO
xuWGIcjpiLaj+w/deMpgoG+/2ovBjfdZ07XzYFK15Wk4olKz5N8jnw7hmY7q8G3a
mSiXzyuvCN1tNFz2NQ36mj4uiuxd8XppsYAz9wupMe5Er2XpQ6LrCMsL8W9KGQ5+
bNaJ9KbVZrhhKhbAtCNVCCapakz8ukl6Q852Vk0ns5mgZvVC9NelJxPvtWmwlJBs
1vzB2I5CYvAdPvA7Ymjngc7qDP1XjE2sJVb55qvo82y2t0+ATt+4+1/mOxYEp0OM
6nblgMlUPXclk+C7XX0BNbRcPr7VTcDg4qqCks4ws/UvPJmqvNmK2I9s80+ifhos
RwHwKcwXRkzlR05YqoL7/cfjc+6Ut1aprPztLFOXuz1ry1xFdJHgwrVtfy0BsbC9
Pkak7vuwO3HH6iJ1d/z6pOlEiFRByvX4bgzqLWzNG/8FALfCMS2ZbNARSSTYj3Bu
8sbcxO/poDtQGRibTfk5WEwpx4gi+249JUQTTYv5UV2LFRWetDx3zaTC8zH/TNXi
gY6hifdCOVn8yWC1jbT/QD0amIyS+74KZv3nP868d6zQanjOooBdKETd3ItxXHps
hXeEvwj4zcuFJpIwfpB6UBeuWpzXhaKr2uz6bfMgQDt3hQoGukgsbAB0E0rPewFj
3SdhpF6aVuOwsF37DceIJAKqmTlse1XsE2vPi3ox8qE1Squ8A5gAhEdMsoOetaPL
0ZyFBOtX2BnPfWY1rGuc/s0OMFdANE0uKli6d4wr1BwbKOO3GVsXQqC6/nx+xV/6
N+QZ90fDqo/bYI3U1LfK4vdMJ4rFc7WN7TAYJdefOdzaFc5ArKDnYl4adTDRlbDX
GdM5GQNghIRQNThucc69pVVJj5FI89Jt0qN/a574saBW1WRvi+Sacd3Ptq6uxpQ6
HyFpbAa/A6goIUYLhtEuUX4sNWADKy+wHJyF7RlLJ8fJWcwgFPgQD0fIPBos5r/9
yQrfYj8k7WNYKBBiL5M+VSZyedAgc8/9MjrHJAzTTevtd2d4FDTfMvBU9D6gcBlI
wzklnRUPq9DnTdhbGB3TyX6kF6P+IeG0QgaIKUEtu0FPtmErtBRL87riXUCIME9y
XFl8Cj4eJ8A5t+vYP6iH4A/S6O3EXgMGiXF+9Fss2iQPO0DObrVC5kgmukbQBPQO
acNApj16vK0kNue151mK59TdBxRFh+IxdICnBL1a6RsjJ8kWbxCSTaE72sHMxcO1
4WMrBlFF/kKx0HpbPBLsGl9i2rGftJgYcK5TdDl0Vi2oGwlBG8SFivP3Lc4+sLs/
4F7h1qLv4rZ0RrKhVd8hmM/gEJiejN8CHpsBAnDZqNvXlMMPIwsr45kw+bh+fksK
HUcWfOOIbdIQelB6oyyIIOUfHoLjlcJkY6Azmak3gvUgB0ujqzpN4sjWBdzrqO/5
fkQwHbWek2wgC9oyvWGnRkO9/iPn5ff/uAldoHzSn/h9Qero6gfSkSeIp1x38F6s
jhP3vmUnLQ45CGn4u06AcMgpg0P/26EieX16M00P28KupkLswfLjvDJi4cOLT50A
SGrCc3BXjlMi7XXihuTKoadv19f2MdhbVDBq6mfKuVb2/A6qc5mdQEQlGViH18Qz
GKF5Ic/nc+nB1H4x4wz+6VLYPWjEXRmS24oV49Km14GsRvpQkql2sI7EDmwecJsG
rNmB91V+IIa3u0MUg957pTnVZ8gVgVjxhNXpP0sKRQar3U77iiQN+q3DXpTHgmwl
bJufCZaWz17oHlF7dnLb7WTOTqsCP/4ya8uCPaHa85jCNpvwCl0tHb4iFgQa1XCa
NQvLn0Q/Zw1aTa/tEj6dzIfL3KKOVJEYZtVShZFEZlpExXLE3hLRwlwBrDFBM5qI
wmjIjG5gvAqpvOdQlGvIYhLmmMpMgsZdNsFwhBzSvuN0y8lAr2BIrryYtpDsMIle
3KNJJ7xLFAKFYzKW0C6X/1XLzo8J2HE0yNHlrk4+F6JfRCtwh7aJfCnSyBYccK6B
SBQA/72Yi3r+cwWsfAQiwX3MGOIklEYBVSjR6I5w/070eDxagg0ZZq0+lzUU8qXj
cJJ163U6sCUluxeAlGcAovBriG4ncGWHO4SNBzS4L/91IxlZoyCvcdex10zDUFip
DDnTk68y/5x3GKF01vwq48WUm19+2Ha/s18nlmlvUQaAivHjVMywUoIKEbjWZAiT
AgpHG/xolooSOdGNjzHi/50txsaKCDTGYqESwXf2HCR7tUiiIDGGqpbqY9+d3SwE
1T5VK7kIPytbU44MpDwtH4lyQ55kONJR2jMnyFy4RvMrBmBE/XkEUl1FLghGy6I2
0FuP1DotRc24Nu2mSWR8U02qAfx6yjerT6hBWm436uGLsaT7Hie5S/erEgcw4Wfy
sVIUAjCdww0MBsE5LYx5ufGh0aAWhlQJhH1UCwcxtO0QHI1pWpAWbzYK+WqyUjrN
P54Bwneq7wbKu/vPR7j7fe4fveE/iKe5usYzYPXwDKlbu0roplsEkHNk8YtypyUX
EkTVv0e/THFJhxQAz26mGqW70lForFIdPERuj5TYRFTIh72z4IbFtcXw/C+kTxG+
kvmsYq/SecoJ2WoWIYOADsLRMQjIKKWhsbnnjAN6ievPs6YPJ+JW7SfVVHwea+Lj
bIPGB8/u5Tbh/o7o2/n49rYm1pqNNxfW5tSUKGHmMS5B2aQhZ0x6p2IqHvqGlko3
FadQeNS13roilAZiecZSyee1ppDTd6LGMWlki0YSyp1ftcBAIVRdibTMcLuroa1R
lkt5ocF95V/1JWzklwhj7at67HxkrB8MYC4tEL2XE2LAm6pHVYB/CgsWEk0AP99a
0jY5zSDYPdinYRPdobSSX99GJL7MziILm+J6T+Uh3FJXOHtmJ+tG9Sp6C6BCbm7j
eEH/dY3Hfe7/AT/VI7UKheT6PAdSh64gBhpMEgl2JAsVY6BvKQ36HR5LbX8ov+gb
SOjBeQrsnx5VS09Kb/N0mysLlyLk7gZhVri4P63kfs7FDG7at7IAe4WOvegf9rcA
JeYzWFPqxbTogTS6ALPXR0om/F/Jcya2ViCSMW7Hs9+29B3uxfRyHW4M9+mvl5Kk
bHz19Yy7BfH5opNYGLMjimS/kxep75B2a9DnqyuQzZ2/oB8uFfeY67hsSwMFWx4f
XdoTTtXYpzoaOCTDzkK/86a7CO7owV5QEMqAnO8ka60LCtgzJluUg4frLpQfQMYn
8rDFRPN5Y2ApchPtH4LXKh0qFNYPe0J+WwT2OWzSeMi+dJi7pzkRBDUdKC2JHJCA
4romTBH4TP4Y8GDpiTqhx89Cfd8mJHGMBkFKwTVDcTCmyehvvMR08LuDwGQawSIQ
NZ8GmHyYZf+rOzaTjvs4SxW7jh/JyHsvm4PA4hrrFvVNBLo/Wy9P7L6lQNmkwEVs
8sNmeKNXC1bOu7q7DPenbJHpR+qpGXFHr9JXJvSXu8ZhM1o7NsspwxA7DvF7OSkA
fcRbbcVKDHdYGxpaTAA8HbGx6IMaMeUwXrMH4lu4DFkqFlJRTfyLYjwDr6yux/TG
wdiGuUI8xcBBw8BiCiGY5z+gPoToSpuLyeZTtEngPwQjDtlsBhBqKTQlNjn8Ej1F
m5RHM05yQ2ZkiKW0JIwoa700N1kBMjMu4PP4P2AeY1b9jRVcC0lJBE104jkpsq6G
k6si+gJQjgff3LUsa/lI1zlHillhQ2QW11r7rHW66hWTYIV7Rmx9JoMoDgSdYRp1
p/CRF4ach2lBqueyi4+NS193+gOEYXQqbYBPqbLOX/UNiFuutVCIPbyVmY43l98L
4bMfYxUoocPq4Mq6BIIUwlW01h2Z4Kk5PqjB/zCkwg9cCo0UVoiKU31dhOUCHD/U
0IUKKvWTKxmcUd5jEQgPl7Jnj1TxI6XbwXbtx0ckoMtrku1d437Yb6gz+25MYpSo
2IIZ6RQzv8FpVt6pmqbTIsJdXByFBPzNs4Dz4NolyTWooSBJmpzclriZU5Lw7TAt
jOpWXBZ3kOlz8EcS3nIRZzwKZgYAsKuGNTQI6V6Aot0eLPlNwj3wc/dC7h3OUbmz
9SsG/WkSnrWtueNfN49uA5ZH3wrLEdzDb+jB/DGm+xwfnJLJcAeMXqHxHLiBYZzu
av2JVumO/RE9GK8dVwU+5NxCbtegukLx3VkETuj8WKaCIU8GVHKfXjS8H+bw4hb4
WCppEf6bLZHIOx65eBP/khvUCfP859/rYjg4BtSyQ1AQDlkIxPRfJ6UNZfNkWjvI
3MFhY41HpnNwD9mAyHu0kxBkzTa0I3q9OgOqleb4UTLpHnVz9dnGfLYxpwR0c7jg
jfJ5cv00aD4mbMmJAQwQqi1LvbZ/YCMAR1EMZYsJHVyErrsCY1iHUnfR9uuRuvO8
J4kK/LCaqDlWbPV8xfpvsmILqE3GH9v9LbOYn8bk/2e3R5cmglm6syd983/XHb1M
da80xQ2V4dhJONlMPyqNwj1X/YNL5WKBc/pBsGD9LyTVc4pYmAXzdxWnMjrwXRvv
qOPbCG1jMhQPS8dMX1h3UpIHXYYIXsFy9yegVy35cnu3dYFXsC1YwkCVOklwzGom
Fiyd0dSdg/o4pv7Eqj6qJD72mKFlcMx7rkK5+cVV5yyoZbduXlyoSkYFPVAClfva
QClUDXJOhVKuyvb7rgHEBLaJ9KvR92U+SIwutW8Nde+c5WbDHXIS6nSRkerol3vB
oYY62gEa2x1O6t3CRE2n2XSB1/86KVe/krF4tKPxoRseleiSird8RqNHEFKPYWS4
xiZMqXcqUQo8jzh1juUrcXJ+FvChfdoONhU5SlVMFkuJbWwv4MSaqplnTXTBXK9l
IeuD8Z76t1FbcaEKMQplZ3xyY8pZHeIAb4vTwhxAkisIlLIUp1HC5+/zvqEP0FSk
nrOhWr0xAV+zYC8c3iEiPEkjzW0LIDydSLd1ov3Jz0hJCWqGX5ZPGLXuJVMAINQt
U4QeHlqV52HSw3N4KXEvCY1Kya8xjH8x4gelmHbbj3RwN6ESZ92HIck8SBP+sfr7
qwCDICRvOYgtTA5S+eB8+sLLy8khpiefQhO/616fhxG3f4hsx9bSDvyG1sh1E1DX
XausLQbVBnxIg4iFMSVGZGC82fPQZNNgiwH71oQVUNt8PNmlZI8ou97rhjiPmU8o
CAyBna58pZkqJlG//Eu2BUJykNBsyJ+V+Fyij2nffnNKkjOt50aDozsIV0jtv0h+
DoKwcprus9trJLQDR3WILLTf8f7/0mgR09c6orhzbPTDPpLtRDKklQHxPY8DnHcI
gPe+VCaNWtpDMJinN3uaaa4p8I+xuLIWSt4cl15BTtXjYeRMJMHmRbrS4VLyP9Yj
coBlrJjJuwTKSFteBiyWh+QuaemiHOJDXJi7S+zDl/LgMVMdrruasRyFzL2CJ9If
jyYWOpl2g2oVg3oXcTBHE85JYDh80jJlJtHinu7DmmHJohkJFJTC37asZqwbYZlI
KUXSTPnX3n3RPV+CPDp/r5x5nmwTjiryqSQJ0xOjjlCp0qojfthszdk+DNlbPQxc
yk1AgIrgqIfQkHgwaeMsT1Y2FT69NYPtDWi0kox2a/fBMFmcWGiIGaN4J4Qw80V1
gBUP7H2M+c+w+HB94CBnJZUZyh4QfxhvINtOEHfTCD6yTXrLWCjmUr8UfiQgkOUC
XA3cIVICOo9KpZ2n7fFNbemDXDIZU8Ar9wRPt1ic8LEoonwQhcJPDWGY2N2qH+wE
e4WdN8mfO74/wPf6eS/0RRXE/v0XIoJiW6TzKonOYh11OK+0UFdeHiKzjZd5jW7s
kFErHcuH7dlEbHure2/3mIwixnoCVFqGp4ilhO2aR/Gv1fHBAh0OwUWZ1MwlhC2e
WQ4cVvP89GA1pG8hQ7halFEGzHxlXRa+oRPQ05HFA9zSWr4EzWU8UuK1plw/mjL3
TQE4QjAOOZFAGWPPgbKStLFYWAkHE0mF05KbqGmVOZsC+C/8oOjcsJrEZfIiZmz9
UIroz3frNa/VU0QeG9c9374NQj2rxSuTpUFex7mSJDtsuaZ4nR6cnNQ1/8giFOhA
QD5qpIzbI690aZVAk3abeNIq/K6Jy+Fro7xruv4FBo1FBJxUaLyLqKBhGsX5fDTo
hVWnSxD+6BN9Ck4jcL+BvmNSU7w19wXMK0LbEXikDHVjmHyoxy0YLLCchxtF7IX4
UOVFJ54UzvF7k/xaYbINyC4DpA6wVSfMH7biEZsUB9k0hv9bswSup62QY/BnNn3M
icqoAaegKAL3Tylj5la9PvzmpW7jsZTNRF/OhE1Nb69ZAq2dllSaEXNZ/W11mj+K
isfRDjjxlF2cDhZ+HghpH2Uy6fFA7JUVvbL2hZ/C9EqZFiWXYim7SN2Scptm9Mk/
+Asb1qpOAZuf6EpvHoXp25lgz/PTEP4ndP1c4ZieAoAQePqui+gYaPwVaWG9tHPP
8ZSp5PIqDs/4GriDqN0If/Ws7fhProg+dqvm6hZqIU/9hY/QWktiGzPe1CiH9AlZ
rKBgRv8wDo1FQxKiRkBCedBemxhXchcCpjMeGO5E284Cq8svR2+/j2udnI5p+vFZ
raGZjjkeXGxZiHwQBUMLmj8zrTIArp4PVppNZX3nYcEuHe3wPNUT4w60Dg+tvo2h
+PRtWq7ATXy7FMGjrPRcRaf75kuU7dkYBS8VJ6Vp1l9zt14ifRtlm0F2Qg5ieK9M
PvQ/XzHLFptkkIu5IDTUVg1a9I/mw8RaVVU/CYaRgcQQ2jhBGsA8Vp7u+Q2F0YUt
6cvOF4NNBQbtSVmf/UdlS3OpDPmT4AgsV/CU1KPpaqwS8rKatrVqBZreDiA29EBm
qPP6mvQMyMzj3POir3trsMXjKPekoeRykBygaLNuCysp7nQ+U0gc/0pJA7Mny4yc
BJgmS/aF+idMUBz7Bhx3GnkxmHfQzS9I/6QAt19TqBtrRQFvV9jOxFDnWYprMacl
ooU/6N9ZUOudg58BZ5Mqcho1uGyHhTKKvdLNwRzFxxSY7zmtPpPgw94rMKOKSH9a
Clzk5l6+5BLDjYr2ov+wl+USFr/5IZeHSDz6epyBlvY5iXyJ1nyyoG7KDpnmJ2lF
GdAEqU48les/2Q0tG62fiaZVKcnb1Y46GlcIYgNXNPMx6gYc0ZQbg+YQ5tWTWR6p
glqGddYP+Za5wYoHKdRDsEJw1vOnMuhy7+KfcKvOMQGeZ92QuywYJYtMMi9Pkbft
oJhXckh+7cg2/3xknevunaQNnXWe13o/dqJT/bbpfCIjbAwJ67YS0u4K7i6HBnCl
9D14uIYWBhnGLfVSGeQgGLwF6qLIPIFEGPKeiJ9avB6UWHx4unFTEWX4UoZ8rzHl
Htq2eP8R9KtHlqNy4bFHH/2lKGi7myw0MWYcRUIixhiKm9R+/mJNOntXvYZXISl3
6hXmQErI9+a6EFL1DeiSIbC44LE0QVauzxuGBRoM2wm8H6sYkzXuZ7r6O4Raaouv
muAXWuCS85w96lse19wgRRkVyjmKlVWiSZLRtKJXNrpZY+DSW+80WKTTFsyALP4+
uDd7OJqG0kSTulGdpw1JtemAQEFLEckUm7QS86rQwbg2K14dqXJSgbcGJ7fVsGnA
MWqSOSiWERUHnZxZuXwm5kDSnvFXhd1dR47c9jcrarpnw1zrnZP4V6mK00x20W3d
rumuEMsfXZwfOtGY9emsMhm/0VdF+a8PZTNpArAsg12xo+BOmeDZFw7NiZ5csulf
oLrh/b9jfLHZOmhZxk48oIiyAB+tC/LtMjbtLaFa1iVMUzXnU7Vu27slvT+ZOsae
2zFbFLv+7XMM//7DDchDzUn1QDHw51Gbo/dwFqSocuqSJ+v7FfzsghaiJ5qEfgII
92KUy77A8WBtaEJwkcN34l64HHLi5/slu/SLJoH43KucWFnIyr6xBt46/enKYluW
HEnZYeYrtmAH61Lr+m4z73jTNGHLxIk9cj2urnT3DfC9SC0xfME4tnZcSXWG/vRm
55arPpva9fzFuo9dFSgBy6uyKBdDp6ZSTMfKcR8hNc99tIqxoVOSrVZh7Huojns9
d5KnTXoqjN7XfEn8wqyyxLxTugkNv+i+DlBPy7wc/BBgWpTV0TyX4JNWjBsHxP9y
Hn5DUDaTf2TMu7OenRzx9qBSD4zEFEnaV2nWlKqPL4yB/nUaG+zoq/wKwiS4Zb7K
WwdjeP5b89xdGHY212XsxQ3IHdmfXTVsvhT24SMwApGRDntY3QHgnnotgpgdM4/z
+e6YpFu4PtJlid3Ufdh0anps/RqYmnEulcFj1CxHhf28hvPj6Xy72pBdFaygsmlT
yJKkuhvxWCKQqngm+COWwbmD9+BsFcWb/ekjbIwEZmRxqsdgSjLxC9KPbhX74xR0
zJXTG7diMW6gftHQB5KerAxeUeQWKSTQNHUpx8zXiyoEJYvm/ZDVsCXxjvHsXBfk
Ku/kyiz6+atK6/DQZsQcbhJ16ixTAfDrNasPOYJhTp72X07XQPe787glKg6AFpBq
dYRIJsc44uucHxgct+5zwO9E1XsplBAZufm4exoWY4xV0Bea2nRCoKLuetsYiGwa
vGlMvS/O50CbJsigl/SLi5MwrCFyh3zPogn6KoExHiLawZN0NDa6z34N87/hb5wH
qQayV+jrf6IJJgpK7nPmr9QAvWjqdGJpQljlfOx2wA10+BYPhPmvfwqOW/ka+/Fq
D1zSAsgwnd6JsFZYQSBIjj95IcKVumfW3Gds2IYO54K1IArkninp0Wd0hUxxZpxs
g0ZP71Wk1uIpfBS5AFb2R1Bh1y/ci7L3B/IoLAOE6J01OpPyzD8yYrWtRt/cjxC6
i+4SeQxj9V7xdrRDi5vw5XivaG0qmd16eRcfovfXuPlhUaw04TIU6hos6Cf0aecI
bVrTFt65w5iInsqsEU5ukEkyKEj1VJuggqEwzxEdS2sZWNZP278KySvr7yKA4fwH
lzV8mWALwyUkv3zcQGihO9bsGDXOVSKlzZI2SFddUAaTIqeHziXlQnvl2XfWZ559
A66FaAnbT6EMrWdVSNXirMaZTvGnW1U4cAyzDZM6rB5WzvT3mT9r34lASfGNZHM9
zke061MdPaTVs3ZNIsbZ9Ntb27D7ukGqRqxzvl6XSt9cXRzH9T24XNVIdlkfA+Ut
zQiLU+fH0ywAJj//lgijmt08sBDNNk6S8TQj0MipVYN14NqTVcPpmnh0F3mAMnCI
3jxwlx+xt0uJdVACyjB+lVvixG7+VQI1pfr3p+6TB9zDjBr/2/J7rx757fyLcxUs
tmKs6ZyqHhMttiCi7XqGJcXSj1Uf/n1Ebv++Ar6IpWU3fKgoM2v+yNFp66qmuWxY
IoJ4SFO0+MPyopoWs5gfNLssqhQdkDRKhjcR6LH/Iy/w4Z3FCOO4wblocq32qMk4
QqeKAGioMbJmkr3lqhBG1gDu5tm/vMNKIo6KTwc0TOu18HH8WoZVmTVVkT/Kv6au
yXYsIZGXiKq8h8KKFRr2ezssBrM2cLDbpYT3JgqyEP4rCdV3pA5oC3O1Izu+nEi2
jLxTmFIQH6wv7Itmdp7IaLD3KDxbN01khAiwBzvv/1dqlN5QjfiVWZx+y4Qf4mY7
3Y0FxpKB8zYQs/v648moLCYCzGbU2vuT0QfaRWafhOZWsqaOCbobIbz0hVM+Wu8Q
Ey8pqYG4AhR2d3pMkgVQKk4DsOija+FqSXwCCbk7Let0z8TvPbvSE3GFaenKYSyu
XT546s2sz6qJGTbZlgd5xPIHCLX6EACxx2e8RE5HZcxA3whrdKFm+/Kl0vSo60xT
FD/a1YOka9B4avsI4ycAMaBK08tI400JAxVPiSl3bllLarpeCK2NvCx/67esXYW+
sb4u5tHtlFvI2N839vm+7FY6eARLZZ/eMEKlmuPoFEn9t6Sc2dk2G3VfqEK0JfTC
oCIGfW4TsGJl1QZMffnfY7hpY6Ryy1h8UmMkEXOQOi2XWmUViSf5zsFjlq/cQGdc
zJsN1qc8LrrkqEhafCerAlJwIXy+lWq2hoSmm68gyjiIhCc+zx2lxZl+Eyv01/NX
oxLR5HZ/d30MbhMWfoxyk0oiaowxRGTS69x/rNoYHokoJLVgRP5ibVguCu8opWl9
w8s4rSFoqUo+WCVpkkAaAiSMttVvrE1gtNlvKQRnsEZqJapTbPFCCoVP+LclS4MX
xSJyfoYtdyxDLuQ0DKal/IqYjEhh6y/7vXQC7JElwQs0BB0Zm1FEsLIOgAks0Z5l
g4Js67J/9uPAsA7aYBlnAeM70p2/1zRkUAVT9Iu1AVCkBO7Z5q2DFLhzIRei6RWL
a44Ar39ESCCpP5y2XI+cYKxGREHFlywFreZLewcps5PO3zy+gW3nppmgXVr1ZBNE
qeyEGLMozNgBWEET1pppbpMoQf6PV5uB/rKTpeNy9Swb58Kdmyk6cr2StJQojAzS
CLj2geESMAVWMG42aZbdyIZwIAIDBV3onIMKPHXZ0IRdX53ah5BpSRpfrLogldJ4
mIp4JVNXqutlOBfEiC9+KG/KYxU3N0TN91xO84gfgpBwNa6yNmEDTqFregX5slCj
RZokX68P7Zg/XJzGSYNVQTRlDq0BhgYTlRBByUM/gDRh2UQ+gLFRi2BRLBBlxbOq
IFShIf+UpXYFSLZI3TnmHEZtmb4PNP6+ufmiJJDePAefw+6gsxG5wBcxJYACuu5T
MqMNrnieVBJzh8jEVCcEzyP1l3+zLIbpktNP1Qn6jNvRwUsoyv7ia1rnaBlVN/56
MBreh3sUhTalyEEaSg7rjHnOAViSK/accg2HjBk2IzELgEP0qKfXYnZq1huz90dF
qeVhm0MAtcDQAAU0sTpHN9baU4zsWlJkk5cZrGnWP3BZSvF3eg0APhFZtTlLkkYw
QVP0R/7Li98ynm/omUzqDFQs/xeHjzpPRMzy2M55IqYQPmW2E1JLV4JupVeZgIMo
CMeAqmHh7zCl454aTT7JC79GWLUlP7KibcIwstb/LFKo+rKYcZ/4I8t9mID8YZXF
Pdk2v5vrsTtqF0t8ILXjEiB9IiOCWJISHLuX+8GijEIu0jY8s7z0SSpzi5yCOA9S
37jdL0prcFkV6I6zgvy8fHFnEsK+jBxgEOrIM4PTJG+WgIBwvhUjvb4KUIvfCzS3
VM5IklOX1tdXUa4QG+iQWsO6Pmspi8tyOBipvI1Z8jM42o/BMJlT5DKh1VfMTMbl
SewQWQLUxqR9lA41EM5z7nYVv5M7Z2az2WgZNe8QRbvUD5BeDuZ1QwnAzOyAVZwx
YJLMIsryDktLNQzOCqnyS+njmvuyxBH1vXv+rRq3c+EvNNdblHuOv+XbrR2/uWvJ
qDnbz7FoWVJSEMXc4dreINcAy6juPG96lUje/yvHTPfV01/HLbE3Qb+6ZFRHgGJt
xdaHR3L1TmhTj3DN7qX54/hlGpaQO1qH4BDv2ufqItOpcTbu3CRrTTXUb7TakhAg
0nY1xWm1/W8rla/gFRSf4bXYImeIhS+AUzZCAG3HRg5esHUKqoY2bo+ZatO1FXU5
34jzbnixrQw/fUR2Me6qqgKrGvqItbzTjZIOfKtUD73c6IqU04aUk9oYu9ng/xuk
Y+lbI50CJ3m9dVarhmRxHm3HtoLloVhspqnUEgVDTLMxseHLIoD+PgBPWmfM3YFg
e061PBnsmxhd9M9Bh7XIG+fkHDbfOLuCLJMrDMYaQUSqd3KXuVXYrelS7OMqKzQ+
/S6ho/QvDBy9b3dE8VgTXBc7v//Z4QoLQQiWf2TSW8fpTXkoB+uOzjfpWCPVYufo
v2Gvns5zDi6hI0EsI7+KFoEkjU4QcFjRh+FmTC7SqEcGXp4g2zpRpZTf6CFsYf2B
yYPJjd8QGj+aBhNXbubpkl6JYY19EAzGi6AiKQGCyxAGkAilo5JVa4peFQmksutz
3wsMDjRqOacldYQWFw1pwp/CjLY3l5Mr0qXDz5uuV84BWpV/dcXUhewaMjfSiPxI
gF92IUmL/WuEyqKINYZ3SuklyZizW1TB5rzRjnTLGLjm0qBtirKo/rWA9quVJFFW
1ICrzCNoOIK0RZKnHQZkdSCPs/gTMUOhw88t25DGHmhnlFgYOjnwZT90AUB+FXAx
GKwvdV6wQkq7Q37K+QgOfPW8HEOzkf0kAyahKumGxSnsh6Cg4WoUhRB8ETvwzf3l
HARyT6Rfr1qaMcuwyub3xJtXglPbtK3RhBpSUULo/WcPZfGlyccH7mJZaooHCmJa
AnQtR8uApyvD3VvWjVPdRImUXtlYo6sXE2HDGfuJVumfe5/+DIk0FFr6jMeEOfRi
QeVn3feTCqipL4mvGcZwKfP8Oy8O5/lZPQpKq2Z+MhadinlKCC5TAWiyYBZnGK/m
PZLEzhE64Z1JdCnMv1ZhH8yQK7GGy2xm/837tHSu+i5s/rO3HGtyF6TwrKN9LJtU
OXvKER5Ae5ddtgak6ls56X9NJu3wvhdR4waxcD54C2j+AG9FizE0QCCc35NyU8H6
dja6F3Wzpy38ZAkNXw4SiO3Vi5uxc8GwlKy+rylMH4wzvxGgmAxfVl+kUm+8JpW4
MuhPyxU0bCti2iFHvScRhfjvvLL0fpaD7xWsCdn0NVXfro2NiFgOc2be0rs1aCyJ
1PyK9XSMLiqO3fCt/k1O744H31HEueYzhkFhGS3EV8T6Nsh5gVMaqrWnhaH52y3o
jPBLX+H7y4Ncqh611EACorM6WLLRo3djQfQhgJoQdvexwz7TZBlVNe1snzu/LjaJ
Yqd6Tf1TvQyOmNLJ5ZJH0a07SJOYt6cld6DCvRh8eTBBD8psQbsHXRi2mlw+aiUG
HYfcmk6bNbDB/3D8EKK6AeLNc3JzdqQHJCTyRF78mFeIgWq/x9RV6EscLGK00O+B
zguG3JJOfyUAqW3zQY5XfiBNTuxFd27dt05AbF+H3gFhQuBoThkttltNpWtF+yK5
2rnFMQgLhhXOoFpIqv412xpl7x8KBRj3LeJ+AomQVpFknnIhXZX4L/kVPWsCJ/ix
1/+mY4OM85CXGuqd4bL3IhjTlkLAzooU0BEuIKcBg60MbxPzoTR0zeJROGSZiCu9
Gbp8GTUwHmNJqJsMVW/CV8120HuwCn0otmvqyMro/r7ju3lzaNvNLHszzU3p12wc
/XiT75PLyb/ZDLtyb6WIfPnItHKYOPDOliOiuJhgjcRU9KMhc1+dX+ouwGB7f1gY
zEvtwpCEcoM9Gcax6+AvNfWGKACrPIquqYzuEni40CI3F8PX7DKE2XJZI2Go3WkL
XusicizK+74aPpkOJaBeD7llz40+ZyT25d3kG20rHNw60Hlhi7k2zbBKUYxJIdrG
4HISZJBS/GdlXw5Dg+7/54trKM4h9R2trW9YEziEoYiX2cSTcY1cipXkyYkOUBdX
l+zl9oYgQE3IFwTuH45vMyOiQVzA5XZaO1o02vnzWFNbSTMG0hjcz+n13JF/roe1
T/IEQOAhesT7A8VO2l2+69kbqUbmhmks1DTvWGAoEdBHbuoGIrB54cOk7ScFlMiR
ZlhG4D3+65CvGy5NB5V91lPt7KgaGJnmuVoq++ApitWWeZ9rAgEv6SjNSQidPbfi
YuHsCDjopA2OH1pmaAYlPn7bTEAHto8t/7eYOLwUmoYmle9NfNxmIgfw4lDlyfIR
WbAVkh1+wd0Afe4TWSKj21/sfLnS/LTKfKZxOuTn88hXbk4mAOVanaB2XJFtLJCG
nMx3KtB/gaiq7UWbKD+uK/EQhmpkiypnHVEtZs4rTiFzxwbUfRIHazSnjXtEZiac
6adXsIPTIYDbj2Fe21KBZH2had87a9eCi3n7+5RaUXhTjMPpSc1fhed5+VIBey4x
bJFqyh/nzCOFlPEXzXwHYfILpHsAgg0o7gLby+AMFpc1q3g8cjvyttnzZSfcp9qO
dZIobUgkCzczHZkwKD/dqfISYclzo6DOOxyl7sT0AQQIm6OhkXO31LLR62GwnDxL
2ur0IA7/sig/hZsjppxJ7BapjWuZ/4miK/eodECKhwGc2kURgfN9cdv/YgoR0UVj
BMExLEGqNd5GTvLn5HURhHBVTUmF5jNGecqryy2Aj2WjOzNOVi/Nin2n/zAtVa6m
C4ii39QZuY9tMqmVH6ls8GZMnKW7yxlb+6jOA9EaOeDLJivViY8G4XgT0d9eB3IS
JHEP5/sm1hiOea2yugsbRiVmwCsrBfuzSXxsNbhu1BqCLT72Z5Gn2Fa0q1jFMsGk
CmoTnIXJa6h6rXS8497+3hU5S+ZjIAyi/zV/nfOdH6pRZijBB/rb7QcOUnBX6YGm
/6oG3ztfjPzOuEMwK+iq2zWkai+lu0a4jL2/XpVT6yhDJRYQFCWUXNO6cSUB3Uls
hMS+7Ttj1fv0+W5jyasv5LZScI/C5a5rdDr3BprSBtO+qHQM66renxf5jC3L13n/
Kps13aWlg8mSZ5Fj1TCOe14XfKO9QHFSDwh/+ojx9Vmd/0+cAgILTj3JEgH0ihdy
uBv8BifsF4O2h/kX7H3NREaGjOMr697V7e2LuNHuNXl8F7i+Z0lqG7CR5ei3bWWV
HJNsux9e5y21mycceickzxSFvhmj8B0SiwrBzeXhAnyreTfc+PALWZK8rUrw3x76
hdvgqCf6fN4AdPeDtG0IdVTdesPr+CQWWTGn6vZCffHNsxNAAwRrhaSpCvDLys7Z
APobTCas5BMOaomPODSO0GtqKS9/f04v8W+qNsNqcqXC4Bf0S8vo6YHjsPUWcRAT
r1xfzXLbN8UZeReF5kBHNsKTJuubT9RLEpzQBpHBFM1euv9rypQmz/7HYjbpp/ru
H5Z8MXxBDuRPXHDLriBlyOV+pZMfQsP7Cw4ERlWlK5Y0xpzjfecdU11fT+1u+4ox
orvaG7rgmviRDJ4e5nMK9spvJXYkiC0l2cjgQfH6rCW5ZXELS/El6Z+MMOYclRHP
QdDQ9e+9QsdyRbRJwYCMzYbOv7JT7dUkK9xP4SpEGiwyAeJphgh8KsMyxNIR0CKC
jmeAmdwVRMcCiQ31WQd3mTy7XHA9bo/yLpC+MmEGT8LjCOxXiT+Mh9rnD2//iPVv
h3SQI2d4/bc4dY6NRoV+s3wDQIcXK9TB2ULaqDiFksKcU73Nt5SNg8EyrhmgJCLg
KhXzkRsYEvAZxxJxIDlUld/STfvfKfLkeFwOCm2ZGIm8PenNlaQ6vl9OWtfjCZ4P
AYNlN7W6IU+zNs5Pd7xgg7g/NniQLMLx+LYLuCJzi/vpcVO76gmXzATlni0BOHRX
RhyrGXW7bXcbHj4nCnU25wX7lqMhPlRNUhIy3onn4SW8cNYsqW9FUSz2jxnrJwBp
lR6mEojtpM1w9fM6jUjUmR/D635L9JbAPs0a9fn36EoVb2s7PvPJieWMTwek2cnC
OkuJbicuAIVPimRJydqqi+HvTsrkRK7JXZFJoZimXjFCZV0AI8ZSYO81YcM3FK+E
03MgCWJJ4Zez8DIXvRdYP1MWMbRNmELcG7UCAxAjOB2FgwFBkoE6/IDRa+lBmlZ3
3wGZhwTxeKrekrq7YU4eUBweijNffb9igoViR5MLDzWtG75iCm/wHMtA5WpIhotE
/BMCWwsxrPxuVhMlhLTeHLfVDyx8UgcdXOipvzkHLzPSI7OstDwBqufzXLJIyab7
7GIVCtipINsf1ZJLltV7xkIuka+ekcmYLUFVvgmlBYNQKXHBg3TkT7sKkmLFIe8c
23hUdvSnqIBHnICsSD/tUJ4hnAGMQRhtJiu2LRsNVPAXzkeApYjWebGtZglcRmp4
cNrintRs2P00VC47GZxmxeo+w+zPrOfFLf5Zdu3+x/31ZfS9GxMoQgMwkouxCcP1
/S/JSfHVNW4Q2l43AMm45ulpjlkOgnwK42FgQgzjIgPbXtBpMxViMawijjurCDcL
/meZoH4YZL1AsrvPLuylqsy2hkrMmYab/bKysa/U5IwS5jYFxhHOJqw5wNCErhlA
wtMnglTdgfayJF6+nqJXzd/rrRZr/47Wl8Clo1YBN7zw4qIArvvMfQdkAcEU9gaA
W/q5tBqmW0jvM5lBHQnQcU6x/Mj9OXrkgYS0Fc2mwzPDTwIZ0pRK5LeisuWTo3wd
+nN56c3JrU5DeoQ5JhKSE37ZkALWwdTa2TS6L6H9lmVRUnF6UVwMvZ/DayT5CRod
9CjwjtP09pCpopmy5Kh3UjLyh91DwU3Eg8zILKci1qg403zE+AB8/jDVwRMxU8Lt
QyxkaEVcj9xU9KEgMrZxTyN0IvmBriJWxE+cVIcjtJtrt04U4t0JgTiV6FD4tym+
qI6xk5JPhnuQAxZctZpOjgxscumLUMhODXH17RaydZ9yKP/UZhmjB2eKG+8faaE2
YwsjiYPU+ln84V7Ugx4u9KyXBOfm7/+SAaHrHRAdtrLSx9Vwfu2PzyfFmsOBbZOB
Fpkvw3K3sWmJ8K4y2orpl+Llbk97I14eohmHh/JKcBJLkVJfM64fHS/gXty39wHM
CpsC3uaYYbVrwtajfMrfcYDjsttnXdhnEMZCNwAILApHQHiJy30YNZkULLwTIyeQ
50F67sunDDSCLCLNFilXZVWsT5Xk/TRT/z/HapOuepjS6mD8GMVlpXTwOMPkWK4Q
GK3INk4hlIPy/6X8sIaeM5AOQF3AicmdZK4qDwXhOQVGh/byFHosQBMfIe2tb9V6
C1Th+C2SLz/UGL3qFv6LiFFPR5JVBwqcG/16oLM42wcVRaoRXz0Xphxntm95bHSF
kwl4YI4gu93NjB1sLdoop3V27Sniq3KB2H/pjrAilfHOu/wpn6m4DdUj+XcicMnb
EDRyDQM6F8vKUbY+bYvuFyFyB4C/+WyfYB++ATAbQOxArwY6x5QyOloEkAtTpPtU
f95tTBAefZfRcvEqFBAKuFFs1dYpl67A+hDW+yCxuE6m/aMfR7+6rEEVczuTmeIv
b4FFerx89GksiMrWM8+5kl7yFCcmtHbcVjsQ4coDRjVKKgiWJsXj4pHtjJVl4A8o
j1K3tQsCiW8yLLnrGw2JvIDdiLm2QagNcEAsJv/KK8tsrEUD/iMkLFNHI4pwX9+b
WfqXg2M246DzfS/TFxQ+Dba1Ly/wn16EYu6OjWsaZyH8YR8FVgdoyA7NGLMn903h
Pvt/kXzFI+iUA3f4NL+mYrdtLFAELcY7v2noadC2jdwpc6g+04iV8ScqxpBjvOpI
hwz4snAQERJOEh6csZNOtwV2W9uH2Cm6tpdMp69P7CEU8rBYsfi4wzb0aB2vKN63
cYc9JYeGS+Ky0N0Fgwk40sG+ggWIrCYJF6fIGBaGA1o1brZpRld9t4A3xmYGbJW1
ux9fIAzI3OSe6B9dQnv/seeNKUpG2bEr/iFgiLisQ+yygvgTFtxJ0dp3aqa2kFAC
60I0yjTxEXPiWQmWilhTuAAcmbLpp4FdgUgVQVCXgrf0cHgkzhoYL5HET8tMiPT2
KsQ9MC6NL/Amxx0P8Jxp4/TgzaP9KLwySJJbNXVUq6RMVvf6XIGjvM5N9Cvqky1C
ywdKhN8/ZM9gU2Ggxx9HNPDq8gfSTA7ieO56RTWtu/YrA8MPa/QlvDEGDTOYHAUA
Xe3cuGUHHeB806EGFM9TMURE0SkOVohnIX6dkxNhvIvWcjmixvXrIaLGzQTb6eBJ
NNI/P5ajxxObBw9Vh/Bm1lPv40OWwt8h3HiGgsvi+7gNX2l8mT0lvlb9s1NfoN70
bDfaV9TJ5oAgazQvmIzSGzzkCm5firT8AkqesCcVjYCEWkHa8iguS6aYXTzbLW7u
23sdLTLhIWuzB/EeWPUGXIlSBWtCPlf85D6qHxZ2g9PznfM5Z7AepUTxjLS46KoA
tejj7V5WeNi61EKqh7hMpvHSQSNXSd6yhryPnKZnweHGKFGXstL8ANHtVi2oY4+V
QElxComWGiaHIduNCdr/LeDMR5PgxATLG2vxvPuqZoER9+IZcW+3SZ99yDWLVbSp
WhvSxz7x7CQyWEYe5jOkqevg4+QBxi+LkwFEQ2k3BAtnRZ7TWjz2q8MSIIj43pwF
1VtwZHQdn53HmK5gL0If9RAlT2yx01FtQVfhMognrf7A2NjlUWjozQXXMe/lJDVN
dT2qf73UM/DRHRtWZq+ZahJK2rJ0dYGpNazYIbto8weFsuCYiYhn/0Jvd0QIDHI+
rqW5UlGDUoEpQWcjQ39/FV4XxmUojSH1hMrClR9vH0ObtXxFa7nde8zTkeTaoQCQ
+4uHNewp2LPsCpnNasV1qRtCmVUBW2qEW1DWTEc820SFMvzwNzBxMF0nE4LIENIv
P7JfACVMApaQIlWwm+a3On+TmYH16//JklO78fvckMBMpsfoKbFJM50XwVhAWsoU
O5lEPo6EzgDMBbPMKK2cpFM98yh4DmTu6OHdqQ6rB8imUYMlP2s3sRAkXR9Jv9LR
U67xEqseg/Qly6BBC/E+XzSxc2ylDp629OfcioKqt8Nuc6BCgSzgTnnwGnQMKBJo
yD4cBzhr7a84TnVdTn7VCq0IL/Q32gdBKHA1oZVd0BY6We64HTvsbLSwVoDRo2Ho
wBqy5wvU4G8nO2FKMwDVbZd/ib+5aaChiSU8exqny/Xvibf54I3l3ph/jQ5Bx3/S
kNw19Gb8IIbKE11+7iKdGVJT5Xij3GiVWJ308b15FYUHx1xO4yS1AhI8ILaMSLQR
VcFT57zp6KxlWBBPxBdyl6KXB45a+iZzPR3KvQqVv60BbQs4iHz3ptWRTh4YApJk
8u83ZzQU6xX4miuiyn5tRRPSy9z2Xmt3V4BwksSptu2iOw6tB/0uY1S+dH/yiaed
Nl60p6d4G4Aib7RsyHRnNnjG5U0nin5RXC00xd/AIRzfqnXlzRikzLJ3KyZPa/h0
ds8MS1KPWJQJzMOlRG5PVIsM6r4zbjAeALhtp4seHTzFk9mkcakpFWaAmizpm+F7
mlXDMyLFIH5ATTbKtz3vHClxJS2eRhyWQBiCOZL2tb2jtr6Sq2Mj3gcfgtlPpMhF
xv4EEzfaYLlFmg14J3YWwufSbgmDRMS+9HcPi+jGy/zEBTh+fM9/03OURjXzxgU+
Q9SBNtUKGC0dfWpTYEU/sUpICAq0kbANKgn1BL5Y37rN0On6n421CM6NjPclcxOd
QjjZQ1oOPu6WaAac5Y1QgOSDad0fc2AySfYjQ3qnOy73KDZDAS/gdZcyYl5Q9mIb
XJr22DMMlZ5hH6UeAQ92ELbsONBNcH7lNjtUpnZmRkhKPeXdYr0v1MZpJ4oj7oGW
/mWSB9qQyOZ2nb0R1U1AFHVpmqti6QLhWWzEX3LkGiPDNZ49ZSSd+cBil6H4UpAy
Ll/x4K3e4FPxcwPRW1D2HjPWXl93zO2xThg58Z/+F4LB1yjMfN4vwUlX4A1ihNsE
zKLVbLE12z8Z95BWfVeKIyxYrc6F58JpEQlcJOe2EagU4V1d9Cy32PfGO034t8yp
rKpPPVdPSp1ULuwlx2meXt507xlNg10LZCU8kf4Q8DFDOjPzxhLajcdK0p2etlok
B0nP29mTsWhObwYQDAvYEqS9ij8EBmsmqzZ2dlMzOydxKt8scuCX05oyqBChbgve
kpoTid9m2Hulndka8EFsST/MMzgWlade28dEbWZ+RStew8dGP0zb4FGxEfAVNRwE
8M94e1Nxu7QoWvqY/aRc3XmoosQF8563k3SDiFHJ3sjBhVpTC8VlqGyZ93cRliod
Z+uUh9HF6NBL4smC093OA54h9TlJMv4pwzmHo9HT9H70+bWTwaTnIeVqRJ0azMwc
HGlIjlpegdr9P5+cQzdqfx/vJjLK8t10YvJnZ8oTXHsYu8cvTQ05kJ19V4MYTcy/
8G9IK7+4XYmBQZXnbft/NwPyFjHzaRPjm8YvJlA2spFvhjlPzyg06kxYTUijmhJ9
oqgWwacowjJc05hH4MM4ZvPVESTmPv+ibUgAzTfZOO6f8MuaDPxO3zkVzQz2R93F
L5i6KJ/R45auIfXrg07/+ks2CL5XCbPmgwmSs/tiAK5Zpo/PzENfFaOZK8m7xLSQ
JfnzfgiWFG5XTStcf8m/vxFJjNNqKKtxYJDrJWAQ7jO1F6AEJZaEmHyrYGn6KoTD
druvUHaTcxOCVwHJt7de2eof/HdwRCpu8IWiWDoNxY7gm0J7Y/3JHGHXaO4ifNCj
5g12Bqw2sp7a5X3YU2jooey9epRGM+woQQZGoQRUqfW2qIs+lnvcdzPHaq0nFirQ
PeRaI6dKoLs5pLNVG5Tz+lPlk3I1TCd0Zd/MPrAIIAar/f94MZKdADKcEk7g/SSI
c5lrPYyAoaZVgnm8preuCvIe7z2a++D4KVmNSXv2I12mtBPoUjLVbj2GiCIwjoSF
cwDWxrE34w4bpa3jIBdudOXwZpwqWPxMRcLM/WvClO/AQSbY2AcNKSzFKcJJ8UFa
9+DfkKbf7bTK6vCQgFlYdk/xZtJU3ypIPnKvVjDdfRoi9tk+FxSsoltb06ZgDkXE
aJX/abVuH6hQ8Tmurn1k9Lc9NMCMm2IjWFUBfsudcbDFiPssq8jFNAQjGNKryY+4
I8Vc4duDOGCp3Jlb/8miJhb+4ziYx1EzS+o9+Lo8IyEt6o7CjiVQrG3zjohv6SXr
yguGvD4CLZvrPNvbHQgWVnynlil+1zqm4KIxeDokw0ro3vdc9Gub2Lkhz/jgydj5
8/ozgw2laHvfzanCt0WEgxRHuan3lP6ZywgpCoZ8xMNaLnauzGx+jRIZehufYmNq
Njm1OfvFsENa6RIqZAZQXi0An+OCE5j347a4ztvsJQqZAeN53BTCaH34YOIQ+Hvy
wx36prB6t8ajo/wPzHnFMcRHgrnSYG34MTCog3DSToOjdZQukHUtHON1O+ncjY4s
HYt7LpB+ZOyZqr2HARESe3gtY97iv0fFH55DT+FxzRJ3aWlp51UlkQM5VsmbRLco
vgCP9RSjH8DBxh7cCHGH6CexGIjkm+zKkukLm5VkoeMe+X0Y1OZzwqZWjCkS/XUk
kpC2VJ/pYBb794RtlG6lnCX33FNVC3Zb9bxdcXolRKrf9kIM0GQeOB9XqLJY+n4I
DkfH/pdQxKM/MwA3+rgzmicGbTKE67Sni8BaWg2qqSLLAGuJocy+5I8+3WMrDdu4
eZebfrlJc6amO9UF/ZiPGemwqL83mJpLDJlnqJtYCFwv9JbV398lUCRffuXPq0YM
MZ+vZuY2oHPd9yLWHPL7BKORfwgS4xutDFRafhprwq+bT0rzWHvNrmGJurU9aWF7
nzemMB73GByPMNP4fAh2EyhEvbB03DbPocWQdIJBuYRU+d2hV4Zp6rRzZhbM20XV
LAPb3pMUPvrNxbcCwkSufbcqaKOLrt/F9UrhS2QHSb6yZ7kUcoyC+IqUovEho+E0
SXcIui3QnnghVH9LhEeVdCqdhv3izPWQ7FWjEjgu/07nUjhdSfMNXO0C8Hmy3D+O
kin/otIkGw/PPkmYVJPBXHF/3WypsyMTf7xEj3N9cHtuzrmf3Ra5usE9S0tFNJd8
1a3ry06hnxo2g/WASBhrCt/ty5CwKZjz/MoHirVrqz8zoQpZiK46GjRE+g6DqlWJ
swnjIFbVf3ds8DSIix39JHxG1rRHjP2/KGZi/sXfbWzPkMBZmM8tyAi6DZVx9EsQ
Nw4ZKovjn5zmLW7aLjIf0ZYlSF9tTtuaPbmsxUyJD1CYtRVnr3uJSsxAMv1PAS7S
w5W5EysJ8dodD8jDWxlkK1tPeiZUidrVE7yroq6QiHjEUfcCVJox6ycDwswZdK7F
ol8x0IVTKiVhKBuUFFoasVhb0EgZw+vAxB/qaptw09vlY1avHPdceHsgHC4E0P3M
K2Q4GQxnl2pubPpLkEeKmmoAsyOcNIcjj7VonEHT0UidCIzstagxHF33yfb9twYs
Xx5G0vUM6J8tsTg5YGYAfIjBFg6nXRZgC+ur3GLe7GCAlm7m+HV9MBzJnVX80/yN
0LOrmLkVN6HB6SZI/NwiXrzi7NSMS0MGTcXc6bBHzjPBTE8SdVbSpiJj+QeLTWot
ega1z03aWDbey1NR60zuEz3zUc9wBcEjZbr2zI0esccqv9uYt9xIFzj8lE8JpXh9
U5e/K0BJHGKUx85110+QvNnfeAVwZe4K9TDWreCfbyhRp4mR1f1vFJApZXsqDP9w
d8d7d/k8kZGuFLDdFyXWSbI71hK6L4rEGxXlAyueMtPe+5hoIw7VMNM+inqGwv6j
8t08ByDK4imGQ1XKTfnccsagKkUi6ujM3vHiWpvzPjvFfquh98Zxxlm6IoGrW19n
CBWSD/knPq+ESH5eTMRHySBniuc+2HlvWuFn3pLk0XptOg7cTe5bgFlorDw7Fsrb
NbVhwH+LCr2puFZfFtpjXM40IfnsuQFTzH2aQxEWtMAxG373itQWL0OdtC3bSGLg
d/j4jM/htCo9zGUMshTmbAyuJkUrSE4dPhW3RZC1Gc1qpAhD+rFLviR4QjDKTAhO
lCx3/5duq3eZ2NjBoWSLpoRSsVGtVd+jBc84o/OQ0MD9Wapc5204H4QEuy4Ts6SW
PIynukO4mmq4Ch0Zk7Uwn3gjlISDfrb/QMxXn5YpH6MK21Xdr/3CKZR1fwOJgUVE
2sgJyR+iFQfpmLeoyg7pqhe8blY8G2UKgu+WGnfD4UQ3zQLen0zKxxsgcQ3C/7o0
p/Za89jwmI2RE/r/IDW19X3a9+BPtwpg7MMZLKFgvZeWaDDTC3JJgHHI644ogxeH
uguwtawbV63UEp0Euar/qMt4B/7iuOAxfwy2gdTRfewGnyh3nSZnD8CeQWVxzwIx
Tzy+6/tGDkWZjFTIkyJ+jFLhj1ohCsEoQawvSth1glq6NzgG6d9CzcSlyA4/JfcM
c9Yp/2saHhWMeCV5mIubOv4Lhk4uQkjqDZaNUcw8JMpXtSW3kj+UrJHKc6ZFy7O8
670YEzHjD4AcIjHIW3dV82Q0SMFW1y6YA4mflhhG4M+BZUeeFn7a09c85s+u2GUr
/0n/1SAax4+q5l/m2tJj4ZkQ6icpVIeX+LbV/1qnI2KpOX4prnC1lvJlTndxA6m3
Go8YqCCXVGshDQHQtMFi+JWYSxWC7DcxZlerPZvVKhqxRSusJTnEx3htVT0S/vM9
r4v3Vqind8Uzw9khIFQrO41hQtx7XDaRpS0MoaSzmJYLrItZovHFKNGjvidGyGLF
ja8UJYhs9fixmc0fgs3ms+g25NqJ0Yit2Ye7qpWuEcVWXwVGdcbMDfyNrv+n8KFa
iuaaD92ER0kG1NOqS2vL6yvEYUgEbQol8d01HnmIY+dXmSoJBOPw97uHc/F9sbmw
g+7KS9PNs4KQQDmUkfiwuvp9IX6b8UdJJViqNEVyaO+/mPC29widwwR7OZg6CCNf
BMd4L/JwsnakDDQJkursqxfYJA7H+tX4wPrLDHmu/ztj9aY9Zv00iBo+YjA9HMsl
mS4jzys3k3Bh3lFyKfhbScl0UIlVzg6OCfKjPYfyHD/9C+0YceKkNKywQ1/d36Jb
yLzvXS84HC2UEw90+K7iBgJyXnaMg7qhY+tHOXq5P5RGTT07AANfY4WH8ByqK0dr
kBxeeOQZYE1yD6IQt1hR6nwB+DB1axIN6BTQ7MZmmbT0DLO0N9F6aGs0/qx/pqB1
18dkqZoXiTBMlzQC39gt+voBeCsjJDleBlv0bA8hEwQoVmhmhpMowfN5qQKH2oLA
1MG3qPwyMRDGtIGP1/V23qRGQeQ3GAxC+mD9V1bL3dWmwTsSEEV6SHJ44cVVun15
jCWN5zIZ5u77MawQIuakJBuBjpUENbIq1x/Krp31hjgQQX13lTVU49zm3LXh2wok
lb5Z4W//016qd5uNbEVt53GgOC44A0hYBPIphHGANehuOj+caMnswCLW9hafWOtj
E71Lt1xuWwOGKnr+Cq+CrKAd4X/6NfrHq1wOsQDgNLclqLd3oL2mNdknIxyLi+9O
+3Ahsn3RopHHP087Dfvmko+Eu+h6wumRd2QkpyqSwN9nopGzEx50Ki8r4ipFehxH
57uiIWxqZGFeIv0rd7NSlfA1vrh6YFzlD/FnXL+bSVICKhA+OuM72wVuSpoV/9ZZ
AwzI9cbm0ZkxbJE6335agi+XkKdvI/W8Efk+/cQk9wnF9mzDIWgmw3eOpRfYq2hK
X9TxzwJdaCF61XG8NSwyrzUfurP5fThrOOKg/RoOABMAnxUhe3mqN/d/1gtouo6t
GU0vVU5RQBxPTaJxsiRuj6KCsVdhQcdbZTj+GS06qwqhg2aJ8C3aM3yR5WwYASC5
5kjdfRFISX/x9QJfchx1CLmwF+WKQLbJMwkYa/TbQaMHBGH/9lOc8IhOAcBaKSqa
zWG2PKPVzc72bBmzO2gT87+9MDGzm3PmUcL2VPOQH25u5Pq0Jx4bbbB9Fy9df1CN
u27tBTW694+4/qT2tBjD73jHTaisnMi0lmXTfBxo2+z13qJt+l7HxrQsp/G0WbUB
blbvyQFggUbC4ZkdKPDqu4XCvL5WgVcNMdfci21n1j8nAkpGE5mOO+LtcaxYO2oQ
g6j42aqzbx/p/QJv7osz+LVqsMg3R76DSkmpul/E//Cxqq6B+IvpSHXdKtVtexrA
nq1tfm3xhoU1cZzyp8mzNwjh+rZvE1/BA1gj91v8SifQ+hYxTTSFmOH7+mCrcNfU
84jLKLLmQYFRNOXIsOLjFc357Ak+LLPjuPV08Tl6gOSE46aWyAK/qDmOAP79WK/i
iCfnnQOlu25bzdwVJOomWhFcT53m69zdL/PfRLMa6YtXkbzGCSLWRhieEBH43PGX
mVGRtJUNOFKjXDGwiARSVWCFTAQMWIZUzmn3oqtzSDAuHlEJabbabUVnfA6HRKkc
I068d2nZI7aN9hxg5QwnLOYyGVk5lJqi4pV2Ofoq2C5WVQccnuHBVTXageF++6ee
THBdBNssqf8/DZEZadEXP7aPR+g2L7KbrflV8Sn4bYT7zdIdntQ5Gk74ffja8QvI
PWC66+x0nTwzJRpk5J3rGprXOObHYZs5wQIYbFd0EVDysRuTpzqYwLCUSPm5MHGL
PWHnyjkUBQniEJr4PEpIO/JwNn+gVXx3bZOVAi/eqpvDSHLqt2FOCWRaAyurnaeN
xpPLm7GqtpplrhObJy1/LCoXFSpHFjlUXu6Bc5H8C4LlvPbPJjHq6HuZ05RIJf1W
hLLxTSB8zaIVH5Ky7Y16feRCXFWYObPZftj8VMAS4CCsp+MBROBjLY4wR9FmCwF8
wVNJ7GQcqtHp23hh05y2W733/d2kwDVa/FBnWSUiwOgX6J1xsc0l4jasdV3saWOb
Xs9rQNOau6cc8TwDofc1ME9NKb0FF6nZdi4oD9GeR1n5DVMxl6Vn7GOdrePh4pPf
PgOwv6gXVSx0lkgr+feqlY4mL3LAQsSgsGp3zt6S5+qa+0igX/X2nn4eSRG1TbMl
3eTiMa/yy2Y7cU/YT7eInTVAb/3PlPj3RmC3E5js3+yFVcVnJXvofPxDfrjzYb4U
JfKyx5Uq3DvCTbnzntnqeivOksPQXBuT6SIdJLXIRaUsgL6zMvUTZ1W4o3RuBECz
5kVQJK6nielYdcHCUpZ+dVPpF8jq6gZv3KLW9vLRmZ+v3N+sb+fK1kGIQ63DGZT/
Tyq+2UbC6EpbWpuaKWrtGaV5pMTTjBS5hAFjKx2Gr4Xx9UpARmNOcWeOx3O+lCGv
ktLkMdck7/h33Wsz4WTy/l11otkPVCd3jMgXENubagDpH1aLh/Y1YZ/rbv8vQpte
rLTH8SbBEmeerldKMhaoiIoofADCqfM54RzRJPpGuSGz122hhRfYgHZQuAV7Ya0v
MZ94H+9OKEmq+svyQBA6Vwj2i630OBiKDsIhj1MIJSXBO5NR/b5SRZlPMyVhciLK
t4L5H6a/CetYqz6C0/NPMSp4m0MaGZekBJqyfK+Mf9cW7UR3u5lX68669+Yo1D9q
yPNAc6cNkEmdnqFN5er1OOUB7SUeS0Q0ooHveHOUqiwrmxqMvexNCmV1y9tC4p8G
ukgchgsiCY4w72vE9MDEGDgxJQ9grfhP7p7gBypxfY/h7d0uGxiGWQ4O0tlTNpDv
g19efJoTZBe2ov5xqzjx7D98tUeBoNX4junuNodsf5DY+QobWTCcd+LbO7ox7QbS
4HP6JlQBm+1EGf28a9qVuFaF9Bqpas1qcbszFgB8wQ47FqqsFGvnLKPZkOEvPhDk
xiLDMHqqOnpzUJ236drWrvI40Fv3o3myOZPATU2Tnzv6wapr2BnlOtpD0uSzCNXx
picucANCybHShtSDmuBCbVZ9Uy2aVqTsWcoax2SfI0mgvFtfIkdDK1cUSLjnnzAt
GALGreD09kopqSfuPqH0tl0mV0QxSi63754018u12n9kr0ZYE66wTbDIqYFrUQXg
LrCT6J6KM9a7phh8YkId+aZU7TbDXLYb51mZKfnhyABsKVUtkSeeuJ55X3O2BXX2
i7Xq+RRrLEXnyQk5z0jWqQrFNxsSWPfr9i37Vi6uob5sxNnSzA94Iq1QMnJeTXLu
wiIvb90kQB7jXczekHO15ZpTMsEJ/nT+MZ9bnp7DXq/48g9zfrBoBsJ/6SnqU63I
fCPGMTZd4Zuk8XS/EVbg0etR/lJv7wd8AorU9Kc5RDDs6OrV/MnRzwXqY1zBCYY0
fUDcrXeKCwlOBwU9XVIyTPPBZ0IImNVj9so1o1odl70LMnpvmCmJD2uKe4dokxpA
tb/Pr4hVquV6bTYIqqKt21dX7VObiOB3PWOc0u9iW38vvTKi05Ec7Zw0Y0c87/Xz
EazCx2oEeCmsmaaKxn4XUAStJdGXoZ9Wq1bBw+f0r43ImbVb1AzLpN2+sRXNk8/Q
OuUe+Nc4BLoqTZCuB93Px+W7cWgRVvPCZXG9fdhQZhNHpHGJ/eW9AXxOXCFTyRXI
Y+0sPZ26fmddx+gOFQOQeElocSDT7yoRrKUeTEOztJoqxg76SEFy66OupWE6Ndby
CJSL2OhQT1+D2I1avy0Aga7xHuP69UIO9hfeB0kRDdHR5CWAzVXgnSkKERr/P2pv
1fDZqiDVv1+qAeykjDodtPuI3sL6c8izgCsjD/XqwY7cOi2DlDvSXxgIWZAWeVfL
Tf2MFe5bO9HyFfbV1iGbjwC38gwGO9lvkPkhBUb3UD0hbg4vh5Ahzl32o0AGTIFu
jVmGah5Sm4J/Gg1G/S7cWIuMj9cWNwGizEN4365m72C7c03KORZQjv7AzGNS+cru
WZD63hoK0cD4tRSzZSPCscczZ+qahMVX4OYkykmKSYbSwjW/au/BkqYc7NGvGz+D
o7y7fi0rpCkPxuAbEg7wn2QNfiizph08LZk33+P0++QqBBsynQQk/GBkVxsRdIT2
MV1dlpOemHCKRc5N+brSZ8vAOIQyaYNt5nry2AGSPHHi7jVDgMMyYAQ3qsIW/gE/
spSWTR78VzXnrvWJxQdlEPU0fNNm+g528GeRgK+OKy0q+Px/DJ1bhKqnAwdhjfGy
2vER7a9UpyejSnC8egh8WZausx4e2T+aJNO0sFv0N99H8biyt5kBbiJPKcy4GlmS
sEhbzUUTe+zX9UdpQv0IyWC5exbSzmwrsAyna+6FgPvEk6l5+zUpDLB3s3nwKNjl
TiHrrmi1wnFeMPgvvi3LxxnRws67AzntdcrBDuqEq2t6Y8AlPSgc7O/dB7VmTcc6
XKq9byCm5FdLaAyPkShbQ1IYHNdhKmgAMicgBAEz+tHI+sdzxHl0/oq/5pCH/sL9
8qfCYaZcwewCA9pUWU5JKvwv1llAltoQhE0/Q/wEiVr/FuoKD+Dq/DsefyH656Cx
ih2w+jzmRRuBXBDGKkoTyAmxUr9JJGUHfVm1lcDBQrEzWTXu8e5Xwlnf5/jNRNG+
BLSDhHUqHalyIWibN23d4bfNzMKRVHX6/V3l4LRzEsuAdaF+0RdPNCH2A5ap9rPG
tPSVHAN/FQDB0/kc2ZvjnxT7uqJYoZqUuWwPdQHFFsZeiP0Of0uzyAt6UOvSbK1e
1jyJuTw8i6kTrwFvHkGZ3wbCxJCwjY5o5lcMfU1AO+82jCsqnwuEu5idxONZuMl7
Jfx4PlsHRj7T6zNS/6OzamOb0FwBqs9cI6usQ9XrUvq0X+hmJ5pHJaq0Enu/zvnE
E0MIdQRisOqDnkBIGRueWD9bgKgOKHpIuls3Y9o263vqJcV5cD0foH9XLslGX6d0
+0xWnbagdpMaRPzLjJIlxwf7k70DF73oi4ZtC4YUF+PEKeobFYi7PFvEeoX0d0TZ
Fhf11ZzPQz7K45MMStwp58GTw23MfKgmy7sLfpf7ioy/L223Dei5QCrz/+IUZ1dU
ExCQpWeHZ2l3dh14bm1CFSd/LhZhmbdDuzkS3DBsfYztQambGGd0jGKonNiPkH3b
Tkij3zQn/BBX89Ton0qyUgWkJydaTAiiBqmFf3VQhgszxP6BLOEj6x/SO9JWV3KL
SMgDqa30yVSQ0bM+hxsFeLkDRFdH1DzS9sLFPNpUW/aJfao1pZcgP5UidsBrsy5o
L3j7MlggTX4WnFvuDFw7ZZKkrteIIGicJ2TkRcWX1YhxnLi4wBSoiQLs/jo832D3
vMQQUeqfXyBI6Mig+SnQk3TF9Coz6El4UFMvkgCoFSbmxSbd3gIBY2VrWSBymKan
YC2MCtkATT9xFsFTfmz8PprLbnm9r42x6mXi1fx7CW/6CI18SsTyQih/DDrsR3st
YCmbY3STe7k+Pr0Tsv3SclRAKquMtHboc43p58BtxsRWaIbPzc+6m1ZwI51+p3ia
ON6ufrvK5DXLWPBRRXdNsx0QnJeBZT8dbchpf+YXacVAXijOcQLR+9udp02ZG4wJ
38IGrccw0pQ9WncwTi+5cHMh1kISOLQsGtLQnp4P2tYaTaJ1mwfhnZ4uStUsqC4u
CFnXv1Hf/wyAnOh58pN7uvDd7UmO1jV4gI1bu4nqmm7Q4e8pA3NHeZBvcQqE0jAc
z4ImyChrLH2PRRib0i45z1bALp6eLmnu7lbNnEtIYSGEeKwgdxVvhh1M3uqZkHCv
PaUTWka/Vx9iv3RPcwxpo9ZmquYmdgj4Ny2jixZJx1+cWoYojn+CP83jvjj/on9I
p30qYdwvNTKuNxDdv5nVNVkJRn2EXOIuIQjGOrIQSogcDzSYuJ/pPBsJPpgpIRZB
fJoA+iS69DZtWHe9THfl3/qUnRFWdHP04cFCTI0ywgc8tT+zydVvyEizH6IY5pf9
3u6DxXIH9m20RRaMH9Hyj6ZMeliTbRbDN5kRCb9K2rFl+XoEUFKiHVo6l/zKMaWc
0QGQFxsFZFz9/e3reY9lFtYbNpgvdFfIrl/0Xo7wqrrMCMlt37mw64AXIPh4M3UR
5IH6kVxcaF/XKMgTjehPMB6vpXSBv+9ZJzpcxG4jTqwIpsdmv9i+/5IjJP88pjLQ
LGDfV31KFX9nlURsQgCEJIeQtzw3ZLQjlYJ5deEcGVIFf0JNv4IkDWaro8vz17rG
qh8P/PZCMkDmHVMOHXKDkZkLvBzi+RrizwSCthCNotXqpX5O7WQlLulC3qKIhqkf
PEQvRGtT5gMUVKDk8Z/RMGL7PW44lg4hsOUWa6/Er+lp+k0rqwIxJqYGZvI/W7UQ
/H+xnRc1+X+Qhx8nCfJK23PyeTXOYhHZWw2BwL+lXGIXVmK6gIxY5FbZOyYwGXiV
EagGU3+iHenLwyLH93pQGsMH3p2jpkDho5flLnTu1ZjDYLN5nLIiMu+1oJomJr2W
Smw+Xcj2S6hjZHzFIJVGNfHY/TtPtX3DOriobEv09TmbgKe3PsNjlGk8ClBrWrcA
zBzqX1c/RLwI6Q4mpurOXz2iMtVv80dCHS7O/vIXYuSIFu+RpSXcR37r2BiQKwgN
ZqYK0lJX7jC44fdvTC2CVqVCiAYMhZKcDqen2U24OSxWAarSLaFmvn2pKKt/pELX
Y/XeVctd6ePKZRb6H/04JMdZKmVcdwcEMBZO4+Q8WD5uvsV700yVRNFXZHa0IlPA
WUOw2Vy5WT8EqAbGTTMQYBoqj/ZlM26n+pb18u2Ba2ER21vd1G4GYmr6B8ph6gxe
lQWHtVPySqYOWhF/LhYqwOwTz/isCEOD2GDnW7ZTfTsWoB5EphXM2vBuQH+ZUZlu
VIE93t/nIXSLVgSmXlUn2cQ+zbOGkwUUDOchyROGKBUNW9+DdmLElrAtFNCh74Sn
Up6ZtTQYN5iPYOPpDuHwnw/xe8prFURXT7l7KaE7KFtkwXK/qiqGbliHzQy+vABT
s4ISFPh89CfewhnfM4wuoZ+II8maKk+n5VjgkLoRHFlg1GHDbel2BjI0uC84pbdM
ZAQp7YJCJl7DEzfXnQi67F7X8+mYc6WZHd1yjYuMssRV0Hc0WZMd6QSDGFvYEx6D
V6X4WtWUh3RYiFcNXgEMMI6+OJMUvh4cosFeKfzvOMswaPtnp0MwZfBGf+87+33b
YM+Xztj6X/BDCH0Fshcs1BmR7p22TdC+EmOXjbeoRuz3711ZtwD/dLYrT/HnnTvU
v93LtGG4463n77UuwG6VXevoDnAj4PQBL6LYW3yRSyoDnvc8qTdJhJwsU9xl+vQI
/2NuGENCX5XYfacEKxKM1lc2H1t0zjVPTPAhmajSwMt7uvlhwzaJHW7P/2V41dQ6
YOpjObcbx20CH+MtGhfLLpyiWvqMKBI+NhLVqTL7uaFjpepSoWh+7FX1NlvEEcbV
8LdCqaAv0NyKNRtQgSMZ25e1bySJKl22a+R6WjAPX0VHZAe4gAFbt1LFegc3FzHh
fnXyQ4LujYKTL6oUvxJrfjHBVDWeRdODAJYTmXepKwJjL3nGRmVkOFb7tPHIx26t
jMGmER8FmxW9av73OSf4mtHtRJcsnTGllw66Xvte2LRV7NtMNK3WlwdsUk2oLg+k
rZPdalnTsSMl3A8Zw2tEmV0NyaPW9ugRQU/ZUsqlAugFI/XQ3dAC24D/uLMVppHD
8flTX56iKHxy5pdhKSr8LjHouq5ceBgqHU/Vu0NUoLEdlLp7eHQYu3z2fyGv8RK5
UO+3nQHt1/EAp2ru4VNUCCrFy3mLkXz3K9FxDa79tQUMwwv4xu2TErVD/qya9ry6
3VC9+sa8SxuaWuJjyzJzFoMriSihchl3QAdiJ1BhUdj4oJjZvN35p26NpxnLM9ub
/sv0exQUYHm1a1vYyRtFSOqWHH2AI4wzCRyO2qLDMHoBH3QUZEzZqrXvxXK7OczZ
GDN65DRfPFcEBmMJC+F9wmhNeXzeIkL9qEDgN/86tnbBpxNBIm2fWqI7GL4SK8yT
DgWdI7uVXpYY5P5UxZovYuRCfgunnsv6XPuCuZCRCuSqt3fWmEwQthsjMqK6BtKF
E4QNoPf/btBX/suIt/irWZqlMi7bijUbVkAhDsttidr0tRk5rWOHoqRJUOWmDZ52
X46eKT0tK8hXYMTV36Cs54pMnYXFU6JtmBM93m2AwSpGgc5o2JhyqqLwmfx1cnHN
T/RAc003p79ZM+fdN9M7A+kQFvt7gX8FKdTqbKSAymdGLqcNmgi+W+j83JIZktUp
SgdF1ZZ06XWb/aMXsB8m2mXbxhWeCnaeuL3yXDDWe565+lBWnSUnvHz8WfBpFApn
rypmcWPm0qQNh0mCDCO9Xp/AEwHGB/zdoRsqGm3KB1S/GWc4HV95usHXECQdWssJ
XFQJ6bEHDi5QEzvOS2Np8/NEp9nWqzYjdqwfrpnqco2JyyxKC+ApyvZ/ZzdSMP56
R6LhKMvG8t3/eUuWrYP2RFMRdESsQfZMRmPaqgkuagSp1DFi/0kutU2ACcK9SBLM
/ncN9aThDzavSlaU2RqQzfUXCi3oUm2SNzTtLQlmt2z006wn9J+pL4l/KWAoCfzU
Ru7uQPb6cjzf7pW8UaWv9hibX3LrjYdf1nWH4h+H/aTDPhodZtvTKDR9gGExjPw5
x9KlmIKAYJEOLvUbYDnDNGZ3YJ5rX/LBI1dfNxaZMmy+TN58srlO2IUsUcdsK606
lrv7sWhuez2yLn+CUn3mJMQdO2qAu6eEDSMUxDPr3fkrK9f7Oz1rQeIJhACVIeoB
MfX2FPUuLgTNlQFyv/Huvd3Bg9XKIBVUp2/6ZwouDIEd9zQCEyyDZncFGyttfOtT
c0WVXCUssSr8Ap5/5Sopqk2GDcEda+n6AiNjZA/acQSek+timu+l9REMD9QR+kIZ
GdhnBmHikbudaukqUNRofmFrKlrrVIgAjeaLreFisjQakyZjl45NJSkneT5aiYbH
/IvcCu8pDkt+M/JV2WvMaw8e08cG3xbtJwbDrz8w1kYq5JF6JFuSvmpVRO3uKEKY
PqqB4SIrirVzSXvob56C87r6YzTf9im9VrR9huMUnpEXSyqjq7xTqKgb2U5YWAtt
U+9UOBYTeqbCwZXWZqg759H0k1IGZSr7bSOZfLutBj+iaWvfPwtPDpharEIFSeHu
ITPrv0nrRxByzCs1M7k0p1HNgL+/pyN9awfC+0iBsIQHfkfVfOA9Bz+DRBHjTyoP
KGAYjRjsp7hHW9gmGzMeH8HIb0VNT3b3jhvFk3ESkJLQUu5SNlbiS8TzSknk6+Pa
ABhjLgPZQiqH+zGdNhmMv6KJ7/acSQm8UyetGKCPltzJYi1IErPFs7hwplio209m
nfOWFQcy0TPxX+5SB9AsCsCoMvQvg5Vg+Y3X1X15rmZZFjZLr6ISXB82f56CGl9s
F37XbdAAPlXLKTqX164tQ976pq2AoxDCEDr8MPYKtVfJb4K9136Fp8uciYCMbJZ1
C799n7NvRKn79Jw8DK3udFIZiQC6Qj/SRmHLrzpJcVSA5wZK7iUgi6WT+Jp6078u
hnefjebsSJHuMuW7zAKLOHE9Q2THvn/nCZ1pZRCI2M233NdP/sKzHQRBYsRpo+ww
PWLeAyjVZX/hjgO8bOKzrD0oqLKb1uifZiVwC3LzLWNLqJ0KXKzNqVRD2lzhgvRA
Y5ANc31bN4A27oZyEYFKcLAeAF3pNOspBJJhMW1qUS9vyCyt48/+cZCNj7Xut77z
ZKv09xDcPJZ0MK+AOdOXxwmuVMzSpw5giI3K8B6ByAHzHYqIieePnPKCMh8YqWjQ
fwbnu7XjbRYa7c2Xmok8dsoKKras55wm0W6IwQjk7eHgiS524ST0SH8jnZVAkrbk
UT8hbhPwyaMm5wSTpGNxYzjxD7swnHVOKZTR/4R1cDkg0LffOU++w1IT0a0dun4j
8GpMv076+gQritq+BNmDDvEmSfS9enADQeTw3uIi3ZSyL+BmmGDtN4/Qv+exLDj5
+P/5nnePY4iPYDaik3YB09teR8CidAk2C5E6ctgF7YyVEPuASRrAxWvPCVTeDwhF
Mdps80bctXT+5PC98uJcPC339ygk9w/hi7ih/cfbmz8xmt4b4SCeoPc3a9kWINyf
iCv5QHbPdepDscG1TIVvR9NK+1xas4V8umj1cZkYARpq8guuNujBqQMa8Q8hyapi
nsx08eMEayp1w03kxEI+TDQuDiGcTYhSQ+nX08JeZur8TMCahn++QBVZydjqoX2Z
qlaCF/sndVUqaqEFGaDrOfUFYLjgzN3iuuloarb7TlN1FevPGJVTzOYxNfC8sGAu
EYLr+o6ADT1W6wJiYaSmUWB/oKoKJFG/+8MahYUybkF0adey3lvuU0tZ/usj0QtA
RNI8mCUI0xrWus/TrmYEV5/s3CC0jmGHjsjRorEM5kiy0ySK6EduKYyQMDulHzIC
/7B3IVMhhQji/2+SU6nuR2FXrO2AlP2cPwqpqPKKBIwvin36sDH9BM9PryRtqSKl
0OIq/s4XL49JMnNmMSMs887kMKfa3JgGOS2Z754EiQ7Cc3aeUVycoskjgRwWAOPK
y5B6lLkVPiPABCxT0tyOGlNdp5DG8QMYPV8M6XhnaLwkzlPvzmkEyiyDNXL33Ztc
Dh2b2zZNkXtK2dwvBlS/Ye/MaA8VJi9BbJzpwCfCtcRbr1bJ/JuzAZxh+XM9cw4I
nmwohzHfSinoCH2d3ZDXgu8/MMFookWCpKjZfjou9GQ4Ysv+2bmv+DT87xmjwU59
aodNOYjGLLEgS4KDn3zCRYJivTbQdcjFKEoevRw3CUAhXjzaLQREFpPJFvdBhobo
pQFqUpWKdlZHeOYanEADzMKtcMnJOytCya4ufMAY22Cns//3agX0YPu2GfiGoGuk
0YYI/gNGgopzfTcPtsusYGBdQILlR2BEsShH+5x4Q+dyRULVCQfolZbEqzK/KjY6
lD/X7nA8Y6t70LQ5dXtsPZX5CfUPWSwOcWcyk6dxT6C6KsR+3JYgBvgR7gfptYaD
U3AB/EREAU1jA4bS6qW9ZFrGCGnpiveJuBMR2RVcaUFNeusNNbhYITyiTKxtB9sB
42Eevhyi8mWQQqYUMQPE7qPcnl5t2BU6EicFXfQHDbY1UGIor+cSpQmCItl/543R
c2AItzcaIbsOlm8MAEEUyfUnqLvuoNfeDrCP9vDa8IxTt5I+qTEPWQMd8YODXMFa
EEQRUTDEUtFBEYwAyq9xO+4VxbGE++29z1bVR6glFI9gfQtdRj3rh5l+yOhiG0j8
L4hzNIbPMOugSEbsMQ2/3QHSfNDU4b0Vu8OuDNeafaRrspkxJq9O67dBbIn+0ELE
5JkfkKLKtaosn8oAP77NerKbJJZUUtaJfktUTHOnyQNAdN3HknthyedhLsS4o960
Ngvx8v/+JeWlrMGtVVePFHadhHFEKpVPTQe70hS6oGS2QmgoB4QOknqStxo4/QGh
GjE7GbTYzRCjW+uAhRWpLVfe/nDz4rE306xI8EXmM6f2GhtuB/zPHSBw+tGPvs+b
9s92M2wYVYeWEy5gP2c8tOfY1mbSYJFJFd1kGGXsBHqeG6/UINoc5+we4W1aab+1
tvxBG8Q11QmzPvGZ2SQyBfIibix6YF6BQmht5F4CNcsLJ/8pco86XVh8FsgdwKk/
mOK+8dAcaRteHR9PEzKhJR9dYS9VxCQ+0JhsQFVGz0wgEebWjPEYpNXa/osmTICX
2303T1IF85FS9qWwajBAsEGinAIONoDt1PB3jceyK32FW1XpFnBtZeqpXPBglIm6
ug3v9f9mIZQim8fAcCrGTalqHoV0fBHIa2kS2IKZ8yHGuezmdjj244AZvJIcE2Is
xuj1D39gS4y0qsOUaM9N4f11uBS1tFgitk7Z4669VA7HFtRlD3cAOld4aflODQg7
SHvXhE4a7R9CFIiHlIt0KUCz8TgDO5cBClUzbkWp2DBqNkNmiY3I51B52SbQDMAR
3FwzMMNDmGaWGBr8Te82/d0xQY2I38vL1Vzv/bD32JY1pO3q6jx9+tU48BXX9dfq
JyYTvwlvvbuOF2zXR43ZpLUrwFLUHAT3vKRSkmPUKWRqNr1oFtY3J6Pc69cfZw80
2KShpkFez2KBgpBiWj3ze49UBT2QPbhqxFyNX8qihhHoMDPZXZrfo9Eijtdey4pD
31J5B7W/U6lTsDLMRR7FRSjCY7NtqcSbYptINxpN3JiIMM9B08STXrp9Fm0wbmAI
RP08R3c9xZBwRgT5lVZvpNNAvp/0k6Fju5BbuGhVBOb5wGWG+1EsA+RaigjhZNxP
wz/azjGssi2YhVJYzHx+WWHqYTtU3eszdmQ1qzaA5xB6r2ABGtAqFf9yA3iOjtee
iZ6XOZ23KCmJSoJ0RG1wZsNYh6ZMUV77NppW3GwfpTrDd8cHnIFrzBekrqJx4U29
HB5YAgFuED56N+S9RifqCJsen5iZ9RQXslmPiHG/LIWIuQMUgaAKlTC0G9XGcmzL
TAi4gQAaAi3x5VnX1X2qeiT5EZiIGlJ9LsmhlzI2g/ejfajui2JLpbsyxyughnzD
dW/B8++V3irEa3Q5Gb6/NNCaSOX6wJA8mPALP7GRruS9rlL+6LRjWrjU7n0jlI4D
0Qm4aNfSf/9OcTbYJ2A9wHN3RThUCpAN86563yv9cJ9nOyyy2ypdS3uYlNFyqNGy
0AiJ8zikDLDPD+eqqu9DwkCwtq8lG2nF4qVOuFOG/Qo4woeKbtcq2GMj3lfAYZMh
SyDTdX228/oArPEw4VPso3qt+oKQiYHSAhiJNn/grCwk0Z1dZNhWxHUnP/lIcy98
Y1Ba/Dm1sgSOeP4+v2l0abVj4Y7+QvRIHdnHRiR1p74/KNq4EcNI6otKGS/lj1OT
ZYYQ3FRlBjQliB73J4yOGE9cXSTp5c/Qh+q/vbMKEhkBNfxi4jwbCq1iePC/Mg4m
O9pb9y4S96xYaFev47hgjQGnZJs6b8g2XLMv2j0OlhjfUEAVEJSmfi8aoSHAMIOE
P/+lAi5NrzkZS3gS/SgEGM3usvE+6RjU8gu9XzcU+kCcAwdPZAjwIdOV5nako2Oh
Mfo4Ixe/CS0rYw+hwfUyScu3brNyvvxBQnr7hZzveNU8FxCjuTySi/ggblUedpHR
M/s6uqbKJ3FoHO4qb08MvMJTp6TQOGooVVTsb3BiUAn3wWUKYiXmAmc0HV7OkFNs
AsEfJ6cN9Y2tNJLiVW0ypcOYtWchnXNDEcsGwVWoniVKovHClQjvfnV/3x3Vtu2A
65ENegQ92DbeI08IrhbYNfM5AqCS+DvzEW1ksH/ZV3Go7Mp+JgpCAXABwkmfY89H
1fiG7bSfLe2S1kFSS1OmprWyuSDHZuOMleW2E9UtSIxkP8drQKdc8JrSx1Rmwvke
FvlWsDZYgHdp8LYC+/DoiAEBUTa3P5vjp/FyUJFmqXioD7xyWSLCV4PKmwQoELDD
z5c0fVaxO8G6PQp17k3y/2DbzyQuL7k9s0+CQB0uB7uTGb2iLTisHHKBgPAn5XAf
tbxDCDCAK0DAsT8PMOglYEKb7hFqQP2MEz5ykHBncTm4xxSkEqFtvdTOAZMDTIjm
xX2zqDtmToSr9kjW5QsDLbWW/zLAka/bsdi60vZEDsBJt29rSwMg4AOpGNagz5z9
Dm3gr6tF6MgicegBlG/G8eU6qXy5LrGObl1zw9gyCRaoZOwO4p5YFmzCH6kTl7qc
Ew7euPreOgRa/kGRhi3cxNpwbWQxIsGlAraprpE5sXKBLJ/LYrBR8DQ9HkBnSYRq
3nYQuABlQhiQfJK4WHu6gOYpxVQsWx0Il5Wqe/EO96nVOV0s8hxM9jyOnClBal1Q
zpxG0XaGBHg5J+cpz34t52axoFbVX6Gf7tqKJSh0wNSk0y7Ys0qoU8sLdB4Lbzl2
0dIURE1EkucamCeQjq2so3HHFqHoDs3W/UtdHe9RfbAIyrgjM8076Bq9T14gxz3/
/mBJl+WFbCodw0mYwPBz15NIMpe9Bo9xtk4dEXoi1kRMNDNUzQBjVcTfzVFj39xV
F4/1GJbuRxgW7M6qxnQIdrvhy/Guqi+8EYUGtdCo03cjbEiu0LBikI27Eydhg4GA
LbDcmcxF2qk69UrecXvXK7zh3Zm/v3BwVEKziXmgNRG58SnnZ+hxX3iTJORbBvIg
GRPIuTMGVBPM1ILUAUsIoB/mWRIQIrovUfPq8wpUE0vOn7wZGysLl3TjnRlImh1s
lCBiFi8Q2xhFAQ8krsmM4ykLehuzw8r+M5A3UfVURHZrSL1Mq2+lv4Sc2XRoufKe
JeTDrwU6+m+eok9UnXnVAwysu6Roy4PuEmqC91qr1Smts2+s8wURq4qE+h/IscB2
MfVccX8/80YHf2EHQ3hsVTYG15sLKSTysbILgOaAmoPryywWDc1o5FgjJSwkmIkh
lZzcCGROOQs9+BmoRLbCKehHmqRqvEEvsb8SRkdBN3+WrCRc5AsnhlO23tLrwtd1
wFG8p2I6oA+6tPW8Y2KeDuA1dQUTjIkhQdDzPBFV77KmegewSWh3LYcACslam5Qq
8z6Hdy5yP/yQhOP6eNUj1kf1yfPJoLh/vFFOtQwhBvk/fk/x/cl/KDZ0jsOBgIn4
iHTs/zHFry44zB7kJhiEPV5LEU2syYeZJdVneAW1t0AdTKfELVTf05/sBopmiD25
JsG8spj6hkqpc40WirpAXXahVbnyYiEK4BFLOVQc6DSzvs7FAY6p5ZepU35ED5ZI
mV7PRZs4a5IL63Gz0zhkvemte2lIHf0LATeWHRFBMQ/Xg0gA/aOniLi4j6Rn71nm
vEGTnKrV8Cxf2/G4YskrngHC5VGZb9FgqTtKz1kOILEe25KYs2HCBBG316sfxOV5
OKXYfG2w9rOtHxGXIypMzsntpKGSm6nXtCh+iplh6Tyyxot7h9ocPxGmSwHiG05a
VWFtb7cITEiprQfC2kjn8+uEuhoODrYA1luhneyHLV7D8M57YJ0AZph9e2+FEWZn
R+3w9r04trZfT6ycQpvnfKHKAzTMlygopr5cq5RkdWE8Wvykl6vomKTbsZWUhueK
2qtLNI7b4UMwL88gDJbJLi3oA4k0DGolm0uxopqFhaaZ49vn7qquXduaZx2lVYCb
Dolhay4orOw18zcOexWpI2UhnRazfzuPECiZPDX6xXepu+e8MXfWbirdBeDGog2x
gISenyUSOO7qPYeyxP2U2vTJRBpbJMd25BK7DZ5jUmU1chSv2taNJI1Wbfwfcv0N
NEdgxKOMcuID0e5mbQgPpm4ncE8JJAZosishm+tDX+dfUqjyUZw8dZmz6WfWDkzJ
gGEhiBxQ7NCPtKYh3iibv6C6lIZVX1I8sGE/8qtVo31EKxYIaPOcADfeE+hrJ+nr
L/qyaBFc/xHirKRAY/TV64awt6kglJrpZlYyAqK0DkLw69u/3lUnj7wV2ge+ijxS
Nr8v5SvYs4vp1Ga67Uj8x31PdgO8MOwKq0Nr1Pb7iTBoxJNaE8jqPQG/X1I3KqEj
mU+20avbp9EtZ6nGtsI76vn242tT7jcy3GlG/jPWuoiimo5WFT7I9ax2utwBaGNF
KtWHQ8rdnyUpFAo88oUImPB+YwSN8z9RN9KJRHSMzWmMwaNXWiCm0+x4WnRTl7Kd
y3rOmCB0NmPiG8i8Ti7b6Hczsg1GdxgbO8030YBclAFCRqEXfcPBx5AEYSsxn+SX
tyTe/01pV2i1wtizazH1tWn4tBE07m6s0iPlvjYcwYYyn9MjtbTDL+RWgfhItuQW
dJ/SwbfVfNyzSFxAgVOh7u/OtvexN8kKsauNP8fMSkkJ9mRrfoQFyvaS6tP2hS0h
kP3+HypcCpU4+txbB6B0TnJvTrYCPZli9gp2mNXYsE+TKgVJb9sjM7NkfLYTrrxo
g8g9iBf9VWaKlEgDmzvDClGrlTWb0TzWvnpa1R07lsPDpNJdOQe/SajiFV14nCGn
wRYbXWeQ/FUBILb5BT0FhAKujcQuZirU5clkTHlOhG9n9wbqN7RsIX/C1zf5JFLi
ZiV+lwaLkFAawIFTR6L/flG2iaF5HfLnUio81AmHMEI51mAoVBefbfHP0SyMf54n
kwlg6riVR5GyaX+OiNb3R4q44PrloPuvrSN1C2nXjEn1DRSEdquJNlsF49Mfb6XV
pv4q3h1nfyIDyaTAAtCJrcWLgcZ+/GKj0+CMaXiXw6kQzS5f632xBHW1sgvouNf3
aEEWZvXWuHEHqa7w7uMYS0Tg0ej9k3cUW/WsNaXHx3osqSUbdzgbUqlN+kdzOxPk
8JVI4dAosh0+LOQfwARqC2n5E4dQfCWEA7CEul5IwCCQJeuTHf3uz23ulC92C8KP
rAtKMSCpm9WCQ4EN8hex/neDTtIjBXioz9Ev0gyF2gESTqLmvYPawdNV4JQLBQTL
Dkr7RvC+9Rv9X6ZpqPZ6RxCFVapMLSQvyCPnPZjbFvmoxVTOvWr7FHyG1q6f4xLF
8hdPcOJdPDYmyaPc/bxIXbNgZAw0zjV3NVjKAppJUHt/rGYcTXxaXzv7tWVddu4u
3ybgwTpJIthFXrrcAQjF9QGDn/nva9KOMtgEM1jeb2tERmZ9bUdxtNaWVy5cj3xP
eoIbPPkHIQxXKEL9ZH0SBeJNd8zMClWogejuFl5ElQxUlHmhjJErDSo/woZA+Xqr
z2eLVtHY+Xx/rejVJA9Znwp/wyVdKTX5+2GfiKWaTrzka8WEmNkJJl1cd+aq1uzw
lMqQVRpwM6xWacRy23avHVnFGL6kQgwZCXzwsfoM/zSXYC8v1auD+DJwLnZlEEij
PeIr60v3ORtdPTROrL6flb8TnrPMYjOCl+uuAUTfiF2h4DTnTjrqQq5oNVuE6R3f
hKobDNfk19E3L+peYm5P8rVnhk4e3OIt9SOxUwxEqJMkrkZL2e91fMyo0mtViGC+
d1k/5xUclIlIp0m1xpT3v5aH/Qt3yB6nwAEHPQrWbeSdJB+1HOsJE6IMyEfJKMW+
Yn/lKPqKYx+tRkAGCqjS1jXf+hpKyjD2wV3ehEDq6H4bf5jzgsbBVVaRU92W6hKv
tSJfXFAAIAc7xxaiRrqxkDhxkl89wmfztOfVvAD2HKiPJYPCm4VPdSynRvhyHpBw
5+iJh1atVFtT06O58hnuOsnpv38qiQotfGkUHPqvuuzEeKZgiCH0TLq5n/+SIKJZ
eiVGK1/bybl4OlP9CY3S3MjEv6ODUNvxOzwaEuM7SDnq7bEm45H1Q2cEZSNhlmlW
+wSiMj02OXtblg0DMhlsDqD9Ml2jRHTeO1QJYIHi3w7F363hF0EMmOx57p+LYJM/
r7XIfHo3pVRYuMIESxWJkTFm7hPy2uGtqLT9QAcp2AGUtMLC9XP4TkDyWFydP8a4
KOxGV+Xp0TZ3ASNHWvsMM+z3g/nq596Dfdvy1KGSweHI9VTCWJDAu0Pfulpx1lM+
ZppR4iC9qdZW1GWoRgXGv6n5qWj8PODGehS2Q+4fsEu8IG6lGMDmGRie1xJB9WmQ
IbCpeQfC8vGYzAaY/9IMmXTeEMiKuNZ/Y/9Svaco44HGWYnWb01NKDNJPEcQyX2s
Mn3UIeSvb2uM/4dRycj3lR+gTUrwbpXoHUEec+hnIIpNVBEhmrCcQhvF14gPFyk4
jJ3XuIlol806lsdH3QneNxCtIrHdpPH3l3n5rQnHXgA5Sq/0E8ZjaNEyWBqhJVIW
YFsaGr1o/IvhU+NM/YhmmlkfYRqMZm5trkzZRwYIdN+mrnbBLzUuLsnOxc7tT3XM
Sg/GpVXNaEvibufR3+nVhNSg8/RDBy9r4xuhjY4tvH1xzJwZL8uH/pS02rWaBxss
UZUkxu8CYaM1vWGeDaBeW/zsfoWDxTmG4yJ9n8fegQJKVxc+gRkOIm2XDVWSNzSa
4pcMW0rnRTlOpKq/4Y7JBlaW1JOUQbVR6Xpi/O/nLc549lW4kkHmeGIBJ9RTOh5G
+kcP/0zvfX3Y0RiZzmKRpPuaZEXXZCMEISHNeaF6aJ/9NmRkeTflLrdszsjD2Smr
jT39OaoVBmkg+WJgv862m2KCQ9Rluj82ZwBP464PG8hl2cPaWjIhHzIfORzzHddH
XdxCcLSgxCwv2dZeUWHXK+REYXSEsc4GeMv2tC0AI2DsGlYNSouhg1GQHk3Nm4xy
ld1hMambnLm2dkhGTqoKmL03vsgVdRBPN02F1DuGm+2Lt8ok3vGxEW8wp+FAlqit
Hdul5k4JF2+dpfoJREhTrn+VxyHBs1ABY75LEad/raVVpmQTs2un3lNVTbrM2KQn
/EK0SsGJQ4/54awnBvqOnFpSOpy+YmwAfRmNXK8/rWLX4LKX2vs00Yf9kLm1Hkaq
T6kNkAr0If4KEYl3f5GFG2t7DfotpvNwFwG2CvnwVx9iAY4Aws4DuNn/z45HiMIc
4aeAvnkT5oQnkX0726ObowNljbuQgIjhDSDn0Wfmm1s+7HZwVid7PEUMVLb6nKa2
/XpwiwulYsrvwlPiAaMGmHaK5M4/XhF2N3ShS5xhYuVgqXA/n9GiJL+F5P/nN7A9
IvbgI5Baeii4Bw2zsDldUjpUa33ULka/Tu/O29qAmW17hHF1e4BOGEbLgtSFVADw
yiDxh7w2NwGWCcJznt/CDEZpN8sjcS5ZWDDA/vUpj4w+/DYf9Na1wnrJZszLU1+9
C5ICNgDji+QWIJ3rDZlIuPlWT9THa9LDGDiAiWxYM/WDwQok86uLqKSyrXD2FT0Y
eV4me7JkMct6lrRrKcMQr6SjYAtjcDSlUNkBciigl0+Ungfp+6gJL8zde0Pu+FzO
IPIXqlbDNU9HneENabVIeNwZVpoKwYWWIU5s0qWuOk/iDvgLISChuV+yq4zoI9up
r/Lpg6P7yb7eHkGzWQ3NtGQuNUJxHLaLGZk00PqzOCgWXEnpO97TQC1/Ex/NTIzn
nbpP5iBtHzsg57T98A8IccMQGoqKgLBkQHJcFLIGV/vk+sHc9rKnjuiU9hvl0qdQ
yAu2PxVRreT8rNLH3ZmlgaqT7/pLGKNaHKZA3yip1OBAYbz2wTKbWRWqSB8v0t5H
4sE3R0o2QM4mPfjAmkDCZLiaUOTe4WYIpCsDF4uNIWEdUXnjIH5WFcNsOyBSz1im
//QR7P333DEc4OrB0rEW62fweU3XUibfo+KWZIK1q6EzPcQe3N4N81ouGV1nEafY
wkdVMcYtw4WO5e6VlAKEb4yfNhPJdZs0WODEI7/FYjb2V43o1pH8a36CqFQL+Hfv
OvX/RnlKnzDF0GcRE5oeOzWGM27/2zQ8s6D9AxYv89HGEtYOm1nr6lEPVO6xmW+i
0Q48WcFSQK+4djoQ1RRf+0PbwY4Dk3d41pwJyA520pl2MT0YKwemEWkWGChnfIou
on9KM2jv8Ixpi7pHAa/22o6rJ+ARXNjr/aT2UB1u7h4ctD9GgFFRxV/9n8E0xtI/
UPVZ0BZuEOClThpBN1J5a9hqD12eA5GJloqW/0Aze6QQ5S4vE+29LnXngciv7tmv
k/6DwigmljjFDF7UeY+B26MrfOUyYT19zsaSwX8WpLk/wEqnoMPfQ2uBTqtHtpTo
L8GVXmqS9kjzJHmyPVUHXCTplsyGukGaQS0Gz37rPRh00TkfzjDa8he3c8JORdM9
igb2nB2QNCowH9fs+/pbJ+mAJfhURu5T0EdYhdQlzNjglXIA5Ayb4eW4FO1Gy7LP
Sasm3lpGARfDDU1USna3Hf3OSfG35u8yyAoOcln2kIftgXlNjUrq1zIPGUe7mrQv
8SMbZTHtSeaNB6bW9G4r080est4HEiySibDm3psRIkHhsZRwd37pGmf3QrkiLNvc
IwhxZL9375iz2aTzZK+xOw/SftUVLmehd2/aoC/Obk6kdYjS8VbOTr+y4jxVkCBP
fQ3hbjhcMLiCSJCX6LdJVhBheyL3rXkTHQhekXMTKZpeH95/m8Unmbh3KybxD6o/
Y+/YtPKR1KXYQdOFINHnC+PQmn67633c0X0loosL0HEw0KbFTGbpsWKlpE6Yq89L
eubMOGUbzTe6ZUWAAsfWFYFdb+vWXDlTME6FI6RO06senMt3Rp18pK8ofUmfqmhG
FG+QehDXY3oERBi2sOPMZBbyATJDZFMI/5BOt2Vi0Nh+iyL9pYkmOVI66wBFZN27
hSb3myjWsk0Ilyt3ThkGJ3SyIPd8X4m3bCYqo4G2i9EjG1nommpHhAa35yxW+OmX
8AC9wP5lT5chomLBwLP/I9t6kZIeUlZcKWL6bg354iC3jvtoU/Dj2SCBSOKKYe6p
YwA89K4H9O5D6eXliMkkEwZ98D3G8EA5gQ0j9yKR6uhWNrXDjQ+amcheLhkSa8Bs
Ube6jifwafgUTKXX3Lu5j6LmfdptHjpB7FYij9DbXPonrwm9f7/aTk/9ZsHq4jJ9
BHffoCcoWKYwjLomB6CGWB+tutsWvhSTW1RhhgJ1jrXLuCYA/ClbpzEm5iVY0gIM
IyVkMaflsc1QIksfq0DOwIhgV0I6Jv6ftekextet4C08Yov65v0zaaW5J7xAKj7T
3fEgwVvTgmkaSqP7VYn99D9fTnKaePHPP95pbn4LUj/v8mgtnvUXpuUODbxSNqeW
R7CUR6jF/ngvdNP1SRyx1tYf37XlyRl0fj0CuR6DK5Gx/5u36tIK26PYDZTP69Uh
EjoFDJ6G6volbMaTHpsZ3YSYtO0Z0yGKyNg/w+Aso92SpgVhy2kT0agEUW6kdmfP
3P34b2PnyKjgTXZUVzSs4/+4tCUUiDCu1ehqLfm86cvUT5KjPs9JHbDQGoTEYvVC
GMoaoa3zt/nYAk87YRrfRVC/r+2NIHFrjldkFXTGlnIXUTCHGP15R1DqVVPE8blj
Hg1rnNW5r7Dz/XSzBdIglcJxx3EOTmYlwryElUzBj+jCkOlT+xJROzbmOY8YZfby
AHHEavoo0saDdwYCfvO076f+AW3+Co46steBrunPDzWjxnRRgSsabOiq1CYXmR8+
bv0ArOwl7Dyg4gKJY79ZdvsVH8+I0Ophrhl5gh1lE+/rL8N1kfEplthdcA5Uo/z8
BYxwc/LjoBtfyN0rSuFwQfQeYTVOg9vku8t3msCbtk6/d9e2d+ikdFmBxGHxO3Dv
aYvM9jWJ2KAGkKdyZyaKnQGTdTKAmuMZ0J99DFoFCe48ILLurjItRiI1V5B8TBhQ
XQNjUXv2yLr5IqiIFwzLr/jm0Md7p0CeGGw2DA2MGUpQlYSIhJ5P+NsvyklA8A6v
XAAxgHg0LK5FLhrHQU6SDVhaKEr1vw9kRgGH8OZNyQNfyTJRGz8SwfURBikQVivC
03NbUNf5RfXPwQ78jbxJEFfOyXqCkqkM4ktJbpEmxYX51lIbl7Nr3OV47kXmq9lR
Q7E1lmSNguQNu5VK9WKB39GL3Wgy0JB4LyMSYaK5kvDDS/XxEOF2Aqmlpr31vb0F
IXxtq0wW8wOifxrbkjLlTfm6pw5lGfOIykoOpKSUCNJhOzz0S954AFOBjaD3KDrP
wfjWbBUNIaSKGNrPbaqgwB81jMSVsYiCz9hIxucEmBNh9hDfEtSBxrMuTpiuW0Ux
u/5mlcDhsBXaOqpXIN3wYj+P7VjUDD2JHKl7qHAQOP6M+nrBA/oCqFVWo3bpbZiX
tGMf/d5v+Y62YXgKXyyIOTW3N75Arwucl6ZrqreK6Au4wK7f/gYq2pXuWqcY2Q6f
ilDxT4LyLA0dF5v9KEJCdMC/Gdpb2Mjqq/u+M8de26J+83KOOcf9QKClVWQ92rh9
QIHDaj6b71sSVb2QgT0fKbZlX8cWa4kIFtzChyD39ijL4GotVvEVcTzNGdu2WBT3
zdZDVG+598dR2VWoEpf06r71k2vi0NsshnEKuMX0wAAHMNqJNuZtMaunXMNUayk7
GcCasFe479S/fKs8QLREFij3BVfYaN038nry0wcnYrYYUjHH+7wABywdKu2HDS+s
aHHvFrwUZtqvz7KIVHSZSy+cr65poXmcoRvlioiYkqi9naaukyDOOqCQtIEA2wNK
qFzXWD+Ao1/TgzAi8UEUOaJmLlmbvFgJhgEq2N87FVbLHRznM2mwc70HfBsnn9bi
CRrdgxtJcHCdAl45HnuKSgOQO2e+J6w5NjXOpR+zMrip5wWGx5/oWxUOJ9MwK9wk
Fx6gAKJ8H4bQZNNmS0kdo+ubny1up0pryiQK5d48RS6d1Ag6caWnE0qxWRnyuKdf
V5h7SpzAcY7Nu0ZRr88Q/fzRdL3ejMesLNKeA1acHYLG1ApiKOqv6h3uAkoaNiOa
Z+FyhzJOA6lxwwWaGIOv6idSDuXaIAZ5nroU+yfsxaAmSQI9rRNjC3JV6SlbeHLk
Z/ePghlTemYNOHqMOPdF9SK05YQf8HLRMPIxoMa+zbDCJVfelwqcosE2413sUcCi
NpTGE3rSxTgZuPMdGUxD1Y6OjFcqgCP10KoSnT1lu8Ch9o+p6OVFVx8H0kI9201b
hI3KNrP8Yehqjhwlxz+HXvSEX8UxJ0Ug+hmuaie9m9mbw03G8AEd2TNG+5THlkH+
NsYtl+SZxvgt3UZgYHyL8HTQoSjCsupMjipRRcLwc5x/rL+SV44ybRmqGszCnC7M
pQnWlI3b3h7aO/mjXdp00Zg3JsxvFqRtXflIS5m9V4UcsvxnFXZIQhEWpy82WH47
QnyBdSpDSoynmw/6djsFlHnjK4pu88mEFfdj14dP55Z3cubEJxEu2RWTk7DmAF5F
Rjx1mgSt+s7sC8AVyOzbdCLeiQiQ3zTnAu82NY9kOKS8sNCEVtvpqZLdTI3msskL
B97JlVSy/+Zeq1vjrMXn9djIecRLB+jYfwR67ti4R/0V/y830v94OVzt3ELJcWGf
KM/keImYlDxM0fH7pe5YJnJhTNOPGLH7bdZF1B7sRvyLizUyNNxeKYYzX8CtubsA
cl2qTqVkpZJg/9uoH/t1Azk1SK2NwNzqVf4cs7je0BaSKVkrgzdEIxtbfCHGDnaP
2frQxfcESdxjQ8XAGErX9mFC9+yCzfVr01pek7ayeHNEYsVjBUciCLUuYUWw2kOD
Evwgl2wpf0md2a6yThmbZqBi2EdA4VuQTb63cIBGNlm84BShsdMj8opub9iA+3Yh
9jGMQpgG8wERzJURhCnMXhvc5ql24gFqPmbr5sYeGrhoBqus6RTaCe/xtHR1yahE
GteHt9+Apoz26tsz1nlErOKPDP6sqhcyHk12GFuAkHslNMtNRRlWUeoWcvgYpLfQ
BjEvrEGNszWzQfIU88NfwTW6iHj+ajtlOTV2xfWQ/fDEn12OaZShdaPUo5gg9819
ogshJt6QOzQjnO6clH6cEi9BuOk9lNBI6LcdxazSXCX0+ClJ3RO6Nwr1Dn/5F+Zw
JtHelkVmkpfh3pgt4KaYPJT8Ev6Mw7LpW9nJhC/4i1Am60ssOD/LGojy+y67DYdA
/oz8Ic5VSpKF8QL5RfkM1xub8VaU9vm/NIVnBStrLH/0asJen7oHYFbynqOdNI2/
h6Bg6Z3fon9KS8cHIQD+QmYVWbLpZyZydwQiO9VeelvGS29KVqVTrcmOBfq9l+3z
M1ZilwyO+3R6DE7VK7FLkklc3DaKAmzLe8qOnFcjLWrH87m3meZ3dipxz+XGvRCo
FyZR85SzXVKuf7Sm16ZGBWKfUlBGGDhOuibkEvJ01/sgJ5SNueQ4PpSbF6HSCYuH
lMRFUqH3w56e2NM2hqvu8rSjkE0EE8T3CaaA4nW0P4ef4eHdxYHudgUlC8/2sAHw
S37+D7tDG4omG1l6jbiCcglY6q2T+JrP6HZELTN+s76nplvlQZz2xFGgb1wZXqZn
M+maluQ6wVgc1sq5FZZ9kucLDvW2mDv5aTeyUTL3mOTyCTZPxBHx4aRLP63LDfgG
dBkXIkd5vkh3DhTCeDd9qVXZWGXtO/QhHuhNFm1/C6N6FnW/JI1MdKR7gpoYr/yW
JXDXjcafKlfzeM1jBHEvsgZZUf6c+41dNicuLzQ72PVaFtHXP/N1Zjg71OcTuLS1
ICEQ9NA+WgwkkGNxgfr1DqEsMaZ8Dsl72H0zbsgDdaTs9SEAOu53x5tDcW4EF4IX
AhkbPV1hCXIdYSxtN4+AcdVSKT+d67GFJ/J15Y7gZAT0aYdN2RL+TMwUfr++PiBv
ieG9CgDc+Y9VWdDIaaBZc37B1lHCv35hzgKV26StbHahuWGpB/CcqadWgusNkljJ
3MCGcePbnApdqq9x8dSFKPldH8ohHPx3/BXm/R4U1LWYa+0TvLPMxxdR8hq2Lixw
TuIzDynZ4ADj/R/tvQGycJA1xkjVvPCqVYY1DWcpR3Fr+zG63xhqX7V62GU8J4jl
b29XExKjHBricLj4RwcYrAGcVrxHxlIxPmKzVMHWzY2PbKrBmhImMt+BACcfQFuq
R8Htm6Gxw1hhk1UzguTSqeG3dnkZG93vrUjFmU0HzXdO6jHNuVR+cpTMW3ebf8OX
1uJUpG6J1Eri7HFEsqNMiR9KMFGRIk5vKKh1HZ9/YWNd5YL/vs8rUNQkkwDrdhbP
78tiYCMVgs8QBT3d8koFtgaZpjIvmd4LCkSj7tDKqhiQUdNSmo0Yn45lTvJs4tpS
HQy2cJwcLsoTiXUYIElED8Qa5Qk1YgbkqaXU3/QQTC8KfVVVa59Tk40v0ALsufv1
VnpB5RdSMq6fRCoWP6oMlfjK/s5qfSmQLjLoGjIzMMdN93tewrkIh4ZbXlr5Hx7u
KwYq+V0T/k0Eu51Us9zCvS8c/UMg+msMzvr7bbrPgYREyl06gXh5cTeiqPfFqqmN
DC30q3plGd0RBgS9pJpa8YSe5ySR2FmuW22Q0qdJWTft/yTvtwzq6kA4eR/Mmvit
rsqPkxdsqK1XlxfwDfRRuvB0W8hLmjNr1V57IEq+zp+ATbO4L8aKsQT2+C8mfd+U
LbpBF+XQespl5hdwoE1msrGNiJ2R8eyYzZ9g1j7jyNIsviTGLrJUfIN7HxnDSvYe
gCmekAykPGo2yyY8mnlML0jbpuKUn0INl+vCTQsW4Ax05Rwiim9ZVD6C5KiimPzX
znfVbNi/Jhk6fRIEt0mpw9hJ7wAIO/gaRLJhQLapAm9z9X/6i7CGVodqOaczJ+cA
ISrS1LovJ1ROf7Y6EltJE2xLJj4KFWGPcTwRgoMwp95JUq4siW8lseun+QfSLr0K
RtqktyxPaLsY0b7SDJxJhB8vJQvtBxp9h/P+KCEDfgIjjrpQ93js9Jd0VFqa9CSp
crwJcT5alUDpSmHS0J5f5PlLe1JU5fbbP0YEpYSVO03mHGsUz1WMkli1B7BfFYLD
zsOT9VyN1DvDjlCQlbKKiqknOogUMzkSAsVHr9ABdRSU5wKi/pGh/3uD8/XinA1L
/rdDw1fFOJtzQo3JhkmKVyuW0fQoaBx/gjMCX9Ew6Zi1OfeO53Lr4BaoVGMkIjCT
K2eSxgpEOC/X6P2XH9SIUzXmu7LzvIOTN6oYWIY6VsyaHuJy6FtVg6cpQyKsxMaS
r2APTEVRV6IWrrNbOR5BOczZgsOjvNx15/9VQCrqdXUVN0kROrEr5acE4rj7kLLy
tL1enuuxiMn0Xxiv9pvIhHAnhVGOePHb9cp3YJwdCBt7+loS83MBAgxBtIQd+gu9
3OhnNyOCwucKQqWGV7fIolZbkAeUW/BTsrD5t57VcdCzqC9r6U8xZy4JuGn5Kavq
ScXeV/4jf+40RfuZj37hRRJFAGd2Oo0TDnTmsOMZtObJHazH2vFYozYBRjKRswDX
ls87hkyPmO6as6jg4o79Gh5nUQ0Pus2YTgpfViMxBSCW5Na8Xpj0nyzj0dOuV5Ui
KY7cSwYlip0KVadvMeFucL6jfAvsSZNnJOqJO1nZ6/k4L3I3HsmNU+ycSOt50l9c
AMDzgogiMihVtjjYtXP85Edkgo1rnMt8LT2+qVtUe+uJRXehFXls/EK5JSFcw/IT
6gl1cCTFPrS6v29U5spL0wG0SikxSEjihJy8EYPoIwbqIjKHHmnLzN6ASiSh7AxT
odBTogyhkSOKyZP/1w710ARnahJEkuaVG4X0Oj66d2q6PFa3/dD9PjqUDpQOmYQG
7V3MYjyYmaPViwP2IBLAfN6ivKmQp4KMOgqT96EQ9aOr/6Tg4LE0bwkDU1qXseu6
64iEcx5wgH8oW+X2RQzH1tG48P8pQL+VgeF3LV8xJmK/ZVkWInqFPT4Q7FKewwNX
YFYKfiGDBojdmyfQN/WyEzv5DmQCgH0qMux4WM/fAP7tUHzSN5xLUz3jKxdUcuEY
6paJ2SBFFXQNt4cdms6P2m8t0fAy/IXdhwoQZOUBfTSvJ0pQIfy5oQ/iOSPAxR95
eZj+/X3qehFpZ1kuCmp1MeLrtM3i9D7LwxaTgWzWMXG9yrB2fOTKgHIVaUZEVrtB
thpHXvyilh84WQDbEYkfbpPaRKybXgSmfSYGzy6IkysPggwrnEaWUXJMo/SIqRhU
o8mzVrVd5XoqsFkETXrpikvrUHYTVVXCUTm57d71PXFt47BFL4Hju66qQVMrD0NF
Gm6OsWfANMy/YEcsbb6p0ZankaJOA4jEjdGIpmdKy0vj7RRWyY9aOW/EV/h12K5E
BS1fBbhBK2rpRLIJ9dVUt52mzsmk/nJz8hi64BZOOvtTK9ygqyT7IT9mMUgVj1Pq
PPvOGBbLxmZrVYXUnMFJubKP2ilJrP3ULwoexRcPokDAndOXw265cpEm9dTyjKgZ
5+0Lsg/Dc6/f0kt1Lw/oICNUBiab1eyTZR+JdwvJXSY9QTJiV51Ci9JQt+NuEa8H
9ATlkozm9HcJOYIqVAmmtVEVL3BgDxUczZ+4Rqm998NlPq0ceyoO6sMqA/iVAANX
gg+lBWMs5HVsTrfkM4/H24R+z/1kQs+zMTdxFkiEQfHliS8++tTiLhZap7wbHwav
x//ElYETbsqgAAA0Kxlh4EMjss2olO47mlwIH4R6xw0jX1sqbrpDI/wdj9cNvQib
k+/UcP/XbXxTTDYsqpEc8fhK91yPciGefVDfuCJgZTe6OZMUoXjmjs6jU2B7GukD
KhCXUXg/LuS6XNmz4S+Fr7feVVvg2cXCg71gdciQK13VmWFKBRjQL5d6sV0TI3tS
rX8yyqdvulzpQboh5pf+IFZ1TZTFob1VfKXiFhWfRL+jx9HcjSGzN9yWwpwMxirz
s7sYaMtZBjL94s1SEj4maEpsut1vKMQEvPOMPHOgQ54pUGldCHa8pzVQcKNGXu8g
X5ay/ftxm2+3SJc/IDygX12nE85BN0LcOT2LakPgrsW6Qj95YziW8NansHN0FihC
NdVVr/ce+/tca8RqfDFKX1eDQtM16sIZ+nJJm/1spb5f84EqhWWNiPoe2B1mYmXc
BV6rFFKTAFxALrAqaA3lZImNuwVZUWi+y+DdRICbx/Sjn8DfGloehvBEiKir6ShM
USsQV/Eqr9OvoFZx+qX55wqPbT47AJxeMvtWyk4PmRZ379QPFFSxns6ENnf4iQER
msOXkxc301tgnAAHadRY4WoXYRjpuUjsW/YZ6SwnvBq4TIYvwLjW4MN0FPDFc1NZ
cDQik+tqek0Ov+P2Cdyhkv2W3XCEs/aGAmC7f6yGaYMATwIHOPMcXT0lQ9K4gkdK
biNXFoWl960MNlrQ34NAFURrirJfU1NVwf94jlS1Yh3CYDiQE0k5Kt1Tn4NE52ZG
wp3VpSCd/fHnJCSw3oBWsrcanobjLGCVhIceNT40vn3BSJROU0rLvE3np/iwPBft
yiZ7hGVIuczTmLqmRouvjS25OG2Pykc7SsvuW4qv6SLfwcJ3GVC4Ml2Mba1QIsjH
sHYL2TW/a/sCcBJW1RHwxtbx46ywuZ47/NqpQy3ZPceFy5vpnDWn5LuZnvOtNz52
HglL885hSgvONK6wQIfXPO1pKzaidWVAeg0OhS4ozfEqDeoJdGrCSD/r4mBj/Npx
TJBeUIfmQnL3rqcG679V2EgefMJ88n6qYCV385BuuJG5SKw+zHcrxoMDw2EOjcQR
O/fob23wSTrvWykYVAkyzI28LtETj79toUx2XAEV6e2Qi3m5DKOr4wjE5cKJtY9l
JlxvyEDaDF5+zmLMy6doz+wrkxVJuMZWYK0iqIFFg4BV94mGG69fkvbcu0mMvmxR
dqv62EKs5HUSRL3mAOZTejzU3llBZYarDInUUjhYRpDR0GtIdA87ZdGGJMneCYVp
ieRLaQ6TaNCt9Yl7TUhbp8aM21s/pH9NWhDlxdkxSvUJu6APX7nTMJKLuIkCfnKl
NLdStsmrihQdIphVSXbIElOs3HehCK1bb9TQd5ivhTr+IJGrjbXx4X1iIS4Xis88
s6rpgoxjo+qYHLjLqpxoxadJfAf0KySuccD28h54zhM5WUza18jh+ozFdaEZ+SpK
CWtNWaBb5gzjUzLmWhH6V5q+1y7cLs41n3Vc92vIETxhf4gWd+RD9o6AQcv6NtQO
VmOSgzBYwPBHMko9AbOx+XRrCnwNhfp2fE0+VnJmTSS8UEHNiraKggmjUDPEeCrb
MaenLAclw0jVdrUO8CcghQRHLsZ7P29w6Q+TR7Qtz38nb36VWvEag7/r1G2fTmXl
JWvxkIO5pVxLy3V/8wf0X9L2rxA00kdrpKTKFwa0g+HuJC3m0BPMqfhZpN3SJ0ne
VasviTzZ0E92919jbwHDYrDEyo2AOv6Y6UIh/EnPwWhgI1zeRulF0Q/XASrfpabl
VqSS/gwOLWEWYVnafLbYSm4b+rRlmbtTK2AUSinIPlPN0kG14ygDyGLuZ7J0JUO8
b5RQL38FcZGl81S2ac/nbRn+QZc70p79j9tjenqvdJRt6zZ+2kgCjv8XyA6SHuE3
qE2Cha3QU0+itnq098tDmG8m7lW4xlUimjqXzqeaTAaPgnUMK8TLAMss6qNc+/MJ
BD5Rh1elf0fhqLf6MGHv0d0yk/x9lwjTz19MXy74LxQ4M6vOEMTk6huGu4gPnJnp
7pTmSoaF0Zt0B2c2ivY1xu2JjX9e/eOyZRwHs906x9X1aNpm1loOXur2XsiQLJap
APrejxlQeNzwQm3V+DLvHamoS/5xW+uXZE3RJ1ZytpbblYkQV9RqO+H0YsshtbfZ
HkcQY8Rsr9A6wa6rteZ8THtBkOASDrXo581PmXNd6xPlXPmZNw62fluKm2pQ4Bof
2k2eW0Oyn0VqVBm1bDknJQ9T7FqJxLXSXx0DmZU9mzVtbhrgtQpQRjp5gUqTAqZO
o3hkd7CcyRJjl2V/SFIwa5dh/xSckIFSaTM9DvMGKdutd+8+MRXv5yaosUQwRYUz
O+7yCcE1DITfs0f+n+eXGCjEEEMy4oCQrVyj5JqhagKr/jwyQ8Xkg3y9QH7sGkz2
mpC1TvrgKXY4BiSwwbY3rucnt3wvIokl+7raGDMZW79wTjMq8JwZgv3H0IZALJAH
CNXKDTbnPP7VY1IMBgF00zVoaMp9zsyjExQtHPAq6jldoYgQVQy/246oENVZ/3Dl
j8H0P/CiENoZ6o53owg680osJvJR+rESWHEdg3uAgfbbNjxFP9WfZjxXccCedq+T
Coqr+q4FtxtZ4ghV6UjWiI3IhUnQ4K82aTpHkAPmT4RSo7+PUE+r1kbiUCM5ub2j
3OH/k15AuhdMLxqQvN/4dGJUShig4RG2Q72fQnsBVoqveVnfhoUxK36vSGjwAgFE
ID63tEPDppkBzdRuvK4O0JotoXt/2uItA/8EdVJs5ZJCDSbupG5xkE1PCp620SjG
zJb397bCIculzlRCxqWwC4hU1gTRajKpbAEVSdxmw5lyx1+lX3FeBBywnDe/sFQE
KTnhblDIIhrStFUIECg4i6hrQcIoM9ZvgI76tnPw1QBgzJgbqyLS72J9GXRfBHq6
+kyCpsLSz2fTDIbDHeiLWdwbRNqwFfOT4toQLFJtid9HDcnzc0cXlGkY/sZYTEF0
uNOoxlQ5pgPDf8OjYEHuFRRlrmh7rUaCU4I+UCcvVpsWkMZV09CuK+XvJn4xgLUA
KdRNVVERK9zPMzMMXwTliniZoQJaw2TML14l3MNy8JPa4qvcwxlRqTHxBIlb2+tE
ZsPpTQwdd5ucOe30E5OsBIWBo2YmexRkEYBDTW8vBK8/Rm+ED1Fjinc5Cl7w0l7+
oOhjKjGCepJ5bLy4cjx4MjASUIYplqvaxK0s6KlUAwJ7VT9WlmHM1nwptpJeC0p2
xMo/y1qhSygalzXV0rfY5ht9xOkYQcVoyX9xSHi5TtpLGHpLOJX1ZLADKYKjKae3
23SvlxbfR97rD5MDR1v/ePEJ2TjVZS8hWg554RF9+xoqyF6GpUdEFjBq8Olfuhav
HZcwSbHnB8FkJvQ00wwcl86A1S16QmpGx8RiObYHKMDsvVoZCxcBJca5d30yZabJ
PkiBBFrhNzT1jvPRgFJiDTw0HQ2apQe1vFtWa/zOmCmNnxiBTNBxR4Rx5/+Y2OXB
B5Z31SKTlMqNpbFUE8kjo3++mZnQkSTVxTRQ2TOMEDwgEi0wcrJeaFbDkGVl8Ej8
W+ur/2SKJuRqadN48etAbsDTXbZqaQKI+P+rWVA7kRpR64wT13B1zVXXcssBw+Np
LzT+YYlPKZL1gUoJmYfQ6k8XDvciOHrZ8Sd0Ve2ewEvwFWS4B1RQe7uZF6EOFAu4
sC8AEwh+GbUZhSU3NlHDowE3ggpMUgWvQxYlHsoktd8GgOXi8hW39/0nSM0BNg/+
SVBNhvMsDcwOiQtc1nCIBEKIorHFl7nUdyDG6TipBqv0v7N3j4ZnzlHim6M5uJgD
klrCp4DoTwDpICDoqY7/aBwCro4/wbtTvEG5eRHCJd1DO+o3CMtSizhZ0Hjo0VBR
adIV1NxKtrQhRlXRr0jJo6nviAg5r6Sgsxj1l+AWq4KZs1E1F31rPKrErdmMLQVy
rOjxbobbkd+E85zgMjjGlIJMeBRMENgUZbJ6dolt8DkSV3HnZneJD6lGqML4+9er
lMUeearfbxcMST3VxOgZUbl7HIfrTbEAFXVxyEGBs+uTpLnAcccq2fj7S2q40D0E
4MqwDxL0ugYLOaW8N2Xp1Oe4zhXJAz6d/TXehuP8VbKFTCzEmlOCt1yGy9vx+GXB
kxW+OKqCON1pGUS16Q/sYAcOGCLZFeD+/hXMF9mTpeIZfIcjTRPoRvhqPCnzy2Hp
NnCn9DsxXpY3OpjbF4yTHHJK9uW7Q/pIccnWq/QcX1hICyFLLiMVZqy1W2xscUXn
28Gw6PZpDj2xl4K4tnDBjiA+kgqSdzaycKklXnTZ4mS2BW/8tNKLUCJZi6LkchwT
x6SL741WM+FtJJgdbRFECbxAWHaqadYvyqfzsU9nvKdx0uP8waImxZ0NIYHrbAgI
44TdU/vl8L4y0vt6RkcmeoIOCrvp6qZbX6hVXGUdLWM3s3jxbsePunGSAqlVSmMi
+z/D71CCK7lrasj2OB9Nq+KF12rK50j5rdM/KQTwYxtY7qgCElg2va0bIS/tBMmJ
F1mBuV1sA3s7y0I8uSK6EbvLwRwSb6vmBqlYaX+6owK8qciIRWsfykhYc+HbTnDP
yiaOGypXJsdgRUopM+SEQEBi/8m658vJ8kBfQI0mFJS8417KTMW3lzsCwrS+wv0N
54zuTt+eaUbtwwuf3cGsSd7YzEds5gup21AADxdSSbwNRrzBw9PBQfLZMjVruGtm
nVTZ8w+WuZ76eQ3Lfhz+oAGby9ZIR0bDPwNsyDv12518mCx82Yo8y51szGGQkBxv
w6W42sZyRsfZEKOjHFX7+tjoibOGSGclzO1Z9PRXhTHftnabVTiicJFmJyAnkdcb
BVX2Mq4FslGy0ot3uSTv/Hb1Lv/IAw1lcaMP+Z+PHpWO66VPevRcMBbJdB4/rjoh
yiRobj6ewn0lBOR6fygThKJN2FJQYyDUL2m+/0g5h0wAonfRTWyiLSe7RWFXUnrQ
0gt/MCus8TQ4JSrAyoLub7+og3e3D+o0k54Xc5wz2Jlq1i+Joni1+bK2Kw3sBoS6
N5UP7bnpTdxDd49Wnfkx6JFrCFKYiPvmuakR2ugIKYUsaLs05uxa1oEwXNeHD5xG
/3OPEpYeZgBRbUzSsm6UepLd+sE0sLOH7PP9AaZ3G4RDFiuIL5cqyI+Kmstrhwz4
P5rRbjbV7x1lQ/eKwd1FcMIHO3VrMkb3byY6JS9cwNmsYpkC2f8lkpzedp9q2xU1
DXxV6zY0XsDsw8VNUL5hia+xxHFxUqGzyIPNcSFc5i9RSNs40kaq1Un7YHpSD55w
ByWuhluJhhBKZvEhbyLgqZjhM7Y7FmQkMgpe/BQwjJpfbI8vtuVJpXfUwxZjd0wt
slv/vrP4CE2Mbyt9rcPbykDHqMCdheqI7NKUMi6PmD9dJV0xmnIsbZTc4ZInc/m0
vV8libcKuoEgB8RzM6zWOlNHursxEbYLclkAYyaJJDOfp6nydi3Nur1JVaPLTFlz
iMghG729017262ZCRHfepxtvfHEctbTv4DWfeZKSzazcljAdPYjRjT48y8RudTXB
biKlBmqjaMgqADY0p36eCMntGfUwbxu6Ql0hwxWnm1855SKxs8NPhqK2TfBwjsWd
ep5tiB0xaWUGbjpI+tNmVx1nU+P0UW8yNdJuy3cZL525+RcdcJx0XjX4AbdIDHNf
7rzfMA+eFKlPfipzv3TX+irJXtiNtSiHWpueYOHJ/KhU8hH5jtgvkAOe+pEz2bEa
+eq3EW5t8FMkZ4a58TCkoU0P3quRSHGKUOqJ0F8jn2LAK2/5qlxN8YO2tPDkQlm+
JDVVDcqNnUsfH5t2laigeafmXZ/0Mika2qrP/nDbh9222Pc4KbKTlU5InqxiOYHg
6xoNPKw9ZNMP+E05c5i6QEYpvmlX7sc1+2XnDetZUad0Wxli2ey4vZx3sZPdsmIa
5IV7OJGrodAlmCAJS6KH9unkds9GcThdaERY3OY9bVM0hruGRNnWR+1UGIhdLtNk
y+X9TxtLZyZ/YaCBiXalVU9Ukg0osYKsD38+RGl6aUW6JaRz6KDkjjP9r5qXlKGl
wdXaO96nSBH8jSqxgd4L1qgA96q3Ri70FshDAPtn41DBFQwJL5AkXVppthlXtQYB
Qqm6zc6EKXeUEuNs8v327crizcW8adE+fQOqt04+q/S2vrnvC2qDtnQfb5SD2KO5
8HaA71iVTa1ZsGFLvdMizdl5u2XeSA5FOfGqwbOWnxzCdZZE01K9mfByEqTnfOyO
QY/f24y5fuHXxmnk1h1DZtToukDR9iaHAMqjj/M+71R7bwlJ7BVvYT5q0vHoF6Ls
37s8AMnk4io43b2KdUv91czy25QDJBLRVdNC2/Z7fjjF8MQQscv53BH4k3FF4/1a
LRzkKuUNKgwtPnQPZM91Itfu9vq2EwRO6dm6kN+2kNROcJsNng9edp+njfBYVW4T
Xk3UVU5uc8+rGwkUJmof/Oya5TgcZXDOMg+9dcEaXCCPj3c/VRn1j/tRn1yGrKpg
B8JqTyB/F6ZDkfTQsU/HRyTEf7Bm2V6HBv9/wOxNmS2RXoK++8GSSX8XMQ3mikp2
SD8iAxoiSjS5zGN+oLM17f/kr0UugXpk/5FO2fouVi4rENh7GXz5CRvAf6wMrXrr
9gKsODhqEjZKiu9rArMrwEznU2QNAWzssoL20ujm8Be1hb/ulQ85T+UGcBioVHVg
x/moV05rGzxRVvISc1oSWl9Mmf92GxyNiKn6iVEwIAI0jr6xyOjjJWGTwqaI8Noh
i3iDolas0HZ8JTmK62poYGWQOFonH7J8c/enEXSOns4BhHj2PLtfinGzAbA1OTGI
bJoIlk+q2Qi/c9J5cDDmOL4EMyjyx52CpUh0ZseHczmPB8RVX1eBSoXGuvid/xla
L7V6u2qu1eweXtWtCh3sY+q/iBdVvWhbCsWD28T5nf6b9n68fZMb2xAIh7uEq6kH
bYyZ+5hFJaPikx75EfaZnB5KJOa2NziK4Yd3t/IHrIPSvyFs1TGgL6RbYBTsGG1O
3cxh7OH2YTtBs2YjEs0kfZTWEMhopUhxDMA9geeKlyQKveCsb5s/61nL/0IW7Elt
x/aJWcrYBmkMO9I6Ib/HOTRlQmH3+8o2JU0kvI6ZxACXE8U4cqEAO73lpLUHdZZ6
81U9pwAD0LUUDWPDfU1g+OHbKqWKGLphkrXNbikuB7tYjyybZZwLnH+vSs2078VS
NhIuMWPQhxEWOVLdza+FS3Qi7mUHVqeQZXTeNWqQ7nu+mLQWJ8EhAGrPVQjHDaLK
4i6/DyUKBcP8rU11NhYElUGZOA4Pb5x5cl6RqP0Vd6lpVMUGSvHu4fJTpt1klZlo
QfTTGb6ZE2Vq1db85ftDXavrjOBDUCr+WasK4RIxXraM5J24eMBUlqoQo5D1ktzi
tiwdPnsuUETdA0FrEy3pOPMqvqGMInQQpvuf6scxu/8riX91oREKB0CBeioEwTty
myHONU0BVWs630t1wCAQ63aa3Azzh7cA4b8K2W85GH9UsmOnkPakrS3W+VzaT+YA
VgXqVp+rCnCOSYpr16Cpj5o1yqEgwz+zH2UMBxnZCzq8E4MwsXu6ij49exVcd0hi
TvsyW7EU+f39tgnhv7Ed6fELAFYrCelsbSLtDFxQkViqDH9F/OKJs6FO+2mDV8zh
O7+3vNZd4mziUvq17raFjoBpINB5HvNGrVYXMMzAVVhnOc0CVUuq18ZekFQGBru6
YBwcpGuMJKnVPGV5IrnLosMPjWoRlUjFXd/yT8oTI2B4CDpcRc9T5XPgv74pN2o2
tG/wUzcMw1AVLC+ygg7M0uhDDFjZErTuLeQx18ojw/JWZutrzubLmepdor8+GCt0
iV439QcU9/RNazLF4SA/xwlF3SRA5ThdFik/vrmyHoJG4CY3qVJ10ZocgQbUtccL
/P+aNT8Vk3jAY7rEDOOWu5OGdqYKgMrPsDko4mBa80AvxMmLxsNGMak+IdQcq5Tl
bfcePx9XedFvTOGxWLNH8d1yFFAtT0/4ZWOoePmWCXiVRj/oPjyrP4zAg5NMKhKt
f/sHnrx83DdwPyNbOO4DprgI8Y0AqbnS957katEohLbOVb9cPSJLp0EDNuKAwlgU
ntRjm54Uzlm11+WWoLO8sCV5/xdLJUUt5t0OVZ6pFCB/NwHQaivYo6CnX5PpiilX
9O/TuFID8UtaLRSeDGeqGHFJVwoaITk66jjnuLc9LT1/34952T1hYFWoeGQZAU42
Cb4x2gpeddVQU/vSe6u2ycvCkhfg5cd4uLwXECk/HTjCg7RFtadPeY62dC3PczNo
LgV+Gv58gVGefbpDph01qRd2+bIb5yBlbj4icwtyfNVzWPq0HrWkRAEY2tRRh9Pk
jhdtkNrfaf7AJ+7BKqnjN6NxbHVzkOZztOOIZ9hzk5FSZWFUM41lTjkrpsMU4NFI
GkN+TEKDIEJrmVVkNEM6VXjoPtwWwjaZf9LxQKjAaFx7tnicd0b3AZk/6icRmy/9
YAwK0jaee9Hhe9CmsjB/hW/BjvXJeJAthZGUqrGs2pTFzrV2f/XKDLlfCCv6kIea
hsuZBn7rKXUo2JKfeam2fJrwjZXgQ7JUqnHXLxOWmb3/tqXipp88QD0RSr/jVixJ
59nVEw6TVaL35HNJ16+PKPiw4XAstJZGvUUWDiRF8Q/ixke+l9eypHLZpPblYlJY
mVua2u2ci/6zknavAZYUX9nC3hSujncRN55qrt5XZeltbGUTHhNX3i3szcxFH0EA
IEO9MsMYBYmMWWvF91E3RUVwEE0iccTDb6APCqdFoxHgHavGyFMLPa7H99MQ0KM4
rLWDxYHTAmblIiboajZ6vhO78e7gI9f0qbfIRKOJwfMzgckkXAIGiF0X4MmiKUcR
ItlxZy2THcFBy3BdMwW/sSC+y/vghT57X2BmQG5HEwgNwl/QmMUq8SGidTxCkmtF
5vXYK2ONLlYvJs/pXxzGWcr/cYyA11PefVwCw1wQ7XC8qt3ZT6u4Ulr9AhdYGrff
O3NI4+MNPuDoGwGjM/viA2C3vAYRp4CtVwIo+7SRj1aG0usnMRZOes02e+iZunzo
34skazD/9Dzvyj/rj3bD3vbludvhCb5bPlfWBZyXn+Vp94y9bvpCzDUnmEl2eDvg
F2joKq+ZUOYXZ3Erduvo4naxN9kz2n8FX1MX6bMaqfLRGU3zfTiE0jd5PoVc+cIq
7M6c3YL2pmCG/lvRhY0V/liDhhP9QQpY+24ofGfdL45CyxiYt3cmyCCz7wwfyxEk
JKVb8nDo2jvtKlWYY5o/XqLiyyfCjhq43c/buJaLL6OMhIWmeHBaHhxOJ3nSMFHN
nczrOcOQXwZ2k8Kph5RBEjAPT/nPsNOozkS3prBQo8+oKgwRLU3PrywgSNNa3/hK
gEDCpJCuiua6WvSPRamUazxY37j7WoXpht47nTVGWD4imQ3YD31+/Y5o/C6fqzvw
EiJEYLFUgOsFdDyLdUPNVnagDvsaduzk5p45+PfIYz4C7AyvSCFqSHFag+Gn64k3
xEUje5HbJGqOEXR0eCYuDwIcw8KeDtw1fv8ASnRSmYiF4aFbdJ7kHz7F7QUwio5X
BhnvDO2yUxOxu988ikjI0yxEPDYgn7b0x2jV1p+3ukMz1z4OYsRXyYJrlNLX3USs
9OatCbsCF9ge3Sk2dad+JtPQf5nFSsiTeXPHtfFCCSTegeaqRAvMUuTYC/ioc4uR
e7SDEfhQO1pbKcgUUmALLMroufSZiEnXQJb1WTjibSul3cXk6hsXQkE3giTzBtiE
TZd/B9LNh0Q7suh+0M99uHFoMnt26+n7Wvm78iyD+8vFvtN9y5VQmd981c/rvISi
vrgPmt+lmKkTyeO3bLbxfLhZegRslRmOVFI/BYXq47FlQJ36GsvO0SH9qL6C3Q8f
vbBfQeBHXO886MgOKMWTUmTpVIXLtnpnx4y8B09/hCQjvqKXaUGPiZt06Wrulmd+
VIqxN9p0U3Ac2aCQ/zmGzjgHG3G72V1JIRuXaU070cfH1PmMWuJut8xqNLdTBNmn
R6bRJg8IRFBusGSD1NAQE+ZnTHdyJ2V7LhVnNXxzaU5R/aVCpRlruobr758VLbLJ
8RD8+qFRqLXgF8kCqaapfYM/9fVDS4AOTI4z5nyBgDIOj2+zN0D0M7zhXEYzKqRk
hthQb0HNHhzkM+y+ULeTyhLzDxCE7Uuh7EJ0R40Zym5j3tMdaO9LIJQ+7N7e1+T7
7iRZZ/mw8SRE3iEedoIRHh2mbtjXiW3Dl03vxOmu6zE5duGCfD6quSLXQXXgExY0
fdkvjEhjuTAf0Rd5M22PX1C4TBPZrdwl8qUejAVy0nTBUolm6SL0sGlNYoDXqLre
ZyEDSPY3aSvOdd1BJStkOCg0ti00gjk2Je02gNCrJc+/eglq03gFUeqeDUns9lJ3
awOXmbIuUJ0nYQG+BuqUreohtLAv7e+bgS4ZHB1eOFkzdCnaroGf/HkmRkR4lqhQ
W7Wd1RSMYnj3XLFo1DOtU6rbRmq9cxzCVRcebUZ7SNDFtwDQ8xGFePmv/s8DsztQ
Qq9hfuyzr4Ck/3IdvHYeiR3/tVQr8nTkiglUUz9ZP3fr47Gp5tGTep1RABLKoula
W1FStL8LVe0u8rn+GjxNMl7MNVeqZft1N5zIN6Txd8AaaizshwULjy4YjNwZfC3a
gatrFyVOo9FP/O98hYA2Hr6Nrd3uhQ0Wv3ngqYTj+/1BX5ZbS36FSJ+oLmkhrPE5
1DCYHyaxQDIxp2Y4nex8LmXQYpwRON0It8oehiMJFNDcGoMdVSdjNisV3s6Zjhlk
D19oyeqi3UKKN08SStkYrwnJZP108wRwwiOKTiSSBIOEi+FJpYyLOycybvsU1rJw
g0PaqDTK89M+v1/li9uQ5tKCaeSmgUU7doSG96tUn4XlTnh6Kz8f005P82J8sfMB
D21AQjiuB2y3by5R3KfdbATDJUnxHQnz8/FBYaxp8LNoB3txScBEBjEajOS+TVAu
TG7ufMlkmRv2QTnfUiLzTJ0sW2vTpEWmALahcN5N5ruf75B4KbAcWc4KQLRYRYZQ
TyGW41w7qOxmW8w1p/BELpMC7akkjB9NpJa70d44Gmh6WqqSOZRNRYZkGbGjXUNv
TYNfMj7trLuieHBMJBvAqtZSHD29LJBxACg8JDuavi/wv1GJfPbr4kOMvohJKhoW
SNoob0sGNyPSIB/LN2qhs/DrX1aAC3sOfxePQShdQxYOK/mhtEhR6Q4DY9RwQ0nK
178Vi35M5/w7VtA7sX65seD+b/y+xUJOwQjKgTt8kAbrgtlA25zw+q8TFZWixnvK
hJTZppwaxhr69wZUIK8nUGWjgzGRAwkdOuUVtnTre+jYDZpuvsFd6qOGQpxA7Dit
mR0FnP7kkhzOT1GFB7mFc/HGYCGEmswJQLKv0gzDaWgFznvsao30v/w+GfIok4cP
KhlCb0PpipoPQfaCANvRgUtrc0AABg54raLwKIyrd/BYugfR50vmEUbfZmilVwfY
CwBipPFTxAOSvDD2XKBVmcFesIf6WoklGkEE0cFoyvXEOEFPUUg7G4hUUf4PFwDQ
RSen90Vhkv+KgxNIFu9tnvb+cEJW5cpeISssB6GP5qcThjB/nQ105aUdHPlrnl6M
jjLrj+ikgc/OkFEfMx1q50Muc8xSYpovPrfl284sL7Hj1Q8U8b+/L7W/z1wqkHuv
lEMu1iy5gR11PbHHQwOBeuh2taKfG/QpfWqoDAlmK00WZ7RQU85gnwYwb3OK/CaS
YW0OG1P9v2OSsWD/W0UUGgeMdJHxrCzH4lHYkMRFqCV4+DaG6/1t1H3+/2J1v9kf
sohzM6H3kKrncyNjwgTB76NeHjhekPoXIQyrGtpAEbhpMixEDiST2pAllJjuBEOk
ehfgyCxxeUw9EMrSLUGfNSl7uNVpfPuWfc0RR8kOm+TyiJaqQ3JW2Fn4BldNvcxt
/nIJRUk4nq5Ls4grl9nEf91OBzKIrzZK1uPyJU2o9nMbV07+AfZdozzfxSkKS6W/
ZyZTcvD02av5MDAfB+xtWxk4Yd+AqbCV1M7dAvVcAlB3DgWsDlO9R8qfFVU10+j4
MP3EffZkOGYYHi7sLugv4j1fvKXPXdmv5lkcu/vEvrkI3qfqNg+7SCmHz0GF7Rjy
4rnjpbN6LOM16cxhw3yH5S97Lij6H6tm+6Tm6Ltgu8yRQYDYhS8MFGkmDwJMR0R5
4bvx9VDnQJBjxu+XhIRIjGyeQflCqP+kN+tWlf/aOm+t1MVu9kNqNO1tI3td/sjy
+4MtkCpfeBzS3CQGDE7fhV5WyXEGS+5iOm13nmsiNovtusJPMH/OT7o9tXwVN5h+
wX1ZTHm6gyZ42IIN7L2cXfph0SSrxukMzhYIGjaX88NNFfNX+wHk9XuZm20W0Smf
oTCd9lSWts2CHpXClaed0U2UsRfpbd+OV5mtB6VYoCZfaGuXBj4GkdIMckVoA90l
HXzVicYhXBM4zVWWzsj/ihQAUQNf9h2RIktO/R4vj17YAP6YrVMJJuUuakBeXG6y
ym5aPvoIJX0eroeeaa5xggCBG8xHysRENGaxV/LZqtDVesf1iTff+xsvnJGS2dcO
Xd+JffBu34pVTIYEhJTP5S7xeyh7s+ENnxGeNSIwxCmDjrDY17L19zHUAkTmryGn
RT+PZlH+kh1dJzdCqRbKKjs7+8C2+YGbk0P6SMM3Y43WjQfnYMCQed+TOf+AOm0b
0VoYhONATeWF0zmPm7fle8qL8DBl5it4GzAEg5OTxmyd6AzWfmyU0D6MnWLXeyFO
9+ryfMsvjKsIuPwcgrulldSEKwxd+TLvyzluF07LMZ0nai22qRxe4KxDC+tJoJ3a
j1xcl/c7Ityadb+psNmax0PPKqA2LoOykFRTR8xmxomHmSn4WR5QKpIhE/SXOpi7
eq/DpURaG8aEEXMQ+POJPiPTneAPak1oPmGga/DKr9dEjNiG9FhmdkaB7vyOeFC0
cucb5AumfCwZc0HNSpPppOueQ3n4as2sN/WxC0SidwAipV703qfUYvI7OfvXqJ2J
+55njmsWEAMtAQANDZiV2GoCLSXI7lelEJz+7bhn9lq3qHauoBHY7orH6d3IzAQY
UFYugPwFLUNOQeUmXLdJs4R9nYfapCckNwbK+dqcYsQ9LqIjwFEWoeWsRWzsdP+q
924xRld+ReITEoB6NiGZ29JBTJAPusFJLJo4gxzKuJaKoM8Uol3JDtcUUCu7GhjK
9bsjAfcyJ8mX4vg9tj4KTmMBi9dC9ejBI7LPasUJ8NKwO2Gbw1C2nOaPOq9Qjvet
cNNraQsh7WlCqFmeNoRgCkcqs8Tp/o3FcJg6VfZJp53sSEDhmL+bbG+UvBYVbGCT
nPgkZVmgrwXUQoLIoEQy+g+JsqsWJNmT2kXzLEX8uNIjv6P/eqMXaK+jSPefDpeB
13W1gJTX0j+gxH477uuJnscKPb/rUCFijYDUEVtxD/fm4J6VaAk391w423vu7lDH
BHpN/xXAo9GXzRWvFG6I09cyLHjjC7UchCKi84Ib5JKD0729Gu0Ri2xfEjoQjgCU
G2CNPCWdPnQjCjzqdeIv/YVrNw4ytMl+CDeYjeFObNE5u87SGT0J+awOsFpOFmhM
J++Oap2uHUUPME4SlWTymEooObatsBDdDIskLgkOMQ7fZpb6emQ4AxR9MTNM5p/Q
xkRcNBwkCdsVb7n/kNd3VL6iPpBzBICOkivvsP8Ke2OI5+N1Ptu3W4U3DQbkKZkV
6M46MjeBDQcnPAui72Ck/GYiqB6efcEQFN0E7KKHYeG30RH0lTtM/hyv7ZiuHK7/
4vbscuH5voJZUAsMV+8RZ/YX0qjXSvWJWkA925MWSEnsSTNxe+I3TgYoIx569jL0
Csdlc/iW/ED8Z/jqcrakAQWnbtQ8p6ajHuohdIuIxJghVIcrHY4p0IglbV3uKVCJ
WFkaRcMveo5Rlg/wWNDaDf8ImC9Ii6rszPR6rwKNecfuZNJ7umj9sNE346cgYHft
RxcpjVdoK5wbcQ+8rROqO0nLaqPdNNRO1dc6PPFw6ODvLFAAkEurwGlSLfKe17iE
ly6J3KaNRDItxFGmtTlGFVP6KYKuCGU+1dvlBc4AUMHOtlWqRXbhsRmWwteX/tGB
auYvwHyC11Svsf8aQj6qpwyaQnrXGKZUvvunDPgdVE73iGm0QZaJeqwJKhgMQKOr
0hv/Gty3wYdCF0dZXqldxh2648sQ3ZJSUOwjg09t3AfADXDdzMSwRjd7M7y3345p
2Ff332Rdlw4a/62sWh/n6VNtTRScrAvHpXKIyG4pL/y65P63jBP7RptttuQ9OYLP
1teIPJDBhVMOlWq6fkKX7pAsPURCSodLH51D50cZVtjqVjvp8zNTabPktM1PrOIW
QwupWcjSiRzfrx6ZtZiNgL2GTtVFei4/XB1arclcAcN0TfyIiwNXop/a7QsrPlzy
rLyDnqfQzJFB3nF3mWNoEEhSfbqigq8IbXqqv9kAJnWZ3U/loXg8U7ctBRZYqCRQ
7a4PJgoOPAwDhTOjaL4IZXpnwcMRMcjE/hcXI+jDrf1y2q0ni1PyhcRYQJD+aYq3
kUR/p+oalvckaVBV3ii4ynKWoI25U2ryJzcQTDl5XmwDbk2/EFFNX0HbG0o/rw8m
q/omdItPMO14FQjDn4AngPwMii8pWvoyBZKv1EDIlVIdtkYepoMJHzEJwMilZjHb
IB+UHXBOunc9cTVNUCl4dxAW1dItH0ttgGjXYBvpplALz+ZTurhaHkT9nsC65jcd
IsozvEivChWa/qB12xTbfSnhPOvjDVbM13CSEofY6clficC3I+o5Z4FhPiuVhj7J
YOHqHHVD7JEPcWZ7SEQ9njDz2cT8NRX/3Hu3ae24VXOdR2gtshwQVrR0z9NCpQeh
ouWpM4fg/Y7rgPhxIF/4mzBlgziVjxT5lRzxTzNk38+nsLJt/28FKBZrjWdAbQXY
+H79+fZKb5cRIzpoyhZJqX0uriipwf+7Eaf5h5PMk3pXrPifgp/1V7eeJ8Uvfc6K
dOCVUpweY1AJxvihc8IAR6TEds416QJlY8sGLu9Tde+ysHtoa4cI9i+nfoeO0LoT
fsmQMoz6Daav3teCLSfREUYapn4y+ddgAaA8SR2QJzSrdvkw0RfWOf+VIA77YyCx
Rk443AUvFBIjlbsLrK/kns07v3U7SkeZqfHIClT9pBvFl22BjcSao0QXIouRIEjP
3BvYWKKdCJjwxey13k8RKGI8KskpFu01lHbrQD/VyponuDaUAc3SG+upuZk7fLSS
MQQdqAAnpljp0ZIN77HwXMUte4r1jGWZcXJ5Py63V9rc8lHYUOjHMqgq6TT0YlO7
eVf6+wtytdZUf80yXegTf7+Ef026+3a+ZV3mZeJPZFGx0V9pDsiBJ4ogCw2KowW9
27V/sjPr9Xt+HBWqGyW4sxELA3MvdrLr2kYB2Pag+qWQoHZJfgi7x/hdZrmC1mpA
xj9glwqG3rkSsTjhcyb8Ugiqg7eT1KQemeZdbb0D0hGy+oAy9zUR49XvV1f6wyog
+2dZBseYp/y9wSri1zRH+Zp7FwIs5uheEm4mVM4NV/AE6tig17yRXmhJZcdfgOqd
CE1LG89XTwAtXZBmMAvb9YWNJSfcdrMNsfSvDZ0MZDW9byjDwdQNETMuhnwrQwTn
k1yiRN8WpofxbUw0wdyDfc5UyM8+w8CRfo9jxabbpEAlGWT9L9nuRQPRYPqVEcXc
fNm8HVQK8ykLPhNlkLWv4CAuQbi/QIeM3gtZ0w16KKYJaRtg9SXTyCjiXw8GG6UJ
MBRMrRCmN9/9+DpoP51m9yoAgXU1wYJpZdHaXIOU4y2qTSIOKr6VepGzd2xyzuRJ
I/Y7BTrVQoitm/fx60j19aocT0VGbE5wmziPvgZteFReZVfrCr75UUpr/D41PnrT
J3jWLAAc47Ty15UueKu7n4BOrhrjtlIQ6HmaGXjNz7ueDbozfA5efdoPACAwgbaI
1e3DKSSDP9QCROACdKhiJcu2ylOUziOwZwsfLKuJ+cTD2iizIKCYeVD07YIO71OM
Os8z47sMoFaWkRN9L3cjUPQQnAr9uSFpYUjC5NLRiHxdDk3Fb2gMwKnEk/OHE/2B
4vUghjxN+3BdjLhjHVT6BqjoYCtZFtQSESUW1ONk4elMnifEtEs52l2AnFkwce+s
fQ66GCr/EKf6fr63OxgtKggaTcESU/WKhBJdgEoLffdezBqOJ1Sbh7mfJmVahBJ1
k8sJHAQ15/CntE+VwUpZ7Hg7HhCbECDoiO0yhmr4iM4qyXHkzVvWYIlayCce9TgW
MRNE5qatO29vrE6evQrOPZQSQPqpkWhHqaRjUOEzTF9UBEJz9UygGAABHDnUuTic
e6KlEb/samwiFdQsAdcLCHyHWoHYI77DmjTM8qjxM3rEgNoLn1cPTKKiDczIrswB
fMkou5wUroa/CDkPMqyP2YtmpAPg5EhVYkRB7NWP/oj8ULjXOw6qrGUseQCh8BIf
Db8yf5/iifU5p7wkgG9mFNSuaMmIEyk6i0ufz0/fBtK/GHmAfjAy/qmBuEIKbx71
m+ffF/g3utfk/XeBEzY8SSBpHLqcx/1CeKLAYMWDCgEQujP/+2IUwiJ/C2H6MUrm
2A1NDpB+c3qPDzRGcYM4AtkgI/DwQAb7XHVCx+zgrczE2TJAa+KiAHwD/ggwe7zd
6XgQ4F8YT3XepueaLmjpcvHgZKGHNduIcijuF5xdTNTsqffDiuaIyzZnXsu6JOmd
GDAjL/HUESc9FAvoQ4Csz0gPVyPwN9nLqZiVlMVddJ8qWE2jP/vJ/5M/AXHXhZGi
h1oQdilKBEFWkhJ20g+th+Jb4j2CkzUGiR4eMgJl7tu/H7D0ST6Pz/6kSMhrSpI4
zJcqq10qNmLggnGzpqbGXD7kYIUgA3V+cSqH8+HbvDWVcHhZC0NLpyBBDbRG9jFe
LWUsmksxLjqkuhtId++FYlsDLTc9FQ85XgW9YHo0IDc5uJxT+vwN1wIbHCcpwKEy
PcE90nXzLNHg3XNf96VYUbC3UKYUnkpFG9C+nqCqb3KlySVJUCwWWTP+wopcJ0vM
oUpFT0KrDSm2iu14wKCECGmNk46coAsmJN1Z+YjVGhbNkyuUjTBGGzOSTusO+GSZ
Xb6DZtOFbfC/EgUaga3gexVtIgfxzs6iAvLcBE7BpJIbWR5A4aL5/b+zkZCRGuD5
TqqczhL8aNppfZTVX4rNdt/DyXku2gpnwaat16DElzsPegm0XhhgQwzXNy0mkDJ/
Gi/FGCG2v+UKX6czzQVXGMazk3Kp9GjLLiWUqE/KAxe8+2r8+GcaWoOobGZ3eZLe
VBcNGoTXLYkTNbVqlqZgdsgy0KviskFGTWV10L5FQlCkyg01xPdTNf9+Mzn2J6IJ
OC0MHeiY0iOGubPMq0DF8W8ifsIUt+zhS2soqG2F7zPwCDMHRLvS6cIPpCLGlE96
HPA0CYEZmk91xFnxxzbi+5ATkKxU2M9mOP+eGXJ00pkvaAaVC39QAqctpyzYk6dE
/Xl3nA1VfWoXZQLTs4IQ9XTEpMb3U/Sbw38UlmrRQuW4M2I163Y231hshoo+G78f
rJ6dxivgSIK7n5nfezT+26QyD+vLBW+ilyylsSlTP3K9aYe2FElHf+YULzlY/8Jc
C0Ps93VguonCuCU08YEVKYsfAwweoBWaT5KBhCS/L98LeWHwX7s1AiyxnVP9zziJ
8KOCt4D9OaRuibwz1yGPKgoxUi3lQKg5DbbRXeGdJEehTSLyLq+ZWiVGtGtKMIFu
qAEXoropphkF4mcK7NinKzqXsKxQwfQ7eU4ACFE/DxForFThGGRkS5Nd0wSZeYHn
/jrGWcpnbPfuy7lSbQBwiPyoAYXk9/Yi95QujInvxHBgbyu0t9N6DUdy896RejzO
hknxkaPi1RtBo3MjQP6KVJfPEUox9kbULH6i2/FE+JBHuc3565QeoL9LbdtpQdNB
B2FQQ2/iw4dw1ElvSttV/x7sQibvjlRMO/ZTI8qp19hZHokHtngjTIrnVnzBlYVm
xdoBnShSw6rzvlvgd2FFbmKpXWnCi4rEFXU3jRLUH1pPa1+upeSdCyWdDRo7G6SP
4BdZy6hhGZdL2dtunjuk1Ms6sqW+TonsfdGchw02nXxOIeIOHoYFGqlJHJSf5+zW
gnLhT5dCe1V5KlTJhge5veIKyj0e2tE9qvo2CLpSE6ytXmco9u3Wx4XjB1D3AAnR
udsF+i+k63K6LaAHwb5ONoC6OalF81FjN8fWnlHwD0WMKaZBzMQtYA+7aLl6XFJC
ek4vHEZ1u5xKPOueXCju0eqt6Qw7pCIJI6+UPv6tUhU4ITYx7Oc+mrxTDmnxuz8y
bTXb3YcPxG/7y9Qhj0pOuJaOj4UMDWCzZBl2MPJDyrjGpb0jUPqStvTtsOUERNCy
/wWDAxi9dJlKN69gr1M0IjmRdbuC3ZxI0D1c/mVXqIrNjyTVFUogjEtt14enUvwx
u/3z3SIuGtcZyGdS+Q3jzrJzlzCQQhmMRevuS7wcXEIv8VPMWGNZBD89lvzZxVfK
0e3Cq6AV8e+X8vMWJ8YMLb50XSRFgVNi8uukB32x1FdR8rixOx4iNhhF1Npz94cJ
xmD8BfXuW2iV1FN1R1XgUXdcUaTxK0lTlnpfeRhqqCEsIzGHA8XV0el8AkpOodis
HKEESyqWNfYEdAA6OMWf3mhWIN2sLMxjLcYLUrLafyvWaq7r7FCwPdr3C1LL48m0
LTdlyDoN+g99gZIYLmD6UX8PWJF2WmnJyEIU/zFpOjgRLF683qCTXmzVGyuaGZuR
3gSDbe2PL1lrdNRopNmAyVQkmXch8ND02JKxnM4seDUnojZ7cwJsn4DZDRlskdtj
KBbXHtXGI2PjduigRZ7qv80bqjlvqCwu76Fou1CesAJfNbYD545A+D3CH/tJeGXF
oRRUbM+Sw3kNAfhf3ijrgAO9MkOC6pMrE4/lfDplWXu93oOYwlNkOAxlnccMpkIw
aTuaIrO4cczJL5F7qb9SxIahBwIHaWZoOR/kXWLmh0uLGZpl4nX1YUOq5dQTeLu9
oi+uY84wWxAmnqZTGd5Qd3ysr7wPxqB+fSGnlTH9VCjuQz+pwhvbBxPX5P89cSL6
RX1JBOzIblAbz6KrDmlqC6SLYBYHbL2xeFkRE47sI52sSys1+F/IQFGdOB0qXZ+s
h8/IC6KsOOttMr8NXnLPZV/KmILi+R6KR1BC4qc7Pty0VEyB/1XS6OFwISYubI8D
I/eU79Grd2YkCYesl+/h01rUn/0g56CKXwl5d2x9A87iReNLEL4+HxWHjj/srwKQ
B28bQU27GAJEb+lGUn5pnaag5aiUWeUHGhx3RtfUHOj1R0ghX3ayEAmMkWY44NNo
Sk6gaw9V8aG8kANokCSPLg8FybQYw5JsoIDyGzF7WR0WaF46IZOp6GlA8qDb9ig1
g+vkiv0CnxJHjQhusQp5DwYz3UITksc0PjR4QBLBKqqfnqVqjupoHWjaKQjY4M+F
K5ToYhQBdYxdmgLS1O5fePGJCieTUAMea+CsnbLbIQbPyDSpavtTbQG50tfkG5j9
5WJfPl835HkFsZbDKZt8gVxBSH7JITji81lTsrMNUPr/rh17zY87frY7cW+0lHcM
Y+TsmMWPBiZ+0DNVqBiW8yx4pKwMxOab30xr56yFY6iRbrP0QzzrNTsP0J7f00LH
o4fc3pDPYDpMIz4bCApoBTnEdnti+RqB8Ni9y8ZtDXcKSo+vQQzJkoCgDbsARcCM
+sO4utiZ5G+bnurl8g19ADl4bqJsleRF9a//GcCvEfOJKMJZe8xMIar1YatP0tjj
ZgbWfCV/uXzCOFi3arxr8cJm7WuhXidC1t86fP8YY8te4boX/uaVxAjvrLP6gSLB
f31bB+iFeZ6m1FQa/dZTq6sGDEqhnZUO+MaXXxCE8LTDf7T0owrrKM42Av/SVl25
hjS1cQm2i7LeLawAID97lymVfKfvu2YMJCVnK6KR4DqZi3ZjEdy25enWu+Ml+SxO
y/BB64M1Wh4yGMJOQp7CaAAAqndsrspcwd35CSxnDk7+urn/Y1qJHeQM4/jrV21M
tQl5CoKdMhA3J0xJrlWL83sST8lKZ9f/hBoYBHXQxZA1T0N4muYmsRsTNOD9PwM0
wdVgd6H+wPnb9ugfu+EM92+/1Y600RkTle9aIr8YjzPywYN9wSFWriyAa+1AZzZO
y2CuR/6Crrfjd6sB1iKbTxGSkJrDMwBe79Lpswnrxp4ctBomqMPgEK+khl0ozQpr
JtL4/iK9EtJ+bO6mtmoB4yDaucVUAOaovn5JCniX6GZ/8wy2d2vrgOyCG9tpXV/G
OzPJZ8WkrK/cQCaPi7S4TAzsniimTHIzJo7gMwAzfgWIiBxK07eAPAB5nb/SukmV
nVfHDxYptWF8qlV53cEEt1uzqh6FTrpdEJ8ci146i1A6kLdBZkBUXrONoQ/naAaX
NtjLJuRIyDkFAmnRI7Q9fhGGvPQ3KjZ+pwSOVT80UmpL2jbzZWX2oaSnMCBUl6IB
tbCy+JzXO0DA1xHCItXZ3pJ/b9elX4fdl7/YxDRmpQZrZrubQdrOCXCEET8BoY3T
OOABsV4UPZ3atDn3UE8nLCTERwS1d4PufnJ7R05Y/Rd6nt3eq1lJNPoNIt4ypEZ2
0iQrYk+XKAzJp4gs/iZxuf9EZNUpLB5aR9cJb/OlFJLWATmzjKcBtTs7FZN7VBbA
8zR12hV9U5BGfPkeDz+YAgZeRYrHHDbme1+sAAxlzq1ixD7/0FxYCj74uNscEjyX
MDxnWOJVQ/lwSJkR0kppsW2K/f+tnFkngyfTLpQwDBIBYFmVdNZoYtb+l5Xew/F2
OejH+Ioa58AXasJ690mbkyM4+n7ccKFo/60HZK2YJFWmtpeXroO++n8RHMcAL37D
fLts2+LgQ5aceTrUl+5zIzsVhdxAWGPAv0ODyEOMaFU9OdO+zrke7lgpq7U6wCbm
Nd8LQlUTO6hiqE5bk8gSIXhXa4+g+vs2crluDc7mTvARn5iVU8VMBJVJxIWZCxbF
kaFAiZyiaGMZbIoqf+PLjZC8p1WLLV1HHYGMg34YfOKNL76/kij/GGvj/enEL8s3
sDtT/iaxNA5drIVelenhpfaeXbLqQYjfsRtxqBNtGBVkF6RUJgIiYykSjo+O788L
88YpZJd26JWM7tCONb+EcmX4jQDwNmFE/gaoAdNMWMO+IuUzB4wsQ95YRrvFjBXz
4FTbG8mJYjHTUx8HZMcHjSCkxuoOlI81z9Hy+vva7jAHz2MFx4uwz4/VcuaS7kmD
xU9lFZacI8f0kR4QbxbTJUjhqxUTpM28K5zGsdVq5rahR4Q5M4E43Iqey2IuCjeZ
VQWhvJ1EbCQYdGaZczvTbDANegcPNG8hhfmdy8RfeEjTfYXTxV1ha2NrYLZ0QDYf
nYQV3pvpk4e8f2hi9xRTk2BvNsxztZveBtuMQDLpexttRiiWK1QKL4Es7/F8Al5z
5XXUNOc1oiBPg/Au0lLFhhnwPoDj3pcAiUdmTZG/4kVPYn253lUT0D1NbDuQrtA5
CrmFhHay60fH47kE4/ycJDRFKbPra4z+8L8HtVss/ft0KJiYrN+K/izvtl6e6U5g
Wkjni/csQ3gvukGzbUPe+HEjT7MuOPJX8HwxNiGV/cD3KK3+Vmube3AGd7ei4I9p
rAdxWyjxe5XerHH90iibexEXFhZLhZUAXBVojmAyEFxwBlyytGXlx8v+Om4Cy+ph
YMCuCU5U11OMRqE+I2AMtasvCbvkQBSL5ig92yb1mtAxjz/ipcbGjNc7Y67yxwNw
/po+47QU7ekjvw3vNqykxUt8brzEzTRW3ZR/5s36g3JzKHnCxtY0FQhK8r8AcQTH
xPLtCeLdqucTgWK3IVBQYDT0UqLiUQ2et1lAB+Nq0sbH4OztT36QD4K+uG4462EI
ZgwdfXqIUdtOhpNYF/HEUD+2NDT6rxC4JktxEKsXUkMXhmtrSDwgrOR3NP7pEzrJ
awmxg5LfSDjOnORFkouLF2fVa4uhaE4FE/xpKZ6YxLvitVji/X66UMamlLo3F5+h
6bH2YUFW6Wy/jl0qNpOSTE7MalQsFt81AHZU8iQkU8VN2H56himKS8FG40WPLqGp
TBYZJ9sh6vdffNWid6jBBFeBHabk2/OLqf0juLgtygjMI4a2DFoZfCmTFwapeeka
rUypFZgaDnZkb3NIxAjZkpgKx0vX4T44G1x/Dw/crepvPo9mRtfw1LjSVVAIwxUz
H0sTcDmbLOK5CdGXcg1EH+5phZEzEIadeuddD1y+kD/M4AbzTdWed2VURlLaq2f7
K0AGSQn2wDBjgeVS57G88O/DgMwWAH+pG+LD18ixOp57fyYpqm+D3uA93EYDikDU
KjD+GwPePXFv+0KrA3K8Xt/8JW/yPLMDyEwH1wKVp5kXApNBwlKFo4nsl6tSauWN
OCeNMBVMo6lyOxeRW/c82C3wGz3HTJTdSAXmuifboWvtlqKwvhiUNZonvhWnMEu2
l6r0tiQc06QCRUiC+t4jaBK1B+0Oc2PeaDB46sPvIj6wACsTXc1OJEFYYQ0yzFkk
oJIJQem5eWpddXL3aQyJcBdrEN/ZdMKqXKQNcs4zd0IDCQbvjJTh5zEg9hYJnXTk
W8i5OaFvgy7MvO2V+HrJh/RIJBs8M2GXbda+S36sOEFlJG6Ud/dhG/h7nviwsFKb
xmRiZhylZhpOTdDCxvlIyow64UePFjfKs2lkY+yPrLRpIUqo2LeYxPVUOEMlWn46
rw3KvjErj0Lv3BaAkAJI2sBcVxFVk5nE6VCBgBKUBMXGC4EvHCo+gOs+fBTRFWxq
JM/zQ4g8M11ZQJMEWW61BMEWZhSKQKy0TjmD1gVKMirFb7vrWd+Yr660HbhC8DgP
jc0LC/6UCpGJQkQhBV6aTRnAS+pI+Fd7Vno/eBYKAoIzsZjRJlcaGxcHKRFq1uqX
AhYG+xdv6ebT7FoU9gMZEM+1jl9fqt50EX9Gx5aVNC+GjECNwDRgvb0MvYTOpdy/
6W5SU5saOH26iFZzBVjgAPKoXtK5XXVQx8d9rDLoF1qYDhvH9AyXJpQfWdFb6tTR
4S5VSJTwQdd8IMuuq7HBAEr1NJo/AMkPK+A+5reHedIxgIDnWIL5dfoK+Bxvka0l
fSJgPXgXmMPtJAmTVvB/3vdm3x7peVJpO2KrxhbeRjEpmw5Gcz/WMwnSsGfBAKOo
v1PT/iMpq4F1G0sxNwksGM7XYqcNUdWf3hi2APIpcUf/A6dXfWocC+AnjVvuJg+M
TjsLabJnlz08/5P2DaPBlbDwZ36nw/VKCah+SN+UrMxbCqYzOIwCTEZlBW4ZOalD
NdggAN0n6VESaROYYp25GEPoWxo40FcSwKHfgWWOe8+toZ+Q4+qFfZASOQIKCiwS
QI//o/T6fGaLKMfROr+pC2CHzY8M4ii4G/mzXUu5zJud7FsKKghBrKPKHoP87GEH
AkAaEPLb3uSuad0F2k7QB3w5sx+qhJgOpMKnO4o52hkMFmHXV4IPCWioMoVRFaA9
B7+OG5fby0/uIdfrBksyqPGjR00TgtJTS2YfI9jauld1LMacScimIOqOeiHdZH52
fJ71zZNeTQ7cGEtq67M8QxpALGEyHasrM+yUdMdvEyUkTumpdXTJCVewHP3kYNqS
4J/bA58WBP3i5fY33QTNTG2TChEJf6Hm/CtxatiicD2e/oAM393bkNZfJSinVJ3q
tr1W9L157WR4xA48OilJ0tVEHMPTW+IUo2HlZpRVYCzcUk2ncvWpe+dIeg/4/Lk9
IZEK1ZVbA35MXyuWE/GdEII6j6ywq4c5lcB9UviPkyDrtuHqA8rF9itkG6zJBZnq
d3CX7kak7wHQKJmRkl0a8QcMRXsLCRW+tFAEKt71bmWGT76zQN6cpvf6ua8S5D+f
3vFiib6B+ShfDgEGxAS4z061plmZ8lmTk8YKiUc9zPipm45NPQl4cXaWOB2HEDoM
jIyy8JqIf2HceJJ1SUZGzC/45wc76ASYMDRk1Zpwf55YxLo8Pw2Xljn9mbuMO3j1
mBwkVqxqhzFTsY0FsJKhi1LQ/ETWCPQRxDztVCBBxSEv9DzYcyoL3jvrqDMV7pqE
MSKkYJRRsEqABi9K6A9ioqmmWNZoA65ZW1t/nY6x/WcyAxMYx4f+PU+J+G+PLEWU
8rq7EAe1RH1pdgqpZmwdenysJ0xPImbi4kRYTRr9jlnIIlEaDoInXdSwuicDbajE
cr38HRwUefRTaIrSfKuCCJ0So7MzDmDraL11MgF3siqmkOlESxluKNtMOymxMjFZ
6ofSOkcwmF/IBZHBNNe0+sz8V4mC1BtbtwNNgcjBz5s2TeBV1LCwoP4ZWsLxXV+J
jXIzqNDyH2YlR4E02tELKkvEC98ItCtPNWWqn6TfH/xbmKjY1vH7mteZwt5zZRyf
pmx1EE01m26TrnwxsOUfCPQrjRMi9OJn19lBwcwUlQj/taOhuBYY6hzODJcvv1Zz
2I8iA9kvxC9gPuYCm3FLMcN9OOM17nBjqBUdrLW23tNGTPhoNisxgI9Iwv8JsGkS
P5k3ZadMBdwJFS9Xe18vyMHjEkzUyL9BhYD8slGu1M/gHtImchthpUsqvIVikow0
8Ae+QaxhX3ElAJwmxvSWtgsTGJvWD/ZtjpUVUhuTUOGKOLy6zw2UKN9XZ+N01LBB
+VDYLr3YLRXoVcMaLMbRZD1jUSR25VLelInvjkvhZIbmzUmd1skxX1rpJR0J+13G
bJbyhmVQSpPms06iWhbw/Oh4ITAkVbi2oymq0MqlKCUqDHPTvXac6Ns6CUm7Kuu4
H1Gsm4n5Gc488KHffY6JCXMEvZfafouiTRigZCIBTpa7wlHPiEQLTr/bCWVg8Yg2
K4KFCvCXLkiNs4FKp9rXvpu8Q0T1gGXU8r8h3m3a8WRNSTTsfV7iCFely+dlNdq7
y1oZeNRNflWUgNw394T3Lwp4i+3yDfZ5zVXQF9HKfibGeGZ8P7npfQ+1/eMqOoi6
fS+YvB9PHUHFyK0K32JSAhDXkQ0Tuh8Hq1o+4HdtXURh3Pypz4tCNrehkITmlh7n
+BqNNfvWXDAN0WhFhBoR4J3NPePZ4+/TW5fBLFWQc7W4EVaz2XVu18SjXlXVj3Rk
FTcD/IKyAS94gg7h2F0Ks8S1vgYt3SWe4cEJD0M1Y5N2d6zP61p/hIMZnDlvvLGR
FqUS9gguw0lfqHb6xV9ZHcrqwJg2QUUuCo5v6m4lcNJZDhRGhI+jyircgJo3XH5Y
RA45KPXFPzG9nDml0RVou3tKWGyj3XAlrQOv7iklbmPbv5gDkeS7wysIRlIr/IAW
M+LhARJFLeeRzIQujLs/gdgNEoahoa4vuhcsXGTcrvw7Iyd7m89EcwIVvKj/IX78
YpiiEtfJASUR3IZpl8rA19VZFhG20SrJdc0vsVbn7HcIQI4HaKR1PpVb0n/rmApS
6C2Q3fPJfb7CY3x2wipPwoubDLrQnJ9gauOmCE6kPJyL58inEWERijxa3pO4L2eF
GuLIeVKpYyjUwuOgLJf58dxbovX8SJWNZLqyOPY8wijuhHf4B+IbWEKZAFQnlMe7
7kWBqAJjjK5nT8Ez8Y/9jHLSWeRfxyu0st+61USleefT1nonuQvIhCoH3PVbWbn7
jb4ZcablObMy7ZIAaLMQLZA7mKGmQsJHQd/8e6AmNbVzTTACL5XGeQsp7q6YP9rk
IWUay/fujzO3tSbgYJbKeifS6JqbL7RNa6DCjKqSALcMu1+9HZtZF/7sFrQtwbPH
CXqeLCCbYn7GrYoKWTVWWs3F0mypNA9KB/Ba3Upo58kJkUvbKprmBi7sSZfTKqxF
u/Esu2hhZSJkB8Lgnx6sdW9Khv4ViTmOXtdkyfI4dIJh1Dljua9T0OLkvrSRAL84
nGu9ta1/L57bdZ6f+iB9fWY4TEeXmcoHc8hbI3nz6pMa03639Vvmy3W0L5qLwdef
LzqxDxlIC7DSwXXQK5oOLpp51W3G45DJLhMakwP0+8H8imYOwdd11BF6a30NVrtS
2OwgVMhZUt/8gdjiAb84TG8Ar1OvruKYpb4wK8qot2a/lQNopSidIBXMk2M7Eg9e
fDiGDglK6ilunc6IExuCByd9882JcoSeIz4Fc4joKLIGN07Ja9wIRLzysWIOJelT
yuPcwQfvOJT5kQSV3l9szVbsQjd2A96jX+h/8GE3U6OZ0e4vFlKe7WzMTmew8m/u
9BZX9+6ujh9bQTsX+xnsSKbLPHMphKG+5s8DMNqSd94SL8/obAp+hI/QAi8LfjUS
v7C3MgvVnKO58c3lmNlJrYF4e/t6BHCq5xgLmLt7ZsluAlsBAS3V1WVWwyJm0mlW
/WPkFbFDFjpypxq1eaYZ23BZCRNCawiT9vVEvQ7PJbrEn76+3+EoOWTE3AqiXk3f
QMgAYQ4SkyQ6FNaOMUXe22xNIzhTm2SaVWkzCDvRr0TJXAgkLv0hc6xhr3y2IdbJ
WtLKRI9P0yYkpkJA+Kq+E5+1rUA1apGRxwKG9jbwj5N3o5XwVu4tq14BjeXicDAj
8GBywzi2dS0tVrx6CfFUWY5DThIte3x5XqmwGw/JWfKpQWKCt5bFK4SmCEDTnvAU
07anamt4LpeLfNw4e258GRojkL0vt76DU16uLAkD84ccsd26a7q4xrqOY1HYiK3g
WAfZubfK16ycz/AZqgiTuqbbYJiycYvMqmIA4H5Pak2MfLSwOcP1LVVpnvHFqW/f
SYSvB13jPOfJ4kCfM/l3flm1CJghbww00F6CMHGSKhXU1u7akyH15NyUddgwD299
Wx+1EuHm15bISptQXtps1lcFUS8LrRLfnhUJIe66CWPlSDp2hA6ymMQT8ulFwqNG
exxHEN7pIyPlQc8NHcLguKMxFCLPB/8NOX28Ht/yX0GLWDqNAYD8ggwaDI620R5J
A2fCVLx1FpvtwtFcSy+BTkqx6GSJoPizk/aZXdoy2RTTHWkjj7ZgrSqfXQ4WsSDV
r/SfXy5CxQJZ5HzHNzNwq985/8xLUtPf3Xq1gZ59eg2GLO8i+zT783rOIIFdh6iB
1aMD1YE9YeYIX0FpdXu6sdyS8/xib2vHGwdzpfYklWDBDYbu8GhcvjWtGiHfAwos
92bKBT5YE20oO20HZwWtb8PcS/HckBGFof+fSGZmw72/qV7coLvJtSmyRmTTiFPT
q8bIxumjUQ1FbDnkyuAKuV97URjxkEM98iFIgeXOhVB95FilqXg4cb1oVGo/0/Ww
BvDK6N7zXhw6Iy6b0hbOI05S7BWDnx8vTr1F15nDh/7/DF8gvl3NLtdpsj/SnkpG
LhsARRv2cSWR262qXbxuv3HkgMJ9c452OYD4CWJ4jbeYNubbWc6gk/lxZ5vjC9SC
nJTcNyGkOs55szTdVth8LQyWoFJWDYBWGrExauv9E3xvrAmFEBLSHLVESp/vsEbW
DPLNXHy/auMD+unWlS2MvBHQuWmeqv9DwsZmRn2DVoC98ziUEA/LG497f4y2Yz6g
pgMno4AAj6ApiLSk7EQB9nKY1qKPj/qkASBr9vE99g9yFKZCetwaIvmec1MYzHmm
vwOH37XicyKzRSOwYvviKn0FWLaSNople5ohUTz+xeBxUCQMp+wVOfjDIeXZyrUf
qSJx/4JijLS7NSYAlEnnGbfRmgDdJa91C+/NT4aj+f7v5655XFePa/vL+HJ1/sbX
v8Wlr4TKe8MZbjX1P/b2N3LZNPgMCMuUIEFa3FSz09x9EnOqoT1J/+Ea6X1H9sTy
M3bOFX0e57J3Vi0e5Rsr1McCk5NB5BDa4z/R1SOq1z4J+oera8pA3GD///UUx4AY
rh9B5a6+md5E+odjKXDbN17f49V8F4Os8eIBiSp5pJr88BtOQsD//0231E5hrP4V
9GGy88Ofly954lmEGBj3wQIizuw+qtBQ6f6ovDlPLBD3z4Xrwlu0JmLUzASTN7nb
fzdF1B05WuUFcldiok3ht+xsqqqPFm9JtoVLMmwSm7VedUJ4uvQVHC/y1mN0xyfP
hdWwEgL3J3YYQgLSxRtnJTpQetPuEdamvZhI7Qi3W+9eVAAXXG+8itmH/20kR67S
oUm2iNBuGT3dsecQdSt1+ZR6g0tEDn9u658mwYq3ms6iKmabkWyELDDQbP+pjKyR
kx3kd2aZmxMwj/LdsOP94KhYtqk1/dXVB+uJ6dhJsiPy5rRT7bjTrO6a8ww96cdu
BX5VJHb9h/p75zMja9opwWXSJ+x3TYYlk2o+FqAKw4uj85r70LnsNY4Yf1OB6LS2
U3Qvo6I5bclVCuFzY/tbI7zss4rWZv493IsERiLhvn8XICkJ+OGWyFcEpaA+fNEU
kOrZWLWnXhmJ8hcQO8T0NFKXY4ZIyBrvL1poeZMxtF03o5Qfy4V447erz/+0cgjW
PmNDRfZOQb5X2AoNqjUpOW/CMojnxJwLFX8tjLttbIh5GYOP+5swJeqXJ0czL9h2
bkMAQSV1z+m6ApoddxNog6X7cLtXMuAduepZB1hBsAiqFigTqx8nI0Lxbew1qrx+
UKOQDdTiUOi8kB8Obzyq7fLc3/G46BgzSDtoWaPrOR4OrDZ0hFY+EKh0cH6dQlRr
w4cuuRKjrFkQneweShc0qy1k9i8AMfFiy7BmExFRDfOqPIWpAB9ebMRs+v0AEn15
UFgQkdgln41L1rNYy5OxIRRURr37/pNiRmmb1BImapxP1euX/vMQGdFtvrcDkgqF
b/Yu7vcPWcbRHtqqvk0FGT9XDgOnXG4YiWeVucwMKgymslCd64ep/2NyV9E5nmcl
ClsaQUpIu1qDUAOXvmgDkL2sBPR7cyKrKf4FfWcWoWFPM5M2QyNxb7k7FqZznNwG
PIXdcmQHni1CtxfPNcJ3M84fbq/iK0Qxm8hp8KrvRdmwnN+iM1KkSeXLls0+oQe7
5VveGXSS3ciXU8ptbrzYA1fa0XPa+4CZSZsPPdATvBfa3oFNenAxrYtl9ZJ71maf
GriGX71XXx7YwGB7hwh/67frGW4e4l5Tb10Gd8cV1aYvyWjHNNVOgqWh9p/4hWRZ
dxvS5YcW3S/R9RpWRQamhmTBe4rpQRg7NoADY7A6UX4vzydm3eGBMpfYNVCh25zI
XCmqE2wvUAORswmMpH5ZG/HTQIKfVH469aVXCxbCkn2F31JCSd/IjmHbn2nHlOai
Iy0vrOUem70QBW5oo66+E055/TQdrDt8WckRi3Vo/GaJaO92f6uuEBzWuRe5rjjb
z14ew3nsb1DRbTJqBe4IqT0mi83fMjKDAGAphKbGAuq54TdYBELTokJGQ+tvrjud
pNlag2jg55rmvB3NDtNWVJ6hV4d3dHjZbBk3Pa0fkYijp6h5E3Rn94HWy8yPoDL5
3FhLU0XumM095342ITjbwIk1gFMJA47jTd+lSbQ2tVW97ULCXxBPU6huYWs1oVed
3aIVVbOlvR3fXPBQ5bj/IDZ7abRZOE3iEOq/vrDk50LhDQK0d04TKXzfTmOGZ2Ex
sssyzKEwPjRfOK+TEB1SpyCkv4uaR7X6/G7HJSei579eKZaFiocJgkpgcgCzLPKg
/TUl20BR9vCBhcQjK5b5c2kdlLlQfZyHd5q9KMlbXPDN28qtjXwjkBx12iCcz4nJ
aDdC+KXavp/lVIb4jPQL32Kip5HYs/dUOuwufdiITQgYSkPXW4v+WPS2kvg/y3ju
0SIy4bwqHe8CgjLJ14pJKsPneCzjLooGnRRr+Cd8Wlv4AZcciA7OO8eoudk4LNMu
FYFZVKY48HKlSIiaA23xOQuguHd7lAGDOlZI3Ry+klCTUtWpCkKBcaA/OjSEwl1G
tSiiuNuhyWwqH8tKWKbExIRQGWhOFGhX3AkgaFCKmyu6+382rp2X8YSGF0owpbyJ
bBTgj5tG9JYUIVNlpmzpuMEU1WBG/Tla7elkhuOj016C6VlMipIMtRnT3iCZYyps
9hcY92+PNVcoGVKYI4bvY07blWsTCgyVt8dkTdd1CM6CFp9rwdEezaULNuo6ZUkk
lSuo3k0wG45B8en+zf5sXs7bouYLkqWzoMQ9n/5Wjp7svmchaAwlNJ5JMgwAI4vM
cHEvjRqbiAkbnwwC4w0IAL1oJQPdsGhs8CaFcC1aigCvuabPt5KSheE1VfhChrl5
NVrC74sEWXznBeO1J+jhmVU/M4l1BZB6Z0OYliaJ2hS4Fcq3EBcn9osRYPOPWaXb
sV5S6f6yAup1oSKtAi1+h8jyZuvTz3Rfuav4MndGfxS5mexaoenIlhw5eawVCSbe
vP6s9gH/q46gw8Yoks218f6Y1xkiNfJ+ZslBSjjhLo94JHjnHN87NZF/t7r2OpjN
J/UIsT7W1dLkpmUr5kOe2Q5w6FHBnTxtdsr15FoIB5HNsx75XHU4aayYfD+LVnje
AShT4YiO/zxMsQLTPr48ljiuZ9nUAVpyvC8SCl3l7TxacC4S5c60LLi8Kw0FlD+0
jc6i3nt322mwREn4EVcty3aN8Wl9xnqgWAikdsUD64i13cyZWoWPBZ27P6TlGuQs
wL3waHN0G7a8zO0PN3+xbimAbmLyT6CJlAWTS9vcyd3MKqLorZi6/5DIdRadmRs4
Qpvg9b0JWIy4dnQWpFcMO+Rv+a0NZAfrhXvQFr1VPzy4jzv48KELpGOLrYAqOfop
grviUYTGv6B8+kVYRngWown/iKJaXEB+uKH41sg2pnWPU1OOT/UMMcLCgRu8xn6x
ALMn1ZkHSBV+yuuyxb1PW5YGj7/oXwDLDWxkhw2SHAKJlKKOSheZKLidYDqzmJzD
CKRBUuMmT/RdA4k3QTr7ia19Ap/qZFmqRKJ5oQf9YrZKuoxsqM8CbMLhmPB0jSXw
vev/lKHhxVkrviygfN5nNK/SA8x6hudkunZOj9T8ocETjCd+zxFV8Mk1DSW9NgS5
83xqB4j+A5WXipaMQv9juMCsBEv/79leox6jn/6rfC5iXfZ4cLUjIKmvwm8fHAHU
6lKO6lOmJ3ACqVC1g4uO/2f8EUsFnC71oWXTygC8UI/o0TCNSuChjq3UTErl7T5c
4+oeE8J4Sj0UTn40rRnPjek55+hCs+53v0rxKknmZrQonkHtc+rOR9CEqvuJF4Co
G9peI75KYxtZ1REaW0lMnHSR4WVnydgNSNBjkxAEEEIwx/N3qxo2whaGmYZFtWb2
hPz1YVi6LD/k0r5AbA7MA06EMNGExaYeikj8lWrq573of1Tl9B5KmoT/GmHPTvSl
BERfgrZlisVbE21HcHKzBXQIgieYdPKuxn/K4RCF22dsA0sdqhaFioBSFNsP9HSg
VNhib6pDSvaCSbGZHnWAqjYt5tecTh28rL+tx5YSLXSixZ7NlhHh4usBSGooCyxb
sqoC8gADUR/ypbi9B31YUthgxFhp55TxaY5H1WP6faArfMCR5Q3Yb31V46v6qXVy
u0Nyf5S6OBZ0O/J/672x9A6/5Lh7GAC8ntm0AqubGpK/yCCpdCgAJazc+tIAPMrD
SiKZiMhEQk83QgdEhKoIoCQJ/yFeJMz5A4al9THL/UJBfKPh4/AiN6oPHhFjMqLH
9Jad4XjC/IzpCMTlJ/kRkh2nrPVMHo0x7hPSTTWTETS3LB9xIcaatz7YHTPlqh1M
MjpyNtb2ImBvuUPKpBy3MA6YoHTrcTv7ZtXTqJwer+dKgjLDT78cwRPv8yLcKwIn
CMwj1JwlsQY+3/onB4+oOVQmVEoza0DG10vqJgx8I6RNYq3J72STDINsc6EbJX1B
f6AIVmVU8d+iJdnw7KxuLlMrn+T/gNEdUyxKGW/qWNPb9AQHNAp1X5BRXyKjiBJ5
V6lgG+2XVTiODISWF3/Mp1Q3scSabrE7ZMMdn3CrC0F8HVcWx7KUEMRoKjL28pK0
/QteUcxHa0EN7Ur/MYCZ0QLMW4kwhMGaMB07UIkaFxfLafTCcP22ZY/lYFINq80H
NfBZ9miuXTAp4XeKeXw19hZ2kTU3MRkUQgCiGpvyrfvGiZhxex6+Ow0up8BDWPhs
+YgDwyRw6HWRSwnFB/LAiVlki2g42E7q8vV/MP2Gyt1FYfUvPnqX4lxZNdOGTcl/
rE48cR6neBADwwETWP01/yEx6qGVAV82iCQPaUL0j7W7mhqznYDQpp2eaeyI7qb2
7jYqUCoSErbe4JUlGEMlLOhIJUvKiKkxRHOflPykZOOtXL/u4ovAZztoVoF7uJsP
DacD+/DN2nESQSRpl6yH0+tRwyLX5HysPcw79eo/Lxj6Px2UXZA4Z2RgXKk8sv/j
63z7pSd59D001kVZP9eDgV9zcdWb7NdUqscHPsKMD1eqw59Ny9K/4TqxeC8CC4px
MWx+o1QvyDPnAfZm71GQMM2+Zt2Ob1I90fd+nSvffhbsD99Footcdq0qcc4ZtrX6
uSNfuuqLATT9k0QCsysXUow4KA6PN6/5nzHbq/WHTWauUP8oNF/ngf8O4a3seqT/
dQqtrQPeI96aJpHLMd3rT7PeWVvPP0Hpdb2v8gSr1aJ4wyQnYdcpZVJf5ReSrtOI
6AkVplHdzI3nkPOpTIRFefZlCH/DHkDvUAWnIlxaALrIsHx35TABGGmeaMvJy4en
yXCqGlx0+GkQpgzYWLNXXKhPADdHf8K3/aJP9ngLsVnVE5hNRadGjyxL6m9iJ9QK
rWMshbCyWcXHzksW5pV28xwX5ubLL5QT197fkOJrgxTdeZnaJJMq67g63ATYZVaM
MTcKgwijlDt9IueOHQGDPElGLujkRqUvUocohK2CaPPOmQGcZt2DRd6mrZxz8rze
iC3iefayDL/bEqLA4Vcr0kgJIEbtA3gb29vSerCvZi2d75jCUH97x+tooma9O4xS
F+1ATKhHHpRWnCh7NB2QiM7R8kynE8M7jSI3cso7UEUKbTQmcC5WSyAeMwByxAJg
ZFRruiR41odX0Vnn3RtotGR0fRLjE1mRWpGqOxJ9hBqTsmFLk20qOkEmaye3pYbC
c38dVppjtalyLapXLKN35EOupTSHw47k45V1ekJK/waFmnSM0HUn6HFJLf3UsNCU
I/rSmTN0AJ7XAjn6pfHGuydIXg1TNhGR2g6l8ID97GVmibrfLczjvtb/JEMwVdYM
tBABNSEvfPoLqHLu5XDfLGnVUVlUkXcU8zp3LwDFhlMX6U2rWj6oNUrst5UkTRQS
kJC4gwjVD1MEhrkqRYfPi29K/4TLc53/54Hi1VsfJICaU9uci6A+aU39u9a95Spe
lBVBYinpSkV18UIH40vqstDVgYAW2sOdqVOnyH95r9TYJlrp9M6vE0/CIi25A5AH
0BiFmC0fPcJwTuZho3TO9V9gb/paonvm9vggh0JnIUxIwzbl97e/9gP6pyYk6Ch+
9Ku5d6aI3qA7S9MmhVjtggyABcPY3bRNlhhMpLSE2kfXWoWI/qIpE3gSTp6CcE1h
yWqQH4hNsIuSfOV5g17VooWwY06ISrTkJI6KegFPIrRQVjSZ70lEqD8riMYORZKG
sNE0KhsW2/y6OlM5iAyvABLrys82spPCFVi0oU0LGLnJZigN60YcKlU+scf+O97O
GCs2OxA9YMOTlwFCZ+SORZaXSyAhDGrwLQG/oRFLbwTfLvz01BOhWrhSUbwKicrd
ubH5RNj0fWw2cLyphotwCEkVaW4Y0UXAnQH4VW/linSfgTqut5gKAruZ6QDAodI6
MlvDrkYGJtPvuvWMr3EwXbFxWbSjMb2WmGkxeNYqdf4H7C65GhPf7i9RUxLiF5v1
G1NTB6SwKHJUvhziD0+KRq28PCuvaThVB/xQSsNQQXivSIUUxCqM7l84OeI7viw2
bHbnY+Nt7USM5L0lRglX7djf7o2f2WGL2YnKBiY22UpazFoc5+3oAZ57jia+xSew
a3GaXnqI5a6hEEEiqtnxQCiOyoCsmRp5ws/3ZyrSGV4vGvwBuaWbLpGbeQnP69Ta
3LSr88ulKsL+huDW81jH8f867cdgjEgdrv2aM2/Lg4gNlfjlOcb3rRg72csx7UjS
UxdIvEXWMyXfelHGxcEk00VEZz1qzrNn92ev05JBjEEND+MdI80r/+1N9fid+1Qv
PeK9ME82hC+HtawTJOKoBXjT4NdNBgCGiBAno6CWKr5DFU6I7k7FmdeslHnCIwqg
z05p+k5b1pOvmf+4YthDfeq64G0Gc92cBM557+bNmo+HJdQ0KKJkN42Hmf6g3jEl
srFgjTkk8/eSsAZ0VESbT+rPVxWzVMQq3Q7BY0s2UrZ/9JzcevN8vcNb473JUEth
u0KfDMGL6NxFAf5KIZ7lKvUpdXL2WSqR1bZ3P/i/hqJnt/M8wocgpsRzFsGEuv8h
a6VszQ0ORrZ0l26nbhDMDmEcNejecuYo2TpL9MoHvHDhtaRjeW3weSXrAYonpaTZ
/n6LpObghTSHF92KqI3MuHBl4utWBB39D8mUt+fxbTJU9E6BiHAhcHyZgJdWxwaL
HE0FDO4e5591qxiMzRNnCFim7VYJTN4yPjIrlyu1U7KycnUj4mtREMjSU0Uf8eyX
Huf/3UW8pgwLs67tu+Bmc4U2HdyJO5/2jQBxXgnA21ftq45SlINeEs7xrQGhziTS
c7bPdI8LImGL69akM/3/d5r37XgSnyUYImLOIFpHkFyHfzkev/9PZa8lZ3AVisnm
7FQIGT9IK5nIEZkRHnUYtx/66gfCTB1qAAK3IgNW/lTwFdBKelcmb/4NNd+On/rE
kQw9j1l+YD2RLPdE5krcRoWkgvLADz6gtmP/z5m97yoyiplWryUTJH4MFq15PDxU
oz5A8KTpRI0uuXn5ROTdcnEZfWIovpei7o8yWMjGWpobypp5dQWQkeP4q5J/mcuP
6qM/eefSxRoeVg3HiMBt4SjFFpCZFfxrMPyN8iwJBU2FEUNs1FaF/P15fWLjnZq9
hepOj8yxP2XaQGo+FcqN6OlDHDnA8IWOCK8FntVC3UTYrHB6m/ECSdyCARvdyziV
2RlZTpe1HkUxBz9lNhYzU/qBbY8yhC9PSNhj8kSThVlD8mq9PVya/QiKxNuUMQ7U
AfS48ACDoiuyejfiAiEA6EZcKCFbhKAMBD7p3952KoHMyhbcFAnTDredZYe5mK8/
sYVlnOnYkCUsVhM0NJS3o56llF+IaFq6mgnDy/W8ShOrBGnqkYz9BOdDBjEExSl8
kAbuIiOoOwPJuOLS+Hr4PHbuAhoUm5VqBiEVsWZBoXeBbfFwJafareKxsd5p37JY
P1rAFPyQmYvmnGptpu896Xutp5VM30osv4aI4S4qd+4Rh60AAxYTSqErwq2aLmYM
jrlHGH1pl+NupElIcHGqBBLiu2ATFMqFsw7/0rmHoeyYOHk1eWYbieocYqj3aIwC
pEVGqkOEn3SSMxUkoa8q5Sig1UK+Etawe41q7qSQOEH5TDy/c4fCeD6C+eFe6sRp
xYcEx2XD/1x7E68hl6mNK5f8aCt6td/b83mugDjwu+VjVwIJciR4XxRTrA1HwmFZ
8VxHZ822SueSNuDY38mnKoeoCHVP/A8WVYfMpP6FagDRVwMAfxFNQJZXIvn0X1Ur
rASw7LJenGspzzht84JnawqzOrIRT7cClYJRzv30OkrG7b0Qmx/DpyLO4miDCkbj
Qg5i39VjYIIaPsj0zggRI3V8JCQgNBD6AffS5RXfa+/B59KI7fJXaJzCnZgAmnua
tl5E82JjCwaCFKaryQQZwoLGFT0Sj2kszajnwDuy+6ger35SxEt92dC1S37+LsHU
yrVt/OcNupjtIs/GOu1IldmPaqhSdSmqK77zYcAJfZZQO8oC4uuRsb3gf4e7DCrq
V1iwmsGt9ZpuB+3X4llmL3GGhe+CT40hQK4BZ1B3oza4FVasYmh62LXVyHqZzunj
dHCR+mgBOF7rpgb9rRpMGmv75sY15HvdfTKHuH1cdxOHaJ/Lj/c9l1ljTbTlvy56
H7PceRlxdc946WkSJmfJ8rjsT8qdN3fxn6Zo6jbviIVHnChM3NeN1NNmpQO0GVlw
SmVzPeYCQ1ysYQ1QJYHmalH9I4+fOYHkcjlxkpMiCXUhlWnw01Mi/lIOvp2qi/UZ
HyQda7N243McFaVxuGez9yBMgF/dGonz77az1pCHebla8mwOoX53acGq2iIyRBMk
jSJ82dKPX/uLTxH6DEvFmLpL4zc+fBEawY9pWW4AeUHCyOs4JEUnxijGLZy/SesG
qyfc8g7MV6ojl3v1rr5rhzyF7Ltwgkwdv+8qFOTQsEOLTBF/oFRLgpmx0GD7cHik
yecagrUG2q6f023BmbTbTP9gfFEl0uS3xwDO1ZJ2rfeBxqdtL5HyK2mEuzVsHU0S
2u8sDCqhBddJVGGkqWJMYdf6ol/723W0nV5OBpQTV0N2Bum6cQq+Hbw1+8SlYHcV
vjUtDQaJXHXXZnddFb0IjZ2jp2Ai/HuB6l7ij3uJgCKb8AzcHDSzew7l93a08shN
C4bSDtArJV2IAONPGresG9bNqzSMCmY9+i0mhmaAIfBDHVeGgnCxrWdHA9ZcKfoR
oJ2ky1A2JZ3R1eTEda8/OoFbIIpZJ5AOrO8BJ9pj8TxWq5sbf4gmJReFO5eOmoax
zJUBVEpLOyU49KLKgp2ZWWyO9R5hUXlN5/3EaB+1wEyf5aLGl0IRoOT9xYa/6MqX
uz+h5SnlVuYfw9AkMJbH58z8FJrVhenB6OAKjd9g7pd4/Z1Y0zwZDaOjsk8Tp56u
PoVHGsacwp2CduC0aGqjHw5WLB1Fe12aV23XTqrNMChnPgY92TD1Hj+KQfgE1efg
leYWVSSBKupHQ+/Ydk3uxASzI5/lWNwl/elHm6dVNtXHEIjyRNKCW6OrbAeNpHz6
r/ULejR+QByeCjVPbJpsYFOg6il7HRe8kPpLCnnurXIoc6tQ8s0Mnji+8uYlSjax
gWzpkcvzNVS+QMaaI+HXH+kcUsVQc6KzyJLINcQy6AU7ZG6u/4Pr7pzQhNel6Jrl
rRGKUoOjjdn3ita7p0sLnOsUJeXJqo629bXsWaPfnr+9Wwp8l6q/SLpr9wr1d2/h
03rJTmvlc8vDxRYS5/eMH86HP/QghBYbvBhqRzJv21PNP2YZUe6zh9NxasG9Lc6d
nQiN0JXb6DsNDSCFW9eZFQh8bAX4WiVr/dmjkbpZpOeJANNhgBuLQgeEHCPNTYCz
EyuhX/nE0uv9LotXuHAeGkBfcgKA1zijTSiEjnP6nxedB7XxLqmLsOOeSNhOkdU0
HqRhmDyvOqb5hGANTijXUxP7uOX4CuG1NoyjvPmu6NhN0sYz0Sn0RC3aeXSotRuh
lCnE+z5ugtBhQIw7xa4vCtn7URfCf/Agp0Hf8fEAKYChMx+cuSWXYkaakkcQpbLI
p0k8teQlM16tqwHdw1PKm0JM2G5i3KXDjC/F3DoqwQCfUxZbDkyysyaBYnr5ANGA
iigaHCynTJlnZRwrjSk0hFcSYCG5c5YKIOyVSJ/vH1S1Ns4QyuZl1cbB9GYsoqcH
gfh2h/uPxCnp6bI39c13C9qRGUD26kO74PuwvgJGVB49Wfj6BQJpQg0NAmONDl/+
5ujuCYnew5U2VUZ/rNAJWESsRNR7b43LmUJJrZiNMItEQCGiU3U00o+XvBoqi+LA
f90+al/xBavi/kd40BWaPeSnfdZpWdlyQSfxjTJl+eb0H0dyAbOzBOpiqix+6u4f
2cAJXT0pUQVii4+mZt39eWaZ+5zszFQq1ZOhnMBu7XyKt7KlJ2Z2PwLse4AlzYr7
JZZUoCpgVy4DNhkjeM4m2M+p1holTwhE5MAPUHGUl433ZVbnZ8SZ1z8hfnN6STrm
yPbDFG7LlSXulzib3TnZvQrE9Ak2n4cIKi2dmoz4bCJ1roe15QjJzpzwFCJpekKC
l3uSAPclE75THLMzaxJwUWxQ/CRBEwOaGiaOHwBInkkx7tptlOJ5ZANKGugksAEC
N0izlmEyFeRPUDWxwWjc7hEWYZ8TJVsKeaTmVKS1mv3We5aTEIMheyW4L0eaTvdY
40uqmSaLCtR22tdY0WOJhLaDPAfZP1ghl8214p7x2ysMRu4OHBPDzp90nPclTIjm
oFAkSrO3/4ycbPRDcn4RgGtWmYCiASCYeM+fDxCXD37FsrIKQGk9ICG25Vda34aR
FGascW0FOxq2SIiKOjDDBa+tTOMQS0u1XZT7ms1avnr1P2hW4fxf6d+HOUrO2KXc
yBhYveIa8o/3HV6dYGfbe2i78SxBYUUQp3etONrn21OYFaJgDCiKg4h0LUa4tCz+
ssZs2+IuAl3pinNqWjSxetbKdAoKBxpfvXYYQZSujzPtO+neATUXDEOHnl3JOzpF
LkNDxluK2Tvb7CtErfi6LW6NUYmM8/igl/9x0JLXojyBvqDmEo/FLnPOH7cN5rCa
Xs5TttIn+Ub3qJ3gkKOJOskAnk8Eew477P7dOhnipJow5vEYY0IPDQK3J6iEUa+O
DM7Fqo7nUM1lUbuURNSpxjOk7p8lzgCVOQgHuvSaiefzHeyzSjyl3qYjtaiLcWCF
mZrQ3cyRzwZ/mkBvVo+dOqZpTGVWOzCCrh14rPEDs6i1fs4LVdXuFzmTYllrXIrc
P3VCqMvNNitCK5ljyTVLANmTlbmhqybIOqMpmdxDrZyY/Yn8kMBdNKo8Tfkr+abv
q/XVqapdIOaLz51S8Uza2wzvw1VBV993+U8/ecLUfFfixYsQHer9+A+cARQo2VCY
9Ali0ZEbQcEF0QDLh9iuAGrQYzGP4LowHRKlWKL3IQOStTQM4YgZv/yjOLR+DwMW
fhHbJ/y9O9HrdZNGW1KfZVJvVLwqngH0dU0zIe8UT1NjZEWzrUjvDsvax6plfrxy
mMXQ4mM7lcpxyxwhn6Zu/200I0jrt7nkwkJQfTF6xt283UIdt3sHJVT3xWnj0rEB
QiP1LGkryW8XVk+s3uRg6JL13EADPq8ETxguFy7/hu7VmfwJroytY+2ne515cW2M
kEJkXMPMof9Hz54CBnYg4BgPMPWsOawyptHuMVSJ8hyZ15+2xz2/rF5D37w1AbhO
fjkBw/J2dfUNpnrdY255FdFu5KVQo1E2tDU3x7k3D1WsFZjub3YOTYyBLmvpzI0j
ksgamIudD21TEvON1EHpOoQkw1PlSNAO7y8TZI3+r2wKW29wss14+IgNdxXj+V9x
/yrv2rMUvHcfLDxEn5E/GnIzZAS0GuVJZrqvxEMzQl+RnyXBrEhot3u5lYitrVvJ
+lJrzCL/k4OgAn50V/xgC3XscdiaGccVVuU1gYGnP9dTTZod0Yu0aHLC8lyZaSFx
bigdsGroBi3NijkpFrdl+Tyi5abOTXMlo9hkNf749rtx0uKYa7SqZ30ljRCqxzvk
hYxb3tvPC9q/6DNYIJ/xDR0KZWpms6vCOAseZedKXGi2znVHyIS73Qw0+mYUduB5
5Bj5xjHoVEsrwVbn4tIDWSy9sSIgZVlbL8Y0L5OAog93y6HnzrK5gHcNj6L1+hB7
OnkpkIEqlgUTg43IawD7BmkAsQJsGErXyugLvkBgKFQzYkXyrw2x+BhFefVZROw9
9F4SnSpbkTW/6SCaZUvqWkJ28k3K2wBLhlpFS1XOrvR/suUjqzPyf8JH5aiL56h0
A4ClAFTUMCLh4H/xuey5aNsxUokUm5JiCfs6ChYxW3CZlBeMJVfh1a+zWhM06XkH
bE/CpfDHoghpJWnz/ma4cqXUeVlSHoUcehQHKbFDNxCs7Io3XGc5dVG924vqrDTx
/i3F0qWjINznLbmp4eWbc8knodmFikxFo+ws/mF6XhMHEmPkyRJaEM56xjMJMD3y
QdFQ1JUMl2f6SRX20TcKP3S3/nEEmpvYeA1Qjmcsvia8A9vHYjKURacN91UQfAQ9
N6i5sjGmHzORtjHQ33FROZxsourFJHdknM3noHs6c1FfTgGt0WO80zBAgbPM1n8j
yt49KSFwm1WD/Z35C5U/S3XEGrZYr8hKtxX3/NTJGd/7IFtENRawtfw/Gu1t5UEf
g+yALbB2b1wiDrD1r1+xqb0vQEv4616Bx/fDqw3XTsiSfu7VwerU7HdcXs/SpgPd
RQ/Dl2PVqlYdes582K/Qqw3X0grl8Jj/vVvwe3KiQQ32UiR0RDIBJiaFJlCTyowm
jOfmEwyWXFMLZ4TWrRS8yzHHgkwNdKkbYEPD7a6QFWPpPeEOiic4I8Rv21COBWM2
Nl1FOCytfj9ihY2sxi1u2FHeQQ/+hEE+7uwOaRaL7jTFPzM1SBOP/Aaos6eLqV0o
93Iu6O1GMYeMuvY4W8iwpBWGMNPxzbNkr+jIHi6SQPk+je9CvmeBu8D4vzQVV3XF
8OfJLrbGmGT4DKkFSZb17rUNYOIKiukFIyfRmzk8SrlhpNqbOsuQHe7q6yYdH1YA
Yu7/J72SmfQrm5gR8yZzAHf08A6ITQ89GjhdNqTaZntJhS7k/p+jpH88No5vURUY
1GObtjWgJgAb/FMLQ7XN6NDmvJYIzi3GhcwCMaY0YSuWVLMb/ldzhMlw51rYT7to
Akl2Et59Rh2mI5EqlOqilkArhgnULM+sC7P/C97+s5iZvn2D+114vfrpUVv4dplh
dFyqFMTBLVAoJmoEyDHaZ1Jj2yrcUU9qlktnOlL5JptAJ75y1jJbrxyO3M1suTav
n68ogmtoU8/JI0K9YnqxLH9sQZISvvwI3lDtsEYYNmPJekPaRODZ1/YuG1hz+9u1
KkFp48wZFOIQefefWATVJPqXYCYAxZhXvurvUC4UB4dwjn45XN3REONsYVa73GKi
g/u8K/2yeXX/QAUUgAaKJ5DPyAik8jTyQ2733YoVGVmqkJyXXrzLfcVPQa54H2nA
tXWweCN3ziZe77IcJ0wzRNSLdJGalY+gwg7QiUn3lQCqOQ3IVyOc49KnnuV/GJvB
NmJUKE+bKxEAaHitOyPWFRFOmgVOvwwNY+/Jl/kVyK4IbmJZq0ZbKXHH2CGN6feM
LATiRZDvNeRTzp4knCUmrkMzj62omMNdEouJ2j6AbjO5lJdLcPRzuS1o+b75qnRh
GOd3ERBMXaDPZ7uMjohZagWI+iHMHFqa3Z1bv5w3hjS+e5gWJ39PytFrAOcgjAkm
TQE6EwztffjT3O3mlk1s+WXIsFIIFYGBFKuvpfOmU8S6IdwtuJNdQxziaUtgQsf0
nj9yi+Bx+V+87dchioC+TT3V1xNHvStCQXvrYfG9a/6AeQnqeAMBcBVaQQsX3y8V
RR51L5cNTfdXxtaV21oEIsnMYYTnbLMJ/zlJhcJopsO861qpBaDkFhbRu+49h1WB
TqipaCTfanuclKakvlQ5o1oVJbmU0Rzp+bLvj9i3ZnaaUo6hJVA7f92V7BNGRN3k
nSajtIoq22tNIZ6ARsFjG+MXMGzvWuoBOdlxRMyZXEZ7P5h+4fHykF5eC2dAmCbt
tD3Ygq2IpkEJ1pnzvFAa/kvCT+grHYZMbACylSvHWKTO2OGcw0j4t7VRi4D6HR/5
fDZXgOrKsNlELMK+7IizhIX381I8C2/iIwHXCCOZtweMgBqRIfhSYWNTYWe4lhOD
Qe4XC4EXBKc+47MyWGUX6yKz4PMgr67tse557Glix2vGvymjOu3hPA6NSxVPuCKw
mmQYhaz43WBLz89hJ+BHCCERGPabI30rcxybbtXb9E3YNA7TuvWR+RiphvtKQNjo
ZE4aPEqGD0M9OQTZ+etotsYLhdLU+ea84kQT4AfudtL3NgWWyKpVPaTr6PNkM9tg
Sv89HCtIpXWUW4pnBegxF19lUGJt5aHTkNsUr0bmLI27vYmNebwtxM/Zlatsl1yu
QDxzAy14ZyZ3A8AU8n64nEfmKb259N54D/WdT3HKZtsaiDbAAwZ2+5/vRs1lnOww
M/vFjJkW2AR06FLgKTP37Fd/qbSS00NU1jc5e+Ybnr1lI1fWJK3FeTFMpJWMq/EC
mGMh4qgcMVcHoi/oPwu20y5B7PDXXh2yCRDaxFkz+OBeSFzrwHH2LzoFPVY3FDXA
B9Yh95JDAZNqeIEL9LWayOLYiNzx4Os4nlp9igepRsK1tD5EQye9g5fztSSddXg4
/F+SIPayAMKWnuHw8IHfObNw5298nvPh7T7l36E4sN/0kzDslCFWNKLpu5FM2mBg
RKfZBcuvZ1Y6h2ahZn7k4ej5FLxGSFhqIkixkQs7HJwmF7X1tY4MXXtK+Tb810vf
Mv/ZBgfU3mU5dfFzvwF+TbpsPwf3oDIVaUBSBf0IF9cJ6HEJnp5hFlpWLEb6Jf/v
4VgnAoVY/F9/U4GPqY1ckzTQRlbiOTCe5C0Vos4gZQRen5EAk/mlesfm8p7j2lIM
vMbjLkfhjl7zSvzEVArE/hdMffMxdombD68DRSH9mbt25sjJFwNgoEulxEF0Q9E3
NbvcWNtuuQ+TbYZpudXMgsQdr9AEtsPoSyL2PyznWjFYRsBfjqs8J2OvxUneWP2T
18y/9NHGL7gbAInQYCYx9zI2JY/pnbc5OifNT2zPPUm9Fm/vJJYCQhzPnCsDwm3g
ERqBwZq8lDQaE54vgxObo+rdU2ndg0nxYvnBAq0Voqtsz50OmHURjICYaTYHb+yW
LIhYv5h8si1gqW1WRniyifjoyklovAbYM776RqTMy2zimNkTCqyyF2TPE7zF2a72
CHfzfq46OtrnnmklZMplVDn62sZq8gEGP9zrzeuhjbLY3df+noDLpHG3HrxN073w
wlGa/PaFtIk4YIs8Qmb2w6U6VntDyKqoDqhSbyNcHhvxyYrixrTRs8XpGTO7fdOR
aDO7VQGb+Vp7hDLbfjEoGVuh3QHCpK6U2u5lmOmOzQcYPZFAXuYy0SRKjWmlXP0H
tzl3qAFhxVLZd3hFZ9mskE+Lw1ZIxwiPddgLNzoM+KpflvlyKeRO61NVfpKOgP1g
us4pSGjT4YG9ixrwbkTaKfKUmlBUuBa6xEJquvxICSIJKKV2GTX8xw+OERDJw+F9
3+L//8Z6+E8sFJnEmWQRauwgSuUD63QQJ3DOkGE2pEh0MIm4haY6J51rtewVvGfl
oFj1GbGg783j3Qc15SmOxqbhcKAX0+3N29nE1AUB9bdXJQmwFIKIAFuFcSqYQkh6
34NwPhOYgOq8vjQBXYsQRhlvpou9t8tFZvobFQj8GA3QP76W/+cJIiHHT8W00GJI
gcP2bQFjbghZU2BfEwRAmOclySCkyDwnVLR7Uz3eH3KfWmFhkIAjWlwhZoB7ZdGB
9Rd5DdBjI7EegOGyB3NS8s36AfH5DoArIXUtOLlNNxvsthrUulhStRbXuoiQsMA/
NP+sbKCucbieP9w+AOdOhF9eSTe5wEvSGxRoGmJNx/LAVO9MvAs+YSocE5KpUwXM
kUQsTCxNFZhMn77QnXAahA5mxdmgoW+DONIqKG7cBJ1BQJU9SO5AzseZ1ac7Ttkf
xCyEYYzQov06MZIDbFalAQHpJvm3E6Vo/egV791uYYkoPJqVnr444tuBujeP53cg
CG60Cdp9Ry5ZGLnUOYvQhP0bj2FBe+g3va6LwLWtsYkNSpcdbAHcHPGmidjyY9pj
lHC2JKYenfBr6Qy/Dj8jWj2bKA9qt2FhhL9922hRXe/a20jLBzj0xV2ohqc1QnjP
aqA60RpgDggIgu8OxRRPPMdDH52g8kSM1v3J9kWmvFY9TW5E7/NVn3lpITIIiZrg
RYIr8QGUZTJaMW0o1LxKDHyFzz7Xs8C5NOd2WLoX9cALjMdPi2jChTFFGlvNJmAJ
Os627AKIxeAhnhimED+jVrdV8YFwMqztO1G+RbHTAKhO6NFyeE1V/KtGfUaD0nKE
J8S+7yn/BuoXCYOQA4x1NcHXgBv009ZZWCa4j9WRFL8Li4WBmp0SjKWyxmFmxpXG
L3vb0GNI1d3g8Z21N1Q7wWfG+09ynYnm6ub/Q/UvmrGp7etWwdTroHKnb77Vags2
1XMVlXKGPC3ZrMoFIwEJ4zzclZfy2tFPxB8LKNkeq7uMy0SRa4gHaukHU1kBWbOv
Pl4gDQ1mJ9wdDJdxCUgnyoUuKgtLS681AMvUNmXdE/PA0EA//JV1q+rhistPG+5v
xngitB5gez/KHPY4W19ShpHkAUOW+B60LMyTrBP/w87ohZEdvqqjFauaX6zW7Iyk
1KIYgZV4qI6HcgX+mVvxSdeCi2XSwkl9GNnEPQrTKmRPjQt/Tf3XXTf8xJCn3KYt
B9e5MVdu20IynBMGy980mYzwUcA5mtShMHkTTABDxnTBJ+rmo06uRJ/bd7sRnyhT
mB+vhkNSo1TcxdI8ipXj8LcbA39LCLHm112amPwC7K2INQGxx1iQHfK97F67IGso
jLhOWnx/dH0jlNsOrsP8fuMf+6AWc9ZEmnvIv9+lQx8XEsrDcDQpPktkijuTCCxH
3eUa8GNzXZxDV3WwPR7gbyHh/eUw2DRGsw7PVHT4/K0wM8JMN+lJwo//dCWsmUse
RItaYE4l4D3Lrogg/ysE+SIn4iJHLvZobUwGCmdY8d1rOWeKZfUC2AKLnWZHRff6
TvGQTOMPX3txfg3s4wzkeXJJ3OCSEVZQv6FRqbkI09zSzHjSx3Q8aH05Otxkgd/J
hY7+7sVX/7Y6pntUbIa+LhvR8mLxTutV8RkoPUzh3ITJX/po8ubNZGv67Khm+pg5
rjvdRxWOUwiD6av3iBQfdduJTPsjO3E8Tj9yrMzs5kzBoibNz+RsSi348Inq0PG4
kDVa+Lb1o82ECUx5KcWI4bW312Jn5X9YgcR0iJozhxOz/+jy47eHS6ri6wZiEOga
Go8/7YDua+2wCcusZAgkCAMKJWO7ltLve2QDEvYqWbVr+gzgcBJ+VUso6keMbgwu
3m37dFAq0xbtXxiQxNqRQYfKhW/X8wB8IGxrq3v33StTIKZ+Awy3v7A9Z5xE26KK
GFOH0DS9bkHXiLABIGqTYULRayyjCC5B1I+q6KG9c4ebYgjYSJ3ZGJi7RlEHRVHU
8nKW7NS7sfxSaf/BbjLXpJf7hCM2BPWiN8j32lYL6EUyyNk2vb28qSNrAJ3dvCZw
mB3Bq9ZSqjGDol9w0/qqFN/J0d7PMXA/6AMqZXqbK+jl1RP3wEuFl5EyjBryIMIa
PK/CtTftNJhuJommrUS9w3SgcaU4O7W691MKOLTicgNZlqQ/0WgiOqvACfsOh4MD
N5sded6fdQdtvv9rLz3cIUQW14O1WwkoVerXLo4L0/BeE7Ri3k/eFNAPIzHjmgLv
hP63g4RkOk+ktDRzae2OmmPQtPFRFPK2OVa2F8UYFXSdDWAdmu4BOBooX5nlcu4E
65VSyX9DW/u5jWO9fyjAZKp/BLb1KB8zEi2P0fee2NQpbfunYKZka4F5ZLgRO8rY
XGVh8raDUQzhFwqmtbSHv2Z7ccO2hW1Mkx/hMUVwmbYclbYxCr0k2P8DOr8Pf6Ti
mJB1+L9DEoSm+wuBn+Y56LSPpr2f2b+jjQIZ6eodk8ilc/hYtzTSpE7X9o7wAPgV
7lTs8N86qK+nJhuGWnR49GBfp0RNIZ1HjBh0nEtVBkQNMpMupM4lHsf54KnABsHm
QHV/8qfB6wQ37jK7AhH9/oyXycveDaPo5Ggpm21GQDw6vbb4sdBK66i0p3DUaeCA
rHdZ3pLpNRveo6Hdb/XO7bLQDXto52ZkA8P7tJvZqViCpgC7YE2CVnfC/SKvpBJC
2Aeg5QeYnsIXN8NtP/rJuS7F1jG8LjN77Na7ZWh93lhfgevFzwfg7HmyqImSEuko
ctdKp+3FwW8gtreoCsrNmlnx8cKRP4cajwNGLv0Km6doqluwYhLRKA/P8yYkZZw4
2OEXxZIazAnrhleF3Eq/IGg1Vxf0usYgOtz5CeHJx2FHpGt2lUJnEabinhUPeK39
jnLxydAoJ3s7mBu9GfvzrbRaQeBwXQ9L2wNo1dw56vKhteP/30WaFWbCg7ywFuJ+
f/8ptiIgtcXuO+JY9wTq+9yzkxcmgqufQdDOoGbuGbZJn8mJS3522FpcMlG0ipzf
CwO0Lh+mkl8G9nrTlWo/4dobOLLC97EbfvFeisjKgbFfkei1PUqqYMcj93NRV71b
5Dsy1V/ie2Elg2rNXwA1ILwGWyt4ZHPzuvUwsrqVeVZ4A7/DsCNAs1Eead7D4Y6v
uixFrGF4YbdgdVCu05YiwPm5jk+683eoKQSHWRWQfVfgboBMcq0GxBTwGDwVsNW7
+ygEArpHKoX3WHTNG+Zt6ub/Eh85YhWFBohgf2ZB6qzV6YashHYDnfwJW6wTP8+u
2SQOKhJkoYQSvRVtxhhDvCvCmh0sC6nbcm12k3r63dV9Ze+5bd0Td8Gl4jqrxGWR
/4i2KEf0wM3w+x+EUQmnhfJwdYZ4Weca6hhp+78UHPDHW+SjiliDQL8lsiLhKg+f
USfRTICuO/HNe8WSpT+qg7yz6UAyFOelfJVfdpyH28F469vNO+voNhzGx7x9SVhR
8tSVB2xlup4y527LpGyXn4Xee5e+X21SJsTCZsL9WLUNMmJbOTQc8z7m4gZXPxx8
jOxRBXqfBv4EIJYSlFTDtIREz5xz1mR9wQ9EECBZ/tZD0PQAfUqzCUvkmeMKBO/I
dKjmpq7Jboqk+k3V/cN7OoWz6+keBcPZqAil0L5Czyzi7I5NJRgEaVGqNYlKYC85
q5+2ZKxlbX/p1sizYAWxLcLO/bUp+6ZxvebtSB583tq/VXcwGXwZS8tI25M/9LF2
xVnUR65cFfJtsu/9kRz64N+0iEpbUyknjCukHVYAivDQT5TUGmJUkhHqR4saj01z
bLtc6halYCeB3xfWgK8VfFPSeZtyMI9Zddn+ii5oxc6USGHyTYtwRqVbUb5MW3b4
psupmS916RKWrs2SBGG3P9tqIzqZtbA7WAVpgv4pBLtzfA7vT+iFn2ONsLPXbRUJ
wvSgQJnFKPJXBV1fJw6WxUg/cvNNtv+AQvJeQTpq8WPe5QrIFv4AUrZ2Z2mKr09m
4HYjl22BHP4f5SBJ/WmmoBrdT7CeYWZSeTSBSFz6O80ThneIQN183j6A0Lu++Q+3
jBJyxWxdzTHyZhCofr+ZAaNtr2BssHUZyaM57TGQVVg/w64K76uHVjY3n6fVz7fv
OuH1UOe3j3IUwPKBjdIktQ5gWWo981gUPZFxJ0X/ZZiEGP74ygIz1lupO2/DMlhz
QlTADreHRVqJRIg630NDkRx6AigAA6k3TdcrwQQDblF41EwqR5jJnPpJvqvQCGps
7XCjH+d2FxYqwhcS5FoB/vNZNOKODxa7QCuvgUDvDQUsQDgic8l6gELn+FvmIDpP
Yx5+t+4i6YJ1ziObj/grYF55px1VMDEZczy7xjI9W+jlnxSeNlAnRdt5y0nkiXzl
NgF5F9owKI5r2YCsHWVw0ZXSiYCOk8ahoU0gohk+dYPywaj3SbDe7sxRVRQ6jU1m
8+ViTulZXWrnaR3Gz4dELOeSxsaLoE1u7LoYV33jMIMVjR8PDjmtQkly5QVZBeWC
JfVf5CVZxLosAfySHXGvLDXMX8lB4nf7SfBOdcrF7KXjwEZPyi1DrjtnewH335wG
arSywjA/cejMQ9tomtnQcf1KvUepZULjhwy0ybEM04iHhW/1Jn4llCB2I4oEnEbb
lJn62FrgCB73X8L4tNqKPg+y59VETc/y3BWLy3bgXWzJQvAWR8zn1K2ANr5umWqN
92Iv/hRUZkoWioqRjcXUnHpzknnUkTvjjVd0HWdcwkJno8i54DFnNrVpPdaZr+OQ
1pygwnAYnjyYu2H6UK6FQgjt/hDNuTIs84q72Kb850yZjPEkbFlAlXdsIOnIZPxM
xfLW8orBGKmAlGOXvLCYUco2hcqpKk4dvSJcnySgOD5QIZ+Pu+oS67ONXox8kk7w
LMv+CZHQt14l7xBTgtnyDb9UzfRK410zc/DLaWh/f74zq+xP01iilkkTRNNOiumk
VI+iW3Lprbg3SM4o+s/XTHNr2d8hYDLvUveYrdTjrbrGDzL5LJ9voMQKkDkZzfjZ
0gVPePv4HEwAuAlV4ZH7UkKi6L5l6AIGRlqxWzeHcLSLQmOaq7rrpIQCk/ARpNuG
eiMBS5kJtAv6ZrMWnu1EDWt51KHqFw/yJdZz9IQ7Avq0vL750yJGoLITDa1sCIir
yM6mjEgC6AraO2nNtNlJ9mKIE6slBRuHMJ2EcEqGlJyOyBqRXkOln7MaBluSDLbX
REqhyXn2p5LK4stZw02Kdri6BDsTAAF2dRZuEdPoeHS8wWEDvKZBba3B3pabKxB5
U+arm22cTyFBTF/mk0cQfneDdyWiua7dXkY0HjtTNFlCuFhVb+p4Gdavm44QQ/uN
yfSu0xWmCpOguIvoR8iUnoBmR6t9KEqbNtP3CU+UxGJ+aKyv4+osmZTJqSuunddB
BEBETXq+1eheonF3WkF1ccRbprowHLsbjqtEL2WJYtVM0eZfD9BzX8lxtsnbCe7X
3yWmC/Rt0a0WUzwfvWoxaYm6mv02gVzpnwoaOv+mt/jMKAJIsB1jk7MobuVHoKBv
65zOYmtIjdF37Y2t4q8S+N+1Q9rpj3Fo21G0D47FIU/5EVkjKFf7BZ1AyB7TKNpy
v1Um56ib+5yAKROkkwS/0j47yCUAQtG7Se+qfXRcsM5Qji7I14ig1qKiIw1AJ8QT
dFCMCutD+1ZhQnswGgXhC6El+vjEty/ylc189/iXFCUl0XDmtF4TwZnSzaKHjjlK
6Asya2zKPvKYyJxnd9t2qA1WqAS4VLEearv4bLmUd9YhUiDxTY/4JE8vRN0nBYFG
ftFv5XRpYxpAWwO27cdfy7Rq+d8qKuhffyACn3N/PjH4J4FHpLFbSEzh1bvDrGDj
k+zhIJqMgZzfdjoAGTeqARl+oqwgUqm0AjXTzQpkYFZDuFZSUMPRWVNwIxIMy234
V2x0/A+nMaN3q+4yngsQMbe15HusHw06+VO8uFV0hYquxdTdtlCD1UrJLKPbNZYK
8DsVx1j6rSbH2L7FMW9Ki7rp0O3clxOQAfF4VslcmU5vmtnzueYXcqIHmzDKnt61
5EVP41PbRvjoLd1lo2cXftFJ5rkZgEixsQP939BC1VbiRKfMSsdv64I3UGZahIGU
2bZYqyto8xv91IgHjqDUBJ6FKDascL8QL2DesER9l/t6zl/23F85WFgesmYKsfpE
nGJaFI5k49PGGaSTlfYCwszr7pXziZbIj1dRtpIhizo7720ftfZlrCyHfeceVeXK
v08Asv5fNQ1tQ2logW8XQjhISUALOPEuV/dIPrULPBb929ITNAN0V3DiEH5tDCFW
risT0AmGZRMKohPFTm5hDrObok607693J5JPEdrshsSFEl+zgZr7aStLeUq92HKu
U7WfNoFl6QOihK5d46t3SATN4sb9eKuN3uwITMe1nIljQ6o+JLsIPPlnIDH7NKnL
+vugCb1qJnA8fYUJoSrVrtoftmBYwZjMuaOOSYYNCI66D5PWlIfMuaLQs8xI5waw
XNMd4q477VvHbA4mAPfrGVQhZx654iUKatCm225pRmszCctILlQ1hM9BpJP8U3Hi
h9/1HQU2+wKoBr2N7i3p+wDobS4NnBfsVnjBnyTS+c87zY3uV3wX+wt28B1g23WZ
K5QASxdUPSUOHnpShQKPWi38jYHgbdwnk/8DQWOEeSYTv13+2X3n68EiK9h3ZTga
FfX4UmtgeHQa3hwWdnG8cS89kGzVbHawPQzfcDeXJ/ioyEXbTKnNSzLRIAsJufq8
vN4SNLPJIZkocvgUXPdbyEoblSJF3ngyU7/Xd2BsoeFRPMpDOXWm+Zntj2qjulzj
tIBGQ379OIZDXB15koGNHZoZYZQytkwV+xHBdzqWw4TI97+chpqDyp1mKPxtch7D
+QzKx2MFlOGaVM84FqDhbh3xnW2Pfpp/Ic8+EgtfLaW7NW4Fc7DeFP8ZLKGZ+Oe2
XCRIbpk/VXbEuPhGKe2ZNElaBWxf6/A9O4im0QN2/xr6OIhDrxrvWmLp3ejtn1Oc
EOrOD7m2GULkTMr8R5SX2t7kN0LrHhMDXoFOBIbGExpTb3HYbdb1UrxFFGJ9xRkz
JQl4aby8JUvcVyKXQwlw2y7stkQdp+ZF81JEL5H5J3QRg9rk0kUhEXTuhr2RM9/4
GVx9O7cWgo+4tUmpyjsCuPqqs53rwChWFYt5jNrwEJ2+F62HPJp+0oejW9QPHRG1
JRvgAOc6PDmcAz3q0zXADM7L0rZY39j/uhA8UQibNIe5Mx3UaanmPBKLyZezdMMK
V20Pkl7xPoNlNK5i8z06ObvPTUnNzbwnnI9ORe/2Sfc6ORrKNRVV0AcNZLrsGYom
hZC5Lf/xRO2mNKzW6MvrMsyI2SnEoPC6MYApIzNpcBaWQia5AljHhDJ976gJvBwL
wVm9UdehJdQJw7GcPKaB3Yx6T0RYnibPdGNY32RmwxOTZ6QdIGC+ZRieckW1oJsX
mV4SHclQKuPP0xQsZX/yorI/26+kdH8G6CvqkJiQDuTsBXB7SDtIM+mpQ8QsbW1g
144O940MGvATZlviYYUz4qdiewUmNv5YnV7aKh5glmH+Nt2rCQPViimIJLAuNW5f
Pww07d4e+T7evfSj+bNDi0GZmJAyXwWUy19ubf/HFZ4aQzXCbl697B4eRyLimWW0
Rz+3m6MVrvGDbRoGIx5yMDVvILdMdjtBKd6Bt2SCp3U5emyFFHIyeRwHxbfjA5rO
iqrmhwi77SpoJse1Ia5F4gHEtPuF1+/JqUmrm36fnYWbtWing8nCjuNQ9qkf721u
Tm8SgJguERnBU3wAPNd5p1Vwq+8wmnVnHKldg47/go24NDZrHKnFdeef08Vwuiss
49iFOqUWXJPHhaJfJ/VqAGa3bT2Wpwll0C9YjOfndpu/ICmM0oPSOoMc0/RWNdXw
jWcXujLGMJyRmPkUzm0XrPMZniIFYDibED5BSQOpWhpHLRUIfjNxngvBJ2dZZUm1
f3yamgQs7AvoSE5OwqVJeXVOFx8vXtwzKqfDMrrusiaHSZPg5UCHTeRqtWv+qiTU
PXuLCxUKd4BuW2ANwp6takvQMfKpCS1d/0VsWRhPlraUiKrhvyruIxqOUCUhzm2d
hjXhT7CQlOgdSyBkpr8P2anL5Chr5fRzamsESEdEQa6pT8xLfmbfwZqamZ6EFhaE
2hrvbr+3tLtQuE2fJp1lcuN75XRObTAyOn8LROntjhuATTneftbS3al7UKZCffE/
z1Y8Ya/9Vv93x32BR6Q7DlGGLuyJbBwPlFinU+i+zcrT55WAMV05VcECMcgkr2id
3k0SqSHA/XKgzXi8bTP+TFP9tFSUWR10gQGfl9tPz73vaW7wv7VM3u+0Ns4c17VD
2PacLOhMGMf2LuWW/uBFBs7hyALYQ180oZc8zDiZiCRaOOmPMFKSm4pa62HW1cnl
4hm0IBcnYAHnu//HInbnlgpmtWoE5F70/XUJHcL/byCiFRABjIzcBUHCLs+G4Mnn
CqMlEXOW3H3azUmhDGT72A/1No5HUFmx0uxJ26+Rg9EuHVsGmCCGxTQ7caofMtAa
fISuWkK4I6f/A+LcgS/zj0ntrnzTypSuqyovyOAfoxFZfYppd8BLSNE5H3chV00Y
XJfLMUyZGLjo7ez+Tx3pSXtrrXzy46lbYL8DWba49xhOK3fWTt2JHFhFIvzw72hu
ylmoo1IkykympKOgKr1inp1TB+awRjVuXWLisRt2u8zSvo31yO3PY8tUVN1QXxNY
LQFdHcMT6m66QiwzPh6Tm9kQjkfWRe8exjz6xlYqej9Q87x+ISru3m2ASCY8E1ww
pA7yr7NwTpX3B/XkWooJCWdCPR4rUMZVC3tC1v4H4wHmxlzmDhpA4i2ku1DFX+WF
dscn7zFQGY+1nV391IOQzmz7w6aPSqhEMw4mYqFfPInkCzOGYPrfmfkDqiVnQOiy
WI+GBfgHm4yaXHtilaYTtjIsCLKKj6bnbb1IHvBFKv247tW6zki1I0RzImtO4TqA
CJi/aZh/5iOGcLP+yIV0BLYjWcWwo6RtYm9owpi2qwOX2WIWTkLCef2jini1Dupk
x+fU0YSqFVYxJbxgZnibrjGvbwJBSV24y4mkmv3NgngCeuXCem5GoECgE891pIAS
bsaF9HLZDG7tA5l6DNX1+9Gaj6RQsEJ5Jr2H96i4xw7awcf0c8CVqscnG5MaUrcT
WIPCTmHSb+mAI6WF1zUGvYtRbF3zCLG/XJ5xBhl6JHFRnXB+eLZJxxBflQhN3ZTB
E2wk+J89W1Ga1nLmLSWJc91wyPFDCDcr7At/9WYoNtXI4g4K9YI1OEDceowAuueD
8roBWK7Pd23N8FjrHu2+JiCeWPn12htFB7JbLK6By+/y8S/dCxU+1Gj23lyqAQnO
JGk3Mf67wvuGRktkViIrPOR55mlbCuPbaPUaDVs2DFqI1lT/NWlPUnoqiCWeGed8
R1x4unr4FgS0/cMKqMxG+WNc2jba0/IMnzRRKHcDVC1aAiYT7uyAPLoIphIFPNt4
+hQVSaTaJ6+RmAH1KFEebF03IOxLQdPn5UPbIRHgEhXkMqgr9c2KYj8z01fVhq0e
oyFGcLx5dRLTAbKCiREI3G2ZGzdE9C53oYf3WXUYmacErGkJpbCqVOOfKiIBji18
AkH13gM43WouqFsMmPqIfIUlQQgb9RS3UW1nnRYW8z5imWcdx0p2STAiZipiBzYp
qA6kq+eH6+Dm73JEvcWMhfXNYf2X2BHMLrXsWEatFqs2drV0NJ9bztExIAifc4VU
4twbUzO2d9hMRef5Tk/B4xGmvoJMsRx1a7Tjkl8QDBoIYFDM+UXARAcXXaoJTrwJ
6s1XKCbfelEusSF31/uvdeMjM4dcQrSWItZswGotW6Q+kpIm6I3fPDW1XsLBA7cl
NRo9EyYGs/NyRQiKFVHd21nYniyd0wbz9EE6KGKQunsiyEMFOMbLZ1ia/xEITOgj
iP6jBuSEKqhtBkwH7IBCWc6BBZKhlKSza3+W1gcpSkdwfYCSSDKyTIQEdKiSbeAz
iW9pF1pU7iNpYE8qPkVQlMauHm6lf7a/TzbarAO6tSUJTvf+owbm9+0EcLSAnmlu
gVr+U3+DwcJKnUae9pYk8VjLUHvHF1RHpo2Pb64nB4nFglEiqh47dHN0r0jevq9U
6d6A5DegbwU9GZVfcVmUwf59fZeyibiDxJrAnIeSVYqWmmrbyYbHdWbSjSKtEP5u
AjC2d2HoZTBhq9NInfN0y2VTNd0dYIS336OcB5YZBzPkr1lnIX47FRyBd90msZCj
wZvorOxR31p7c08+oLTFaiesUOShPf581V1HqjmmZfWtsw18EogkzBvN5+/6nzSG
GlH9r7bStEj99Z+1xI/87L+dCZwSsdQ1KQBYYlBS24+SCku04VgOhhsLlK0c7Axj
62A57LoAl6cRQgJhIVN3Pba6Ym1X/HtxMzToq2QeRrcBuxQ1G9LzBALf2BjdoEHt
iuwXx5fUPNb9CnNfwkbVPUvxVDBWXoImcQDJvmmBYtrtlAxsrsvYX0VcRoFEjbtv
rfLHsxe1sLaqhmVSWcSNGZyJ4rgqLzgor0RP2kz6Pb+q5vdySbDowi18SklSUFTV
09BQgkRY0UIKmYunIC2399oSr603C696TeM8UbyxpPwSMginfnJN+CFeOTxlMHET
lLfOppCwy4N2It0r4tAfBRnJH+Pestf4YOakYttiTCXng17/DI+H2TFuora5nuMM
ssEvIu+F81xw5htcnzUjd9chsZS77zEf/otezQy5NlCJ5jel0NeESI6zBR7CMhYt
sA0C0OqaHXj5JOh0NgGmC+WVGMlea14UQC6W7vuJfOrxmIvW/gza/BxPmsUBKfcY
ncFqVuL69/DicMTZbKYXwY0KfwFTon+tKP6hS34XClQXrUcG/SLSxWcdiQk0I2b5
RlyoXiJth+sIxKTLPMUL2ip6U9Ye7916m5PuQTDKFpErRuQfjYdxSTwcXw9loyC6
RuTuBcQj8e1qc36TKhSulUXxvKggzmnR9OvBC8xwK/8me3sDQX99NTaUEBdjZQOC
GvQF2H2VmmdbbB5hzi7GgIx0cMcJhKUw2VUttR8fsePMvp1gM2TcnYWT9lYmVrRE
YpygfNXt8HBmHQUz3tgw0eU6NarY532ZdW9UiPCfOh6atGWWmhTib2aE5fIXNABF
jYAjntob6PoFp4AiD1j0m9r1z1bosH3b2an9Apf+3PWWfB0GfLb5CShoer8/VoGj
dU1rbQwxgNXl9QH1r0B+taQns8x1fkxclJn20hsVfChDGEqc5/RMrOZZEhvgU3qn
S/h+FXI+9m5j4EKTdCGc6C+c622FanM+jY2+WbTiQcLhWeBubcStRzpWZsVzeViX
bBcppuOWyxhqctvydZbHePvBBl0SRcE6vjz4ftnEwCgiedbm7DUREe4AkniUEMU3
1ODSa2BhI38ECMOMqMSCd3mGk8fQA3kMeDtY6hYeJ0jOctWGF+IV0A9QLIrqPRkG
9nPE/aU/NnjI+dGUODbTmyYDVm1cJwQ7zhrTuypi2mA3j7uvpgC218kDuYmy1fcB
gYXTIqZBVwY7Y3kgzFr5TmEAgYKqbw3vBgqfJDPvKQjJAlGrJnbsnYpHq40FUbbo
nJh/o9EakxgZrYubmlu3jSDJ5aNxRkS77E+5Up+ms9AZ9+dPUdz1gwJX8txd4gWr
k7N303jK5O8nIThiQC/U9TPbeWqdBvFC+G7aCUwDb4WjiWmI6imy4v47RR3Ji9Ym
sNL0hxLjH8rqqR/2XWLROPBPYBY0nvs1el6lX/Fo6PVEgdyWIYyLYB/w42f7oq0p
5KWFNcWmPJNhRyXs7aCyrYSRsJNvqHtFj//3Dht5P5nu59aZzoKoSLncmxhHSGUX
Y0Qa/YWBitMGFOhHZDjRMxaXL4Ar3FciV4IiK8t23zXkBi5nvvXDsOK3cFQf/LBq
Ha4WfGqaGXuORJa1sodbNsKW/Yki6V9vvXCJSYNyde+cpV0fIbymt/lruHuZ1yGX
kK289wHG368tHpIcBHx7Z51INlFiPfSpEVvHd6MDAXyW6vQB9gjA7Nxa1OLMVPxz
hZI+9jEjF4L+t6N/abvFkgqbAfn7+1eslnxZmK0GrxSg/fmZo+Hu9wKdHZC+5coP
tOV/YJJzxSggpf+YvEqaXggq9fv+aa6EUnR7khc6WoErpr9tYAfljd9duO/K5Aem
iydlSgHFKlN1t+vpO0dRyNjyPGlhKBuRYS6hRbD/3tdTUsnbpz4I4QTRHZ6PKYG4
Dbt1T7mMhTLPN1giYGXaKpqo7uAGZBVVd/Eyz9mE0LR2HPhUZRtjGjQRg2mfl5ya
M4VEYcosg9idYgpQUol4OTvPrpNLfDspeua6Rskd0125aM4tWWPI35St1lqAH3mP
pqdsKYtP/zolVRQynz4XYmZ+x3YURDLezITw1nfjWDESx09w7HeSyxhWjIULWl3g
t4lJaNd8rWGV4Kzd6z6uXqqQ2uPikePYRQy1QwnEnexETCEjPbUSiN8KFx2draDD
8wtxeFZlFBXl9Iqr327N5A8z5HHliKD9vpe4v/Biw2iWmDTHyvwVrCpPPfnztK1d
2nDfR/dcMXe+Tv1KE9r5YdRr72umQeTZy8Adj6WOPrRnJKl0S4IwNJ9VpMfUxsu9
BBXBnlbigSRzpqPo0KOpTr/soYsx3JbgwQHZOeKkD4N2vNdyA6NaoGw/lxgK5R/U
gBDyLOa5/417BWq6J5R6kB5ABvalR+o1lQ1lmzWkUFVe6yt8Ut/z65oYjzlHwPBd
MCFHg6pt/RgPQA4JVkkqwfFGEg28zwC31g5a7/Fh73V05RG1SzBuLYCxrFQ+qmqD
dR2Ef9DiNy6cBCv4Lq2beFwW7cFdzIokSUzL+iftM47I9vaALDg9+1GtoCdtZqJA
4RaxSmvWLOI/ZeYtiW5y1qgPMwtyLOzwyg2he1v01zZrRgLqK+yaPjTXAn1Fdeg1
kvK4UjlWRZg8iRizx9v5nrnFm/hRWOXqeQswj9TB7/9fh622pnKBK5XtaiMFlMur
tmB5qlwrPvSrkSBW0P9rAgYFhFRSR8eaDMiX+11Ahl7qJStMG8+Tj5Auex02KfxL
cWs80OVdQ8lLtkacyM4ZYXyIen6k2JCbUsfj3Fv3Hc5AyspXkZQfXgc2DF3f8PFQ
GsOuDdUIUGv1HSGoPt07lT+1oWEpIYVRyBP02v194Q30XXihTYQB7nx0fQjfyJId
acMF7n7CK3kViH7dgX+oX5jH/pO+9bZ8D1GIB/S9UTicF/+qiHjy85Iby8WomGTW
wdB6ZqG6Ez/CmYCMzBS73xoTNMb09dPDUDOBxMRi51RrlVDK3IFBE/cNN4xCHyFB
qQjheLYB5Hf3wy2MAaZK3G134RWJ1oShvbG7mbG2DDhuWRSgJ/L8H+bHOqYIsnGg
XX8HgzNX3pBPNGudzU3KBqsbmXlKeQW1g1TilgPagqTz4yj/hXFWojeMqU7re1Kh
nWBLs7QHe+u7gqIPs74zslTXHxqPM7x9RSaJdAv7deWrbSkevceTObbjgNvVfELF
D2A8VR6JL8Ro5jemahGPoqgroN+86Ut+nRue+9lyu10hqLWGuGIDxP+WSUCVqjpo
DBCg7W9gCy99NSwD/T72Lgjy46rAuNVsHra8xcJnXLTetPaVecaCcY3Mgi/rrP3e
psgWlqW0dghWfSiAXkDnFL1WOGWJV7sOnH/V/DHzfZzC/deifP06U7m1dwI6fOrV
Ku+GobBW5RVHpgIJ7jv3q3fLj2o7UE/do2x8WqkBXztIgYJtPHUgcR/al3Sf7g7L
HnsS2tIvcYcVbdTVCFL4qs4aRsxN2iucVF5vzE4c7l76tIDxMBnTM8PkUifBH0zB
w2xVri3oUpgTjClS0/NSsjswIqTlGHx181ul9loZx1LANy73EIpRfAruupkJR5qB
XZyP764VdwDRz5vuSWcGO2RZoT24GhxvXRbm6T9jBMY4KvZ5vizZbHykzsN67ndO
AXpiZzfHtOyDPc+ABgfOYD0KMCBpF2W6xFWeB38zNck7+6Mbte3pOKgCoTnboJUD
uPYs0+eN/HKKBLBrWUwpYSbWhBrnEabWfFFDus5vAcIDE6Ds18egMWEn5PbddiJK
j/qbekcDqHjZhpBNZ88IQFS8pH1uaci28cpwsevnCT9DhjDTTfYfrRa2YYnWfGXg
p/qKS6IN2Vm/dwh0EPBu49SlyM+eZKWx+IR8Exq0gK1qfW1IzOnU5deXSl0xRvkb
BIFZxGiW+YOF5Au73n4h0I3QCbbbrMh6yrc2+qE3Pqm0sIoSEWsNF7iqJCeLaldH
/dqApm+bmBkE+6n+2UyqMHm7zfVHpRSRbX7FTuT59vyz7KBa8pxFKTDhdn34VaKh
gl8Ccex80UFTrQvZdXmVe7y3fNUL62VICqQJn7dTW/DgkhlUEzy6lVGM4K+TGRTt
X2RaNG7mVDkPCV+lqNI9q6Pacsv1c4jpAOcTj/yvf4dT771vUjN87NyhAGQ9YXa+
LZp+7uYhLliPgkxu9FtXkl2mR6YuBTp764WV+xj9mm2j+MRveqXh8pWZoEfuowYC
u6tCt1d+yzEi/uNwA5FU82wE9/uSaWQPjGtFiXVwmCFZuOpnLOw87x7E1MmVNTdA
oW6/DB4vUwCJXHZPa0RuREdewlGF6ANRogWFsosIs8WhIkc2MYVYboHTgq7Rqkiz
1e3647HjWLNIrZyXqA4tQ64kDGVfSsA0HBJEF/caHO8HEl2gW7gtyEPvsl4EF1Fg
nUElabMUfGwUOSz0qA6aZ42wpDr7rDDpYiFT+QSfoyHJVwaB14UPeFULwdiLenjy
bQqMIMdqwzjEyZIABg0wGeShTGn4ZJrP5i0XgXGbQVyNk/nCRgURf2Yf+nxHvkEE
+vPYWGZAkOhsxfuWKIQJiGUckVJAF5Z9YZ2XZ/bTIGgwR8QpGdAOVYvKZOIJH8MS
pDhuep23OOuZa/XltuSldYJrLf1miCgK1NYui2rp9JtTR4iFlEwdmxwXMmLH5+9C
UbUegsZCem9sAN/UBYu4uhDK+ve3u5UqoAJGrTW+LWBOIOUkd+pUglPwq6tisWlI
oTzq2CjXThQ8o28cBTKRPqE4aH0N7m4IEMUIOijb4WiB4R8h/VCdmaFGKF19imPg
5wMekCnS2qGVyS4/Xw2qyXWAvsQhmOJRfo4HO0nf10+Cc2zyBkIeRlRuxjwqnXzL
eMqVaiER5CMS+S4ZIyMgOfowp5UGe5dWJIXQOFNMFux1SFEYWEwK2az8A/qwwes/
H834BAujuIVHHrSiJqpLA2et3xHjmaVvDdwIXbsiH3zkbnqlzrs3xRJctS1UvbrP
RU6gIbcJP0py+XQfWx37iaUEnFbdLzupSjD8nuxZmciVeOG25xzW81fqiV22WaiB
sqbR2wAbEJ3io6oZlwlCXqBOvvSooL64OsKExEnwidGcbOI59mcamct+g+6zD4Cb
wUuTm5/a2lMkXa4IIEpdMZKw/m2bz/1EIpbAGRARe+ZB5fG9x9yWi+ZFlRsQ6rLd
jmDXBnUVNHV1fpOschXFKpQkIs13v5q+mOewJN7DUw4TFAsxYXfrPUEmhtbrPWfk
ADWxz07bQRlin2btOoKvI2WG8O+RIATUoT+UT7Dv9F9FafBOSk04N4gnx/eDn+pO
zjObyTJGOq38nv7pPpgLSdjBFz9ulZobYPTsebnWWO7nQ29BFDn/v5Wg8ah1WPgw
tHTQ063CjhwmmNzBDstvKgCD0R9D+3mvaq+5JoNhzldKmSCvTxYXfDcbZM6S4bg6
busbL8vnBmHqaMWGTsv+ZMnzYhUhaYUbhS+P5o0W6PLYZOlLWMtlJS3VFShbltpe
rwevJcl2dJz+rzKDia1WEkv27RrZSFAwoHxNGUdU6h4TyEwKXxVZ0ftdnFJfNhPP
6sSqaCHRs9GzijouTB9cfZFillMFLALRzUQZ3meV3bszoSqpM0OSv+6W4cqVyFda
qbTocAIXJkoGlxLCUe6u5l+BhNG0HteQz0J9loJY2LfNpJoKi6EuL7gxW+bwblHD
sQC4/RCJOz+jBbNFq30TEWRfUhquFfy+l3vGnbH7cUejEIhh9QUY3OA+6UXAqndR
Y38VHV9eJ1mVzZPImetffnk492UZO23xkMUmHQQD+JtjN+aeesV8jASwJmZxOfCy
kwrsNwzfJd+A3T8xGaYDG6cFVvAs0jAmdfmMnSJSCtKSGJu7JCRlsfohr9wKXVla
BG0TbZYaUk7MUdR1iTMLV0WiNBtvLipMTEjx6ZCilKWnYCveW3dD1TOoSIWi7MVF
JHznrlno/sOF4jYGtTwH6rgtAHH7BFy9MoUpmhvk4Gu39l5F1fwh4T7yk+CzwSye
xNFG3JWPP4RYI/1E6B1bCkiqcRVhgUIFe52qWnFPfyhQGJM+l4QwBim0JizHC57o
qNCJ0219ayA25IPgx4Qd0NPLSowCi/4OD+QOUI8yOj06qNTw/XhTjJIGOC6A6Q0B
fmdzItr0FU+pYCHBRWrSIBlualL4xpY1Z2XUC3oOMfijeh5DKIERtff4E2zIMr3I
upyn+X+ItVVv/eeonWPI02i9Xkmjav5ufw6cLtPfDy+iVf4A+BgMjqDXLamGdaMm
69RygZWgfnppOjb6Tk+FPgXrz7LpQ5d4+7njRN4RMELhK5eWoWPZA4UIOkMPH+Si
jLK7IU36YoCv8AARKzCv7DTQhD/2qSd/H1LbBW3SDI/QYwnCeZ5h9H7+2arSsRCH
n7BJwB6Ytyhtdhr0u++1/R9t6V8sdi3K6HOJqhr68x97CYsWBnLrc4mK008WHARY
sk3zXApgBQg5hKaM7QJlDCyolJY7Jqe2IOdh0yELCrpo1paNAc3sznxgo+Qpx4A3
dfsvY5Rm3v6FTf2ora0hQDb/cVXEYVLx5W8E9N57iYdH6ZQr/58pI2nTBcNhpZ2s
t+XHKOYcDa1cvL/B32ZPRFXC5kmmMVxwjEAaivHvKnqJPQ5ciSkArnBDOsQwhU6K
6XmJeJRkPtAlEodAuuG6DMOzJjY+dCRubwp9XWnRcK6we9z8j/5waaIEbHcCrZoi
NipMN25gcM7hCkoz5OLnQTQvsGS+ew8OmYidx5hGWHoeOe4hvzPIjnn7syCYcHwE
hQFk5fixTmzTDD4yX2+JkpcrOn9x4edMZpNEgVO3wVw4XI1N6opOETKdxk+f7rvi
SCqwD98eLsefAhrrvR32dtJg0H9Fg0sHaB/TvkMeOXutK6q3uKgaU4/R9eoPlBCP
41hBNptEVbdB0+oUDPPMbY3VX9RX+aun7FeFMYVWz6UdlNOCoDpuNAI0Q7oBSp/2
C8Mqjy1EOn2v/R66+hMmPaJmjF7SoPh1/IyrFweO+wf3tGsffv8o+F2viYiax79d
KJ+itnj2U0F/1CY37usd+kh2c9b3vT8EmH65lMUooQ3Hp6NRlRWiDbz3Ajk3zVns
tyVK29Rqq/G93/OnM+M1tupJvfgNDI5Rsa7/lb93KukF/O67S0esrEuu5dK/4uej
RqOGUQqfRtWULxcsgU2Bs2nfBsdgQwvBLOhQvg11tztixLz/19MNXkzP8HFQljuH
jnvKWYVFjj43Fpzx78aYgRVOzhQHoTjzZ0lFWRCIF7G/umzoaZHhlS5VpPTGG3Sy
Ijvags8j6P5PCpRbnrY7t749iizh9QO9JZvJdv6RyAzSvgmy+sB+SJcMkkWhEU3y
ZIJjtfuf1wwawxJRCBVEC9J0kn8IKEwuvjnXeWC2MU+icfAIxM0sgXMj+uEBcpOR
BSFabjLtvKicMCIiXNIHqFyI+LJCJHAMnpGgal8ciXlPbWGrgZ9BCgcTYD1SWoJ7
vElBvRVH258iae0lqUjHMK3jwD3TeXUr1x2VYxmsss2djV3a+OYDtMky0J2JlxmS
wUHKA0P8cxdoI4u1OzvC6WdP7nwiD7CH+XB487EmnHIk9XhvsM/yCqtL4kMGKN7B
pyZDPMaprpy3FbFT8mGke23eGRp+iRGQJlWxU67rvoXpuQ++565TYx6/YT7e5hs4
cpZluS2Th6FmMRm6MPLKKqTfHrU54Wg+l5qoPQ+gAEooKCsShuwG0kjk/1OSVrNG
+KZBcPtKKicyGPdJ96lVuD54n886hfwyFd8oWlut3S71EFMT7PZRrvFwXWSbaOc4
Zb+RHxhALGrBD37IcSzABDz1TqxLpj+fvgeUEz4GPFYKly4MZDGWnQXpJVNGZZGl
jXOpu1aJxBh/yyWbZ2/ZAYYu2F6psegi6uwolNn9TcLLlUPwdxt3alVSB57Ba726
eb7x2//G4jvHv4FEYEbiRnAgYkmdcncI2weHHQ2tM7v400q6ndV3XidG0E/jw9l+
CzQ3E/1Mwzzv4VmycgRQk9sGo0IzCsRIhFBe3Tn2kHriXkcz05pnFAeVOkIR0vuB
gvRXtg41Rg3qNun1Z4e2jZriUwAt3okDUnTn5iZ1N2WK16YCvMF0JHQ+nnRR1Xer
SumPcM+wdYqRQf5yjI3rFSbj9zj8tvduVmBSYOKSy4ZRiURqPe/9NxeTwpo2rTW1
cdvVMx5YLU4PaQlpkuhRD97XA2Cv+LNfJHAoJu+wc0Z9gY63WOyNT6WaYG3TLXbV
0MEHt80Y+evZ1zhTP3zIxEF8d8dsvAVdoIc8Yc53keTd5lCJV+o1uIkvfYg3X1QE
4kAjLLGvf0syMWTCgglRlePf0L8F7YYTwJRNPWwQfiZXsiGBhxLRRZu0DzzOlZgE
rF8RjdtHLHr1FvnM8L9Jm3Gbf9cjd3V5eGNKWMmOk78uWhDP5cy1S8P96AnYELJi
+Bi42Ot3p/YcrUHej9W4GNnH/G4ZQ2CRWyM4I3qNxaMh5kZqYAfXZf9elpFlyu6b
TDirw8r4RjTRcHc5BdbupPKWHBFMbtCDCIIDAsw0n+eBkOq3aI5z1B+Vgp3ZBb5c
2bHjWD4+h4/sziCEp4Whug9y//WfwJj4tb+M1ardrPYyp9BxNGVs/iPtYnGsSjcB
6vq6iiipP4An6alRaLlVj78gLtp35v4hWE2dNrcbrYxyHL5NUrK9c0Yu39oE4Ves
87WfeUeloRTY2SqpP714YUvp9kk9po0SYyKdidOVvX2s0Eoxynn9cnuE5vTYm6mW
Hb9PhSubehH3xCWZa9eNZFcZhXa5sx4k4pHK2K358Ecfi+oqpXfpm7fH8+KLVgig
H+6B/0uAUR9w5awRYjAtCvWyTUT7MkMSn9oEkGRa4fI4PnFQ4lt5TAZAgDGDJcNs
4f7Kcub3YipTM2abx7GVNhJARAEHUcS0dDRLPUnuTX1iHNJ2Ek5SOTLn8QAo7Tfb
2djKpE/nGseA3cEercWxtd5FFDeV3f/3I/OWDr19eYI7rfk6utdULysqttKfGyg0
pkeWd9Q93wxiHIWesF7HURDo7IY4aJBM9vitu/osY7FD+Tp7Hl8Q1RQS9p/rLOK6
1vHxkIGyXeS29A20I0yfuPc/1x6V0LNfldPKEEiu0NYqH56Jmf03X4GFERFhBlKU
0QTet1eUzbI4J1XjHw/uxa7jx+9oAcC2XHk7dEq1zWT0JPXPOxJPy2up0CNc44fl
q2G8Kik/ieeaJKo3XurXEVLdbi0X/B/HjCsGaF6iHFzmlxpniRY9yMCJyOTwOZMr
DgeRnMKht7yNvs9aRtcC5vTcl5Pa5GMvrl2ryQEEpD5MuS4KO/cqGxgjSSeCOCvw
LxUtAcQ7qXj5CljjDpIBtABuiLWZPcQUwqhLWnnamgk+/q9tJmifb62Gtv5EAKWA
Lc25yQ2i6CKM0BhkVPFbaeYJUoB5Z3CGtSsOXXr0chmzyW/npGZ6n6ht3XafEnF2
Q9jOnfthw58i8J6/fhuVNSU84flZP74qkP/TVmMFpMCHCSK8cLRPq98bF7zGvJxP
T0eifOVYnh3NjiWWzhRlFjbkefQie+GD6PLICtZkeuIbZKdRGh6G2cGZC/cgc1tF
Uugp54/xCJSXIT70ClZBD0RrUlrkP1OCBwpmnFBBHD34PIg5p47Pw3W2fSVPh6v8
rvn9AwjV5IVs9CrxsPd9oWlXy/uxLTgaSDmyo+DTe83FgrX6/A+7ay/AufSGza7J
rWNiX68EqWQ39WKTY2Ct15mRpydkBvCra0GqHjx/aIcsL8e2XSziEacrFQ0N5qBr
dCWBlzxG3xhNFLXcQ1Z35sMJqhgmuMGZ5JmU1i/gxlUnL8OkuYCoxd/zSGo2vqtI
i3iiXIvuzftGYltcf/W9QgdbAPQDbpm7v/luvrqVUVCwTUZqxDyU1RWfK+bEDy7J
Jpzmb+jTfnZZRjKOauuG99jdPtJd/GSeqM5EUgPvKLoVLdm8+hwkmhJ/1Swxb0ud
OoqvzU/p7cNPLxmMowVQjTubQroKW/ecAwQTWy0NCCgYMoSl3I6lQQCsI1efVBwK
5JiAo7CnxBQyXPRhxdKb09Yfqvml28WA9pKBUjGhEuzL5GYkIFK3+vq/l74AKi0B
pugMaheMEoqn15bd2rpQ9wJgjJypOSywTMuEY03x4b0LjA8wEDfrrNoEYHxy0eFY
Kq26NDP4P38qxnlbKwZgvq9I/ERcCGNzXXEMgEwMTToIoWpNee6Y3erIB1gWKTUb
OBKz0AFyhFJjtXT4Fzx7zixFUA/iOdKnBCpynnz8NIlYrgShFgP8Kme3xpo5HEVZ
NZV/pMZbLXXj7Nr9LtXqzp8T4teZHYcDGvkeTY7cY4rxjxLU0NXKeaf5GrbATrTZ
wTEYyaByfWXhBNBOXCKA/TUSu3/G2+sEbq33Ejiqz3Fs04Y0cvVnIMFZC+x6EM4r
PVSjc+2/pu4z/f4fDqY01MDJUj6ZwTxYWyxDK9QgG5vf56W3U4ROO2Qo1M1zrf99
D6P+Mtb4mLgcJ/PQdhJoFY8Q82y+8TVVY/KW6POfZo+ww6bCtYWGPxwzcxyoVrfM
xfRnd1Nm1HZmIpoW42d48qs2h2o4/k54OCyy5mExJn58p/Z3qkBtrczhdRTHVM1g
GXIBttFdIs4Prq0ro4bY967hKYe/4ZdWXf8xdEPOQuycPcz4G3q+kYi9RrY5YQYp
HvjD40QJSS97Pe+E/zpGkjldJdEr8czhLzcqk5Cj34rbKGvZN1nR8L8FpUAO1j5+
RNZoE7BnGgUPAuYqt1lCZRyB7dvq8A1SLO2NL7RaeQBDzxdbvS7LRS8FVv8BZf60
OnIc6fP84m5FuxfZfkQgtP1jr6BWCPFKtYfUIR9TpFlt+Cfzrns1EIAkdvw+pZCU
emVFBnKEGmX91E5MsDepfWazmIt2f6GH3nxikkwlCguaSl2FIDRy87VuQyESl4r2
8APym+1Q0nlOg0JUfv6Gf9DH++5RgOcapvNG46T+IlSzHeOMJ+BIpjYuF1AudMB1
iONxLKSxdSzN4ZhsgZGpUKwep3hFSJgwrUU/kT1kyTtrlnTvBgU7T/h0gpJotQwz
YAUHjHMUW4H0MeO4NNANLq6kHKOEacBYVJBwbEtBOZENGvTMsJ1yi5Q27/ooJRiH
HP7lKBulfs7LtQUoKosAq3ZI3CnVKiAtb/0c7Z+11l5CrvMQWyuMVlhzzfGV9hAy
ToYkCtrsKy/yG3lQCDgJsHWuUhPJLE3P0n9NRsMtZoBH6jTdefzGmTChpWWtLGKw
I/bYMbvVHRdHmhtVV1KFPr5qlb5AZNmP4QcpXcJz8o/se6T6XitVPUiYG7KCOBpS
JuNBSKHIjysSLE+wdWrhLdBT5U/iK0wM8QanO3B0IzqfOeCb7Mug688pZyTe1+Z1
iKV2dix47j05MTNrTgLSp6/akoeClmyzVMpXWJBd2I213eWWLoismTqKar9DgK0Y
1tTUFaOIdyWirgB+Qj+33Vz2Af1/X+N0aaGT+4NldKAQLgEr0QWvn76xgrWDEgsH
5+6VEkgADKiknF4HleNvzfk1x2x9ZxBfBroWFOtQ3Sv8IdMWOYC729OTbSlEbEsa
CO4Sky2UwwdKsD8rNT11SOnJQOP3ST62fm/7cvRduieCIA2I/s6/n7OohYLgw3Wi
w5EPzZZEL7b12MMqqCL8JlXdfwyCa255hCfyRj24TrhKmZ5Wi1ChAgOZewEXezL3
SA3jPcq97EjkO1B3YCOP+kWW6nemGyRTWwH9BBPfroOPA17T+oIcZILi6V9RX5iS
2HVcwpYSajOtafAnO+48SAO1DMCdRkyBRLoFAUpYVgAYp37pnsvNnH1m2W5W4OcA
FgAt1EE31adkyJO73ZIaAlG94BZPoR9sdulVBPX3LbU0V5y4fDTYDO1QxFwScq3t
QU9LqxQ5cqBpCivYlgAT7RXlhE5Uw9eRVHsYZwziIt0ioMVPyFtbQBhvJi0Ao+N8
83An3qidncGtyNrs7zB0ltWHKSR9Tn2fcw6A+wjpYpIc6FGdglSxkIrT0aAu8jcQ
+OUnTWIh3tW5iU5daynJm6H5chUbIyENWuwvNA7Nkwy2n3wXoeLDv+LeblHYlHyn
AJqtY/VKyAycg79mkhOYgLy2Quguo3FaIsfmjVmI05lTz1cZzN1KLlI77amGMbBW
l+fvyceGmrXusi2IlpN5NmR6cjxl0GTpOKSu2m94rG5uyFMVrqw+vqTG+basHv8+
twbOxH+3VR9WE0uCLXl/EqsSNKutAq460BzsR8zG77xjW3edBpbf8Ljp1M+RwjAI
iGhQo77syfcx5LDKhFhy7NTSG3rHm2SAG20FRWGFuxfJrXSeQSrtH4sUgjxhF5Z5
+FXhduYU8DqqBOo2sICGjOVC28hvdebqs5veBxJPqYeNQYzjYxE63q0Yzxcnk6YS
MCN/A6t8mki4FYRvGJVRQhXObCWk1M/ooDhsuW/FEM7JDBidu399GaJKNMTMzkuh
3wQVCjCZbBQNMSgTSCt3JaRUHyls8YKKCw0WmJukwQv+GCDyqrc+tGJdiWRlyJoP
Qwq9jPXojUb3FWgCfA9tv6/vBawhWyvo9PKD0UmPMXmu4Jki8eV62HfuLPd9muVU
tgyeVueZG2T5xoElVxj6P0zjou7Tf0T1t1dgq/T2QGacq8mzhhqxLuJXJ9+C4cnD
15/h0GKT9M1DIbLRoIkCH7/LDDYrt8S982SuW5uCKSdmwaZHVbCOVkk9HsXsyuP6
/iSnuHwrvbZknWGvHY80eOELnIRpfLXB6fdDR+EjpIqTmFPwnipciwCGlRAFV/3T
HKeB3UcyqFklwdeGI3jCeFz0tS0PPQPCabfpHdmoPwB8A/hnRaSevoufKpo7DVWl
Et1ZtBCjyuUbHr0pRioExLtIN8HylmUh3Z5wvjjM/iaBqW1JRv2uwmqAABmFtUJl
fV5RNcQ9UD5Qf8zny5Nn3njzpsSIWudkkg5BEM1a9QsnasmW4cFVjMLXS0tjfV3s
nGEEMhAunF27YHHFsQSgM9eRm6AoxhMjx5+8JyEP4OTNod+oogP1Wa3Q/wSJjj1C
4UyuwJxTh8HIzZWVJ62es5TyEEz95JUjvI1ZsMN7R6Uqe5qveT+3t+k9MEqbJi+R
ByG+DBoFJ/hewE4dCkPCV+S5pOLB2dI8/Vk9fAbJhdB9Au488EO10j4ZCa86nEds
IIH48u75QPPFu9vHFqQbW0t88hjQ/Nzoeyc6ZLibJpLsRjHoJPBx1RJVYQHb0qKU
I4yfWmrm/P7BPJ490t+hd/g6HmzA+zASW345sYF1m5TnBnzoDTMgvd6tSGjgnIuH
IC/J5yU0eejo+Zf0zOziCNSAa7ZBeDKtPz96nPsUhYIJwEmBBBg2vm5oWcmnfoUO
ce5vv5GmyojQ3qcf1cVi+IMLemhKWMJeHNyi94VP8SIXvOiwoJE/gsf6TNhOhhTT
LoTkuWhSeSh2zhTEw5AWTVRhIrGT3bKqT5g59Xz3U2Y6ITllAyvAndp4zMBI5gW9
5k3HWVjQHkQ+U4yXz25nS4PVkHuAKsEt2fymk+NjYfStDff0XK9N9xT8R9Lc+L8p
Ww1Dqwy8/9SjLAAbRBQ97YbTTeYjogkAddSDqmeSnCbqh19Wn2ZI5g5JnX/dSgIa
kYNa6m1DD0MhXG2CpZAKifP8Lx5bFXjLSoEfloph8XrQd8YDc/rOQgBrrn4fNBLv
/qTM3gZh4qU/1eINXVpUZsGP4zNVu2giSQRGp7lXW1Bvj2HQNWKzVz9ZAl4pvsOy
vJQ2Z6vrE7rOMvwahlLTyZgxSJc6Esb+w/i91DF+S4g/TL4rF77zp1PXa3hpQ6CI
wvKfpx23AxYqEVoLJpCAQoJWo9JAKkWbP+8f9woPoyE2F8Mt8p4TX95QyyQ1vzhp
1LqtYex6HbmtrxFfeAPrncgePwIObezUwSPtTmBCqYcqnY4oTNxufoa4+Xqi/jfE
2u2f+ErN53Z3isyJENIi1tMqMANFFw7qM3yeL/tVXJ+JHF339N5+rhTzuhDAxwQv
popWxtOVOyTAo5buEJHpdxVl2YZeXwI4qADeTCP9Q7FpBk0Xlvux55y1RIcChFQE
hhwKVrxaQXkuilk6doZydilu3O3EMmf21k83RvfqHXZa/lWjIip7jfLzqDyzLeRQ
6GR/Pm17xcMaD39Ndv7I0MXi+ZApE9Cqd7roko4AAWUXsLsieLuJG/9LWEbCgtGh
ZQe8kIrT9NHLIB/g/8oK2YS6y8xpHyB/dN+ZPx9i3NdMsXbmiT+9EUytfqK2GBSb
Q1SvQc3hd5YpfCrLk3ErEs4OynPpqtQM93+DJXPmitHxSDRcwk8Bb6dmg+NVYgsf
uHCOqfS5mnppAehwMXp1VmgONu00GiMOimvi6YCUfc8fkkGLsyK9fEUzg4PR8Y7d
vp2ByNY6ArrAub52fCZsqzmb4/GcZEEe+BMVJbSKZJ6JQac8abfDv8cIfs1NaSSV
2RYUjgu24UvhMXTBtMvf2j+te1roAR1SqbSTMIDdwLzfNyOeRruv7VVUUZ8Ia6aT
hQkD89UnCoZquD9MVEVs8G+DoX4AxKHoIrISI9KDfKFRtwmNp2MwEBl4T8b2vA6Q
fr4oufCAC3fSbKn0Q+jp9+qvofJ5HOeyyVHA7VVzOuEu9KJ6CQjMHwYm1xvnZCd2
XaOsKUs+1ZP5ePJymx1oNwynkzfXMcGxagI63OITrF1jQKvaTavZqh+EwJu0qAH9
haYe7kL/ixBOBEUh0YRdJKPFa5ipet3c06CIEKZ/lotxU71jD4fOFf/wfZ2e9Vmn
kGE5pTxj+JTinGmAxJ87T0+aAKTwsIeIdsV8vx37g8SFHFqnAYnucNlsNuhdI+0q
VXcAnwj3GKMXYmKm5l1VoScYKK4m5zFJBLUIgIYu6rT88LZAGyk8+B8ZYEXRXfKX
+iDEoRRrjWMI8GHnIP+ksC3A/bY0AkBSc8i6WDJwel3A3ETkqGA6bpJPErW6cksQ
PscIrkJaER45gJx9c0g5sEMfKWWz1QTLLg+rmGCIGiDhiRYRLREezeagQsQwdwl3
F8cEotEXLI9xLutgyaEGgG/PYrzCqBZnbQMiEEjpBJ6f+8svoz4Aks+pB495ShRZ
2NGo+Dpd1s1vh2A/3mtJyhyv5puhmRO+llhVyrcFjDoU3l52kh2TJoMfX049EtEQ
gyNY6w5CTq8n2Cw0rcrw5uySOH+faSg0X2eCIw3pV+0kyVzkURlh2plZELWQZBZx
CReLoEsSURcZx9Z0b+9mPHFE2cZN+gMdUN0hYMwjEM3mlnVoAELgLFMAopbIrwOf
MGcBuxKnQkmAf2ML6giQv0L5Lk/71guVNeVBTfzjZNqAQEONA2PRpRjCe9AkukyX
PBZ9/f+OII7m44Ror3S1bepCFTI0mPG/VmDBN8XGhrAQpCC9oCSiTkeG6D8L2Z2U
+4HS9I5OItaTgV58k3xeOJz7h3HfANgiJUcFzAeZmLVDjV3GB03JBDLFqLOonxf5
1oLdfBLbn04Mn3ByCCvN50R+ZSK8BfPBIo5JAudzeBdVMyF87MCFxyRoOxCDJRq9
5JQrhilQISLKr76aCdz2rmm0PIqm+FBez0a832mH1d/clqM5LXiBlAWkNGDR3HEQ
F49JjQdRP4YdnkLIvjqNy0bHur9sF1TJsuPtPpLlZhTpcfhhMyQWRCwIbwOGvviE
DmYYR9BB/Ak6iN9S/zgCVX+dCC88nT0uFYSBkwkygS1O5/+68ttZwvjWbe/zQhuc
4hdQgeb6/HpUq8P2qKJdFdQFArsPKNuyJbE1tmdhOHCdMihgjJKjPsvWy8KqDTEj
kMoiU3cmzpoLjOmx525ppBosWewHtqQ7ZsZKFMVj3v1/Vqi/gxxv/qw+oBrsoz9C
ymFsirw+pzmnCFZ6u0+69Smd6In+C8WJBqYGgpMIWkhp1HtiNPfDOPq11h8i8w8l
evtWtUR/1MLnxD2VluSo4/2kaHbaP9Y/m3VqVCioqpxpSiRUtXsKQSGwp1R05A2T
Ls1kZjDbXwbDmA9i7nV8jNweaHL6B35PPUNzKtoZ5cjHKkurnoJH0mTSKw8JwutX
nKFwHD3Wios5alGCf+wrBa3Ll4NoPUqF5eoqChyPEtQzF2MTIzLOd/RQE3oe0Z52
30v9+B0nd5Ce5t0+7Ba/lNGxvjUzuIOgzgm2ZY6Fe+1E2HI4Q7QhvDMLeN7aRasX
/UPeMVEuXpINaD8DgvnnQ45sTJZkBKOlRDPfF6XYros8m/hFxRNXyKgVVnMf9N1J
8ia3UjBa/XjHvZ7HnxTeh32rX1eSrO4+vlQa9DwyIgJZCGI95jCrrTbsF7p5xpV1
mMZLRf3x/Cj4MaIKNneb1exK8DxbQ4u3Fqpk+mm21bqM6glbzQZyngXb7vRXFybI
YR7u08Ohx5eoIe3iDBTGm4MA8fvGcG2+GTbjMKFLCelJOp5b6qKwPkPXz9iHC2G1
rr0xCy4RuT8WIS17xxPxaeis5/gj86guX+RFGa7cZyFuEnIL3/Vzl7yDLENKHLld
IaJT26e2LsUs3c7LmtGXBXwfkJMWaxjgElovvKVNcpiUtjx6jYtFQl5XsGbcXKUT
5ZnwP3BJifsmu8zU9DtXMiucEnBW90OFoKdiuzbozuUOy219WgCOtqnVQAlif7Mc
xcZ6GeBETXbbzFvW4Sn5TwEdRulwCta8M9oom2r2MiU6TNHBdWeLct6Rqsy7WTFp
Va/aXUaq23bxH8VUrSvyx415ToTbgIWhzFIZumWthtIvqN4hayv43YlLPxmt10hC
Q4q/O1qb1SntW6hpl6eDKHSq4wzYhUhRD8TT+eaGrHssHQuI/Fn0aSqmRJQiAa/t
6dXlNv3UikGsCvKIbU0l5lKD8Ifm5/yyMkEjLsz9caScAQYveHEFjWnZ73/7ELyQ
/76dRtxZy6rgdAY9VwajTgxYn2Ff9+PyUaBEIrOekJvWGWPvHoP923WnLgEIJ3Sl
5jH1BN7RIFHtCve4jJzTk/del9Bhq/VeWRWYpkMik4CHr+uLdRn65FtRqTEQX4mD
A5M7FMwcNuKTWORcQG7VrQ8/TakSTlQfDua1kjzjanFGu75lx4+6fwHkU/1O5MNW
q0gAspPQ7Ndy6WXndfKmC1THMD9Ku/4bL/hoP9LgD0XeqzUiyWpSGTvnrqehMPA6
pNQLkHLo+2j0utfCZcLZzLNoNZiEwNN6uhtw+jZxUWePYiHUWTIcKTL0i/NbbZLe
M3cS89p/KSWXmrJoxb55GkMyp2VWD+S9Z9j9pUXO99gJyR0kPRnHDKYoN5tfe34N
bVwRZpDfIEcXqxxtcEEY6oAgNu6Jst+6j/XQ8M6q+Co7lrO5ZjJdhTt0PUlOhboG
ylQHV0a8cAw6D2lxQz7B88hxxpJ5sULH61H40byLTSY+nLejTHPJbGFvie6eU/7n
sOGaFMdyekcRWWLziXdVGqOMbcwbPSaVfELMAzPbavXhW4oC8Dz9QZrCufT1BZg0
TGcelaAMdjNqHNiqsr1Xs89X1EoRgMR8jDFYf6+vLgy9SJJKcu/KnA2W5jE6bLKN
oKQGP7CzdUao+h0u6bpmh+w2IDs3XgX6tIowEeyQ1fstOpo50VkgaIe76z1njFXe
R/bM/1guXiTNYWXU2vRYYdV/Gpm90ntkkeF3w6NZb49a7ME9pKDQQyovaekuwNQX
Ll7N811AeOJX0bh0Wx7fGxyQAw1M+1AhdQjoRj6lX/uo4FZUyDzuRpaRVVUjgFz5
y/4i6q9UemWueIpzxDy5uRPbLCYYUNuYC9Z1OPj6sCtCFuPaBkTVM0Pf9kF53fUf
GxjUxfrraa53JTJcNMkBd/fGSXctKLg7AHZLye5htzZzjCWcRBv6L/l9m5m02Gkg
tlqlQ3+uzqVDnPDdNxvM4aveuEn7PE9+XImTbgGwLf4TkYDwDk6fQwNMCwVXm87p
MoWHNz8SQGDzA9JOV+RIqkp/wA/ku+dqzjYpR2WQlLirzljMxojyD1KIgTqgxtJ4
l/1LsSQwRhGhVum0fiIuthS0PbNJt0+4uo12ozko6moDFkSarGKxwRxyWWPCSMLo
caVwV4WQ18fZ+wy8WPXZjxbO9tdKFZ78v3Wwp5dYCwqSEnL1xpWF4okK0CaUbS5k
+iZYuWWEhxCetGP5hviloc59hYlxoe7r4MgJOWvbuka8WYNUW0HuF1x9NKjSakLc
F3LPvCCwFlXU4CPq4uJ56as0OdfvDH16riGBRwuzumtaeG/AZn+InY9MnnqcNPpW
LmTDMzDKuo1RkHB1TtzW54Qz4Tv3qDRACQkKKLUweLsUDuNpUjp69Dcu6FUuXSty
DJLlbKcYLW8APUDOoObEknl6zd+G725rKRoZrmHXHJCX1GYi2Zw5t16T8RMdgtnG
43BEnsifL+agnVlSmxwRCvGTLu1FzqdeaP13NC8RwDq11gk2BwzYUQpbfzBOuL33
otEpjW9BGSV2veAZ4hZT133lJU2lsKbs+DDjJK/AdIiYWtbwfnOjoLoAJHtZb0wu
vh5lmcYG8ZEw60VGtK3KZg58mzk9ThLZm6rPm9hsEGxUiWPXdvmFPsGZbPB5WpAm
TpvKTMLnBGD+UFsQTNQiKgderIH1uq96yeSYF07XlEtQHQjFiveS33l2a0iOSY7l
ieJzCkPcsHSQLZOjXAXFpLdG6yn6+qcnmgLcj+SY4LPJltWk44u84VXqxI4OCYmq
Nruhud6UuAsO7rZkvhYgGy4CCllsesFBrd3qUztg339VM+Or4F2RyXq4qloNJAPp
IOBAyTi+6j77VxVvCpSf64W/8f3/kQnwuA201dpP0kstc7/bTzfzRGhcHv0ZTzjZ
DonhLc4ThdPzR2hXzBunDLbA8IGCwXOSMJGLSEoww7CiNgUAUYpIoyuDKFdN1xCl
EopCvVld1MutMyrfhyg3bmzBuWC/JFDGKOBinPB/z5fJLZDDjx29zG+t0bAMXKEv
Vv/tmFoIz8dhNC7Nj4FLe84QSDSR6EWrplBTQK6A6lq+70mqYpAc2hAqeiGugybo
9tYXNwOGlJAq9sU/NeWCw7Sukuc5AeKhco300ZdPmB4Wtiq8vz3IKmafV4u7gh+K
sZEGb2bivmSoc5FO9+Zf+arbJi56r1W8JU0ZbYM80RR19K+BPSvkvprKinCyDSX4
o9zSvgq0gpTJ1FB386slTfPa9Y0bXs43WZbHDNoaKLCNQdVYHAA4P80msHU428LX
O76fWkKQm4dcHdEqqBPEVZV1G8Prp9pwCnp5brabPX4/InAq3D07ORWDMUkAu9Gt
PLwNQT88fI9SzncvUXv67WvuJ7evSCTEIFXJ25KeSklglpQHjS1ypykk9/XbsSc7
4V44SG3jytzUm+sr8L+itqJOk27ZTvpj+AxqOSLTrFQjE/HzREDshd7rdUB0I5Mv
qO6TXvMtObs+wLz/wVLeRq6lJNwhwbAEf5uYIbbEpz+IuqOxAKcJ0qDv56PwMkUx
pIta0oZGkTTb0O9zeQWAo8tJMgUuElRG3dnN2R6Z3+apI/oH0M8IQtMDmZr+cwJr
2SAtabbU6SOt1AU7KExsAM/emSx+8tpjBMAKm7ieUlt+CdRUlebU+rXL6utQaSOf
wjuuV7amECGIeJuxM5TdCYgtzC/KGf1c3nmAUqJlzUBVPWBQN7o6ijPa1RgAbuFc
Le5Tk7stl0b0YCG2wLnQKn9qtbxOWl4hVOS6a/MRMlRIDO+XVpFffQIL3eKLopee
NDT67L2rBm+9uXWgMm69Vi+9V5tk38sQRea/muTORi53SKWgJBUiZSDtfhGwOOFV
mpMxA0AJ4rdgSPeq3hilKFVDJ+oE1N7bpg2V5h+X6uXknBMq6LNXHPJVuF1cQlou
IKp8myLTUIkou1Nf4DQ0yeKRiR9+uDZJg4oOp+zwT6HVPB6PxS2OUMciqT5UM6kj
lNmONnpI7IN3sa0G6hYhsj10IXFdMA+nXm5KGTaMVW3pLreBqdZiMeuRpAyVKzTM
nqwzhsZEERzJvFn710F+LBrNji0EW4/sC1nUon/pE97iLo8Lzxhbk3KzYgHzZ0jh
FrURTI1EqNg/Cmv2eYN5OIufSCNAFYkNTWBPzCVu+mui44GYth/5Udj4C67+Z1Dk
znFri8GF0XZZKClxAadP+ScJadO/f9vIjx6vLp5bVNPzMNGpBwDJlV5mpctuHyhb
jZeOuoc9bMcqPDrYnlT5v2na4WVGszAPJ0maVUWDgKNyqofLvvLTym1HO5vCThVB
Y2QDOhH8huYw3jFsZwvTGh2NsGSIGcdu8QmV9Dnej4q+AouLtTsRYikNnT/xuPpD
m/s/lq8n2rHdFINcnkJYWBJrvzPCu8GEL0nNLSs6yuhTlDzk1pk1iFKVrGt8vm6L
cEYbRF+sv543lqT2DlInueML+zFqIPGWA+VNyoQegaa3mDhCLPTuiWOUjP1dGle8
P1bo7tBdBV/UBi6bdukEvHg7T7dGUAg5xTEsfJna3ChNrwQks7mRFH6nqhJ/WFlJ
nEZ7MXrrABFHTzhkgIBakZTRwZL1+Xlzd/xNjtXj0RgCeEFchabhAjJolUXIhWOK
bnfCCTLQ+zWtCY4EAPIXA2RQdL0JjlHOkA268pjx+dIZnH7EfkOrHDwwg/tC+mgJ
AvxMMy1eB3BF/COm/xeLGlqpVYEtjaGP68jvYy0uiU0wDXNgldTIUhNYy7ETufIF
O9UpbJ+2fapY/iTrpdKxL+UsRfMSXjolsSAVkCWxc+UYKb9ThX7F1AiHFPoOiTWH
GnkzeTJq0wgvTuXpLFZOMXrZ4+ULnh81Gbb2Lyh55zyaK6J4sODwLiaC9N8CsU+p
36uwADD+9VtR14/fz8VDVNHUdcKzN9TZS8O1B1FZQmboHCBHyNhw8uCmwsR8vRIf
1FXOQlIj0P6Kf4X3ba5zwbY37VsR9y0JXbPyBz6twhu90G5MVFmXynbWsyJ03tJM
W+t8zgfKZsExeBZSHpj8YYf/V7fsNihtLnvLQXWEwMp9PgfazEZyKGep+9AWUVLs
IBn9mfmoqXNIpaGOp37H614iM7QngkX4rbuCZ9mMLqiRrtTOurX9GKPe7wIpcHr3
UvhVvgV5Qn5QYNVfmTfK9pkc4ci0NunJ8JeSiKHvuoaeI5uUSfCiV8QC3bT40u6+
f+Coqe/saN3i3WBSt4ji++aJ7sqAG667jCNf7+ojgpvsW3DfND9HSIoLuz637mLy
c39GY5D13EBqAKkCLIRGvJS6TaG7qfIxugvQVOF/2BHrA0/MoLo1nHTIjy0L9w/X
1ixlWHPJ5ExxH3iNKgb7p2gKOWkgZvYt363yvQmqErcKYzCr7jAZ6Y6LyIe0ZytC
cyKKiKUkYzm6HWR/GwWVKbwq3cHclU14uYg02iw8v1Kw5F2VoEN/aTsvj5YSJpPD
E8Y+0DGbhlavlnt3usyVioR+E/SRW1GhH10JJBw5Zk2H65fDeAuHqnIuKRcAOhKs
Qkdgq7vhTrctmLQYWxSYaFZoP6JiWvsrr0MgntLVGUPgui9564G5vKoc2/V7L7pT
kAelBgh11w3h6nKnF/VNZSHVitrfLhvg6DTQBd67KptaZMxTlRlzHsqCPH889pqd
5IYdHjt6pagfVXN4Bg2izyER22W5S0gNlpo3iKYRmwS+YFJq+P7Wgd9CPYyaqcDU
sNQEcN4fmDkknzj/jucXrM10wgNVzeOdc7eaO2xP00jNV8Uz3weFSLRinwz1JG7D
Kvne8wnasxJY5xu6VAL8KlEJjgi8zdsqC2VM4JzLCcUf/u0+MTxn7zGGZcZRk3JU
0Ia3dtGbAHpoW6XGb0OrCGi0A4e9MWRsycFCdZu/NkBJ9QC+YOBcUpo0/K0wvmMb
QLqIXrksQb+DcUHgrT33EH3W4w33apfFrmxgxFaKr/F4eeltlkFcstE1W0U6Nai2
qo0l1vnV4PcY2DhwLLbHPbddtOmW9Vg5d5dVobR307aQfe4imTteRXGUPi/khqyM
sZzCfyFSze2deLD3MG2cgMbX4nJjvQwQaWA1qriMyoTeJI/m7RCYN3EYAtQ4qKZY
b/XTtsI/KwCJKGmJsHzI1dw6hRzdbiOJvGWDeYNAlueYOnL8MQnrWWY60DmG2v7z
ZyonMrFN816l1AON2f77e2s6jPlVHV+h2gSgCk2usSwdBaShon/ujgHw3HRVWxLt
VyKMj4wfHi5lz5CpTKMgJgG4Z77MwqVOUmF/BgpbwtUwpCCD/GkRxUAf0k/K3jcV
IIi2WARKEWgxGZPlXY22aFFSCIclpyf3g9I+58a/2vvWclpD+jfeYrw/TR6TyyjP
za3FTAnGPtwwIX8h+R1PjXFaUaKLPofXlm0XLyFiiK/ior197YmcFGBfWbfCIQNm
bSnN3pzj0Ql6InJeqmNeQQZz9WAxLgYqgyytN0KSyZoy9sYBLek3EXYwAEu1ASq+
1MlnyGZUf11QOhaJaVmZ/cJ6mD9o68iI6d1oIeDy/iuTiKedXOokERk7WLZBjO1e
FznbJpOAR23C9ejVfk9ZSQS7gxrbrhK8ql74aFB72Gci9DHp261S+YTHelch8VXA
lfogEeNWtG/L0ZhrwxBOYWCafNKy5tjoVolA1PhPFU43wIbSyIz+6yERdTrUX9Ah
Y1xW7OesL9QENFdeL62b8rfgp19jD3HelQ2YajDtb5/xGMONJjlAtargu2wz/hS1
GOsmyqf548ork/Wat8snvyHuPwFx3qwG17T0sMVlDcC0u2uEjvcTo5YetxUO8Yd4
H93E8kLp3EP7yPlscU4oUD8+v2TpbvcwvIY/6dyOTtC2I8lkO18JvA7/xAP2nEoQ
LDmgHRjaaW2I4uuE54xIZxIUmlXIsrPEEja3yB8HYDww7Q4uQFPk0u6opj6g/cW7
ZEkjfVDUr7FisdJxQKyU/JAaRtugnCgF7d6NBDqTWBDeR7DhOhfT+0iQhMfv0QZI
/gSuOWfFxH8RpI3HeHi9dwtSOfaQK9iKijkTPxzzDAD2AqQTvdE4S4aciuoUUWQY
X76J0soF8ZdDBYN/E+lu/xlmswPOKr3aEZC8iTT3XptcRtufQlLOScybaBywOLp8
wmD09g81tePdatUi1UvUtcqPgBptibYMEWyy0xesmkX3DwBJUbekn8OXJR9mPOvH
PqOWgDNQLtRhQtPDcxTMvHmlB/9/5iJ5qerac4FtrHFnmxDBcIyZcXubdv/fOfNg
jmps/lSQneTbcWXr6XMrc9kKPuMaaR5DjDiZ+CPNI6ciHDUw2MhXEz6JNNq3H3A8
Y5G6xdGIWojpPDWo/AfZPdgbVaRXzokYfH7XnUePE+V5kqokAamv57STmfgbOLla
yI6i1vXioK3vwQcGlcpz7amu543zPyiw2aHhOpKfeUnD34+BXHNCOY8VKwm3UL48
cvAa6Fw4q/O/fQQdEsKHwebIoaS5dxG9ZYV5s0YT1Wv0aWEWNXf2tYb1dSLvd1Np
vgo2HPqgVxvaJE5Ttl6lcIe7/BFLgpe/cz0n6mddzSE3uLCOdAQbzXit6EbwBybr
HeFQfgJ1oSnf++KCTwXj6TCU6ihP4RfukjS8/YDAu5eo0JmwfvttqPO8OgIDDv+m
oq+jIB/HeZaqBTQk4/ExpSdhFUzqLHwe8jGmcIXELxkShjpSBvnD446NtPDTYWPh
xQcw0/NeK8Up60kpBumFq783GqvN/9HPW7IUumh4H1vpjJE3WJMSc32qYvL5+E9T
cimeAvnIHzykdcpFq0GhDkaTjPuFOXMkZZt1txiUDfAf41WT0YaOTz6OD8AWy+Y3
QKCInE2c1Wb/nDc9aWy2gpTFsYCYXHrRtQUD0f+VmAtZJauy5qVKimCgXjb4DUyM
FlVKplqlrOm2cTRYjADW+sPmDEYcfluZ4uv11cdr5vNjU3tQuj4DXw/MtT1pvMGi
Q+a6VVj8rXZCFGSt6vFVf1UXbuzNcep6SJPN8qWD/MOSFGDBaMg5g9p5ktX8Xamc
Q3vULfMjuDdgdMhMZBpwE8b+0VvfgwE6qMg663aPfK4DQzUJMxSvNQNUIcoU/Nh4
ykmwzbFagLNFkM4Yq2Uvliv0oKBG8/kBUYPn5SBUEtxFFaLmC7wDlnPuDJkDswW0
h807o869tg/8FiZ4U9GEQNsPXDI6WbCcKMtAvs7wRJN1mKSIQ3LZAh+YAzd1tfeO
vjbYRozAE9hDwBHmHNdk3j9Nf3z1ZXVpmVXa3uPa5duZXpYskK64NgyaqE4//7sq
9bpqSBkbX6pJDivJyPfLcX9MrwciXkLn35JiRIApYoyHzjwBNL9ReUmOAd0kfxyM
k0/epe2EnRNGNcSgCKhNNv0xsqV9nDyrPdZ8cQxCL63rL8N9So90bJ7WV6vGPhcS
kp9869jTHKn+PpPcuaCN9IbhXUvOZ+JFrYXq3/wSrq10sGimRWhNJZDAf44yIrX8
ZrBOkXfSXSrx7tqo2XR3bLfIi3vSxIuY75J9FDnNum86D0D0kQ6ad6SOwItepZxG
cvSiV3jiP9NvWLr3/erNyHNuTZdsbvVLjL2QsPqNikMJF51UZpabjWp193/DXOiH
tPFDYRK0O0QTQ1cLVZ+Ep14w5sWRGR9sHmkyhD9KhCOWdzuzU8Iwidn/9Uz2ujrd
KF67UAuSjSrYXIo54QeGeJd4jF/1fjx1I9Kc0eBboDYSFbsMtf/msRCD4lXdvd6p
9ZUSdaDgFA0E1tfQmo+Lx4TAvKXmq1ofuq8YA/6/xat3ybPGczqYpyGyDZ5+owsY
WvmUyS/60q4cl8XQbIeL+2N3TElJz3NwkGseLSfCKIpi7YHVfdcyUgNqkh5i6bLp
/cbPDI0wV5RTeWQe8EFGOFvUw54SeQshCLPOko0WOSn5+QCDCYH184AqdGR2hn1a
44cLNfVJn0wSpZ8hCw0dGRiGTz3UZUB3Rd4ZCTLqunca1se+9cmkwWrTkxRNsLPV
kWRYJQoC3yY3y7hU0l2b5GIcVEerpk32tPO6fTbuoPKWqm5F4dDT2gFzoUvxuKC9
J5Z8DsfWGhhz+RTjSIh0QlE4Em6DEkml9l7ktA4sF1m1Z5vyXeYXymylLf/AbLA/
g8YjGF9vW0CU61BDo7XEUdiyeEuMCbykWrevm5tEhXnlceXTzFxUddron+FCBmMr
nF6dk0KxsZfXTuT4/gevNoRVn+F+eRWDJEP/Qs5YlmGQhkwaPzFiNlU0Ku75oFza
9ENED1mAhezFckl06wI16NDcdJFldmA/vOakEGtR/SkknQvcx9FSWOj40/DZZdMX
LFRXEoagK7lpNDTSOpIYEOBPLRjf4oqIjFm0zirgOudtRkCcBrgJZVHKUgUNATKj
1MyHaIr6FNPAKzdNqxuIUJsfE12CROTfNXuNsE9HQECWsPFXOEXtNqTHF3fA72gt
dIEZeIzTmWnAhM6fLYZL8t4Og6AataLDA7exHW1Xu7SKe5KrT+Bjqrymxmh48qQq
vASlGAZ+vzyVaX9p7ArbGi7P9NI4E3QZOp63gRHx8/oyR9eVhMvB+OInzfoEFntR
pX3CQcq1boLmA4/+RtYhvAIB2G+zcC52DawcJDWMgQfuAf+KUhQQjF1kPok0/BvE
CXj/efkV2jpb6+ttP7L1Y/RDbJy/JS1cB9RaIqt4YT/KDQBwnpdKVmfdod55KuDt
01DLqV8YmsHpMY7eNTEZQodPF9zqll1ihpYRZvQBW7IzQMBsmmicVqt32V28PGQO
goNwTkNCUXUqKPYF/Wnt6hAPsc5OkkPGlJyaSdMyy7GZabo5Wu6cQCG+blYYAj7T
Cc08QxIeFWjN5GTbOVVkvMppfsqIFpOgn7F/Z5yppwoiIhs3Aau1VQj6mIIaXlgy
uhFRfJ4+xC3xBtNEuN8KLqfK5QpzlWyrRj5VHxtbmebii0O9CTuM2GM1z+xO1tsE
VYpEXc32uD7F9UxzE8vdhuEdzgSQ/cuG8MdnEkpjkvV00ixq0wUkjtTw3Rt+OqSx
HfKQyM5TuAdJ02CmoYFd5G51p5Q+EeTo6cEtIXM6LrLYAz3tIy/cU10wiXWefEhL
caNGU7jpwAqjvTDALfAV52O7zVkjpwgfuy+Kgq8bv/ETyIW7U0i+L98xF6gqbTMc
X3J22ce0f3ql7057cP5AGHAX9sP4loJng7mLKZBSp/DN2IQFf/mAbzRlAqAnYTFn
nTBxvj29v8I/Icbqp4a1kz6edEKm8QyccaVQEk7lHQke5dedaJEbsj3J8K9vE/u0
omu4OcP3D/2HmTYJf/nobuxR1/1sy6uUJ5p9VGO9bBdRofrIofB4dxwe9utFQdCp
lAX6pZL1K0gkEqbzgirUHzQbUxR4jv6IUYboDK1nnEQ1HMM9fL+xMGwsgd++2T2Y
X4vw4SB+slO54DsCZyu1XTI6C7wfqxmO+pZ/pvtpaK4pj5bkcPoAhUY76OYXri3F
rXNmjwIEydxDSdxxgMMcW3eDbXPbh4BV6E2RSVg39LdVKxSsylur4MJremZjYYRN
NkJH9CqzADAVR0CsQrz6FmQXUbCwHkOkue7aCAkAsAKaMHKtBnPPQh3U2MFoLCtm
9ckJGZ8VLF0NKMBSYjn4CdYz4UroJ4BQyNKuoeGCLU2xJ8mrr6sG4NfNsV4nPsrb
sl3+67G7DyPu2qm7X7aiq0x4oUogQEV8LeUp94Ky21MMv+sshN7Hprh0+3EGeOCz
RzuQ1RhnpNCsnknm81fLX9FPOGY7OWOciLuBC46v3Q+gGn3pN7Uomxyf4I2PDpur
If2aez+guKfbXnH+NSNpixdS1DQcw8b7iqbUkN4PWAb2irhck08l+f0JWCAcvKNl
f0dFAa0duXhcmFYczk/QsjJt9elNg+JN8aHwlaa72lryX8rjtxITmMMzPPcyY2sr
Zc1yfbPL89DkDZ4yUgdVl1oU4vt6Q7oRrD0bEo+MihyJyigcG6yQryk8RKIEsfFq
36yO8ugC+ELSzecxz9o1Dl8/aT53E+IsTyzdZGIQmj5OVeuegAd8ENNIyv5AWJpk
qhzAAP/fJyxkZAR8rwOc8GGPYCRUct4hUAEGhmiW2c5P5lg1pIDHBkcvsGQbkKvz
/xQ9qmFGxjhPuVbpyEXKD/T92i/il7jWfVwK9ldEXP3IseWY77lWHc19XqDyfcQ8
XRTdir3T6Cc2WzUfV6KwtV4X7v0mln37FbHbR9lCH6zL7HFzt6IPaadxK2OIRBkX
eIjox/k51WErDVgKSkaYCzTbNmsyu9P6BF2ViVbi2J53ttwOR5ObJ3jdUzZsl899
ygNTkT5pfBMjNTCS1n7cl6kSF8srniJgf4tMy2E6Ie9HsDc/zAnCo54qU1/mtt5Z
EKk6yemi8eE7795fwYKBx5r5mYVKdBe/50b52dBzG8hakfHMYdLSRO47bnIGB8Sd
11o25a97GNPbgBMZ4lvmbZ5fHGotBqNBgbrTAfdy+Xgzp6Yy6yCkeZA8CCQ0jRGr
Gag0UXfiLJqWAHIMqN0aAyNIl4q/PnTDsf00h46ibWhEDJh1B1If7v5SWiv3nGum
yy6ECJ+utYdYdVkQH65hs+d+UGBfdl8Jz9sgik5IBhvyEsnmusO61tTrIj5cTafl
62TE9RbLk3Q5yhxyC/ksUYzKDuGHMni5dQDzt4lg1SmLcnI4JmN7aHfBMUuZPBD7
NKvLCCYGO9S1/m0g38UOwrnOww08F23W5UwA4AR0FVlDcJoty7AElMkJNdu3qh0w
laAmzllusUiTD+sFIWrLORqkOE4p5uanusG/JaTekS83Kd6NZ0e7YhvAtwqGA4cb
p5SmPkT1NA749Xx2Fzh7yZwMlgfJvkFWFgKpcrWDzQIwhjMVSvGWOj4M69v/saD6
V3DbpzAR14J5Hzvlt7VU/c9rXcIlXDcT1VfFM9r0j9DKM5Kcs1x+uIiNzak/RQFw
dc3WVls8D6UbPUTzx0oE+8JSoEd1MM+yWpytX7pgnfKo0EbvMapZv5WK9zEa0cQU
FmAIFilBpmdX1TwiGBou+8rx425MTjXUMRaxQuC0XX+wQfS7GNDhj7aVxklSOfI8
orMiKdiauaA/pUuITVoJWdft2WEaUVWiRKJK6U5XQHqVFmBgh5WxOIzyPDQ5FVY1
WaEm1y4awY1HhBhPCBqyaNFBwRP1MlObHUr8QxTQRuI95WFLLYdykzOLxOihA1Aq
qlI85RoxZ7VqpZp31wfY1PYAdmr4QQ6xoIcTQbw6E0yb0r3pKszD6PVeutrojlg2
UfPAAygTg4dSCwYprLH2ZWgVwWAzHPQEf9Z6J396zB5biD4kCNnfy+rjkBtoXa3L
s8SeMENAr+oc9vMenwkKjl0BcIFijeI7r/PIGEiFBkg0C8hFs4BgMI+NFtDn0kMd
Ig1mpPgOqvMvODA9uhAkhuR5uEk1lMywFnO7tbPve0eUldQZb7tlIxLxnSh9hoy8
0nGs1OPH6RUTGDInBhiXvvqtrZxAzneUiK23UGlsFN4WGmdlLgRxSbyJaoWhY+rf
TeStV1xMCuMI2AkOPZDj2H712TZGBJEZxYuFo4+rTEqe2c56perc+UDqu1aZGmFF
jze5H0nO24XrKGjmGPdzMVDNVtOQe4DRx6foAQmPnzcQvTB6pIj/TICgKAWvuk1p
3rJlksBsjXqJzejAt20rEk5gQL4TPF76eUlp5ApqIfTIGb78Bb43GgE74AbBQAfM
8CmLTsgwZIEBm5ICX2fI/gxF2KzYbovMfPN1wicVGMyIwxv0WqF75ARQmT/qIt0u
AsSu9n9AgqSp/hKF1cb8Cq9tlDD9YL49V6OBFM2ey4LuX5ydfFnBiyTHC03e1Ufu
5uF7kC75mAXRjviR3DqISDmCujgVRV9nA9tQrp8DJmG3VQJL3CakjXm3er3zuQf6
o9V9Yn3ISiv0CfoOeUSEYRW//1ZnLoVA0Z4zPPtEHbA70G4OAs6eFFocFZ5TDvDl
PdN1olz0+643PQ9CU4eJTfFpa3kDmFRnVmq6lYKx31sdiV3Ij6HjMYaWJxR5jaTa
zzG9zeabNUDHodU10RVmcaBlLfXVkP0xHCoDvz9bV7y70UPWaQOYJi2gjEoqqONW
RWe4SKNTK1nsqWt3tOaTBTMRs8KAIrZ/+Pj9ornjF6sdBD2VaVIeJyiFX6S/AZ8E
N+JsjTZRxcMQs6VNNkYB0wxgnCJCaocT2uaN2mafITF3DC246FWslepj6K6BVk+m
RAUa75He1Fzy66i4fzzdeV4wj+8vxBvd1U2xEIm9km6vfD0xAAMQ3Q0J/G4CbM/5
gagPGYaq/RQvmxmWIX+lasPig35+gozQxEsN6iswMmVkT5zyIVhHX6Me4jDDeZkH
UWP6vwLwhCxWt6blF/DFH7/m6RuZF0SzcirsMGXwjVeslW5k0pJiujeGHLww6JGa
hM2ZzZTX0ZVSs/MrN1I2nnQN1wG9L4xIPzvx8O0SZvV0UDcDW3aF8TkwQRbFkfPC
LX48QjrDYcRQZgYZ1zMGucI6YXFvQHYk5k1yt5Wdrbmr3Hw4/UbMHjHMDzZlUQN8
HcXzp71FZ8leGO80QQnynN0RVMYDeQx37dXPnJq6b5jHFLz9vvf5BDA5abz5FvS3
o1QeNZJ82S7tyHUBoqaBPwFmVLKkkNCOZz4SZ2WRiT4B/WXnhFsMlxxHRYmnfkyD
6vNC0GY3M12WYtqoW4zMoyt96M4uxRRHXATql87qMNHz+hgfcu6sVFvfSecIpYP1
I4rTckrAiLdlzCUgggYy3zhIYhrT0d8u0NHOmH/b+kw+35X9Y0Uz+pOt5W4X+jwN
eifFLE5pzZQsgaXBqMW5YfmH/kVXfma/CC7KRXfGf2j3hYIg8NedR6F8rDJQftdy
sFjeNDOF69QrHfkOY2yEroZ2RSsZHYMduzc4ijYiI2JYk3628BgMA5P0MV5439oX
ph6FXM0Ce90hfDxn98O/R6GxsVhcpVTCn3e4BBbJzhJSRuQC3QNAv89qGjuQ/nr1
i9Fra1S76jBYM6ViO7tp3RSnWyZBrAiEFE4o7KPRH4CEU4n7AcNzN2HQU0TYVhs0
hWewSKs4fq8ig8hSMpdrSBsbsRIaWlz8Rb+oNZrI0ydh33NhL1t9Wjl+3nhsgN+s
ZHlEvS2b71Zw/pLYSxYSYfPGKbtbg7Np9757ViSVU7G1BYpkxeT530LKN1M/5+f0
XypNFXbhoK9DjndpuPP0Cjz0DPw79Oa4EyRL4/vJsN5RY+6uOLTuC0XCtsvKhdCr
NDtQiZjlWTEKAwWeLJELgmzKmLjX8hkcKI4H9rpMqIpFfeGXGoY6HN3U033EFXQ4
sjIGhE4MWi9y87d2O4+mMIIi5VcrIhHdLDs5TfmxVv2MB3Urz8GIVNB9bX1gEnbz
bsKcsG4bWTtjIKqzqbobJKdziXIE9c9I0J3XUcBFaJz9yMf+IukSwmHTJdEeimaq
zLTMiApo+lT+0tsF7QufjPlulaRleCu33FuQ8m/wBp2M8tuqCM8G/1Ypjg5laBDT
3Da7Fu1ito9PMZqtZ0LU0Qespa/r1kqDlzgUeroWbXYET1Ptc1fuBM6JKHMpm4hq
8KBj6Dv+2WWYWi5SEt7/6D5WgYHyXaU9lB67F6J5bjdJYNnS04fQOomE8TVHfJZD
hzoB6AYpluysCaRGhnF67dM4poYRaVVT1Lt4KXcfOj7OFHvRa/WmqYluOtpwchJb
AiQUDoEIzZIVznWux2YLa4wbpD1gVRPumR8A+icaWAHlstDgCvZ74NxeYI+cCRnp
0zISwb5LUETuIhiTJ3ExIPbG5vmH6OtXng1sS5cyY++EcOfG2RO+OAt3jEWr2hp7
yBn78i6RyWcwbQ0Fl09wqg0nBZ6siX1Iw+LvsJUM0TpO07qILXDmNT2xh7PW6r6S
3rQCrDYl7Wxt+9iFP6Cc3vIJf/uXL2ifV5l8b4YSUbWX6/oh0FP+ysnz4h2juDF8
VPw8pmi7m6EWc0F3bfNUW6qfxZqyLdYnU5V3NtQsS/tGROBt4hfiAu8RZIFFMi2H
drPB6OYz4FnEpTYmMc45mRp7sHMou/Uq4F8kglJdS23OIMvT4dKKue3ONwMvBKzc
9wgOl0u1hD8wdo9VCnHtF5oLJ7dd6hehTttGg0ayn3EhKqGymOBOh0OIbSTrzPWp
v20MJFSVolaNioIP12dsNk2SuqR/AQgMuWOYqs8qJP21Jg76aQfQl7/D9gITG9Tr
1CIWi0/SMJneCr8QeOKJQCTccG5qftYlW+egSu4qTQXeuTCkry0uy/Xk9ozgiKe3
1E2kTnjJd6837M7mmcWB17uXcGMewb9qsMDitRtYeWCdTQBVVP/UDkPmSBCXBEhS
UYS4Vyz/A9Ty0zMqEPVdujSEl2pss9YASyNJ1oH1FzqRRWqdxd9d7xXRrFH7i04N
C/Y2ufyC6Vg3zAw9bUHtUAT7bxfJ/C0E+sBFgnZpTESZ8YqwJ8t1oBCGCfFHZNxO
8uuY0NgcwPT46pN9KdzTspsK1wy1ruGA1K14FQB5Z9UxjG+F7ci9JswslfV3d4c9
vhzmambDICtJmdJhQbieGCBeRS3HTsE5p+MyPOxmDbcv7imPntBAFWljUqP2GQRw
8QQz67vnXGCGuiQ90TBWQFVzTFdQXcR/kP7l6VGg6sxyPxmAZHcy6BI8DhtCkvop
EOynGJJTEuX/lua9544C0Q9P51Xc8qujzfpg+VIjT/Oq5W/XAvPIkKP3RScB/0vB
p6IB2zNUo8sB467E67kDcM5CsdGWLE+Tn3PwE1B6RZqKf7rNsrZuuDlKy323f8KO
UuzOGqL7X468e14b9/8uMce0kJ16Pne74ZszgLG0K/XYN3XdkpiDvFVv0hUa9Dyp
RkuvEwT4GcPG+LNa+p00WyNnxhpVO0ve27XlYko6H5lHHie7blHx0ZRZKCsWp/8/
79/8nsZy1O2tDb0b9wI4TwKkxY76uNoEJIKhNZUWAOhM643NPpvk0Ghhmi6m9WuS
mr+IF0cJ+/6mt0Lr28AUb0q4TjUp2l8eIDHv7CiqV0z29yxK6+zFqyIFGM2dHS2h
I9quS7tgmLBA/4Db62Jl9B/J/86RLq8yQt5PZ1wPHsHxvFD5DCl5G5sYTHgp8tgQ
upZqagvkI7Yv5jBHwkX4HMRcudrC1IteErP15vOfF5EnmLhsF2pHvtZatY+j5PtV
jca2G7cKb6OxZi+c+zH8jqz8ptzlbYEB+E3hNe99/D/EgB7iB41Qln9M6uxOEZTV
10wjO3+pB2h/zUiuIc3doqoIbem6B7dSKULXd7/glPZsI1qep6R4ZkAhYB5vaLFG
A1YJQ5qdgGCKj2U8HoWynxxzqk3Oq1398W+ugli8vci3qhEcLeFtF/Qwc1rA4DN0
oYf+QlL0XeN9tyKHreZbrCBk+kIzyMPIEOw0FR4Jipmy0S3uU4RA9j4eMMTiwUgO
585PyJpoesZb46B1N093dAbgwzwAeQgiVI2MSAGgbykgcW13s04e9kWRM+EiO/hd
GmohBv+8eSDjHhwemfL3O2n58KryZ3rPTktSY1Ye42LrjF0jr44mPFddaSuOUFYW
BX0yQ53Qbk3ENM5LbnC//NUENkkqve1EljDbT7MXSRFFLfhzt9MIIBlkCTnT0hIo
ptY1ngTcQmZrlHWaI0Fj7qK3iodKbKE9DryMweuyplmBmZz1xyn4LqwuvuBsUqYv
MvZVupKwsohFWdFFVbmj2HzhXjJm+yLpx3KwAGi/h+2FwntLcZntdUwqIgR3SvDs
zzAfhgM9P/50ictE9C+KDbNQa35G7z/pzUFSahKtlcgqFKQtEMjcUL6xm2Y8z6Ng
uCF+QbjZc4theGLw7He/Cgc7SjTaAg7ZbO67QGtV971qDGllv4sQW5t5u5LHL+Gm
ieI/r5bD5QnuJ7JBM6ktLpIeUVwce9bkSntuknWJjPub8H6lXK3NHBqUYkP5v/a+
bad6Q40Nhyqb4KzMVdoakVe1Wbl07Nt9VKQRJ6bDyfVgfXaegj6kDrXQMO1NqGFd
CyY3Fcrn35bXRXFOwLIlKvKx4uy6P0a+1LYOd4vOrHHrE2ynEpL+75aaKmarnM7I
PiSJJQEt6POkxHnbcklOIEJpI1b7TwcFX8klHmRIPj9iyUcuFoADVF76yYIFRJQ8
O5CRTtpRPnfQzclO+f8/j++Vblnx3IYhskcjjK3p8I6zxgdHhQUQtmMZYqFiFLXI
DN0OTsogkANzy/Cw3pLHVuBIie36R0YbUx625ANTrmE+HFZc/GUCMm5Dt6ipDMjn
2n4qs8B3a99A+uCrRK4ywCTpDXhpHSVvC7TrFJkfDhhDbayNjfBBTUMtwI0p59kp
yoEbZ+mc9KJmPbQ15KXOps85LJyCtnqiBavQEfYEtlgWLhWyunuHQg7/g2FPbIDx
pL6Rs7vCzaN2pJoWeUqyWiMRrPSoH3r/muZ1371ACSaqAo2oEV0wA3vfT0ZX+gN/
CX17+xVXVDD8hs+cyB974xpYgbZ42bS6CmCB//aeix+uCdL5pYuPxUajMKhpOGfB
Y7C/i/cwmJc1cmhr6kIMMNHYHY2dQz/3MdOVOdtcxF2Ipkk1WFOGCNYvQVEJ0pAM
AFmRmeuuSVbkE5FrkAYBio/klhx258CtsLQkF8IsWaAWFjEtPiAecUua0mmv11ZD
XSn7Usxfq7rSsMxU01g3rr+gdweLUapvz9ASrI7SXf4Zwn6uSB62UgpBYHNdtWZ7
NIYjK3wgRvxKI+wSGoTwcMVoZiuIOBOV4U2qHNo5Nuil72wm/CWWdAOGgzk6e1ep
hR4WL7H6sBPnAlcn0ua8xvlnJ7BHcJwR8nRcqYJyk4uh8YkIR/ktVrHkiZsEuLaP
BKcSFRLUPC4iF5zDPIyhKiuvfrQtJIB5yTS2xur6k2cXny1W6dqkf7FR8iQRcoZ4
2yuFdM1p9Bea5TtKha4bUbaWDCeXL3JyvZkZy6fEuO9XznLVCbtIPhXl2OcjmvuK
ur7RAbuv9Z+isp5qOGAC9B/IiPBHOcrdmh61aDRZE9azhVUaGsFmKavgZNcW7LaE
o70Qn9Qf1+JMgRxf10zepR1exMNOAqA6umnBj04CXbhLll+OA887TI6kY3whV+RU
Bn/ioV7qfHqYKo/SXyNP8bh6jU6MgrCItOpLD/1XRIjg/ZgmABVsE8CJpCgeih7v
fMbpE0CGVVl+9PI8khGzFpE55zcbMjN8lU1MIc0rYTNW0I9WWUvTgTbeS0nJXxeD
hmqJtOsu/mFydPLlP+0cukr4j+ZJpoNwB8k4bYBUjKovQiKeBEar502qGEs2rsgL
gO5cldfRx3sytfN/os3q3Cxo0ExQ01Zbvk/+gDeUbdPnMFxjNat64Z/iP/RUQ1/C
+34plAjxsn54L8a0yGxCC9MPpFqtW9OOhx5hevS2BXftreJHGFTJnqPTvL7jm6nc
0vMs5LUZHlptmO1bxTcoxgRunS0tYU5fpVLBd52iX2yLlTz2aj0IH3zMFpgAoF0s
2E2rTbsEpjTmhccvF1hO857RHEtHhy7Gf8WvJtOWhUfdjS1FdYaT81Uc0TOZLIie
Us4ptCUyH4soNLz9OQxqstC7bNzGG5zBOUkG+MZijOsh8mkCBQlfagPrtWS+eIXB
t3z/DylVaAR7+ve89CnmJoyTsUbRs47GkBHl8h9EdY2A48KFzT1a10bviX86y7Uc
Utbse3i1Dk4HZysZfpGXDOzSOWxBEjYtzrb8ZQJV9jm2lwdmDlkU5uyY0pAOiEON
83E3/cjzVw3a3q2Bu3RHQ4WsMTQ3Pn0QPJrEJTesStR8H1DMn8alGALXEhhOPVqW
TxVVZTQQjAJBudwkGcnyyGeh1rtyMJ4HomdDFynplO+5q/x92WEjYtKIrypJeur2
gR6VxL6uK3WWW15sZda3fRVZj4Qdw84WrxoSnP9bOT3m3t7BP7ac1L3Oc6wgGYm/
UyeyjrL1n5XfdYbvIsuRMfn5b111Ks0Z+MPz2fN/c9Pg4+BeuehiLFAtwvKhKQIB
dkHcK8cM+JtAzHQf0sK8jmbMp8AcUnV7UT+xjkFhK4IhqQla9kG4J63l2Wizd8Sz
bVdQ++snOnnRgsz0WCM+M60/rD9J4aISGLgfev9xEwsi0ZAQD+Up5eiSqoneLbyl
R02UOUh38ZGEDeT02TaVg+qlQ/GVNGXSepFwisyj3CxX4QYfs+T+XyUgmO9Is6F3
zYty43d0MnEiM1RCW4tsNoAau9KG2wlVUzwdy0GEnLWnqzG09lnEyN+aanmDBdva
hqf1fOBYmbG0PRGdqdUVyIKF6H0081UErkl8Ke9bysBy8Ko0GrMw+RHW4G33N7Yx
pZ7AuMSl+4/nWNqPw+1UvvVS+DPusHy2zk53QzinpSJM+VISaH0k+y9WqMRfxcuH
QXCJghh+utW2BNGKKYpsTK6n35PZpi0EXm0MptnNVjone2388vGPqmwU6UBVDERw
xDeSqkioxUIBbTGeccqSO8pE2jSh187HJV7hVPEEe3ODUMn9nf0uX7NYeLLZJ3AX
TYXM+4wCPmyPkh/Pgv8EGEbjKqI9JIJxYlqgDDSGV9Nw1dVHryJ1sFl7WlzydwEz
ZXjGDga7OCMO118QOGsPhpcrG6wlbG9iPeTt4tG23pQnzrwSgYqyTLdNlA43E+gV
MvmmCqdgS+kp+wVJ6uBOvySkpyPAun0aYEcxmYi2qlW6fmNes40xKQwm+JhMc5Se
iXr2rqYFuDUIpY22aiKTgVWE65iUOyBZcLyUmx7k5YZSQDmAnBjyOQNiC75K40km
5bFL5bx5WRk0CuqWnmvdUo5xWqsQdNfb0ZTqZ+eSYfVpuaO4LdUScBC8ybSSrHes
ek08sZTcDv0Ue8S1h5RL0zfa069ZHMwLoDCWaEMXRKTLXW97Ei7xy9J/pM+ogz0s
5ggaw/dyoJ1nrDeQQNm0GfJGrPPj98pKWCLfS8BpPRcsoyOaACuLoaI8Ui1Xiczl
z4/+d6eV64rMCjhK+ky6R9yviQmp8nZIhJ0y7b4n+LEFrwqFw+kwqZ3WDHyvRlZX
GyFjaXjRgDZMkvVP7YPMHcmWF6NBwxlmWV3lAcYjFZCwybb94HtP62ZWqwNSy3JS
Sfd7087qcNp1J+cHtdGZuWfaJeHYlxTAMzTG1VYH2bipEQIxySIRlf+hp6sCMDGQ
Dhnjsm/0CqHS2M25ZSh0JVxQ34NeZRHeSefmojVDgchuMQgRuaqVomCdDT1sZ304
h5pOCBKs4b/J/F2Ffq+CawL3rRl7RZYmtlEGB6PD+cv0HiipJ67s/NzMPRkTRzlI
cw6BXQoxkHIAQbPubshfcYPPj1FRoydE1M69Lsu70LqdARunvACEJPqBTB7Q/WYF
DlnFarMrD37APJf8WDO8XTxI5VSOiyjOUitt1qUPYB79ObuhXSSiWF9y0qzgImzv
q+cNto3MRZUkMx/X3EeAiIFNmBRyXxbcsCY9YxCIkYHdP1lWdAIekR3N/slHQwk+
njTekxzlXorNuX2e/dzW09/YrbeCbWSKsxwb4ZHUCUJZXLxFmKconLRPZNvo/52y
JDGkhLfAwLuCcoS90KDHKk8bPX3bD0LAMjaqUw3I+Z9b4kJzzxlD3ZBHMWsX32Pa
0OR+7darBD8G9owPCGt+0lP6HaHpqtP7igbNd0U034/OvF2lJtqC+XxkamvqqWdv
Am+FxWRQib3XT3lsqwTYOA1dNuMNB/TE0hyoYsD5pHE+qhW02PSVE6QnMEkcQxrU
ODGt1zWFwae6Jtpyxc627I+zh3dwHvYGPnZ35PYmNa0VvnjprDU87bf3Ti/NZD2n
qOrF9aUq4OHrHd7P8Qx9V26YxdPoHZYj+gEDs/zPVLfg+83xu+6EmTgcnrZrRIIl
5KlPEK0rGNi0H+Mf+P8O6jd88wk5v9/uoQnfYniz0mF2w3Pex1IULjPVHyz5SKwd
zvlDsIFzCk4wGVWGLJX5ovFYpqTfMsw9Yx0xJcbX2ZNsNXnZiQAKzGp7KCs5cyH8
tWmPG1wqP+XbdMlM1kV3Aakp5uk687SWZ3k31diq6JvWXMxCg3s1OCWV+7zBUoOp
o8PseMTzDOdeYfiMkve3QTlF6iUYWhj12oh7UyGoyBY3tGPY68u6WXVUHL5svUYq
a/c+lP+O0OCPjI+L8XM9AeO7JtgCE30YCIAS5oxYK62rrq6WMwi1//VUsIl5+Mby
5SFqTg7OUvkMB4wUA7zLFUTbozYEZHQrNvw4yMkD5FMXey/dCOr9SE05v3z7dBkT
zgQJZ9WqQRWSLacYp+E5uegzAWdZSO1UfanAj/XhVKj2ntxvvXLWXVhojQILahDa
+kVvG4r0Xl42YKOZqmru/XcLLqj/JAqFZGCRAoxmGTkyO20lmFxYcPH5bijSE3Yt
7szPCdwNcz6rpAk7MxiHzH3EINMhCYzXEkAuTj6mOrLhgpKIIsY63pirzlBiyrDU
QZH3m7RkRALhIg0+xUsTRhRj4gNN7+hLvYtdQ41E4DO8aKDtL5cSaEXe9nTkDlff
WEugEXK7HaX5v+pMI6XSWdupqVq4ffJnUNv3CY7hDsFhB9VjoAT9rmkabz+u/gGt
w1mC3BFGARbodk/9NaSztpf4+S5VG+bsZhXliAH2MWYlC0KKYzSUb9pVbcb7fIaR
ues9Gs72mTAKxtr2UaBa2RPIQDVEfbOepV6C6N87gAPKfB9e4ldK13aPMbrpWTUp
oF10oVivurnJxYzop30WWhMrLzmk/PA7swbrXnrstELmOdM/5oVfSPmJ1cJIlpcZ
YrMp51uQXN6rLCgQJw6Dxxh7S9ephfLXDLqVpzCaE3MizT4OataRrXka1kQrWM4h
olScTW6DXLkRr7RFg5ICMWnbvKruWtasBC5nCxg9aAW163Fr+bUTJo15xr2KF264
kdZE1W3BpW5IzcsF1VBPD3LWFUNecfr+zyXGQsEgk8kh9SDc165zOde2sfPBCdIO
80ZDv2BjgXqnaxXgOxZfLWfI6n0/UOy7Yhvx0zl+gaR9L8WCzuPNNlBucypPk0k4
Cbm1bN9cY54hG5C+m5c5Fv3ENm/yibVzaAqWG9qiZXO94LbNSj32xejIMM9e9/PP
QBxtGapiY+cgbv3FabHj8Ui9mDShh1Ndbkj7HlPYpSiOYN29pvups01nO1Rcsjpg
nqPxCDTgoR7NeLFqkvGRVXA4uMJm0rTsw+DXnlpWX+v5a3b8pPM8AYcYLz73xJOh
NKK07s/R6NqYlNu1kRPMt9ByEVBE9Pd7FFNM004u32cOmH9SY8G+4tzP4HtO/GPz
RK/+XWC77gJBz6X9QyITOCeDJuEdqz+MSGbr2lanzwJFly0pE6KUWoqNyuqLUmO1
k9Ns+pfBj9BPVqC3fjGdvNvrLU7DDtwYjgXuUSWlr7mLjXZYQo5aUHH061yVreOF
8TIgFC+mB6DWgm6rTDCLAzlufqftAMoMbn5q9NbprnT+ES556vt3ZBqlI5PsFGud
9YcOOd6e8ckSZNHUPwPoVWC02B22NiUkNc9VwTJRawsbLJ8d3zgDxh/THBdkubm6
V5EePU6CQKrbawsTKC4augG4shQzd4uQEpFTnW1B6JPOlyllkkRkM7mUJlcvi1rl
1qwDOaY+YOAD9NsEEbQBftC1UhMJH/X+CUMGgjaGTukDB2JUvDWZSS6zLyfBRALk
oEssEpYETwzq9+KfQMCbTmLhs0U1diKRKWyYOT3cdZDUcAtxnBcC1Kza00hzKWtB
wHWUgpLDuPjZ6Qlw6dqKWFPNTzEneH5DIpoh1j79XFJ6vu1FnLNodgeaS6WYz3te
Q7dfsTkv3vY4v2zhDRPzzNZ0WdeB7mdDBsNKgCryBGq8Xb8ITpOVOH+jdeJ61NH+
NLSmrB3EsRjiDgXptEaTT3wSdG6HGDn+Q0LfKWR+dzXsYqzwj1/ANC3hZSaXujXE
6AWkyJd3hs8Jg6e1JJL2LJYNyFMnhrgwepDvbrtOp3bv9cYYZYFRtAkvwxZA96YR
j+0OQ9yE20SwPIuOKoUaPbTzQi7AhZ3ZBHbNqRgyOib38HAVTPGYTGbVVN/0M3Qk
lM5sb9SLw/HJHqx2ss9upUf+j3h0CFdqEKnuLgw65sjTH9lr1OwWZMIt/Bszyh+c
ORgQek6mb6JoHnmSRNzKTNXulB4hVWTlUDz8dJUghzHb9q/xXW1BzWxFaSybJ+3z
rSjTDWsGq/ty/S/x+EP2fQHTgf/02pzCYXdMZz11/nJ8qmpY29/0UNlWIVzpwo/M
foXrOHHATFmtLgRwh3zWgNhRTJpR5YTRgX017nIaS0VCqh1rDqFA9VT2/JVFrKhG
QtL8t1l0NkoreeCZkOpPWGp8WX/r4QL6IFWivZC4QqAzDAGFOc2Og4nLaE39KfH3
qbmzuTPCIEOJjT2gqTLpHfF1kwSfWEXraLd4Bs6NsVbLrLbLYP4icYzKe5zOqhG9
UeySZouql8VNg1zuVixMHBK79ybeBmwu0gxn7JuX2pCBmDuK9V9tnqYNnzBkPi8I
1v3AdjiDNGWiKurjq2dCVjNLDXLC7B/Vy5Q8Nl2kYlHgr1X9eRV6lPL2U/yCJvV2
X739+OKqoSTf3lBhrkOupTBkGyR1hUFYCcFRaknuN/yP6FdNHnsMyT8v9IMcOwhm
vrETiaBji5DBtuqK/k6fdpdlXpUx1FOX1TJ03cCEJYLx66V+QtGAIxUvLsZqBVSc
GfwY9CinJ+ntrPHrhg+bhhF8C287TFf10ENI/xI7MpAKlrXz+5fhNzMZ4qF5x+FA
W3g17lOcff/kFEBlKHpTRHZbi0pk1qLrM5gaXyrHMP4TF/EMGrPC6Dr6id9iTMSp
KFdEvJwHIdsrbOaWvtH/ce9cdZdqIZeXT05YqLe934uBUeQy/nz9Aa0+f42XPQIJ
Wuc4IMifrodbWhqIjnqEYfQwpgT4Ff6Luz3opgIl9GFqTXksxozk2P0KV9qRajT4
z3dMeJRizig8cPEDoH48gJXtn5ubLyoehWoCNLZMNBYkwClxHGsi1KmkX9Ko4mSI
eNoA0cde2VhjMu1n93WsEZt3Wj1noihJs5cfrWSgR88HnVgmlWYo6V0Wpkjm2aaF
JMAidk2iDPIErq1eI7VDk2T+5BLVOZEljU5MsYRehVG/4sPCevZW9Z9svyEAyzk7
+W0ihLeNZcMrUCMSnInDJlqc0y/mA6YRMROrf9G7WFlvFnyfqFf8nGJkeNqB90t2
LtD8qiEmz4Fb5FCL3ZJH6pxTvOkk8eKFNmflkRn0+zrqOoR7qgQvfShZ/PcL2R8N
S/kHt++EjscjbmJeNvvOvQ0nIsxhapN9xKFVC7J8vb/RnpOLbakZ27xek1HeFH3o
ufy+Of8xx6bNUQuW6vrMAZwFyQ9hCgU0zJtwN/ZcwwiQ7HwU/SN7B1KOCVcDTlki
zNEPSMhdLNQxIo1RJ5c2527p0olte6fQhU7TVyB/duFQ0qcoCjVxq3vRebblVbKe
SjeglL9tPhzDDtx0MDwLz8gZ95hDgX+umRao98w3/ExJqku8quXeaNC2mK2BzJhC
hB6pBCokHUWe1vLDhv1rBNCPjKT1KLeG5RVW84CqXkLRYYyT0v8H3HObjlxZ1SbJ
rqOoLVmcnRw4fTqZ+QPxz7Ail2+icOo/c/EJVCxH4ESQESnFvJJxvr4esdDQ7Zl5
p/mklgOPKV3vXAi2tyDKY7xY9mGJtjo/FEjkFI2E4siYGHTBo/9FEIggSsPR4tSO
7S+C3598PQiWNGvw1K7UJ8ct3G/176ZR8xqkcAKwqrdDra4IwEAG96l+miozZtp7
PFi+kUsYwUaTRVHBu3U8CVKzo/ldq+3V5R4WMoKFZdprgeGyHrrWn6CL/hT9QNFF
7SCFfH+2Dxp7IhM3y1UmRpNwtbojUXjf2bd+VCsdJc/SxGbhCXSixGyPM/0a1YcX
RBq1n1fryHo5Ts07kTTGez4ZOo/L3y0JbIz8V7gpBaim1ZE9PM56PjOyrU/ePI6D
7TuHxSxWyectgcTa/vy3xPxCGgRfoNGRbE2/+CFfQyVydxaafVs28Pnk8RKpuErN
GBy9Rs4mxEANVqcBofqb6QEOB6ShDMo6j4qxPZOBzFVBit30fBc/hc2KbNB+hV21
VmkxS6/KRm0I/T36F1/imxa1nnsaIcI+JHQwunsTJP5zjlIQp/QxuMHZWbWnacbO
Dj1bl48CdGO1LPwhZTMlD4oITWa1LrDdkd3Cdudcw8oWAL9RVXkCS03zBPh8eGSN
dCvlcL4jLbywmtqq0Vdtncu+3dQGcdFRhG9qQ9EzXI7WMfHJrcuk36mLgHfbPB/f
v+CsVoSUf/yrSOuwOx1lAEyL2jjZVyihWdmL7lknhMuDVata++2sx8M8GxyHtlJL
DE46xMxPZA59oCWXZOgzFaqUdjFfyVQxX4D4EPDPLvkUK6YF8ZrERQ5NHHRjBSHu
m70jXkSGlOmoAVrWb7IBNqoq/DJUHIhRpWGc/JvpxUL7pkeoJ4hwOpzXKSdfLM4i
pidzV3DQ1Pjmc64XS65bWMnIUwuFAiMpPRMXNzhkbexSJAuauBvdAUhRLrzOxpoQ
vWttPBfsoEmoymnXfwxx2wBmdzm2/H962pX7CNUsVM0FwwU5W938HIOXxXVfu6Sb
43Ugam2iHiHVDdgH5p+tUIvjz+NvMyk9GsQfFrSV4X0WYyJXzYRG2IqiuhE9hgyy
1Bcj6uIyXM62XYrw0C1cLYtzdsBM8bTHsb8brK3LKcLjGMAsQb1FBNUUawrAqcT6
SuC1y7xaS8ldfEAoZYobc9YyhPHFajfOiyX9VHZo4lRdNwNYxp6qpC1VWKuAz/QH
lGjpzPUceU3Hvb3478keLa9XfSHjEkztfFgNDztOg9qXoj8JdMtyZmpLr6QD8Z4Q
kn+w1Bc9exdgK6LaaabNbcB6iBg/6besRv7hQXSENli9SXTJYlBqNrysQJQlLTQY
fr4jKwyRKF2IZEOD5rq3y1ec2RJyl8gF7ccnNhq8JRyY/6Pfz1jLmu2/gowIxVxb
oOt+lDXm0IAtdiZG+ybeniqfUMsxKs3qxzjXno4nCRb4NfmfI0m5JvZVw9ukA9V4
BsHtVUyyp/1HJZ8fOrWr1CJvshpEcqGnW3N9Er/hGL0RbNZfAVR8tZR6JjS+3AgT
MkBtqhofaw4+I/5Mg6Q7mA1OpcGDl8E9Ym703QEXq2UZ51e9bSLcHN9bDlltxLN9
SZIkTyvcXQgdrbwKiUPWc4oShP933S9t/vLmip9sipJrr5q9OT/NFmJLLwaPDYsK
YElDw2gmNF1j4X+e97TVJINTV4fjl5gR0rVQwc/4U+Qv1buvN9bW+KCqBnJtpEVL
EiBerSW+YJjLT+go6iGpGjku6axxTEGLzDIwINtDG3FDRuHwVWSWb1xttHaTcCQo
XecaoW/hdijaad3X9t65P7CGa0uvj5qW71pET4cU/4TQy0KZb3m3fdNyS2bYbbdj
ijmkpaxEj+oQc97oO/Sa9PVxCZKNz7eCikfUrAFMmACiOM5TwUyokkGXTahqwujq
GDS3lcsPGDr21bULsfHojYgxOos3YuCZlnl0kXNTYZQzESJZFmGSYyMCkFEbKo+V
2pQgJP1vCf7Gwxl+/f9hhyHFx7S9UZFvKR+9c/c8gzylROSZWqPUSpSCQmXrDT82
ZRpt3LVihae+Oc/b35HMLtWe96SB4rcpKcLQRREd4bedKeirttY5Qb7RACRN1TNr
ISWoPFP99NNSjuCl5HfZSfk25qbRp9QCaFY/a/N6qJ0PNMDId0NVKP8T3BBy+CyO
jjrpuLy+babUPVszNDJ3xx2IV4ZGLk6Thxnu1H4scMnz6pG9omPqqYN9nxb9x5Th
9lT9y5KBT6turkbSNpKepsZFAIG6YP0YZc2updA9vKepKRTDvxAgiHYvNdp5XemZ
Y7HFGxDbvht/id59LQf3ljKNGAKUFuROUNsNmRRmgV5LvPP0QpleEP131zwqx73j
9BLbDEWzt8akQpL+3D8H2vqchLVwT4vyI5VoPBSdCvtRz4RH9j2FeXXEGAGq40ep
GHe5VWo8jxqJ8P8MDwsWHkfGd9jHS4tQ1eK0ETSVAb8uZD5CwxviEDAVzjx908tD
NHBpL7CO0qm0qCc3AMOGRrk85/jMENxjqi4OkKhHUcMzVP2Gn8R2aifE1+lOBLTF
y2IOiQ8HkYtBOk/vDmtICLoF1EMEvHD693TlT2sMpbyqc6rAFHKjpAVoVEgZuyDk
gcxj8UiCaZ0r0nK67FEaa31kzqoxLWT0WFqL5T4iHoq9epYHlQroie2faqIvL7bI
pRr0HZy0Q0mjK6okYSALBQtiUIuLNWawsGQsHlIQx9gpAhdd9fsAd1fsS/Evhnrv
iR+iXWMimN7nRzeU1cPg7/wd4rYMMXy5aHqpKpYtsWtP66vk70EmSE190k53Sj4g
TdB2b0hrtbvlgAmSXrmzI13MdSWI15HXDwsw/hP/51vFEEcXrcnS5JC+X3Azh5i+
JfxljCxQAjnlRvlDLixmtLmrHA3ArUpxdtHym1MZC8zCvBuHkVYNcPOW9xJlCoNn
/dklcbacG2gS5ePFlL802vmp0BYxihH2pbmXjfjugtIhKP6zqGSgul3nw4QnpgEK
pZiLf98AAGbBinbwLcJBkse9abdRWVRjbKG204XYw1EbL98obJcUo/LD04w6vRuC
rW6LlBGO7D9rYZt/Rlu2Xkqs2EP4jbOvHAekYAFqym7K3ESJy7nTJxrRaks06wTC
m+Vv5Y9eNWyyOO9w/7t+46d4pGoZ/zIcr88I8uJT+i7vMfwEmYWjSFafdImbG7kl
Mej+rBg8MbMU1TFS0bhByIKodqMBo3nVc3gzGf2xuH0DQ+DoVfAVkf/n3ptIItFm
ZG5xzNK1SNhLPkiM3FopGMU3kz2FC13G+9Xrm4xOk6TZo8R7U7jAfxB4MARwsdfy
wGfJV3/9ka03ylbTWK9T9nDftlwgDIYhsl27nM6IphnUUmMtfba0/YEZ8GytsaWx
mcNDxfOV4cgneKGQdoPzqRyHPwhcJjcR4zd/R6Xq4txIggxhWXHULdYxcF5DvWDk
kvpjdJeUaZoW3667USvW8K0mKxCTzUDG7z/T22k9Kybs0pfFnS2qXSjGQF5LexXC
RVPDV3g3anm84RvOz975mbYS9bOCmiUCirJ1ZOwQddasC4efDRI3Nj61R/RTVLYx
g1ITLcpmLq9Bv8tN3MKhP/OwL9IXDubmXIpuis55YhHGFcta58yy7i+TIdFDS+5k
XujxKOMbZFJf6XZDY1QocAHGfpytfCdV7mV50M9kFtopQ3L51EgJR8DyY7EshfRE
BLI2K6Pn/lGbpWJrckoy+sh31WrX3eSiFmdPl+6SPdMynH54VRKg4BNdwmegsrVs
Q1VauZfpnafrunaRE1jhvh62mB/8HuidH3PNY3WVTEIZASU83WVWGGHfGq2O1UUi
mtmo99udjFPSH1CMAWb2pBLubG+iHI9aTLqsxnbT/qLr7F3WQt1QYQx9W2wQ+XrD
3zN80VhaoGMruWkbh+7HVYgQF3plUumD9ESzs41yWBWovDh4ZP+tZPH3Xni7si8N
JA9eMS4zDVsGydz4QSl1LHMiUFpLiaZLwn5EywSCuw6vx5kNm76ubCT2+u483kco
MEAHTgwezkWmzSSi6nJevUt7oY1yYi3GIWtxfNxNVxUjVIlv4QN2qG6u6IAxDdvK
HRurH/OEP5ax2fYv7hnkYgIZScUedgttZiTJkZWFE1eJ8TkyAABr0egMwdy0+3aB
5CjMhre63FCCfoitNXGt/n9fO1EAQBHg7Hk1hCOzLEPZl5XYBmk4zANEzz+n+rWW
XRb1nxmeAmbSLY28WpeVcJeERJtFcfWHJOc1Ran0xU5gMmzff6zFduQv5KRXUwHU
RKP9zpPdD2WVwW9b4PjLwluuQlhmfantiny/i39woPx/Qs23nReBDTjhVEq3XFEU
gMqE0mPlGOCrfFR3zloSyXOL2lT5Z08GToStvJzg7fogjq8EcIE+lrYlDg310hnp
UV9+sxAyefRNg54XGCfA57/39qZ+A80jJ602xMo4pMcJX8xCJeoJCDc5T2bd4dOB
4uP8Lp1obV/PuKH2temkqUbFv3YW9EZgcs71nxt9PdLm38OtsCA+zVFtS5NhXfug
CIYsKxTaoTeI1ZbtNSLWDSlziQ40WWN1Ddkmr/2NTNx+Pj35QwXj/SO4K8DoKAIr
ZX7Jo0GrOKQbOVpdI5KbNVKMlO1zXNOkIvxcDIeiCdCZ/Sqz3scXTjisPKfdsqdY
PQeaT78GCSUGJLm93Yastc+UQoEn8A1wqeMunXZwUaWEyR8KBqGf6DayAfGVCcVZ
CwqkhPi2d+cAzbVNCPmQH9r3DGiNarIpEW1TOyyGuOE4W9jbhTYyOpPu5+e2jGGz
j+cVEedm4cyOYXxC1dOxvcMtZNXrtRjsIKx6zIHuMLVOS2754EGQtRq8Ey0MWF70
iN8BHgJd6IeV6kGRxysKTyRHVqYNGz47EsPJLdTTJUhgAWs4YyESdp4MiZBtsElL
6Z/QDqN2JFGN1OarVuDWgwEL7xkSW+TUGd41M+ulKD7VNeWpbflsxye+nDP8KbQV
x5la7Fna2GhA2swgEt/bs7Js0jmHljaP/e9NyCK7F1Qm1hxWcDGn7HNkXkJLzn8F
MEqB5YQ2BsRAvkcgleykPUgA4fbVsVKFE9V3LfTQ8VnDxwzb+8h/lZe28iA+zOMB
iG0b4Rxn5FeoHqoSGxE9kDbunS6N9QYaVcpbBDXZyf+79ZxC5NAz8UJ4siEn4gYG
7iB61SNYE/ofurlNTWAec9AGGDoxU/v1+bNv0jtRanWsVKlZBFpVlxZJYyNkrlM0
GkugZyzkAqNe82/S0kO/YA8Wo0RFRL6OYCZNlZc63MXTyVD8x2B/euGL0lLoQl1/
xq3hRaJ+cZMw+t6/B0uLEuIa9TpW0+LHXhbDYAUW/Zi0Z4pbHrko0y/jWwYor023
loYFx7z3NSU7dasmTBEAnpDnv9XyEP+xWDSY7QoNqTV6UzT6rO+DssK5rfrKqGZ4
xOTdlIlECjAjeHd3fi1QaEd4vdN3bVp+XIME14w6IOqpFJN6DdsNSUKfYiHsiGDq
sp1KwaFcIFQ2+3w+ZBVqWPX6G8QQoJHcXhjXN9Ar6B6UvH8fwie9zThL/wc8L/Rl
5R/MZLxErXW90BSjKHU8C4mBGBSKEHN5lRBPneTjKn0IGNRZHgm9cdLyEocp7kkK
Y3fOP8UZpYWqjmGbfL8U/a4+y0aQrWKKq195optu3GvM40DsZKLVKPcLMimABBRS
0wuLPezGwviZwLgUCILdbsDDs26EPnjqrQoD4MRdWQMQYYyRA2pvkBM8fsxOqW/E
Lr7BFvEsqS0H75MfEgOCK+4Z2AUCfEHVoIQpW7IWdEWn3ihPyJljQ8PDpbsX8/HN
Op593RXfRZ3rxNTIU5EVCb4dn7chzWmwOFuoqlb9cXRT1xwzbsR4UmmL5eAwFO3/
a6QKsZxastOPJMNEDaXUnmfuTia394H/lS+MxMBAE07/pJ+UmEkNdS4HI+6Nrtsm
oEE86jIcrmfAmm6jAiLs9T3Sv/hL/2IyPdIGn3cpz46QMLC1CPv18bz6n0yJQAhc
vL2qH+l1YWvgIRYqf6liovqV7uoAGl/B4bIlAjM8nDWLx7t2yN0NKGq8yB9+HrH6
LgH1rZH3RkFgFWL8xpEhG5xbgJQpynwGdmu4YZmIwuPciJgqOR/k0rRVxHzSKQqS
AYT9rYHbXNpb2is+qfsYkSbHKyGYjCMsBFE+Gm5VSpGALImJOFYb51hNaVQoxsAA
23ZvGc53AFFu0ea/5s31jZK6c+JJ7sf0UzqjYbJPFdOpGpIAYxU/UCWSnkZBBwFJ
mGZk43MvzyRS/iznSsBfjbIh5+riN4eKK9bz9RrH9/mvw7G9Ya602Y08f/eFSVeL
FFcCq+zNyFV79FVyVqR+e1N2LfaV2dA7aLlj1JVqAKMZerELnp69irf3sOGW4cky
B0jROurGVthaigDP9G5SaiVWqpMRDpINKPFq9VP5JnA1618WCwfd5I7vQcIZp5ii
BmtfpPB+JtT39dCEsJVD9d9jPPgaV9YfhRqm0CAty4zUiGBGcOSvCIm2ntsPNBe0
kf0Fb32DMwSTe9jMhZW0ftZXcn4fY+3vVqSn0jn+uCtGxmy+kCkYdVUa7UqT4mzj
SONsPOTU37lOOzFO8vMFqaSqfrQPiixM/c9d9Ug+xIriR7lJxKHLzpTnaCprm2em
dctVcKZMW+pn3zExCAeDf6dZzx4+IcdN0bQxVBVGPveh2tnHQ/iTbZZwA+qt73IB
UyaDmVlfatEsV6ILWJsE2XJzB97ioVMWdLKZKUgp2UgTh+Veg2jsMeSJ8m982fwI
BLW7wsD08XVe9XwfIsqTvCYCiP5AeJmZJvim80gWW/Ce/JbU5H31Y1DVCnWUxeEi
de+BdxO/Z5amTUqs8Xdz/Y1YkBQ2GMXOA2sZR8hYoX3/35sQwzWoX52IxgGkzmFE
LhvWU31BVetHM7rPdmig99OVNv3hl7MGi+4NzgzK9Nux7IrUGluVRUczOOMo1G5w
SpQlI9NQfR0nDJL+86hXZcxh2yIOmBt96/n6+hbVcpedZQqgjUbaUUDRHShoVACw
HPIAEMtK5eKMWpobjasT7F8aAProhwgmusRyhdDNjoA+PEoQ639FPptIMsvwa26r
Mho7/KTwI/HOF7T4u5TQxZmNBjCb+0uIwkisO2gPTwg3omMiuaHJJGMkF/yNQFsf
Ebd1+eEdbIgtp7pOF89bv4HqiBqhtRM3w+dKfkdk+6hUHDO52j1wnCNSt88ONMvg
nzcWhSkMW9Xh13szA94WKIE8saSJzOo6OkaVT9oeQdlB5kWXTgAk+KlTPU7C1hPG
nltCnk7Bm0vWjwYOV/WPA29oNvTnbDfDB/K655IhqTgSmf9O0GLLykbEgVqqPCOs
J7hF52vvDkMawomrcAlHU+v1PsW2ugZbf12F7tBl0fnU1z1/kSGCgP3Og9Qe3Dz9
wEcvaWcxMLNm3lfCoA+yecWK0TZqSq/ikrXkjA2M0oeSwkZ9dx8DDpeMdGLsvZte
gXnmXh85vUzThK1A2Z4TG5TIQADy8WosY0PbywF6pmOAzbm/FPPJB8XSkDkSDD58
r5gFvjTUh/uoS1VyjoOMJQA3WWpG/WPR/S+mKaBQ35UnYGGImTfSn+hRAgseE3ey
UIbuDvjc9Zld1fSvuMv7gDPQh8hm5U+YMoCGEpSmdPYUBpRL7jzKRY2ss0iuyyM3
1+OfOYde3oOKG/haWF+skeS0cE4hV/21BZHOJc3PGoUqeFv8E+6H18Vtocnasuhj
vHFiRd0ZMBbnsrtZ4wmw1GIJOtWTPJpLyr0YngomU6kadoph42JG8PmNhQ0439pe
jhkB378LV7z0vCpmZVYSTxj0KTuTCTzU5wFbPI6uJthUuOo8k2h3S8a51NyizmUt
vSg4c22cwGuI3BUXDbbxjIezgxwil0JmJ/upfg+dwzstNZvLvqIF5PIvYAzNxAae
K7QWxEJIpFfyjvJo99QWDrke5AfMt4n46fZKeqJNM6aQY5lFhjBfRzKFIVqh69jA
cC7XpMfHgNvdCronpzOCzCTZdT0/ihKaNO2qXRh0+HrVG4uVP8ggVc1y2Ky9u59i
L2AGUwIKIDpnXsFz+/bAlWbsq8jl0WNrrYpGQA4swHRpJDyYOIMcCFMAsYX19Dtu
TnXvFWLozjKPvvhtyLM9dKDuxIX4X6NCiL21Itt88329JSHqb1Q5rAETbOn5faCK
F16k95DTkzZRAMGoVp6NTMIrdvTvUbCe23fJ4wWN0YSo3Qa/BIBmyK9TSO6B48+X
Y5FHSn5o3eMIS1ylba9JkKzHE94rrN33A1Y0WTi5gj4TMEP6wDIpwWp8jjE78ku8
tM7UFDgVRewF6cIzn2Oa5F+8N0mLadR7SDhyiyuYCPWChrchOe2LpWnoUQ2zVRuu
2HkSTJMUpGRUDbrBX+XCkl1MP37kiJ1ymolDSGLiHklqWC8Sk2JvXYL0djEySEmK
jUhzg6axEGXmBGr20nRc3r83ceEsU2JXKhxSMrpM53Pnuv0U9Fydu+9u8zAkGRPo
8bWFVpCXUcXugZrg6sOD5wJhBPwe593O3LC2i3TT9M6wn3jw6Yzw/RbIvNyGWUmL
9GiOOHnIYR4lpu9FDRRFrohFC+GA5z64UM64B4IjrnVKGGYob5cjhM4joCSZLJ2C
oencI0qaY3YSy63GXrH2o3bLc6F5tjtAPe8WHrrW37rOfIJMZVhCswl7MaAIaotL
VQF4TzFDtxE/Rge82EtMIJDnf5T3xUlE5G2qKALBMd/DB1JR6mYfv8SeQWDumX1C
nybKfoOvx/8q1nvHt87xzMShZ0maGBb2L5p7LEMYehshxwjmFi1TtXusOi/X29Lj
O+fRCiF5p0x7/77EcsPi6N9xpvz4EoHwFJNo26aYRmvwp2cLrDuIh0pJDU73u4uw
131pcuvPIs3Oj5K5YnBb1PisCS7xyHE8sswIJ1Jryub/Uz1pfPQNxAR1wx19Drf6
I+af5Ps4rW//bDpWuWktFm2W+5uUHVGS4rBbdef31ObY+grysPshhEzX45d2oSBj
JMmYCiKq85f5LP8dMWvBZO3ytgHmZQ82UZ1BoXUmA7fr0mXyUEiIX+KzLPjjx3LZ
W6An12gsdjajWTNJ9dwJTT899a6VlsMSCbL8/1jRFDZP85q5zX6VuvTPeDXcXnzT
N0hwcl8wmoGWf1044NpmyovcfNGjYoOwCc3cmUcBw7XX2zRSmNG4qwEuaYpM6g8B
gWlO5LwkSGZiiLxMgcdPgGTqhF6YF+9JDf1GdVDiEuOk6G0m5vGOnPLmDnplLHnd
yIy9XxJoYi9XPo7r7cN0Mcp5t6XQ6T0DjwIpACVjVzpwlFoFvYb21Cc7JJkxgKFm
r7Xnu7Sa9Kmd3wZbsV/PJK9xp5W2uDFKv95Ss4mwaa8ISR/e9bmeOzyVaE7EYPsO
wSU8Eq6LN/NHlsnagKUYGKmvW+q4QYvZSG2I/rCGDUQSGs6pvarwZmyhCvjBuM7y
bVGKHDPeXSOpz7xAC0Uctgterc/JPcovqG0lBFmU9hivPNSHTH5DTeodVn1686vu
5t1FSaeDJ9KwZTgTqmOaH3glfqb0FEklzJOFA4S05X0CQ1/KAi09QpITbLS/m5nu
G+YQvuczcy0AkmFJLHhonF1LoTGmXiNV3l2WUAH0GznIwVVe+CV4lCZhXhDryRNe
7Dvx3GgPBzb7pGoyRW7BhKTzbtCzJObG3gMcP5i6/95XX3c/U/RcBWyuYL6VY9dl
VgkraUnArpc9PiEg88yVACxVkNny3VNO4JD6YR6cFh4Cz0bLCsLHXs5sCrV0Wemk
ETXyfdsiZXmuhyXbiUr6DtCcxsybZJheSP0vkY4BPSps3BdQNwBOvSVPSOsPzK+r
+srHewMJmJFimDYLIxoz+66nBjjTI5TYV5NdLQX6iG/ya3y7dIsdShxJgXo8gbwO
RQJZTfdm94DaRS24xOTAywxkTBfQNYQpmKQYPLKThx7/fMHE3p1EAOhJC6Ql+eVK
HtKJ38ncS7FS567d2ndbs17BjdR/YP86UpZGcqHCPRimohTNCD8wQrfKrvAzuPAE
SzkdhZZxvGukZgH0PvtrijuHW09m0AvDzheG6+EoplGU4VYjUGpdPzEbuYLUtYbS
IEO8VEoJNIx6pqRa4h3gngO4jbFtDyhASvS2c8fNWZuj6wyVCDzrYZ46IPUY9kwR
V3WdJZMmQ58eNJ3F6T8Ah34Iuz0IajiMWA4qkkRvaN9+ZykR50e54c3AIi0aEcI9
+q0Ic1wC9FQ81g6oe2sq3TTOco6jE8CnKah+gQTZD2mTyqx0Mc5gHAHZHAxUlez9
phnjOLePJ8X3RE9TZuE4kqMfsHld6s+8GXLDv+w/P4fubQgouMlg3tGzNW/PvAfT
eHhl9ug5PnpJ3p8dwtmo06ongYtc49rTtfhH7/WnTZxQFmikdCOFCs3XC/xtq69L
MhbLFeCiZcVgIGcPZgQ8I3v9M/6moiRKJL8dKMzwELxrgtOA/ZGOxaN7eM5xspzg
zTjekP1/BXAnQPUaMbyc0g8x4DzvBe9ayq112b8H6na/PysYOMsQzYWPWAt+Dx+Y
szOM005sYJb6gZi1q/BFzLU1ZEwhtMxDBWIb0qCpRcNwqr3bj1DDZUWGtqcWz4Up
VRZsWfzT86LAKIjMFvaB2l3o1Qinmp1jpUCFZ2RyPT3swsN9Ygw1sU7fg6MIMFk3
NQgOuLJaJftDgSUWMONRgs9Ihat45E8aA9LgkIaixCjRFZJIF8I391qBREzOl3q+
SZhBe2M4MA96xQKR96E3sn4GriWYa54tO1xvmDEVGymvKFJTxVbqYcvYeVi0S9RG
GCmvbkSPHVtMszy8lqjy+cYvpNFcoPj3CUOFDJUms5D67MT3rzJtsXSTFyhjq0Yw
tUOQcuir+ouop/tugaEmabIRmYG0RIR+C5Q9v9Ozc5xjdZQ8X2aGE+QvwmgfclXy
g4Ws2QSLy4oUzH+uQL0bKXKOzJ7GS6UwWFmWMUEkqDFt3/BVeNbI2CAh225k/q0z
bpuoo2/DBDTS6HpzyHpjnA5gmlpUez20vS6aHRQbPCFIJf5Fza9XS6o2ypD0nk4x
FzYez96ygKXHjpbKXNtYOV1Abg+gV2F1b5n6aO9tcrpvrV3KKOt+2bZvyI3hplhY
t05UcBR9FIkZJxWeSsvxvIm+1wc3kq8BxpnKziWXBVN435S9SPMQG/M1JwOAQ/r+
XHmTthtI56xmaqqLszhVQQeE1yyduJBCoXY9dtMbdB/V0O0XUff4+n37M0Jksrzr
RV62rTj/pKw0vlqXl1dye31uuONeUKB9/iioTsRNCzL1e5jBqnKH3vrJOJRNMWOh
dbVOC/XPmerDY6eNF9ALhACoKFg+L7i/ssbXt+m02gPHJh41Enm7VDi0KET5zXsd
vTUBK5fAPBdsJ2S+TmVr782Aj21ccARb6k2nbyFKLFuuIeuHJyXlT3Za+bCcIiIP
z6wmvw8z52PEcKr+o2djgtOVi1S/xN5eY3G+mQDnsurqLWa8NBkrG9wrekVH/mHF
WZWeFKAIbKoUcx/9SmhCiAErQbEn5yJov96tKhL4kQFn+xrhh8kfT7I+VaUU4l5u
MAyr/xq+WIabUqdAaoxt1LuHLktrv6u2DAOPu5UyDjJe8WoEceL0F4JYtvgEqNwK
6s9gceFXtxHdrl1WyBVkTKkhqqN0+O6O6ghyn4WmuC5au0UNmjkheOl9Jvfb/2/2
UDSg1KaThPmwQoqDzwmsJeXSCNe//4hCL6gxqiO+cOPDPM+pSl6c2X6zJl+H81oE
XorgY25Ax8aTDGaQwcTYnyCuot8JNXwysz18CCmHpHE5vPMWSSl5WJcw53eRPIPk
sc5uIRYk5qElA8+GEzYkrlsxl3vR7wremW5mhCgJL594sJUHT3KO9mcZQ6amvbyg
j4GSUltsQMs1hD+PAlLGYZiUJF+sUd27FCV6pToMEL8bdVyYvQL3Rhp5yQRS+gAA
J+zJ8q1nYogy5BgU6g8bg8ymKj2t6kbmd3+tOhzv4lEqPdmGirfKvP2p/bcM9elD
Pp0vWl7ko7sgSX0471ZYzUDBlAHU31VlA8Pvu8Xk2pBlkiz1Pi//N414ulSBNYA1
GiqrUe8FLC6Zd7uhgENw4GBbuqn07RhLAOOPujJosY1eMHyz0YETYgvuiypO7kES
PE3EjqML2fgtYQVOi45yNFATaV1o924mg3LESs6dbkVOXvwnZRjWkvZteTBq2XWC
wTlP3hKVGZT3SddX/UXOCvrQomAZzR+MoxC/k9+crd+Pv9afwA9K8GyZ6VLxU4mg
YP3cJ3+QL0v+1sm7cdKOJey/kr2jYZwhvlGoOSOwhQIcOrNWZKs1k9yEu3mcS1vn
KKQFHU6JZljamhrUM44/VxmdRIthohMTvlE89yNuTlf2gne6xyOFbJKymVUgbizj
vAxRSUlEXhY+BPuKu9T38sii/mqUum0yrwv7SqJIH+MGN6VX1WYE2iIKvulzM+rb
cbFlqoLMoSOD6uRLZfefnwNZaLPqIIRAVzBifZ1qX/4FdJBbdssOFIe8lNS0UZut
QtncucvlYb9QxaqhCEAQapaICwWV5LaNEDIehM0ZIZHVFFeQQkV4gFxPyLFTJEi9
R5xMvPrBBTagkv4fXLLNFEuzilXnVMp0MQaCHxzE9Gtrki2H4by5tLbf0FgXk9V5
oQ50He6jYU3AYgEkh+nGnRmc5bsx5KNDyTVrTM0ObmgTfD30lekidTU22Xp+M4ns
14SFUSBZV5lmPDznTY2AWNVbwOwTXcWQszuf5PaD786aXEktpuDKCgVwv9YPYPzE
s1P4f78E/CvkaIVDr4zU2PJAu/G4SL3kPGAW+3QGzyQiVkJPXa2eYIyH5QPuiK4J
Xb2gcxTgul8058lm+KhfHS/HkZovuXodVBzQ8gC1aEbotM5NPvj9x5dZTAYrnrip
UhxNiU+Xz6dioO8TLE3PKmGjv3HjVNUsfjy62KC4JF2Pf9mEcfW1s1n8oXLQQfDI
kyIDBr0JIisZBkG4uqrZmeBTTkDQpkYWjCXc0kFXjh4Qve49NWSEjh1ZGuIHxp5L
PHLV3v2jLlMljSQvCglML6pOnB2Tek96ZKSbAezmOIDV1HnZEsVWtR+y75LGH0xD
ZIzA6Wl4kCrFK0ajSxSahl1dihw5nnhfdgjoTlorNZx2Bm5LcGjgox+ty1xjUD9e
WMcD/20TyAnu4imLXPKB3PGTFZMWYCe8qenauYDLmx2BKkE87eF/CFHDwUFWhNfT
i5m8zsg5RVJyiPv7Z0WyotcfB4JA0viil58r0Zups4i+xLv9wDSv0S86R1X1VAnh
CrSNhRRqlP6+u5S552ANmaA3Htj8QBvEQhKQWSECu/o/DOrBK1ygFLH/xKDaBObC
MdTAOvko7GNQiZQeZ85x9cJyT1hhFhH73p/nMd7DSimSoiSOgizFIlngvHvXSD/U
Z5Lv/lQsKAykpBrwaCks+dAiyy5jmvWGvVHDnKrlX7IotUAVbM023S6V3FqDbfVs
1+jbs/DnNKLPA0wKE92Smar/UlVyq3sJJ9kxByQJFS+T22xllrltZrSrWH7wQtrQ
ZCew48z5s4ZkRFOAl2kJzb06OgSDYF73YGLpl4jZhbinU/T9UV9MCixM1x3u683D
GR1laChsk8i4cR7CB4dI14IYhijmYJHCSWhQ2Y2u2hj9sybasMycqfo+HPsiIVNl
4US9MjMIJGbpZ4YO+9QADcvI7YEHtBfu01r4nuMHR4/oYbaODD4CoLehFerB1A/R
vZ0TIEnJeiMs5UdpermRSRqVSEtUAuNUhogByHp8nF3AuMc5IuzLy/v9J6z++BK+
KK3dFKUaPZ7GYqaBvAFKI9H6BQALt3pPPIORBj5F//XrXT1VEqlE52SHu6jMYIFf
niVk4/2uRxElALgSKxS44uvycuWYDHHvUEK2/SUOmMAFeAsF5tMQNFDAePaN4z+j
6UnguD3M0FtB+zg5Yx52rMFBccs2eyt+ZKTLtoVu5qS4KJg4M+pK/D5EmO8NeEnl
f8tahezcA/TuZr1m9uOLY4Cm+rJ/vg1YMDF7cFHhE41abP8f+Nm3M9EAW7jygWdO
wyAiC004v740CCKbf18Mq2armaM1IZw98zLtmwtRuzZaDPEGyVL4ct+5IfvmaQwW
ErOSl3mh3ESfhpy0gnD+85QizG6GgDLwBH5YFSJUXEzMhLAiIwF+SF4IzFZnz5Eg
yMmrl7rCyu4M3xGmBy9PfSW6wyfL5KezO5mz5mRgRF13CV30yL/kZmH+0a6xpjO7
1ryPICVDEUFUXl3qsb12M+JR/xAAynmODpCEurCxLrEyQ9S5i/JYek5WFOqT2DWz
lSdctAGUO6ZGqNut+nXj81jyqBFCxuvvq5beXw5VcjosRL0pjb6IE03qPWWwyINB
iJM0zogzADjWvOIKIjRtZBULdys3GIVZ8k/BNk7+a6JzUWvNJnUJ7S2FuF2eLT9k
dK6j62tLff9tI5Xf8llwcWWNJCmZIKJTe8NyWIRjSEGMCf3GdYPBHDwWn0OIvTGp
Zlucm4vX0Lz/fXvw4h1DHvwVDqhExXq7xjtqIHrqRerK7cPrTZUO4mehQt52l7UB
7mrjtRd0Agp8teMqACR51jhDBGAV0qhFWccsNe+1GRUFEgAKXVGJQ4fHKxjVF9KM
GGhopiw5YzbPrRdhzzAofGiN4EN/6sKqMNoJluLDLKly6qe8yFAXmVtCHplW4VVm
3jG4Jq/J3VcEt7fLGiz2wDP1NSaFzRJ5uzHDCAq/Myorqgk/NUm/atmivlD8cskt
S4nrnEAwyEowy8GYiR0kIo5Xe+CQs8XZwpZ64O2eBnXiDPharvXjcCRMrtTijw9S
lFifOsfhJtpG649BxOJKplrVx0RvREuylPfnsSZ8v7QWriKerms3AoqeVIYNdC9y
F2Ck/RpKrzM8w0ARhqIdcVzNmk7Y4AFYaJzguFtuEIH6j8ynA8nQ5NarX2RRLkDN
2TQVP71fkQjw44tUsYKR62ZiNDPJ9pQp4oP8w7pYD14aKBx7IoFThR4oeQWNoIBz
MJsDAzhBXVGKGF4SnCs9HylSxuRSa/+9JOXGN/IXz6Z1KBSAZEWiJhGIXGYsohEw
O2MYJDtczzmH/NxHcBTMmFAiRT4Vkk90XCpFWs24fTmoi6ILVf6XXsCBK0yzNnhI
v/OczghdvauNJPFP+tOTEVuXEGmq4UWPXw/dHk6VC5esd7NEmR8ppKYp93a8l7Ch
a8sxXKWpLexUutsseQV2oHP973AV+6CaXS6bO1hIh9QZ62unBWZM1te0rurV5tPv
MjCPmZFeIDx8CQFmdNmPgZZL/0bN9uyzz84Fp3FPl7wIZLFVJhooY8f5Hj0uyp0e
3m1J7P8pTTaQ38X5lZafVzKuRR5+XS+yqBDbr2Y/3IyW1QupD2u3TJHOZtwQsW0+
J8W+J/hgN5Gl7hoY8wX0sbATvG5H7oYNzibZIUEjuCoSuMu75ksyM9hEA7Trsutc
6Q/8r232AWVpJbCL1zw0T1sR8C4kWTrXeuqyiXIMUD03rNmjpDH5RRqxUDwzWGmM
zQEkaJEx2u1wWjHJUZlvyfwa6/Zs/f3WP2LO5NiLLANd5XfmuG6Qk8RuJV1bNWwJ
hufVAJ7dw7l0Zl95K55a/JJkAnQW2xdNW0qSGeOgP6Arh9G+a78geTLKsehYq6vZ
WgvjFuHLtsqHwUnKEjum+60HIij4meA6kmJYoR5GxDs0XPMObTMUYqgMw1eCn4xx
h+9Qj92IwMAmqsms6/oJwMGYmglIK8iJ8NKX+GAyGy5lc1qrAyD7fn8aNhmqftba
2HnFgFwudooPHwUHyOL8LWnxLSZtytOj7WvdhdLwEIU1xLqrVA2vTJ0UffqvzeV7
QXB49rbnTM3dqWXzG3o/XohF/Af/nevutesXDnAl6e3zfrrHZ72vD+494tWkiy8g
zvuPFqLe7Fca6+qb7dGLtktRZ/u9vGGaxPGVE0xn/MV5MOQKH/vE/KIJ6KEtkjBP
t2EUzklvNXrn9taXpP6M/kENRaPvI7ZGzN3m0ZcEFtpMxrSuY3DPs1VfMswZkheR
sO4oj/l+8rXT2lLH5k+O89AfZxxuUxnPVRdBazNs3yuhvgsT6bM1663DGyXRbhEy
FRv7kDRKsZ4/BpV3ri3GSY9pCQcSgzI4XsJYzRfx8lew/69llP/ecGv8fIm+hNR1
Zg9ppHH7hcoQOnp07ZYiRoE6JeFx1M6P9lKYfX07S2rfft3q7iL/dgMh77tkAoXQ
gFvMtPwpQqq23cAU+2ykMVlNQR3Nba62HCqkS8uu7dd3zniTMloy4iGOvK50RKBF
UWvGqBSSauJtV+1pwjTLylb69dbJiBgrWq5NNqimtrosd0NpefXSYg3tsOJWjp1T
zqGoTiqpe8+rUFYU4y1zesS9QGXCdVae4vsH+AsXEtfrVPtJuaE8KsoYzJagjNpw
3GI6d4WNGayDY9Gqk64q7n+weOwf4atAcVA6tL4Itay+s7PtwKOXM9ehQOXnMyEJ
LL/pGtSI/jWeGT6MFzcHCrdvUO/ALaed+/Wi6iheuG6sp7PuHoAfbtRMGqKsykea
Jys1BQBsDRawDGTjqUkfFo/PMgCwjNgvKL6UKV7J7wO9YLUwFZ6kD0gpvJBtWqI1
a3HiZWcMjV5DwR4mxruOW3s3U7/IwS8UHwaOnpkXm3yf2NAc928P+OlX7wYU5g6R
lQR1ISNnEF19UUO6q5rYfRDH+MuAKU23XcJ1WCRIipxs6ZEbRy4/K8rZ4J8bEMLs
I21HWDS6M11D75IehhFlhfypf3B289BD2DumMjR/Yle+VCBAVYzhECaiFeb1vFww
b0fmvJe17PfeIna9ewtoeNCRO3wet1WV88IenlOiD0UVuWSTjS+88p6UO37yLs5w
CEMUCYI3NdQgebV1VOUsZrMMzZX8dNrGUhWWk3BLNiV8DGPthPQA8jdK37sTVTjT
ik/S7sr2qc7o3SOcxUk2yqxDmov5RoK2e0t/JMvOSPDUSrt8yy7dySBIbdi++uqC
k2sPVL876si4IdJxC2JVGEWx+ZP7OrZrSBikuMrjn/EkCyZS+cszjYayMxrbJYjI
4ibHOqQV6gUOIM27W9d8kCVK8SVYNHIcbMF8ExmewJ8T6uNBBc8vqKLXQFy3d2Rz
Iba3r+ywo8nl/FToAamg8ePYKDIDT0siKtiOM63yBfG0JbPkRGpsrpTpAsf+kpAQ
M1ItyhCdkwkEvOYsp0fy2BZAVCWKCVGhbVavvLgLw8J/APqZnUvj2zCrzKkpK3s3
hvLo3lRPr/a2mIHl/bbHD2VXZpJLV81u2SoewqoKfs6apHnIme0sSA4foz2gE5JY
2Y3hGRIEj5/Ri6spLM+Xgh24kHEgAdfy4AH+jZB4SWnYaEV3SZhlBsBP89kBFGkV
TkMXCXzpvM3KyCg27/VbGDibZ2lT7Zafpq/A9MUqVaiRMclgBVc1u4kdwXiPogCa
RlQvLjJxl63LsRQtWpeyR7Vw/nwTvfJphI4GmDrUB93H11Ojzp4N0/17DnNJ7rS5
BMr4YX1+pnBHvgol77UGXxvDrILCsoXqBOQV139vDHHzqbkGWZrE1J32pTzO+XT5
PLuuYhzgvW6Y2rbveIdg/IWZwxu2db95Dc6BL+O1pN0EmHVHNGL5RVp0+tu+RD5k
jXaB0cFJWSvuWk5B0YVAtE68GkSco8z06aYbknTFRALBzYRMjq0LrdcuGTyOCf4r
qGcH9ZYcZZFtfQ397n1k+9xpsfCKyATP8/5Nlku3oS+UPo+7dTyCo42odQI5VVBN
kNKRw7IUr/mIO6mwjOzM2S+3lMQ34umfXal9GOlcxBGvZMI6S1aTPrNqeaLF05LC
v/+rm5fwHOVlc4qcRLUaUQa/neRjpa0fckPF0+h+MF7lkiSY6fFp45i6Quyki8EB
ZwvQkG5tExU2PFYCpltY2Gp7HBJ5vOxriHj//Qy/tPx6qB9Of0nmHBCB09ze0V5n
yYCcwkpk/Z4+oq+QKxA374r2rlVu4izl3/+TkobaZY3SADjaQXy+EdNVXz+U1jwX
GYJR0sjgfuOh3JkQyiyTDhI7e6xLePUD/nb0n5BvydkpLJ33Y+m5w6kyp8qYavnE
ZRp3nw+APHQ85fxVjznCVwE+IotIWWWl2chJllzo0++yMDqjGFM7RcbhkNoQzoFS
lwnlEftnV0MDJEA4eOaK6gRCxvGRpA/Rafun5Kmjlckr1MJKRg9ofihjbIzV4Gc0
z21S4opgxTIs3qd5p3hswgdNPt7oCzq7Jo6N7cov4UpUoKR+IJeF2LSLAfFN/BWL
p155EJYUkv+YpkmPxbjMx07RrpANqoqsVgePx/sBcsBTLiqvHeqabNGQJ2SA5vVL
RsjHRtBBH1UV4hz2gsMX1CvkkKgTrZD/keVB49S7B0BR9mtqslAKFMOzAxcooe6/
ZshrDsawhzJEEJ29Hqcxz08Gnqv/CIc5d5DkBV76mHCEM1RIlF6fynl6FWl8DKSQ
MUVUBafyg9f2GeHIvF3qMCYQN7OOl1yNC2rB1X+foO43m7VxjrAjUEiurfv93qHD
NwtkeJQX48qcz8yeLTKeBVauTp35gMOyLCUixki0P2BK9VyCLVWKNmrUcPJ+6TmT
FxzD2rgb0faDIDsczAsm9r3QoaHaQms3/ezOdTzuKM1oWHErH8QMeLaXm19b/U+/
xQBtgkYfN3zhk1J6pD6Zvqzgxb2ydVnq/Z9gM/SQgk0AVRTcC2H2lTSJxG2B5+GM
JQVmz/joyBNytzRfPyuQfaRimUir5qKVRoBqfKFDOWDhM+keNilbRP+8GSQnD9ht
pVrcDhDolwaqhTdkbpzrVkZJ9oMjLNXnVK0itZSQp8aTPmw4zPfMeuCar9+NpRPz
5d1ngK+DfiBfuEqjtX+Hrk4BhpYIE4gHuKvAfJ9Enel3MYX18JR0ZEqUrj3Xv11W
oNkA1oPzCdHZusahbukpfaKUDCjuqtB0B6+nvEyQwgCT82fKDysm7vXtHeCn9d30
M7eK0O5MQBMVse+OBEXVXeYUeF/JWDU9tX4/grF9OLHIclMqIaErndTMTQAm1JQe
0ospedI32sq7il1HRYFdGZabl3yeAUuQCVJTHLCmZHHuEcdjCccTd+BIpseUZmgW
bSoaTdidU/wAKuZULkUkAfNzJ3+LEMLsJl2FQDOZmyAbGbjAbFMSfbwgDwaiW4pr
jr3jjWFjcDyEun06cjm8hAHlirng4qEQrlI2tmEUrgKeAsAlXVMllJ78FyNgTsXx
IxORRXupxJMfWGxGVRkEPUOjbyc9mREnEx0C5UuprYTyBM39S8CC/c+Sj5em9+g0
Sy1EroFgW8+kubSlNjEbuhiovXbErWk/IEvE80KLmS0LOE13PKHXUaoSKg1vaLVV
gsBnam3rXqP4Fcaov4FlkZQ/yLXXlTkKThUC20Uf2LIoXn/lUW3RwYxcG6BDzAUo
alVP8UGaLo2y6/O90lL4TveAsHoks48riydnDEL0plKTKQypVjR0WI4RqQHMiAEh
fjJABDvz4f47sbCD3UpB7ADJub1t/gBfsfRBB0LdA9zkRtHmC0WqBcjLaImMJIx8
9KjakntYTAXLJ+gxLARAwv/+Di+G7wB9bJI5t9vWOLHUgvYEtVcqEhX6aJ5DICf+
866EnUYFf5XZmL302dpbAj/qKPLZDlhaB9l/65PileubQ9TIIdnfHo08xBTV+QBa
DoHZ5QFp3v3WStmES1R4xPAcp+Y94frJ0TZ+YGnq5FVOkY0uqb47EFJ9SCqnF2Vo
GWBom/nkeEhX/iYQw7OZUkGdJZ2nC7pP4IUAL+Rtp00VoIRRu3aIBUbIdFJayGIN
24km1jlHP9DqlFE/DGzh0lGY8N7aFEQkA3LeBV+PoClNT0qxr5JoFhL3hIb4QzmF
WAw95dhqvCuaTq+p0wVocjV5dOVIwRW2L0zCScWlIIrpqTaeHAmVPjqYno6iOYAa
RiEzTdtJW/5X5oQ8+9gpxzhXr6TlqO4783aWhihdwmHqq5+bz1n0f0ReijzNtOuS
cMuhtLJLFlnJVyJho9gYMpmiywMSFhaTssYqOIDO24dpfYzEsQhrIu0+jaW2QIc1
q/xzBENGy1uW1ums3Mdy68sPJp0FppE7h1qsqUqSrsLvhlK1jRztrOIRXKPqDUhf
4YqrgV4A5uxb4ROUSlkf9v4HToBKyLsjEaqmLljVrpIuGEzll/IZULWqKITGQKVk
7mq8Nn7TJm2nM+pKKKWJcynuaPpAE2NKVNnfzJWGWK6Ej9KcdU7V5svryTxV0FQy
Ikal1DISU4onNEJkvTB8wQN1yCBShvlFPm0uTBR/gkTkg5eab4kX8PfGNkg8Bd/0
H4yPk4Rd/HzANzh+1EmFo1rMRfo++hphCqN6LzOVMI2qlQEOGJhQ8E3MvHgB0Xna
1M8J4oHLQEuMgFDnXF7FecEZjXn0wOdmHqhaw+hwXB1l+nSIZc5ByyzmShZB0WGA
K2nUm+bGjeCkUREkw/2YJEIEenHo13GX3nfx7KGSqybhUk3TIXjHQAuE0TjmG4BW
JG1pMxZZCj4ZN0xoEYvE5Z7/wAycVj/bLu7k3JPA6T0087ZIQiOqHOzi5IYOX5+H
GzewZIcY6ZEurdbZ7vkG3fh6IMV5Oliw7Euwh9A6edSsNaEKDqe2ziTy5vZfl/PM
1clh9AH8Zkv13+5oJ4rnAgdnueX4s9O0oYsufLl1IAidlZZCmhJLvsAeyUttTGpJ
yTj2cfGXPTci6ZE7uyEDlzJTCk/zqob7IjRqngekOQ/8w3+TdsDW5n8JaicPlCVI
UFB3hZlN6ZoeSv9oGTOi/eAKoqVoboHWgoWl5kmBFVoTmCW7iHsQTBGzi6XZsyIa
i30GVB2wArF1nxoR9cHdoDwS4Ib1z0cu+9Cly0sb9m+iBIo59y099QCOn1MNEpGd
uoL9l3vu7uZ72xCs3uWC/UZMN20MLSChXRRn+pxumHrrscoPQ0gUobWmEUCqKF3A
jLQ2ayx/oSoWyOUjqKyLMdgaaLDpZrTZPxKGbSH88XpVldOV8amwRtaT30IRDLFp
Ty0gsBbRaTVU8UdbD4vrZhEX9M0EwcLX0BVEoG3F2Z2SjLzRNce7HrzFRhXpdCtU
LAeS+4ksSHxz0Fi6NBKICRaziWYfisolJnFPybOqnufWfOf/OzvhTn/ctEtJ0c8L
N10pLuVuznphgweSb18n3tFegBHgS9NtazRNEg6Dt1f1r+SPBsyafXEH2mdWOGFi
GhO/MmEPaLMm4NxRTfLMlq1gcplnqVH8nfaytxCuexZmNpIIK1lhR9YewVv40cL6
fcyWUfPalp4yItuvU034jG8thqcNQ8xrwTIQ81lYIGbf9xem8yZPlJupo11Gx7xr
nUCATj0HOpxZ7cxUvrV0kgHfIoq332tk6h8aShdzJkA0/Pj09TrA4KaRBJb9U7xm
Kwz456HtNMiN1UO+WWFK4o/xVmjYJGLxk85H3p2aQB+G77U6KfKY3v0zKLfUAwwv
WKfbpoRbIJy7CvMgolRDzo8itsvRIdosQRRG531/dDjoPdraXfUys3US3yTwMkbx
lPP1hIfBMYnxnLCbn4n7gDMWVZE62zLNshwcSV59mafWPLM6b6tkVCmBlbhRwW6R
aMX9+S9sHOfnSeQWQShsKFx3BXNYr4bhZBNM24oPcvu4rirka8LKVrFaQEl8E7sJ
P0K3walmK6FIT0QUVEP3//HszPct+W9aQtEl5Ani2naA45uvdsgo7K2rwGVTo43K
C85iyC5e7dZX4E/VxjC2hBc7gnVB8OrJLa/omp664fKFUP8aEiFYJjwDx7AeN1Ll
1z4ZBN0UXO4/wqPrZI0UigVusQ2WyS21c+yxJJLN4W2KdVKibm+QX3tsC+JIJyOu
/XsGaqpw2OPTG8OoNl9F9gSZkFn0cMn0lmrqFLA5D0TpnQu75n2MJa7zbnaQqMBR
12eyQId0ay36u2b8FE0Pd6HiOULzrhod3ljuIyz8QdMC87inQb+W1PkU8mpe7FCC
ZqlGw98E5y1yhXPgzqj26aPk/gJpY68wKJ+J9bjft34+rozERXDkWXllw8BM7jAr
S3eZ/Yx3hwCXbpOO25rYWaB6AtEDi77bY2rFpLtNhXT+uPFOLborjYtcEz8/3G3x
wuOam7pX9yXYgYNg0lLTvYw97IfO6iR2CJjDMjQ5qBS3oC6f8tFAEayGLbKUsQza
CB2HE3W67GDyLpgODJ396K+pnHODvrL2QEqRHskDm/3P+svp18PvuctbvqpnMatc
i+Z870gxP5SrLWO5yPIag1s2jmxc7oy99+8h+efNNuRWUybdMFUoE1OQsjq4HGSj
PlYU9xnoQa0Xg4X9XZDqDPBflrqU3wh0w9pJZjd+zoPmihPS4GYsBv+DKc7o3Cs9
8ROOGexJuVJ/MXZhDeZHc/GbrWBVvnEvW6khlSTfuY+S4D2aYfHElEQtSdVglnfG
21J0M3/LlrI3nyeHtAZuEVdf5WPUTb6OXGbr+76nT+I1gdIpHzh2Buo0rFq6R0qH
yfdyAU0U64QfK4eYmtQbO1DgJEQBgBVToQB6OIw7pNcG7hqNTBEJeRi+cO9bQvU2
C/w9mQpPqzNoTNT1bOEZvIhCxRv3gjyFfn4EhxVIaKO7QQ7zXq7RpSCeYOYCfbE0
Ea3N1pqOPsaw4dmWYyrC3SzZNLdUy7E2ZsncMb+Qx9Be9PuBBfERm62HcSygUYW0
5C59FeUDPvFM3OtnAz0G+LECYrm+qdoaxtJ8kWbrE6MIDymwLLdcnkm9GaQNjzfV
3OpFCNmKhY4r/LlpwyGk+TeYr1a9KfDE3sf45avfhoxqMpLaXPzSm/V/lSCGFG7T
s+fB//+fEcq2VGAhi3Lr5UJh5ZnlUTdw3ziM/F5RqMuyGAWZ9SHDdc+KgDIjJ4/q
BYTIzbDhzyvSIOB3/7VxHgWSPOw047KR5JUb0OqGO0/W7QC5plIvZHu/ns+C8gsl
h42iuP+Kbp/TIKf4C4Mw4+lghlvVK19RrEL7OAbC4wirZc2MHhia3y7FfpjPgHEd
XoUTIAcsWuHr0mwLGqXcyVvBppv7nfmWD7gYuhMEQOuTZTVh7+Shyv6OQCcsIPbi
j9jYNLwO7NqCYcvUKLTZzLf0Tu9sbfTD4udTRuox5qw2LcDd4pTBwJEXyKWBOlS0
7fwSd3wcaOoo2pgG+9Zy8tTvJGVtCIMjSF0+7zhPyIKlE3jr1iooYhDOyVmxBA4U
ggR02Y1rFlPbCgzprVdRMBA0c+xdurwZUWXHQ3bXjfoaqoH2FXL96JIaJ8m6e8CH
edkaH89CfwiqIg/Yb6aNw6TmQJLdsKrWZplNSfx32QBFE2eQEcvTWAY1wiqG7uFc
juALb8IaQPBC35iaFxZVtnvqZcAFSWdZAO2J9dhLo9/1pAXTyLLfbT59DVfhL1A8
zVxL9HxHjd6cJ+peooKCMJrxRfXFWeICbOZtO0VT04OYfwKMut/bzUpliaczyKKn
wYSDt+uSfvwvreUE5IcIBkqHgf7kvpmN3lUbUcNnYq7r+PNHLMV65d0tWgKqJP3+
eDKzvtbd2BSwUpJAePLB7HDTERIQW/IzMtTENS4VS073Y8nQJPwfovUwH2eTHMv6
4ePeYyYVw18sj8KEf0DkhVAVtvCeqj4MNvTN13DM/6HawPa92md17aOJ3WJCDuR+
+5Q8FR3ufuOkozzkYKUvuYqwappyg9OFGB6aWjwukxHxJhvMMUhSFXnXSeR/1arC
nz9Oyuh/rBMTnJ27YLzeWZ3KXsGgUU82VzWiBv72Nmg0xQ15STgA/YeONQBmFe0j
CECViQCxEa/ITKBPiQF8iANu6SNDz/IPxdUMS5OPErr+elSNSraLEhUfXjq8EoVo
jNcdhuSc7YW2QYpurnBtwtsPKh01rUmHVnVDjH498gWqezBRQ3O8t1fdjkfQhLTx
vfYVx/KqU2GufnR/0kLKSgapS/TPM4/03vgy04+fc/Sr+YkOP5ynYF3ZgrB6EXz/
mu5NjC0FK6rW3huzeTBsMzBGgVNoKS1DBG3xbvzPNAGM18p11tOIeOAKtwtqR5mi
olXiHcfQ4BZ1R49MKpsB4IHlmHzvRkX702ZbzBh8OLuXYqlWCB/1NT1UchZ56dIn
LiJ6WHGtBVqQlvIsIWfHjhMBpwS6jI98dqf/dRJRcX6O3Rv+lge6T61V6dodvM5L
Wl6TC0s8prD9/TMX9FyPzyBEalQyetqxg4sDMh7ZJGGTRAQTPaTkZDam07ksL0L0
3vwcN1C8W4DO5sm0iFOOccwbr2E1wDvgCI7h3emrap23ARxwqY1eO7NFGJjbGpvP
6mishflfTCrNwdRpp8uyzs/4KQmhZdGAGZA63toEDdMQpA/nlzbNzBYRvETmiUYE
70iEiDiIq/ic+7VqkVY77hldsDgg5JmAHCYWTjQe/0R5kEESQcxbuPCUA4qYcJyk
ZfA8eI0P5VPwdknvsebz7YZPRd0FLDBR38whLrM3kSnzY87HMszUdgwDlOwwuv1I
jWpmKn1C5WrloOf9a9qONbbfPEbr+jlJ63U02852O5mGrLNRgUOvmBkidC1bVMFy
KLIdxcHmCDjdi7LmW5ed1WtqOh0oz187zdzpUE1Pqu43/TyCiYLT4jWMMguh8w1N
9pcUUBybTzVLY/0JrfroicqwZ/yl/wAylUEg8A4b2yOlunwOqE0gs8QORIagACaN
qTiMPFyNdgbvHnFejw7RdJBGIi5+K96pFIt/mfebuxEZzgp25/9aV9u2Mt/k8OCG
8Fm7HsQxLsjXHVPZEqnXWGc9bSXx3D7zqTbgJtyDgiO1ArnsHtrKv2kKUNs9GH0f
eVf2VWSFFLjR5d/9jcYPVGPE+4EtUwcwNCbGeAQ8pfVxQ/6i6yRLXfXwz/nkN0RS
rkgFizIT92QzT23sbWru1fKHGzTuDqHTCB+PfkOBU/kr5Hy+flRszHjrMSBXr/5B
xTaMVATEalo1cZtuUTyOB21M/irsTZTrUicFa0tBwPW/RWRc34eDUF3NlVlb/Adn
9NZ3GvwVdCx48BbrJykSuyP/rhYOOgTJn6wgmwsmabrEltwBV/nl+RM/ujftCZeQ
W9pOQfF6mwCwZEQltEWLSl+pcPSDCrug843OksaWU3CHtdZaEaoDsVryL8SL84dD
maJzJ1gzwjikl1yD/PfWEgvmOGrJl8u6FOgO/H95w14noItM3NJ+XimFCTlW2ppE
kKzUmhIOPMCkz0MFsXDLHVWSBhk7HOUi3L0qbhC2Olwj4r4eB9LQXq9PvSs34Wo+
zccurYl7z9IfejjSV9Y5mVIdc+P26ed6VHM1LEs0qIBezV6jmf+lm/M/8bgHwPqP
T+S6Q/lzIjhHgfGFsiLO4VFVkzLah6IIe549EpucNp062Bp+o9nbZfZxJEAEs5xO
eoHFFZUGFS/wqMOE5lSbJ5yY91HzyKikG7FrWElihC1vGYikQNqnmxS7KlFP4lgF
zkPTENqkwurLWddy4ASi4El9KGomNo/3whSAuQNFxwQY0hgNYJRwHSoy8A3JfDn5
SHKowxOI4yjdQ9xQInla19RMi13nPbUjGc33JD47d/f511az58HLgwbmNsu1k70r
vHCPvFNGwdIQfzN+sThJc76Etn/6EzW4jyeT03dmfDltLzvYtBiD9gQyiVr/PCaf
PfSeLAlObIj8DlCYe2m3WHC+WzoYRPG9cybLyJJU5nDdabiiKu3UxOEl1Y75vHG5
k4dANUy49Df8uFttC3lwYmofOTXaYRb7EYelThG53JkbHxeTl1auQjLLjt21F9ds
Iia21KUcvstynZpIocWjm+3ecaoEih3o+QbjH5r1eMiV7ysD/cilXu9ErgWbYSRz
7Ofui13tvkfZrAIrLTdhvgSfHT7xnuKK2c9Qe1wsj454TMD8nS5eW/8hD4M+LhKi
+pagr18YjPJ/LLvm9MX8Or1SdBdWvDRrwrTbotLqOnxWe0IWSjpcec6kjamYktiS
vpwSMRwAljbKT/pQ0m0nV5PWgsHB3+QBZlE70NdgegxXIEzDJCWiSN4w3qrXoPQc
eKEYV3PdHRy0rbgL94rclLxY81zUcF/ojW5lH9XJ/zf8ftYJ2Hqmuwgt2HTXZQIU
cpDzx15AfrpZ1cbqunTLGOkWFh0eIss4Hni4wDjt/uTSZ1HOWpTZqLPlAf45zvLV
WqPZtsQ3bhl/LKlcUBayKaSrMGBcmozCWdZf2Bzpgmo6Wz/HAaHxWtKsA4I0aV/2
xPokU0KpIo/P+qPGQXAi/QHUQBBjOHvwgB322M+P9AfvFYvmDbG3/n/i5yJtKPkt
fuRRpiBJEYpD6uJIeDheVHKmZwW3jDDCv/6GgmcVqs+V3+74qwQlpvV0F/8tlMu3
JQWFv2ALkDpbtQv2/vbIgPYXrQQ85g1mHUykoVuykOUM4Ou36AhCtkZ0E/PuFYir
eqZHFOM01VVdmLyrzu/1S1x8i/2/bKOMdYIR4vYPXJXZ0MS28qTmHiikrksr1mrU
ISqUneqLSkCJmwI07feeF/dEtfGKFR7NNBZz3k8L61dgxXroQKeGG4e0TQpMpA4T
eipy8ES2qgAHuIrRAWZokdvI2nQSjAukq3D4z8wZ0vJyqgOu24IHt3Gd9VSk9rGc
3U+EEcV8ELszXQnejE8Zx0JvTQlIXAVcHpjKKClB91BkLJ3bcAPBkbaqxF8AGSB4
xw/6DbNdvkzvuGgq8RasMeGL4yoZnQOZGxu9YQghpSN/vMVtNO9TfgljV/j1vfXE
m2BVvSOC7XkFva4KspDQf4nthA2ykZzuZg7Gz8Lcz9h4qrQElC3HCHeR4XxLSxvc
D69k9P56ShKiaGk48edL/mwBzBFRUZyEU5V9pCFoP0WM1DgTxPJqlmT0FzaNXKhq
hr1xiz5263vtbo0GclmVxxotYYwmBVd4ciSHJ/woEfmZEiRfkxaLO/sPGuhFdoak
cClCR56zS75QTR/xbTLzm4f8ADHWvbIzt+tUifTizFWX8qayzIk+OXoSCkcxPJyy
N4dUIYSKvMw+6oXd8ahKjRVI6vjTleypqDPhQ5dOMEUt6jLP3wE0NQlshVPjXB6K
wYRgBWQRXcgw98rjoW/18vZLSj3H5ariGAZysKqo5AdD22cclVq03sKTWvalr4vE
0D57tp7QQ0XX5dcjvvHvKa5dAAgKJT/aOT6cw+CcJDiebGWq2nOZzVTH63rMY8Pe
XexTouYFHigx898aC00y8QC+EBiLBYGWwUo7q6lDPMcHGE9q37K9HvzqkWnQudyt
wgCyQxdcA/rDgaQtsKXGxNGHkXbOaW+OoBGlNub7HWog2LPmmf9pibDKgjqe3Q99
NHauXeZ9GG0LPzatpjq1CSBeWPJCzfySoBz2JRYT8sUjBeA0GGRFw0AU5roJc99B
iSijE7mkEg2HQVR0ycewUkDqoXRJjJNIbcKmfI1BBYOIsH/Zja59YaO5EMXOHkQw
PDheMHvzjnwlm2NC71XtTFklOnyBR5sNv1wEq70LCKX5N4UtPLdGJwS0i+dUX0CU
lKKZLYKhRBj+6v0eOae6exrgpfptpMXRgRWYNdt4ohqUDIHzfOCmw5Mtb0kumMxA
HQsZEBj53dX/E1FFgSDSzeA7BNE6fdsVRlsxkzdh2dnI5z0sWTtRM+7Sn+hUSwfQ
MFcv4+uOm0/gbdumNKEBHPsb9MunynrcCtcEHf+gzcLEcGtGScAo7XvtKqf+eNu6
1f3okGY+gQ0NyEBDHNCTtbDYQmAUNYXMF+W73HRnkezA8zswu/pSK1h8m0sBATRp
trefLopGIHGrMpl09TYpqf1TtraSBtQc9ufj8xi/PBFuYbSUEydLZngRnceeu9hL
pyqRXDwseRBsjEtCqVN/cPzQBqKNw7kzBAZE7bbT0Gd+eQdiH57K3HDrhpFJMIFK
FQ0JzTh16U9d2KiO2GzWWSVZ7I2lTE13M4tmwL4Fmx61RzqxpW5jVDyoOKkS4rMX
3hQwNfPIwNQHuhD2+WQ8DTwM/be1OIyB+HhMNMBnehT8dkXi5RRUpm1mF14tdIxR
vu6Y0k4jlyXI9sbik+Y4mPYSKUfimh1Hv+fQSef7WIrPCF+sllH+XYVWwOl5e62G
/0fGyV6rOEBk7KUf/1rzhn2XMHjlEwE9m6rFFC4uvVsnou0CRADSDff5+HdzWPlb
IcBRLqOClnYOrMfCMbLOG6xSyPE1tyyLXTiumkwxlHLagK4V5qk+sPl5zdRayxuX
u2ea1SnBoJCQySF77pnK0uMlqZ439uFk01LXO4mLj6bpZD+c8LnElxdUljuBspdJ
pHvQkKt5ZrsnB145SJkApLwnGU8O7VoLPujtFDykqIDz2uXGGBYeuKFNyCWh+WGo
6zEFLT4aTgJNqWfLg0oqHEhuxbhu7mVFPU9sw/SizPA7CmTmLLay5tql3igUHMa3
notKXhJLJwrvrxWZq9DVDgv2tByZExIew8ZaNVgUSROS7lRngCiUHxOnu/+VGGYE
k11vrg5ha0BHPkTEps3KhGANXlBI8/O5FOYCzvO/t+JiOnlGB48IVfOzx8RGlsez
AI+ZF4ZCMAp3EUcCANyvDramglZL0vCqFcwv3n0d2hHsFosFz8jBzj2/ZwrlucOu
KUJ5B9NTOGyavK6Zi+zK/7k47m8uF/LGNT5eGLHE9euMbfd8dR1f1aNaMsYEq7Rz
dOndhNdhdximgkbcCUUIr2L2ERV9fybAJW+vqrQQrPBJR5bIdY5WiD//z6JcVvkG
5Xnd/BBwDMf3KftPctatwuQyiUdhEFUdVB9+Hbbtht6K8RSYVAT/1hbAM3Y/f0r0
JMyLyx0wQUoBgjLL66iqo87M6BfTryJvZ/ssqna1Ir4/Tb0r7KP9FueLdXhWtvTH
0Vi8P3j3c+qwuQqKvt5HGVpk4hDZdKKK/F7n5F4VDPiLm8jzO/gzeOo8WXfS60R3
oDBp3/I8ciQbIu9UUi5yuBe7jZkWhjK8ssbyB6FuGcCQcHqc1GNZSghXhT6NH0wO
7dFcyt/JMWwiyOwIMLVTyPQb4rmhgSUwCxD89e2SVtIGyORzw1moiyDbM4e0XSY4
YiI23du231mR7BYqDiAgATd4CULorOYg58FZ8Ce0vlLD8aKE5AlwwEjtxXq8Kyq1
9SfA/NfKKYJKfcXift0aZLu/FnRFN3ecGQsludY8ObPcBwtT5eI1v00LWkM04Bqe
DwzEop68ZylXkAVtIsLoJvpP/Bk1LpwBfOTFjyz5KqzKro15SsVBn5n9yzKzhOUu
ew94RkP0RRRyK6X0uRC1o4ykkgyJ0ZYaoXax1OFnRzFlIgdX+6Lm9w+OX2jhcaip
fyrUEGJqK/LJ7J11hWmO02ey9dNLcPtBk/pWCU7BBpekiSMG2ViM79tVyWI+B4Yt
J6tTX93egxfOUBT1ev7oJwM4vfjUT40TyO2h9sPKngZmMwz1bW9qRbqFJpvGdwwV
q6mHqINAqBgnzocCvr84KVIYaMWnxRSaiHKC3JHR0uiQWY/s68O+5YQv/FAC6i2Y
7vdlOI8+YiRwmKyvM0LNN1MiYORy/sQUWo3yNRIlqJDiR4h0fHfX9s3+lyszu8O9
wLVbC/c1li7dRODKEvV/8NG4aGFaONxl1zHjY4pH5l0WUkmtV4Rb7Sxt+ty250gr
50SSLKNcWMb7549r8Ssfne8htVwtpAF/2jBiTAWLzo1rNcVNXKMnCKRPvOCsoLRj
kKkk0WnbS61LqfRRu7fS3y4dyrf3SPRASJ/SFdBnBA8zJNRpHv9jNQRIlzraO7eN
6DJs7Tq+IQ3a5MilyXIEeFBRdzxMFZvFFbceuvmrXVKeClBgHjgGDKHSeoRhTKXT
ljTRvCATx5kHcL09LZ1wzsW6Tzl1SGU1qv56EZPE8tzJuiFhdggvBUbsYmSWa8vT
2ofSP8XBdqpMUrOcnMoYqkjaMLqsYB06ZczFrCLSC0IcmYkCKR3pOEpEAQS+j9tT
HxnOLsvWjfE60RbsLP0tDwSLGwnhEfRvFcXkPc79aqkepqPqvo1bx/M7vjc+pDRC
6EsTCgZAQNUdfY51KVMDxOkA9PTQI9+qFIkpDcA/YN1MKFGkH8MAnu1w6fLA0RFQ
b1vVMJbc5czU4z60gQIo/Cp1WDHnL9VxMxxqjxLi144iUouw1z87vKI2rsvasJpA
5Ui/Aj+dE7hNW3wZ+bFUCAnogEk1RA3XglhGjoxSPx68LJr8MKF52dYEqmf0jzMv
CrAkSoTV9gSIr40y00jAlMHvrJeRn8auBG/2QqqE1MNZ3nEf715HnmqFTx6pPc1w
9rZzkuD/pc2LMyOYlW9m67bMLwysCQb4FTC68i+yFsnuODKF/MPf0P03risex8MR
92elrEboKuqYh22+0xpggTn1/pRWVbaI5D/tlSZaQcjq3LPxduqQ/kzGLdmt0ZoX
KW7qddKjQzQejokPjYr5hM70IzhpCix3voFyyxisKGouvrydqfnw1jvPCUvBOjMg
Bu7jcD509XjXF5w+e95JLEZ/7OY467QbmCzyzLa8QyWwaL2uZsCkBSbkNX4Tw84X
pyV5P9o8fC6Gv0qyDlXOCusoS+h+PnxpjoDLPReX+ZkQzAE3OniK1fxVGldxGc7Y
7Rdkv2ovHz2gll34dPJwMteFh8H7Zsa4QKh9OaZtkk/K85MRi/8l57hYw/JRXGOP
XPy3KmGnK8tUtg3dwjRkUP18Vha5Y5sWwi6DeVCyYr0nG+IsP4Ku1d1DRiC5QNMT
k5AOkSZwXhf7IPapMK+h1gxDU7GNxnEKglMYqxnzqEbnUos3XljH1W0AmLVXE2Sr
aYn7fzCZZTmKXvEr/Qc/SB2pqSMxFYG84hHxbaZfZNMzJshR0UgsxKB8AXs1f1Hv
5nTRd2+s4iYu3joqTMyXDLDCAX4oeuMO896hfAEUiGBoP/NMv6wb2Y2DL7wjMlHD
BdfL8vRI0zqGyg9iDGX8MMp9FvZxSKZj1MeZqQM9R2iAbMttEdcCTl7a3oIfEOXa
hco7Ia5hconw9S6H2Ap6Nt3gjbaglkMmXuCQTWW05F/iUBD/BLypkEbqjLkkJNiW
K3FEAleMQGOHkvpS6/gK7m+NNW8miRUNAhWCuX2ZzU01CylfKqsnORCGQlgNNMlZ
Fp5dt6SYuYVxCf2QDT3vzlsT6VH9sfWaap+SwuzxsRkTJKFICGcKh1Y53BVVZJRt
xDg9YuyG8ABuDoO6vVF63vAV+MsBy046/nyNaHBb9P1jswlWiZbzm/0IFPp5oiXz
TRT6Z9G8D4FWaOrmOXLuxQX9dCYFAWdCpNl66dlQNehRBxxjRsPu56zatXZDoUZj
3erh8NFwnTFp5vKlOuEmu3FIIYUD/1yTneTeRpSJ5GxgOZo6ohy7+4vZJ8RCocxs
Q6bvvySRo4Dq+1GSbUydOp4tBeLNZQAjYEFBOnfLO0OK2aDuqJW/FHJ3iqn5qzIf
8XiiN/XUeOjhYdSCqkNScMcRV2MhMRPCfvD7sj1lQ5BLDyD//feKUAb+BiW6zwVt
IqAIW0gQEu//sLQ6qhBc+vEp0iRePf72qBaSn9AmX/F03TCtrh6OLRD0qP7GdoOS
Qfacm6Oj7CsMdFf4N9Zq3zVkSXya9Xcqs8e3U2iL1o6LEybo5zwasUW26aES+B02
O224wQozk68fuVXrYEz0pdJSkn5IgbA2r/qEdAQ1R+NZBKLrGG3fmQcgeO6eNFWd
xFMBAUJ4fmOzNGNyl5joJZ1Q5SjVErw01KPT2idfCz8GDy7a3rNTDd3Tu/UuLh9c
/ZXdvS/+WnNrUXkq8ahTQrX+SX4A+IIK2uWQPIxksVgauyIBNadFVhyfaehVq9iS
IC0SQO1zA9ABLbZLwUmeF0+X8TxtWWVJO2t2sCafSVkZprp4qVJUw30ItpPYXYsZ
4HOAuEh2n189QlAZkSZIdtlNdv9D422c7Q9JYTzAh2aMqwJIocP/De3i26bVDJgE
PShxdG2/Y+KWxY7F/uQ5u7qKzYbWA5WA3LriOEdMFAQzDfKjgbhiuRAvPCz+3T6u
VAsgGzHzfyOEJh9SaGHypMtZWuIrfwL4t0ovM508337HyH9Q5ccY2oN5rzmhUTcp
qx0887ccMCK2gAhcaAy3JYnEmmMEk8/qD/zEQ69MAchTgAbk30VUOhgpjz/dN39F
1YFTTzCUPxRCJM9oQPQkIoIi/PfU30T2NsM8cCXiFPAWwrsz1hQqnw6JhWGnCBx+
MX5qOzBzYTHjV6c1JnsxtBE4DbfjKcBXznUkltvBefLKP5pvBObLvYkiuYGKpTEX
LtQeGqqJV1SbquEIHCoUfH1H3Ku2kcEXz4JKVJ7M5D3LmlDYyoWOngeD+ZJwSoOc
OpwNMrdMHWALbk+MkPRLj5HiV5WOOurNas/ftv6G919jmp7dTAqP/EMVmYsTWrvB
V+noKlVM+nHUR71Sn4mGz81FYTsqibE4xezybkQ55+Cv9nd9tRsKMefOrCBS2Unx
oyk8ASN8Mebu7qIlX5BtD+uQmMUuzeMuNbDXj4c7DknbHAem0TxWPyYFH64QDVwU
fVWg7jM1th0krfrdfAueYRJXV+m7RoKRvPPMx8ow4etkUEawFE7kn5FgjITKnCdj
uN9dbUeMXbDCpIlPeMdgcVjQb4ZiaA+aeuV7WzSMj18+6LMuXXa2RKW1SEVUfoxz
XgD8BWZsQmiElb4dhW5Q3OkSS6wKlNYcy+KCXPbb71GqFR3MBxJtetgZNDC3W5PL
Mgf3TtS7gJ2fEt0U+NRg2LWK8m2KHiNrFs0kHva1BLv/yEtWfGlfn2UPhwoZqTGM
p1ZpvGqrpfLym2zAYKqnCYwOvv9JBLHm42VrqUZ2qwuXe/zwmFZWM0GpmLPI8e69
aaTCqCeFPBAl2Vjk2FGss9hnXG150Z0zWspr2K+nPGU0iLjp0NRK4HtT0AbZV6Yx
sN/MSf+tHtQn76oq7SIBYtEkt2BMPSrO0tZjZk8E52dNETvWvN6T3KjFFwDt7S9a
FQSsp5EnnbQt3nCJifzGfofq9gmSCvDAe1/iOANXN/o24JnvsvH4yxfIcLnBHoxU
bkovGG6mO6uRPGVhnlVfZ+zsT+TP7j14RhwXWOtj5U9t+Ms2Em5afSbx+MfQ1Jqx
/YXMNOYTEDrvQRYI+njKUpPsSpZInwXyT1SgDA0BS7BytroCiic5ZZt7uVDHQyb4
SJdoZG84mvsSdoySsnxQVRuX6644mHqf2UUx+Iul63EKr5BLVnbSWjKII1e4zHt8
VcKPF8raFAY78ao5VFZ27AWfRBxDW1GCkZR5FwQQ5ZL42vuKDxv/LpFpnGp2/f4L
qjDqcjXNwBLjbP7JSTdOMpX0CtoqAEnBlM639Yz58P2u14ipuZJQVk/YVYFdQn6n
kR1MPw96pXVyILiGjVxzE9Ku0BeU/2eztA/tcSCIMOdoIVqVGXuw8VyU+aGsfp3A
Ygh/HyZD00pgk/9xrEr0//mcYh4XzYatQPzT+mrzvrqtSXR5NSm93G2YjZ4ixeuh
EkuqVgUfw12wNQAElIDYCTpnYJ34HvpNh64ZMCro0yBsVmVQJW375SmIi16147a2
/UJjwpT5Zh6B5mNiIc6ynNuVZwBE9KoBt/YFt6UBtVpopyWlSxXPttyvhlmXp3v8
8dBpGaRRYYGb9HoFHyTBZWEtW/RFYnjjXw2CUE7KwCcli7wytfUUaQAAEUaUI05m
iAUVLQH5svo3PGU5QjuJXWFRgC5qwJQJg3FmZgV6myoG04mN+4t0IDLLt+7UwcCG
EmWiRPZ+81T8oxs8LfoJL70vGwfM4D8T7dhMQjWL89Q0JZKpz+pxPQRtVeQxIAp/
Z/HFUwMF2h05nXe3ZJaG/gGz9onqawFQ5oB30FcIJ8RKlTcU4EEYF1NqMN88BuQX
1J2kcQ/hKZ0UErdSm6Xs5+JoTNfO1BeZDivYOBHa0k+v9b4QgZ2oDm3NK7khwOI1
+IA/+ws16mREzj+IzcRveN74jilCOWO2PHyjh7+7U0tX638WH/GI/7kyNtj3W+BC
uWk500tOWiJ9cUSmO/ON+hkCgd52GlIzc7sUBvGFlJI42s8Sgw6lmxxtczpMmSul
U8UoNiMozegL9FmG6HBbXxn/ajA3pGUf0ieoq7L7/7wzwv1bCbq5P8kFyzShZVuM
y7tmkTRyDdH+DimQbgqk6ou1Gl5Qd3ATM3IqHnzeWHbr00HxPc3+BznsGzDdt94a
fGJ1CjwRiiswnzyPDkWcM7yZWArT6r2drWCzCaxGVyofM0R5ovGayuysawayucwM
s01J7CnLZxhHw2aQuiblJAiJ0r809dPNnXgCpgJa+l3qLWJB/kIJv5JGiOtltCGJ
A0ZmqhQ3BYKpsEJEZNrStOShHSdhN7p+NuF5w97DzNxlI3LByOc6r7C2irbzDhJC
+DqX/Jap3iU4mjXVwOEPCFMetnQf5v+ijuXwnUzHqPbBKAU+U+uPcHEu+4vJtl32
iXHCHlAIMBeT46YdWHlt7um6GBpvUD+f7vCKKa5ccwAnK4T6FcppO3W+47wtFsuX
9gIIjk4emghBP1NNGscQsl2dG4rWJkrVTFO6PktwlL7f3FkoNBgSRkT1D1lSlQzC
p7IHb8KcVyxoKhUNHAkcF5AjUl7eE8pWpHbbrbdHUnIfoUZSdVSYLRvuIy87fi/C
VuUS/REPyO2if6BotStSYTolwTABIVAUjl5MFg+JWKr8CghqkSzbMjsCndtGoek0
9T9Tw9cvbk3SxSmkfSJScu0r+xS+08DpwwuEYCC3DqqLWHrz12J7yl+gY1/P1v6y
1A6OffAtl9AQ59PCWmp4QjcDD8TKaAZuH78zMaDnvmHsMfD7TVFF/i7S/d42H7Sx
DfCS9QyW2Pan8bkRzptgpgxts/ufSk9wishTxicIKax0oAK3DjJtVaA3YshOyoW6
ygYpWeIbCdohf8HG565zWxkCztBUTW4fGAzDee4c5F8rMQK1PG0yBUIj2U2V/3az
OWSTFWsb0+Ut4LSTnegLUQ6PZDBNCu6CVck4lfef5U7Y9o4/GGyItGH8UR4CLj4P
e8xx/DFd7YA7ylTYzcxWpenpt6u9VUIXVvRkoptfk2hV94j2Xp6HrV386TA0kpXZ
QcN++BsvYsJY8wxVotR6qIot4dLWgAVRHdKdumac9h2BErJAjpKK6rhbPvNmmBxj
yOEqUQPB7eeIihBl7NiyAcPhZaZI9lbq6DePel2jomRh9VmOGvZWhAftWjf/Nq8h
EpX9YfYLVFnqVtGTS4OdZLKCq/E6DZTD63Op6Wnh4oJrCu76sVzgLnA8ToKSRyT6
7Qn/zy+XInYIYqv3QyBx5W6Fq/PuSGr6O07X5dvqyNb/s+bB9knRa0hf9SB40kJm
5DiSqhZyik4Jx6KL7RxAN9W9eFu+PQh90mBINuddESfSbnEojo5ZhL6Xaqu9ICfP
aYqhZQcaNuP2DDfXEH2sFBJiYLAJBGzum5fJsPLF3Q0Jo9KV78rZcZq/iZS2YZSE
LXguOHsmg+er1OiwovFrtWZwZZY2L/vwcjYH6ar39rcM1pF/0SLoyBLtfeC/t6Pq
WrmtmqBtrlz6kM1kQPaB4ocyoel9AxjUVsG28ZoMGbLYyaBVz2wEOac8W/eRhRgh
Me3mj1mqDYo4aEk9jsnLBxQUeKpuUgSXOJ2fxhYWChuViMQEGevgPJm5/BHWNmqY
VZ549AqriLGKcgFvyql/1v+dETmq/xRtGuUCX15/UWzbDEYn0DEjsg9WG5wOELBf
rBShUBlHAX44egWQQQdGS50UJs1n4YeOzYlr9VAxhT3wDuRSt5b+55hRpEISaaof
LcDXhro3WC9lefyHh+M55w+WuuLLN+0GwtGolWv7RuGGCt61n3EQ0gKCOqN4Gq2/
kqCGmm6fS5KGlCEewtz1xO7Pm7M9qrlon1LPz3LZTlNTITtKfTmSmYdBVAGixJ9e
uwxCqljOchefoJ6WopNXHXp1jMOM+QqX+BOUJLay6o63f2CWChvJ7TBuJQzVJI8U
iDyphm9sf36Y7nhsZ+CY1h5Eu+XEszt9N0i86VNGy3ZOker2GR9oQVDXWDa8nk62
B57OmbZ4RbJRGwuWsF86Smd7AlHseACpEJmOLw07hnkrPWeje43LcPmeyMqXBw46
YezwtbAPcaAf2SQwz3c5zRoLAbIn+bi50doSfOPL6q/G2U7g5D5Kj8VeqZQGnMmi
JGmzK5/SkuobxC94ilU0rPoRjLIUuNOwQdQwtJdksx0eLZwp/Ey8gI+aQAISqmJV
Rc59nbl//ecj1nH+FNmPsFjZGQbg7W4Pmp5oc+ast0CS5xASqmAhKWmN+qlEfumK
NRBQQNGVANl16iKcdlRUt4zCJmVjra9nkhRatWxh4nKWV7UzEomWOTQizpjBui14
NraJJyKYWm5xUIF28uIu5WpyZJhZwZxySaJUIG7dX9c89akRVChHdxT5IA7I5rNQ
kAy+q1uy79whBZX9xUgyyP3hQ8em7poji1q0NYI3MeByy4+3pnD9OeKQIQJNWKai
b3qLWZOiowSaO4tnsyesXp6D6FFcDE31EO8jOT+8k0y2sNHJl5buHSai0fRD/HVx
3onbF6BrpVgox8LFU3eSyVQxEphouxCW8ud6JA72O8Tq1gkVBfgPVwFW/y+rrazs
iZp6UlPRqdXmucQzswxYF500ALPVgpFN+M/yOk4P2qmF/FfaXPNMOpKN1FKmNIWf
Joi5erY9G67eSFeF7m9O88sNrBfu8QdbicvLwPvhphcuUS/BnhFMC4LSORwIvJkM
MWMv1ktqWFWyzpusBn30YgruMfcovDxkncF1qTP6VjbJ6YzPYZw7owMeq6m/DdY/
FEUzgvO0FGvAIehgQ7QVaygTL0KzhqliRUAKX0chisBRrgsYvElp1LldS67DhsIZ
+iw16Kx3muBiET9bDMUnAjZKdn72UqRQucOeSkmeM4ULLyFckQoEeUGhDppsxVD9
RSg5xsh96+aRBnZow+tMgAazVDs5b/I3N4xRzOLRGsEFEb95fxiNRCg/C2up53SM
g9m2sMNvyqUeHgEx2/tpABR+IogxUmkhq2dWVdUiim3TDE9sdnVVEZbjJwFjCh8A
/E9o5vZ8C+2J6lGpGwz3kF9xUx2oXtEAar4J60ywDOOUyR+qKpC8xINeaeikMclb
cNy+TJJRIlYjuwmdjVGa28+mIGuCNp4kZAMFcl9FJedOGlzm3veZqAhM2dqZz6ua
eQmhZMxxQyDpuheb8yEgHlg8kWj8T3w70YXomH208TlNz2Qj0J0+RSwz3U+Mj9Dz
5IKzzx3tQUt7neTNtpNW8spwNwzwWxBJ0MkoTXs44kt4GBF2fSa2I069Sv/uFjqD
Jy2Wi58QnXh8hJHY21718ggONn6xNPRRBgM2ZSOxfiZt3dFeoGrVnSMaCKehvMrn
/bMS8f3yYclEtJ9Y816unxbKNLswkuNj3zGZJ8oIRn1tlSqsg/q3It0DCMI98K3d
7bPDP1Peq0BK5Xl+CLj2XDQMjsJnqGi/YLOFKuP2v4VHD38arX01DqJKTcRLKeIY
k5/F2NgCQcCpqmlIA/Im1LeYZU8b23DSGix/7yAsp7k8ulsLZCyqxsyfI6AyZ2Z2
awTKiPu8gsMqLCQjX9d98XeqngCA0B+ysELw09NY4cIwLaa6kZJLg/m1E53KdwM8
UokCaXRVYZ0DAU0fUmK1NwSb2rAMwDta4Zye8VnE+aCVp1i3iHuxleamZ3gxN2S0
Fo0QxC1l4BJOSWTFOVLvZ4W7HnlowuduHM3zvARW/kZsFhL/4blE78MRdP1+urv+
ak7Lbsygql4/EcynwVMGkurUMXnMDtqVGSoxcmclnVo11+k2ArIaVylX9XLMNgsh
oij3nGA7jtBtkQx6LNDNKl4yxFzGMSrdCh55W0D9w0ON3OWT8hXnD+cDj7Id3ELq
tvrq1SCsoZ+4HuPgOgGEzkyuRWebUVaxkAr774bqmtG0+TS2Oi3uz+kuMeI513Ch
2/CAYsexVY2kJ23Mig5gn+CJVHRsCIJ0RaZBIT10cfenOHlc7x4zQeKo7ItOEdbF
9cpxCAMJxDcL0Lf6QnxnQqUi7kPr745QXt4MA7NHeFbI815wMTYtjWRH1f8LrHQb
SQfWHz1Ft4UUvveIuJjOV7sYHvtvy2IBWA0sDQADXHtPU0snp/GwlXZRoIy0hwV2
pjxmkEVELkL1lRakGcWQ2f4+JklWPPR7I3dm7ml9lbQ18NsLjwI5FCUZ2TIw6cUW
wgu2Nz3vg3GBiNuJzyq4+jkVcAmUxwt72pY339JoECnp+ELZXIytKA6zkuEBrcqx
bQokVSLl4JBnB7VufzD/98yQPc/NMKcdhpF8o0NkWovXwTRxV9YjjQrbZWTLnNp3
p18gBwTj8yxEML3DLjmzBcnQeeyUAmmsvME58xh3b0fpUl+0PD0NJ4G2edA3bQM/
pDt1arp7Mc3eolPFdpxCjQFfw03JZcWa9ZmOZBQbAvBVavN7eAUzTP/0caUDk5tM
rkLr9FTBGSsmp3s8MQGTM0YC7TcVDGo8L9CQVLlS4XSx0euGIW/4GzqF5Olucwhj
j17LyyZPLeavRZKBOKAhjhZVdysbaV8nfp5qp0d+ppbngnbUuXtA8TuH2ybIm1Sf
gNLKxoQK++7j/MQrJgIwhoBd077StShebXleyLwvGGuL7PZ5ucUQqPGMC4TJ9wrP
CFsbGWnkp/kxNyKjAKPBUYsWWKWc34Ylzv9gqh9WHVIatU2Erz7zP0vO/eBeJtu1
maNXrpiLGE8eK3pUeS6b732HAgNGZTKhp/Ea1DfJ5ojvf3KWu4YUhGzlUhtADVhY
m8uHw7kVA/QnUZL4OyxXl75u87+r2O/iwqx2AA9kZCuVYS743/w3/R1GKLUV4Txe
B6n/tzMohnvrPuHtQtVzaW4HwygyVeFd2Ib1unHCNy2bK6dE4hZVf2SGhH8xTnwm
Ojq3zoiENB3fappqZ9K2bg6DxopywmpQcrVoqel5B9zSZIu/jY3B4Uyb8r6U5Gt2
Qvzm02LeDfnYX+79WYKHhKxhoVbItBv7VdOVUsHcDfvtKN6+25Aoe4wnpH7hxd1n
ET5JOEnxIKwr/ODokoYRaLOOcrwomhAn/DyfJTmEkcTp++FqpaV6h/3KUknamvAJ
EeVkvgJ2A6G7UuLYPvrk9dOY7ENjRUqueQC1QP05eXzAZx/pbAxU7ngdXGOpkq6J
Ow+l/RpXnPNGpOBhXj/U9Tbc1nWppogZ5891btbcNAcv6lcGZzUGhVpBn4/rFIGB
uJZA+D51RCqmKqBiS8BtcoMeI2ItKiHVXvoZmCxqkNsI6Z5bVPOaP4m2rNH2mAEx
SnGsEUYUOZmEJrK+31AzJUEdP3KFbLpTGcSPuUutS4b17pu8fxcZTPtcW/+Ey8us
1UBVVG9eskNT60KDhHyT7OOLi1hmWYCKYAXlAMWfGViAVdM3LMPGDdIb+C7TpdRW
0jk42id4d0v63YA8PoRtGtKvifnCpr82fvfpGd6riT2utPDeoQgIKggluc73wgKA
CAL+IEKuBghPas5WEN+WmBt8PgeieFPUYRSDyLwMKuLROqNQBP6L6km+Fol+fc+j
Km9Cm4+q3wDxiWCv+T3u8jYH1anWnFsdnw/kv4HNGbafDdVy5WvvnUs8AVIVbCFL
K4QzA9S9W/NiA79a3kM94MMrgGI2O3PWOY3hD/x9mOtNq3KWiybfXc5g/xPFBhDE
ouvJpKtlVug/lazZoA9yVAF/K18H6TvWQ4m6xEWdMHZlRf+2Yu7jZlK7KkhuGgjk
XYTZStu5FtA+1lui49/rDCxKTD1rxY5Imx2KfoVBpRfHieByOa5GIbYcj8zON6/C
r2DyVoB8nhZTKyb2oRL/WUDD7OMAqPT30LwsjE1Hw0dPKC9H+odjKKZOVboPSO8a
dQjmOeyYNtp/ONAQthnNd/afeHcqt6zKmv1zI2tKo4G5P9bOMY6SnG9LDfw8vtk4
qtRSuVW1oKkbGhbj/dPgfL15KijbyUowqiDa14xkvCiZt5TdJNA/F+l6G0iRkvmp
dUaazp/rKlhUBuj470bsGMPJrhGf0MdVdUnxtLVUYWK9v4lyRTA47B9k3/qwcZgB
BSgBZGu2XGi98qYJOWJmYTqy5yOM8woIugEYHzKCdBgQZm72Aqzwpn+m1iuDRilR
cmPuB4A6Ebc+Def0m2j+WZ5mymz84rSvBKx/tkSiDJW48rcwlmp2GIYLoE2fb9fK
rYEH8L6LacKI/cV4Vz3J3g30vf6w6/Pv19pxNC0wdRIGJRoffqnCQCTjydLQo1KM
YLjTw+lSeA8JFAxeEoioQ/kD61WKQlAgQ/1OpMkobnVri5yioM2VLNy/0SWnZlyE
FaREulGlkWiPFlYWYgOwrNOb49kzOvTH6qvCAU9VJgARN/Iefjc3v1t8vKyOLVse
mE8qEjt4XU/5wmjtU/Ph1HPV/LkInDp+j2lqc2l/lDCpqxJnpLmjhnk3mGD7OFAo
NE+mGnrcqJDZlqEIjQ8uyJMcePEe4mvPBq+EADr+SiBkmln9+lEW1jjfLE0sqooW
GUMfsHNhQxMCMxdkQu0O8LNSYgO5QpgGwj14o/lfv6WJJ5iLgORxkyWgcOkzbIaD
GLMj8syWPbF+0jhsih4BL5FT0U7cpuD4ST4DsrSiOIzxYB3LTjmBLmmvLqFwRZ6d
a2PoVXDm3jC5LLqsaNzP+3BR6lh4+wVFtl0sGbv8V3EQGv3lS2uNMbvgObSbf5za
dnF2kcG0/zTRdnbqcM/yQdiO1dtq41TXAHp3tEL46yo/f+KkUIijbsQmRaTDzOzo
+w0NvuVKLQdQzs8OICFlK6C2/q/P/l1mBbcVq4l4Hi34z8rTdl5Vh7LgL4ufk4GJ
mPSZBV5AiJdpezwDECgIBHlIDyF14+LpglRYLS3Uf4QfwtAaYX6vyMhEKfdP/VxG
XxpcDiqVNwv4hbwWTjxMZ6sWPlP9Oy/kEV9jgq9Cnv1QOZ0bof5T5ZZXjpaIx28Z
i/6BUTjWR5cJ4zFMlGU2Se0OfDvNd0CgMxeXm6CbE3xsU530/4/lbCn71SLKuouX
wDVX/UOvkXUPeHUFSFeyrS8qsuEMll5ZCtDnbx9QMcMavUK3Dz02X1e3LjwoO6NL
aAc2w5xxzq/N6R4wW0HcEcQcH4i3z1+31QLUpE7w9brZhWE6echg/IMtECyklp57
1bACURUjNwPtYLLv34fkAa6Paq1kdneA4gOx4I7OvKJsc+OWjRZrp/yGcEs6EczL
C1BC8+9FVYYKpxBJFeE1nSqKqEDzMp2cZ8+W9eC4IzwaCWw7EUXGoYuyO12r0+4Z
ZWE0X8ZITVxoTm82NXNj4vSzp5lAML6GCfk1ly7U/XniNn6uYYIBIxRhinCPe+SL
zNSpLRpGE3mItpy1YgJVD6lBcCKz6k/+2RsMI1xo//9aUFmh5CIJKcmrOVW+rJMg
YkVqVzd5URECvv4iSHY+G3KP1aBbuHWQaxl2O+QjTIrKqeIR/cfJTE5JQ39TBtPg
VZjjVWuEjKyICeYoKka98bsXhozLkRouon4AZ+cujmGt7IHTvMpzpDC3mxaZab9+
wRwWCBd4GOkWalODiElAVdeOhASz40uzMtekv37XbL++MWh6T40sAVAY6wC6SktO
ft8sIpBYTYOYM5rXkHHZ9wI3EqnuGjz0evzMnuCwC52JYqrXhAjKRk5q5E6fUb/7
hgipqT/6C+2MedZipk6cXcmOAO0E0R/7h612lAKhZkl1BZoNy4p4aNPFbJCJ/quB
2D5hPm8LuuZvm9rFiAPT/b3fD5UZNyEpy/VokNrf7kclnaOCp3PM2vBTdO2DKqYl
Fac7QJLmaeFzksBjIwTSz9pldh3dlxH0bnSdLdvEOBcABjWwiT78lVGSdUPsQTJa
H9+XLiLl+OcNdapyOLh7XjluQjB+Yy8qpOeZQuYxAUaG+2OeLTyeXUyqnfdceSmo
lMfEcXqpBWRpz9a6ij+RTzU8Wu+YgrvuYhcBkfdyn/Vv39Fy2JZT1yn3BgiaI1YL
sFoiVL0SnYDvxmSckC1Y3lkzBnjvBKJB10O+45Unw7h0abKj3sDvfLLz3mDzrRyp
xBSdZ5xgDUSH4svPFixGJCM8SKedWOqPiAcZWFI4jYuLgxRygQ3DVpSb1OqbxF/L
+C5OGYBWn3X3+VL1L8juO++LPP84AVf9gVRPeKFq4aWPpwiG/akgLYmYzJnhbZAz
M1Ak0937muoMeMJH8B5V0PR6Ey12Dwu4OWYgWg8SlruYKc1K+AQlTWbQUsDV4YCy
BVt2ughyL5qrdtCZE1d2FKLaJwdXj4E1Vzx1x/XOUjfFYOY7cOYaGwHu+rE8sTkx
rlaKqXPjKN+dwqTZBYkmh86SdvNoj6mKnUtuvHRvlW7xilaz/4ydIG7T9/xP/XbN
5OWAzm8F/vyHxJ5q6pyiAiInaIU/RMYbN7QLrkPo0HrMhzS0uEn7dg0JcghVQXQf
f1N61MPfk4oCSdKZoXO62qLDZk0d/KJNnq5HErw4N3EEQvu/XD++Qo863T1/SICU
PvgbisXNACPsi9vLg1m8gKRJMrMab0YUhbNihk+YmTABMhxxQdXcQbkINZ4Aco5M
e+9NXyLfHhIZSjxu9sJ+XIduDeXEofy9pGTLXcZ8XbavmLzMFDZ1zksRDj4AlCLa
AYepAcPkmZVS0SLkzrcYex/+ktxwesqp1Xooqw/gAoMxRSlhY8TXMiX6Y1rA+/kA
VxPxP9W3HWPGUpzPiYPRvg4AvNgEs1zSaqvFNZCmsWrp+ri4YAn2KE4xAwTnVZFe
BFQXWvmEomtZZ10GSjx19tx76MOsxE7E4AACN8477JnN2lIgK+s+zygo4mLTIF2k
fXopks6vexTuTCafJS/GQ/JnfqzEBhXMHny5HB/i7tY3nAlNK/YmpO4G1QYH+a/j
ARnFSN2ZUK+WJO4MWn0d88M+E8uv8/5uPpi+n5j/cIlWhv3aUsuvN3KMsp886qlE
a/9OlnkvqZCfkFAODOQqMva8z03O+UQ6VmN8tpJhZbrmmwMrY6lB197Hr7Ws3Vim
wpfBa8/YuXr4IWQHyx0la6vez4zTe4PrsFr+ToLGTSQuv6v+pxEb6JDkHYWePKNu
upd6WG7ah65KAmukzwhwYW7CNZBwdOF3IwETkeQSEGr3yMNinslj8DjrUu3JRCOw
m1xoW7qPq69htk2fAxHzadeSnDoSqlkMOcSKgAAKr9Mei4uNAJkYzK6PPbj/H/j6
T82S5npfMnPbrI0UDVOvz+4FVvQ1hPGvC+f4K8HwUB6QzS31XsjeQBdDg3XUl/y+
v4BpVZIPko1OceYnbH6eiMDNSw9/5Jjh8V7NyYSD85zXr4U4vgYTj/zxtt3cbflz
Uf7WZOC2TFrtGoyrYoPEB6WftCmWAD59q7wa4fI6cDuuXt72vffbm0JBS2MJG1vs
3tjQdZ4R1AAXWFcRT8DsN0bQNnuOmnyrrJCgnXbfIo2TqpvaLCCFMceoPi/KrcBb
G2tckBMIrpXXjh9Mw9pQCln/IIBJYtbiRwKFUM9WfVAK/7MiJmy2vnkusYc9orfu
rrf5eCbtjylbs4Ysq19DB4m9hlarKy6PeATj7QJtyfd+Nha8JlyIISPVdsaGYuU5
xJyXFg+6/LjNaBnJbuZV2B5Vn85ZVUSisCCxY+uuy37Y2CLSz5UZNnbiwyEHJNI4
k38B+mUhwQCLAvGS15YMaiRZ57x2DyjneU5TvPraKAijL38ARxN2PY1qq454BuAJ
QJw/MN7+JrQHZXGy45HOOOXiUsHgugpRKjvjOFWCt9MqEzCLbChqO6Zng5iqFxER
lsH0PtvtRCMMr9tTygBmu6WxhW2UtXD67YSsRnNXx5IZM7qD0WKsdVhEkPAc1u9u
k7k40+pEZR658pAltCfzAFpvaQT0thdQiE8Gpvc8jrUi0dvm3Q+etjo2mGc0z3M6
EQtui2LgN5m1jSkgTETUvAUhcoXiclzxQoF+SMkRVM/zZqnoGHDiMGaqIIc41K5p
82LTmbomTmQ6dVO/8itWJie3s8qQsHtK+3wx439DjMNvBVfvEE68WK3Kbp458/fQ
pPhIqH7akOaebl+oskRzZFvI1QQp+AzrK8SpTQcD1Nlry0K7QTXoZwpEoIzPE50N
p0Xjc1huUbICTB1vv73ZzAPVAHrtWguKFQKIX/dW/t/dtlV/kz5X39KiBTrar6nh
uCDuNgZvLeYmvRgUhbjA15OTfnIgpFuRw3wpNPjlHJ6eQdZvUh8JlDHVzXEDD3aT
U96hcdzTkJOUEyAM6BK1UuLsn0L2tQROEIC98eTCKJEu3uD1n7Or8VfPfztbg6md
tM+NkO0B1vcc2tnovVxotfINpzw5koaGY5zf35sgAG6y6SpP5SJPlg4vLyPS1egZ
Wxs1xLyvtxIIOhQGPUNeodSFULcTMosMwQARF/WGGssHp9aKQMTkpEU1XSCkmf45
/IDqRi2M00Mp9O/a8s4I/HRBeOsp/TtL5fNCxh4VTE2dk9PuuR2OplufpJGsoerW
ZBDeTTQY9h0eHdek8W5dYNXHygQbSursom/41WNOupRuzk/xkWDexM/gBoXmWAVO
TpIh+JJD363ltsKsSknaMdP4vrWsn/+3CJPV4NZtZVwa3ACTnOFCdx3kDyF+LM60
Jlmesm+qLLxizZFRai8NSkqigXbVyiJB6Z/KTZZ1pacgjWzJbSMEmhCmt0HmBIfn
ex8zqT/ERP4TosyUJsa6R1EP7fc9kyLvzefSs/kgfPcLm5/mUqXgYOy+43WjlKuS
YC0WSgFrMv5SkMLHrF2QQzQyW3gcUUmTnhJZr124uncn+W5h43gSaOfh+vLD0IAi
AuVU+Xbdpu4nPCtl3DEC+VfRW+YguMyD6nprkMb7GG0rjnqtu3guMcWe/JAcupUS
YF2w1T7fJVPIXpkcIBEuo6xO4A6LH1aUP9p0k49RGW2/Q+OI+0Y4cKgMGkIS8BfP
JB06L54NJxVXcnfAg9IDTysL7RWXyqxWq4lhEzVy5BlMbjhruMj9fPyOidaL54K7
MgEkoQXEB+cQMNTPnu5wks72y5Jqk2qpghVYumwcLxO0hY5f678oJT0hHNZ9SEUh
TmvfwjiQs6Dqh9Flig7Z3DHy3JS+sCOPTLwcTYlASkoyo/hSCmqAjYGvV9N4vaSB
crUvL/q2awNS9rm3QhbkSvNNWFDhCN3p1hLDrzTm04x+a5eycmqXzrzjVAxB2UoE
KOGcWR/6CEhlT8e+n7+E8/Y6mJwz8hSYlZviI5R1gQu2+syDwZzTXNDm51OVhsdK
hyGvElsbZZaTlhXHeH4rhVR8GgVU2PFuUJ/35j2dXzxFcz1wUK1f4FJpRc3TOOoy
jMaLb5+xnVJvTdtPyyiLNcGiQ29tE4NEFfvX1oP6g1DnYVQyMAwQZ7r0MBeKbKRK
kgGnYiDUcJc0kqw5t58wyiz49+JpWPVrHPx+TWOEZtvpA7q8EXP1+D7wWjR1gFzY
ts4vlpFyQToLONuuklVLie3YkmwV5dZDUo3mFRLukHI/duLhNVlv1FyzHrT/ltgt
QAaR/lkLGEx4LG8105TW6hdnzdlIBYBiJz/rsksG5glbnDOke6sEuYz9e1O9uSDP
bpkfd9+/U/9/dyWSfljgSyBvQYSaRH57YfTYJOHvn0aqJO+jd6ftUE5YufD6Ut3M
g/ID3nKBgmtrJERpsRnJMyAVZvq8zXOjsQKcegnEs0JvFa1aSoRx3h4xpVfYqghK
XXgJDZH6LRLdDP+g0SP6ZWAeUKTe1nyzwzNGIp8oVgNVg8zu6x+BtVVCw4ex2s8B
sv9UFD33EbojxmwACUddNIgukfyNuzk7Btte4XtmZRz/Y5IzDT3t4+qdu4VbYeZv
LPViqvtvNJG6UIs+jx7PX/37FC05S55moABcLtISAkyZuZaeZmCWtwbkSgfAHGRs
VrvyAtAUtpO0XVr9pHO70ICdPdVSYbdVcAMfiQq2NfJErLeE4P7dtJBcg4ro+4vo
M5FY6wpbo2vMKnEk/sVQHRqe8os2eo2CrSuBXQb2fHuEP6jhbWAbZhWg44xZtLMr
+LlTyyj3qAN6U+19afiSeOxnpfvvgzaqEpUNhoR59j13ksYMjhwi+X75BC7zjU28
qJZunWhTkPbax8oZVvezzktiAyK11o4z+ilUvCVjBfjLm6uMEW3xlp4S0tOOkXnt
k0o4jZW5OaYJAD+lSucEnuiMX2n6iBaZjQ00niqK4gCngZpUj50FhEf7hfK/qdTF
T9+lRe5EY+vEnzSZXuADzDKv58FsLhBdr1V10UgxXVXxHwM10YGz4V7/xxt8+P7f
AeOhQ1/aMA0lrrsT0XSrHZECQRKT3O/qBoNJLXXE12b1D/qv+FiMQEUKGZ+qrTeC
05ZmEQcrZPKxcZzU8dayaCVpeu9e+5oGaPk5sowisO2hEvwfRWAiBlZVXG2PpwRT
Jd06IVZcuInOdGTRwXdYY4+f/iyJ8XfJ8yawwqpARofF2Im4IfqYEr2212VtREC7
i8l2R3A4RCi7ualU7rSfNIS6tytR/BHLRATEfCqhzk2hPeWsbJ4fx2QsibdjenJw
ig/l4y0Qu9kwk62HVAZ0pt+HlfetvfDK61vezIOsrK7F+P5XCIyysa1UIr6cz/yk
bwtGJBK+ovnzGZQJXlqw1K3+GmhBvm6WSqhzceqMLslEkzd5D6MLOQLMOBAaTcos
f/u4YQ54ae+CFO7X0evqrRXEUDzH0a9C8O7it60RARv6moMvgMlIBxEhQXQ4rnd6
aPnUSH+NMmZ7Mt9+69D6hNPbLGJDTsbprm1CMGDhV7lUZ5O/k8GIiV00O0Yz/tkJ
OqCKxmov24oEYjCKYSVrmLMcmMJnRac5pxL+bQ3aUyvAkUXWn2hImNl8TYFaldov
hp4W0zVkLVuBw2O6nip+w7h76KanaVqpQ1EhezfF3DNiyWPWD78eDcQL/0FDz+08
BNxG/6zcNMo1AKz8FRIZlWpCvMg0HPs4gH8dgg7Hu3LG101PEae2GfxbGp3EMkeb
Sr2G1Ftrqzs+epvDVhbOxpZr02QuWhVPTILNv+P9OAd03xJ3BKloQhxgbvbPbJ88
EmtL1FDReA7qOD0kQ77WDSuyb6cC5SRsqU7vcfbI3iOn9CWKMzqzQXBoOdXPX8Qz
s2JfTJtzyejdz1ex3gXhNGl4LZ8C9Z/PzQY+Gb3tO/s0/mHwCa0TEMLmN8fJ+Oyr
g0bK1rUlm5B+5qawfb/R5aSLq8yl2js0kESSMt/sh6DJm3heB5Sf9GEGOPMCtRCU
2FQLRPxv97hNX8cqX9pi3LnK/BYUu80M2oiVPpHN+QBInGNmSpyUHQ5GtKbl5Dm3
F5vdKtuvROmtrf5c1ljUhAUd3wQN6fpPphbDdCLVxwIwbLRQB34s1fpWyO+9wr4r
LBjWpVtitCrmZ1u64ChT8LJ4YSHrD8MmwPK7pkbGP2iAu7KQgsp1VW6JjTcMoD7G
T+nkLpjDktxUfNOE9s7crM8r5xZdyYsbTo3AE/hARNgV4S19NVKTQA630E5JXci7
Y4tJ5Ex5xuJ1IFzvllQWLY6aPlfsYmVt0VcUJMFoz6UFZwrtz5m7XLL2gAjeOcbd
KEfIq4FkvR8xLVb25l5v3hGbjByJZhHlue7Hv/MXm5Y4Vhqp0v1qNP955hh1fdUm
ssS4H4Js1Mwl0a+WOIEGerBny5sZeoH9hmRlPnl6nH3O+rtYRlAE3qxcahhFJQW3
ecIIkbOxEEwQo2BQ0bXygHC9S8alZ89075YGPNDmQXHUMDuVbVOBqG9T8H8CK0FY
VGWl56IT+qMQTxgDshOg9yHt3FVuNkbW5ggc0qN4Gln33yVOcxrXVvKfaXTs8AC+
R0BW8hh0wRp3EksS1Z1iNmBB3jVUCZwn2V7dKqTKLLQiP841tHMsM29rZgxRdr8c
hIT8sDZmgDvBxyR82SZPhkM2LH87MYnqoov955jexcuPa6eBar1bxoE21OG2Bflf
wu6WtN1BWV1dC4Am82L6c3RyQEfCril8tohH5V+tbB8lS2bdMzGyQn6bhpvFHwip
jsWGtRPJ0htj9/+i0nzExlINtn3tMSkwjadYjldXPle92CdpUmV7/ILBpPc9Sd0L
7tLWO9GYsUzs/iJBgygSjv4CGebYbuh3mpelRSwgYs8KBBnKlUWzCqp1VJgIYdp7
JUWxxAZHtNBWiqazVT7q0Uul61o9hZXkQy93f7nf1U+6ODjWuDc2IylXQY1aKNJs
wYBuUCtjzXc4apJjNXMZnnE1Odk9P5puCem/gOo9sNpA6teEbe+RiDRJcmMk/RyE
Lnal7cGX/3732gI8ClBNgicIcZUJIiWmmougrcbgK3Zr0TP4gwoqgAN/XnrkdaTR
YtzuqtkdPBVPDa3q4aBqFRm+YoKRAj3sF6aLrI7um/QjCUWhtcGvxE2n706p5hwF
oijsvlU6G7aP9JacC7JBm6RbNTTe5BhwBz3++QyqKIxYWOda47CUyXmAVzDMUZSj
AW9awpjwkHRbGAvOIk9NXYiiYnIGexNLukSVM+3IzWjhduNGrjdDcaKfUqI7/90N
iAubmujdGZvwK3sKXhl+9+Xbdv7L5TX7kBIgFNkqmYIKSmR46G0AGL+t5IRLCQFK
ogQcyL53Qz8zBVH9/bTN4WsIDFBzZSACys8Rx0x844qCvUYf+IKUa/o6KYA1m8ZL
bZAgfSSGMboKgzuygSitndYC5TSttr9z6dNkJzrZmmg0ax9Ay0gBxYCuzJoKqdt/
l8ymvNKrj7wK+MzW7wFwKPcT80wFaUTihCxvhePdwSBpdqpue92qXETDXjy4Ei6H
WOoNMHCSAzXUmjPZVS9Ju5qrUYcTg1vYzuu6Y7wiXh4mnQZm/HuSiWXnXkv31AFg
44qZgR11YJ/3L5QdIfWb2JGQkIAyYD3kFMdu6bFvyb56sYz/WJqmvja7AQK9jDoo
gn83qSqhF/FxbmouCU4RK7cxxGj3cbiN6Yt3jzs3JFqmHe9ZKNXQbSujqOWWxblW
+WyQiValUc++IJi0d8nXkpcxXUNB7Of77+jL2hYXKUnUFf2LEQPWxD6MgnOYO66S
EC9+24yoj5XjiKNDASQJ8NRth2foWFEHVeMPxv6yv60QwQXzDcdMH3N8O+Lt/1cC
yMh3wqYfdHo5j67bArdO4Ri+dgmpFWyCVMCPsqrFjJ/nyVQMVa+L1e6O5L/c1u6H
wxnEivCeYEmHQBfr0BL6+vdiLY8YoQ01tbVGDh+2pIANyNGp4ZyPeCQq60Q0eF3g
Ik4J4HJ6pc5V/sl9R54E+y3D70OZPsfhO+VKon20R6OGtoaAq+QVAdes3/woAC14
gKNftA1dSmyfRDKg41szp9KQ1nCK3gKtgTw9jZZlJX8bQ5JD8EL2yvYjbfpHFONE
vc78Ru6TEcwmOdEq3bBidMaBeqyv38eL34Aa1+z9LT//EW9sGU1D0isqfHktZy0R
5kRv+hdrfU1yySGXaR1AUu0xx8EvBIMQrn0Y3KIZBZxQlUFBLvJZrP6GwaRqGCMq
j7XYIYZXa0BKtfZSe0kKvfjgE669/tznsMmm4yVk6voEEOsjAwTY0To7IBjqc88+
Xqm+VfZUp5byvxel5mFNEjQ1EMAqqeoPWgwxeGvvOtpHtYVduRcyxOec/FJfGGt9
85Y5aJdq999k6kjmuKOThU/PFTlmfVz7p30V2NpQWe432NUasRt+Zum3NIppyiL1
CWSWc5o/2BJT8OV4mvU0yKFgnA1ZkSDs8ClMYD9YXt/7j+VwM39jl6JhcFX9opFp
t+ZYUiq4nUfzVEM8jFbk0h61HqVAi54HFu8u6aRaUfsBhCQPWFT2pXT6mmoQXla4
8b4MiGpyviev5+0z4V7U+nbKif15JYDBOXuZf/PC/pjq/kX1o5jbSpNAzC7sBZH3
qwBvSnzU5lSuaAcKmks4AbhslSvqJjVtnnoVuGOBxzlKapPNCXK/5SY5lTUprMmC
HSDRHy0YkBnadKesQyQ8qLYoJIApG/FWJbCPZWd8//O6lL8Lyajui4j8xJDM5PKe
GB/XunGrknKlDfRn1/H8BNjRiJN2YCOx/dyCDCzZfZPYcwbtRU4THdnDo08kApfZ
kUlZ89aN022NS9XZESY/8Pv5+/4QkTLIwjpg+PBF+IxYvoz8nltknRyfuTkyRqXA
Umm+UmTUmQBoI4EGk2+PBiftiURQNB5+xuj1wZqKVO5WznjxGe2LYej0KgsUb54i
eRhKnGM4oTl8KrteRE85mvAJpqIa6P1kirwE5e4KiBhbdW+LrwgJO+rzs872FMdc
flfGnTFUIazqDszh5wijIGF0lDYy7lJD9bqeESBAyYUBAUdO+/pa6WVAJb0NIYoG
kMsEUSKSCxMh0vW+2SASiX/2Ty3AxXZTzbXDT5KWnOEF7HJO+IH7Y8uaD9VZ62cN
ACrdd8+q1OqvzzoowGTuxR2ewGtzPjoMjQ0+JkStdgZHD3anXfeZpVZeTcQ0dtNh
LMBLkA+sa0IP9xWcTInr38G7Q4G1n4BAwBD2uOz+0BmTF6fEDAn73nOtj3ROezBY
rvkEG/XsO1+uQKXy2YvUb2PEdWzrsqKikxI2FAa+QnHOVceZ1ChpCZXDMM6v9aHr
a/mtAvygBcGp9k5YBQahkkuwmra5w4z+BIlWR8Wz0sd9aMLHPjd7S/BniO/4MVKk
rOZIUCiSs0vGzS2vgZeoYcDF5cPDKrzoprNGiUOvi8CnRKYkDlm1U+CSDRLZy+KN
FDUdAceKfGI8j6jA/Xju0WuiukMAz2ArvTtcDTT/hZQtxpSwtuIUvccLIQSuVmRQ
5O/EF9E0cTXy5H/brG3T5vgbqcNpfO5M8YMl7T2Cjf6s4/1Ty96u7PwY4CayeFmE
SBHMlaoeQGC8Lv1j4vms5QDMF/MQf7bfoxOQa6MNVPD8qm63OKJNzLjaKyMArO4o
8/hXSUKjqs57cpzdGg+8cM1mfNyLHpTtHbOxqiAdnazCJqgX0frUhP2SzcvCMi0H
4xPL7x6DJSR92Lm+/Ka9bgsPIi6VprtUnf2DLkZaiJtr4L6Kw7BXBmcjNNMG7nzT
cZohQwlOgZmh+q3IPq0PuZKrko8t8Lj4vvv8lDA+PqAVhtQ+fcgF6PB3udAKg0jP
ZajmCSyRqMbU6WFTWBPrAKXVOwMNdFvgLqb2o4BWSuohkXpQLEh2LxKO/CH4SpG0
Gs9O6mdh6c00HvMKWVd17lwu7l/Z/pqy+qllGkly1ksVG7agexGD0V4C5KXrjdCE
nvXV47yPiYCGPa1K/FMN1DGb7ccA9v2JcR1emzOTI7bDikLAcX1hTebIlQJa2EQM
5DehawI2+2h51TAJ5Qfg3PlHerh6IiX0H4Y02ZatX1opG22uCtnaUH02LO9xr6f4
Om4wAkkxpD+ap7oEM2LdA4qZjsYXga4WKr6X4JOOqcS+4MqF0OlkYLJv93IFVaLW
Eg5TlFZwYv0KeJpZrxhHU5qZg/FGynVNmiNYsGZYHVVQKnsmtKaIkx+5FUcil2YN
KWeO0ZZOJ1gd21bnhyoSNBiHy2mbAx3dap/XnzSUrSh2eUudS+GYv5IPCzexbY1W
J/Xx7sHYnhQWrrcYE21w6FEyCrpPsi9iFDdkhhBus4GTfBscPUM6QZOV44+f/EVr
buhYzPP5WYMCWG3oUt7ZsZcuQT/untSDGQAJCNMi+dOhOPO/zPZRDyybWIM0HHQB
GgYNwV0+U6cgZwXcJqFVCh2Nfc0/5XQ/wBF301O2PQfdNjMRGin9e2rc1XMvcqtR
KfYeMMNF3Idn8aBjeU8mlQVkMci9Iui9idfyPsMiJEE+Fkg1tlJUp3bkHCfpoxjF
45T1ztOE7ABsgpcFmSwOKYI27dmqTvWteGPj9AQajg7Ffik1IPfSnXFk9Iz9dprL
x7eboJXEkgmeFQkOd7aNjoy5juQQtKDaoZvSVkWr/pTmYCUxosGJCD9rIbucX9fV
lMA5gKMLIEOmeEZhKGrBB32Jhh2OPo42PbWIR0bMMDn/d/ZtAWNScReDuZTtxndy
Olmnr8shJNnDalFhh7SJQ6tqiujOQaiuN5NPGyi4o/GE2SevvmX/qMFmjzkTdZRH
RQtM6m4X3ghKiCPWtHIH/OgEgmHJJz7LGjWk1IjozOe2yF6J8iqFWBPF2OwgoAjj
glhBPubgw5iImOK8G8CphNtVPjX8j8hsf9JN3f6+8YZOz3RDSx3D1tAanGHZ0/Y7
gbRs381ge4SG9qZX/lYDdQVii/4lOtZ+dgSa9DjxZH52TBvIVqX8CunMFx823W/5
EuIhBlrPNCalYeAUXXEEEffpGHQg85bZOW9hfEjhznNGxLuNTwIYtvSsnkiU9+Rw
HPdYdx7GyQaCIlqoM7DqbE7zbHI16P02g/m8zQhN9AsLmlPTPdD6PrSF6fLRLrNf
JInH6bdzOM9mouQmQUFWmlGaINS7HclnBFw/xRXLZj67/05FB3qKVxHEWFxaSTd1
E5x67S1UxjPMe/6QfAZMzC4tJCphvWTbtr96doWYODGF0/QLz+pSUxd2A+DBTHsQ
+AcoDFz2XuGap3qTTvk94egnAZM3nhdLm144G0K2cR/o0h+F4fW1tpJu3A/7To/p
JDoE4wa2IEitvB97odUCNecQZiKAnK9zUjo/NYt2SFAuiXlO+bhOm4aSMYk4j3g8
6pbmNzcIuQUeOQHjocYFWuPb/pS2Oi5oE9/j79NpRxQ/oVVAURgFFNsyytVYyBXz
/lXlDCO8hzOORwpMtRlwcnP28lMW2xlTwgpmACits/I4AMLeOYCjap1WfEAHOi0K
jgMV7zej5x3EwqO+0qhWGfYRzO3kT+MgfdNS+qr3lG+FZBJHS0E/9iAUG+IdTgXf
XPUJ9OdCox7OxaEUyvQNkidocG6allxk3+BsxnnvsyXe5fOgEvl+vwM88/udevMF
wzWO6i2yDcWV9WGxbiCyM7c6zCs2hKnKLrBCIlBv2Md9HpwGCLLdymek2tQ5u3E0
Gy+UX4qbI8W5Q/dq/iNQ9Dx0pHybBInZHkTmbQkogJ0fSWltngtFQoe9g1N4dBqr
v/B5ugJmXVQNiYwIMc5bXkQNZD+e72Cs+L4WkBdIVLyrAPkJh0z2vy2jh7N20duN
oKPQIbG00RjnP1Y9UqoT/6G1AGJJ/F37z6OZ6MqXVaqtFmJEwu0JtKcJ2lRLDJU/
wewBQf7UeiFc3SRgToL6z+JFyKmK7C8MFtChWBe2niMrzn+ENLGX6H5OowreyUrQ
gyuuYmCraFvwXOK8AXjcNtxTQj5rYhKnOdsPOB7ivgM5r/Oagyd+rWExkgIzzHZC
H2GRJcaZRStP0Hc7BEpoHne8mTZ97uhFfiKg/T4OGCo633MkuIW48iJ+5KZ7/LdZ
E2ZGG/G/A2FulxXeTvjFTFcLpKSlpMfj5dpOz0qumo3fS0m8BEElU9sgf6dGdIeD
KHL/Wbze6YIpH3xdkl2zjEJ/83GEO5Uzn7NpvajnXuDta38wqgHsQ+UoC811nZcv
dRKALq/Xq7DZuFJaUeHgWIP4BpGC2eZ/VwePOMiJH+J9QNpc6lIfqLQ8ZryfR+Z7
HBtJZlMBr951Y9PVhrnVln3joWlYH5ZfK4FZONzqQwsct3pTkz0BY/I94I8UYaFS
YnWrM4HhrKFN1tIv6qdvWxd47ad9KRhu/OdQVPK6XNnYKTPjYFLX5QyBRAP7qv98
7Z8mWcAvITTIp7E5SJL2SdqsgMo6CXVI9SxCH2oJLf2/Be7ncJxYKYvHRW06fm3e
a+afHzodW1R+MoPnM1nDdVsUvihQqFIf/S61GWcXXW6Vubesx18a+8I6bogWvXm3
3JOnFcem1lxGyExBlJIxOwh/sdnt7HlVATN5/wq1nCaJyXeP84yAbyKIo4spvYd6
YmQMuUGdOFvZW/T+olfC4XF/Va/mizq5zDpYvNI4ylric5/KOifLI48u/52qZSWd
BuJwKHWBSfrJGx0fDmC0o1H0q4as0nxz1NKtHjWk1NDpft2uVWmHjAzP9QjcSUA9
Rf2zEz47S+klCFPcBeQ5EB2FvDL4mI/G8idchbwUevCT9GTLYF6Yi7zamtQNMNwz
Rv0oSf9c04cvxP3oNJlTUvlGxBziDRFFHVx5KytFKmi61ehbUk9aEGMAsilnFuz2
S7p/ZAaOBan2uBwr7tdvVNSb5dIrBsuc7w8qtMOg397P3mAXWKINqO7OxqMj9ldv
9cw+gdAbs+de9hwCnOByS+dz0L4fpfVwsmNDq4zGJlpJyIak8fdj/JwZQW5a8NWx
YBGh2RdzUx+e4GCgWAgzDAObuMNu1Fm/bI/7pQxvtzcB837q3mbeFDqYogSiCZ9w
FFcT0x7ANQpMvDAtD9vwrdeHLPBnyLb99ebm1HcRjqKD7tlU8vu0RLR9o9iorEN2
HPfAxsZth/fQYSQSrW2veDOr/hytaoeKjBYCGUSqLBXRXbrl3zssLebBcoxxC0Ju
B59jmGUanIfDlzGQRskfrtJFQJFWtp188cAyj5YIg3+t2kbZ8YNRkC18dvNqYDJf
Huzv4bqLZ7KwOH06Im95ZDJoh51rcb/K0NGotDS/LOAixUmWHtB0vdlFG0KnY7VL
ANBUscfOEtWQmOd3xxYgcr3k9zLGBDozu6IoRN+c2gTMdPIUzrHL0yH1p9/gInWR
vSUETYdmDLAyPlh+pUc4JsgKxSh4QVcqXbtFGb3tdvJyUNTYmeqK1SRueMqHI/Gc
w26XVZ/A1qlz/lhzw/1ubFqiaTxwWsWWD74GrCOjv+rVV3gHksJblrD9O3bT0ksr
bVvVRAMTlND3hf07q/WY6Yp01mVU9pJPat3GliyNHjZd6RYgZuzL8nOBdaJfS9ek
Yj57l0jzVJSectUVOCRSpykBhtDyUFrI25ZYdPjinPLwPg9nXgJNfCzlm1v86DGQ
mP3h+bRn+37Vc07a2L/xsRNOPr1v3PU/vTsExmobKJnZ7juhcL7XX24Onq7KHP5H
FFamwq9UY3f6ZiIjgWG+BRRJ0ITLBpI3wnOz173ekuduleCZL8SPrC9Krh3br7g/
Q9rJnYA5cdAgVz3WvmzySxnVYbaqP00mqboRMQJ4NnSx7qDfHRKgYx5YRNveAfg2
Tgz3i59CMglmWHAJZ8CJABDllWxX8i1RR6rUAQR9BO9eLdIcD8umwBrQ+DktDly2
suPMQZFHQtCKQ6yckhKG4ZjwN+S0wyRKZ1FI3Fck/4wQDUnT3OqBExTSDGD6Ctp0
faTdxPUKE05qm15zkEtgY7tJJxX6AK/BVLmOYs/fk1EDlXBvbLqecEbE5LMwOGqK
n2ncKi6kDCCY9/OKpHVbl4DGoynRsGorOOz678axyM5MkNUtOg6PBUBuQlrCIW5O
Dgemi5/g8Qk8b5cNog1O9phl16Q7PQq3OCzrdSRvOPt8/IxJ4S/CHrSVKXhJQ0jN
TQts6GisFE+2Py69Te8HzwuDPCy061swgpB2qYs0b2YI1e5Fny0/3uNySEBCL5N9
sYCVEeye7178QU9BaNxDuscPBaWDnpFC9MEj6NlzfEKbIvsYq1euOxY1pF2gCuZh
fIjZVlusM9cmPhLEYx9mkPXX15wNBwcnaAth+DnvpNru5MUK9sFxXfWspxbvv4U2
zZUhq4E/ZNiUWOcCaklaNoZqo8R2yi7wVYtlAjdLJAWlNUvX3s5WZ2D0hzRK3HPa
m9XEu9+U3sGPlj3qBGN/hqQZENnnP+qWIlg6jnMguwO1YsKmG5MxV1OyBb4nUeGR
VtNMlmhCRkFh5oJwNCnv37jWUKI8LsAAK20Gjrh04OReIjCo9IjsjDkz4usNIVk9
Sg6rbZIh5zL3CEuv/4GoTY6I1r0VZVDoA7Lwbf85k6b2JXqvBW0hZcjFS5WBH2Pp
JoUDccwisFvp1yop1zglU9G25kcEFkwa2gumQZMzVUn/BD2wJL3I0NpQppfAK17+
5N2NJ4MH1Q8sPCWe6q3JgtCu+eiHYl+ABG13jIoa5SG8wosRunI8Gd6TevgZ2eLn
i5QD1MynW2KEeLT86B1Xakt92GYlQLB8ijJeSR1DHgXGO9HXSlqKi1kgzX3+TgV4
S1JZalCgJLbsiZJOAKiyoNxWzB1426Qb6itwifRmp6gnim/Uup+9+X3QRy2zZvuS
OShYKOG+mhIkn55GCblolRedFu4WT3xjEcKkm5mqS29Hg8FS+GZl8Pnmvff+E1GC
T04E0gfg6m176dGxGh1HreqFBQTv2qasgTsYwwYcmSud/uueIRb4eAR2x3h3rMF9
/mtbMjWmyNcIEOvJYN/PCsLrPU5DGDHqIBohnBCJJzPq+aBIXbhd6wnTCGo1h6kD
KmSqSXq3wIJvhKWF2bLznSeag1PzgokYftG72xHahnDXz06eNeU2OStDrIvjuH8x
B73krUEkItPplH62p04PNyYN1EdHZU1MK/Fx+DVut28XMKhT+OEkbmGOA1zGBPIN
ukwB6MEcpTMnSxiotLLa9WHvRy2qxKVtw0+59PDWVxdSb3qPTqC5B/mb7+LuYmdV
yRiUKninvj1YppLZZ3eTklSzHmn66SldhKT4cKjRGqyigwt1XEp1IzzIuK4MMOf4
yc7YimpLuGAjaPe4zIU4FvhfmT/OEELcEdbm6SK6WRDIG1ilHdBpoSszGVPKIPCb
Q35C/dnWK/uPDnLU6cfgNVCwlKUyRzi7BbKhr6uLY5wHMhcovDRQgc7XR99zvnWW
fl/WW3L8l9pBrCbumriIS+aYV5c0CxVyNDm7MjNiYpFidh10Sm15eK7JamY6yMkv
BXn7NKMyEA4T3lAlz2XpldSmf9iqTOuI6DpdAUPFyso8xV/Ki9nmL/hcWilDHT8h
R1BnsYPAsLqMYXosI8+S6Z+Pg68UcI7kDouGlituToXjURAe6cXjJ/VfJN79IeNM
aTH24dpoWdklTs/KdSiXH/XurS7NP1xN84pFLu+G6p6Ghe2RFmy+0+bcabPNcsHI
3wcfC/d/3YPzbLptbt7axmvFIrEkMlPEafQ1r4EeDKjRda3Dd/BfoCXvHW9JgfcL
vmd/wMu7iwaitMeKFbBV93pwkE0iWpl2vuUopVfrj5urZwgg088mOVWZy7SkyffB
Hx4E+DF1+sk0TsDqBpKqs6opKqqqpcaNZodJ2KhwqdC9uT0r0Ctc/x/6BYKUTYzP
uJftX+WD6VwGeSfkVmi9nTJMnOngou/WFGMp1lyGJngshRo82nWQZmV0H1li4yok
mFYch7U2pkmd7di+u9+OcqnJUUmESQ3Dz/6ROHw9FI5SRnBsoCFZQCJ2JXFulUVn
/WIViVS8paYhOtL9naDzMyV8Tp7ssnPYqHPd3v7LNhmDRCuSFheFVkwhyNAs56sp
XNx3pFKwYtUSrGEd2puSWtNryZBnzcbpwECOyIsfF/3R5OIupKy1cks1wB7D1114
+rBKo+U7agMxnW2JE/S5wCVeUYjAT255VNPExLa1kpIfkaGdOMvDIOSn1qQD+SaH
mDAsW2sbWNJDkY3Cqqq1SBVM+o6wDGvphaMdQvf98ia0M8x27RYiU3I+LiCurkcj
xTUbo7e1llAkGkkHC2NbBa6dNkQSW5/j5oqegOiFSxJnBlrt00vkqmBP/0usKFgw
7KMYV8dC1gxlhrnH7+vDaCnrnBApXPNYdeQ3sgMOuHUZ9C+tOdz++31Q+67Q2WS/
kpjOo6nYO8zFChFkyxjg5JAyotuDKlJ/wQuKO9lTweh6FIl7JyBQRVr8fnu7nYrx
xG6Ncuep03OiKR3KUHQICoKoFqbKAElC8v5vS1Ro8lzJFs6/SXPQWS4sWpFdNTto
waprLSPX9guUJQ6lpON0gJGiK5fJmPwqlYLLEmj8xU5idokWeEG1ZUFG6i7JiQDt
o/GmEBJoSEgYJNUsrhbX+LHpWFOQb58rt7txIQe+6yoE68vk4gctIkAE5CrEZp/y
rAWqG6SU1kzXiS3pIX+gvkKq3rOABhPnAZ5cNTxklGc50gv+COq9F/8QZbbvkvb9
3bzUxOhCZSXxVAd2h45aZVRvWqFlmkTjuvu7LfRn6/oN7+QM1OILZLwtZRP9tLsy
CJpDJyVw8lo6HY4cH1EIO5Tkyba1mVpRzHJ3gTcw2vXu2za+l/7H4y7cK6ff7jHE
/9lQvUzcMHonbHBqKssaMAnQG54GA2FLUCvpqVCfw7q3WINJdliUI6KGPa0nYB9s
0Ozcvotzk1fIXOO0EOq+nBPgmc8psbjw/4dIgGMRKyD0EGiu4MTy0yPfO7s/QxO5
ZVYgFA2OHc7v6phJnlbppbRPg2cRLu5ZPSVeR1sFq350OFnJD1tSAQru/Hh5VmKl
+RbvdIARwHVpEg6ucDdziHac/FpFKeUx9T7WS2wNLFSe+rT78jJGv/iBtUJWijnr
EMdKVUiLnR1oWOvP0zWXWZLnj7bXYoWn9xfz5owGpHVjaitymib1vDGSG3zPcYl8
M6sQg0a3UDY/YZKbQp1kY/OOZmnPar+3jRYPDqp3Q7illGqNpY5uOxOtgzNRuRbN
l1jyXHQBGvxjpxCwENFC46W6lkeYpt7TBlyokWBGqeD4pznjXGvarWlgH40SBzA+
EOsp6FZK3WjMJbYH7+4O6tw/PCgkMA1E7ELRblkeTV4tGHdbP0Ys3w8GC/xrbdj8
vpiIBw/GVT6dv8v2Nnff4x2V5ldQZMwqB53NG3U8gmv04RFyi1ExVjeD3OTBeVnE
JL3S3Wn03lmDMES95Efn/CG5M1IrVuuI4XxsqLsx081yWD5NYlmTMFs0T+9akehI
IRtSHrlNa7PMm5BpPSMeRKLLEB4TIMzL9e3cweiq2DE6UNCa7VMQb4l9QfTkGvXO
dvuStEVTZelGEfeXNNAV9qAE6Ov6HJjjibpUqo/sL+velxfSDMhd4THulECs60Ad
ZTscqBJ+CHyyZcQ0ViBVf5l62bZau2IeiFT77DUVE8d4JdUVnaosB7ojo3M79de0
bh/1Odab77T6NUyiV2tpI6jLYnMZTUpHtz/F8vDAqQlpFyH+JKGPQLeE+/T/Ch8d
3f9lSTpqWRhmkyKEtYmHZOrZnpfN+5VoHJaLbnojK2xURnjd39Gf+NPQ2lVdV2ci
mOWzGcunq+5RLGtD1it9D2m5SfUfLypB3LAiD/Sm7abYYS0f/UxXj6MNbpU4y63e
DgNKrbPECHVBGRGUqXAiaSA4IbHk7/8G96qQIhr+laHSTWy5PwDQvfVj+EgmP9yW
Kkn73jgbkT8tTL4E+NPkGmq9rOmp58vzGc0iT6mTssmuv5gdSCBkzJibV5kxoY0L
8eHXakInNvJypm1fIYR+3m7ynvD4Gzs+5IXG7+5OY59v3HblUtkwlx1f6ZMM0+NY
OkR/upp5e8x2v8cR/REbNPWkvfmot+RN2fql3KVoxSc1/qJJrHX/a489MJO5vsgF
VNciZt0CikEN1P0ucg0y8VElYxO5vmGPnBhEe+CbxU1aeOjEt6k9gzgzjNW4kVN/
RugvQzPs/Hl7FhS+6BSBqCj+/qF80Z0cyxfiCIGwal+orLFKatp2CRuDNVzdl00y
OI6CLbku4LOxKOhyH1knCwU/0ihcnZ4byC/GoQc1wwksBW/FJQwchKEpZYDac23A
9AdAqJ4Ew8CwqHnIdfLS2c8D3uzsvYbOO4SH5gVsrQMnESh6NBYxfr9dtf/OuRix
+CeY++sT6FdczjcfgTQRbuJw+1cuAejxvhmxpMOJxK7m34xiFz9VjGnJdFwTKHpU
oXQNqoj0m/Ui7Psk3lwUS+RHG68a+BjRvjB+cOz0h+0Xiu5A6gemN+lumggmAvaa
vflHv2xiY18JJXuy/nlu1KCbGeImzuwkQ0V8fS/tZ+azI2nCi1VRwtX+M3FT84r3
srT3qzzQtZwz8RpfHni9nRjLCThkoaXQQHfZHws3qE42hScejFeASDuN5eGjjtAq
ddEuHtlwGT0yEILylL7niDpYVaUJ48gjPmAc7a9p3EhzI9t8PNnsDBgl1UTQLjrb
ivfYQ/kyZDLFx6cvu5iWyKIrsSf8KCFjMzdt73JwRcIBCt4Nu559D6ijCmtkS8Ce
MYw8GGVFd9ECkUmxd3JxBdgj6OemePt/IQbKJuT1PsAuYZT6ip+21G4zT696rQCF
CU5kr1wHRnfRETa8/6N/6d78+pMM+neyTk9KrTDElo6I5xEsfBbuccy90HjTSdWf
Tc76Q3kyE1XgkBSlIhPFQJkFltHmcH7ZKTKVDITMp8F0lBONDAW6Aqq4ASP092UH
8eA9r409lUUHXFsA5izglr1vKcgnV9OQYcIYE/JKdUzcibXk5erchYbTx2iABwuL
nukKuH1PNS+9wlFFG+yjXX7wZYhauJNxKXT6tR7BjkRR+N2rK5XdDElxrDK0lDeZ
l25LZmqDEwlDsO8ANDnPK9e2SAe8LtE4M21ydzp6QyARpfTVabJLiEhK7MJCHNrH
/8Ym8S7fTUSR4blahH+p1Sh6OQ7aFcJkMxNTDPewF81twCiGPMXP2bLHn8lye6Ws
jEJfgcXHtFHY1WsAs824MO3HCgxmwTIYw53uAVf4/S58kt0VEc2eoLDCZRh4UrSi
DOkHhBHec12yrA9Y4Q3ZIrAjgC53qfJsAqCikC3D0x+0EtREupw+PykAfyLZ9xv+
7+jjlrawaBSkTgECEtDaN/n1KXP8dTf4zw/Y6MFKm7GIcEpGxJCzLcMpuRPXPJvv
H2R5BDnyB9Jz2ruv3Bcva6CNQdiz438zhzZKx1L3doLrU8xpPguVtrSeWVl5gB69
ITh3CiyJVJiydNduDmbZEmABOJogqNMTrgeEJ334I7f1c5vyAjINlLiHDDBt4eHo
N/SvT6SzDEuHuqfn6WNMsGsU2E9RpSvDbCdWyqZ7agD3LcrcQLYOXvGSB9rwdXsT
os4XH8Z8i7QrsMPCQxDnWiaIJ07G1lCIJihPkAXKnIFNop464ydBPTp9ey/aipKp
08MJnyFHIPWnhgQCB0Q2hQhEG+V8okN2RAg1YBYpriD4cUH5VQOO2ynHFfPVasNM
5TQoHTI3USu6oLVpIjldQYIPM0nLilcUz49nr/tErXbEqm6DKKPmZWwFNgm7+2hf
A9iUf3L6fbiKl5mi1/tWTARfUtqn6A89WnuBLOw1fLcGFuqo9ZQXRQF+QtFid0dq
21dLoE3w0uW5mAr2Rl9g76/VONNUmw/HCYzwVuxZx6vRmKbN69W4lambfsmNIi34
0iDxbg4mzFoVzwLYFeezkhchl9eQNjXJmyhjnnfV9vLiEVS3kv5Qxkynh7DMeaZM
DJmt/qTJWTplDOGhJS/CRtxddGn9WH94rsrEEmpO747wfn3kjAV3rVOQBWX1vyhH
qhF9rku56atTXMoHSJ02MQSZewchjGYrqUopMywWOXzp4we2pVSJUPbIsWl7hGpF
fJ9/3FMmmn/hT6VbZYDRai3jgbfa3EH4QfBIvZ0ufqQpVbjZTf6IylgBwl/sMQUv
/ZJSa8TzJmfMA0CyWK3cJv6k5dAnMjGpLm4siA3o5EuKs+2uQflDzF9hJ73Rs7go
E74cZR2GPn130WUQ9L1Qtdz0KV0QH741qtQxNn8YWuPlO4LZ2BQaSIWMb0zHp62S
TfiecSxOIAvAnoTD7K1sIGPHZ3FLd9KNAV48oAOTEm7P+8DA9ezQ8NyM5TVzHX9K
zDLGGcBLBlDGZXj7Up/xW4LrklpJ6YoavG5odeFlN2GShQ/2z3Waaxv+5UZWBChY
f+jtD7U1OdtsN/LK2Ro8aT17A3vbMvc5Sw/Tagn52j+njhe7yqys/lkRqnWQAIgU
qtZHWffxyFyNXw5TnMtYEPs2Dmyq54DBNT0TLeqCOS2JJ6mKD0rdTeoZV0aunGsO
yDlruu6nn6RsmSoKp2ckpI8XDoeyRoDTHMbvezi8dkPoL49O+8HC9OIvKgugyy4h
gP+9CA+/4a+xVFey+IONzjmVG554/ItTheBpcH1hq1iMm8/sRjw/D6t+Ok9r1w0u
PoCc2sonwlEUgcSafvQ8PlH5H4953eptb6mJ8XpvG5Ng/LF+alpRITZSnF6kkTv3
O+0U/CQWCt1FnjwR/625fB2PwSJrFCjxq6Jau4wwBjR89XFq1KznSgVzxc14W/rA
RuwD845uJ5BlwNYKlmWZzzWUmIk2T5NOPk0m8Fvi/A0I6/BQjpmRiYSHuLEJOfr5
28kH7KAOZBymEm9K5ayn4MxpQugMMfcWJDkki/2KZHnS4ojgD/J+EuX58naoQf9p
9G+WNBX+jIjMtYlWCI4ULhscCbmmCMcQXRRdR4acmzrd9ucTcTYiTmbWe0iXVNQp
OqTZwsjIFuhqlfJpF9D/ksoUiE6t5kbuuZb1arxBFq58Do70VujNsqU2QGAV7d/h
gAHg9D5l4qBgVoRxTYzIhqdeIdI02ovR4bMF7NJJ+rCyEzxKVA12OYhJM30ndC/I
IbjdhxFsHNNG4XsDHdTplptqcQiE/Rl0JnTF7EssHHXVJ0yXlgNSIcByk8jQXXGr
U6G4pQ8I/gwEkx7KSrZaluZUviuxA50hbm7EIJq/agsCtta0OrFAM6U1VlEVeO23
243kcXvlwyDRuPSPkzw6CZV2mYiK8ZwIFCqbFGYyvJH2yITSHMR3Ap8XkohOMDGW
U5DGTFYKuKvIJDC5NtZIwUNT/xBttOLISk8DEHVtGoynPjdm2f3E70j614Oc3pyJ
MyI8cPd1Wnt2DpGwoEHLjdcz8+9ihkxES+fKpw2RmML/wjVKCcqQF6Ew0Y1ro4/x
9sWLrcwsMa885R4fMOT1mcVvMuc+o4QC0vM/XoPm7qUZ7W97xRcmf4CTYG0u/NK2
BWuQUTuZA4caDCilVAZ5bA4RbU1JijzLL9+4jt8Lljn52T1c2Q5tWMYfgRLbpEwi
r0pCfQMUk0F7nhlgQAh1h/PzY2GgxfvBO29ezRaddfcNQcVJgkG1IMgX2FI6ZK3v
A9EyWz9rnRZzdhBg7Lr3Zb7zOI2Zam+uSysOM6mlhisE8otR4xru0Sq6VAatk4Ji
Rx2J+KXC+D0od+pOLiayumOi6Uhbl+lTKK3eM8rH0oiqPx46/NA/JHf6eMcnf439
Q+UgZZLOqq6xVEaEqjw4tLniQJ0l45i7B/g9aJqsEBEF+Otpd47qkZqpCY+CbX9e
LGwck+Xmw9f/RUusLrCqXr2jtGTDAMY7rlufvR4XYWRcNBGA2O0JWulCYU0JEHCK
ZgPaDRiIBFFAtz1Yi5h6Bv2dB+bmygRnlifB3NVHjnVG8zwzYvRfpsUxB2hC5ZWX
4ckJEuBWHSjUd2Od0fjEA0ZlurQ9JqQ3wf5DgvzpmAQy09cHnwatOQzUpxAi5gII
qfdzqc4tlNmXDXBqdPJZwQc3zCWetic7zIxAtSBwoOFl7khNCyvrRMRWaF6mt8nL
EHYM61Y7s6MsMBkGbM+jdWDT4WVSJ4HedNI+Guc1r+VmDRMrqfF2xvCpheKDZZsP
IPhWb4tl90JYJ9swygzGURE4f53FnE+TPjsy5xIXRpZjoH0pazH753gZhlhXttUD
q1ypgbwH57STm7V1YdnMIae/vTG1rewvY6Cr9Kt2cU+Q/z0ob6yEdG2z5KGnPOkR
wjYQ9/ryww57qblGAV35x2+lg1x2tfCNf18Wnu1jyK12joLgB9B2pQiBoFyk1hMd
SlH7Z3+hTBA0m8LW/41zfHAAab5wQX13o1k2wiRXvW3/vNC+wZDW7GXbHJltt9aj
lTezMC5320vDoHzC8EwhGtf779cI9PTnAyQKgjvrz2vxA51C3A7j1IdekEJTKJKr
Cw/xGYSPloSr1BgA8YnkWOVBTAqREz9TXvMJqWNmUFd+2jpszPPT3n1iD6M2yX+5
7BNiU0175+gd7IkXr0xCHk6Dn2DeWFiX3DN+ROwz2GEs8DjQBx5961Q3qMWT1idh
LIIDt2xtcsPGpjVPXhyOPzNyIO1/Sp8mKBV9htlS09Vg7oP4lv3rBpUtSvUgP3y4
0X47hRRbd4l7Iv9JMSLyGYSGWImkvwL+5HXlVwFcclpK5PE7yiYDyYhodCcjcBGN
IgX++oS1psPDsFMZBE9/dUZtg/Y2BOfS9s7Z7IeMUj3m/69kgIJCcrkE27CjLnDr
57c4RugzXItjVxgsAdOV/GTXFrYWx1yk0GbNVRnsz3FFZAY7pK7qHO9oGjoZO+jn
xWAnu2694Re/4v2r9NOFLxYMrqx/qGB63hkYLSAH5FtziMniabu2fPwnQjgmOZc4
JFQqTlMuIThd+XkjSL9LAdVWq1fY8v5SbY0ul/UWSRr4BkoO70RUje4J8o5X9rt2
BTWbD+VAzOBiQIlfSynzW4b7wYiIlNfxrOOmYY7xJmJgTy/EPaxiw90ZrqbRc4rM
9+ZoqFGb5gJtBKrXJjHZVgBuAaLT5v4VFOIR+jfakkgK1VF6fMMX+dWPu/MaglTB
TeTdqLhsMxRshSCG67dEsBlwLWVDziK5HWwur26ux8XiCY4LfQaikuMnmjVOT5kJ
TS28Sn1qfaj/qm24D1KFmr8SI5k2DIZ8Wn8wtorwHewZU5IWlJoVmp6BIw1MCBnz
nqsnf4REZUEkjX0kNboPt/lSajmfHDKVphu7WCq3zo1W/ARIBCqgmsmPooKS7HX/
TtL7+QRVfiq1wGwVJeK7WWU+KHrsFrD+eS1ktBa1v10qCGQXS1z8FukivCkwSS3G
KQVkFuh2oGNwLHychxqNl8M/bFkzjnNwTBe6lR2nFgrRz9l+JrKmNc6kop/uz1xB
TAzuFfpp4/TDA88Z8uWvLravGUy7+PvYMlDAPqRfIOVJOxDPn7O47kkUpMJndEli
lkHlUXkH2vy3nLsylqXl4HzyQs1PgqdglW0I5B/v9NmguWxo2vXasteeoKia+fUa
4ecwQNrLaPDpRDYujOsnXiTSxWEKQahDlUFBXdXrEFLjXmTnlyiCLuiHGm8SWMDr
o7HLpRseeB5byg5tNaKS/qFwE83El0UyZNGPZpb6u9H8BHYjPw5v6YyIKpXy6s8q
rgNtGI37NewarW4uj7Cqhkz42Jxx1sYazH0SuryzFEwycMcdvzzabkqSSQUPaJ/W
/GxPq61MvJHIfL+GNBWir1YdN7y32HJF4usre2SJG/3bIYQuc5TaKRIJLrgQ9wOJ
J7BH1M2O/njokAEmdg7J83USiZtq74R4Q0Rg67ChRJFSJeUn2oEjSZOBXxR1mMwR
0M8LtJ9uYhbX9fxXIoMwnreDwXWsTHPTBGS60ofCnyGFyNsu6bUifnihnZIs/Iw4
hDqVnJyRB23HMsKbzlciMKQBqarZNcDAM4LwebTQDx/Wkrru29axzwzrvKPPJ61z
LIRkMDZZnlfP3HqUm2JLRBLsCRYPByCPOY5e0300DqBQyJqgkS/zOhCOIvIxgv3F
KBABiL0nMSVcQoQR/tJTz0QGEcrhXsHWxFcfM0eUSNK9QvhvkP2Jlf6N3J0kcYtf
fkkenCpbr6HVkR7HEHaAiVnFPfZD/cs4I1XXfjoc9h32RyOErlB9lSvNLuPPhw/C
tzBVj3/bawrKLaqvvu9NR2nVd/buj1quRsINWWsn/1Ka5JEBG+FV5cvXblaZPT9j
I/vAzNbKQd3gJFFEsyYrsg6j8IIkBgTjnSt170oTv3Tti84gNkqoBLjMBBip0Vlh
Hn/w4MYs3enXbFJibXjSOHDsNR92L1C83YYF5w1bD+uao5kAleSmVoht2vypRpB+
lSnGXy4wKVVHGgkwFO1+xBRfD0bvBYShzpg+IxVqlIS/d3fYWyD8nCJspmFR6raw
G76bk6vnxWmUbNw6/ToAHFNX/aCOrtHgWcNiNAyDhPEY7r5qOUKoQvYkLJAw3O69
g1qhDtuhqCebY81ho3u5CP5xUhInZbrHGyAoKiWCWqSnZiDOgND9uHu+n0zSZRH6
QL5Zu/FdUAKZ1dJZSWV1u6FgmcDlUaI0E4ZBIoUMAtBNOkFgKjioniVQEznzFcig
zRZZzZK4la9dSIt9P8tqGp4uNdiDsyzqChPSF0IUCFbM0EdRmvZurl5qt8j32Ib2
vdPzm85WFhPFjrxoJEvNTmf91XK6dqncPPEtXSsgy42wZ+p/0GCwc+YDfRZgOfQU
onYpssSKSZZ/Sr4k13hJYe8BPI7J2a5H5dnyhl9cQiFkfo4NJlmXNN6y4T8Ii4aB
Zpf++aIcElg+oN7ZSrJMlpmdtY0naHjNFvY9PKql0YJW2anC/UPBDuv4Igl0yQ+P
52+s4iyZfRxuuuP2HD5W06Oyf36BS0aMLyS0vyh7d7lCJhFSkyjCvziedz6ylkg7
HetNTNpbFP1jk4vGd94+DnpGKes+kcd0uPhP//QKIubmaCoMqbNi51BDUWY2kIE4
4hmO41fvNyM0UPuY+oKLmql+LHZ8eiPamM8IG4o9v3TC41WfIdz9IILQXq8w4Zq7
wVx/HtOgqG2wSkGsT9rCA7kYxicMgsjxRZz5Y2E5/34QTVaIzsoZbj9g+clthx9a
ycbvdj09uf8ssCYNIHMiFO1i7mgPd59lnexA8STcWHqpaUbFXU8ilyzDZ7Na97Tr
barHmJkxLDWseukb9pomJJId8qFTZbHPCzgTDxLe39pbbLF9JK4nlQfiYVtw8gzW
ycQEDnRHHt7JbPgHcRLlutKwrRCCf2hrVV785mPntBHK99OTn2coqiLgHsjYi2he
4tyNtsH70Mhp69ZpR/JASkHW03QQnFnar0yy8e/yQGmvW3if35F6mJVJacIOfn8O
RVKH8ZSQOHMp7t5B+90UtmAgcUi7iaK+8fGxGySsAF2t2UzB/ojJi1lNU1ot7BCT
/VKEEAtn/+Gjul7DLtckN2HK3JuJU8yjbuYnSSQNRAZA6eWaeALVCqL8dD27Sv14
f4TxJIb1H99GZosxAWzcu0PteTaalJXwJrOsSH7uOiIUq7PtH5F90vFNGZtyJspM
2NDZCPvieLvL+tVIRDuq603WPkvFKT12uk420MGM8zI74IoVdip7fIbaReCnqlUL
NEVOZPKfCUngqbj8fQ48XFr3zL6eCwEY3kTWsdb4MqX/DNWQgu2Rcxxf5SuK3oTT
1Z1eAYJmWswVLo6hPsJ+nRXt12hJNE+xuHGtaPTtd8ZXKI6yqw02TLp8fq6GouTL
Hu7zXyI43C3HIyMP0bZRzb2O1VOhnQBL2T2XrPR1Tc83f/cVwDfHM4/gYNDE42z/
0YepnqHPGgfzNJhgzuxsimDIXyEk3WQ1GhXzuCH4RH9wunr9C1FY7tiB63hu2Xxy
oawmmSfwJFnQpNCi7yesUu4i6547nC8fktsyauxfMCt86q2/+JSyi68bwCrifqm8
VZq1lAjWuUDnvKVJWvijVK/gWEeBz3lA4IJVGqIVA+Yp3hLcWwEDemLQf8GeC5GX
8FPIO1ZN/QCp3jJPgCe6jnmgh5QpzdADk468ic5EI15tmXdQOvmLauj+xQ868ePH
A/uZtMSEjhB/CLrkC/zFC04vkitJMO5o/wYKXqlHp11rsdbnA9sjVfaLB1sRPg65
rIFucvR6SRok+I9ORj/cE+hjVUgQlKmui0/4le74deLNG2/VlXAjHmodJBCCQkaQ
X9JWRRJL7ewkCnrnPL2+y31WsodsC0Iq69OUK40GGE0YVbXOETbdRUwblktN2P1o
5vZKfEcB8HqZ0kkbeo3C3vVelOL+Jy9FPgOnrHmzvBTjZCd39v55YcGSNgak5bHX
G6AwO9BmuCGYwfAE0MJC11SB5KVCkPGBjCTYfO/BTkDkX5pQberfSC5bGaD2cHNL
BJ+Uq9tNKq2muJHLmhFZfU8lRfVAeHxr6VRXJGuq0KYZuBS7HcLnUc7ef17E/HNI
TwHWU80ABlN5upT9D7sFE5FDqV1oxlewuWEXQEUfRw00Q1RsdYOJZVIvnq4ghjmi
oyJqE0XM/ojT2E1NsTUxptVIbmbBaWa9yXHvPkshVp4X6KmrQI1Gr2t7AePT/P+O
Jk3AiSfRQi6zEt8ChOp/D1mntDOPmo/8y+vlZ0Q0yJyKLPrLA3G8rzT0cPSrIcDJ
TSoX8aqwCTj25DStzhg3SyZ2hhEi6doJgxjv2Cm3UIPcqXIt5hIrWIxA+SovIGmi
epd/cxL5gEpYmtRQ3d9ZoxPOGQ0j+g2uDmAyCG0IY16+YdruaA6cyQSRzPXflEIy
fY727EQwujOTn0w8GGXYtfaAWL3MPX5+Uir8hIQpo0uQ+MyfXVi9I0Uk6UBypKE0
7RaoLm5csH9Xlbd/hQIfIeFIoH0cXOOJIa0mLE6+Avme06VPqhUUyI7yms7Xx1nI
MmyHFmGjF/nOPp4O61t3TaxRE8NfFAw2Edi5cnxPRfl157BukXNrL+hVhIkUbnYK
2kVU3dTvcGPDI5DB0cj0elSJ45CZn5JcJrYfR7a85kcFYvN8N11p5iESATX02cOf
3EbsuuGJFx9LbTtNIyEu1jvFBwFu9uAEyZlYmzIsbSkS0NkM0iBQUtRZt+oFVNVn
QLHhhn9gcHnLt9t5oV86r1JR4BeEYWEt/giyrtr3AJYD7JGYW8NZHDgpiZql7tii
wXuuZaRiPzYhJyyILPG4n6tG6hXmr/EmeBM1fcPP5gK7IQ4m4gpEJTzzqwp/Ij0i
r2aX5HBUUdIbCjDtlbaI7sH4nhw9sQHwAKIn7elc9ywhSGYPMRbFQ6+bqgve4zxg
zQBNxNAPUsIFfxnz9gL8WRWPc9/M1MDfaqLOTnVn4lCY3epseBuLiFsjzIgXKRL8
vwoaHnh/TGmozl9A3Xvr6dTntnZYWof2vMTybzbBex4FJoBciIGMZD3vpAj4R+oF
80COHNIwelEG+OIi30GFuE1gEBRWE7Q9qW/FXFG4IzjAET0dreC7cBrfnPxD0nji
EMJ4Jk/jjN+RRG631jGoQ6Dd7scMolFNBrGAMnBWMmQdPGXutU2MuVhUGISglm5X
P1QMheriYuXf5ClStfKFr8NogFEYe8PQCa+0jYRCMapAbxuzmTZK+2n9knFWTu64
BsR8LKjjMhJJ9G1Z+gW0p1mvaAgtBxOMomcLkRQkWSTtsmRx9yonpWiW42RMUips
H9yB6KpNE4pohDqaIN4TQW6NeyIIkJbSbJqSJpDxab2LOxEB1QSfJlOsTYCqFbiG
TeeKVuavIFmRMAnEjptVlAC/6aLbdo4SZwqaHlPwraWGAE0mI4rG9EbJBpr5NUHT
5D+Y6A5kruk+j0oBUpbLgRzeguo56LLurWE+rLyw8IAKfXf4cAQHKaK4XUVl0zDg
XGyl+EgoDeYZbabcCRbYd7bvvDRcSQSwkoW18lI7GBqyGURb4XWGSO1+mapEuu/K
NE2dDxkaoISH0gEhvYd2G6N/Em1R3ABSD3KkSMwlpRG2X7F7IsLyF4kHqaW7zGwp
NNPJs0A2SQ6xVPIZSnT5HdZxJIbK6SpZzTSnsm/s0pPArBf8272eTh/6eHFrE3ZH
afk56q/2QgnZaMT5sLLtjqbkTconkD74WhG3mf+tRgwVVcVbUjQlM7fS3f/ovI0J
a0Yw7sBmwoimafxoGOS6u53Z8QrLY2NelluPe+pHPws0E1wpi+VHXDAHZRk9LPtW
MrVMOziiOx6mtgW+ni2Z3SeW9GYVV1CrZXk6umJljleWSkb6CMSPcsHaXYEu6v8E
tg9DsVTqDeNc1Qu5uetjEWZsgPqRAPtSGJ7GCFmggWiwZVJCphEEm4xMQzSJgin3
k2toQQkyyfPx9jx1ppPF8zpvVa2b2WjxMp3adIcNf2cD7bCin4gN1Q5d2wq0dEkL
rNPXwfUCGkTxYPjtl+drlLqZrWsvDWk2v0+bfnLC/TAtZdfmFXCvV0qZVL9Ks3dv
stj7D5GiaEWwbR+GO0NRRjWa5BOUFr90sAkyFl//x4750blnyYYC4NiCzXZLh9rL
5eFGlqEYo49fbzSFuE0mL6MjHSAdpfdn0BMwEFCvLVGCkpWNjbwECqa2x40xg+fF
Zx5GBAmmJ9u0ccWxMpJB+oZXinxC2jpAB+XvVpDH/lhVFJ9uqRjbuQpornu0kREC
Yyhk0ke69H5caBRZMErPhE13RJf3/zfdg5pcOPvXT7NdNxAZG3Zl5mXsvzWrdNzk
VcEDcDtyAOAYOwj7cSwJXjCBemy+HLC8B2MIVc8fnnkytZ1Ul1mDDtCsLb1sNPA5
DyjkiYTfTSmQqR5J8PCI3fW0eFvDeNJMwN3pkegyrde0eOXzRDkrEQ/YE48jsoZ+
9WCqwT5+9Ph9u3hEDbnoeIAmWDRSpFh1BCT/SQLVj25EZVLF14AIuKGKPa8JoRe6
k+D8sYdu98zs6wCjgRWNguAltUJmh5NwRlROb1zLPOJWzphCpRVN2GE4F+35mRBx
HNythHj4BPuEvmN7cBPlF+OQ7PkNbr1+Uv+St9gU1rO7ew8ivXW9U/yqqeQWYVR8
mzRukLJHqce4D/agBs0VFIcICVJGNHSNLDcNfJT4VTTDnE51Qm7zLzLpOKItmfyM
McW0QFSQFl0rKBiGNCEiqhQw+5jgd2COs809j5ADEzclKpSm+tYvmQK5qbjfjMRo
W8y7X07i7fE6NXwul1opiiHgOPvPXbyduhU8/BaC3vaKSURJnvR8OrYViEKNbJRb
955Un304j9zZTJK07dHMhsK/0B13jw9mQIZ/eE8lmhf26eoiyAe5InuO1lfttLbz
7+X9pONonkgK/ZoL3vF+K7tphG6ot4crGkOm/RPTMi2L0RLMCvDF2tBOijpSf+rR
wUmv4HLQ1LKa2KfDBbmupEcn3bbQ26Qt4DKGN7Xj93TryXe/Tp+9pmD6u0vMYSeF
OtHHm8H6JJI9wTKSdcMR/iB/RKzkMRXgwGJEXTMsXuEhsSOmTmaL6jroM1/CPs+H
DwnvrG/bTyvrzLxjvtPGhVL0oUfVu1IQv2+9noaDm05cbqMddT77h3NJdflJxD4s
ThtyBS7CfW3NFZy9sMzqcwVO+DvZtJnz8AnSSsP10u+5ts5kY0jbKtzfl2u60cs0
+EZCKcIsChTor3oCZEl43IjFyeYxvxl6h8yN//99Rv/vfa40g/AjN3aVXPmApiTI
3ycyiubzdGk8q6AQQ01jtx9EKJvtIIF6s7HPiBnJhZiOXK/+NIM9AO7FIH5fTNnm
hz4kQ47+7l7vkzatH2MZt5iwqFfjpNCmW4PUDZADWU9zXH+hy+VTbonxvQFmmDEw
c7k+vTDZ0a+t6woyXH/jgStG6nMVZJM1R9HKr+Q0jfJto0HAaPALxs2IIkXAVbYB
Vq0jAIgv8lny9acBsQDwTCDnM6VxjRjgcrSYmHQIF/UVgvKML3580j+6wMb1INGs
3klixT9pH9Ud/UI3/iNNXs5bf89TMBUwUIqPvDTLiFSEKketMtCjDlf/5XpnO1hc
DyvDqlWfjP3lrVo2WcEl3+BGV8oy44+u9dJCHVOwQcdRKxuFwDCYBq3E6x3/CJo2
8wy9uGEiIj4PQ0l5z5hKaDMJ2UN/TRsJgCev9795FbfwvAHqR39PIgPUZmNB/vlv
jJXuOnVjJQjYs8U/GpigYlKPsORhn2uDaviyUt1e7aoHOFkSGGZtfccrMWXierkW
i+N9fyruG1ZL+WxIpFi6k9QD7m7wLk+QmetSD1PJD+mtVEJP1pwAlwNHs6EnZaoc
UM/NGtfB8G9FUckj6UbzpBLcS1bgxNErsjWyVURU/Vyg1atW9IGggP09aTENiIXr
+1oJu6qzBHdrtNYiIimJd9PUkvbAmoK2cdAmp5ozJZN36aHWY2XO3PxP2OTHWZal
BEvPmYtro9ospOFbsdHek/rsT2vjCmKioVMzLZDYDRFIUhIeNRlJVEsWWbYFqRwA
IySe1vTc0n7iA8zT+ru5a9D2ofc6QNb1snVLT0783geEA9QUCUHoWa2A5w8G0cPN
RmlkcF4o8dQ7HMlnCpSCEMZjOBtYpZGVKGm+tsd3gvGqGlr37vdTN9NsWTqtynce
bUMlVrefvT0WtMTiDgOOmwoxUiLH613/AsuWgdpCVcDaUEGnrzW3R/FFMWuBXvnX
rWqUampbqOOAu5n1bgI+uO/8MkHS+0mqbs4e8HS+Yv8+Loch//Nhf6LYRn59q9e3
vSf45YX3AjFUaGTKgo2wGCtEow2IT0627KzXhfHliqNOJNkXk2gF4wAFktpmxT8i
SGZDYArGws7y/4FRjAl3yc1576wTzwo3p3pA5jdsUvCr1/5BXykNx7cC8/ZpFqNy
vO7jUf84jThsthNfAbC2XKuCze6ExUl75metyTU/5WojZBF0KQoPimI5kefz5k2d
wtS6pqlreHPd4kbzyJqHYPLs7C4jULesLPvyxiQUrXOi/uRcupNi55UApNaFmiRt
cmMOZs79oJNMOT4jmfCjqRWS9YrknQObVkIHCEtScWVRq7aHPdSuYl9KcVDC6EwW
FAiarxzLI5FR1fKDOe1aquyEOiakLP42YVxJwhS7UC49gt3p67ydJrb2NPBwBdpE
TX5EsDbnjmezUjLZw344xrTXTlWAKbuRV+NDNC9DDu16uWPNFeUIWDGpwc2j+zzC
RuxOQcbEVeCdjfn4nXpf5/lAtZHRX3IOSha05AokweZpohT2mJ+m14Sokah2NeZc
GHXFcXsp0biYy7ujhQpggFJD5az6xbhywD6maVbRF1cQVPyqMg4pzBnjuoyQexdK
7Wkc02EgDuCA10dkvzINpD3srGrG3my/ecu6y+K9sPJTBoepQScyKCz2rXiOK+lM
3BTtrtjb5NMKUtLeESZiVYAySmHg44gbi+540PLdKrwt/r9OClXioWyYM3XtZj21
AKO6cQekHsV+eXfxG6GNKb3i+R0tZ4U8FrTz2SN+0oCElo1NxHx9GXzq4PNN6ix/
ZFQMj71DEuPq3JmLdxCc8of6eUGybA71XRnDDwnl8QvhBeumuFHlJRlNsI/bQ0z/
Sm/rCdJo/6GUILzgg+Krl7a62yun2T50bi9AV/FUT80oSk6LzCOZPIcV7Mch7dfm
e+BJceQ7QM6+ygvUL2UFBYtlP+VMG0+JRN2dsZwSsC47LyAhuKQeScv1NanozprD
xMbhCF3Qy3qg8lFb+PPRNtsVT5dZhVJAKQBtovEtvC0qZ9IcAhDDXiqxCd/Mg1v6
OgLHZEgVfvJb07hjqKfdBBrmmBx2CIDimlirXT1MiIaWmAeKwTydA1EJm8cklaf3
np0L+TW5YRCF3zuCgpa3hDJlwWo8iECIV08DaEacl/Pa/oEW1W7Z23ctbT4MIa4r
GrIkX06l4vPldMim7VBJ980chu3CmXtC2MlellKRtvM9rkR3Dsy1ULp5Sr4hUFMW
7xIgkoGFnLllOmA0+roFFW7cg48dPtSEppl/G4o+AIItQMn2K3O5vCgKwAAfAnU9
EuIjCAHvXVTcOX8nZjxmk/sMyYv7L1EZtbsxRGi2C8RSC0KdYij47FeJl6fj+YnL
h3aOXMkjwaQmH82jcOuGGIPsK2o8LGXTNerYC8ATvAu1FIk6f6SjdI0Y1MRjqlep
tryyxcOpzCz0yhObRdunlVJTrvANAKniQXG4/Z11oADJzRHlMZL0h+JOeUwuxi1G
lGu16v2jhWNWfcYwnP2QDtnpfN7ORkFCaz2gxrlYqK/nYUf+H2ta3qwhFtTyc/m3
VQZWOu3bo9jJ+IuJK+FTjVBYQGnHR53dyZtEzNII0+x+TT9GWGBcEVoAJhuYEmpS
vSK4/Pgw4X4dLgka8Pkd7Jd2cII1ex4gzlSL/f0jWfWSUvgesG2Q0rolgI3t8Vgi
lzrxi6OqN9AbsY6PsIHYO+iOJQVV/BftVEjEP/+91grvYT/IUsLfh0O9lraiV2Ek
vyX07mU8G6sJrlKXd/rypDP+XCoS4Wo3EloXq4eBxeRljzVzIvGXxnmYLi3+en9w
dYLHZENmElvwa4ecFsydWwgJ9AEd2TO1N5sOaOr0Rpi5PEVdtS6dN0pgMnSGGMOz
o2v9njAM3W4sx6rlUVYUVDw2aUV+PBWZ3XIvax1isQQHRuCwBKkIu691IhGvjhml
rdJguYg1SDmOePOgLC3Tl0HkUydYAxq3H4SS9bx4zzBALe054d4S8uFEUMV3NFnM
hrd9Cql5OiayfLVcG1K9Hkpno4OcqcNMb0mJ6bpDIxv3SNnCMj8pcM7lDX9uOSUa
L/JkW1l1A690qD8FgpCEzZ01R6Mu4n74RrzUnZS3arPThm1/cK/m7cp4JurJkR5c
3MA9ki7SFVZyFaXORdk0FgtxC/Uozo/IzRtbSJXjMuhxFA3VsmLeC77J66cRO4J/
nZiH5Si+D7+YU6u/WZlHpOttM620ZJG7PnTH3WGHpv/mVAAAJR5aoO6DMYx7u3jz
XTAdJGt1mHxIVp0P01ytGCPtZzAp/jEWnx/9OAW5S+ss1Aj/SpsSU2zK1vV3UhDQ
9ThfGJxgyWjYCBlntBmKGnCTFDidsK9AUYSRpcaq1Ql8bFH+wa6r+28fMZEbFLXz
8hvKdwXO7dtS2K3aEAIv7FbeS37t+GSqrp5VN7YAumTcKe93HKPzEir+TGGg+sbP
7PXg1boWGM0nLd7+g9uHv0S5uhwTQ5q26iIzgM8MRgZDlxe+1F/MqmG6pI/00HLs
vPQ6N1j7MboefQ8WOExvME63TRZEFDhb8fPFlx9mY4Aw43ZSsyZkaE5qN7akqicd
VHgH5HepENfUxWpOkEaVqxQ1MSvBys7fnd9gKB6CMNvhxaaVI3csZx6HpDY/rKQy
3psVKjJTRqXyPUtjZ6+xn6MkJNlpIcRa9LXkzKggQew0otDCYtoYsUnw+/Z+soqY
Rg/t4nZgrHLCFHkfIiS7phr81PB6KMNRNetTJCfGWlPzOQiomgVmAnfn37C4quAW
c7umY9XRYbgo1gf44ew71FYiFe9NDzXK69yLRqLA4MfoYs84ZUcIdUG6rVM6zg4D
RKL6lGw1Udqaq3V3UGc9OvnxG4clz1D01XOXh4Jk/lKqwyLANUMgAhSawsImzdJq
4icJEq+keDOffVDbQlJgnuhc1a65ef6z7m2z0H9rCph1dN43oI66wXu01tIzJeUw
ye1sprJOu1Zuqlqk+flj7zZK4MVDgxnQKmiGFcvS/i94PL7OQM+nqZOKks8j7Xec
3BLr+19dnhknjAhXCjy/H9In+HtLKBfomyTZLyaf368tKruHhI+NB70QQZ8Gkpwo
3n3mCIPk0bEPpn0mPGM4UkS1ICFYsvgYVcWv2DIy+2Q370Ebe2qtAdoR92vCGY6d
HU57D4JIxfpkVhVenLcoNrXbs9q25qcLJAUEi0sE+gp64AEBh6tPl8RAFXsQK25c
JbCw0PdGMawmOEG47D+EPVw9O06sWpdBPMDN7HeuxiX1Kf+H3Ftf+83EzMmwzGaX
ToRGGczKTDn6r/UHd6J1skNFsgQ5D+D+Hw3qFOmVRSHxbJCJFqkTmBNHLD/cb0zb
pt/jX4jSGtK8z8Dv3k51uadb7JNZhXvUwre8PY5+vGGWXGSDZU6X3d5E9TC2ig12
WbU/qS4QOcmYo+dqLxJqHvZLX7W2a7zpRd8pcZPTIA/q5XLxb5sXsZPzoOU7yF8O
niWVekTLfBRLk3rvZLkwlmAwaD/dGCOTsqwBoRSngiKunbmBuEG+REpt5ITM81Ag
XgQtnPRBATlxF3LkciISNCUBKlOoSrtrzaPpPiBBofnsg+8wkFVy7eg7I1Yh9wVL
7Vii0wC7+be0ElLhNgmx2npfzFGSLvmxK1EZM52JEUIaoeTZ0dQMj3vKnOg9MzNs
0iov9qw8ZUajNfZsm7Q0z9OtnPzgnKH0xY2/NCXrt9RWUWTLCR4YhG79ZT6AytAQ
CGejtFJMBngbMXPAeIEqScf3RvNWsJ2RUu4cCPVJ8bo9t9SMCRgPfArnIXEiiB5o
ChDt9FYaUdGuc2YdQFuw+ZfiL2V92SqKtU++Q+FAO3J2Yxxv9E4V3Q4dn+HLnyew
utI0LAR/K3xfOVb5aFzcHJbUsNAUP4qzZ4bU8u6sZ8GBThDRT8K0bKJuFKhFQg2B
Moa3lORJ8BiZSyfTfopOI7d5ok3j6CKf2XUt+yfZUr4EKproqXdmybK8rBxnSqnn
KR8nz+AbqNbo4qTUhrEngs0wqCa3+GjWQEejAtjKSXNB/tXv37/1gtd4EPJSVNaY
AnrXgM8ZZw//zrr5Z2I3D7qlhdvrXtsGkExMYoGdEhOX3xTB+KdJrH67KDH0SHRa
zPABaoU8QASzWol/28vBfzGnag+fWw3oBvOWANVpcIh/R7qsVoqExNCv87Pz8JAb
uWkZaW//fHmbh5K5tC7W9qHuYrtWAmvgTHNDcCEIApkZBVbc+Vkl8NH3R3GmvU+l
563CfkEpetvSnESm2MqieaECmYYSEsscTnzbGH4Sk7onIPNDdQMzbUYuqDSoxUHF
paYiMFi9fLWgapyExGhBIm3EcWQwsQLi1XI77Q2GAEjLqspoFtifv57N4Y0/gexC
Zw85TH3Np3CJd50Q1mT8ZNEQFtqLo3e1V1851eK/ecrVzx3FHtjfdKo7Rv85/kKE
gpaZri3RRbuwZYaCja3Yt3J/+GjLWH7qajjcVngglgj4yemrgdOEwv3pvC8ILG60
DxBE0/PzaNlQJJuMqWWxu1u1i1iBgxnVFkytup9dW+jY6qg1/O0QXoTBJwr+IXR2
s+c3zXDQFz8yr0lLskCALP89Nla6E9Ax0RhkSiWINL/UGrRDbo0vZJuclJFHePYn
EhVb78F8ZikNfLY0fg/xlyCIr278E1h5oDjeTC8bbbBAclDHpnqbv8WP2WEsagXH
GUNXu5/bGgd4MgF0wyvaqn9Yh9Jx7+5dBcRkdbRfrNukertdw4eNHA5xDv65MmB9
ZP7aIediJ9DU1QqzoCa0sZUT6PbsNResrw1lCQrBeyB0OCUjvS80cDTclONhbWP6
bcOjnQL8Rw04m14qgffI9b8CjyDEpdLaM6JxXc/HSwpGfi8VLxgI9OQWXAnoRQGC
/g9gq/x9gQH7oCLf65j/Tg1q4bu8v13zP7Tl6MFs4v9+2i/4HbdzGpDeFhTRxYRX
hjV35XsvGj6wR5ULxcaHpX85EbibHLjYotJy+Q0lRGdvnwWSHJdTk7LH3HOJstCk
y/96S39qyYqL9RqwE+od8nlcwYvg+kuwfoGKf239Tg/LIYInBcB0hPIP3eFdJkNh
08qEXVwS1Il503H4f6Xrx6CZT72LnajMXMYS/0nJCpJnfjLAKBqy3vFBnxs2HsDV
VAR2FvCvBAR9wv41KSVE8apmz/LAc+5gkdSf4rtbubfYLPbDZNZzfwH8Io/d6/7I
CZY21CkI1u7goEu379c2TPR1FrGxrTAld95RiCKB3Qin4INdfL7xIRF8OD9GwSSV
jb0pZFugGCbEkIUBHETv4Xldd7P45sUV3xvy3IthKV15ezOFZL4j/wkbvHR6Zi2P
xSQW/SOaOmdWp08Y6XOgo0QdEigcCBmcruHNS5ZBSrczlfhn2FeNZKp2jcYCdot5
RfiH0sXm9SdbW2lRf3IZQx1BN7bxJSIFkbRdq5uJx6AMJVpX0e8VdGJf+APOHSnu
9baIa2TNZ1MfuOumQubc07pTb+Vfokckz0d5Ba9yzcrmC1SdApewBcRCcGtRYmv2
JKMWLMOEPoASQSqh5dpeKsr5rvFh4qvbRfRTqCfDS/CX4brBMM7BuYQwnV98PyqI
LrKv6YD7HXczCzfN9EQVxGNZIvPW6EN8TpmEeUvemryNHTanX2a7AkoZW5p1f2K3
3DsalXNr6EuNnkG6RkeUciNVWkwS4H8RwQZdaOusSzcA+67dBLVyiWjAHDfzihNd
Om/tk6H4LbgDcXM7j+v+oata+ti7BlyfMUNmMY5NdU4AqFlvJmzzSmVRezfKlLWf
pcn6ZQ9/3zKFx3/OKdLU89yaj6ytMHHCdDl9l82uwdwjFkY+Ly13My5qxO13GVmT
/zcciscaIVic6PxwaCNdLTC+COE1eIAf3cOxpD4xtAs6RYCHEx/p4XY6oToFiQLp
QDY0MUhhC+ZjGuGbU+9eLC7BwTFM6Z9IAP53ohjmNyIEY78L1x6TBFbLYtaQGo7O
Ldo8Z1kwrhTstTqP6FKUXNH6fuP2fVerfW2fKglI8sf7uDdCpBLP5mEDiWUnz4N/
L/FNYL+v3n+2xJi5CxLvV4RNYryRRpO5Tg3cg0kGMChtNQxcDaFYHWm+acCqKAKG
gAJ3qOzMmNXiHkVvuewaluUsX+qvAGt7//JCDXJX9H6yhrSFh8PZM+CtkkRobdrA
950bfwk2lBRtc83tPFBxSivK8QGo2GYRoXpAwGB1XeOiEL3lJQPPcyGP7hQJj4w6
8F8t/xCal0P28n26wadJSodjGbuCZntIvw6La58LAurGB7gUsUYwQkj2UhNQo2hJ
HZbAixjnL7mECwGym4jElqszWpPOBhBFRxEi19t0C6w8Fn34F99iMfFEZYmqSB6O
afdhvM/5/+q3kkKd2IK4dv1ZeZVwo6YZHpH0mZ1Mz6E4Mwg+8iaIbq5R+ldHoeBB
ck7ic/1PsIDLnTwpZKvMGsyKfFSGhHOI2XwH4KD7etM+dfRYGWKuWAnyQQmiT+7Z
w38H7PaXCvHnOqu1e5ZnjVbGFBs6gyJpRdO4rY/uROi3ZPsW2+HdK54K8Cd3Nloy
RMvGPr7y15I/l7PglFF3R0UHKhF4z2DSoCojMnWr0gawJyMgF/35XboMpU/2PzHY
RDaWLLikgc+U9Veuno2LrfsMP9cpd2xy+c4SORYoYOn5ycluOEzxeQdDbTntSzEM
UBuVor8rs8gmvNE6acm0w2MIimHCT8vnKvK1mxX3kVdq+qfZoHGQBsLoXoM0z3HF
hCQAaOLum7D+lH3DZ26VqRVYllL95fSrBKO0e2O0JA0wBjfQIHOYF2Za9vQSXbGh
PCZhIsZ5cc/WDoE0ahCghwzIp2mF6wC14kzRERxfoYHRLZgYOTwT1zm4U+be/tZw
Fv+oQKuCZ3YOzC72Q9S4SfFu25/k7WxLmNGpfwIPIZ16QijZP34Vsy2XZyOXA8q3
fTmuM5f3Ptze7KrM3g9/pgRKd6flQ3jwCW/okSfaqvS++8oJ/OY6cwFUbbvEMlEe
1F0vNjc533s5/LjiBVdyTcm9jooUGuSMUlWo3wJ9cgI+qpP7g4dyzTomq0+JQqQx
+8A5JvdinYP02mldoU3/0tfCowbVZ0eI3VfRw0kfLzJHY9+5gAe1pq1BLeZTpuKS
xeYJO/ihiC8X+URIIdLPDxf2PpCtqNnylbU1iJOQ+BkzjVepFGzhuW2xMQ2rZd6t
MayNHLbiX0IG2k72DIW9ZkYNgD0JCryeSV1+c4PIHfFlo/1pO1rs5N8hSJXLsmdh
B/7lXMZ7B54xSAgFZoQgJvxCvRbM2Z4Y3p9C6hxtGoxaqidRWjzKTsBaL2izR8mf
6O3/S5q8m37h7BA8GtdTnI2LrPc2gvgSOpLDwsb+S+9/cYgVlK+l/3cK9/aFkWHI
z7q8IlxF3lZ2LBkBS/8kaIyAOOUBmmbaHQO3JmOykcPvaEIjmmWty41pEk9ZXELM
1EfcXOfUycNhL2Xr+bn26ta7b3K3qF5Qat2Mt5wPOkbkZKVnoxbO9y40TT6/krI0
WmFjq+qxHqrNeYc9vY1o/egIn8a9Ai/bS7HAGHglXWKYPMoDd2hIMKhD7fR6kmyn
Hdx1ZNbqsmubnqEtLR/ga9jKZDye+vmWwKP+c+MXEvMlUsPPMBpUylKNEpBtFf5u
HGYV8SKz/yYgrzSDwvfvRWTvz2WhpTQ34I1o7DACGv3ggvne2N3KD+7CEHIaeYWR
8TRjd37pP+1yheMTB2Pmbe/WRBzXJSu4CClvDcWtA6gtlaEWQ+PQFhnaWeXXvnbn
3vb/31zJ+miMJJMsNI6sYz3uOAy9w5bNyKy0ayct24/NiJvDwmweDcScdhW2FbXA
zPubnKZ7/MhJapTl9+PZRxQAWRg5ED3YmRoCOaS/Na5yW9n7Ggi48n7njP8a75T/
zNfHwMGilwYLsON2i4orr3810gXrPElJGPVsdWthJZsn8+QtiB9WH4hNJLT7+O0S
WJL5xRDsyaPJy9gSb9UmXccs9neX+1IXOT6icgsE1zKi+TUi+fHkC45yR5pG/9kA
jdCDOMwdFfgn0zapJepay/6sYzzDqcx0LlyxcEiitHMCUD9HsahFJYQkZvsckDcg
37n2wgbONBfM3WqLDqTpECRmckfOYV30eM/wUvADbnwnjDAy8pK0QEn15eGdGDYU
/Lf+dSDfDfAdX+Tw8ynzazA/uu+FqtQmgonQqO6ElTzSJuib444osx84rhdRNW4E
5+C138tqNkl5dX537rlt4vIty6aBB0778jr2d+YqZSDInQAPE9GCifsr9jR8TT9c
QKKlNZ03MJi9j7ZB47KiZgajse5UwVG9vqVhFnE4lcP9klSLx88LlZ8rqzZMnOsM
SKWgQH1O2488A8e8E1ualCvAy7V3F3wXewwcAQTH7mF23T0Tt3vb7ftptA1w7sMA
6CJ0oK/YL2PfgB+MPpL04s0V3HTjShmj1wvsOxDE4gxBGgB/NdmAFc4mZYYWxx5o
sYdHN7xfMpK4AlHcfmyqduL3zG7cmZUq2+SU4Dyas28O0S+/Mqsccot6Ykrt6KKt
ZEaPRJd4g2OEUbPj2bFJjKF9ZahiBNKpwfjjka9LFNydRSjKInY1lmqoF/NG/uOz
L62yRNrNVZM5/1b1QhoFHWolT35JPx94vFj02e8MlBPKFiTEBBfXPmbX/WXER+Ah
cy4X7lXBxF61hnSzzshN9L7I+9vAoGjoe4u/ioKKGnQ7OkG9m2+MDhusUhhwA/xa
K04vTLGloVQcnh40m1Dw9f+dzJvWAZfxfBFvnYCHDuacs7o8p6iy3jR6iTr4ODvG
hQ6p5eGGoaixlUAGfykR7+mIdneTUBsr7b32O2RBbxCNZO03jbvOErI9fmBP+taW
CnqL+6h7O0FewYFN+GX3NOOAIP6L/8FBID5MIEpeu1DMEhjzz0eJ5AAldfcTwCzQ
6Nres+xOYouQsLF/wt0Stg6u3H/3rKXdwb04EOlyWMe0egU+pEb9640ufqSBXd9r
RZEhSrnuYdp518GNcuRQRJ55F5CsCjhRGBiH/YFF2scoEz/AEYk9iiYA5AcmXJMs
+tsYkqDln8d+g4VFCx8PsxTVMFcEuuXqwelVOdSX/rtU9votUMjobPW1Rjc+8PWQ
a8DldMZDEqmWUgnQCIjR2MXWFs/OAwWMyghOKmEWElhxZljsj8SA/e9g/ba3ANGj
Eb4eIFn4ieUPAUc8YD7j5l1p5MutRTMtlYm/Uy2jwH0hs8VjJatMAdt0SlSfG7+S
irG9MDOiswAoXyAYlPPgKwibB43PLaWiCABtWDMHw9NaJdkm87GU/OcA3Ry7LROu
n/zDDiU7yQDdOhQgiE1CFV6q2cVrkMqor8hpCrnRO8xyOy1A4PbwEqWhliGQtt4o
yi8RPioc24P++84lEIrXMroX4iUM31WmVBNAxE4wiGVmd6enkvl+8kOZdSsCJivU
GgJsxHLEdkHQXPk4vP7dUTqlIrDCopLRO3yc2NVCzyhcbcM1DcOlTQnf/99ggMdY
4x15yivH/Fuo7cYLhAKTHK7b7EMhimr7NCFizGFHeHDayywO0Y7Z5rubO3msudSR
zg/NUkZrtTCadX3F1SPB7OrVgEVacuYU6qGgYF356SK0Sy0nTvoVsHH5f+/FmYUP
D5MQ+3se8KUwwC8A+MzW/snpWfz7DhcY7NJdjDwnF92zJm3Y6zyaNi7+mfEKus48
TkeqdQJaWBqOo70LhKA3SJrN94yWQFdz8P0uNDatqlP8KIyoq6cv+NjhkggWLEbp
8ztv/PxHAvUBtXHzrg4Z/B2CGBxSMR4oC7zAHOTQ2l0L/JBQutde9heTbhz0bGqb
K6d0OK6/8ERDlYNXz6E6ODbnDuYj6lk5IlWd14xdKvoQpJzg+O5xjuxnXmr3b6kZ
J6Y1eioL8HAsMa/4IDQTEtCQHMfA5zxuP6BnSQBc+NbdO5P3tpBTv/fhFTM55WfF
Mh5M5HmJ9cajEoats//Bdr09FtwtPfnCB1SMxJM9bWeyTt55w/j/hwbTYBynfU0y
6OvmnJOGNbHmVxkhISpFJpmLgUliHOTIHMm58msnUicBj59D6zFqbJKNL4UsovkZ
wPnWf765eOU+OvC1L6eVngFkIyGEHriGa0EWfAchUuN29QO8g47/A8GZTuFWhluB
v4akAlYn4edSxB+ySnki1niDg/i4rn9dVIG4yDikGvW2D4kYrU3z4OpLrO7g+Qi6
fNegpVffF6HWbxXbT4rtjcC0q+QrE9iWwX8rcJ0g08LBHcfX8Y21KTUfBDG0pG3i
wFj2Ko3woN6B5NhKtJX/vZw2hSm3VbOC0P+07mGFBaiMXRyXT2tdJBrf4hfrKlG/
ETDl7UnfrjSqBs+DORkOZZPLszlY/sEe235DcYkP59RSSgqSjYbWU8Ch3e29iyfT
nCiDViuN05f6aoCPnSs8/WO/2Cd83k3vrIKLbnqMrg2Ekf7ytUdjWxxzbZSZ0pig
yOn/e6g/BLJJYucVnkc9UpAMu+B2pGX/JS9ynPA++DrCvjWqBRWVqJXpKSlgXj2J
cpElEqK1inJ9GsItd2IdQwIWhHHnX7h3tnii3rVxlq0+DXfCvJYmhM0PYoAzwZgu
AB688L99KltxlnmigQ4XHsjahczcfrXwNYtDEOH5Md+Na94lAhSK1Oaw7XsvoRgR
FZiWXIlnL/NNYw1rY664mjy7kPkp1zclPp6pqWEObV+Z5YuVbAPA619NPkA5zqbL
C66Dlstd6oHc+CjiL8YfujUqJ1y0UKTa8CcYySGJ3w99U6tTvaq/P+mGm6uzkNmt
Y1M/5s9hoRNpDY+Cvo1oPbuLQWeTsu+j5W4/T84yBXNYfGTdu17jZ7T3oXmF7sG5
QQKHueimr5eZmL9wACElcS8+3olrjO/Nkne6SdxcK4aXnFkTGHDLnzdhG2ksUYkb
2NVTPjTZjxagOAS0opwlhD0bJfn9oWdU69RaCVAOKJ/1UxGs46PxoXnw/i04CJSI
+K9wkT7ul3Sz9xrZZMnhk1TItbVZ5G/iXtPgcmlxVD4FEgkRp8u5RSwu6cXaQ364
u4gWID5afsNSFY0IIzkQPHdoykU+zzvRJGp7L4fGDbtNx1d2fUo6bJfBJjG2z+6C
y8sA4mCi6aD3d09nD6w56eAGgMagnanGIN3xJBRHS25YWIOiu3K7zRXTN7FwyniH
n+X+z4mNrcWIVA82rMWdIBoVI0V6s014ttHp7zsO626HbY0IQQbXMj+K9lAxyVR/
CnPby+vd4EEls/yKF7zek1Mzc9nFfggaO6q0kXmbtnc2HfW6O/HFBu5LeoMEpNmO
50gaHZqjm4R55jlYSNV9r1W+JmlVxoxddT6BXEF5xWwLqwSEaO4IuaINmYK4+a+g
2ld2Zbg5DPdjgGvU2XQjnBfXQEGSz1dZjsXyX+873fWfeOnaZ2DLsUdy6mAAQ2YT
RvqEL9btO/1ogLd+KGtbILo1WRcCCFHRWTcuY3KNMmX47+vDg8QcWTsLMG2C+RcZ
pidmwo9Kn7dwbM5yB+nGBDOd/MVLjoviKdPljB4a1no4ZSPUqLUstXDUpZEonsq3
NbZjTs56UTuEaBMcgKRe3sAeIhZZ4lSNz6guTpncwDO0o0YmvNM7ZZ1xnUGdek/T
m9nZbQAzT6lvrRAYS88B6eGEgwvBIi0AeWGQyU2q7GgWOZ0KT5CKG6Y98HqZI+Fs
ktnGP4R7xdQelKVH8DIqCydru0Jq0HYdLdLEcyAJ0BCUKyNxhhOrKgsx2j3DIFTd
Z7oBXjcvRyApBoYTFCgqGHJK144QYGq5tp2NFz3x+Qly2VsbcHQkg3XeQbZTn+mb
2nHv+bWnbbWMZb8xjW6+9eB8K7lxO7jTrIjuAGqscU6jtqHPyJt3pe+twCT+8r1r
nqrjUPcnpN49C+VbUhiXWcYkx+UNHre7fGdvLVwe5jqg/ZOrynEn3+QEEwIEBDEk
iTpKUOmjelcME3oL7okWP6cq2tAR61OlfQwx7uO9iXMHGgq0NJ5o7wfjY9ExfIOd
k/q61YiL50zv+ecuTgDUmuM73wOWIj7jKB2n9xXZ3YjpeXP+b/llQjvZALhx3cic
+xqXLUokc0SkNnr/0Faa68ykxrbRmEBLE5gk/zbGSpFnV4gK6XiUHnOrTBZlXwIi
dyGPVC1QP81Mv8/wYi+htZuP5KtrtjkVtXgNAVTgQCa3bLL5n2EApf1ooPjDfyd+
VvjLmHQLcGdOrSWCj8jmRrGHbV89KIDCye95jWLO1r9x/k4h711gSCZTvtvJ+hOQ
Hg6iqK3tAO4djLzf6F6HW0+2d5ToWROU9+Nr0VvVv6dP0/BUT4JqZLfaUsRSGP3Q
z2Ochnbo7pXaOd8ruKdACoQ1Ao4iPOjveCDlJISp8Y+5oE6OVKZkMvjBBlCxJFm1
qPROEHpsK7f+VYk/F9MUPj+2VJodVTejxArcUL+kr9shp+z2+7ciJ4cdQNqOC5TW
r+9Xg/pOoRBAao9UJHh6B1mOPEPn2v+P4cyU88UA4hIAS2S6zjcJuTVqjBbHWKIh
0IeDYB9uAYjuomu5GgDiHKhT1JZVM7WbCPH+GX4xDqxR+Y24yEh0vqZF3bTY/WAr
C0NoAVBBCEJ3qpD3Ocf/tiVP4az7aVphQc9+VcSgzono1tMCYVdtGjFBHI00LkM3
UlZgikca403mb15VGVMIfY6/RdG8LMRxFzZeanE2B/Z/kGq1wOoSxs9jUmEDbZi5
VKXaiLqmb2mQAQvj/CgdLAHMVs1BxnzmF9Y2TOkqDEDTTrCs9f4XcZf13hYpDg7b
RW4BeBFIYYhVHltaYxO2/SQCAr0euyn4/0xsUEKdHVZV5fO+0ljzfhfOBj6u5UsT
TBvYRIA8EeVdG7wULKCZyVxscEeV+bvKwgrN83zdFpVI8+PhNB3LuvGUKmmGF3zk
L413tISkTC6+04BYLOmLBUvUsmipb5MRrdt8hHFFZW5A33apuaQIkThuuUkHXw5d
xZo7fUpZOgqXo6QsZsoWDVHlX1nExbhgsT3q8W+6O0IMIvVrUqQN/fPQJQS0x94Q
j3DtXzSLGphL6C2dbmf/t86qZ+YQUNyU36MaPkWQhS103/FOMfwy2fCCG6BEIoOg
C2054aHjgLwTMXHQZh/p76uinrIg+825p3d38o92+dnVF050fuGBsu259cdlnw8P
Y9dk6qYAeBNPqiMV8mIEI/h/1Ak9AmmRFf/tmMzh9sza0YIIHeuJ9D9A0WZmf12T
DtR1CICfEn1Uhfq4XM/Z5ZFGE3yRLPjHN3FsQjQ7ANlgtUGVsm5C9PD0buYrPP14
w3pPFzPJnrVlmjRdsy0rtK25L3YDQ6KmrSain0RzEwnWtUNxFa0lbCItpJEUW/6a
ePg7feJTyTs9Akyn6RfWIvIduvqmisAHBXM6LaX1suqZ40DR7i+BVeYDJlw59tgE
PuPMVGJ5Or4QP3y8Ak04qaDTdzL2Cu0Ejtlx6irLMohVPT+DajyPGLbe5dzbmQUJ
AbPWc8NpvcmXGMGo7Xu8DAonYLKI6gQQuVpoNKbCOi6R8Rei2N4ywuRGMEFS+gaP
CkEP1gBbe3Xw8ObRZFtk+zw2TOiQ8ZY/Jrex6+/KZ3tqkpRPOQ6NB4fC9X13Wd8x
anOjh4MziP/PoD4q0WD69I+gGKnX7DGbLAG5+2W+/TWFYnsd+X23o3ZT+OeaQ/vY
+So7KIaYhsOy3f68/aEw94LZoF+D4Mzky0dcg7ddu0Z+UvB5ZOuQC3jgW8j7FVzY
R+xr/BEa5r/fe2+J8G0powqfn+wc32uSbOk5+Jff9iyD0fPXYRcVZeAfAT3l3MCr
28lX1fMMhScQ/4n/hZUIVanEuludS8hXQMJVLSXMB/rV+ezbkLSHqwR2Jgyn7Y+7
osTvvfIeRCkzQmwD88GT4W30I/mPcxMgOAcxPxHWPlHL0H8PNEMtfwjUbGApnyKJ
0/Scnj63Xn0d8iqaroe60bUn5c4+ncB1H8Kgy3zrpvl/o3yrP3R2EuWUQkCBNSBb
kv+w7HGI0iKsT+n8jyzOJWdkY+79JrXCA9GFYUdxdWW+H5Hzs+OYTdu2OqfBWWqX
4r02XizHNvuLl828oSWPnQTz/dxw4qp0u0haorEpF6UN94TRZfmD3TXzmLlfPHzD
coz/Ek1noKCp63ks4h55d6e1xOtydw3ciIfW2DnQ1p+hJBJeM/VAKjXmJbM19Rs3
3I8tvpWtJfqBCoReaCOvi07u6IZBxlbi/0MGG+UB4OUCmJKoANl9YSozhwPrlzZ8
9lEwo3F8UjQekm04xeAPOuHAl6dwRBHdscgXckuLYZaWMGfA8IskYHcJ4Thzx4IF
aIkXSvBW9DDV6ybmblq8EFKiQ5SwHdrJLo+qSHDkOTHeaiUYaFcx1RxbuTEvcbLg
aes2cek/pp6XDTO61Nk3zkwT7OfCax4D7NRu2NUEVvzt9HwnfE4sbERg3Xaj0tQP
wzmNjIrJ6VrFDE754+nn/D8fIW9fbcMpBdV/wblhdG8VMkEPcP0EL1SNTBvThmDL
xy5ZtLbtHClVSkfmgIHjI3GewpgELf1obPzPqkwYHmngw1Wk3WGdb/cEqfRxRiPk
wvkpoTODsff8U2BFbgKYR3GweDRf91s9myZ20iH35wURJHt7d+IZe9Y0Xb68XnWd
7gsQE6O8FENlTbUPZOFY1lNzyg5fUnnPhuDWHaSofuwndaWKCskJywgSBHAYSHyr
3rJLuLwn0HrgB5C2Scz9BnUVkNHTQ8DxlH9iQ19NEEEini7j9ydRVFuBe7o/bVMT
vS28F2/VyoUb5C9kgy4+Nu94NCtsc3OjPN6A3A8Kq68Hph/7u5XJjoba1RgbpWJ4
ytTG+EEQfoUuXNqNKjyw/BvN1tMb0TO0ALyjzPwqWKgEpx1WltyWii9PKX0IrmEg
C+PXeoyAKSoSL+qx99rbDVgt+voKaDNuSBLcyjC07u9SWQBPUH+Kk/adjteFSQPi
ckN53zMddkmf2Oc/MEOK/h79LBYMaqubPo1p9q2O/ODjxLx/FoSVyIAQkRdh9WPX
q6sRmxQZ4xjlRk/iJsXDHbV+WgvDodUy/WqV1Jz4IGxg7M8WERnxQUK/iaQmY5CL
KKLTIhCZp3INKvGU6RkGK1V5Xgp+GdM6tcC8sgJZaFo98rNMmzSXSb1ZezKzwZwW
gwtnAuuK4MIi6+Zl6vSjXQWrEt+6RZ+ke/sqS72k9kOvM1EU+8C3SKKto6UFyzX/
4B6EJdfuEyNvcX7LN8z3EgdJltvtzaEhlx9sFbASSu913TK91ljGHr20o5f/Y8rJ
OdAHP0Exykr11UfXuJ5mtv6bqtvM+2vb5zN1yoRq4ornAdh9H3h5XS1FNxZaED9f
Pf1AhvSJWX89lPjY/P7c7XsvkV3hxdMdABYuTPLw0Z8IrK3iMMyOR//nLD1IRyX+
c3N7U6oKxasdKGCIQBQD8R/dkWHBUirsXr2aZSNKOjaZSnpEfcK09N0tE8eF2gLX
KiK5p7Id+/qpNw4236IkaPh+dDLMFp7ck/BJnXj/rGh/9PoSlW/WOliJy28gx2RZ
0+9Wl/6JBP8EUu8Nh7qwW7wOmcJ2gl4aWkj3KUGWkDogsefTUKioLw90tIG09FJT
BfpKGRJoCu8nlfhuKMLs7wMXWBY4KjhaC2J01JgiOx72apBhDB3OMjBAIHbVySOC
Trbk2VQITPVNJ9eU2p437oo9dHRoY4GwViJyAnQA49kMIw2MB3u35HwwFar9xUT3
9ykboeR5a8+bkruPlYt21KseiCJBx/aYlmA/OKPVo24a3xC8C4/Td311tSlq+uT2
rmaMyNwKq6hJqTcKHdWbaLBuyDyniDaKPbtTVWj1I76bg6qv+nGIMCy9Bj1ejA52
5Wmm7EEc2QXfejrg0ABJI66dflG91Tb8CW8/oaWy+dSg7hwi923iuf3EDb9aiZm+
+GJPsOLWqD+APlOIV/Zo77FrYBg5v9tZm8S2tVx56WZZ7YMz0cZlwbEnGkaYKvAq
vIZmTuexTPxxCy2fWC8G9IQZ2HFgRokyXWUik2M8ai7iIZABaFl0vLwTHIKfUeOx
8cvwELZkqZAsEEuBzwJjyCEUjfavSO55ns+oWQZ37KSqxLb2oOIOuXvh2Uc2h3di
uXvcFqcx9COyW6lw0eh4wP9iQcCusZlXGRE1rHOGL2TfE7w7O6rCiIp8GE5ZbArP
puJEvaKAkjbofRpHjB2pvWHAEJDaoeTFM7nH2VYvANC0lV9h1uwDZG2t++8amXKp
XlI3YfJqW+139I885iz+EcDFHBpKBoq7so9JfnKVyzD6dJkD8T8F5CvbMF3UsSdo
kyNK4mAkX3Nkg1HBpZiW0M/Z26QStz1ANavOB9+KKe5yW5GVR6/7NB6Pcox9q5qG
qLUciFkLuC1liVxtFoz8tmMmzJ1LO2k9zIH/hSFEnw87fPMbeFnPAIkg3wpxoSKY
h1KBY4udTXh+nYyNT9dIhVp94GynF4MRD2vEzURMSWVo4kpzuxgTVnTQYO11dkJO
zuz3VOFTEMpcN1qDcU9f6EakOhkJ+WxXLjJO1v94KOCOM4Ga5965yoFleiyVsAbr
rph5BYQiW9y9uOcKXghzGfe+6Dfx2icpR1H9sVOGZgNBSyAgtEuX/acnYAqhx43B
RtnZGAmLvHUTpW8wN5w9BGoTTPBcVZE0bEp+zFI4hwAxvYg8j379jVoj1xHRqMK5
ST3n26Xt0v2iov7h9Y8x9v6wVbTyovskBvj7ul3xTJHWzAPEkIKsRT0R+WV+NebT
boObuv1vgXwlb3/0U2JjnhvVvPU8H833zRh6IPbMfdR2jymA6u2u8+pidmBRlZg+
geMj0mVJcOLvOSee35etVP19uvhZE4rNmznpyjG7L7tExJc6ZWJrT4LsyVhAXNts
ev1Teny80TWCCcekHrSR+gHQrx4FMqkairHMsCIXmCLAgdQP2aI0M3KlQvSNNLxa
loVq2OxFi3xz9MbH1zFrOP+oJRTwhUrM2mQX6UaVPKVKP2R7qO4sO8HqZF89RJVA
ey96PsShJTNCnIo2taOvDkbLHnKl5Fr1Bf17nZBZyhrYHKs144/MngZDNAUCvHDi
N+IWoTp+M7aVMQPnYKh0mZh2dh70qXEk4e/2Snbf4MkJcFi7qcCD69pf07yvYZ0k
HN1NkAlLDdA/jeoplOJACYrjbO/PEqzYTLDoVDiyagJOXN/VHZMI8S0A71ISTg79
m4E9tqwvwv/mov8JgVCxtT9N7R6mYWTo9DIbreenxaJDf5ZuBmtJGSlmDavZr7Hy
mkwXuwUJAZI5xyspgWYkXHijjKq/EPqjRcPD24NrqbPDW16imDMnjIWRRTSM1kBq
z/snOpSv0MbjV6mku06DfM1advPT5BqvRkllvw5B3k1LH5CXxOep7LoKrrr0QsOS
q2Qrna68UK+fmxJzjq5kaQbhNFEe4JE2x6ixc5uYRV6tlmlJ7TjUirOs6KQcpD8Y
805sRSVrOd0KB2quTjLkTwrHluv0jfbQVs3vDWDuMrsiu3BrkNniaGlhaIasQw2z
TQlZ+IgKyUnphH2775HOh81LM61WAg6/vgmvo8Tc0A+6XDm/6pf2rBGJl/Mtw7yv
VsVDCypteeCvXWWg5TtEaRowzgz4OEi52RUMrS3nKZDnk/Luug8trzoqbP28w51U
FxrrwRV2zeAv1lmkbc5Xp5f057sBAwBQZ883JCGEbUkNqMvZFl2k7J/PubN1Wb3D
OxLVgL/BfoYIZi6ik7fsEiQnMGRqU1U9iugezJc7Dbg7zpadcXgKPw2sUtj5LC8o
Q5M0ow3F52zpulcNVm8MegOxOPSg5R4DRWeX7rfm+EaRX5OLPJswg2lpXL0TQ/B3
AymCtximqYW4SA3JULQXI0Dg42+hM4UNRAwmefJi+Bd2XDV1XxfnU41XfGCMDNU7
8lnHUmlpxXQeZCf55YUU6bj/dMhdbWQB/07wwZOMLd1A5wOm3gr+4618xGQaxjmr
pnIkc+9lua8Q6/9TdFYp0g0qZe9XR8X2C8uvxXoQl+SpBwXbL5uu1nQPHhp/futV
AQQcW9z0k28BpH5Hw3DX44ylDbwDUHIS0BiLj9kZPd3eGEvIpuqADfQhwJaRDiuL
v4cncR9Aa5kiVu6pZIuTCshYfw6yRraicO2qlHQEknw6+U7gkZawZgiIGBskwox7
Vg6yNdBXRVmN2aEa30cjqmxg9qQWWvk3lHsSu2MypVFNlOaDAW0sHgXGn4Ab8VMO
F4SiAaH58JPXVvOfNLF4fN1HdDj12BYNIEEWiDGoc1X1zuxaUCGa0yLjPEBHCsCI
OV4WU6TEffJWBdLVbuOfZpVt/kp9wisc8+l/rXw6vQSZTIq0LKlKP74Jr0ZgkWu8
fGbUzf9fNg9+1TIupUwvvldr4Wvo9KFxGsbX9rU0zUPbp1AVzNzpsU019X1fYO1i
DO7BmcxdEEs4tsAE5PBhOkcArFYRftGqtayo0DlEoqCoGvFqArOw7fqNGIWghVfo
DIVKy/OKoIf3lq8EX3d9Bxj0dpbHNw/CjA/F9ph1dLxvslNfG28tTREzqWm2dPrZ
RcO7LM1bM48TQ8oDJ8JvaFi36KI52lyB3nD60heERZJnmbvnG3XI7KNB2fffAVGX
Iw1VDbGVfBZlGrcXDWS2aAq9AtMhlV0LN8qP5XdU+Nz+AM21uBpr58sQjo4aGuna
q3FF6wmUBLaWVoqGuYgTK2MKQQlrhMV+iunSLyhcv7CA0v3zFMBQiRvP7VgNdS5l
60ZsGXjwhaN3iSjPcYL7j38Denx0LJRaRaDiCnH310ZJ3UWwxOgtVkDTqxnbDr+x
Dm62lRp/dGFGhz3YyZuK5M4LJriFR66v8wuC12+V6hvn/maZjKwYouxoxtCy36FJ
disji2g2EH8DUG7b+HYw9yp/KC4Ih7IzWCs7UWqq8oswLoLGZLueT3jIE6zxAqPF
4Z9hO907NCnaq1oXHJuyk07l0x1/aiCR8eOJ6445791ynovyvWr/km9WJjX70HKV
fnEWLPfd1FhPlT1BaDar5nWfWQEddFUbkwiGGmnRVbHaIgNPho7vsGi5UKHy80X7
FUxKoZjAatpmoeWURPZn76xgver3XQDOBbgMuQ4bLxYb5GIMdmaZB5yhSD44mbWP
l79KSbq1v33cDrddEf5oN1YoqDyIsnJnweuPqirKb0G0MyrqWS+ekFGXSz+6laNz
ou52RbzftD6gM5nee4JUcWCoVwhhYY6W0GK1VeWdggheKe8ZwLIHfKLF55HnhA7u
2X1vduXCSV6wWVmBEiPY4usslUZT0TAxZxVWsBFKEkgYknHVDnOGVli7qdDI6iUT
XxD0QkKBqyb/6j0ImdhjzCBiY3KqEl1hUd8WTvmfNKKIcr70rSvUJMRGJB5hGahj
zFEy5uC/AaBRHUnsfm5xS2fKM50PoYe3GeOFOMOLlnpHuBaDzJSWoIlsRlAvda8b
ZsOZ/ZGymr5QCCJM2B0kFC7SBqhqn2hNcEEwH0nutJ50nftgcLojsR/Wspiyob33
PnMoTsM56QxLoAXWu+egv6P6OJnY7sm2KpukXokcN20Zc7M6YfR1KUuTLLXNBU7X
Q9oRzzQ0X4vCmXW3a5m7I6Zfci4ciP2ywFVxsL0eMAQSQJLW7Z8B5FvMcaQrPD/D
NBxKDHaJ9THJqNiCUK27KbqwvOHiTJQKh6s4y17eeTNxVEoSfFJ46x/Uy9m3uSwm
15ePLE19l9XW47fmIcXH8VCpn2f4s+hysQCir75dZIm8rJ7jNMq/UKq44vJJmDuD
MyCejOItuLD4wNqiCK6s8tfLg1p/fK5Ws7+Q9/Z2ZOXdJYr5mzEjfnD3NTpzeBdE
RfHyqUhgai67ABjfW4auK6Ug4cXVFQjkCk8YJnnHAG8zAQNkeo1uvN3l62m3VdOy
RtBKHt1XJf3XxtCl8LWWg+OhfZRHIXg+JNHiQwivWQQ0W2J+Tr7SV0ozCYF0mTEj
a2I8iF1/YK2cwnashZvbx0Da8iUp5aJEQLGwNVi2Ex5hbK5Lw2P1fIDH5qr0Sji5
L+h9Io8EppPKT7jLu9huYLljiOP/qcoI6Uv9789fImqNL2oxdHinY7EbGnojA5dR
CPI9LlPt80jO+IR7zaTuPtGdeEOcTqFXWdjSkHyLvYmZI2OJJfGCY83Hmz6kp/j1
fuciFR+3KF2hWUQIJzaYrDWvUjcWy6UxJSRbmw9XArr0ZKB0Te7jDAXTK5qwGLDz
ECPNADiTsQe0TRtHa/g8VoquhiDvSG+AYI6RYq6p1U+O/OTuTAvlO312Rr/ADqNe
sTED/cj+NwSlBt/zRcGvIvtsoO7m90cL3IsKQQnlXNuX9pf1404SyamPqpFOA0gf
yH4NsNROr9jxiJc30eNuRAcTs4TQStA5u/CHOMShLS76NsAzoryo37orQhGZzID/
tLjgw/o2zECVgDMwVKSq8TkoSka1MHr2C3wxzp11JtGdHIUky8GaM6qkkBhjFcIH
JUBtrZc/TQDOSHetW22g8OB3ApdBhgvEWyvWKWgdHjHW6iOihEPIJkhYfcal5ge9
ZlCYEgMsEBYVefu2PLFwf2YEV/wwhi8NZrg9WRNoPRAQP6mxnJ/9BqH/zFc7YIsR
J2TdDQ/gP6nuTEOkPtj6B0TSReEUqGaXdMVLu/yPPtoO9JfRrXICBBOHmCkG45h1
OjEWrTRf6nH+EaNGwRs0bxqFUkznW97BiDyv0Nier+xE4wG36r1Iurhy18FSXfGZ
R2o5tz43ZWVasKXskFNmM5RrM2H1O1w9mlxOzGQiALjyWtA4VibsPOviEdTu82aX
jUe+QOseH/LyOFmEdRTmC/UyKlgoNHIDDe+P4o4qeP3L3DIfUjPsVYei/z2+JJvn
M9NFJEY6MEU2wXHJd5ac2UmVYGa+p+UWVHdEoZNDgagN9DAqmC21fsvh7tjGCkkI
B8CYnXk28KxxigRLArWio3FG4sKjv1DwTqjCwbpcO7MfHFR/r1FfQOTrV7BrbOTG
4DU1qmTkau3sUhFb/63mzsrTQoM//SbUtHv1Yz9oMM1PYwTn5hE7hMSiqx20UPOs
xVRUEnXNnnyIZRt2bg1+f2r3zYgkj0s9ySUoAuitn5+tob+xne/7fill84/uG0lD
r0m3Ua+/JMujszPcOlkDmQCMPAD0DcXlM9BgeMD7keAAWf8MfPHLQq02lD2avIAj
1OAw68tgCQEQQqImarFaY1oN2JWPUQxHDXffiImpF3XTwUWSvW6BPZu0TKMI2yMq
cI0Tqm+8+VHgQXbIzczKGKaCZuP+pomfs/XvvvGNJBe6HiaPoigEQLVrfnxfxqBe
U4yNi8l5PzkD7ANF4JtzkM67QBMrLmNm5GHEb7Bs9Bfha31snFFPBoBoE7SuQEOc
ALy7cwTzDkeBD5YlEhU92edg3Sa0GErf2ottKeTH8dcg0Qq+fQiQTNRjYzNzw0ds
B1S21dsgfkhTbuQFpDCwAY2oILMLSw4scf98wNQqyeUcFWs+DHZGEUCcfwqyWklG
1nYllsyKdukj5TUpUKT/O5xkSGAqShwa2WASgNIrGo32fCAzR8tiy8QU7uWnIZrS
/fdOmD7zlKCp3/OA+JqAyYQzciXL0aHhFVqBLOtyFsQdKLIcO+jzilw0acnZvl+u
gBlh54BqfQn6QEVa0ZeYM5ljWvTYWRoAsCYxR7qBgK4wANnQiDeNmalKuMVKsNB/
1jTwVQkLhmFDbxkmI7b+MP/RudhC6xkB7KcahRehFB9h+SF5SNIvq2lUfPvYAip0
M1Z/qFYjPCX/CgBw96DV2AS5THMzkRITvJjBGHIXgguTkW91dKuLfEhVRk/uUglR
F3T0Y1ueh1pYJcApUq6t8rZ/y9EBTbdrDfNeR3+rw2J4L4vzzWtsgNOwk7rls70g
zYWiCmkEIyt/Wu/xO9JQchdt7Fb+bA//vQV7sOTscZY8KoxrVzV2JWkwSb5bTs4M
8lvMe01SgaHrpJWvXOLIXtNmYSrxKn4s3EKtbh/JYiWKsixPVYmk8tp+7pz2jSGs
elyObCZpNgwyhD59n1z1m8w5PnE/nFnDvVgLBkL/6DAj7dCx3zDPaPMJGyZSUztV
ysC2Cgst9OwOMoDDOCXwYqrr+YtVQCnUxnLQJT4SUBcYRzNtvktDN9XJ5Kt1k3ic
DeRuZKiU1lEmbotMgXiFBB9JZtfp0yG1J0dHUf2ca5dpRz8+WlriCw7ybYNUzjti
1F4X5N/z7XRC84uSGsLqTw8nUJzZUlBUKxAoC704cxuhbGJ4FZGjOe0/DGRxNcHG
m0Ai/ONpvNtVXyXufrLQlBxHUr119qpwkEcP4Q25zpkXCERJQTQtabRHOtkG4wi6
oBogbkf2XEs0PUznNAqIiJPnKASvOY5esONfdwLVobNgiC0o1n4taDHFmWb32IIc
H/u39hlggeVjf12BREHGrbzMcK0dDL6uHfB0sJ03LcD7pJPA6rfpb2EY6PdmgnL+
B2UBKiMwp6wdW3uwPyz+T1pbp+mEqlya4r5G9Px2ESDztwA2pmiNwcYtqRmihR0p
do3y4ofPdDP2UATtOt6h1tebJyBJ463Lf/t3OBKCTXcoYeHBJhZnuCqjvLlZQbWg
XSFPtEkMXSAm5l28k7slNnwri6VIjdBk9qAfWsKhRD+FXVxKjRqgPelQ6n54+JbG
iaWhfQwohLOS58WndlmmVo4cEApmCD4ISOy0oD1K2zKenUv+SpYtMrPopmyB5Fh5
8ckSBR23HmPdUOAdfebTu1Qii7vX9Ei/qr4m6tGkxdPy78BAwzw45RSFmXRhJwTL
+JcsYWeB+0SIsR+3R7wPgKypXl/MdrG7yhNAS/sxS4mA4YOGem+p0B9sXrpUmhJX
Jeb9ygfY2lAmjGmzh67NOrDxtJDLv4So6d3V4vnFSbE3El7X0pcLzoALp7BUudQ6
bMozoIWcx/yUPMsJe6DZJHW4b8waL5lcj+TZIXgUYU24i5aO2i0vmGnwTz3cvnC0
K64CSh/YAmJJMBZakuQFzBPQFn5AIpgLS8y6pQztLYg9YPbax7/57mvSr7K6Lye2
a/rPP0gMu2TxOAtFC9PwGfJue+OQkDF20BpL3ppUDnefjhRxiLeebc/oNLDZMCdn
OBi/VTroB3LqB/4crZ+qUXsb5YYgQsUgdwjwVm6tcs97LtZ0ujIEaCWAgNNVoXOi
+XZTGn9IqMITQUCKOwrUycyjHrVHTFfsK3OE6L0zqnitJRk3PyEs6VOA6Kzk58wt
1nn4gw16C6LqclqCSEmMSvYt6BZ+xmpWGiAfYGpa+P8hX9fyDf0cxJ2EUFcBvSn9
iNJ8M0x1fxlbBAaLuepHu769v4W90lv5pe0SttmWTPWbJv2EMWHmYG2eKchO03K0
M4yXTNn/Evdp8e688xogiZbDjPzG55B2N0iEsvWx4T1xXa2dfVULh4rCWEOePI6R
+QTKJSD3uYQMBiwbxH/7LINd8V/0j6MrvCUpwWa1c4IHlzqvWy/zwYBN+OiJ1yq6
wN6f80yUoDyriq7+n8LUjHZzVC0bZlvHrvLLsvDVXGhWHyZ1cycU0fsxYwJKsyVP
S2lI8HGJ5HkIfSMLTzDsLy7Hau1jj05M4vbUYetNIqtgZKbD3R0Bm4S5esGK5Hr2
AJ4idDK5Y33SvjWPO3ICxJs93lQBKzyBmhRd2SXjBAZjgrDvX7g9AWUrNB+umIdf
oOJuHt9j3nVPLp49lr/6MVGSaoluo41KSod5do8YXhuadb7jmQQvKSO0IPMYHWrg
JdPaab1iIBesCNhTcpwDDt4F/84OTsfc8V7PECbVBprGig8Q1lh+LlNro9/sGdC6
xpw1YSawq4SxmYj9+U/LtWtbOVrT5CVeOZbYg+C7W384eknXXRh6zc4gaOzNEME/
KG+ElhiPa57/4uz+kl4g9IAKiivXWtO/GH14ObSsHRolU3KbX+izjB67d+rx9J9+
RzDDl4Dy9FWpzCIY+cnzbb79Ybf8D7E5K9ZzBnly87dqJ1wM0cP1VF2QPw2r6UCu
B0HlS4oMbOvhTI2QIwOQDQtN7imzoIxaTeNkXl5n0JoourhjZmKvRoeTahkKwbWe
5YSDHadlsjYMr+EqkfXjoxpQNEhQmm9wgQttI9L0LY31xvSa3Ihn3FZoVpPvcXbJ
USORzM/hxXxL2Oo6DNS5OiFWPanfDcOId5juJgNXM1oUhSib3uNLIMq1m6e2ymTx
4fTQP1h2y4sE3WGbr+9D1whZU5FbwvTQT6wZMlhShhYjRPH5rZzT9hg7nxqVoAPf
bjvppiLnAQIC4fhmAXgAgCiPid0SOqtNj08jnIa3XfC0Bq9RCyd2Jw32tGb1dEWi
yUublTte+wZ+hMIOqAjYawQBFWTfMwbshYWMeaS3gV+Nv81g3VtdKDjVZobwsB+i
+lJxU89h6B2ZXKCUb+YhqcuC0JE2cUaKyooOwJHp+HURxN6xfJlUYKgI1BpOzJ+J
dvSIUv37jlXLwt/SaVPSHY9uYMFifAUPK/oYYgPgHZ4wtzwHGV7Xo/cbHShXtXSP
98OgYj6IiG5RlEFHoXGNuCR+daq3lE6sdLrGbq4bqIeJWtzjZdMCfAeB1hly8bUa
1CcFdVnXbKiyC8iKLTNSTDr2JN1gmmKfwtVdGS+t1dsONd9jDfWIsuChwXJngkdO
9+NYW1WkQYl36zyY6bwyBQx0HgM4peU3mUdbjS0P7icOyiuqgzRJL0pQnGygcWv4
BeeHHDk+IU1qs6uxx/SVsyhrCOpaOe8fZShcoLi6nigtDN3Jh8+ZXW4I0JpHZXzc
I8iWeVfBFSenVT214HPU6ltgGTRjOTm8IMx0d7U3HGpABlOAkZ4SIBCOorOUZPe6
ukP9JA5Ps8aq96AiLrlhY5D/MS2golpUB5wAezn0ik3L83j1Ll5iuVXiCPQh+CQ3
BPVnoVce4cSwzQtja4z2SSEwrrTTWd9PvQMY0u3vc18kcZJ2PsihfAOWWHTIpL9h
N6BTJqPqXythBmplx4A8bmF3cfN7J5jq/6OlX7EguZP8EG/C5o9sy3qel6p7rn9/
Mu2SIMjjfyGaqkzm2QWHdJR45wBt3v+Rv8JqOUrfaHt6aBKyKBI3ehqID2t3Ndof
GYLhLQdZpvqGKtVIwO6cKCpokBQliNaP6YST6IauRs14jEMgy925EqpVJAJaxWeK
FAptYdC6RnXTwpUHjSRyyc9V8trX8r34qESz5nNnTTY+WLJcjGShvFdaLidStZbl
52jRezpYBlUIaMyzFmWxko7ksHB7sTYcOFcdhHTvzVnX1oUfMUEyHV3uMJTGbUIb
6Pa0pQpj+418WnUzZEDCe6Sj59TgyChBdJAv6YLLHeAgwZKL/umWiFMwOSvUi9JS
upPlqAF76osGk0YYIT0TvhQ5bomM0Xo/nuFTjjebxx2Q5BbtRBXPInZV5u4AVdGX
gRpzvWwy41TOYpPfCNUG2NOJSZEYEdndMmdJbKJxtvkz4To6VOCpNK/njO70aFA/
XYKdufySe9MP4m++pqIV8gJxvnQFVu0btYRdvaCIsJewH8D9DaF2lFY09Zc5gQaN
sGSLQrnNNTgaTVx+SGlfYSO4mXvdSWqY9beRFlx6U3mxNdO1yd+mp0/QfcchZ0SK
XhNhkOp/bt+nquYlxOR1QkxyoDIk+FrrGgX5KtNpujXA9r0RXnaxahHtWd9TQObi
8+vwv9qo19DvUqQ/3pG1h7vTW6iWIOjouVaL75xGisXwi9Nv+DqfGs0oq0jHlw5q
KSQycgZ7NOKDfEoYaOFildkOUUPrwHNyRgCYyK/ECHnbe4FMvIFQ45jRqCkHlcze
eRaeY/7ZGz1LJnx0ytbFdtlxbyqAcrtAKW9F8QR36b45zjkcVWDvQkRrOJK8FgeP
U4/+Hb5p/I6gnC3utMjNkBhXgL4L6Y4JbJ9eBFqF/4CcAkm5lIQYTn2TnD5ynhjk
MoSDtHOOfB0WBHwAod8VJnfJLaUF6ADQXITc2IXHd5MmVNbWJMfjrQsfOU1vCexC
XeYNz8jVLtNZX+9TAwKpba3PN2P/FJIk0H7O4Y2aw10uKikSEdGvI1Gsgh5P7CFS
klEAX77wjGz/NUaj/x6+q6J6zo7jBbz8vs7EPVZRmyYVWyXZuRLnNbctFMNweKLF
PpXOZz2H9l/11QsTu8lK4btAw/lRVwLpi5Zd7tpljas4L+QkA42KKePHdq6stGYN
XZ1zJz+yc7f+xn1FsnoMukSqY2eY6+ObVExCBZGQKoXhpvpvzR/rSEUCXb2D4t0E
lzk4ozsvdi648aVANWs/qEUoxfNO1tR7TyFlwtY4dr+Cc8XLqNtHCI4hIxCMyx/I
VJs2Iec8FCnlr6hluiBdIgbD47biBg1J4mWwYik/23yQ9NBYJdeZKvAPxEqqiS9U
i5Ume7ZepynnK8+W5XL61GRGLOsGzAytTT8+qd0iHhHTB6287C0Jmoxe2kZ4OoOR
tf3sqmOKA+WbwGDmYx1yDGuK6l71ZqKOAAHAD3hKmdveRNvFnZDpXN8bajBeD0Et
o9bkGZ2HkwFeDe34Gvkv0M/eChRWx8s9orW2gI/YgxCEYpXcj0A20j9ilTViXIxL
5Jczpz6Cn1dnBKRl2wQRR9IoljX2A2GQy1y6cJ+0hibwRLnccsugqgNzL88Nse21
aYzq/dSsbJtB9KnqA47Ds+/tMNXeuWQpq8JXCt7Fze/n+7rpCBanRybqfvkTAK+a
OVR8/jZCJVd3MZuczOm6tBzR7sR9NpvfMRQTyZjp8jaRbldusGLF97sAeuv+VgcU
/7l+V1w59Gx8P0kHHRKyAmrDF80UdiUG6tXiP7xjPt6R2j553wod9V8UWFUk5nPf
+ndE6CirZetavj4KlwdcFmezm9SAP7KCUbLGNuFj7tteqt3V+/0f74fSDnXnqZTi
IoiEjQUZRDQ7WUb2bnEbkoU+sq4nePYL9Hy+WaqC6k0D0sdJl8oVLJtNYvkvPPoR
I0HPb+YJcQWaZDK5TC4+ocluvMjbnsCrcW3qJHaL+BzkffFllMvKzr2VNGGEjcDo
7Is90Y8XaT2ujuIYLk6qGBloAD/jCvVzfJTn0vgYtPC5CU13o3qeQ9Xkd1lU4hcB
TY1CjHcZQlN5G/lMwJ0dKsucMzJmAFJeu5lgqG4lanEDt33xv6c0dp6Byv2YD1k0
1Z8dZlRK5HK5ptTqaceXAHUKJhUNJuE7DLqpUcY1ymi0VI6ChVipmUuNhYO0Dlmq
vJmys9BSsde6GZXvNKD+LFPMsCsqPefJtVOzLoEOsZOw9ZVBoWT+TOQe6BxZt4NH
DoAL+ghJKSzUQymkw6diaQJRDODj7y6DDltH2qAaP1dUet0rvAz2a5OdfImLPH03
vn3dnCcSIB2vpPbjcdiWlAq1Kh1moY8eMCW/qBnQuhpyqI1LCe+dZ3IVrjmXyrKe
0Gc97Qf+XXxSPkPP43ABQkIqj+d+Svt66LBI9qEvjN/VVHzPXCy2sA4bD+KH5y1Q
ECPF6IbAFucQTWwWK9WEucU647zduxB48jFnoy54uRBSTWNvhfOnEsqTB0ZAkrri
KXdKBuv5cNjSk0InyBxbxub1+bM77/640MsCqfDYbt8U4bnGWp8+EgmSO9ouIkda
BNzXOxRABhBi2rkXlhqk7xZF3YHNtYoI9x2V8S8mB5iN9PtXUX9Tz4ozbtkbyPci
dwpuh5m03cdfomyEdsMNKXN3w2SuT/Hso7lAjLR500v2/MVtAUNFjWh5EM6CLAZR
l0Zz6F0lngH48sdyLxQ2mXiIqnncE4XAewoElB9GFfvxBsF3EAxl6/DKMeV3lamF
FHsuLtgywz21icFrSn6CB9SH3e0qEjF5YeocbHRkSTsOlvb8PMtaETf6H1Z99RmR
oLgkd7//a9vZ0PC0HCmHr8nDJ9SOdp62oRzEnC3fjZzW70LglkbYwJ7EQKKZIdGH
cGdzCxsQZ4uCHLrWPV3aGEsD3cW5JVNc4bL79QssKvUamZdBziP268lxf8TegHK7
8w9fuDBIFbm4h0pTO4/on5MJTtC1sv28+916bB3hitRvZ1hRYqqdXSWFQcqSvo7r
0Yssvtr1HiK/mZTiyL/F+OFi1TKVJnPeIw5vTGo1PBfYMrEVDZrTK3PIfj64KzsA
Z7lhQSEFEH/QvmscpEZHwFPSQccmskBgFBgsXzgEVO9/DpmAisMlPiz/OUCF5fZR
iEAsDxVKJZ9TGgPvLnciOV2xsSB7fx7ectwdT4DWWRqkbz4ouGtV4V7aRtlBuc89
RPkUskNc/PEBklSQnk3WW94hEqIaR9Vsq5PLewb+1CBBl6om9qbkbXUEnGUzeq1V
LX8cjkYaG5IsHFvMyjx5t3xoHOOOmVs89YqlwRIKGt2Kfitxek1cdSenxOWV9Azj
jyzXYgHZa5oxEVMEHsDVXttEw37Y1WTpN4JiqLPgDe3p2znZib15ULQPMpW5/PYJ
8hWixFAfwOin6D6uqXzIF3VjO6KCA0IPrvuUQgfhgh+kMfhUYCm8XX1DhcGnMBnj
rXRlSishdPZGsxrVM0iNLAeBLobpfGi09kVGLPrmXSt32qwvk4138HR0XN+Au3jJ
9c13vSuCteQb3VG7uByJlhtvU8K7V59SwtzY1gD+GlQGygfskFzI1Y1kmpR1laCL
DXYvJx4KZPteHowR9fQLGAK5ZZ8lX37ftACPw8ufqgAs/BB59bW7iR+U1cGfrPNQ
4vf+ESOW+bb3ukafM04FB71mCJvRL2hI3Mfc49f1biN022g6+bFpG/zsM3iYi5AC
XumxjK0JbUDctjo28/WjRGHQ28/qUVrm+GEia4LkdjHNzwvrSVSsDkhnmde7pEFZ
fVoiskTk4xGqZjojKmZWn2gK+sanTnuraWmLqk1Xu5toJ6MV8X7qYS52fG8XiJES
WWAAHf7O780kNYE1WARBlIlu8W82Mh/AWuTvLxey9EOr/xoAl/rNhv8+YFX2qODg
zhw/tdqN87EcjogFm4Itq+TsMWwKbAeVI0wrbGiRFjUOEKe5K6bLOxzukbR5BER5
F75LdO8yhDKhYKcYn8zTYhQudKOwGCNurcoVD0T9+Ysp1ICgK6kHTZiSPk1j4IA6
shHz3A+pbp61cqC8WSZ2nt/iljywtGOjroNsNcM+YQzCUOclEvGXngrp3Z2U4rPb
CW2gwL/gp/Gf+e3dil7vs3c0wX5vncRBH5ZPwQ0DvyCdrMV3T5eUSHy3l7fmgW2A
j9LHWDL5qOFPkokSSjKlvR+BBo1E0H597gk7ls9Bbum9lILQ5PZ+RU5qVUFJzevt
iY8dnD9M4TU8SVtC3zUF8SNsS6Yhi1H2iVmkaNq+VF50+j7ZZRVzQuBfrHLD5khY
qNbPynVc8WeYBZEBffFe44ukpTuSCotMSvqZAW+HC223a4mYbtgJDkyJrmdKyGWo
NUtOEgKRZ9BhNfTY53O5KCLVw2oTtfMp0XYypGsKmdQHrRNNwrHf16StVzSNs6xE
YvFujS8T7dM9LUXNLqUBV+W8ewbx99kyTfeguKrf1HxH90o7CCq6/Kd+wS/7rOsy
q1BOjAdmFxUx+xveu342QcHMmNIjFymJ0VZ5vPQYd25UWAOfilwhtxZLAkQpxAVL
nzXlG2P1YaTk+8dE7c3SqNlMi5P0ud5vSBRxMRDDRQdK73oed1fEB+fVbU/z4In5
7hqlPfUUiw+gmkrSp6AyXE/07qrBbmHLY07FGFlFqHupTNTa4NZyYBZfDWZC1Q1h
J3DLZEch3PpZvKpuLvqu/zxVxrTEqL894LjndisXPjulmW0WoRR1m711dbFXF1eg
vg0Pj0k5iRIEJM+epvFbmX/hxO9F+w89t8IAWdASPOIwo88IyYfy5Gwsd+HjEj7D
Ny8NWYeiVXDzX6f0OFJhdjuhYS0Se9AxaFQmucbOWjfExNZ/hm/efhedX0SUNePc
ToxhX134ucb0A4BUDQzWU4z5k7/ynaTDJic1tJDfdgGL9rEAJTWOAL57bxkUvlA2
RYsruxdu3FcyawaxcOrWzgah5yeP96SCEivjHbDMDojLo3WnLDifnEY7/VBNq49X
tlIOo2XjzN8C1QipO+zKXiTWbvH/U49eNHOkW7cNFdI3ba0+h8J4HJeXhrJJXYvt
1NFVstnowmoupZf40/zQJR+2Z6Pf5my4TaQPjuKsAPMv/hyuY4JYmgeCz47zcGcM
alEk2Y096hm7cULfHHACMiI5BeHSikxK9AzNT/beBRGUpuHXyXqZf+7WNVhQEMwU
w+CxKqtD7IlCxg0yCLpqmsDGIcXJxe0ej1E6aX+Zfl7pOEgXwNCZF/U8sMrpB5PN
uyGxcleLGMtnJzU1H8Q9gCnJo2yES6kHqJDfACY1BhhtAIDP4xX78bLWwwRn/XwG
mwgOi5Fs/1qMt9azkwk4/GpLTHcHb37vKV7uboLgxPDW4sdaVGzItr34JY0jvkki
iSlSAeJYFIEaDndlSzPgDKKMOmPTZ5kUBN0yOVMQHlj2TFaHy8XEzCOtn3PHMZt1
1onyOK0tzhDxIQm0lO3h/ftyYOkDhEM1WRFrK0GVj4lfE9PGGiaoxdQEtbaSS1Zj
msct5WwOPTG4JJin13BZD6PBIEY4Uqz2b0/molHEHM/YRR/Mpj4EhfW2l6eBrKKj
4EsviTKeoRNDo/XFHz6yxgDp3LPxmBl0x/cmJwqTNxa0/KFQ6wQ6lLRdbe0z3HU3
84M1biW+BrcIozg54frqWPZ6xFgv3YPKmLtXC7vecsBJ06eebR6NFUs2r73qR+H1
xglaLxhlep3sUNxbgGIHtyM1n1upW4XsObmFpXEP+q6mHkRuE1+GpdkoTDQLRwWh
ye6Ugm6saaLv2nWort4RDdlF4H6fBJhezCs5kM6/Ba6lQcYyFodAwFvypbF8ujzm
BKneccAc4mIwGt88bIvZm/267MwevHffI66yPs8ER8/j2BEf/Nc3NtN1xD+EUNG1
uiEQFx5EYosF6TfXNmTHeoioOsVS/5q19G65qM6+jVzqIbHyvWK5EfzRtCB9W1dr
N15R/a1yBZQjIUCqZRHdXopTVkw+dD4KrbHqEx5eYzxOHvRq8ZjZjmCskerWj4UV
mNreJckQ/upuTczEX6zxkWDLB/ceadlZ9RQkZkhbXnjhOK4PLXnNn0C8v6L+IIhf
3I0LDy62muMfIkV+2sHUdr3YzklOStjV8L6odJ9EQ5fMQ4s8fHQ2Z9awqnnlAho8
fLWAD2YHLgocwWfYIoTx+thlJnJb+5lv3slqZPND6YCNgAt9PNvOKnhf36pDtMLx
Eefuo2xc2+wU7SvWC28pFBKYiKidOxU7RFQ8gKjNajsFtkhL7ST7MnzzLVZhcp6f
sYuVbjNJDb4dzexPTdEQNYt468KSYvO9Vb6gsHOLm77i5lSfVnmqu/+j8zGb/Yn+
nufaYlLgVrQeBacKovJZm6m7yRuco44UsIfHzfMe2lbS5HvIFnqS+94s4HuHsIQK
tOeqKvto+9U2yCfriS1ScxtRdSIM78w0mvTtBdI3igMse3uTJR6G+DVUbo8JJSQ+
CpvuSJI4fYiLBeOuUt4o9306i/pPxIJnGR5jZlF4yVkCGVT5ItqHPHxyG2IUSXbR
JMTd/DCPI4Owgm3CALqUfp6SZRrw3H/mF7GS/KIe9nteC2l7NqQDZHUHbjAyvEVT
opQNqr4kmBko/DYuptoY2ok2YeAOIe77bBWqiZjI47L/JbI0r1L7FuROhD6nY0x0
jDM4NZuuUfTx7VD6b747YbJo/3/jS+DHyUL+2Jahc0ugC3zfHjht6K608a+uBPjO
7yzsDpzpLhWZUs/hQ7ClrXPVfnsyXAGgjKinbbzX662PKiLYmYNNiyLyBo04Z/AL
Kc8H2pCpJJrSU1cCofMPKAiTIH8CK+4TCHg4i6H+v2zyE9722jzv6ipLeH+XHaE1
2Fkewhxu6NYi8yObSsRQW4Lp8qfrgulwA4XkEM5nlL8VwMVV2fteO7AJMZJJls58
JW4gG6wIkTvVIDpNZpCjD6pJ2d3igpvsnlWMhSIUDX0QRXu/+woHxkzJu4Kd+Y3T
dW/L9i/xzG9DBKKhx5wP5Q1re5VRzI/v15GNP/OIwm5NN7m6MXLQlwlkY3oVJeAk
Y96xMrnU37ba6hgnmB5mFwGxN5iX7wPOSrzYM8FaZ2nI4xr65WaO/8yHBAYUDpEM
St8VPBt8XBdERFLNs1fPBc8v4lQAMzzjjsqBnMQjEk6Ct/sk7lJVvO2miAEzrOHA
Mfki2PpyNBKGS8ibol1DKuvr8KrLCid42JzDQov8HJwA5GxaPLUiXSpEXPINE6/z
voNgsBrOxpN/t0k06e3fhN4317thFHGNCtrkFvBWwlL8KKs/GEpP8X/CtDwwkUgT
3RdtBaYlG7zCVfizqN9yu62OG7rJ2do93kAqNKBRyZWqS0j23OwZ7GaQ+z1QMZzw
zqHEAsFRQwNJxzAVqGtf7E4SunWe5562Z01eNE8vIAfn4Vn75NDb63T6VtGpMSL7
AvSI1DhTS1Ny3d90dOgDi8IalVR2ATSSivvwavFoXDt177HrKN/DaaL2KOLDEktM
ZBCND7kMJQATjsSBvgNTn/L8taU5UK53z5BZpN86L2Dr/rwd9XtWa7MTz85dUG9X
UNUs6sJcPtZibeKUaPNLlIli2Fmxy2FHo0MBzWl2cSp6m3jASYr6JX3ORpAC+3mg
FhvnD/SioWNA0rDcGJtUM5KZIwna1MurUsAInzh9pRs9xPzJgk2xJfa+3R92ffYo
nI6gc5IwPKlZQtYw8oygELc1tU+Oc5//yHZw4/PnIZ4oeKX8zy9UghHzbV2cKpua
x7nz5aqvt2CwH/dEETKZmXCVOJykJiJD65pAB9F5nBtT+jd0tEfILVecvEXXBhCi
AXDOZBHHhPh00dkpDfJgNZVUVj6+8ir3v9yNSDfbsMCL7nEfh9Yavuakk3gJRNCK
ba5K761PU48/Jhl10Ui+0yhUuQfPlym7Su0yXMiiSfkFogBz8PhkFR7UGpkkeeZZ
dbGKysPDfEgB2pahD1puxKdq+SG40ml2XFqs0KNzbGmdh1EGex8OvAG188DsdBtP
eqTWzk7AeSNxACPDVo40HhgZZo54iQKNrqapLc0ZIXrck/bs8XNwY7wgBurJEBEf
2Wy50n2daILep725ZsIeQzQjcCNSSjH05MIMhSUHfVhiRuje54OmTmj9z6lRBQH2
1mmkSU/1RV4wSjdtwxYqmkQBOJnkSzoqUreJNSrfwEV39iWCTn4c9Vu7lVdJVRL0
i7drGNCIvLQjhXg1J292Kgr084PVcx8qQ0bqvyUBvu18QuU7QEv59Ma58C0XMkKL
PXVeKkOmeF5oGEH9njq1zSHMMjgwBBE3EL3Dshpd9aUy3jXOZ7IOxRDb5ddyMlGm
eenmdS8h/7ZjqhXIbV0l9m/NKi4tftH6r18A47JW/TQR/3yrqw25RE450wlQRmYM
gVqCu420QE0+Vy81w1qeDcaswDp1Mx/JTjs83qgEK/1GaMFL9tEbi+mT0XHTly7V
12mz/yiHtT0ETBveJbp/LvOLpp1Tkh1CrtF+GQPFVWpGIMzPmUdKYD9miECYTLVN
Qki9Wo5Z2U0s/s3SprUDCO3UesNl4TzT2VovLQggTHtTFBF0Pd6QSTuptrm2Dacl
xBGcHEbhesW1uyfK5LekrKSZtKkoTxQKLbKS68LVSHQ9utmdbyEbhTvNB5EZqR6A
GM6xFBAFPc3lU1DOis7yqosqb13l6aptsvldQlbSh9quC5xOrdz9nof8OmeltnaG
nPWyU5nsov/TQnhjyt6GVQ7oIuJNl7sG9LMase6Hwoj/uGGco5MwEi0lQVbQhMsx
f6TVHTJ8JPwo4Cxfc6Uei4VVPapYhrrHjjLscwv3Fe4vpH8cliewtDZoJGhPpYqt
E1MzXewASHSOMYvlZuPyj5Z+pJEku+Loq9QUhIy0dyb8sRQIWu2nii4cn8nhYwnv
2ftXboEV4dyeJSg1z79u2i/HePQQelvM2hezkZ4VfI7BUyqwkbyynYi3pfSf5YAP
PknlVQwYcjhNPcAvE0L2eC3HvilSGb4SA4fAW7bI7H/HxzteqqknDFREzFtXe6de
klgpdGLd3nNGjqzTjcxL0fQ7nG8iIGJU0f5VQ30UBSrgPpx596GvzCxCbEr8oeQm
jgF7b9JijyuHSBlFjnBPw/1+Axmr7Xo+cqQf4dspujiyKeCcVJSIpVZ2QhWLbmP4
0tl0PD618Fh7QnoqObZBUMB4SLT8ih54oIIotClH3uaZ/vhzQpkn0ESRguCtepx2
3vV5+BSUVoh9oVl5+oqCXNuzTwfhk4n8Ho5qFu31UUjLSgSxTMuMBEb7/emUoOYF
f9Q+BtUIuU9XxfRmGcICEBeg9GpvST95KpE/Via2A3KOpg7A0Gm5x42u0eyWZoqX
yR4teGIk0vZnOCy9RSs7LHQP4+0Z3q2ryCMk7xdd7b7/6VPF8qDALP8nMg/8gRbp
fjIHbqHchKXcoa3ULoED6pJOKBe3aVY5CQuykqAeLMz0pi1+Ed9ppmNLpzBKCH/B
9Whj9Q6NTi6SeevlvXckjdjSPDaRym5MbrjZ+8zXeh1mM99zKQ1qBGFcOBV6EZOW
hGsKYUqbW80oso6TtCirh/XTksml9VtmD9MVjo2ygx/KaeOWUFkLTjLT4GsPtZi8
DtCBcHWxDg/D/b9QBY6yzjKwKxk/oic4t7TB+/mJiu3Yk28b+/dV4g6km1ZWKeZN
YERZzTDz8HptxOJCn0d+QUNpn6N13OyG3mXwCfRq/Srttg1nHFg9kd0Pmfi0MIVc
Y+3peT6TMSCxbb0TJP3MzmCr4Ns/1KsByO/nISdIuwgo7YQWi6CZ5ZA651VcyOBb
kOaoqCJu0nbDMKBDKiySfNiBHSJG4MBa4e/i/gQ0QusZRCuvl1BFGgnsMdu99A4B
XNCIm7di4icpj3TcfPOrB5HrJRbM81CNR8UA7Es8yT5BInszu38EQKvV8D02/Lj7
AsUfri13oA4t+H/PXrmuRh39qAfQEDYUmtjRfXRw8xxpdDMXc7rbwrDnHAzNgI8G
2klb//3IPKCdWV8g85f4cIw1UIOgEpFbwkCk4jkWSFr/geTC3lSJBbTO3qR0taxz
BOIUVbQgEiBBf7jM62UX9/Ih4lfjSUYyyTiL8dY3lri4g2G8ADpJVVhButqajRgS
8jwf2SgKif3ZbZ4pRJY6lrGglfDxRC2KMppApd81a937ZWS488pJlRhET5gtqJ/m
sMH+M3ZMDtUuISuZul3pfdXTyWSUe8pqPyEjwaXEgObJNzRG8LuBlN1jzewREjyH
QsQkaxUGZ9A+YkODVXNTnPExqaX8Swv1kMuZ4RrgD4Iqcyyig0f5WzJqQI5tm41g
N+Rlmu9K85/4Pf24/LULCw6+ZUlCrxJHgAG/zqFYwH1WbQ0pjCeceMa71T2d4BPq
E1mC29ZNS9R2JcHb9CDrQTfKmpj9M0C6mekzH27im+os55skk7smxrsKab+/Q3fi
czyLfadIaq60iKh3CowD5mC1MNhn7xOfVQIlT97P3whiTChwB23KLXtkX/2gYxEp
XiVhMyMZG1n5GzuXP1p0d4AQm/g5ReehEB1KQ69LjYeHUVK99xsxglMLjMyS+bAO
o4h3K3xLe/l27KTj2CDQrX/s5SgnzceHCe6v3rNr/E4j0DAGlzezjI0ciWjtLfuC
yFD28BP7egsciwXqUSy9tp7OXPDvNg8yiv/EsPg8Cuf9DXed+LS69yQRDKilkfR3
zeyzJQbFUsiO6K5Z7FWzwQmK5bKGcqqWc8vaB/Ht8YjtIcXR1D7VDZnkggJJlEan
pt4yWh8u6STfrVBQAOtoDmnNNg8ChIlhGXUKOUH366I7kjQOgCvquqn5H/3lzjqH
zvKe0IdN2jZ1a+MQzwAsuABbRrD3fg7kG1S/qednXTWNXBLUrlvdDTJulmCKNr0G
MVfn4p2pvvOdAKlqk/KXgrwAEUBAYcuhUYUywr77MweGYw56a0T9icjmboNRP8wH
h2jI56SeoaJD4PBv8CwH3i785VHRh0xOyv18wXsGwcaa0Pgdhchx/+N4FWTJUThl
VZ4Lo3esphbxoC6mW7w7dqADdKxMcYdbfoYk556pKghI4gPIAgx/QiMDcTjzM94w
wyP1kli8YvNyw3vKuwXn9/T29thNW7b02P226qkV9vggBJLN00hIEbsA95TRf6Dr
rOMl7SZNkGl8cY/QVMozPeb6QJs0D5YI2TJmlYtL5mUjRI22Us1YvSdAqEAiIIVc
kdYOzkUQZdjBCUsdt2Pr4yLRvizgDuhKa4+MxFY/EqypAwBvkZFD2d8LZ5WbHOfm
pNwas2/E9r2l5cX0Ntj7RcbR39B7gNoLSMj/ynkKca5zxC4B0BYbYrqgNj+iuWH1
QPlKhaBj5ZB9u8JHLyADGxx59B4pFpKY8NSjr4xBzIL5VAJhu1+CP/E4y1FlsuNy
c+UENxCmNVpgut46lORnGL93lc3ZM3tLxCau3vuJzEHiErQaLTHQe/VMypKOtffA
BnePlU2QJmK1j4ozfRG5seedH25pKIytwJN9S30X7iWX82gX84gmsXN6kbE893XM
QQ9dhWhOg31cDiJGe/6YRiXve2RJK45sqdMZd58Wv84Vcu4nzg+vHjDvbka6S8Kq
Qq+qq71ojuHLVOnHRs7gaMttwiSsWfxmb8QTlA3o6EEIOR/0ydRn9RUCpFda0ouK
bG63/1W+y9wmJVFiZwoo1Ej2TBnmNURVU68j5J+75WveBp32l3WV1cgsSg1n0D6B
Ecq82n7YCtQBCgHsA8MxdSnBiZ0i0ivP6+nh8beHEZSxYqFAX/eI77rfgf4+xRSD
cvF/dOoMmmpvNUErNFrMlNEV4XmZXAZ7JiM3hKuDVljukQt0osu3pBkyxw5kNK83
hH0qix6QEmW3RUnWzxALG7g50jKGU2kFhCkIYCxcD/0B+ecm06hCgi9awZTOEFTP
mNTI7pZn9+wwJykRwYKgA+s2FiithM9B61KDDiRW5VVdg7COcl+07zZ84dcS3MeI
7STCJmWTf5Rzveu9ToVV1AJP4jJ2dydlzf6ztXkhSOaICQjSRxmPOL7WUeQUDq6E
HwYb/F2GFduFEaQutSHLL9BRDqTrnEKgiwzP/PDiC2RcTjP32wqQMX7QzJGDBBmV
GVe3wzFr59OP/zRcRKDnBGm0PV6bAnU+a97Zw+dBiEl76yFDm5+Sjy4zlsNHyBKv
opHcb5mXuAiQX2Hwzdg83onTaTkpvB1qfZqtXjVLzI3Mp4R1qB9dVlCgjgxKQ+q0
k7ytqce+l3SlN0EbKs3IYH66O1FhgkqcYlcc4EFm01UZMLYrbueGneLLcCYmumGn
Q+qbyGhkDC6g2fD7wxtor3QeSBIuUYjxOB8rz0z5JWjZkAlpWZMr/G6fI3b21h7H
3jzyt9Au7uYZPN+NrERF6TAYgP7HHQBVwh08S2Spj/RItH35cs5rWTiuOwgVEBnB
aUJ6UO/Q9BeDfTf6GiMrzfnDDvVp6FSwkRY88kj5iPR+ygJBOD99ltOK6VFP+hHX
0UnW5DvibRkNK7XYHsNyspkez5Nih83fEnyJybIaNWh8qE5P0C/1x65nWBWwtqvl
HbBt8GZI8/VhXqO4CpmiiI5wXdYsX19AYUfZUYUd3AJ95V81uDKyLdD4xbh99a67
cIrViguAlLwobybZ/ZHDcySOgc3/4gTjsesgnbfuiqe4bjmLc6bfb06zFCdWLYg+
4GMS3ghB0tJBjTI5B4UUAtnlBMbYdBg0zym3sVoM8gA08innZYrpDOEr6+Rn9oXL
Y6ZjswiKPubYGf1wpYARpXnvsh/QO7jj1ltQRSe8Pb7NLr3yneK1t53KAUHme3wU
1axOFATTpqnLTs9KGzCjfdB5u7IIi/i0fn1GmfQ7MJRIjOlKQs2vZjlejLG2YLyX
cuUlMA+twi5tt0On5yCpoJC7H5uIHJgzvTSB+Y9QXUWBzR6hvJDMHtpUXRKaelCA
thjDe4c099mSS2rnfOyIlxr+wFX2fEAUiPo84sagWav587crtxUlXiRp3HEB8hWK
Ol4bP2sw4NdkFK5+k4EMCKtaZ7ADSeuvdSBQKGguxqdVSixlCLN2MO/R7zp1o+nr
oA+yuSFd6K/GDDszIZf1G5p6Y1l0IBj4wBaynQLDzvWissKxZVzzVy9vlU2BGfg7
d9GQg0j6egP6b0FEr6FBSyA9Ue96B1etGbkZWUqUfjDwgynj8hE04WOtO3qv9PMV
sDFIejwfDPn4xMVmZqPwZMd3XiaGrifYpb+OMK63nSbvMwe868gFNzEoIG5xnxyI
k/cqtTuMjFTg1I9Kl4pyeQF+wqcg1N5T9NiglbMEavXjFLNsb7R3hzPqi7WHGz37
ypzU4HFX9F4nTo3utocb28GzAULzwdDj8uVrPbMIpDUN6j5Ai7rWK3E8zx9j3UCk
7s/OfGzeOfxL42aM99A2wyGkViVrz09odw2VYD6vRsPijv+lqoxiY9EJ6Qj7f3aU
1Ip0CJCa+LY0mpX53PuDR7yGXdcjwtaIIFiJJmRzsKmImALb3IhrrVKooAZlmThE
veCH92U97V77aus8mJz28L5o2vMz86nVmM1USjIxPl3330dX/c0bAnCbHCZ1f/t9
Z/53SzgtES5Q5HUYy+h8Jv/idpEuqa60yTx4Ebzykmhv03+PfY9taRhFOVS8wyTR
tdLfUcF6b7VRjqQ7v6SOfDJ6/DEF7fotf4WThBwX4hlBSEPK07i8jrPH2pR7ozcr
19vwOqGs43xJ6TzNteFYQDPbnji7OsTBvIywqEbqvlLFssMBMdC8afy/i9Loe9FI
uRLQKFe5lLLt5kJ1eOZc3C+3lnPWqJWifWe6RfFYAbXZryzR92IADRCtdovImKGS
rxM+Ffj9o56IZhgAnwVT2u0kCyBf7h6hTRMP7kzdpiFmXn5q3uAWUF+Qt5rvo5oa
KOjzIqTYFU35isWs3Vm/MhTKftJymPxzBF2Dz8OEhuHz2Mt4O7uGjSN/hZjPOSqK
EsEKHkpy0p5fbZNeatbE8aITlptVLOJ5JRn8XX8ixoEq4XKayj4PIRD+k4KuIFPD
NSxaZ89ldhU6oGuzLZH9812A1Wpa3uwe46OsgQ3ddVN8Nv5QBbk/DLofj1TaMvY6
VNLT+FWEpEV6rqop+bMzqgxd3tX4oPH3bA8xoPnrpzg/ZkNNlAB6sGdAIGR0gFzE
ubueSQ/uDE+Tvu0jHX8DTOBtwIH/RJnzW+T57uH1IUF6JxxzF9z+M87MvXWf7MEO
ubu+Pae/tqGbfbIb42zoNkUr8kUyJYGS3Bpe0lWL3OPDoaYAF+goc/4iSdXOMQDo
4pUtqZ+v6P3XnTDyB3BrL0G77IEI1PXvnAJ5f1fytJdDzj6v63LO2D4dTRj09Efu
Z+rygncnxvLbDCjhdVXmu8FdpnIsNPoOq75bZ0N/EFAgGDruj11hU2/RIEcOVt1M
6zFx/IPNAknYwGcrJx7XE1FkqBiSJPo1JRqwOtLrRhHb22g2iTOCEQzXekYVFXAW
XgCD/nyc5Yu9tQrQhOKH98Mh0vXhBHrYbvuZJ1+NevIcPUzNgu714VlRcXjHsI7H
Ht9J+zFAWjuxewma292l9A5mB4F9rQRE7K7F6voofxWoJDofD3Q7o/DQQbTPFQ7q
1fh9DOEWQlFGZurixVHC4LGWAOGPBvQXGgGPaT+SMz6xu93h54x4//1OVMREmhmx
4pw8MXYx9h9d/auk/Ej4vuvYQU2WWA6RnWX3Lgn1ChMNvEOETqEzP5mwxZeHwH7k
/CxUBxiGrOyZEfYSz18SzkvaHdAN9CmwlmcvyKHO6JvvulLHlle45n+l6IRgqs0+
h58HvA7ewf9WOpXn5MfG98dwmSskrV02Izn2l4JKeIsrF8pDqb/M0FajrOKCLY1J
Xv+fXnKnKTQwhLdUyTzBsnzRXi23qYP5MKX5ocD05lQtWhQtWwj0nqVUNR6UhmGd
hdPUbpBgghpOvN5v1LS4tgNe+wgQ8E7D1L0/cjT29sUKULdJnGTdYJKnmFmQ0FhY
a5JAKLItIxPXytXfWYOl0xbrDYd+Leh88r3HImJu7K2lMAwxomqdsZiR0qZj9VOz
8XHEl56C2CWxmr5QEGwb0l2ZX2GyQMH4NCoZniZoiSwIBIxKdYMjBZJGGPTqV/2u
zNoEM/HzTiTcTARr3pTjDToGMhyJ0/KFx0jqSGnz54m+Xq4TPYMPml5zRrFkKKK6
kRdlAEHfD4xe8hpncRkEglaSPpETHm8wx72TjjwYASqpzlfKukf67wK5BTLdBu1X
CkyMxKPeRD7vxzmLCywlLnG+43H5Ji6lXioXCLlFmiVfyPBC5Ae40l0syJEVqrel
3AxIFqhVbwzIjNltmHgs7AW2/TqTE8TbIt8WwwV+6hHqgUTUHbApE+D9+kG95JkW
f596t84obuKg16g8wIz6NlSN9pitCs3FHxSJGPgu0T/nHAxi+YzPAH5Diek2rxqX
rhIj74Tv85PeMLi9QiXG5oDpUgiYZQRCL/Drc6Pnb6kQTrCqwrS8QqCHNmW6PCzp
EqEkQMwrqu24QtOYwRU/34ckiMt527iDZrKD3Oxfg4HFkuna1Qzw1NAjaaiCx3Kf
JDpVII55acHgUCFPFlX//kkzC9OXYsz5j+h4V/K/SL7c9WP/T0YDBJOeOl11bekt
hv/3aItGAfOHQ+pNRDmUAeZzn/HKk0KJ8xotOY+BtBFuU47y0O5knMdT1yIdxKAX
EZWPywvQfGTatx5H0+cr/nq5P6gor5FB764wQeseY9xbnmpEeby8Cd7dCsE7qjdE
wW/9XebAdY3xZD5tA3FdYddy3JI/mgET1zzGvjaeLO4c6QOthdhK1ksYCNbCWZWq
+x1RLGdsguB2fwDN4hO2nTcQvUNv6z37xqxx4e32ob0bYqvvYeV68KdtG1yHr/J8
Wih9+3QDmUS432m4ORWuMWBC1rzoVREkqM09dNpMjQYxk8jx2mV6gWgbu9vQSYvy
JTh1ruZNSXL1DSjbSnze5GCPrLVDU65fuGn3o0YittAlNCs2NPMAzRylFhm2HNuP
ay3K9q1ZngRXaGbgzwDQyE0RQZeBVKrApBjZ6M7p/pE3KiiVmGZimz+rNMOBEvNO
v54GtFmJQhM/oxVcmVXJNMmxfAtBqbE6nY1XNTCrW4KPtzUC6tNv6RBTUrqWP6Bd
5J/tqepYhAySTUdhqK6OrbRkkpJ2h7wAVghCWnlMRg+agU7/yWWSKnBQYpLdcRBb
7JsFQV4oAAZqWicrJ0Zer8vDAEa/DbN+rQe03XK/gGdVVKuvFFnIeAR8Q7TqygpT
4F1ZPs7VENn1SOAWXu2O88pqiNsHI/IraE+dpmdnXsR7vCN0fJ17CIQEjhEb977C
ncXr/3Fuq374QRYK7f7mGQFAGV1qGIRsBvaHCYwIcBEyOmlnG8YsmIyftoWr8iHm
sogqm9huG8jLF3jn0lPozZIdPQlkfF1rru1egEtMINqmeiqGWncLkfOfJKBLXmRj
wfIFOrOuUZzkQCHRGQQTMu/OFwwljU0rQ2OBP8DGbZ8jTc0J/j3ytRnFeUgTwkCC
EuyfoHlq9rPJX0yjoyEwhs8Z0XHl3jjo3+rqaCirbaZa16bttweatnRJ77AVf3Lt
A6vGaDXb3h4LXJc6koS0zp7w4OKR5R2sb2TCS3SkTmlFAuorjuFTCV90H4a86Vvl
ov8dP5cz2mvNVoSkqchOa8pL5l8tOiORPbLB5WEJ4hFO6sSiZJVuU09s+q7cxnfu
IWL9LvCidR1Tm6COudNUZa2QqnT8eeDPDPfTTPL2GHTOFoRMwcGWuc+7Q5f6PjBe
O60Gta0eFIpv7NjMr7Kr0J29pSy3u/1LKO4HZlMRwnzXKB6ry8CyiU142I6HgFvt
I8r6NE0vI7+iL37u1LftJSZDKXBOddoJwB8JevOUWH5U1bHHb3WzhZPt9UQZPx6i
DF7feYSq7b0e9pQBJuc3ugZOKi9n+H1/7KkUvNwoRyK5C8L5eZklgV60vFF23lt8
MEpRK2LmI/+1qeEKC4aycP6Ac/AGF7+ehFvFzH904oIerp2dIwRVyVBuYcMoVBYE
J6O2vlhDjcGSvavbZNKv2Wgi0CpmnQu8bfKwXwgwUZVWSeSlq61ZfsR+iY7MuIB+
2uS8jYN0Grbgn1OZVl/N2LG3IEcMRwb7n2YzZkNHwdZ+DbjISrNqahoBFuPOk4v7
Kl8UO8mwLOtgFtJZRDHYEmh7YD0Y6G5bWZwt5lneHryuTuU4Q85u5AdrQLUuNLQL
keObLyI+ZgOjLAaiWPPUAg7BMppvs+Y3AEjp20LRY7L8mdU8YGzil297fTDG2FlO
aP5SMA/BkRHXb+KxnCv4ENxvcVT74KhOjxjJMyLsUirRRhRPbfNV/LiB0m7aECoe
jfVsY7ENNNdF8cnqOXNoufy7VfgMAnn8B83uX5ylfZLFJXxqOlJunctGO9yo3sdp
Kk7eJ2O7YziFaq1PrBQO1kOGbgZsdrqWklh2/M03JVsxSI+Iz8pu0vZ2JXcbMR2w
mB2TrKkVQlzLzfGW5i/zCy+4ZtS504dM/6N8lM/qx5ZULjH5TIcntvuOzxlL+h3x
06Z+HnsaGG0zM3d1f952hJU3uakUDI5PX5Ndw22GH0zY82Jd/6KkL7qZxJZM/M6L
QbEecCnlGOtTNgtdmyGma3/gVl1gA/boJT0XFWkjficmb6YMe0uS27x+ctLX8Z5Z
Sk5hsnQX47lABmxQipkj8TfbVi2eRWWMhYKmsECvJjH94pFZi7LMiMHdl6rMZcji
I+olOiWhT4pwCSXxC7sAYFEGEyCAw40QdPTfZr1od0rd6vwqbvSrR/c5XM1ZtoHg
iUFMje5K6sYG+2NwpFG7rZ0Coqn0jHt6QOLcNbY5feb5DvOJOdMylvgEoMjWJ1CL
e636qTBqPxDZ1Jn1vwf5SzGV6oOWo2R/YHbs8Om0PLEGHHmksW38/QY5YoUgDYT1
f93hmVEXzLJJFewkUo24sVcNPSUtXSCgwhKYUYjLFrwMxuRlOQ9jvJ6ohneFZUxO
+M7umsHfk3292SvPccPUuLVeNian4gQrEceSo6V42415gU2NcmWUI5ChDgjCUMWG
hhIMiT+7GQts5I1coQYPQi82f/QYdKcVMu/2xFm/4aeZluQQ5Chqh7ampTlubp4p
2uSXQrRTQfQ0KQDTE0Fdl/NdPTiLqB6LnDZ226KZ4MPCI889UY7QakmW9r2McmjK
+K7ubYNCSZHETiflQFqWwS4J5vbleZXy/lzYmywNPunUOAM7EIvvpHu2Fzn/fqRB
w5a56oc4PNt+tjHzE5SNTFB34T0flLbNZ/+DCp74OOumoih7mhZxhmlFmvA/FPf/
JTtwg84rHFeRVursewtJF0VvBAXifgMng5vjCv4T7Fhc8euYXChkI13iEVW0Mme3
na9Lc6ch4luWUlzrXzaumjyxQU9jWL0FZSkY5teWIqyvkcuHAXhPlsmBe8OGXArN
u21d4Yai31UaSJ7dxLqyhVMbulG6uMu4iKzoZeg0JKfjpNQEtiJPsmMLkWbH/cuj
6ty9AZ2C5Tm4hnPPsN0xJ0UusZ9tTX2Fp4gprZrQKqc5JjYAlxKOizackQIF3IdY
jI/0c56YQn3TskNW4dlYjqVZOXX7xtFpI6j/Ntm4b+z7r2tSuqJKI8MpsfRdPfOG
zkVZz9omlS3GNVlSkZ9AqcJpj5/ilMVeOMD40k1SO9ILAG89Ai2EOJwn2EGO5uJM
ws3OajRz0gvh+7AMtVpEn+fMIJHbAWZtDlIOLFZmag9aVZeeukUd5olrfKFcMm9t
yFJB0lHPvtCTRdssGVKngIyFyBh5VFfMyLGcvgtys8N1vZ3FiANiOfUlEGweYRmv
wS8Okn9zj2xtx6VOgHeKa4/pO/mol6WlGiJOEmuUpMoGXOGamMDmHamTyIvb9Jxq
91h0Y7RlibMo30lp/lNjdOLDlWGqnex6B0D2aXDmJ+D5BRM8Ofl0iz0l1CUsVQZm
LiDWKRpupaLLieBQwCKtDN9qZJH/L8xkY2yuSv8FQdV8c77ZWWkmm8QSZzABCbg0
OaC3SkSuWffmkUP8FpmxQyn2LoGhTBREUPzqtnzTDGE6CuA9xWz01ns26AAu1qMx
+1f1ncm8NylYKyb8NN5/QuTr2+rq75/IHPZ7HEgTlcXw4KUDXNsIAlBXVxKyVPT9
Xcd4eVh2ITqrRPpBoQquKoc4jAuwbQdzjCgz0qTWFj9zC6Vhxdl8iP4IFSgWvXrA
85UDTAQpgK4MprpwVRvZ6/ndBoMt443TAdOnM9vLhurq59gEcf1cPyr3Th0sIW/3
NoAdT5jb81ScdXAPcMMIPYhQh+XAOTTYuOaG0Ehste6eIElFA8UDqMSDw4I7aOSR
nY+LS2LNKjj2ubh1stUVg7QAxoqEUtlC8o/lTpO6qvL8/NSXaXsiN/R1cFvqaopg
uyQsk4SeMLYVF//86qvmygmXCryHK+stcYfgjao1HZettqgwcbYFSgl6KAvG3gIM
JcJmGsKxMdYrfc1BNqcIBSMnuzZC6vlCAD8Evcd1LIcvzZBD3SMJ19ximV37et/E
Ap3+9pDcuJZa57752BiPFtLbIQg7a0PeS3jao0TUJV05btvVYJ/WyVTL5gWQ7DuD
i7Y7F50r4XxS4M9sTWtTKZeanVSkIfqzT4FK9ufszkpb1JTYiQrhAk38Lsw+iKNR
xeAyQ/3jiZ4E9LoKGt9aE6YXpnyW9f1nnQgAau26biTok5nq2uTkGuMyl0Sl9Q2v
WF3ZmqPkUxUDIMuZ9g2lzY3fi745q4g8nlliuNf9WddR0rebfHbh+/TQu8mV4NhW
D3Rupgnf//nQuJjdd5J5aUjW0KKq4ri+B825KlB/HJziS+pp5QDJGyzD5IaWmYen
y5m4DdyQ18BVIb6OqKwuhH39yUWOXbNVgowhQwORKlnEDo8bvXdNvv6zgil6SKfN
L0oTo7yH+2icK/SvGJMoWszpI9butVmnXUtoLocgJARWVliKLMKTv/PM39qe3j4V
6wCyue09bFXAZZw+eNd/hLGqAzKLgcIfzrnXOGw6Mo8dpPvZ3FAHYDlawB9ELLSZ
iEPPoYfIMtlT6iR8xsyuDt3iy0cIwj6oA0RLttpU96+fKof9OHojGKywQAL3eMX7
Efpzlwp58aA7LDzRnIYQyw6IyqNW6er5mN2c9aJCmc1+oMtzNE5xvedyXCfz63gE
UsUn1ENCxFyepPl1IWBoAhDIUFgzfMO8KTMzDn3zy7sf9/jW/eSqSEVLlGV6Bya8
C8jHwKFj9Of6lvtDhNNSxiHs6+si4FOEYQcnHpWHF2A7L35wX7EDKXF2iWi7XCu/
dxnjdonBVFd3tYKWqSUwnqzqFjoRsL9tzr7Qqc0/DrqTrTSnHbJTSB+o4ecFTS/a
VVyV4DGyQ7GhRwtGK13UVO9c4oYVA+uyePzn6PEPsm8pVMEW1uzzh4Tp/qKeEpQR
yKiOcHAbWkAdFkShxl0eCcEqr2p+56nfFA4EjV7HG4V32Z3TtEiT6tjSxztCPR/q
ZoEygbZljjtg7W2lI3cbklPwzAavhLkV5la9gXsjA3HWD+Hi1/bIrUKDF3n38ocQ
4fZvXGnh+JSQT16/2Yw8uCtOUlIh+iS41BKv/eSzMGZckMSllRE7S5dTk3jJ1QcV
Lb0t9pURL2kDFd0xHMsgLPmrp+VnqT85hCXoDnOsnQbZGVSDCFymUzRutd/AB9Gj
xvKD+/Og68VovsqmZzjOSvhlVlKeDtIw30fbeumXhIpJUtTDl35+Og9iphaeoDBF
Qyk7Q/zo1+PrMlkjUeQWes62Iwe61MA5I+tGkHQKx7tK0p0PMboL6qSGiZ1ttYGT
mzBqOL29gWCsk+2B3VxG9QQde/r1h9jxC90ynVFiSTpV23hOeVp1FlmxZN531vat
hUF8ZlK10VX9egA/memLwe7cbot6tH91FQRaV+GndJwomLea8osEhssyWlSYY0Gr
lJb/CbtefPjYV58+nBrufauOR5b3qVBPMQsVO6HcmnmpEnh2/X4KnGvX0qYTZcZI
75wZfzO2jxo58w7pINR+2zBjaE+JV+meBQwOI9MHDPsrAi+bD3zlesIl2dhPtL9j
ht2sjO0KO2YKywxn9psRpkMLnxtx5/8qJuQn7xJuXDfI1h8O8rHVaedmWFZv0Sig
24dEPRQL6cD8sPzpU89fuO4crFrP9g6LbYO1weFK15NYakd63neJ82A+/X3b2VFb
MJ9N6z5Hp4dO6V2YiJ5KkmzPXKc6ERyDNHAXREnz3+ZHPh22KaudWG8ObOJpp9pj
U+mT2lfR7U4mlpltCfq2mbZc/e78lVGBNhlmb7UNQsWWgN37/zK9ZocC7OOcTjER
bS2NgDPQEdvINl9hn3iLAVVsPeF0i5rn6YYFK11p/h27bw8fy1O/X3bQISnqMQxa
hUX0UjW6MDst8RaRJNH8KY01B7l49MOPauN+0Pt4sAREHDCYm//Gz8Kn/nfWdfDh
6wV2y0yaNecjoZrC4ASPOzqsI0wgYTRvgC6xLiileVUoE0Ry0yRejTxq2SVSngXg
Khu61P8v7tGSIoY1PmHq/cz18+ewAmV6oBY7LpKVgyJehfStFcW/7vOevDGNMXPJ
A7wt/xibt9HbNqScU0SIHF8a1xMomL8GpNZCMYqn0ekLfoslbPy5tFKtaF9pPyDx
yoBVvZ3GNY4JLAqVlxv81Yn4yQzLnyVJIrMEtsKUeaO+15QnQ7gsq6OnOhRsiY66
4voXss9uKeyoKgl2T6swUOfYESMgMMISnUMc74GMcY7VQEf6ce9LmqaDto3xOlIF
XOl/PJh2eNo/FitApk7XOPqV95AeNQB6NYGJYweBoA9z2o309xfwwMBlwvZyO/rU
mDVYlJv1+0vgZ6kpXFH3PUrMwUxOvUHtuHzY7vE/NNmBbLkwZAwgi+WdUPjo+xu7
X4N85thpfucv++/KqAzQBHhDdsSJ0XpIAGCz57cuXeTJta2WN0ji7z8pYf6weFJG
6MPZSts2A/sI0vSxlOBHvviKdjW3dCEi2qv4FCfopeXbk5vELaDUBLhYFbp9LADb
XApwrKGNFpb4LQAjXmuGlPNxRi/h3XQ8x25psOD2UYFvHabuxvy/SHI2y6++6UIQ
L1Z7HuHhgshKmsIH3bzqGJA0Yt6nHBgpSnWPrysWje6lRDNLXz2BWUW6TNk5FyWL
Tkn2/ZsIe9XKoCQPj6RW1vUtnAcq/nckyTOVhBL1JmwiqrA4CiQLNgJmswmLL56p
GyvxWJw98fNi8Hjf/+3bJR0lddzPOchwiEJKVMoGKiiha3XK9awgdAkhRZXUcG6N
SWbqAic9XP9qDERMzDVKybHqq/T8ZcUjhg5N8QeDQBDp8zI/SG1w5Y/V+HH5nZVk
6f+sR44++w3HW/75SLnn2v3llwTlu/VwFoY9yjgjrCh5zn0JmSfmqkxbDj5loCne
a13HWkv6q2sRbtTLgkP/M32h2dvHx31StBYwmpeZ6PWd2709iW9SSd76eFHP16Tw
euGy9hOyybxmLX4IUYF4288hoNln9jZfoxA3lWAcfvhfc+AKDJPOY6Utd/4jyjXi
g18kjyAr+ktx5xc0HmuCU/tVpdkcB4pV14V/XzsTg/oFNX70lUtHB+0g1Wgm7GPL
wPjPc4qQpcJOg/andlFBTrFJEmaa0GdqzuM6B2qTF8Gw7EazIh2aW5lhFcaUj8s7
9onf/mRYbUou9XvOOMvCjoA+NqSU6Kgb9HNtoDA0dGbEzM/dWYuQgkzqcpYY0dzj
/qctcHt5ERJq+aCvUNK/AbdbzYtWfcmlM+RoFzB0vag+JrVQxYe0c9vxrxl1la96
fCi5ckHi2kHjOAtuSha5VYcQ8PXDhnbTbOniBAgaZjqjxZmUj5i6GlrZTvNA9MR6
FV70uLUAtJSOK0lXud2/AoWptZIgZVhdGi/MIAVPTL01Kv0CWXzAN81EENmaU34t
Wue6CKtbKzYJj/ARhAGFht4jcRLqkiO3hb0wvzEwRSkSp++369CdtKqv4qlsQ1l1
eEi4g27kmwv4+Vhwj3wCtr/euzC76qoxZUXsfVHj9CsVoLZ4ypQYE/spUUC3ujWG
GHSegbp2GJ3YRhSie1dSAYn+xMD7VwTr/E4mhS4pqHap51CtC1e0r31FCa1KUX8b
rNSqFPgScHza5nZp97/K2Wg1Sx7Hq0d6/p8cDm/VU3jwJ2W7GMT3wrkuIK2OpwFD
7DhrBWzcnHzgszjmOWXYmL33k/mR5J/yuks9kgKO/z0euFq7eKqn9Oj2pnNUw4yQ
FfwIPKrIv3FlWjzDS8f+mPInoryX6scWlwSOWXMg7k6CJgXtunQlBy7XJUI884xJ
jFAbxT7cqV6m6LQ31a0XzbWtT9fpXyKw5Ba0svFfLuP8GQ+Vfjn5IkpvK/0eVgHx
nPXs8L9fpvuZCOQrV6PtecOJf2zloa8gS4DsJtagekL5Ce2ejwKqsi+m1ge1SjKU
9NB5f/nxpCKQmukntcBI7ock4G8PmglM9eJhKuWDnpAUfCC0lZFJ3wX7SZgLBx1T
2oZDfQUdmJ2BUdieD1uiOXIWudhqjBi3TevMZjED5NZJs46m8l2Xg4H+Hlcu/xpN
Lfu3Le3UixQzpFyvkrLB6Mw3gQQpZ6XWosV4VDPJ+5lauRX+xlOA+F/k6/CowUPP
HVwv5w4RzyFsRB10f3SsRYNoTpy5b8Kr8Fc94ohbO+qzCl/426Ocu6AlvaIGun7i
7kb8d1Y3b9Sjm7xdG4WqdJ1phX8GLUq4+e3dWJVAeadgm7uao0WV9lrzuRHLww/X
qh+yki5Oux/mE8f0uHoLajt5p7GudmdoAcJ4nuBAR3ykfYcWFLTKM4R1zKhoaFqR
cKzBgkFqQz6nny5LrmqzzaXUo4dINg/dQP195ypkDVX4Xtm5NF58HDcJ8Rysf8C6
ay7AweiZQzpbMMKTIrCsDY8opd6mcobqbG0PE+jsYqQAoybbRRUKXOcz2rbN2ch9
6zP+lm99laUCEE6/I47iZAbILTV0NBGj2xqRgV2DkdrWSZYvHliorDJ6meZ5b4xU
uiSbw6ZamL/CFZ9V1p5Ezq6KgG9UVfZRNF5ebpXOYwhWTzllj8PLZHv0WJHaUaJF
k7uypF1wq9/pY7Q7qqRtgwuLcrmmU8IUvjSFdILNnuNQUkzGF9QqUezNkDSgiZx6
uAHSg0qv/mZHgbZuPCb8eiqQmmrbTrOUfL/m1minyEgkc2jzSZJBRyvin+4BrmPg
crTseEbmYESfnhyhpeEQvcSyNvGQTKu5v1z/L+FflbheMG9J0ANWUVfGU8mZ4Obh
upb6vtTFNHMYCZkSE7WagrAA/M7W5f2Ebxq4Orlq+dBP3LMWi/DwvWxMHS16+jVW
3eIz+cNydZ9zaQSzrIlIHlsVn3UeMadusxNVpJd9z+eDYg7PzJO7QFw4OrDzIqbe
izJATdALFs+6XLbbN9R8D7a2V/YBHgvPXx1RsKuAcWIxMCIaDgOqbdBE1RA/s9ak
WkeEEtl2NjVh0KlcpDmvqmPxv1wNDTpil66+CBGKw57h0eAn3J9UNmgJfkTzzNxC
uCY/YdiqLxkGErIbBnMFXP4sZkBnTOk+TNd9NaO/tq27bISIxg61BDz6zOKn70vk
Sz9irCTlz3ZLLRTwfSDsXJajk+6uYrTepIkFezaCv8STyZuRMETaJcqo6IJdA838
XLfEzbdfuztvuvEZ/rtaa4g3LuJ9EQbdho9vExFkB5E44QjHxHkmdx3w9XtbYPQh
fYvrvXhBNlKXlvQQY+M+FWvy3Efjed47NCUYgMAniVVvzuch8er8f5wLDF4ntY1b
7+IBN2AAyAZ6g2aANUwFtOpzquBn5nwDs6gWyFPgPNvLIZaMYkImUOxwmUYvrbeE
U/MA7CfusHTmkRWbwtTZLSSRsAT+KZb8pPtlp/cST7szMM0/DYYORzgPZDaS1sKO
jPArUxQTvCVVfsT5pQFENS/fO8IRLfSH3ipNO8GbO2dkZ+ASbadC2EU+TgmdkY+5
N6d3oBwUw+umCslMqwvX2uauGbqnfYbAhDd4zzsHzTPOpqfpkiIi993vWX8R3BCJ
MlVv3Xar5C3YOhFsuLMMAs6QA0LynHqNoee1dxsbAHkmwGfA6KYrHBDDxqBupgfE
R8R8F7r3m0AZl+ku2b/6tJ+3I/C9JAp7x93O2k6X5ptT9S+VJnDvpJ0jjgDVJMWA
GxbTCOm45FM8M8lFTt1G9816OJ56A1sbxu/i2IG//OjL060sqegknwZjFuWzpi6f
9YhEh4A3amUeOvEnJw1y/KysoAUzf7ZQ+E41spGeSbWzdj3TNBI+D7owiuE/a3vZ
a1ti6ASFak38DFm7lpcgzM8ia1vcux7f2dOz9Q709Cc6RII2uUAbgFDedkEruUHw
JERdC+E+2bpkpHpyGBbwi0D1fLMM2LMEXqg3/ACBsuoLt15WevtdSkTB3WSDhWqJ
VAT+Fxy1TBpb7IFiKAINbpH4WW7CXGU2R1hUOcttT0urLoG6Blo+uboO7WMCt1GO
nMJO1um0XILSfsvNWnauIw/DPoJEMzsBM7/XpR1/TiYVMeBfRN/cfZSzGoGyqEE9
qQFt7vsHOA1m/IPl9vIBx4cg2B68c0y0LUV7ph1ycQnFUv6dEu4sJzNvCsta036a
ATYV+/0VuSBfe+af5I/U77Jg9IytMDqsTHbAO6jNaUABEIvL1ctZwiU2UGuvI6sk
KA6HRU4B/IWgwE00xTuvUpLrpM4tdwwVaEuoPKftrxT7PudnU3QZ9kSNR+8u5eQF
wIZI9KisQ3gw8wRup6zKw0cSOuzV5rdVCO/ACduOuZfy8yMWPi4d+1HZ5lrYsss1
HJSJXX1ojGHlEbbdIivXtmVw8xJiAGuR9b53XBBd9Adyrys/wz4+kJFbSL6mYEm2
hriBVaR8IGali1kzI69LMgyKEdufa86s/w+vfB9oHi0WScAMOBuBWaUT45xJy/GA
kIpwFYWmqYbMzUT8TuxPbJhdLzjpqHJhSv0W/F9rSVIdcQqwPhWyAwuapBUgipIR
PLSMlOU1tDCJBrT43raZRX+XDnR9GOEsTMohfZO8qNenIf6v580fC3CfPw8NUmE3
X0rHoTDm4g0UkMTgufLM2y2ezvcdoWeyy5jfgNtrsDsuA5dkq5Uu8MA2o4zj0KyM
cF9rmt5UAIOxe68HVZamiBE0BLe//P1lgkvp172jf3OqccRnBj+cVa1i9ziUJT2C
7bTmsCfIZ/U6QYR44oxI/5lcYjAnl+b4myziTeksEnDhLqhm8t6c3JMTNmYvRCHD
oY9PHd3k9cWW+b5voGxGALZP/NYadbnyYbvQAqUKjjlUMU2a1JbWxZjGk9nd+h3x
0f5uqkLnH9qzm3mm52gsRDQaBGZhLSj0nl+x+m5ZlQcln3W8JZjmGgTkSEFwCI8e
NbhKR/yyjxgqYvkWZNPrjh9K961uO2Vi6MbemtWvDC5NrfyswSrfrSORg3U4Kfux
CTYlJqoNwf9Ii0wE+w/N5uAL0DF1b9BWd03x4w0bB0oC8/MdJycMwdKhT7/5rzaE
BLLlWLkZznMPNNfe8SHbnj3FNeJjHEpYyUiX+R5BHEevH+WDZcUjacPM/yCs2IlR
/CVPvW1qnSY7vpXixDudKhJTJS2gM30s1qV8+f9vEJbcUGmlKGe3oJJovpvdgHai
78KYsOZKT67W2gSU5SeiEKk1Ne4vEe+zIKVJc4Y9xGbGS1n2TX+hlaAUDVVZOTQB
LVk9NL/dZDAo1Z5P1pkZ7nz1qpQdqnQ+DJrTSgjLEaNuQHr5tYNMZ0YiY7QZxe6q
T52HyOnWYfv/lEkGF2tphjVhPw0jf/7KuukPkFFXuVOEwM92yOlERjX+76YBaWNc
zOherhUXk/Ofl+5MpJvNcZYX10ivRz1qCrIouX3NMtE2MRnCdUN+mSxf/fMhMcFG
j7fPCtwQovGevfy56SMQtVLr+dmV3HffOZ1keyuooXTiHsxII/z8K0/OcPqujVCU
tNEflQgqwKsS9nXOMT6C2HaWY1sQNV4QeX9Zm8dkQQH80YszMleJOygiyPBmvqiB
dzzkgQSgCqZDh4BA43F+Szfa9yvAboSZtt5laMJP/bWD+Y/g4RQ+l0lbuzZiFlWg
SdIgQKV6c5xFoQzQGKQyt17AKbW2kMUUW9piriC4/LgYASxaN5gAQMHtpt4iZ9bQ
Zxfr04u+6QaLISFWXX8fSfttBGwlPkuSftSg7ahiqebXRCKisE0errBhgvviHq/C
fKq0LWU+2L9yVOPnwZe8pgDA9yO84GLIsZJp/G2M7dDA87r8tf4j57vb716T7bVb
HfcWP9thK/6R1QzDTObAM2uwl5epWSL67+iAuKkM0MHJr2nThTe1fGS9OxeTORpo
IbTVgB/xLG7elv08nUm708wW6bRi7sLUIm0y6pOeENM9cDmgmlkFBBouIk0Wkidi
4uuyAOEigTvTl/aB4e10tVgEv9lsReYdetxPBTEPbhNzmHtN69zvWwDdRXocACRz
leBuTZ8vG4Y2HoCIv9ujvzW/WqPf9ruDjWjOYD8ljnPEFOA5zy7Sqe2KxA3ZTngp
p04rHTwH1IQfHmnIQXEsmKGeVs+ZXN/pr46gkTkiQUDpo0o1HgwVJep6MeXdgs7D
p+tAF7vyMIJCz2QbVklmOOTtM4qq+ovmTGqWL6Pvfb5+A10f7qnrNS4zouMygW9F
qtAhGXfI9/OPqcQiFFovOYKVP+ZmwmUG3NZXvJIBRykU1fElFBhTuoe2qcID5w8d
f7qlGkgAnQM1m6sO4odW0ycomkXzQECaTEzWCVmiLiPuO86efmBovtob3qUlCyQC
28qOa95KqRrR7tJ8INXEya+d+V04REb16U7WciDIPD6h1BjrCeDhaNJLd6Bl5OEu
W544MCj48HeEbP6JyIOSLuqU6vTZnPN6cx1U90rG8PeirVtgv/pLygVkGjQEji5V
KSk6bnWzqYcuNmox5dRe1VokMyxl4zE5aJLEK+ro5GJXyWuWpG67yZZ1/quktYzd
FF2y5aTgtsDnoae2HWhGv2xuRjAJ/J4M8c/5v2AOz0ZPTd85n/lFmtQPDtz1CoKe
A14qQxpeUdLVpZBI0sBvfNKqfgcJHar6AjMPV2NgZrUmsZgbINYhwxWvZeIwermT
YgSBTgOtmmUO6/nYx8nKa0qYEIwSfUFLDajtsOCjjnWalYapBM7TTRRGgNeRsaP0
EO47bO8xyuQkjY0URCSZeLw+7jgud+tqd2D2rGSgyS9MD87sqNPb46ZAWVNDtqpE
PqAzGCaMm9Ryl1pqHv1ozfQryLMbZXAb/ifyLc9MI7nc0JdA0SGranJVgQD65pNv
p4B8PhMUpGctdpXSzsK61p3v0TZkdnicmDS8QEMSjnnLIfW5X3pyLXP+DCnzxUMJ
wQmrcP3rxYvpbtZTJriSVelVEGwR3G3zBTQIdGDY+EyvSLKoBTPRSxjry9FHF5us
CW7GMDpMI6E76ZRo/9Y/d0azQ1QEaKpAjfKU/HaeDPwEB7oI7KPM/nvmtGgURpcY
07F95BE2MVPUADn4AEywUQWqj8Gnpkv4Rx4lYTtsR3+4hxZ2JZ0Ca4dN4GDqupVR
Uo2pIJZCg3N+Mg7tgCqVmcq29YrapzWqvKIQhKGdlPZIqmFij5zfEmqahCanEVc6
dcW6MYwGSCzj45gUiEVhk5i0c1dR2GEx4P+/9XG+vzkMdZcsz2O8++1caEEn0Wed
ZK0XxJhDZNfn5u3VvU/ur7nZGW+R/GTjm0/WvJXNKNYstw2SrETkMTvrkUUcOF3o
0TeYlL2Gni+MTfngD4T1suTuIFo8GFcWA0MdyX4+Joa+Dg/ZVNGcmDOpYb2920OG
tgRotAvLjm6J/2jnGDegf1dGfdttqKUiPzvdWNhKSNnFe9dSkzlIBPpqU1UnRbfw
mXcs10Mvv7cih9AmmRkZ7ZWWPD4MEvajCXRn1OL+XxZJuRl1zcY1sjuZ9Y8rKseO
qLXiXKQULUZwuofC4yIFUp88W0uE/FsMmhsuLFZCmEnMNWMtkawyTf5Sa83sSAmo
U55VgNjkH8FiW3e+xDbxntFPs54uKdjikXGVHJyhOhRNesKWN5Y6lktYVVwUx8AQ
EHdI9Gyq4JP55WPOoMC/DKFGf1e95s9clqCC/ZP/VIIZ3hNsZC4qLbobpxv/Dwyb
LrLG/eCFyFihNPlZMClluxb3gKZgPmSgzre3x9d6RAtTq0QHxLiGB3HBz9QyUNB3
ntt/sMeqtMCxyHFS7ldWeGO2VO3c0iCFGqdCbFNwNoXeJRoQVZYXogmaGT0os/Wl
UcdReEXEK7NtUs2pdCBVt+RMs6GikAI2mxjl/UCl+XpDlO9oWwdE/eUEB4Ty3R4k
gY/fjUpBIFS6g7npeeOEK5cbPWFctJCMfRdolqpsAoQ2aIzMM6CJOL4mBHWsWH24
u1LqnQHH0jdB9hWBtPrAK8kgtg8dO01TPV8/zvrW4lYjObllo1TWHsbQDB/LC8Ny
YcjzP6l4OJLsFvctrmcUc1vDC2xy4oboIxXvj4m1OEYFiwo03ifFnagu6ICCgA3D
ZCp/Lt90nCz/TZZUhPIRfdSa6ZymT993cfnr1tYd+EpIbIsgOqO1g+a7eWsNWJnv
hX4Z0wWUuzYO56GrTCWPBZwfF6cgohnoxgRA7eqz4psqaGPvbanZmv9ao7kGthqO
z5TuiwST0HK/84AdNikrSPJmY8EFVCROE6Fk8nwmMRmAOvN3KHxFMks3YttaW4a6
7/8LCZbBL5zTqcoS9P1VhewmrIhyOJD3h3yGvt8ruQo4lfXjVXDwADXhoaeN1OcS
AHWWqthVc7KZvHZj+MiTc52+ixktkinp4LWQrl0iSvKN8mUtB2LA8oXXoU4RoEzI
NRiamEl+BKMf2yVE64xtF8ClZNz8gUPvF9JtdzFPskMpS0+Wy3mzCrNl3G/gWXHy
5HOxRT3n/83EAcwLEVFLMU0H/gGKuODuJZ5S8E/ppoJVa1NG8tUcXlOWQVBuMjJ2
RsSyb+IA+nos7td9wdHzLn+qU06z3ete/EEGz+43gfjh8EsGtTqqhg1RhnYbbFhv
JvHlqADsEQKwPeenYfnY1mJUPmjQdBAEWTvA15iiDY1E6ndDJylcGGpxPvfJ/eyQ
Hzn/BH5Izp0psLvVo7yQeIms7P6g37C/9cZUDktVxhuT23QzgzOSYaY/JrFgsvh+
9lg5LLke9l91z4yLIM63sShdWYZtUZ1nebBue31ZPnu/VGani16ZdQdXCcy9U88Y
W8mRqGEmcsBozs1OR5wHzngAByZnjo30ECUomFc2No5vTMn6xkK33vNFRk8h1hha
Cwb+Wi07Z58n94C32yofFrSGwNZDiRYgZa56Eyp0CcNet9MZ2cHk8w2668iAi5Ku
Ei8oFAVbZjcnZ2qiR2jgQJzpC4OAxGgVTkN5bLRuAOYYnvqg1fjOMW6LBAaeOLVb
cjBQopeK0irpx/EtmRAR3Kt6BFfwE3XWm+M/+Ufy0Lk/PkEKseII2C2sip54ftAN
nQWRiWc6bQNtZCdx8QONNdbokYi57aZoJsZmtwdQjY1Gg9GIKr8BtEQKHsh3v02a
sJGrJ+2Xytdd7A+DAUJ4rwUJgbm/lJogj5k856Wj/ewGWtuPBcDivOeui9HqpN/L
wSjrhkV5WJbdL56/uh8ZPTKlLamxO69U+0rlSph+9pJqNGWerwjTXfZ35w4T1q4V
PXoeLkjvH8Wwv9rMJ4wyhUzKxBEz6uE+6zPiC9cSFlk2Jx76+MQcjG4udfJnVEGX
DPMGPWD2Po8b2bkb/4tM8QLxTmx+DgODN+HeL+zuEpFkaXFjZYD7fUBfqLDC6VLC
Xnic8nhaghozddBTKzVgFZgJNRQGn5iZ8IVIqU0zs5PTXJwtZvocNN2qyi8Y4CGF
GuNI7N+32/gn6P7jmXKymxEKp+eSrnj965hIy2ENDFrGNtT6SDskNxkFDAPxfR7y
gA6ZBjTQpCwHDEgc1vmiTufqdeO/KTY92IaZ+q3Su63MC9nIiE4EXgWz211qdDmK
oaAjBvvKFkxkzQdR3hICqJmuYxXaPn2gPIEWVs97uN/2B9iNm1KbViAwjcJ0ImgI
nBaQzQJx19W17h0D3iITMMQrgTeIl+oItLzV0jmPry/xtb9Uk5fZjUSsSsj98TeQ
Eoys5Y+qmIqtXduJ2KZJRZSCTXLmEo75Y5QuzPp9shGve07Uxj4xLQP4ZEbgyUa+
FM44zoZAfJsAZo767jy7eHzExuTqumrRnkweeIFB74OXasjBvUEKMiv5mm1U3QMP
j01s6gyIhh6o6zJN+Gm2tnjcI1WEBJzByZN4WwsxQ42sqwbBalQc5XBUsrZf3zNK
lApIur4i6Rmdqk8KADbDajiRuufyM7/kpDheob5e7tl2QpvyDjqh5At1oBio/p0r
ywBrbIwI+ck6HNdn1sdi/tWFGqdBQR7CyhWeIFg64YziD1EBGO+8ZiZzEjX3Ge67
XFLXb3Qp0YmdQQlTXZTn/nQ0xNiP1815Vw38M2ogBx7zBnx9SgxPEuCoibfMtG9q
6q7H/JZ+MG3euBSf6jI0wVb1wyobg2HOpA9PQDLumN8ZGIHJUR/IqzFYMzN16U0/
WYugcmjXUG/HJ+/fV6a/i0fpCtFCGb60XQgAIs8nzSTgCX+59mn6RdNUvT3tF1Vo
TiQx3VBtwQxxvFt8bhSZbwFOv/zp7xJ6wC8AjI63sJAOFHc4Fm4a67Gbtp2CcLe1
Sb1djMTrzbXEoksEv+I77+w/LvTmUnoXPx7wgqYaXPR45osZyQ09hCjSPRlxi1fI
YQ1MBpBV3Otzw3qIeybB1pA9DG5voHtGpA3ApdisL8UTnMXvLqmm/Uidoiy+xye0
+50RCSiEt62dJF6GlPsNsoXrtq1teDyBp1ZNEHwZqWNiIAAIp4Fw+QKOaYePKZIK
7Ptmo692q82MXRK+XPMQoYaautRrxEmJw73/NbDtBWIBTr5hJXcao+qT0UjZb/AI
huutCYbzPYIWlvlQZb0ThSE83zhTtb/MZsBQbpTFeBNg++3cCwCyX+YaguieEkvC
+QOZGNuuowPBnamPGfHbFqOKrodDB9aG1dHIEp/5q2JZXs2vHPLzfN4OQ4+MxFQO
RibkSRJ/6AgUnABE6GZYPGh9aOhHAoFlCJfXBIyUBLUrX9sFjcrQtSGUYFxwL+E0
GOSXpwQfC2UgiQM8HbCgTaDSS0Zwn9bLr90ZrQpXSDzadpbft0slw2+J3Ltiq4F/
4mCnFdvbGmrKHphKJR0vfYhIIM3oYSRdBiYViYrDtHjgkyhVb0xK6KdIYxzlzwLh
lgTGqgoOu0Wm0MdTdrPb2mc2/H1TFxaiaqZIX6ZNpwc6QmozzNTzJF3OzBP0vLS0
HnP8+yHHLabG9wmbObMB7o1AL5RguSSbF6GMjhHhMKLBQe77+BWIzIJDr3e1NxHC
4r8jCmUve11kORIrfeWjRgCoFhEJX8nft4PuSppoQstSHS/vTu4szypdlcLeBCr9
+8FLRKcHUVY/veWCb26GmQcgER+TBrKYVUfpRhb6EifFL81Fe+PIf+4U+WcmF6Eq
xlnAO0K4XGT6UZAiFW2i5dMAJUoITPb1Ln+PZ2N+RKlo9ILpBwnPKFoMNy/a2nTU
N4V6LxF9Ph7exvA7WGgQhoFo4hlAmbXvUV4orQw/Gx21T1eV+vp62bcc7m6jAI1x
whdpbeipBVxu1C6NS3I2UQDxtSDY7LOgg09VDsWcyPvNMEYogFEKuVfawLeUfn14
TXBAkb4bFDtNjruYoFhhpdvA+nvPYx+5P+eNi3K0vYJppk9NFqLYjr9IkKaF5vUq
q9clala/5BB/y4/KYBr9QQHYtgz+8/xdrMGlAngUqp0PUcqLfuhfG4s1QredtiFx
TxYgSCMYwYOgF4Tw2pJTdPXXIRlaYPW2Qpxtfj3cC0D2ie9/wA3Qac/9iKOUHttW
AxdGCELgSqgxsNEwFLL/n3Whtf4HBdkjAOQIN/t4G1MDS8b3fT0wF0FQm0AQSm6Q
zpqVBz+ggV+/dRnHWSV8WbiZO6yscwo4q0Lizs2ZfzPuWiglheG6kSH8EeDB6tzK
t9Uj72T3h5O6Lvsyn2ZfRzT5t/YXu77XAYBnUfyZr/QtO3MfDmdHqHZ6MMAlqXo8
YJeeFwU/C8MzqpWeBSMKsWc5iQCPuy2EL64e5vM6n5q8u56aUEcrfHim075WLbxA
js3ogVrTcJmQKDHD5U5/uts5p6909IRVGc4dH3kpC00kRpF4E36nImWxOjl0FHk0
snlu57CxkyPiIySAUsgIVo/UpbJUO/EclkDg2KIfDAImIn9cCun4nMGBZCp30TWn
KJa1If/KqrFYd0Y/TJAsnBVrGfS4aejJWVz8AwT86veFM8QXqeFexlR150dd1bep
JCTX4nKbRvTER5v4ZDWrckCmSaYDfZeTDI0fKPi/S2dk+esB7HAzVXvD9eATwjKd
dcjK0lP1aK1Srcsp/AVyceuhAL2wgBC9WjXNczWTSsRG/pN9/EHjS4idbsGUStWU
1Cj32hRq+Q8FyFOjrgAjdgVr325e4kir278OqtucrdwH2S21fgVS5zEK8T2Dr4lY
j2Rfcf6n9hMZhJM1sY6aI1OEmTQtEws4xWnQuiEI0VKbwt/wDoGkwvhaLgGW6IJ4
I8Dn7Oh4kGnfYvXnR803uScBtddW1THuDJbtwqEkkM3QFPYYvcyhmvoffxUVj0Gg
GigFU3WPI2TlXZsQHDYWmsPPf5YWiC6+YdCy9rG0bVYqxgGtKCSzyCCxyWQrTes4
jjuEywTXlDRjadAeauvk9fuadB7RtwRzoHS2m3WNJTKrqod+aY+NEgQZHQIUwStW
XHGg6j3suDWBhfhwVsE2UAtejbgKlo3+KGdOluGhMZ7V0X9QL1+Qe510dLrBMBnq
/t/nhqVfTttQaZUYEgzYyZM8iLI2J6GL//5aUgXa69YYQKhV+OhkP7nfdMFynYKF
vYuqgA08gOfXftDQKGNAjUwnvrBEq9cdKvtbbYYMEO6g+MpAggUlCi8ay/oTY8x1
rQ/KH+VVSp7/iw/ktfbfwz81jc8+V3H0cYYNqqCW8utU1mDKxDaXaOqzWpTaYP5u
aD8YLULaI8D7ALRByfiTnL24bT9xVt50p043+y7lCnMR7poUqUdmojv5gQzQiTYM
hPJyQ/f6fSKAfvablYdSQpd7x5+yIRVnSNBf38e+bsfhyb3IRTnEPnvgT8OBtfIF
IgPCYyWak+D4a4D8jIkRGhHfYBPW3oF2ADFr7yAXkAL/JA7fR69xaHZkwklk8aVF
fNYOJitHI+Q/dcyqccq2FnaVqwfv0MCF/BK9HQfPFEPqpRHH2PykmXJJf8MSlK/l
DBTUy3ILLIG/6P164Y16u8E8rqCECVLuW/O+Sn2qCW/70WVlrtfU5gI67ieYgBHE
+gsVsasYV8SHT5EeLAKe9e9tCmepU0TkzWlDKToMc+2V76T/m9SHdYk2gQCHQNhZ
hQpTJTGLeZUzmBgTlMhINBBn0GHNW+VpvqNT+SZKl7x+bcQ12RdChpmAExtNdqDz
dVsjplwvx7EsIjG264YMTvsnDL5DJexSjEruaRAPxKKBw1LsU5w+B0+0cULnhIbz
hpqDX4jPZoh61ef2GggWhjN2J5M4DnQv+CRIMdBT5yhPLYMR2+yRc9hZSul8yTsD
6v4YJWCjz4lhNLpfykcUdBJn0l5GdO/czgqgWjN6ENfLCT53oOF9/MXThBK1kGSM
WrYIcyNo0F/FCa6BxbZX/aU0tli4Qg+r7NfJN1fhRUJU+Tq1uJYtaK/zDk1XJB0O
T2xgGt8ZiMyyemiQb5RrLgKFRPESx2jnS8FzeiOxVYn9ld/kEaGhk2I2U1130sfA
bYvLKJL9/FEZekvHA1lXqlXZJINDFfC3UK4c/t8ZOjzVcx85V81btO4nnqw+Q2dm
FLZkSBf09OcDbUsxNujid0t7ObyZav7jyGfnbk2feDeTaTeVEpuzGdQk2/0iCA3L
Y8YT9RzT0+PFo9oJwq/UUXlv0Ma0t9BjT/eM8uYv2pNcZZA+uIvVzNCsQxqvb8d3
Ngi5mA/tHwvxdg597WqJf/+lDEAOyyVxS1UXRoibpmdVYzYBPUYJpn3jQfeflmKB
pAB2lHLTHrzmchpXSXNFcP9AP3yVPE+kjkUUkSeJtn9tgemmd/4OaESpanlO7KM7
LWu2rpRnfkm97H4uaNR3UTHpAGiJwHz6V7didbqMwqW+r+KGeaGxVUNUgxtC0pWx
wp/ahcteYl3XDU8tIFjKC7/hYEbr86LteIbdBDCtsDFIjqmwy3XJ1ugQNbhq/P0O
QIv9LpJ+aVFxTO3LyTqhQZ2gB6IHmElEcYKNvD+2PxLI23rPp3AAt+1wGP/wco0d
9DIMDZmziBpgx3owYc22Sna3gaQoOppNZf5ezz8WggGw0fRnDRY/y0cg8k86mWl/
HijgRkcUDUhIo3LbXxSaV9hy7cY8cKj4SaeXWXjmpwkfaZ+i0vrrmoMHK1rCtVBW
r8kAi1ppAlkPijH8BPCTlihJzC3qov8SolzxN+SHC7OAsgB3xSoGS1UybeqIgZUk
v8oK5XwsK+geTrCps86rLOD65Tb/zEVEYfYsewyGiCkLLx3te45r3XreqbCJunCy
mpxaoLQ7LTVGTAGQ/2PM5IbxTTY421rYYzIQGhIvPt0KXkZacLy7Tk8EigQaMPQ0
qOZNF3ilRaZoX7KdllYSfoovpn6DRl/rg3OeYWh/TrsUhgsIossR9w583jUDIbsF
Go2CsnZC4cI4hkvPKbL36lGOzROI6hUJhW6cf7oBDSUCRcHIL8ySjdL5aXzazg4c
91U+tziA/3KSUV6JLwdwfUC6OKeESDOZyK/boY1Jf3Ed5O9J04TVKNP9kbbbSz+N
GK0pBsdkYiti1xLrpe+24l50KaRreOVuVXUSvlCjrehFjDzs1r9sIFhEdWASKvg/
b0hl3GB68ROoLutgQqLR8qbmmd18QTqC+J/k9VjfZojfpAphHSeAQWHxDvywkVtD
0qBKXGMIEjdbtrkTJQ+C+7JbowzP1dmmwdRyf8JAaplKJkq+ICI34bLoKik9o0D6
V/7QuOmc3IYo134XiR+KpmB047a17J8WuY2XN8SSYirmGjBzJKBWRs+uAjl9rtDT
1BF8R5tjcZ2Q5stT0NB7cWtixH8Wfv22DDt+FU7UTQ0n1wmGqLlcfS4TCru9Dv5G
LHhCxO6AbXBDVHdLCoa8MYVALwvlkAu91/YjaCVTlbRONtXmd4T9e0dGFUiQRJZl
6Y2QMHchoTMtH3DQGRwHkHV0tNhSaqrFe2VI2CoXH8JMV+WRj2XsTUFeKx2U1NuT
Gvj8bO0jNeZHevEWbeWuuyuh4N0YoOZnmwX3zpidy/XcC8UmZYrn/WpmXlr09vTv
73XuNJVRux+QcEwA5HyoyHj9i4HxqTyQvFbExG5dIU5qcDeYIiQ1z6PB3VhC39gc
j7nC0vI6fkwlIvCUvigVbrgDMv98dja9WzaACsRFGzfQGQScXybr4m4P1/n2JmMh
GEJzBVTRX4iv2AyXZGbVbMY/9+pjnaR+eStgr0yskHpgpj0EOblbw6okVSDokJxO
p9Pc9o8+Q4MOYNY8t3VMhw06ONIOEIvkRlQnB/3HTWU3LqfTCEl52jKzYwf1tuj2
GdV3P8zwKB+yiM74Tb0EgKEe9dFQmt8zkBtClJVGnGg/dKxFqVpOgLB3iTrbq+jL
qWaym+CP9btXzF9vFnTox8qb6xawaYZsnoMOif++4uM7IfgyPsiIp64JM72jXbTh
wXC7S9eIGhUTgNnO2CZfo5RNZijRa94QqYYLNTXlewpG4T65BoJ7emtjDIjuL55u
zAM8fisq1MJ30Mz299ACgO9xS+JIsg7ts/1RcIQaBpxmSLttF9TJBWRJvf/PxXqn
HDMPNJ3x8G/AWrckcXDZFsYhhPtLteRePcj980CW03sotnwwPi03FyZ+fsDRVSqq
jsuXksgqOwcr2yrFQ9R5sg8EohF5DkAVwTIqwZswrhRF3IrBbA0eNdywtDbsXnX4
LXYfRu0HetCTw6LClBQiaCO0ZXEb6PAhsiPOCWSsvsqnoaf17woD5ZviEgUSV8gP
xTyun1OuE3W5KZZ+3pfOxbWDA+U09HgKYieYA6kg9xC/mT/h3K4w8jp2OHf3iHuk
5LlyMPUOtf4Dmc5gZLLbSM4xEwiJ/8Ma6wXelql5WFULgnhYCHZbNQl9AEgYGwIP
LO/+3Oi1WsyUBoQObv0Xjjc97SjFEInqyRVuT/l6U67Qw/nvv/HhjQ4oICbOrxGr
pnwHmZXH8Fs85XPyHmZzsIOGLluZd407Exn49wEhwnNBvgjwrMPn5oLtAd91KcAJ
p5jc4gKkSIdXdajpOllh31K/ptE/gS15WAJYVvYo/zK1Soi7QUMCWVlXQRCXa7iG
uMAD68oz1aKsa2tDVTqVVPyG/3qYcIh5s/iQdxVSLsPzW7H+oDL6X0y1McOthRCa
5GZEFOXvZ6ubJMPoeGyfItOp01LhmmqaZ5QED9L0ejeO2UH9LVVFwKY7dWbcGTME
k/4CmPAKqtsN6WwOpJgvuAbft7kgQirwCv5HWfxkKqputILW4P12WS9rH4SOHgv4
9LtDT0BUgGhNK7Y0AIbOVQa1ZRo29GDeFeiTj1IfY4o5JihH+xgcu1vPI5tW0qS/
6aWkiO4VbFmlkdgxPK8RXS47H4Cwe3N/FzNeqhF+IS5td/9GV/DeqE7mlXd3uPcD
jCfqSTd0NVsU6OL7PfZvM5AJL9zwo7GUQ5GYYFQ4LctjcUgRtXhNWtlwTDy0Xd03
FhRuvp4Je7B/6qujZlc46CsvXC0glXm9gg5QXemWvRB4epeb048hF5aEhoReq0ya
ODRD2DOW15GMZxNMd12px3osvfMbpTjBAY0Ezrs8SfTFOtsONoukm/0/A7MO/HhW
N1nCCU5iLwLBqYozBozPG7vTt+Ml1OslTakIP7K+VKcNHe6oIrzmSlLdXHjLMOrw
PnwFhgGHw2piXzUZy2W+igMR7eaK9hT5AWbzny6U5fDA5Q2C+urpTzHjSd+TybTS
nnmIhqDjnxSr7nInXH3LYVS5XTRhb1LMyfN1p1e04nlAZuAf/JP/KXWgvs2uEH/B
1VZQ02EGEbDBmRyW6u5qR0Fk/LBXayQxFtp5zp/DdsEULDRHmedMmRUzjwc6tW7k
o7PHGlOszNk2ak+e/b3P9+p2xmCDCoVGVbH917fuER1lFLQvFBP5IDiSJzI79gm0
lK5pWCz62b4YFa6rROjHlI4nGJhXnTE63loK+F4dHR/KQklxrvJ/QG5XVWO4txYT
1qGJUBYmT0sw7fIO71+8EQwwIXfRS0jItvI3z7RyzIqhWnxs61oZGqr23/x1UkUl
N8j1TP404K92BXhmVXqYtG2CIJI/nUWg6mCcvftAUM/j5a5aJtfJAtv2D+9gLaK8
spRImZCnJ+b1pTL7bdjWNaogUCNL1swQ9aPDANld8OvQGQD7zH85MQK6j8wuoVB2
9YIjTdYnA14tCiKUJwBSWnGfgoTtmzEbufzL0uudmKUfqDoxhkc6vimzEngaZAab
OnCiYq802GRysySytsLTSV/sLZCT2g7jGbOAZmTJ/gTDAunLXM8FJht3KPkzmFpW
qCR33J5ifL5U5SwFQSx9zoJ5/guvNWOe5MirBLHMYHWZ8oendGo53C0yU4w742Qb
bROB73jTKDvSL6Ncj40bPjzUYRgTPHnyaqBK9GecDHedGB3HP9Eoqch7hTJbtWqt
6vF6245M4DJIjf9uxgYAI4BQEJcp/QuPpUcSPrUPWdSv0nhfY/36SnetLrl4UD6+
z4ja4TdFw3Nr6iyljg4TPL2j/VmJB3dd2Zt2DwJ6t6dFlQIkF0PNlAHZB8HvLtgx
JNyxhAbARENoZ538ic7uvAimFYuwfhLFBpanCwP9mgC4rNVVnwjpxmbu1/YrPNlT
UC3YIzdhz1rBs7VTOTkn6lQb5VqH+S+3zz7lFrLGKvPbfY40nFoLbmFC1SQHKv/1
dbgF9Mw4HXzoLlU45ukR+/aPiGRg1lLIZJxn4QRF6JsD0gxrQMrGpROo6E2CXced
hnojnr6GTK7XqGZSgP2RlUCS0AZYbezTZfe6/6QshaohZ0fPGRYkcEJlckYx7TH+
h9FRLNiq9Fb1CzNsx7xPoXzieILPwlFkqvBN9F/OAabyFiJ97Lrb7V36y1JU+7sT
Fl1h8K3swCB/P7EE8Nad3qftwFiScPdzuTVN1/5t/gtoOiriud8m31+bSoKC5M9i
UYKxrLXvsCEgcoXRAQDJqxqvLqVnn0+DcszJoYgS48yUi+au9DjxJqiQ+Kbl4//N
9RsXnp9v/EFD2XufXkwP3oplnzyu3WKwSTFbe3x0tKLbbz3WzET2eXXDxrumQ/NZ
uaSErTNzQAz1hVe3AEi/7PZke8sz2yXsAsc4jvdrplZK6GaPOIEBFet+2UiYujHH
enUpnMr/RtK9YonBTHX6tvhMkvAwjBvQc37Rzr8Fc69ausvcgL3pT2Ix6zz7z09i
wmgd9mEs6M2Ey0hF8WzR9+Gh/tiR5fWKj8yNEkC/3t4VpLHU/2anc8/d434+0qnK
vwAO0+fh2o+Ifip7/pO662rqCvxFNCfeuZb2smS3UDILM3nRou1/EAr+IA8oOMC8
f+ooRMLrq+D1UJbLSJdbzjpVP42hf2ii3SZKpXdZ8vKKRl0KK0LGXfKKZzh6ILID
m3Zpdqs37hhdwCy1gXNA3TALfkg3u0LoR3OsOMbIwGB3qvi0+zYnqEQ7GkuV9bZ+
9ZV3qyVTPZszuul3N0LE5JlFiixhuivE41psSKz0WPhCRRwOn9/TnQNQHE/WzVbZ
dYA3xg5rkNU42ZU+5S3uQUNd3YvljU+BLPAp8Ti2oCIa0QNQFZx8K8rdnIOTzczr
i8uI0jL2s25s5YQox0nOf45snNguvzIZNJvyhlaY9QlogSM43VaaDdP1qewk0P2v
WdffNmYcpqz8AVQYYzYucuwDcD+Pt5O3WCjnY1cvuHAf1iJbjAKaYfqFyGzzPQCu
2UwKiTndC0jO7L1u2ZMRMoKLMcMA79Ax8XBD9N33m2I6kxth1MiUVDZepntzFoLe
q68fhAu+d4ZMED05zfZWdI0JSIvYayq6ApofLTx9xPdIeHClvB3TXlILNCvZAmuL
VJCwcfCH+1/sYAnHeC0b237RkQYiHTnjsZmQ/+XDk33IkReEEt0LY+DVaN3g8F3r
DYqD8Bf0RTOV9XkhrYjHuLoBLUnagW1uhLx0W2tCDT3tRqW9CLBShyVdFRZ6QOtB
JaAGErwl+k27uVaWfDA37IlO3wW37MTF8Ef83+ZQ1SSzzV5K85CUpnRok3iHYFGv
Y+yGIn2sDyVshiSaOAjLWpvu4LDf28pT8O1vuHzvlemcu3h4Mc9IagvaN3f7hvWb
GoVQUpzq+5biuda6hCUWT7Ap9GZQzitM23ei99lzKwIoQL10iLUHggTg3C2fkgTn
9ozkV2bWC7K+6tAT6q/hTOXURI1vwQA/P80jZ//OQZDdU9tsYxF0Ld0hkyXau/vK
VSQdP8yRqUdkEz+UlqVlpyPwKX8K+0rxg0vdMHErNnWoPTwzCjHeszhNN1L3q7+l
O9H2Etb6+j/urVwqaDSPBo+IqF5BLQENG0+H4XXeQDxrNrMonKGVCTUUs54eNn4l
UVL61j61SZc43uhSUoGG/u4sD1W5vfBWH4KhxrTbPwO7E2DOYS2aDdpeuXQ6FlCl
VMrdc2wnRl+l8yDM1MsHq7GLdTlwlhEmIAjb2JpOmb8ETaEF21Du0ICvCgdUGy8I
/QfYTy2IfQsmLozq6LUcxW8kYOJZYarvmU2rM+zwfPRuerCc1GNANeQMmM2CPOoC
9MR7k6IrnTQm0Eb5FqcXULMGIyS2MAF9FWrXUQ82IjOIsYgNh4FsltD/upVmAKBb
BmJQZGqVYQdvDQyzK9ZwqykQDicivyJpqxyectyFIrGF3NFHCpM7Qsc3EW+bTQbC
FhN72vqIn2o/6f6VdRi+9xRBuIYST+vP9y/1JY4pt89WX5BWXR4/3sqazkCrMWwe
03fjMdDRJ3OeMVeSgAdKGHJhFZssT6U71K5yVQD9UAjyomibTOQSgdqsaYHHH/QQ
tN21WfSXgIDnZUECpbo51dgnarRT06KC3hCKbJBd0QML9uu29fPqbyNGhozTLHEH
uBHtlJ2lDztdxzkv39jAynYkmMWJSbPHz7eIk5UXoRTchm+dZKE2sWENTmyjA/K0
en6r3QB7fNQfawGadnZlxzxoolOpqxZDR1zj44w1WSUUMdFC1t2iBB8pbByvQZp0
7wtdH1XE9yrS0om7xVWgyi7fKASYzKo5hR8KmseG71IzZnLctkVXK9wtEbimyI7f
WrboWzOjaigwRw4ENnmb7FAqQpdu41mGlkrZy6hcyV15UezrpAh8h3EjO1VI1f0v
pTIlkxYFmd3pIr1Ctvn2r+T6ab3oT9vuDqXR4XK0KWxNzYJ/4bCuZT0RIEzM3xB1
0cieNO1h+yAP8hj7xA4ZmIClsfQg/SjL3Y4/CNzzPuU9OpgeUne4u7YSJ1JRdMut
c/9EyjBEnQUBYhKvF0d5sp1RDqIU0VWcLb9/XJ7ikaLF5WRUE7DIrFwnxQpFAUBF
0lB3e1lsfv+bNvGuhiDMuSR/whf+u1Cng8HBRehsOrt2WsdEPf+6gdQJKtAVzIf7
wPedmeF7k11Yvb6XTp9xdssl8bZdokmeno4o7vOFnTQSupMXwY3zxY6Am+ywf0Fe
/2g7sLr41yrh6uNwSBgGleo9iJohTcf+Y/d1Z/SNbosH4lxJxCyQwEK9CvHVneNl
InjdlgdZGcQGPVX5MdLyOMVZl4yJDNobbMLx7RzJrhc879Dr0A7NiCyOSlwhRUGU
K0EpAE1UXLadQfxhKxKVtwZchjO4/2M7mgQQJlzzacATFLPLteJuUP2HEHiHyFCV
UzruVDtB5uoNACliFUrk006U5QUiAc1+3dkmE1pTjYvv+O2cZCERUmeNLA3VEvt7
t+n9gIbxaFgYHwS8FbuwjwPrNu+91fisyjU3tK6x6BRD9G9fp++QmtvFoMd1giWs
ifvwkiymEqhd7SSDtahCmMTRWUdBaQbx8hZezo6aTRxhvdWHob21QJoLyRhhh86z
GWD5ouEtevPQYuIMoMu7tMKYjWFTNmdwdbbj4vh6G2ER4fSro7Kj0q76wEyAmC9T
u5UoSXS6S4bxRpAKiW/wdN+9GJ8eQFdlstO77TPJfhSqAqnm0utxuYfYAG2wAdVo
mMwOZdDSfpB35fMwZBKi5ewFsuzfBMMcsf1p9yfYbrv6I04D7fxxMCRzQPxRuVnV
1xCTVESqEgb3VYZRwSb21tPsqC5+sebRnI6mVOmlDRmWjx6PNrM6bRubK5wRiMwX
sPXu0Md6wq8oCKnAnAunqRush0jAq2oZpH7FYy4JzrwtozfTOOccGvzJ1uvzK8PC
YTdK696T8qxsaKuP1ila0J0CofS9mXrzwJ3y64LVKYz3RsjWVDaEeC//sKNUDFJ8
PtwposcMyUdzzH4qtO0oVDcKjVxtglcZnGNjht2Q7plMHNS2hBZBaatOdgDDF+Pe
rOY+8O6SEhMcFSxNd6JmlyPeopKV7UIjJiCRUjgHSS5LIcHPB+sk9Xn2R/5Xt0X6
+YF977lkO/CPeXI0Oo9SgqAkD+pcj3C1O+WCuEymkiD4pdsd91wdRn58IxGeSPSp
WdcnZGZlo04Io+TCXFWjhnVsfgHeU/W2vWFM2YG8zSQIW6SKDOcC80Az74wTRI8T
elKtv6NRhNUNzmg44RGlmWfO8n4LHn7+FbCtzCU7qQSezuwJYLPgB0WeNGlZqloW
3AZ781kzPSKSQsGTF14u4DZeCmti3ou+HOol43JdxIIA2ORiZPe3gXZRakmEpRU6
rSTQK07iaLOTq0XwV9GcgrRpS8hm5lO1GSLDHqyImm836AzcWbFz2ZEd3JqxnjAW
wvrd4lDukuYR1QXADtripo6dr4HfraixtsROR2vcFb2qNJ+YIkq0ZYmfop/3cwht
ITM6qYdTLTeeSJsEnFmBJUoL489BzXl8haxVQ77piJ23BHJAF89oUXVCf3ZnpIhW
vQ34V5G20BFNxyq7M8u4jBOJ8a8z/lGgO/9KiWTBFHNtsEWkrkaiKiE0P7KKb3lx
03q2WCpUOIpb6N11TezfRQXY7KrMeq6aZLdKMxtARcFx5yEAhBnar4Nl8OSnE8Wh
7vgy4YimP09vZFTqr5wB2nElb3FVBZdc0/2X0orAQ8EN+kzmsJlxzk6q+Ytrdi2y
k59QvwM7VFYCjl3GRiuJMOkU1vGLM/DVAkBbh/DoqXcBOZZaRfEfaz8NrFLozFhN
60OzIhg/wF8e1g7NOQBX71F15/YadXl33ZbI1hxWV0wRgJKgSI0sAES7I23lCyvu
OvFdgEIJwztyy643cu4CxxhmDHpdKkdOx276Q3lPuxBG+RCSvkXj0IhN5ZuwqWxd
521Z4Ocb4T6OW/XjWFwhdiecJgYZdeCs3qD9HXWVJ+lej64v4YAx63ZPH8A7NcjR
pppAyBUKb7fIr29FK7ID9Ju5RZNiSAUaZVjk4mufWISazuTwIPtXJPDBFPN6owgX
eoOkmg+J0bWuEC99PsgPZtlbfo62G/l+ElMjS/goPB9nYbbMh44cKOKyu/WE4m6A
RG/MobiSegSGHX0YgI/p4Y7hVrH1cuPvF1Sj8cuIDwW7pCaW5LBbfhuStfC80pNV
VpokxUZfl1q5alyrYwfhSRLOOCiyaaK3YvHagCEDNvpZDDeoxTHevJcnRHnlaUhw
SYigG8seLa6qO533hNb6ASm8FnAEGmrBS++b25s9+OIlWqjZxcTj6M10ZcwGuOlW
kZYHc3zkc7xP3nTVuoFq7xbcdw9wf2uYeGUpYX/EubmDsVuFJvKsSo+lkVR8LQG6
JkpM6+3QZlk2eMs/kh/8zclmKk81KI8tthbmDS2ompzS1xmeKPGCjO89s+pMdOBg
EIbeAiExfWBwJRmeRzDOqXPh2oZ7J1ep0mc6t/103oiFdoWXoRmE+RIRd5RRM8LN
a3DTdmGV9KDOusyQvKXh1BBTK4T5NBy88q7M76DJaHZSNwivC2BL8g8EtrtTFBEP
20X9LmKLnEq5wZ22JvN1Hd40syO3YyctfIgWzt/DBLXS8L6ScQb4VkTAbgbo49jo
lnkkn30TXsAtnSd16UpqkZwz9M0Lh9FDHa5oot8UxdovLd5D3f6hFwaReIGfWGhV
e5n5068I+1UNiYWpNZnN38MhsRaI9ODNOTm93TTAk4DII3eH7fU9jlarXreZj62h
xk/UxXfLlsNtmC3FFjNY3Bz1/S2QdDYAhNpvjV/GINWh9zrycZQ2h+wgAI3fiDNv
azBPM3Gr+JPCOr412/iSwse5z0oUYarx4fSGCKhgk8v826NSHcNogkXqTunZYZ9t
H8MxM7WvH0K1TXtTyHEjdkXb+waiELHsrrvVpr+b7LmvZQnc6jOA+ZWDKZ6NkZed
Zw4P20C6mdyXCvI8qAhZ8m1/z7t2AHB0BDfKsOgpS92OkmWxV3v46O/w6vO3YhQZ
nAdlkwt0bHv97cY94Uqh3H/ljBuFP+XKRhBrqWFYq0/1SPqxNQ9YjuYeJ9FuSZ/o
q4gb+HRfoXQ5uQ2T/irfGSe4d3D9pFp5moaO7eqFeVOFxtPs92gzFK729g0mtazz
ktG3l/3DlUgAuGGF8rXs1tBKJ7jIdWNefHlZqttm2Y1vVnHHCj9cAK6eLK50ww9Z
9s/r+RawyXy9jAzXcATIL/2s4lwqmFgHwRQWWXnM5VgaZmHTFDZwQVHd6vrwm9PY
Wk/MbVRl9mEpRsFY4gKV6RkzE0CpwDEwlfY3+Ewv/7s4Km42vQYtFqVWQ8j9LSlo
lw9tjy8C+WHx/D6s2ijpd/ayopVMKwSsCRJmLyg/mS8I96jHzw5AvKDZqFGPK2yJ
RM2OpOsG6Yek++r0KQfYLq5z7h96llp1pXbBXPokUv1ViVNG/4wW3GW6gWuT+JHc
AxEQH+Ithnzy+BPZzzML2sOBVc+WV5SGrUXvstMPwaBToQ3KZvNIGv2/xGBJPeNJ
bhcOZK8Gonxr1teZhzzgaNA5bkiqF+SKIVkvj7NqqjoS2dtJ5WNLaZVqMhPPd6xQ
ZM7/bSWLh675l6cdRNkYpTTV+Xlu6zBeBk3S8kb7/tU34lVVbQ7t2mntpepMS8Id
kgHYbYlmIUWZnf2N37BcgjczLS/OZTvhBMt2XKQ1hqXV6F1rDKEYzEMiE+2yG6kr
VRKg+DrN1+k9ANRBA6baRlRKvcmhg3+7EnB6enResUX2T7vMcT/yGK3JuxPd/kTD
rCd1PlcmVq1DrFeIvtGCPqs+hGmbDm7Hic4PxHNXdm5JpE6AVv8hPlyDsWu91p+2
xuqW3On8ZgD8qIqEycnIdRzU+d59P9nSLlYPq4MlVgB9tiXreAHoLADCTRA2uSmm
Wo5foKQCKOJBXtx+bZv/72vPKmDu8nQ7LPXL1QCkq5123igopeWVoPxFrBCcEcKZ
XQvdX2LV52SHTpmAabqHB6uBX6dCvUc0nh/w0/wUZsE8M504hsNTrFPoqLw2bNxw
Xm9i1b6kXmHvLLQwc8Dg4xHudo5Dlin+2OUFV5aVx3j1GCPI4nYJkC64edAEz8WU
0VDBjCMGFsObRQpplRIykI7OgbQqXmkYzymB1g4XWwrYOCqTge45gkXojMwBbvaa
Xi60k9x/vZAB2j9K4vVFjRQ2Aw79gH6C/T+bCGEBTqfE2AltA1Ne72h+h+6VfJYt
XZHwRZi1Wlf4BbqUYk4STbqKAIh5UX/ZEtC8OHLDwHW7iMXs0JKoLzi1LPQ85Umz
KrIi9WIfxN48rTT1LJ1eS0lFVv5ndQKAnuVJWFzQ1yPl561MUvjIlCjITQkedRJj
EpN14YdaYFm0vuq6piQzAtV5lQhSrl0x4Y49R2+wD9YgwP1cUkOo/A7fFz54jeMu
juN+x+7b2F0U6vYhTN5DmXqqUomFkA7Ct901SsUJY5LOBzRwJvc3VqRDXI066Do/
rp+WdcZqOr5hSZQVPifXeU8xAqne+BG4r+wk9t3gHkru/6dlZAhTnAiZODbfOv4I
lvKFDVDHl93OemWl9jBw74Bu93HBI9+G2SbFbmhh3qR4IFWOHjqXXtwA14weGpIl
S85cATFIvCvNLH/8kffm9Rc6hOmAghgDhWYu9cJhHSlbNeS9VDny85B0eR3fyWAv
YpwfCGH1+J9IjA7mM4NM96kCm9rOc+r9MaMu+xCStdYs7RLDadwccvQgkPCv1btk
eyYzFu7A6NsLLqox5t7zn91ytFJ6Ayp5Gdz66fFZi2z+rODNV7NKacb3ELQymWOK
V3p0qXvSzwgHkNGM0eQEm1ONC0CAQh3N1XVwAeCeQsk51V7mJRdNRDaSYJag1kNx
AnhDgd9zHgsJSUIS6INl+9+lpS7B2VcvfLSiHGEa84hG0kwePS6/25yXJzpvpueq
UlkSVTvH+T9yuKAake5aCpTPH2g2lsr+bYXyCjGG26Jk8q7ODqjYy6sFjwcu9wIw
VyTbQCJnf6BxlWJAUY0xcxBL2s+IIixpMZncKmI6o43uG+aVUeRHy8RIvgm5zaNf
+BydwTee5bXX3PJUnoIxdDOtwnhR5/vb0ZYBXp6tz/TxcKUZZRrBRVKBpTE88iOd
wYfUB34LM4ibOUH0BvOatTb5SotlSddLDoy39jny5wV/Fadl36QQrcI7XgFBAMCs
PjaXGeUEJMgeGdBFhMR8plqN3Nnj75LESa4WTJe5xn6NEgAMUvi4XhQatitZaKFw
omunfZCXXblJomR7q2Hev/Req1zMez94UTW3gZ7jKqNUsDruMLzwQXOPzxwR7sd3
Ks57gqlejqCnFTpJu30JSpiCdiHufC8j/KXYGtXQlq+QlBwWN3YnQFgCWwc9HDUa
XHTfToKmd14e5HeHIX75MTfCOsFMWDOcUtdfpH+qVw5AxwD04o7zWWBAvjq+z1Xo
AbZnjQl5k5lZk/VZ8qBCA6HYZ5kEOaR8n/Mc/JWifJ8EU0R2IJVV7floL43lJCb3
C5kf3Ccwi0rRnMn0+J10vnr1COLsNLu1ufnNF9/81zEJ8ky7JNFlNi4+OzTCX78p
qv930HW10eNuVqFF8Hs2ka1yoqF5DcqQV+wPrlNWr3OQKUpt73VOw0sH7X4r95Cs
L1JN93ZEJnSh02Pjs1BXrV+xmzggC6FEg9YsYRv2Mmqqw52glk6peJYG09pMrQav
FkVWqT5i1gU+bg+4J50meWn1KsxWrW5ju0IRYqqRNTmLxZrFsShvDMl13PE1QZtk
I/gM+As07cJUcDb5wmUqjs42XflSGUoh4QZxchoZGAKc/tO6h4nJTeJriKIKrcvn
5dwK9U2fwmRoHkp4WDnhDxgiu5PIpAgqZY+rBzOf/RbOXdj8PurOI0Ip2eBpdI7A
XGZDx2lu9d1K2viiDZp73m7TmER0VaJX2o4RzElZqZQvPDGdxECr7T0AjawI+Xvv
9fdsErF+iCV/io3rECWPiwLOtbYHHDaKPBHF+1swd/9YkxSlBt5SiGG/drzrezy4
LEFzMWm96lrT35gX+0JdbhNncTJhW1OHYUbnTqLISvi2Y8+6hsJ7flncRlh4UsvX
oYjeAiYtzkqILz5zsCrsvKfZdAnDbu22b9QqEQIe8PIgL8fp2wKtRh90d7/OWixI
jX1SikyYntirN3tZYfZruNY87pLEVQGnKKAZu3yzY/xYS0q/0PRHYTGNKX4C+zwK
I906hVYkhCuofQtpcd4AEKI7DgAqIjvYzfgzU3OyqNBapVt5eVjq9G2o85n6WJlN
Bgo2dWB6i6v9C7W1zJox6T1N1IofK3N5B/K0htBE8oEnvFsQhrzX5QVEcscSGwxc
CMax75aOhPz4EPFkAhIEOuJC0y8j/mkGEK4MoXgSR/0qBW+ZoB6BJWGVD9+SM3s4
Wibl3hUlbILRdPJDaR6MvHZUWrOdlSKFK/DDSV6gZ6X10B2vwPFMm28fdm/Pr+mG
M7bs1kTaL7J0Dnnu1a+CbS4QthX1YyMXUWskLHaiHlTcRCV6DF0rLsblgh0drWMZ
CNGt5Bu5hpRrny5buRK0hjMZJbfJA8UvD9UdwtWzqpmlJKrlozBzxRF684WKyWfu
Fze1StHet6Qbh2WG7nE/zXE24V4itLpP3Exbd0aIpHmhbsOC+n1ckgc5CpQI3OiB
wOGT3d5n0Po2AueauuFZJ5J80KMo8WEHJqqrrfGdJWsssSNJUsiSJJ4dt2GWelvk
QCk98RXe2vzt1JkBnNlG62iPs1pZ9dsEQ4ujhgdnskoN3geDjobs5guw0PcypgQQ
QAFsbUq+xEPlhdN1hv9+GLOM4+G3Ciwr63jeDH0Kj0pTHFVFnyiIzWXIxrFvf0hM
Dl58BIskl9bL1ZyD7XFjBX6+RvBLCNyXutUaGyMa36d/EnvA9FB7hEJPXPrxRbvV
TLiCm9ux7qHobV3yYNMikSo1cUhXt3xC0YRwCzsNiRSErLsZkNBLvu482FNvnl8m
1MmzHwTQH3Nf6yqQc6U8RO3kC6997hM0fcLWyCudelhO/Qjl0cMAE4rUUXtIAZmj
bnj34US2V0c16+hiVAS/rYkU6AXqw5G0UWgFsiIo7b1Hpmu2pmyXk+qPkBVfGNlz
MpuyDdiwAUq2wWoNnPkh8lk6tEw/6SqfV+EKjj1EFStPIK80ngJoukk/82xUTpEO
brlbiT9PlA4gjppsISzwimC35DFdNPnOSdZjTvapzwuwaArhfNaqyZcmt+s8go3u
9x0q87kaC1j6pqPoVors3SVvPgjzzyvExqYHSbfdrQLN31/XDMpgSpkMrLER0ZH0
gZFScmqS9yW+vpasxJJ0LlzxgKKz70ee8TFdUGStUD/DCE/VjVEU2Fv11tcyj0fi
uQEfgr5s0JYbaEE2bkA3ON/8Xu3a1v9fXZsMsC1Rd5BqsTVmhIlhiovCXjCoot91
BVnbAwp5FmOYGgV5LiezvON94Tbe8DSypKd9PEkWLkikbOB6s9B0nhbTLvgWKRZX
ZKSslbnqhRLncnmZWAwHNmYwaP+VTmo7EPCiZGhn19476H9Mai++W/wPJymvEv4x
7ZfAf5r/DrU/IoQpaY1da187Hx9rS+I/dtzl0CiQm/G2aur5G/MqrvwROlvm0uf4
9PHLYymOiCZsTPjpsGUpW94LZ12cGnYNQAXuRM3oQa+18EiwcwEZK/4XlURSe3JY
UXNXuZMFPiC/mD8EqwQ5YXay/azOlFFM+NW+Kp9e51T/5qUtsxjItW2nE0zRYY4c
KtR3OgfWsAAsaG4eeI16FkLqG+ARMfSXyrraikb121QomjEOsgz8u3UX+io9yDKw
KpZqxr2KBYM0D5cR7s9pX7ck2UJIw2DcxkCkmtbHSMhh5hNlONcXDw5gaXFl3NuD
8+wVak56PQwQ41zgO9wABOdVMC8Rw9EgWcv1CTneOOXdrpKN++qAMamEgAnJYroj
WTRZjCEQOScWu2h0gIEx8mLqn0kWfOpd+o9q2BsoOj1pLH/Y6dmI0ziEiKr4+VD6
SY9fjV9cJ6qGPO3kxlk7+8qGaumzI91hcrnYxyO8VPlzVV06hOg/XzW28cuO7yvj
Oq4jl2NFI4s/8xO86wCNCFumI0f/PdeIX+pwZ1BFADFiSZSybeWBV3xIZAgKDxTL
LNscO/yBFVf3OG1pIlijWEdIIOLDhliaY70LZCVZgBQH6xr5zHtJBAi3qn83uox7
M02CMmcKcbbUjoFi5umC75XOiSpafmTN3V7cC24uTU8ODopdJVfkdkR5+bc95bgO
FBgjpeKEC09kjyMV0hITcneDSq4Hq0L1fPmumYdorpLrBOmrgLX1Q1WC1zD78cwJ
OxV2AClZfH2KcQC0ul7CYbhNNdQumUNU1XUWWlLGPDN3c8B0In+jlLyAJMUJX5mb
buJKdpDFvwRUDdb6s1sT2yYGvnPah5cnQs92llMTWpKCH7OJIDev9g5DDpGEItzc
U4MdW4EX6dn0t6Q9ILNnoqMDjm8/2fe412TczHWcywoya9GFcYapsQLq8UlMJY0I
xFaBmVF0f7F7sZVxngjhmHrSi2fRHHu5qptrFel3ml5tLxG6vxHgvCoZPjzGoD62
SWbuqUpBwni0I9DX4c7I7xWWQcu74dtWsTFbybi4fO/cZ+hqrUlcaCEsUOu8HZ+E
VbLPAF4rZLmF5nFjRxEH7UBgtsxWwhUMEbQONAJRNUxRdY1g+KHvrPBsrnK9lwDn
rcYsNL6CzNEN8eF1JD2+JrrIyDLwFeQmdpkPm2Z9jGNsNm/BRgBfRrer62tZROFV
BB2LS8KWfi1HPTFHKSlYLD5pTQP7msJi5Pa4Bf6kS1jVRnUDbi1wZQrEA0SeQ1cm
L6rKgkZqdwj1Id5/4al81DWHNoP5Wmj+JXoGnkOSmEt4fFhDyk81DH/rUoqNxsG/
EUE5jgmWuJ4SOc/5GTm4cbqdiAUidMjMxNa4jwozeIKsKDR4w4Z/W/Vv5gt0Tp7j
nAInOFy4fi/vSGUcBNEJrEonm9gDyMivu9DYXtY57rtp26GqfcQ1VRDIzRhBaFdE
9qzN4QpZWlCQnfnir1MDk9uW2E5TlekOXT4dGtOEE0eR++fuuF+P14z34XZ7QlmE
gqN8yf3NiA+6VF2DJtcq628l9d27oqjoouqLJS11UL4QDvwLE7t4SDAYW2cRuuNQ
6gn9MdfnwqaStbCQkuRDinO/KDmampKSUDbNadvqTh79e9+FZcp0DPe3DcKAWoDO
lLrXGCA/StKZDhfuveewPxscVnek+qy8c5X94sh+3qTk+2jeOHaGx5Oquy2oykzv
p7u/q6ug8yEKWd/y7ZA+94eKQG6DIALYnMNM8wZR6nFbrJjCkdtbRSgZdP92iw4M
6IYwHd/hgsmgi2fuH5Ax7Wj164qYPF7nEIho/QOlbzFldQqEI1TQTGGP3UEgj+eP
RfhbnqrCKLiRfTgFOFsv/soRQWJWexohhf42QtfTd5sJYJ9FPifUSaQ/JZ3iXQaS
bS52m8SqyKmTid497bsGASSxGl4bahK+gOpswCBTK22H1oLDWkaPWzxKAD3CEqsG
mzgcbYyr5V3qGAL250V2dTyD1vHJaxcY1V1eMb2KgPi866Ab1rNtIsVPf1oGMB0O
OpPvTgDhe8ngTbAm/XZFHpdp/2yY9/oxqBEKSmxjscGuyglgNb3wxCtNJ3wK5qWy
fOlWnYa4Va9FStvShlpZqzTLMD2Dv9UesoOK5Rz1RJiMGhcMlLSvz9z/1l6B5YMh
czVShdlJnIZ+5p4s1IJDw4iAzyqQ26pDsfUF4LgpuF7Dcd6em70IgxFDDzGimobp
mNk5HyjI84UI+0E+XR64YnnkVKl3+j2S7Zb0K8+3rDpQX7a2SgUCOH5LkXgOofUT
kcdfj5NjWGLSuiUuszwL3S89bzeT20wR+8zgY7en+80KT/pGeqJ2waAAQwIuuwNz
DRnbo4lr2R+0jK/j+Tec9518UszEinrrZIMAWuz7t16rM4G/8cuLtDhEtG/9qO6t
g9hto8yOuHZFR4Ik9qbZheKz72SDvzs7CHl7BsYeypWE0RwB+KwZsy264FUZ7/bX
2OB3ScttTXhK6pA8Vk2Le4ranK3Oq8v0I1LONFOeV0zO1aCXfCFDvz43z9Lx7hIu
KbqlZaXpVv0D2GqKvTRP4wgyFMM7GqyqOsjJRRnqP0BlhqtptZa+JLks/JXNYEMX
XRh/KH3C3xFXY+ojVzsSMTRQQXq8kWXILrjIoPe5RPkOaBpmNYP9gJNX/EHOR7Pq
bdcyYwvkO1mpXaroGzPwBbvPshliXZ6qXy5dJE572SYIsDtlMRV9cT5WEsXXd5nl
LOE6f/JkyTNd19jRwdY3CCXPq3soYkbSnVONUIHshJEyT5j2yaBk35FFttzkME8h
Y8z0iyCE66rf7bQ6pNjhpTUjbn4U8RnVyJnQz4Ni4gTFjS7pn01vP0tvCUMLgmkl
NwI9TJeGbPwsSyz3Fb8ZE8RIVGcphV9XxLlgGV68jRLU5sCUZvwLw9YVmEXUsms1
Bbw1eMCCNFuih9S5trud6dz1gbHNvEI3hOelriflMy/HdxYbhdqiOLIWQR/zCR7M
6AMKoTs+DKuItP34kHJRQNw9AHFcggEZMmPGZ8AzysfuZc5E0N3MfktkX3SH59UE
htu6YrMGIxHG+C6rqGK9rUf8q7/rBP8kVrJIEwwla8WxD+lL3avYLRM2SkceNV7y
OJju6NqwD7hDJ/V4M9crC20zSwcIJi/u1BPvpj41JxgLlx+4Ei6r05ZQwm3sjXkS
J37dKzB3EYQa2mc9L9W/dvdgFvE2k2dRzY69H5VFN5T8N11xreTNTD6H6F6K5PUL
h3lk2jovSFdJHfEHpt0L/vhEvujZm/SC8cHoRMvdh+j21F6Ham5RbWOtgQpdVV7j
TlH78pThfdZi9PBMdnIW7tLyCx/uJTsXa120K/IGLWAMy3F0R8pHHNaLY/fTF696
k5s2LETdhdYIhls8q8hsHBNfB9oH2jR+0XHyvEO85azHI7abFljc5k9hfgUZEm3q
l61uOD4vqErnk9cBi6VoBQl6sezrU22mZfT080EfzohrP9lhStAPtQb6GBNOME2w
ZqrJo6uTvHF3PnRWOEA+LGbubr93k2X9H1zKGJIgzO0qypPDDn8imlhuMwqq/Kn5
if671k+sFqx6e5/x14CZ1RQ1eitXH20ZKg8kYq9tZhTAwEvDb+8pmlgPA/xLSQJA
eL6sxNh+FWKzt5R0AQtOJqJ6oteIa7BukgZSph4FssPl4WX7bpH9s1Pks008g0iX
f+XX8E9gFkmeEPiOiCIf/CxIl50FvEnKInmSXTdy0ptMhLcbCEx+9szamn7R/O/F
E9ZnX120J8Gg5fWzzY/xt1p5i7IDmXONX1N2DV6JR7wOTf668mHl0hmOvHZGsDMz
1Ptr4jWnMpYK7d9VrxfyMDizvOCkflnLGY/4/lQuaXKjcYPY4B9xVizDCG6ijBFN
2CIIMVFzfRY4GV2X8x/zsUv4ua3MmQ8cA6xuPgOE8g7NJElw2mGKZcjXl+xrX5At
+sCi+BKg3vFpQkP0+yLznN9nK05jrxfo8+13Xu2EhiAA9othjUVMzypAoBc4SNf/
Uh8JIFSd3pgGRR1028q4LYP9JdDT8mVIRD952oB+Ofd34tuHdjffcYQdfTvTm/o7
W9Huhix4tMrR753PgRFZP5El+DiQuawMAhr+7haJqVk5j4Ya4kBlOhAkqX7j5Tzn
EVo2JEogkMb8icUr7s6Rny6O0QrbV2l/Q8sUCkxE5yAdU/0V8l0D77Lti/RS5sKy
ThSPcwHL+5XhqbKdn1elqi5lPBfLBU0e3WOBnPT66qS/Vw7+iphJYCHX+n/MWQAw
N9fg4MT3Eui/Iw4BcVP4ixaXJlG9eKet2HdGNa12TFDcr5Gd76tR3G+imHW4PUqG
iDC5FxdUt0OvQvaCR53/zDlaWE9Ch5zrm1UehMaYlohH5Yvy/yt1bizVQORYHoyb
s2XKuJU2Yx0tZrsAilQ1hN65UtdQgY4qltDPXuQCL7u1Ikiv/DjptMqJCRfFi5B5
bfi29op08gkFn6iG0zTFohJGHclqNxrm8kSnT3R07Vht39GuwW8HSPwjI5DiNjPw
EPu2Ox0teVN/gBMR0XtoqlE3YZcOTIHWryq4cGcLGb33F2Rh9eh2XGTfkNFRKMme
tVxXRubfh5+moH4LoLF8EzR84FhGs9JtkcYJoRVBUC8fXXsJq46CbyP/pNdocZHR
c02r2TojnCUthljsOI7uCoTbXYmT2Y8nb+HealFswGN9urtTFzxHge3wPddclSKF
MhA10t98AzTcS9LTu4DBVtkOBLsWF39hZQZoLqJLyz9rdiN932AlmxbdeD22guVW
XMvm3ISXShgjftRTQUrSUEwfUjmRnrPYvHp2vE58lRGe5IxKzxkU619PUWIrDUsc
qWZNcd0mg+fjm/S5u9FMdAtQV7ToN6bE3WbSpP99A6735KH2Isi5d49DaTZVJPse
W32XxBTw6cQhmkecxHW0T5wZ0lLIAZkb2NFm52dEG9Wm26WXaVHzWkrg+OvZ6MrR
HlCsFotuKmYC0qtQnwyP8cIc7aF/5Gykuk11LqA8gaz5ayY1gzX7wWPYe2HdMoiz
BgHGkIbrD06dgJvftJLK7B6Sav25/gf3oirg2/9THF/mDIhFKSPJ5d7dhdroSo/g
HPbAHEmdJpQMNSo/TBWoEawlN0R+6ouSiw0uRuQMzd8gi/MUloPgYICHWUCFnMgW
jmL1+ENoom4CJwo+2hlDlgYU+RpficUIBmdaRmEIFarMWLfeC21wZInxXNoayj9f
Rq/SyxokGQmlXyCUPvPM4XiDsYIcsP8mCeri2G1s1TCGn6k8RmI3+TWSjCcKqDHP
moIOdUk7yIv0Hma5xq1gNGRCD3rxEHkFET3mi9MbLcb20FjY9Ks/eMxbm4TvYDgW
VSwojj5fokM2D03xG6nOeoBX9KdOY/sc8SlLHixVOEsgFomiMS+BNUbiH9ZtZxEA
zoPpI40vBDzyUCBs2xsq0bnZMFIHZH3WQE5NqGSFnoahgsvhpiLpi9BWWr3vNjPj
utLGOTFcvUm1t+ZbaO+/zIpUR0ZDpPmZal2ap95BjD2bTIRUdnWEaygPlKsGK1Ou
S3RGuQVYx5UU0Yb5G2V1Qw2sYYwM2Jm1yyPg122fge7h+FVdsqEp3RMKPcvyt2QQ
fwstCLAB7OB6UunsTRGZsOU8JwZEP3colzqV7yE6SJi3udV4dh/rEU0YiXHM034Z
T1EVSwJf517Jvs6f3M4Wxw4xrfWqUVhp2XBUVKl0Klbe9dd6Ye0S98a9mMJyZiid
rDrWa0id+sO15cc3Cug/pg7QX/zP4mlVvB49U6EFToHDssEcNQpJWKLBDa4AI746
ZSBY9HEcxi8HUibftJnun7QxFmQzW4IKOxXproyxYXc0MPrEOtNhTj5SFNngSA8P
RvpkF7FzzYjcxp5bJqEfwekjH0K/WEu2Y2KiXUPnc7k78PAhnVBQsO8me33Ld3U/
xbPCTUuN221CYDJF7+lVobF3ysNUMrN4bZmaVJAZ0QyewSKTC2o/EYZ+Ak3iiNe0
wP/8iK1E8ixfYqSlTxWb+VzYwy5AJ8dQgUBv6Hn2nK87c8qup75hHKy3zwjQ2H8D
SkHH2+nKL4rvd/zrMxHF4gBi5DPBrbeHOzbJAwIrvV0uMmmW9pXybkRQM9f1FIso
3avbQPraVVIgGsS+q9iRgUpxMeABnWxdfgKJS8+nDnYhOkXFxmbfcoLqic4X3mPg
IciisH2tpH02cHOuzUZDmx2OPQXtSS8n4PrixnEkxRL+kasii7e08Y3Mfqpqgy0y
cd6E+RVaHMqKIRKFD8MTYBrK/TonWG2MBp/SynB1OV7gyyPgn8wgAjiaroaluZIC
+AAH56/y5P14r51p0MTBPKSw+qVDVUcTyGq5Wf2WtIg3DdHF2ofAC5fr86+JyZeU
yfqlffWmboJqPlQppt7q/76QOnF8qGT/BYf4LsTnTyYTi71Jd1pBYtOouijuwkFU
mN+anTABGdHyZnpfa9ECb9dluZ+bIjdR5BT5smfn7gvOiQRFfSOsH7U3pkA9rwL0
HRSIxTzjEfbvoFfnGlk+H6MPzKwelejzags16nxQGkoF/LSTbQ/ddcyq4+SKmNDt
9StR9KIWoRTb+s9Sja0YDStsjG0bEZF85eozVmwcp9xoi7SLRzEW1qpHG96VXPlX
/oA+d/GCbFZu/U5SWvfmQmdwdKpCRbabAnGkewy6VenIATQ1FlarYnV1AvHH+0hX
SKYO7b5JSTlksfsnJ7la2wu2mcqdIUdPHxqzFzGeIE5VqVw1WXJdjFPfi3gQAKeO
rDqQuVDTWfu5WTPuFZ+XodHFiXO7FvbJRdlUPZDnF5+8mj9J3bUnEq4uE4K+C04N
7BzKdCAMo4OoQmGLWV9Ku9gRkZ/UnmDpeUmaZ90P+C5t6/Gi/i9tQnHxXC50tnPz
L8T6ojTwwCh3Jw/wx+r9zvVzKFMNaArpohGGaZzXlTS/4vPzwmUACcSkqyeyeM6w
S35avlWocX7dW09MqQ+IhoDj99lBTmPYDd84TiJsLSYrAdKA+SoaCusGS7K54XzJ
wUvE++JZ+HDVlTQw45qqqUOW864ITjLM5KuprqRRke22rcYZr0M/LcVNUaE7BWMj
V+lBphS+qFyxNRF/14AmfgnDCGAg+tktkFwLLf2AU+ATNAkY8vtiJaWyusrUhGcW
R+6ESKzu7seUWU9239GDyIq+QnL23VbshBwZpAFul1oacaCku5jOBiRaPffSiFWC
72TPpOmJ+2Xn6DHgkAGlSysZ+vAPaV1vf50uIz9Sb9A57Mv3MMIBqywHch/2POiU
AJ5VVMxrufaqdL3nVhSGMFBsVQcder/4x+J4As6MWUZK4itGAneqqVj+HiZNqBSh
mbFAVFP7pn1C+loz+i9IHTUR5f1wxsfcWxO27y5Vp64FyOBYeW4l7u+3OjeWyEAy
0vANsSp7It4q3Td7gP+BvcrAxiCIWUc17NqoKoQ3gf32p82G5RJRXqYxd8Ao34v6
48K8npLhYNFXHAIZhD9KpdiGfYblBKGHTbdsYR9XmypRapfRoHkz1e1mjR8RRGC3
nB4w2VN5++EHVdg2vs2lyKAocXVa7jYsOgxhjGU+tDKmeo46krNtXCX5EwhLXEIa
B9XspUkH0jZ/vzM6P562B44vGgp5cGr1kKkJKt6+OzsxNNX2o/VF6sjOTNroAOKP
FMwtbuvOtx85w4Yo45/te9bEClIUJ11wG7O7r0bHM72Yjzq1Ntk0msn7qjseGF/A
UJuEszLYavjRbQ/UQTMov+j8708LPT7iQGl2NfSLADtLhtlkAKhuNUJ9V2GAZmdV
l1zNWLTO+FGMd6yZyDe2pzViCpZP/cglReL9DhZeAzMNTjKI+/KMk3H2O8mqlO1c
X5EyVlanMJR6JsDAK0Fa3arquKLNnJ3zEwPBQCNUFCBgVwNMX/jncDHvgder/aZw
dZk6bFClNKTTVyzn1m9q7MTs14ANJwS4ykrVZIzmN71cGYbIcgx/AzYOeThbjnkV
WsViMkibJPLGa/CSAVdM8uV+Lb/mJJiF481KwS3Q7co8nVdQ6Fz3cS9Fbvaiz6Ir
smNgZOnuZjbkTY4VHPKa8BwQEitP11zbOzZfYlTdqqitgriwGhy+xRFgER+Ilt5W
G+kiShZ0/Pxnw4O5DgLjfa3zsH0u+z8WV8OpD1uqsr/xdqybwzxakZOiaO6KVJCI
R4jNbUco7z8lPv7Hs1BrJlE+AmTN79fnwUN/EVUu+AXmXtEE0dj1kQsm9BTs8M28
DYjNryE0m+sxFEGZWt7ALXg61ufxlpqgSfz/iW2rYCrh1zamrG/icgbvAi7ZXB0E
CVoge2tLPJHrhm0Na2CqJpIVCnYts0DoHmXGG0C9d/i/dDmqlZQjVDQHr/Pe6wXo
s7cTQWOXUR8xzXmMnO1ecSfCAoRaNXRqGLLXDtGC6i07/wwciUCtyxe4bltdK6g1
kFco4yK9nhFkILyc0J6f3tLcrh7/Lzkj8Gu22sa43DpHtwvCclCQcQDaB6AP1ZRV
GRPbFQYhrMcn/ijRlIKFks5w0CZ4Q6Ru6i8T3g6EUbWK2cfAoXfX495D8SBOxfN8
+QWPXEojDqPcBvPtHtZlSE4/fj9MMVmtNxfKB5D6L/GmhFQ/zJ+myiNJZI/YV5xv
jRL6acWPYoZ+xTgMbZcRLjaNGPJI7NIWIuMZeYtrZ42qMjW4o5XrAxM1yGWdOrc+
TXKANKdpvpLV1rHlQCM3FwUN/zShRLLFvQMNGccDn5jR4bvdvgUSI3/tThlYlFaH
Nyv/32WkvnGuRwmvYpdGn4wSYu52116/TLMMPKFJUu9BaIwRnqpplCV4djhTp1Kd
Q66v+9yIDRLNurkbk1Z4KTRwk+dPe5sNV6dqEgbONt07boSaDqLBk4OOCeSZ1rnI
2ZUhdCxM6jIP8BGWqwyLLqiEwFB87rjzcinndHoBH1QeSyYeJ1QwkJ7x0W9TpL/b
uQVcLcV4AMsjzKJKf8xVJwq270lDqghRQfFg6zhaTyuSIrFyXbv21zwe7NJ/93dZ
aqjCpxCVsWgadOCEO79ijTVo+WtboIcZOHQAutOM3NoL9VXhn235EF/NY6hLVxjF
P4wsl0YF3UPPF24SegJly6gGq6/F1o9qOgfjw9o5uOGQmkZhviqwIKL+pGD3MRnK
Jw42t+BXSngwiKfH/17DpTRooT0IiDWNlwPgrOfQJmFu67j6S5uE/vN0X0TzEqJl
r0b8+VHJYzK7Mpro6Ytp25uicAgH+8WbMJ45qZA1cE1i+C0QL4wRQcZqDQBdfi16
kkDwGdB73a5vz55A07kVyh/8S2ITxJN8JEVQZ8PaIks0Xh+n7Lve70IOREM215kg
0YT6ArvfJXvqEeQ0HuxFddcibFn1DnhHylqcz1Kdsi49BfSCe/WyEsvYgXY+aH2B
zFLH4mzLLFmu1/kcn2sUzFhmqRRmfm0OGNLhoVkzod1xTPpPd6pOXkS2872uxt64
Z9VALpzSkydAMSoOIRmAAOfA5yWmKuR8wBm5MPhhazb9V28ViwaGmIZZgdcMDb/i
79eEka8Urlq5a1FFeIGKgjUEp8q7OZQIjxlAYeP2gwFRsOXq5C6REmfA9hJn4hzM
v714oF2ZhUdheOD9uzZf0tXltXBDUIPWN9eRWtDQ4h5bsL2B7Bx8+h2lpQPN72FO
HQxZiV29Z0+uBLlzTdVvpf2xcL2wPg7rJkpkMl2n+B+M+Z1Jz1vc3e3ImVLVbg9i
wY0IhGN/YUexuuMrhI1rySXq4ycD5FNbfsdUYO86FNsKNkvAKmKotOjmlkUv1zef
A6l3iRAQ6yJ1dQQBu30dECvcy5OUzTs+2IChjId45MpWMJTGHYN44gzlwXU/V494
5+h8VtHmEkrJgxS7/X+W9yQ56hNfTu8Sq8SUDJoPLDnODo34RzuuJ70dhlF2kDrt
YGoaGqcEvDqSxHaJgSZkm1P/nB9rdwZFTLFSgdNqKr2ePgvoiOv6FtbdFasnDZXJ
Gsz032AAbnxwQ7YsaRwVpn1NcuZ3sX7MQpOiGphtC6J2iFOP/ysbTpn/kB2ETHz4
xvMxrq75S+zgxvQPr267VDb/D2bENXh9XE7CrkRj1kqLXwF1+7eemXS2JXXoqs7Z
vZ8soxRAuY+QXhnvM6f7dGMuQJu0AqKdo74jMrMb3k6ibKOxE5avzV77Da75M4dL
wiXAtliswxenaybP1eeu27HNo33NEYWsUNkl6dDcZUaf3v37M722/9hUkrI1bY4b
hnuJZ75tAbv6Bt2QzhXlcISOi3vl5nZBpr7NWfcVB7tNAnqfCOCEIG8Q47DU8pPn
MuyuPTy29jnughxyMfgjKSmTnkjly/ZIYB7tBO93LBpWfpMem7xqdl0OcJr4Pk+/
Q0c9135IBW+9PcotZC7vbKiZQXnh5+obew7XxdetrB1p3kWY8btjh2YGSt6JtpTN
aYjDBh4lV7w8oalzRhA1ExEP8Cz0uY0sYoGj8xXPwurR9zu77QAXNO2YrI+uRtik
S2b5Av1F2so0vASU+pk+4lNZrUaxHj00tcUMKoNLkUnd6y03Z9q06RGf7cB3dmcy
uyiM0z6DgID9mT6hvoxpHAAiZjzscfDF52gopjau7VGJx+HVVVZTEgEEkemCtgNr
Z5jtldywWeNBt1ND54flwBf6rZOsWP63A1nDbO0uUrVwtvS/c+62usJ8Z4Xvib4J
MRx++ld/9VhKQ4CUTjtFhLLR4AvdMGjrv2YGe7fqgkhHyNJ/Un2t0nfwO94tyIZz
y6RP/v+o3zYyYLbqnJvp/0we5+W4yvzeQRyHM2mBU2b5CCnWnhnDca62r+k7VI9f
wpI7CV7w94WG4DjAyXxqiGiOSt2Vk/sCllt6LaSJJyw75L0W3UcV95I5SfQJ1YWd
m7tsSWWo28S1ZZJ7Uec2eJp2FdfX0le+P99bXDgFiU5tsrbN/2qtKoeaknRaBRiR
PhSolz/Adzwv3UQM5VUzguSpokKyZO96eqb73FKhrALFKywVKcEzWumrSq0/OWWn
b+ftgmNatxb+RF0/QkQed11FOK1tNZfLZybwUleEYRHzX+9qckSZ58ELjtQzky3o
AhDiEryuOe8lHYME3AM8NgQLuzqOvpO87ARWlHwawPKOa4ETxEo+J6PrhykC4pTG
z9MSKN4Y0LzYHU/NPmYK4AqYYfm+D6s3E9mDzs3bprO5zodbFWuxbJkkkGiIyyb6
1TCVpLWkg4aYFsYEz37+BxwGR0XW4wTHEXTCBQiIRO4tkPLtm4X6diqIYLx+Bzm1
GrEq4FidHYzVXvsKrVQk226NomvAeiwbO2Ev8jMxHkmV+5JaPMmXpOArvnbvJaE+
upAC86Ge6SJ+h1uH+5hk/SAE2t1Qa0cAF42nxbP1OW7u9sqw+Zp8vKeAbLaDQfJ3
9pgBdB9qQM6eQzwTNTURvnlIIAC0iyrkTkq/y9nEndwZujyxsFaWVNUqWSNJqZnl
WiX7EU6CnsF9K6R9cygGtyeQFgJwcYEUeasH59sRMhzpFDV8iieiKn39wNkhMpOw
MKHRYa7GiGGXgq7zVYxfNAxyoQywK1mbdleeavCX0oAYYqsUysPfrY5W3uUftfcs
BNICH6pW1g8vjlJopoY65dMhgKmfdFEdwUrsR46ErhNLGQ3oDotM6cJhzjcGcMsc
9CnrufpWDnMUXG93HDNPIWry6fiYLyt0GorZ3wJKmZoghYflITz/dITvGUB9N1zK
oOnd7znbs685ksu8aD0WRnUgTOdktPNnW9OwfZQ+Qh1ZhDz7dCYaGHD3aGjx5PJH
ZPCvRu2g4fC6Apqvb69Wnli8WPv2ra92SdvX+QYpWD3G/zmwIUxWRDYCX3cTPn6e
6/y4uvG3VRwp8dOhtxuathXfkEwjyAvboF9rkF/fH+V8+lrYKI3vQtHzxwdHmXRY
JHvMvTmcswAgEYjSSLDkvL4Ga2OzUecwvgkKc0UUSbxrlyKgAYRjV6Ei6w68UDN5
cDFWNGYThxd1OnEXCvaaAXMj9u/TR9FD+sSQeFD7/OOzVH74MQdVd90XdWumgH74
kfHyQX0UauGYkExalHucJS0+yq3VfEDaCGRiMCHHNPGMNm9oXtlPnOqwEl0uLyy3
5jaFW5lAZR3xVyNJKkkL3DCJH6po66oaLJ9gTkIGAlIfGA7+nnhv90Z0H6AsAF2o
xMqzNIE9RRF9079+N2oWkOnrmTps3DlkimoKU6Qu403+7crWH10v+Mrx2TO+ZVxp
uaW+3mCkwnaRcTT8OY95IJBgxdS185BUpcdyMBghE1gOkA5ePSVXD9utREYg59sW
qqxWAxsSdGJanE362C3mg2j/wLumV0XDHhGpdTSZswctYeAmqVDh5smko4OcqVRg
UoGzp2IPhNfhwiN5QRY7sIQacIPkwFjh292efJu9CktW8XgbcE1UKpU+q51OxCJ8
uPEcd9QQnP6zyb3mTChhG6lFKOo2M26wLOICQyEQXGkP/HAYP0ouofVtyVuLqKk9
6AS578ch8oz9v6jO8JA0jTuQ2pp76wp1qr1IGHoe1yq4yccTG4Quklo/fsco0m/P
QKRiLoytd5Cse16N4o6/cFSs1hOb/foNTIlrkOAq/CFtajE6nPELUSwDFB5xdmcx
qpliNetifB9ZJnOH7T80kNpaebMbnY0U6EuW5WQdKovlw3kku/bJVQZUudW2qcMi
J4Kh8xmlIVH0GMoh+f1tyy4qBZkYxe2hG5pZxgXmtYjeDWPD+NOhqC89ALzuJ3U7
22t3lsyqaFmtrIl59Mx4xPqR2TK43zelPuY2Vv4wf7gE8s8uq3b4eYwYtUXQ4hpi
yD7EPi6kg07WdRcYwiVaUR+aixRbye5MyVYDffVirGD0zONKnHGWqgxPWZNZiUhc
oi3vPQHJrivDFqQ9TbBbb82dC16+SUHUqu9CSlOJ489OIw6/y6Su+61XLQp/D+ug
BHXnamgAX/64BteIVk9RFEk5fuy5mCfXgPhAvUCWXlVu23r6JWFeetu4qF2yybHL
Sw5vk38LPVNcCeH1hm3AWuG/ONhlkWT2K62ZEejiiCdlZblBRBWxYMPTXd4t6mBy
nsKkOpSun3JEJim8jYwfqWEkRS2D/8QwUKAZ8nrdgpsCuXsh+0ULRa7AnBjlszWF
wBDfRg5l7wr3CPNFeUAArRQ8SxTAp+8+dpmWVqoUsZ8UZUlhYRXkmxST37Yxq3fB
5PRRzp2Kg0wmpqFjzEBmwVnfJ0iEjG+d1AuFvQW3tj7im5cWUvFttYJ8yp+UtK+Y
QIpb8tw3G+Y7po+m7YbwelBYERRYX2mbrc3ilw5tW57ekgkcwacr66vMMgjT+l/O
OWk24Zr+B6C6hWO1ipJVglBALeB5o2rH6hrj5BZBIgAdVnBPFBVNuqDXcCodRlTp
Jtr7ViTcpAjW7pffkInN9fyNGy5yTDD+Wk5gFeT6Tu/wF9jD2HP1DKAMtZJvJMXP
5JIgLZ1Sfnm0wNz5cBX5HmCm4Vxh9x3nU4wm3Jnrzk2367wXeXPmCqx5pP5Hb4sx
9IlmrfYUSTKl+YgMFXUBGJCeWgfshw2Ip5+fxAQuaz+5vyD3CO6jlizGsNhoJAra
LBMaNfu2WrlLZusPZpr5ZKTFU6dlYGsT3zNwxlETYpTmae6su9O3sOtZwMScZCAc
MX/NlhspKs4CtJIsguXZpLX0r5v8L75WUcjz6+vXd+i4HQkMCssLpBlWIs1WeWYU
uTll8lC2C85sTYqDC2IkBc/eqxy67iZFGsBqiay0JYohwvORYGp/M3nRl2oO98MH
EcsuQyiUQSzu+KTnXuSMNOZcJSDLTB5HCDxVWqbyJ6utzdnPjiOW38Tm/ULvEzhA
5SpffU4IeBHta2WwlqNqmnmfVTk63XGS7WXCPfGHuYLPzV9zVvQNbNpTK2m3lPAO
N/Pa23dw7HqhJTuik00gIOz4kPtpLxGPLcR9OYZThHCGRxF+TxTFP+kSSZsai29n
KnGo5M+pxdJxgb4xZ+YSqBMpV6hPqnRRtMxm6hsT8WR0Q66sQhL9YaF+pkaSoVk4
F6E92z7VxUAr2Rjk09cxFDEU5yj6ugR5eufhbfVIWmkx6Mk2iIxxoplEv0Vos78Z
iaLFSxf5WkQSpVcMalgsbA6LuMrsCsAGKapbo2WxNgviddxi8i+9SJn4g9I/a9S7
N6VTKzYAUJGatiyFt1M/iy6uKoM9TSRuqihFeqdaFRHPO/h0ZpcS3lLx66E58x6X
ZYtWjN5TwxFhNPG1M4x9VkVymZjGLvP5G8kXW4mxNcRqAyQCRpjxHr80US1j4WH/
zeYwRjLcxVk5Faud57c+/lbvCuFgcDqcSIEjoS4uzleUd9Fee5iTsjMMUKyCNdP0
lY0e6UiWoamoR2QseFpKBiovlAB9RILWmh5QQPXNJkXHn2r9lypt3/GYRGDDlL9N
w6G7L9mck21jkOQyNFMxpEiByVtNkhosay4jruLUlRCYkFVlS8PVcJtBGY27zWDw
6aN96stpMCAeNBh3qNwHqZLLFs+fXFllsJFmaHHU2yL6tKxb0VjafDmPcmOSWDXF
cXVtwOjWayOPsTfd3VkMUX0Yk09dXxanHfr1BxoXyQ0pezOsR3HKugU6NY7fSVl3
aK4gTxgMQpBY/JtpikPMvg+FtzZW7PDcn9ToIfVYvtLc8urZSLXt+gIyTHvXDRqR
rGCbgt0eeBVLZ0u/AtPs3HyyYMRuulVlWaIABOdJkUACageSPWP8cEyiKH0qA97x
uCMMaegUIzEFJpiiZY8d1eMnozN/4mUpDk3qVb6BJPotS+Zu/DgN0eHAEejEwlLy
scwZFgVx84hRkPmAOhjhaAaYLTt1tA5VtepMZ68OzKjdL/FsQ2lljQeTPyxvOkAj
N1V4BQComQgIE1xW1NWpb9pm5ho8Znx+Zb3fLONHHtiX/a1TnnNaKRyeuzaD8RnI
pRj7Pyl0NbTVNQCULBbeCUOQWbRf8CGOwRvwLcEJgyHIiDfJov3rm3H0QWqFH6y5
3vW1PeQnMzGMdabgRB5FofZhTnDA9dmGTHtpZM6vIu5Q1xTK7d5XhSp51WA1LEjE
issUtVG7RpasYGgnOx6wVW2m9JeR/gbJb9k2XiIEycUpy/jaTNtCGkqkU5qGVlkZ
B2W7MSM6YZYA1nA/K3IwtWb9UiUIolLrC4sv4BDhuKmQRb1pMLHdNrXU0amp+TS2
VuSMu5nElhXe+SbEBYuwSX2a378fZaUUeRe3s45ABgcdA+H6XgKcwd/HPs0Vxr7R
kWEB9wgc9YGOpHMMH/4crc9Z2pjJ36erG8CwvLUA7JlAOcBUJPJbLCRyprsglSJr
finVy6cAF0OWz+XgtLrVLt2E6dIsYQVESfbi3NHDfji+v5pQC45s3rRh4P2E025O
aC7hIIv8kpsXNsLwiIEIOTypHfN2U9Uh52xOUMKKEqApOroCxUx1ya/mZc4cc+FK
fbZcarDmI6MetVev3C5iSb1nX9IuCxkcMieXM3CqbNq99o9Fy9Qan1JHLxbXDCYO
KdMtZNJY/AGr5guU6g8gA5W4ZUZfCBgxMirmwetxEJm3WcCfYk+OJyIhM0H41c32
6If3Ziw/OhQa72coFriIY36mrXSuGDXH1HhYrieTx4Z66YJkKXDv34fIz12Vb6CI
m1DTwxzveLhrBTBq4VMjztIp3ybG7Q6zzbuLynSKjw8Hrxos/rfsEA83bjgmiVO6
zfdRGbmHc405m7hnjpppH+NZdf12Z2X/m2fQsqBnIUH9tVu0PypsFfltMFYMF/1I
doLe8M1IAv93+5eucFNcf+QjBwVqqE90GOGNe4YJY8Bgx5yLQmQ0fHmg3W4gU3Wf
6/5cnLhGaf8PoJF65eUkygLP2QddCfpu2eXi0lBqISXjAo++9tZ9/mWIsMZ9S6eA
yvYNLrBSKAwbW2ZmHlMYOHm3Ima9Sd5nXCYeqcqKlgy9pOkH0sWrVXqS7yTRR91g
BVc8RQJlk14CJ6Kh0P4l9gm+MheqpsV0YVQmAaWyfKIgNP+LGB5Jdx21XoSUWu3p
nV950H8J2fu0cMPxmxpSfp/6YBcwdLS+uUUPWXHZwGeKVIEzAuFpQG8Qy9FDXY16
i4THnBqoh6n1QhDRXjgjUq/Qjto5oYF4cqN33ifhPtvTS8+gPjcVVbeNvqauOT1m
wNd3LSyjBtM1te5dswPZKX42hVn7idu8vA34Dp4VnhYeE1sMwDD9n5k3U7xSTuW5
w7fkZym9BTpVX1pXo4Qf0vyUAqp5ca75YTevfj770tMvBCQHAFYkJJ4Lc8M3JCBw
PERR/nNtyBtqs9bV6nPgBm4DU6mGPnXYpxaizu2j6o2awx1zhub2Yx2weS1s+clH
L2Xbk+NQLK1ugRM/7lD/BKxklTgr51BAOQJhEvtAOhPIgLMzFMsouu48wZ+maJVR
+TpR9RAFxr7oXqe9PhrgL3z3NeNpyoyXfT+2zEBTGev2L0wPBhpieIXwoqAzknUr
XwYQCNzR+HdkLT0rogSslgafC1KJE6LHFSyjgzGsFOEBCp7YtnkDGhIpV92HUUwb
ylY8Loa1Yl1VcvuBWpInHsS+22szSsX77p7F376ExUo2qkJNnST8yukDRvnXMAdt
FDAi7XNddHNOwAWiryRO5NeZLNBahDCkRew/A5u+fM8IKssRxKYzWM6UmnYl9IMO
jTdbiq1aYS1+WJGNccanH8UVlwCamoZ7Ur9H+jjIq44nJl/cae2gTNyTaKeZe6du
uW798iJeexm/Cl85u/hTW77uQcX3HjK4swhrXpDZy+8VMN0fpY82hEFwc78jQqEv
cg0UKk2UBiHza6dChuoyJpkgnnHYXVGgONcqBIfmD5V5mUinZrCOCwkqtVrKkbPq
cMHo0v9MvPjjpk0KDm5ED3/07PBXfY7ml/eeHCnJL6pplGD3lnP1hgLcL1mvYNx+
ofXUOD0oNr7I424VhS4VWh2LTpYtuykV5v7DVhISItH/YHbyOK2+CSM7BHjwV8YF
6/eUYrguOgC1J5Dn6teMZ/J0ACqKC/xsN/+v6g36hGy9yItADUW4ME81xp9flB7S
A8QfvjiH5wsShAbFikN62pgmOqYe0DCjtRMGTZIJyXwB90vifBNBjucP+uTQmPhd
4Tul6GiaRmfkqLbJXyo48swWpMPUS6UKuyTuFrPkXNd+QkCylxu/vk5/cBTNdq+c
u7vdCuK6uSPraTq6Z40raY+ioAyc388RLjkd23DaB+8Jlo4VpoTWWsG4tsWJ9ntE
XvdUAQSgPXQ8nVwC1AMjCe3sgNK0liILR/TBISW9INGD7jwVK0bAdKUBebmVJbic
HwhtiDpL50c6lf4kKdRSpyrE20lD+Fk45YXxauSkZOhv9/22eiYfW5lDV2kIHhVA
FNZ8ma2k4qL84xX11FaUj16l/99vsilM9CC98jUubswnKP/Ro7PQOXIz3KcXaqXk
PAACcb8QtGskq4n4+hVq4NT9qBLJKJZoFb2prcBu1KFyzzwZe1UGzcBj0ss1j4S0
QvguZI3+qvlRz6gNvyIoRMDY4aC/6fMAZtkBzOGHFRlPSAtao8uztU/U5ZbeRKPI
NBVG96LIRS62H28fuRZnJd0fe00753BiEbJAJjuOSm+2gSnnqE+eZygMvCyG4IiG
ClPTvWcpXGM6kGWU/Wa5O5iuDvawrd56RtWB5KLiE9FuC5TjIUE0oZlMQ8TeGtAc
HpvHNNF07Nlrs8gv+8yb8wNUSeUs/QtveGTTC8xTEUnU9mCZDWqXo3IsFWG5RviS
zzPvVkfT3MQZZEZwgiDKdQcPswk1GLuri6uOymuh5qhenm7944dMs6VmW4rfj4Ha
okGYKldo7UP/13oR2Gi8vXiE/QwVbGORqA1Mx5wj9EPu/3JWILQs6g0w4domktem
69JXgPCdZ9gRvXb9h9fbYF7tSLeuXhNRCGfzHw3qgEKhGqVrJfdvpWrcK5snFmX/
H+V7KWorl4jNuneizf5QqrNhnCOMRp2jZHye/CogankXjO2xgWRo88YSNAtZvWQN
yfFV+aGSX+6uk+mZlYd2rHPyba9/zEKulrWxWoiZpPomoWXW2Djkn9kUQYjvZMix
HI7utpU2DTiLrL6IKHvTbWvbVeY8o/AN3BqBZSFPOZ1Ngcd8FJQBvmRcvnbjHGME
tPweuGWmiF2mUiFqcOxBeDBnnPLJOUdRKbS/7eB1RpnOnJCixHdXTgMtc6S3E6kT
w5ormLE44bB7EXUxHN7u2yab6D6i63DwwQGM1dNrBkEupuH5QeH71ClF8DENJUeE
c0ZYGaAzSdNjv2SBXtQfSSoAnG/PbFxsYgW1LUFATPcHVJBxWSbN6V5wkvam1jQO
Hl2ZEM4ZTSW9x6XOtEqZ7CtPqTceA5sEEWS6nspVzwdtsm4MuV7uFwaV5mnXcyTA
DEJiX9ZOpbOBJyDWIcEES7Gx4hUxvPENoft7Pq9APSkvtiLhcIusqNq6P6bruA8k
75UDqX2G2sYY8VEU737yMsl3Kr9aISZPEOFrvbZJUfw9wefPHK5Ul5sbQXb9pphK
yobJrq1mdvVaCiLDT2fpsgjpHUNFtOcGf3pasonX9Wk5/vB+MFYKWzQghVydcxFL
lYKzHzmUoWHfKQtPvl8fBj/RB7UlXzVEXj+k+eQ/+I1I4x4/RAGAu3OE/hPU1t9B
2mTRW4TDob0N8v6JRSEa+Hfkobs5qIOJA/dxGs5QBcAPs25tpbvpaJxs+TfW7892
zDjisKF54TraC8aIXbEVkcLRLWYSRNoCol/WgruZXfumK3QNKZwPNBtTiPPPzv/L
dMQXC1oM03N+G3f6lFMpykSAb3CGCzuqSOJILY/0ukBDTUC3FviIIiGxOg/rZlex
ddisJP6bU8BWy/7Lf2fqvJuQ+ZhCJqrypR6c483/u0pa7NxKpr7Mcx6/Sm+kfUF/
Jlk4wSWBWvJgMEtwT+zlvuMiEzeKhsbKxWmLBpdaUv2lsyL7yFrSRuVr1KtcH3LC
A4fQOee6JSeI6xd36JTRf92vOZQywwOs/RNlcYRVXji7xvJAz5oIC9x7RCDxrXrz
o/QyWaH6j+cgTirNHTRHKWPrHczeITMWEhEepXLq18gmVNDYP1vuR60g7NTCit4e
6qOkGlGXJkgKlNDeds17QHNFTMX7oJ6DViTSaVdZzuEuYA1uIVIOEIidJaW7Hung
PGrEbhIQvrNYKVxrW3uiHrGaY4HqwLJ9hVZxgpeRSVUK1Tf7azEYHs6trFwHqwzM
7vJe7TvryYa+N0O24cTr5W1y41o2jD+7HbvCjpc9hXB6PpJCaDNbTdJjkbL1Ir8e
b0316Z/gqOM92LWlb9xL5hSX4nUCP3srzyJ9WiIZIBDEdW8av6j4s3766RjYmU7K
N9fa3R13kCwf0sTlXHT9tNshXJmoPRn6G0OlPTIMbYeBCCIzVGfMQFQeRnI1dXhv
my66uqKUxeHsFM/7pmtM52KkaO3dSUAjo+DA9QXL8ZblAGdRmabTkf8X6XsRh1Wd
ozuVCWMLyEpKwKJJj9+1kjE9nukpJ7FInbRRCJ638Vu7KNkitDlm7a54WXV3rB95
vLSlqHxbbSDbZvPmdiE8ewV5hKu6Gkep3HRH3iBsKJunPBBFpdZEgGEhcA/khy51
f/x8Wjf2zuS/Xp3cEjZ7xeu9oyYK2ELfP7y6UxIsC6HRFYY585NDdB3y6iqpnQEl
17pK5LxHz+YCh/iZ8HJQlbzDwfeScsKBEVuZBzoMifTw7uBV+rmDRXZhbGsye7yS
X5gJxw72eChLTEhme0BtqQ86uRgfsJHlRxg/Y9P4J2jyTqIq9GbKqGELIH1t/T+n
87zlanuR8pbLBEBPkhKlrOC304pgcPrGT6QoVFSMlY3VUgoIV1XC7F8HEkSV5kmZ
iT1OuEIpH1txV5ZkcfBDkp2zDXSE2ZGMzhrHsY75dmsiIRrOBpjyKwX0zT8KEnY/
M785Ow6giWVdqJgjh8NUXne6KCtCb6tWQbrBivy0bzuLwQ8iXa2QiHjPA16fkmcx
Xs5nehmwT6kApC+SqJJSB36DHuz28GHhgH/kEfaihRfGvyJqm4X5rcp9aSIHpRZW
hfIqV/06i4fZ8FdZ0MjHsdyEZE5syZcrCSKrDeTAIOueejndwkNuaANqXymbm2Za
F04cpAYCvAWT9nG6I5FUPQC3E5Cv4/AfWlUOGe83AtKC2aR7P32XD3O5n9CbTIWh
bfWyKDmm8hoXWFJYKJpCku0P99FxPHHS4wSoBy3mgshZvVPSU4z3FtAUkFHimexp
EtGojY19E1/LQTbdLKV3ttXank9PKbhA2iDEbzvc7zAAiRuNEZQcC/Q8XSJwaSOq
22OEqYX/LaKLCsVg6iLSXlnLXLdGx0+m+jusmxTx9n0nJya3BIY5u9aNWRblgQ6q
cbyN2hmOd1YFGbDGSVn2c35AE2DC6gjHxVjk9Rs4OAWQuUlpTTtJKxT2+vG0hKoN
jHYv+67nmuYBrVFiMtwWCMHi4ZvCEKZlj1tl4Se7YfHWL5njJ23bQDYHCt1dMHZR
yJZjsMCttnKYTzn/3OF2EbMypmpMXErALK5QIRtebHbgLG39YKdtT3ULP6aF1vh2
YN4MZ8KFnCGzqVHnvJRwHrZS3KDwBVLvO0ovsEkSRdn55FSRwwhBhUtUnmw5+B+T
vM1DsC4kHXodmOg1BiV3C+QhQKofesiDm8Tb1EBTGR77ZFLrVzGCcaPrlzsBdRvA
csJkpX5noctk/iPw1nb0P/Hj3bU2w+Pp4t/UgblxSAaKNiliw1bDhYGd5yNEMyxS
O3s56doBNOdWgSxAUaLSHRhg2TzSzJx1SHOpib2uDO7Of5UnkijU81g78LME1/xQ
iBzqV1L/93agjIsp5rHYVhs6Vf9CDKmfHl6AACKUsXwk8L20WPeCmHonoYcPQMei
B9aR3H55nfFW9u/npn1gI26Q1q6/mmWcJE1ULF+Dx2Z2OXW/57FejNc6g0sgYlL8
lPHSOzbZ/xzbCI8n9elGJJuTuBZGyxbFop6jIgVnc5pDwThcASi1zJZ0XaaWlLv/
0f426v09eyaoDZQ+zOe0yOOHHzcnu0lEEkBUnyBZSscnC9trXgmGJI8gNivllPbk
6ydrQGznqOylE5c5hWLshucGgcOcIb5jHSKzYz7QkUiWIGZP0CeeVU9gq0IslbNc
qug2jsHeFB7gbUvgAlGokCP869dpPS3wU8Nvw8s2uhlOPqb+CiVhIxbQ6Aaz+jF8
Hf1hEfKvYJyLsglKjsf2FKhgaI1MDTf6GZem8CLNNmtPURJPjO4nT1mt/3RiXpKl
08z1gmOUA3f184j4cDpKsdYWPKfJGniZYfHIRfzrPDGFVvMnfiFulRK/xg9LJ4Ws
7LS6L+J7plbNOhEMfrU3w6L4I58GSs/H3ciWyf8jJa6R6PVUc63d0EhNKk5IexX4
hIWXHylFHd+F36pYki3YnLLEWJ9Qou1+rtpfY/CZ/L/ss0JHGFUdy/J732TL7n1L
RnPwLq7OwAFR6SRFjxn+0aguaVp/8kYrfOx6lafWC9VrxoxaASi6UMQpnxLfMnFY
IZWaUPP574YYTsD32PX4PNTzV9mx59hJJMwQcXyO0yVIsc0wII6JkS1MlsppIp5L
ceDdGwRaoZMRrODcAvinm8BxSXMLsH6uI57fIoHGcRHa00etxicy3pTyKM60tgd6
hVHPPTXrF13nXw3JPFcYunQaozSzK04WiBHcbGWQeQs6bXQ4vExySAUYP9VuqJVF
ev3C5EXaiI/wfiZnQ/enlsRi3ig7Ex0en8KIykK7KOrHtIJZv1FH4eZJaX+i0ZCJ
Y1NHMVcITKohe405LQjzlfZ7wqk18ZjARoV5rAaAkf2EqU6P5oS3xRYEBf8HM/rN
M8mwpk9E2BUsrIfWNZcVP661WT1vIL+AbTXEXMn8xbvihHWkDbLwjARUS8ENCwBg
Pa4zjpWC7aPG6oKq8TyIX3SFBNv+XNnmBulWXpJSNKQym2s1Kq8g2nTXN37Kceug
72eC2danfOVr/WlOQrpNzf8PV3uZY3wR1ABRsQ6S9XvFYQtmSuIAH0H1OFdlpo59
/iEHIRG6+7rJMxGjv3iO1obwg4n2HQ8Y37j9zWwAQxixUOPNM60yDEfYD9h0YCmi
XGqLFXIfmsBANl8vh3+O6awm6AgVx73hWOnABTXBhegW8L9Ncd4CyQkNTXMrjT6V
iavHmXKoMhXaOvECUnl1A7GPbXq1H6lbBuw1Thb9EHqE2fPgivZpNGltGVyiI3Mf
PTj27cdA3XbQoOvTyBnvM6vkaW78viDyKRvBm+DkWeVWiiI9m1NhUx9yZvh2typg
U9VR1QSG51IDzdZIwqzoKXbAS3B71fLFFSitTCfxRCklEPFCEPjeH81//NLvKgnK
A4VjDZsWauMNNKn/ugBq6hT5qHas2YVcFrYKH/gombsy9ZOoOF4oFKXpXy0eSayY
YQDU3u3KHVi769fCQa7Vmpstq7QkpCZ3sF86dvsN0E0aL5bayD8ld9ULhcibc+La
TmxSQ0aw4rQNVkWEsu2FzU8MjifBgK8Zj7qsxvCI0P7sJmIUhgvMrh+FV/hwSBej
F1l6vuL7lIQEOQZTwsmC7auVsRy3sHyhbJe3TLeldBLsCdBwHUNUzy9XZqFMzYk7
tpLScK6twU2WP+H8UtUWxn1YLCys7+iUA0C9G9GAjGpaeO0TrFtd81Ag2I41tx5K
96o30aeP63Ok1mr3tcMVfU1jcJiLujXyVpiXdI6keAcAGSfkq4NG7R8yioFGi7db
BudEG8yPTex3dJuIool/yYxgL0tolwIGLAuHtFxm0FAj+q4+3HmgU8BE1urIE/bz
BKOIZZnMNyhyEmrZXVQ/1oEEzTp5Uy73w/ORVikoF3zdveA2igwJa0QuX3vX8BtE
8JKBNNJwz87npOwWeIcgiP+gTynX/nP5ZcwNCh0LtqZK6VB5Go8E3No/x8UQ4qKO
dg0D8jWcs1sOQ6amyfV4xFMAGzQQE6+oOND8E2F6Ymm9wJyzkQyt4cGMGoXRhE4C
y7fiTmatcs11+nWDfWSxWdk6AeWifISEmbVTrtmlCgkPLoFHg+Q+30pWM+sZJ+C/
ShxPycL33w7N/fyHaBqhfGdktgC44QwWYUs23b3j7mp8PGy4VozP1afvRJsc5yH+
4FFmLCHGH2JGTI14ioOhuFNxZPD79Cbbl5I+770PB59O5JaxwFOVIJ5xEokbu+aD
Gtw5r8Sy4aI+JkYQDQBGqkCsCCvr4XMhrYO2BVgVluH4rvDvG0cDRQ4WdixlFR+h
5fzFbrTtrYUJzZBYR7odK1BecKJj+dkGL0yJ5iFxdCx/CY5cJnAU/IgxfkZf8CW8
ltUvWwS6JcY4gPizjg+CWXWtB3Jpjqaa+pHyWP/QbfvKg8gCfDVCesra4q5tGJ48
MRlnoJfmkzj9gBIUy5bMiMigeYb6S+d6LqP4T2mTAJRiQ6+EPpPYRLv0s5qshPW+
AQ5T0Z79P8yNSI7QBtBn2uk0ja6smfd8W8GVFkqNusf2fwzSFd6rbLzZuIJfMIhP
P92EC22wYq0zNPxhZnrqDB2jpwFeyDRwP7/gD1AH2pWggy9vbDBmFCY6tZRE/+EF
qoGrVP7Yep1eNsmRfWAhBw+7pwoFXaMy58b7mT1cAqbfHZ37eZ1byvCzCKd4Di9L
xkslPUs34aS5uMSr49LHJpe6a5b5sWUU4RK0jTZARC4aVtRKMnxOLSy2WVfxltZO
HpRigTJl+shnJ7fwag5EwcCTBdeLD+sq3A7rrbjEZkqMdDllGQIZfOQvkeD5t5t3
dRBxFduNHgkWotK3EzhU+amoL1djkcx4xpAEogbbG8rdA904bewanyvQ90UUH2Ds
Sg3xYdoL+M7wexul4qfyvCnQ0i7eTLyKwURisZd2Q5hS3TK6qf+V6aukbA0JQFdw
EPOvTGcjZVvh0tejPmAKk5CJHrGCwVoyXPUulvuVDpS64Tphgshg8JHRl58Csz9/
eg9emojE3jkKfgruBI/8x2GKuZ2VM3PSkkunDktwRYG/fpsK+2ggeYhL6NyRsMlJ
klOEZwdQH/FqWpebyY9frwjlcJiokR//zi36P9Ltbs8/wIo9d8M7/DBFQuojeuO4
TjtPln6jMYeg5c3DkTZFDWQPDfwZZdszwBpJOFb9WpvZKR/vJ8gjCSRtBY0n3fkt
aFHKwhoXubTKBGH5+wCHBy81rl8ZLufNWIWAtq9Lytt59E/e/sQD1arkvu5Q7NdR
8NrQKryEtUBZqhYEbrh5uJWLMPa9Cmu7v46PwpjvzMpBmLWnBUY5aYY+fRgP9/D8
QEpf/kD55bGS2YrppMHrjA09zoPrMKkdQNYfh6B3FF3sxeQ7j39UZMYt0Sx9qD7T
bNBaMsWej43xNJ1uUGrHwXHV3LeL0YJ3GUFqRd8W8bxxc1gTzaeP8wn5cR+3lG9s
VEtI+VuHYZQJUbNtdov58+UYSI7ttX66O9t3wmt/jnGXMsQT55UfbTbIiVfIPWO/
v3atK9pMcjESI0fLq/ebQL2tYZt0Bxis3yO7K07cnwXyQ1nRRfgYqQGROwOiPtW+
Xg3YZs5UI+AvtS2wJ5DfXNAIPjs8NURu8BH0T/rNo9zIJx2XgL5pjnyINn2nZVFu
JsHGxR/nk9LlnTFr9oRQm98wO2gEZgifeP/Dfh5vb0GMNlC+zMdkbr/9hHAwLP4f
HJM6Bx5qn2oeBp4ozTvCCJHwVvEwTHLjAlqvp35QsdAFKQxj/LdCkZUIVGaA4WAL
Uy4eOXTKZNby/S2eItSKNBMIvYZ6eLTWd1HYb92/oP3mRyG+tHd+fNJBYcaFRDxk
aOcwqHgeXE4ZQb8xJt845UXcGwYc+90OrDzIGWOPmzUBMywBsWJJSfBfw4tg5mnm
zAFzfFAVvJfIPU+zIoN7ieGEAh217IsVnugUf/dVQqi3NDu8MqpL4E3U3wUIvsT3
vW2zwp5RQ183wlxoYjul9xXZ+xyt44pJtJTTfvArIqF+znaaS5shRB6aKQUx9f5u
BJRlXLJ35TlhYXgR+QRt+KnTjz/Ck0ZdSCILTO4doqvuToX4RDteDTxBTjvOpULA
Msm9ZSLQL3m5W5t7K4Ve//F61HyllTyEHhB9GUKzS82ol+F4nkZXRsCpJygdolVX
Op7kbwbSuw5lE3x/KcW8cr798hG1RTa7sa7TAz/JeQlZPXaAXf2w1uJ/tdsIdA09
tZDalGStQELtivFieQmubMrN+LCyk6kLdhtl/rDl/iU3+NnmT/21l2CpH4BnO6Dj
MQTZw8OWRMsXNZDMzR0Yzf9cEG5QKTYHZ6zOTcGGuHF5WbBqTGhGggTqOSIEl5Vh
JnRiY6ZNu/8G61a79Y1F02AMpF+sAxCrpP3ZcSAs7qNaVd0bGpBT3gjGUzGYhZ1z
SV2RZe+LnUXw8/ebPCVtfCQQG5XXhAKAYGC7UF42JN7QDUG/upORej8oMtSLgDTG
Rynx9GCRFHBjxSlLmIzahV/JyWytTDwqkQqOxbPK68qFuwVhFN8Y8GuPFUsBINkv
E7/I+ecWYvXzLpPY2rlph6adCM3WEGPlTk765k6pxpONYBnLjD5s8gnyFOrwr8Mq
+o8zWtbe8gEmeha/rPPBiEkmQ3pgXF51wo0Fh5enSPCUZBD/8RCeKcBdPUOWKRXy
g5TvXLeVRIr0PzS9qM2nnVNmp0xEEF6qI48nY0TLwEAJDyzXm8dQQjSkpJbzDuZ0
5D/78RmvXAZCxMm2qntQT7trha/qWOwRINdI5ETn7MV3770lP/MMNb+AJwkbJsPw
7PEydUDLShG3HpQ7kq7Miq5FTCuUr3n4wJpCRGcboDNj6aUuNxcTxHJaNKkc0h6M
OaANbROWAenWqVRAPJ+w9iBAD51H4cwaoAJ5ns2zBGrMTdgPtV1DhHnSiutjdKQ1
5igdvNXZHECfE7yXhmYo+aer9Xig+FusTRVUrjJAyJh7s3M6lWFpPiYP0g7CMNdM
zCm/AK3czWFQP31PhCY382fs5BnneUT4VIcLb3M6e/vcu+qoOXMl/aAj/lX3Zg77
Xk9ipW4heMQ5fG3LQkWDL/2acC2Rm4cW2LR41JWqTYo7ytTdBZ4OP8LEjSdfANtY
8pQlqldOC+L9/52Lr2DJo+oEBQiRiVnGG5afaF7Xv2K5IqTUnDlFFS31aSG5UiY9
L/hA1eJKTpKzSjSXGT39RdVyax2ILb3GqFfbSybAWkHyz6ywiqQImPniaOpPO1WA
ZLyTGqtBlSCSHSHAao5anueZnmt9RH7dRsUTfsaWYKEzkJpxraH002ttXWm8rHG3
jiTzMZHKgTvAtQSDOi5kZfggKdAZ3KT1lC0l6IHO9JyIswe7zLIxzDoomffLj4Om
L20v85psPXcXnlgvPizO0a6LEM9Az0+2SnrKxC3vXX+cnodRcuxE/AByeG5Fmyjt
snEKI711zTAwPtI4uJeMnBgknmqIJzCytx11wEraIS8xKD699ZZ5NrZjs197NSQk
cfdOoWH1nqBYypSgEWq+21aSsqZ7HX3ScMVczmLmnGtcJp2H0eS4fUntf0IL2eEp
ALzxUBHAIkWz2JjW6TuXyXszhoYx/msocjFB136z1d2Gt4aS1ZhtjzBWgJyFpKAU
131x1fcjnHZGWPabmBVsSAl4F6eMMT1++qK33ymell8bQhTGmvyFj7uzO4sLTlDb
nsveNSNFC1gEhcNmEFP7h+V3nwVi8Gk2tNqaSozKCJbiPBnWz6GhT8fkgqhC/yZk
VaE8b4NABKvOunSCkObqIqTNe0Dm4JUYcf6ae7OhGqbj9NLleshyJE+RXTnNH5hW
0mjXDGdx9a53OEdwQR/8j4+a/4fuDxavuXaQc0hb5Qh88PCtr5PA4y4Og3BJoliV
s6HV1gHENbtDvhzWdRQVXHIvo1glJ7RZHYHMVyXuCoDBk70bflZ/VOtEv4h/4zN/
dlaxkSR3LCbMcRTZWacC/2rAo9UF2LYs0eiyhtaFsvA6W9KLNMzuj3oJmkzNOM+H
9LAlbGbx6H5dsOLB0Oat87kI0WV0xZwwZoIrrzhj8wdfO92ah7vt9f/U8ihoEoUj
X9akEd4wYYYmlUwI+ixdJ42qp6ue0ApZuCLPpWDz2xCUi9D3IulZ7sDZ/qYgsIZX
J33AhNYgdRbk8zSnC+sBh/ggPcm1pmPDzwFOSxyGhX4atO+/Qldiym8TnGX8b/b5
oWFU8KPRjcR4xRD7Q5y9WMTStF6GiajFQxN4KvcWBeaUy2kKJ/sf7AaWXjXRz+os
L1tDMaQbWod54vawnx1Ktt6U0OkQPxH0nxprZWH4ZFTM9U0SiTyoy4DASXQ7g8Ey
V5IOFudARyfdvK+ChRpg6lar0N2f4Bq9ILtSSYtKvcYQvrZ8Hc3dvZ6Qtgi6gDSU
q9bcjdsW7BERbv/+sbuYix0WSyjBiYNKUaLZBqL16FshS0FrM3ASroJ1U5FphT8y
cyZDbwfp74wRXZQjwOJNAq+UYeY2AG4cVGCJH/9qfTFLfUjoHtNWBoxxHeZKux5N
bAQbsQ2Wb2z/+dnANv6SjxmG05JockfktBros4luinbJeJNsCRbR2v3+upvwAWBH
ivvhSxUh61nuyf7JN8MuJTVBnK+fiuG4cem3qRtMJHwLyvb7UiOqk/WwBNEAOypS
228YxQM5pg7FOVvRMI9Wgk2GZ66no8x7pyTGc7QklWyhNP6RcbGoFmbBvTwH5rSj
ZJoOFUewsEJY6rh4v1fnNP6RHooe5WTC9RlyrmBhxkXnycZhje+isISj7sI9r74o
wxkLSJrlmZzOY2A8kJ6wK7dUOYMwa9A5p6lQCP4VE9PSP+zwXxslHFGYpoXsH5Y+
bl7Rwj9FXUobq9MsFsCa8J0cSDiGd4kpxiStRu8Iw6wiIdGPrqMuWRn9vPCuJRE4
Xvup3/qFsHaz5DzexjkranpRBtitj4PyHUXEG25iVB+8BzsVZjc6tkvzhDVDHYMi
VMybXqa6z8r8MPqQx7rP7Y/R3kz6rPlZQ71/+5TgZ1L7v+f9od0wX8MQl60kQgKD
31tHjIB5VP1KZPEMmYUKJJBLoETYGzuY1Nfe9WpIP4XQjZzlljYhGtPhxDSVaKX1
WPQYXp8b4nqrVp/kEoSGrHNST9v250QLmj82cstA4o6X2BfmZHXngciHWwMamwJA
2W5DuskSjP42+UEdBFgFYO1R9hi7Ktp8TYFSeNloq1ORGXJ6R0Yj6eUFpXIpN17a
Lp25l2sgt5/C/+BJvfgmGXMsIInR6aP+RloIFBPrcY9D8FPhA62TLEfRXph3ApvM
YwyfXIQTrwbWa/olA1teZ9BBiR6Ouma5KbSuHYwnoIMsp0w4OZUNgMDCuDLmpVnT
tS2OtEknYz/N3lRoWu3/T578ECZpoIAWqOUkJpY87uHNTzkOoul+CPXeTxfuYXb1
dcb0m7Si4myqdRV/0MM9cXU5pLJ9adDhQlCoyITUZlw8jeIqBn46H1ykSc8Sdxaj
XgYqa8M+wGNB2Su8tKN/9tdPpgQDkIRFaM1+aiPjgGgiYJwDxcspTuNVcyfKME3k
tDpZbtwAjWzljGgWtgpVz8JDfyTZ65vmCzC2HzCfLo5YZNjwcJ/36u6YNvTggJEK
6tYfVY7MQwBBBN5r+SwVk5kSCaY1lGkuUSAXHJ30r3MnVn/Q7MIedhaLNGpVUlEs
EWl0xCwRPYV0SXUJE1XLFAtv9t99w7DervsdwTQNnxh8pp35l+Bj9bYUYFrcrLzN
Pmt11kk8XXNCQ1BSt9rc2aIwe7AiDmvCQ3MdJ2JomzCpPaFGKgNvmARSH6el3f85
yb5qi8Ew2Tm1au3FSa3raHgtHY/z/Wpm+ngOgwS1go4wyaxcVKT07aAAh1YXlm7X
X9tROrNjD6yzvN8ZrqkVEDG7mbHrt8LtoHCjk2hgMvUQ7m6z6Kc1moVcwLCqPuvV
wTba7xre11OBUE1vQf2Q6E4bupbvTkYKAJYqJG0AgdE64VtOPopgTQ+pR2+20B/f
wRSBkK4KIufUo7zmiTlSy57kiXpRPe2PJjKtS4dlMEfko2VuUndirQcY36euH5SY
CCek2HEgw4PNvvkQuzLagO7hbpmsnm0PwWs0UIIUnZsenaOnAmug1kONX1xfss8s
MfU/085IdeboTENFniLLLkCVK9r+Ou4vBbBM+IEQCR6gIEeBifcguw5nTnFus6dm
b38kPU05jCC0gUJrmwoCWxKDcz4vnvMbqkDItRI3Vc8ChIjTkb071X6XjfDWvSZg
uXitUO4OcObR8yArhmOHsnJyqEud7NZAtpASQEa13O5jo/rRzPKseEIXjLNsTTib
IW0q0L/HaEpxeRPOV+j/GY6NjOI0uyDZzstlQRnqnC2MUXj4vM4Hz5/atfJuPFcd
nkc6F9QW/OCM/1foVtJXemGCIJly/nv2oZ1TiZbjvfzTdNMT2lBMNYh3Mo7npzA2
6jmOCM2W0/d2P2KlAdr0FU3syLItfhM0/Sfgge6QUR7NjBAAW62eHJLLHEuhkG+y
KJlT3fY96TmYb/hLU65txCjFUGzbZs6XptP5ph4iLVHnsaXiDFsxixtn3gpysmDj
I79JW0FLvoVASKOLY4ZWsszbM4h83zBgra93Uxo45kSONHnxQ4GTLF3/H5llpEbI
oYKAMJoqcDNb2J4knk1x9f9lcDlsiqVP9HbcFAy7RzNzsazE7c15q2Dg+kzEkIyN
+4NZox8MUPcs+zRqCkhsuJBN4L3MbOpr3ogcK7NXVVCbqMOwjAK32EeBqUqVIMZz
mSuA+ArNOygiLsRHaKBFHsATXxiJ2d+BM+ULgo42bs7YVJbL9nxnl/Tnw0kRnsDE
Urdm1jDnYYJikVDq/OjkHSTmVxi4jD39pPqgqC9wngaiVeF4rFxsoYsnncuscaKD
oEXnc6UIyuQX4A4s3RHI0bWwnI+DHRD0wkzvUjmOQo7giuVkAygTGw/bvoeGC7no
fQwLZQaqBeEsUWJjYQV7fTAF8CHR08EgmkvtSeGv5EJFGXskfGNc/M5w8T2WxkqP
SVgXRjuyAeDw9Gocky1Sr51BWXOYzNZO23jwx+XmyPKHJmNvIhWvkn/W+uhQ/1DJ
pZrSr4CtKkf7W03aBEwDmlZRyj4Df8Zzu51S/RiUrRWm01aIYvpEIjyqBhI1tg1H
e5ALskPeF/j8IuGYYgZed7bBnaoJsr8+1s3ttdxbRBklKfmCu2LQ8jjpKGfGYuJe
RTHelwFL5ZguCQuWeAQIom71KBTBtB1NfMo/GiizkO5vsLe0pPukQfF+/GC3wjsl
nnBEx7W+i2NHzIO2nnFKfDUKsHdPq8HGzUgjlrREMuQibyVmKJCwOTpFp5BEYQpC
5504hgOK4KhSCKuK6Z8mkgp60+Kay8/uc3ubrZDOrkLZofYCH68p7Ovaj2YjzemM
mWTSuqtLgEhIrqa4mAodH+y2+svYSREivMkeGS5VsyBxPf6bfAseIfuCf41woIoq
eNgxq/foACiHBe2eQaKQmLi8afcwYOdJKupAFa8RvfE/Fbmnzyfcv/GKzurcbN1r
ZZrlLZUwvo8pdDndPMWY9VvUe12gMTOvGNyBLMUNd/6Uv7yoULuGcCxMPFmeeSFH
8X17tf5mIEkFFAwoEibWu/vqGb3hamdXMFJEUb8j0BuLbzCa6PXBMC9h1jkROvxd
ufPFy+FaTC20nujn10YsW6D856P9/qKFKJVcr2hypr6ztPqYRueRQwZ0Pe9JyZ3z
AHkvAaoY4J9Q1i+sbrGjzV3u0nMEmvD84cQQ0mHgcF15cT40zHMGT0Tz5qjdXO2B
asGT3GkpXIbKooePvYK7JORBrgLWawCBgesFgi0DFZvYip195VCgSw8cr7xHixyL
XYbKMG5dJ7OAUxYQSGUJJhNkRR3AQj6mkBuq0Rmurole2s99+j4o4MeTv4rJOsXl
sehvhUOy76yjscAfbJeiUDalScIub9Dt6GGRraIv8aCS76qRw6dIZA+oyDQGja5i
qDAPTa7n5ZfBkMWfk52DPfek0nUjI9HiKJKDmi7RuptNLQUMHlNx0u4p352hULWO
58yDQp6g4MEGECn2V87aeHPwGxVtgz17Rq62uqkPwhjJ7deEKx/0nuM4pHsJHccV
L1vK84tp7BQTB5D8mBvxE5HChcSSJqHMplXiKVltuKx0FexmdqK0x7H6j5q0jP7n
Q/42WYldvjq9tgU/Ko+7n0WasL7thSMBYj5uecY/bJT5vfP1va9T905Z8hhvNJTy
Q1qcaxRsPcCVXWsgS0GU5WSwHg9cpUYudXc3Ys6wkpRq44GDFOjRGhmFGL4Oubco
ogdHx9FZZofQRDuMSi29wD7QBGDhsyVrKFVzw9WHGgiiWT0CyGsCtYx13ouXuIVY
qwua85dsk++ny5RSZyyC9tHtVwhf0Ca7TctD3UXU4lkoteTf/V9AXnY8WpDAlfT0
XuZk+YaFWxp+B0gj/KGnywx/1n8MZ2fiRVaatlQY/BS7uPw3nHNUnrI67wp5nr7r
J5/2Stl+CQYwAcUghH38k/+xY7td1uo/MByMyHTmgFhStyttuCXg9cHBGSBSSrJb
tcDtDyT163ivUGwEjXpNG63vAY4uo0xpxw22ozF/dLCRs2x3DMX4MrSBs+QmoNTK
ItO+bXposCmYIjFxA6lc3aMUdvVS8AElr3tb5lQHGfPweReMKLfCGZUjlCSW1Vgs
VFthqm0QNdHJ2kT7Bq4rWmJkZKnDh9t795hB0i6NYt0rjjmlN678A+NNzOjHS2Z/
k9vmGIdtdDNqEKgCHQG7xwD1SF01YWqHb8VbZH4PoyG+jIYmbHS7YaCDZF+TE+aq
t1yS2clFT/G/ahn1mTPtFumsUuyPSKLPiqMAzx+nYcjDBP0uozC29nuJqapY6c+e
rZL/Yhxq33GKAXovOO6q8y0yGAqflTUaEVDCQjBTT8aevCjuFLOnPPdhdDc8sZNH
sYLukicuWScnTl4P7NEWDfNiKk7x5RSAclce6asG8GJoRghVMkB17Nmg+kOfJc8t
EvLR0+kLHwL560MmJ1X4COk/yadjquaV9P02LI5jMbjeuNOJlUHpn3D2Y3D13Sxu
t/ZHZjJWrqZuV1AXOqCi1oi78//6LOy3abklKcwqlyis1BLQ/OHdEgdN1Gj9wAiB
I88RNP/Y92et9mIWT0is3OUB91mCLwFCFLPEOtAmgWzC4yaBPRw9OfX6Hi2Uu+om
cs0NTc4n1J+JZsOWDwYq271RjldbQCuCAT8tPwDA81K5HzyoILqWE/LS3+xfAH+Z
HLFsh9V5kX0/2ZajojrGN52nft3rnx78EzemFA1W9A+uGl30ow8ndewyvXRmQCbe
bMlWKR2xx7vLCTeKeV6ivPz0nIP1a2WAmZKCT0GAkpeVOEWZgrDpm8lfuIqmz4sp
30yIpOy9cS4BNmIXnsoo3008Sl+DCEq8s1yrE2LNDvQlaHkcXhDO/A1+pY/v1/Za
T3/92HWRLrCttevLti7iQSwJ8jVD8hy1dDMY7NZdTHIBjQ8M6gCxtBCRRc2aHnL5
bh8WCy6affKtnSPxCqDqgWDWWsso2rldQHefwLtSh+4UP6CcSx/kvNDUOf59DiMh
oHD4yrC3MrrkBm7JoNTApuB+I9175sTZgtWlxXnC9sJN/4WzCEGlhhpdSnikmyeA
T3l/ww0z6xQM1QGY3PLbi2I2BHlqC1DNvosWFKG0+OKjgdqU4E1OJ41xBf9fPQgt
RQE4fhzdOQmnOtH6oQaHWrmWTWQ+bBmg3AuQxP587jUvUqoFPH/ZFEbGkGTnBpHw
H6graVhDDxX2GwHnB6TA4nBY5+kzr2kqZyrE/pOgX/XVFYun8AFnHa0ddZaJvIkO
5h/cbpajIPXwwSZyOJ3I8ZbJfhVj8n+A9uKmDZ+C7GnnnkOpgyvEMBzWahqQPpkz
64PyYaMtYxbPJcoMfcIB9ejcJqVO3E4LHmw5xNsxw6KsuhvKHTvHvb2n4Tn/qYZT
hwGrBdLeY/jt5ijU3d9aNWPtPBqIczsaQCfctSw8wXPNIYS6ANdz9Ans7XCGOMh5
w0ujx5rjCUIzyvqyso7evAEakv/WxZ9beAjX/t9BDwyxuZvy9xDMIpAVtsr+kcO/
uczH0baSUYqZHQuL9w0xlIMJkwdw5Bj/JOga4FeMo0VZ57dfhAx7OMU98IJi0Tns
qqE/dwjf5PobcUJdmHGi24Q0TSIx6iWPNL4GYVhekvwhdrQ+v4HZ0st9YxPaRMZW
rArMvGuPGLP2dp92GCi1XthqMCWRzgS5WidPgwTPDq+YrW/TLUbw1fYuxQ28eEPt
2KTTVj/Q59gcXY942Oz2SxcT22zx5iu+Kjzt4vGW0LLSZspJHOoktDLq2sA8ENQM
oqY9h/70PGQsyRmacDJjzUryXLTx102zwrkk4x0HfUcNdYO6WujZP0bfw0OEFR+p
WLeHMzO0smzOc+x7yXkvrHjsAR50F4Fg5EPYnL8X910+SMevvGkBvNzPPP+PdVuS
FVfgPYtsUL+gNpC6GKyKUumqTwgQ2pdymcFEN5KwHg57OixmpPAXE+O+DJWkeQSo
LlnPVFphUZ9H4HnIU8k6iNHWLLpjuEMX9XnqavwKZT8J3Xjm8F3WnkESH/lcHfDL
TUIjHJyI7Lx9iiBOedrnD09e+JL7DMDyeqVA0/201fSyYw6c5mywNU6SEiEkf68v
GZy3bfjZcnXctBREqeQf44nocaSat5EKajrPB/AK79STlYXk22teQigrb1NdmF3b
YfhN/Roa8C23nX50q4KD1o4bYL52YMonYTCU4ub/FvqE0q7drB5r6S8yg9AE8xrd
+Xpum7OyAdzAjQupXYTPxhEd/xQmtoebre4r8DGO79sygpv+FM6DOYCLQlQ2N4UW
uSGcfg3TiNQ7tsuf3n39WoW6NZBkKsdz/TLsMymzO5Fz6RcmAYgkSDabKnAqYIpN
tgU9ORjGNztv5xLbw7Zp/dgZsO8xbAXHAyoKV0oi7otAf6o9o5eo3RTBSmhL9yw8
KYkCG6EDxenauyE4KSRuEAqIhdtJLvwuxMNLu5UxkXf3sdqmwt+P9aKxZ/RYBs5H
3DfMDxbTU0i9TVG5FmMULrnvTwEf7SvQZSMonSJxqtF7GWI0qdvb9QtZCHE6aFSU
tnCKts3t3P9up4alURvn2v3ZnbrxU1yvwyz+3ZJGH0Fl5Bcz+UtO9xF99zsVYxwK
IkzUuZmVzkx8kSfggQqi8lqHAy///xcJx1vsS3XnJHOerAFZ1qA6qhW0fTsiokCT
NEtQM72OscSHCYvr0QWgSvjlzpT6yTSKQiUJvFNmm+LQ19XQmlgTLkyeWtygWgAa
O2WIR13CSMa5LmcxPsnCrxZ4qE9NbJluc4IW2mvpX6mrX8+ImdnUOGKyprM2cgZH
7JP7LkmFfKyR6vAvxgKVNAqJDsnkzdXWcCbcZcdki/pbnS/zpwfkUpMYW96a7hyI
yNDDOOgIzVy4zRDDRzNrxQLIuZNo6k9GxDGXCjL8CZ6ec3hg36PS/cfhJ+orTabg
1huGVOvbfj/log8oMqDeuI0ABx77UeeDrv7Ybwuthq/a91/zApMlvyp6hcG5iFrH
iPcEWlXWpWivZ9jBl4rO1zT9LguDkDwuTL2ZKbu3snD8O42XqQEuzyPTBbzXZ0X0
tf3k3w4BYVes3P8zvYrRY/zacGdYi8WnhVzN5LhVEaPJ9S0sy86pKaTKaVvbA7W4
hr12CTb/Rjrm2amchC04xqc0194j+ulUaC6LqUw0f+U/KQk3BgLaStZhlJVDL4Xj
hFzYwAv3oiUSMHKYYSqoKCD3Smm2Vne7XN+e5BEEQw1h4xBNdt5mOT8uku4SW3zT
0zrdxyKkgQvyUYn/kIsCLYuC8epPrmXs7RG39wToLcIuWTAzAKywzfODuWmV2245
/qBKD6FFQvEEBM3B7V/RTIxXXqKGaJG83z8UH3q4GzX9P8xm6fiX8lSQWi343RLD
sMGNH6fxVxT7lueojwcVMsBe3nuS80ns1b3s7FOR8ErbZ+ipxwiSWXy7jE0jNguU
l2256JvCCb4OUJK2DIhHsz+1mEV4jPpI2rWQw5kNETY71Fg8B6/0lt3WN1dCuDc/
fL/3xSzyvIHxtxClIl1ZGeTHHPWtO5hTr7fWeBs+FAuaYA8mv61xiWeycInzpsAa
pqxSiTtSHm23ihOrztzKDGHvxYoZRshzskKJSYGGwJmZT6Vwya+fy7xDHTeBy2Fs
HCEKkA5CLUSUKojyEswyIkxjZeGSj3LTtopB21X6FuRV1gsH0TJJNG4B17f/LXEs
tHxb3xU6CCaehr9nGS7M6CMWAPE6OH5Gz04yG7Ifng7Yf0TsmsUBc3Z/tJvwQyYw
YCf3ElarIoqH0f3ieS8Mm9im5re6pAUciYAoCdGB7k16CAlm/ed3QbBbOA7BxyKE
S1ScHHR7+mGzkzQAifjZc6RhNYE7bbV87H2FuK2bdSVvSG1Jy/3tNGj0134uECDP
HsUWjiUyCIefI5MTCYFQ6CEJ4GzNpgFaTT+HKYcQmgofmaNX6Zlu+5HrKxmJooQ/
+v8ottqfr1kdhupsobUd6+BQbJvj/a0NTjzfAQhuJFWdqAs5q0ZO2Cw3MoX+grZK
ufz1/MK47c5TG6RFqg+z0mmF2wf2zYV2kGwQ+b2KNJSTSPPdRkjeN6ZriL05lbNN
yvD8Ygz2lKrdmEEg0ULkMixlJk8GfNurF4FWGOhk8AhRhDIg+qSCAl6xjMy7SYlU
8qyGBCgiO0FF74Os4SYhFzxAF0sTjxRwhg75m3MTQcfPnhpEn1Iw+CImfWsIRcl6
z0sAZMxh6AZ07ld2l//QqcP1uMU+OGR2zn/iGoyEEpXSmpwyvoI+msEOIzyxRPzB
jF+l58qorvs2K6d8UwF456XZ3AAyuedVQhiC2M3IuHwNMdj7BjOJt9rlnFRpM6E1
TNq0Xay2YPtEHmRjwN+XPgM3QEQgLtPV4nJe3RA58Ai7NbVfL8JYxLb/FtTeA3hG
T8Tw6V5PXRKihocIkWR6A8+e6qRuuJGV8NzwTr0scB93zEmvti6TFOkb/8C6C2Q9
HR0UHqRluRBGBmNbVNDA/KL6YREdBnbzOtVMSZf8rUE/k5X5bE0eECE3SMipuxAa
JbdWaq16bhFVmzLHudDzG5pKIO+k0XQmGuXvIApxsxcMhQ5AGtve/q8TY/XpH/0P
ElzS2jCqdiDN0h047yqr7epXGBiDr5CSfZk35bDRu+HNFZXrEuA+zlP3aDdj8jAR
W6xmlPT6pJ7tbIcnvc1jSaViqKFTIqc9PZbIhzpPKZI+ygr5s+U9nbixUnkQI51Z
kJQtCUMtL9wSI9KrULnTU6qoxq8dzmZ67Bu+KYy+4FrNdHwnqy0NDxnTGusYCzOx
FG7waEBYFNruOXEvC+W/B8XCfOM+bzNPcodgTdgXTBYyTvKQHsKueRiQKzQz87qi
/fpVH9yTAHF7NlaNOXC/P1pdrtRQW4IyvCthHVfnunAnRf1skDWVM94RfvQvtSvt
7oGqmaVXyI3MFEo1CgGBRdEQ4ikGhs6Xa8ctSjhx9Sx3WUSIyDrDtQELYMf153qS
cdYnVYJH5juDg3r+matwgPvuCwJYwyf5DXalBuCfF2go13k0fx/cQ5bONAo+B61f
nVKgscBAdkOzq7AsP1degGDgMlfhJqm2xfRQ8VvnRcjcG1gu9t9OGZBwIQWxXwhz
YRlKOKBFs4HRvlZzZJM+zNF4vbou8m43SKfPMfEFu/tPFDyay0P7sWUQ/6PxSq3O
QlEzE03Mv9ybp+5F25Gxc4lUCefsmmoTU2KeBdQpmgMAAOo01jf1dhxhcK5di72s
XnbtOs8WiYivEO0ixxMBQnVLwkg3KX2a9T5wlMwbmkgNWZy1TkNw3vp3C86AuBcN
27yq2x50VKU9LU3p3tTKH1dX/xE525i6zLWRjNZ4d8OfX4laz3j9bIAo6WNXY00v
7T8mSwMhvOeMtCDCtMRw5BXeDa3dx5+X2QknEpf4Pz2erqjf6eSLzc5C5ZSdAoiZ
P4Ph2K4NiBskQ3Kip9/F9Qhh0Tjg7OGZrbayLeAFU7V0e5/8j1gZuBt9j745Sklf
T3X7UFpLt2Y4DDNyNoAZe9Ghxs1Y3UKllYir+xQY/79rrc4QkHFvLCky6geV/HsO
QgvqYwaZXODC3kw6iNfDFf7zLuPT+mCBX4EGwFSKHsGzhBBIlBfzBJMf5BAbdlWY
jvd2vZs421e/lwrfS8Dr5Q9P2dsyk8sTxY10BNVVmW+I9qxhoG2OBoPXAF76AOgB
cPUFKGuA6j69RglBKWdCMmbuDQrY/cxqBguFKJAozRUjQ74ifiyxdp//Yj4awYD9
lmNzr29JpClfOXAAUb9RRoly9Vm0SnyJQHwELoDHl0ijdun8T0OI+bGaYSS/L+0H
9MBaWpbCnw9qum+JZAUQEAo8cbDEUQoX/POrR4THVrt3uOkvCPEsdJWUuQYnjl1b
XZDZ2uV0pp+uqd2WDbYMS3wTAUimoGAz8xHsDo6y3f7NAzaUMhtef1GygcqTSmeU
CnOIrvYHU5lEWyhp07V3K7tN1PYalnEf88IkXgx9lj12QhTMMCwS5Ahub5qwoCt4
Gsvmv2/iwBN+tOMdpscLf5r2NLUPzjPMntK21wiMBRz+koLw6s9/S3AacDp5VS1d
HfO6mEM0pCrR9xDfeYjXFN3i7aOu1yu378I1mDK9im5DOqCb0AVQYHvmItdYo6+T
ki9uz0cqxBdduochUwRsUHRAOh1vaDN/afm6B07TzwzGjvfHkDMpuOY/7lOXKr0N
oMAa6IUdRmXbLPlr6+BZx6NcVLOIYRQONNDbl36BzdL+jrDN8OtfZw3Y6uunDX5z
cd5jfsBdCO7Ac1YXYpMallX2io//el54wnvERg32pdMsxCjH3HoDdt8MRixaYO+R
ytmIFLHfPJCv4mJVj0jl2oe+o2A/NDidLQzfk7iC8CUtFODlwY/BTqNEiXIWmMsd
iJ0413eQj86mJr6Xud63argiFthFbrsA5HZJekO287XLUDPEpI5HX9+ayh3iTxCw
wSVIo1uIGEqoN39BEXE4xRWImqAozE8rYbuKYq0nS9MO5qumj0ir081UXvvIHPA+
F+1d1JVtKX/Eiko+nIhOTp3TNzK1nHQ3RUMZRH2dNkl4961cbmZqKRlPQOu1IRYK
i9Y4Sq2/YVCPI92FNWCeI4Jo18J+bFX2qpmNQGtth6myR71jIuJKQ67ii8fJTraj
uejOE+EkyriCsl02BjQFLEwZKj+B92oJEKnllObnvNci/o01ZpxMPY8EfGZAX6Hf
Rew5lmT+OMz3L5QDFydeiXZubxEID4zEBjiDLM2TDufeOVnf0Zh1Wty3OwpAOWoW
hTwUNDfcC0siCCv2/e3T6kxE824VihLuOTF113622jwXoK1ylkwz4cEgOr0hG3Da
W5+XQR2+Nsm7/tm8gIm+boOgvXEjMR8C+xWaXg1oAlty1XG/v9hCPwIrmLDBH7f7
u2uHZIy8JjKXhEKs629CquTkzX521AeG3up0D9v6vNlvVutRoBZU+PxRPhbji5at
jAISiIAakKx06oLKXdNA/lXwawYEq32zITMA9wwdt7Dzz+km0bbP1q68hBIlc2Jp
w2oz2hswnndT3eRb+b2jW7PSMFzF11d6hAWtR1gT2JH3IFPeGsreHxXLoxJ/EJGV
bcfCNgJEwGPGMQ1Cd3wxksmKtIZYQXms+jOIiftJdFCqyjMo4/s2EkTHCBWA/074
t54CZEnt1rFivl3kIa48DxDIyC4KV5UpPggBu/i5VN8UNTK8gpBk/zXf6Woicdtk
RFjCim1fJyrRq1xUM4e6Um5FNEP62lDzgalXEKYeDmGa4ylfnTrjwv82Md1MJSDk
4e8+eimL7EP2oV2q1ZsCm+ugMiZfJLIlwUaC5t5qI8bOUKd8ceHaypv5nVYY+wcv
2tF7A34fOFpLYVIRN2PkVN+4JDaPS1fwz6m03ahv9tRJr48FMtuf8DmZbkplseNm
miSsXA0o/fM7PemLvCW/jz90DPIG0Y2Td+zsh2JSgy5UFgTRZhFJ6t97jt/t19kI
/V5Pfyg+CmTeVF0CxzG9lV3OSGITMfhxSSrojyjoXYQRwlxiDnUun8pUNVrqPvAf
5LK0dvHrQwJmMMu6HBHZMNJ9p9V1MaMfk5vaC8HZ1ONhOf7Jz3itTntBvRbko5KB
/gUbP0qd7OPXmY6He9+teuF8cwgl9TFbJEt6rvdb06wkFLo+ul6O60l2e93P16+V
d6+uO4Zcy0k/mx/HAvalfWEXloxD6ZQFkwYQY7cscTHNxm+Q11zUypH8B6QLAH0X
DQO1gp/eDJe4MWMnhv0tXLp+pGhEx3SH3lBGYhvfOMdEqS7O1zarypAhnb/NVLoX
MhuHpROEaYWqjJXL6t7L3IPeYBRKxN1SoU188inup7wEcR4KRx0e43aotxvn2Y0G
gl6WdQD6xZgS82me6G4zvxKX0Ofue+KqDn309/Z7SgJh9K8E07fjhzCQKEdrLCUl
DfMfe2Sp8/Hfjrg1h1YAvTtNsj5YQ1mwwUa+LN17c/Z8WTUrzJTzQpQciGxg3USh
D1mrGJXfboKKmMDPkf2iM9R6vTG6LsdsesUvSukrco/u5B8iqrnRHSlXIdN8+4FW
3KIt6icMKdpfWeh0nDuA7fmoGbc4E8z8sGsRku8IKcbf7jhU0Q2xxT1dGC76XGwI
LG58uT+FhapK6XusExv+TEiAmfIz2/igRYnkZwtXg+y9ZzM0+Fv4gLIQoNaCwJ+X
hMSj+oMJA27t7tE8A0N9NX+tda5LnzqxFJoJzdIf3f+2yap82/aZshkxX1AB2aU6
ni9/JxliSsgwcITqBw0cqrx8o0/h5D/qfdEjBs8bd63QaRADMR/xWjmh7LHoul7D
BWZXuVpVVRcIlWWQIYEYPSM1wXmsHTcRtcec4yiQEVs63pGwqzdzoI6Uf2s5VdIG
zEsmiZXBvzP0Mvc7dMp5gSRJqayEuM4bIT59P5WqiMoYNxtlCdm3bq0p/3mgArQs
gMw/2bwsQ1AETKivist8mGJfxZTjXdroPtatVL9/JkCn29FHgwlagJW+mQC/DKH/
qAw8Y2gF74PqmbIJZBGYPUpO9iqfkI2ph9Vs6pA6S1Ij/UN2eswRQ22IIGbeKCIz
WJgVphGjOQQ3yjzjnKLDyaEub3vnV+WwFmjn6kGHqolShi8GpTTl0Z1ckFFX44Bw
virYo3BD6V7UE9NADbMaVruoEgXamhhLwVmBsdyf77itJzOwlT5/c/Zb05JAvubf
giDpwb4AW9fAgG03mNSPZAlpVElUrEGv4RUYfq22L4w4bHUaSoxXyn46iTeAtwX8
8Y9khSTwr1PmCf1ZzAhDrljYA1AGixq5QSK7Qf9zuP6PoWUUuRiavzNtrcBYjHB/
wjsndUVeT/ICMBijLajg5U/4ey9VwVp4QT0rYe6/TBntU5wRHKnjaS+2LPZv6mWx
xCK5PS+BxniA7+JUEKHQKwTmgHa87tUlrg77lgisOZX/EOEX6DuDHXI3RvI8dZwx
PMs9sLmJL/AaHpMw48N7wdPved1vnWdpfkkUgeaH0bXueP17R8k0bE2NcZDDVMW7
4yylmJoSUxLxjNqxyKOclxgXxKX4d7E+690GCqfDIeUyblIZshsJ41tyQaO73SiR
zuH3IzwRREMzz3yTn83RBN1fnDcxQQC6LhqzVUazWskehVFfOTu/xu8wyCmik6U3
lN/9Y9tIvuUc4zK5cGSvD5RQ/eFeioklnDLG1HDiERDBjuejyVYX5w+QLir2bT03
vY2jdC81uLUpqBABnhBf0agdmsfRvkUoZVnU15Vu9CSX0sc4iUKpS+LMfB1HD7vg
bhN2eJGUCkxvkjkf7j5rSXVM1vMtTgycF8eGr4l133EsQDsaTj1I+PfMiu0mckYd
D0cMX1vTW/0HI8hJb5iLjcGJF9llYs0WvuBHkbAPwjqQaZlcXfBexI+2ytjduaEk
vtY/DfNOi5mOvAwSIew3cl7XyT8iitZYnrGoANPY/yuHsFQXwLGxYw8Bder4cdKC
Ihb8rdMrHX3Mx1gwKHM8AouUObtsY/eNDeWd1mQEaMzkFIwgejEuYCaUo1+X1C77
RvUVZ3YBn+dKbu2cwh2N12eppp3/Y1z5Zkh0opWdIU127Fb61UrZHFJzd4DqFHcp
NIKVgftX/Rfys282AXOLajbi+M9Du++jMApTRxMULTSzDnXyWHTlHg+V19EGmT+c
14PsnVcohAEwC5siG3qBINxKzvb7Jkqu1HjInf4/z32UtDul6Pyq7EnZsZx+9x90
oB6Kpj/3RhXbCY3yF44qoGNZpPN4cwujxc+LlKw7EeGuFewCs457o1dcizBgA+qC
Kr5iPuFBoVY3iwnBnXdGArTJ2P/MHLgPWnTeF76w+fNuE8iJp14lfB4jOT/Y5BNM
Kg/ot/p8s6s4NUOUZcKgoZb86pi3NW6sE+fOg7UvmMXBZrSkAwQKwydnqgPY/kq6
B5hzyrTmgU3DhsyLxZ/FRmvgOdlx/dFCsQKOxFYg9XcnzO9i1QIN8TC/H7805CGN
pRLfzMsThwFFyag3XB2zOC1u4fP7/mMjMeJZTTn6RalEmyPBdXlnNhfWsmgROvOW
xnG8YIbPuUmR9XqiD5XM15raPJg+t9tH/4qAGSC5ZD4xP7NVRPSyHOCeWkF2ltmH
Y9VLqKnEGXBelWOhQSOqUTmzIYiDzKROilfsuSQZ33OH+NqEW5VigP9kVokXDhgF
r+m4x9CgQalZFMt1w8kvyyl1JGJeiswMUUq9OYuqGTif4pun7+Or//tEp3kR74Js
VoKe5V3f+x1i5fcourh36YJg15BZrhT2fAR2kUZsmCZpU87DGMm/UkKgrycOHxLV
R2t2CokJlQ8tHAo9rEaOzsyWJna4jivCHnRsVBlojgwayngClxdUzZ/D/3pAiHmB
iPUeZJxYwpwykmAE+r4TE6nVJjH/zbeFDWuxVMpzVDP0Na+ulv/ZXmGZPdpZjan+
XobvqGO/r+ZqIuLhMij7melCB9oasHau+ZJHzXeEfyw1LYFxqghftlptMdwn3v2i
eXhHjiJ8619UEM7yzwnTfFtR+D/UnO9Kc3ubS2c5lfe7xmI3isFVFLe+oCyV1qn5
Rk2oMrJXvRKPQJQ6FgrJ0knclYHr0ub2wc1Ekykm68c51J9WQP/44N90YjdfGZYd
m5MvuCrvFtHvshjxq6tVOzChYY6xrhGuqnpcVQsTYfynTnPFq3V/zemRudTZMoPD
3OAbLDGrduVit5dbY5709lGImCQeNCPoAwG+YAfFK7NSG/1l+nH/zbm2Wo87ZdnS
LD5a4xKYvCjagt1M2LXLn8vWSj4oy0ZnVtzXbsMO6/N2RjILIIMrh+RBfWW9MXm/
u1F44kPi5+D8qg/thCqRTLcdHWS/pwU6kKWZZk+iuuzMTKNNTnu3rxUT7dBQ1k6D
QDo3PjlGm8kYOkVGC3aadHwu5/gKWjcNtUSg3r/Rt9tBlMXQeLOkYDRcYPyfhQ3d
4lFX+7bHRztQUdCIWmfZ2uD4aJwoaIRDQjRpAw0nyAoaacddM6R4MEv1jIMkLYWg
Dc2BiZNAVyP+NW7kbFJg4lx46qjgFTxD05ovBWApf6aXitKsA1ggo5Am0KqU3kyo
51RE3gtRxGZXsftDmvWBh02rAYzWLP3xB3Asp9yJvW+9tFhgunJEvVeO6WVWKYy/
W/lZp9imMPdHXBg8HiRFOR4tty+///BGDVRuG5qdCghiM19VEBybBf1FnGc3DN9z
fVlbOPSNdUiCD9hdPrHL3R+3xTK4comrJSlH+TKEG4VL2kBAuY0VKNuy3CyYHThd
Te7LceGOrbSiTsX5yq7GBPJTzDnJqd4qsNd7mNvjUGHgVXgr7lNBAjRuGtRjkZU7
T4/BGTjCuchqpSLb8EHjvl9eRmmjMT5hys+IMLqmNO0LxB+ObEvawjhd6CcK3qLs
ipfMrUZEQTi/LynDLxe/oI6Nubq9EGjsEDO9FFN3Jp0mqvs5rCRsVQ7+aYn3U56X
ddEg0YkuUaG+KFFcaDWTj006Q0KLwMvuHM/dYvnst8VGYGWeZrKLqOlx2Eg4Td3C
snfPy4AE1GGt+PMH+Y8CwSdEAMMK/NOeiMDLkGAAdL1/NeGyptT04ztZl5ZjIWur
9mvm2ObmRleGsmbEOZFXwjG//+U2JP/8fC3CsITMCK8yBoVeSNnhIOhh21bNzL16
yXNhUktBIMP6G2I8J1bpmKthJoPafB3IBGsbRD8+FRnbXYucn3uCnIf3Vn4E+cI6
QXW9Ll7+xo3ZJ5bPIL0YUGXy5qwcP7gqp5ZaNUtI8OBMgKlukk2hZZosT9JvGvHc
XKvjhaWG9MTxPVYDc/hxB1LPfJrXsxJZkQjjFyg59LrfjZb7OZwGEte2OMAVeN6j
bhxR8zpWze+pFw79naV7eLFWy5MPYp6pl5Mq8YzOlT47Oz8mS0xIqyHSKXUCnqtQ
e7UFCpzo2Ynn+iShyWDhqhXMqMtQK0PFA81y7NnD1ALuQhnVbIBIZYvboACviCsh
dhM5f5JBRfmddWdoIuNGMr+xBROFxE3sp4EXvqpLxZs2CtdH4IPIx5d7X5Wqkv2D
PCOYO7joJ1K+XLV22NLzF8TOjZ9ORbx+L0DWZspqnMUJyLgbfPCc2f4t/ZkbEyuu
4mqq8gtT96P5krnjlFKemBwQlvAmLqKUdEo9hcJi3OYiQXaCQ/UG1d3NdNECb7Wp
vHxBHhdeqPUKjRWCbvgSxzjw6HODS8DnGV5oGUcrRMld+pnS7tatirJVSsZvp+wr
NC9heo25Ag1POCLLikLUQan1Y+9em9YpeQYeFyzSKNOaTKylhLM2+CbGhN9+UcIN
qe24GyyPvVK6U51efR0jLWWKnFbaVkwWhyLkHFHITb/eVviuuKB9fNyO+IGnhFb7
PezqGEPusJz3iaMQhyaAa03qQ/r5RWWLXSXX+p7tTZ7Gcon9clrj9LGP3hczq9fb
Ef9ReABTl2q3muvxh3sEqMxos1LCdifaawFWaKS+jL3jockybmD0qqikattmYJ7o
DTfMHt0uQu5Hvs7ESIFMW37kfcf72apxKsKxEfE38kP/NhrVA7PAUX/Z/KobuGuZ
kg661S08IN+pkPcRi1w+Wvr8m/Y5FYlkGYVhaf88aK8MqaYqEKBQq2NvRR//1vgT
5nmQqawocz22OmNPScP12O1VqQJeCD/+caioLgBvegqyPTMJpjBoniSosw1SvqyH
oMbuqE3/k+av6Rxtuqth2Dz2Js9kFu+VIKp9ObPzdeKMtj1QMHo/CaIo1n/bF7VH
RVN46ZtYZsrECUI1sdo51C7xClsLdI9jq1f4w5fsMAdB7uZlHDPp8rH53aOO+9r0
uIgnwRYXQ5KwSJP9ph3NHMer+3tA7Z+pN5czRUvlboheDu2Dxpo8P4DMFBNxDBs2
Xr8m2PmCR0azwL8nW1lXdNx+PH9VZ28jiggNnWja4kr10qngRcQANVf+OXsXJtWZ
NQjmprTsi71PI5d9j0lhdW1aSl95FshHWRjuGoBkol5Kg8vkc8oh0ZBnxBJ/S4tn
mTY2ejDmVS4TxU/OpN4M04QtuAqXidgbLqsuondoOrMWr+rOH+WssvU6ABLrDvol
2yVZn4cJYcuEEqoskY8QEMlamgTUJcTwkDcTf/CvdIgD0Z7/sK21tu5hzpH75Sm/
MIVvDp9DtlUoM1rG3HGIF2GBCzWPDCRWPmCIuPWHEjD749UBmvlVmpxIidb4a/G3
4ngw7Q9B8RG4E4DgY8KLGwsc7YNFsQE1/LDDxLqJX65ZiR5Ur4CqTyi1vPoS6c0D
2Be29xHfj7RvHT8sfY/8tAEqj0jF7rLxDXHKGZuJedmjKJ/b8ddnE8//3W/uyp6d
ssSGb/ohql3uFoXyW9luj5xof6Kxrt50fEm4d5rIFGhviqCw0tVK3lUvmVLXo1aI
BsClHwypE0onEhYNwqoQGhoIzs9vLWobAMKdCRWPVnahmT0ybu6QlS6XzQBOaMvN
RJiuJEqBk6/n7wjY4iNP19BAYWIg9PQJa9LM+2U268toHbIvt2yAsgrfzMn7G2op
5HKQ/KHTjve5TOcUHHIHZ7gx1kku9Xi8sH7uu4nBd+YuAWv3FH8Rpe0kj47P+B2g
8bAHWtNN6EkCrmiNRdPmF8GCOyPVNPAShwBam2DiJ6MZMl6Ss76lO3VFHTvFRlz0
AQPcLbMutgeBc0blZYgvHZ8J44SZGZUb+EO/PZXj1IiVLCu64UI2rM0Es+kn/RGN
qtu7GkQ5PyrGZDEjSvR7pSqt29XhaRtniqkc7FRDBlvjwlppIjkd6OUj/iDeGkWv
hVYiGo5R6u4EKEIxnPAjV8X7M+JvG0YT27jIRdKL+9IKR7aAArADqT62Ud53QpbB
sAD0NJ/gUCMlt0RZ4L9Q4ul/TJKUfo4lwesfTiMDPZ/n5ZbMgs/gjwF44/Rqb/KH
jDGXSB/JQb/IybxlS/9r++pGXCR5INE0iGV8JMmeXkGVzYDMrRuDCdeGGcGstlcN
tdgZBflYfSHtCBytSG2VrT3KMlD37UW4hl906BXQCrHzMJEnyZmhU7wDZB7GrUyt
TnoiGyx/9yxV6SZrSqA3GJ+eeUX5n4bU6YGbh8RKMRFyk0GIqchQx8/a/v26SR9s
gd7clIjaNtFBxTUv/70WpPmZ5BNAAK4d26J5F2kDy4X+MqCc5AFZDbnCLAX9vebh
VxS2WFwlb9pdoY/BJfnZTatHSx+aRJf1p6ZW/2+cWIQV18CGSRlzhJGwV6ojOaQd
0tDQWHioVcqNc6BxcZNHlHnX6zioO4vvde+JC1YAiMe5vZQqfBAdOqciCJUDAqRU
hTmuSrOmNeKAJtwCRpAYjSJ9Z9HxdcwAtIaky6LjmLzF+C77I7606xI0Twizj6JY
+KfJupnKfkO02pQwqG3615IIJrpanlFu5j/cdDjJLkPbvdckEXpvQzyXPjAH9Kni
h1fz957qaDtW9O0TXgcR07aYXGOkA3dY7gDW6XIQkQef0vNvEtjjmWZljPEZbuMF
WbyvNRbICPbbNjiWxzSolFlYoTUNjF/I+zg2bSCpOYTPprF8Rm91mRftQ4vh4cfA
23kGteggFW/C5iKgD9NR/EW9nU3R4R/zqa49FlsAO6b9LVYeAHMQtXrp4GGHVPuq
qts0Gpd1E+7way1X6LZg4/42NR4rci72IbdZgt7rqfMnnRbovVVQRkBgon3L4jLy
V+vvmfpxTBR9rWtU0K+etXSthDte/hzvcwh2+caq0nVsCKzArvfEqRgkkzcd9Ryw
Fdk44xkDkzQtcVH/tEX9A2IW31Ql4ROIRV1iMfNleqjGltHx9/NFrJu74em/HPcN
AfXQ3lDkF0/blyFyYOCbhahV6IbMXH6i2uHyMyLptbtHplOp0nVmZg/J/QkyBhqz
aU0rxfdmcIU5u0Z/YGsvEoQKQeHXKiq5jnYnBFyPOcX/CGBxeuEgS1qLxTy2jstA
3FsMhQ1h6QScswD4V+a89Qvh5ce9lIUGDzALkfpigUbOW/qzS8Oldfz9EzBwKHdu
5InywAneEXZGkMnmi28SQrMIeSiETnq7ivwm5tyPVzLAK8JFJ1KzqaDyIsNqwQWT
IOWTxV19qZ4o3clavurWu3NzrPfkOh7Qz/xV9WqTBYbGFDnoSBYVzpmhx1hnuSPE
9mheRkgBgzGrbqAzE59tg9Fx7NbvMeRWiZaPLgLR/kVGHX45rdayJwz5O8Gvlg8Y
aBXU8YZtE1Py1NG57WuqlOaOm+odS97kMGPd2qPJyhTRSWcOwyHkc46ERWNdf+G/
4NjHbMURjZVgMXRBlaH0QICxxVtx74SqPBn8nlj1HMemB78vQAhjZtE+Qm5lz0xB
fmA7KlQB13H3zUlN7oBoMaARdeWwRylyAV5uq3mRzhZMWCcr/wMU4KR4BLh1QPBa
9wQKg0GVduh98zpKAvPMiIaAlrkREGt6k3oQDrFa3R3/uvIG1r+bcrXqQ9sooF37
pHCiRVLqKFD88TyEiz78EBm79vHt1EoLxgGr+/F3UVyp3cN15ao71EdCd/Z56Ldp
5Tx9nYW5KV7wQVIdx/WO+1cR5YHvNivEv2A8Wn8xXT+e07+2kV6SFDAh+Mir+ywz
pjUi9/mqh6UpI2WlOBb4ni4BvDggU+bPzsKBFmP0J6woDWRpPZRQujEGIDlF8P4+
e7OhY8vKgo90t8kVQNCLl6HiSjCgBerAGuDKmymqReTsK4j1Hv9keonWsKid4sJc
+kEonjzvSo5DbtfMKC/jAaHo9ziTyZfSmMSa6NYK3JkWEota8b6MpHzAZuscbc9t
LCiFtBTvfuZAcZPBqGl/wgseFpM7SxteFK99zPFBFt/K0YtMfuVi+48n9G0zXU/k
ru2JgI7xCA0mG1/swosRdH0hkF8rjg+k6hSZkJ7PmDj1OhXsZz9L3CSly/3WKdpa
GX6nR5n2u/EHwsY+Wah/17H76zHcn1eJFyzhrvGaAXRJQaMxxX99wbI2gEg7YNzh
1hCkoBK7cFn3RMkOAqUfqeXC+UOq0VE8pexD4uPrVnrcm1Cxte67bH8z+m62pARr
5KVPmtkgeuuRpJ/xMrb4ZPkyTIgaI8z3AfXAZlcajE9qv5GEEYevgz9WUrnANqbw
kmakP3yHXwVj9J7wXvVqU++8EY1JF8IuaqdYlGzB2n4QSjJPGnfZ7+Umv9GXw6H7
H4JVNlOZwlMTPlGTj3Pv5mFsM8QnJ5B28hoEw/Wn5rhx+2HF+aCKkhO6q63nmBDT
aZsooDHy6mOUHLaQ5X+kQKHFQMcoBPlH0C0i64BhrrpGk54zdMOlzMlf3bCrR4Zd
XfkOHJuarVB8uUawsXxZ+9da3orwIu81SyYhkD+CSQtdv1EIY75X42YTwGeCB4F3
0JalIXVZrltzkdoCtMYUngneL9OLVjLrzMV1+oy6lMFwBLszidd2VO6B+0NSETW7
7N3AwKnOgNsiIVBeoXM34bkMBQyA/lJGm47Y/LQuyAVfqnYpp1i0GxuVQKJbQKJO
i+AhjVGRPNOO4rCA5fikNuqf7HEZSJ2Vk5twHNFmmHG2rUjEZzHAHRyACopV+qjT
4EnjTeNoY770v0ut+ezcArhHLXOJJayJ456Ht9SkiZp4pIz//smyuXiNgphzi/Lg
LpH7VO7ljZF040Y0bVyhkOXcjWKiQIm6Pf33Uq/qCsi/VwCIFlRNQWoqqNF4PT8D
qTOnXrDWb2Ss59tUyF1ac40idkEHIFnFjGB+7i4aHmq2WqZLWA20+hUOqeB14afo
1hI/7IWOS35qCO1zSmkUR8uaB4x9ilNTBuvSROA/0EBghX6JMuf3+Dd8W5yGQhik
2Ntr4vR6L1bfncf73wpIWF7kNrQfKgKUYjIUrOjADckunhsZHfbNE4IZjtqnlxG3
j1WjyDnxEYyeDk9SYmA5JfokPw7vijQM9dQ3MA/0OEPjwpMY9d/XvT14k8kT2xWZ
UGg0iSm4WYNz7dAelAzva8ERIIexgNE7lx2z/lpJhtrqi8xshSa6iPJqVd26mE1f
UjCaNgBsQ1aALi8Lv3naEL/UpG9ybGctic4JX42+Cd/I+M/LyfhPMXRKlELVh83U
CpY/INwXuye04WwQMJrRnZDEL/L3XnZjAwzyTMtRqtXrKxDvtYEhAU54ClCzfCjN
UIQ+hYydKMkcu4h9Bq2LveSTLqrHd3cDRb/qWJYIO2w+ftyrW/mmlI7crKSyxRtI
6EUhf9iqmJillSORiM5+/weG/gKzYFzXqrErdvJYJi9NlQJ+k0DjNOhldECuxpPP
b/B2qfEUHP4E2MoCocQcGn6+z63YWK3P5FtK8nfrKAx+GfS866ZiyfXa1oA/5dq/
2HEwAjgEt9ACS1qakTh2tqPVUAG9Or6HxJbTS4/1JoVbQFCOdXjJCJfXsSQTFkht
PV93XKenJNlBEOd/1yQVIJxUxmMX9l2yR9Ym01g4PzYEIMoCK/LoqjW5o43vF7k1
ooJFHcPYtt/5yVOfC+bT9l5/70fasK51NcpgMTH82tk6CTpqk5e7tBamczt8ypzu
a9B87GJYJeCSvyOgiMIIyP7+5ue7LW3ZG5pgZ9p7UsIvOBRWGdUjoOEcWTAoe09i
kmGROtnvsqNC5CFgAw/dz6lS6i2Q54ZBi3ZcAiQKrWMtSAl76Re+cPVdYmmRDKI0
ja0kI6xN23BVqwBg24Mjg3XeDH+pwsbssM8RCp6y6Blr4UzU0oIX+/L+gfkoQoND
1e3Ua2k8nVZEgM8JU4wSF+rqLuBcsC5AQnll8qVnLiuzcar8QjZsR10c/81p2kTM
9IlPjbwGAscnXP093ucDt0D44PtodCMNhKnZg36j7K2/Hir2imZfQPsWJfZeoUYX
PKaSBHxVuKaqH3gowZODpRBYjhSvywyScs0wJIZCXaMJRpdZ1jES8RhWInvOdG6h
1AxknDAc0Y7EQw4F9+XAZVZam6zrPQ5HwAO0DmpHx4Q9PZCMZ0egvul5fYZ9Nd8Z
YoQH6ldFAXNkjMiLE+K4nqjNJw8dGWaNYbkXW/w7Dgv5jGD880VomeIYZwI4Zok0
qsyLhgWUxu8XSnLUAX+Ws/uLGRx9UYNRXW+5jRn72MKnfnDjBvrAwFBZ4/1KbIrP
GxXk9NUla7czY4BoQK4prISpfQ5nh0b6z4jtxK2kEFWGaUtG+2YpmORVwH8zF/+l
QdJBMmQf9SeltESWdss3zd3rVf6HZZIg3T9rwo0G9h9rI86O2fPUOt2ks1IuYUpS
hJPOOCK+Hl4XokYAdQX2CeoObWxs4MWPUY3q+cX4vjYKbeIAsG6s1h7bydybWZ1J
hAQNYKBlS+wITgJOU4dn5fbnM1Q5Q3LdTf7xmTCm/0Eo20Y34j9yJtjP5IgNgKUv
xsH8a2fMb6b9rzTZ0GDUFzs2NoGkeocAot5oGFQ/QSgqp7ss8dNaTn2NV9IVQb1U
MM0i6NYGEWcA1MEsy0am5ISEg8cj1HysmJzZa0a/yluauDK4/SavlTTdu7MOjsdM
QLdIoWhW10vKKzAUujebDDqGU/311cCR0Drr/5Bs0uMxSOUqd5pcA0XIWAWD8yhl
pRd4zyxyYEGRIUrS7YFzm8V4NjI2Ll4cLA2LJH2JlusHiWEKXGpVZVoeAZgmVpQu
v63R6NPwzMFwF/m8lrUn048ir3XFS4F6cuckvN5PvNn8K9Jen6sYS5kJCrJQ+tx6
taue+tjdAHd+ZhPfNFo1dIZ0y+0XNkuRcxMDcfsRpUXdh5vACrTOV4MH3FkgI18k
nnn/vAwXjmCDNz6UMLsE14/TSDJ0KkCx12RBSG/6Q+FBtsIwEMXrGMbSuS6PFIXd
7VqIWasLVxMF7lCI43A+u5Jxx0jeSwLDLH/a1cDjDWOT16V00pFT/iokeP+odSZ7
0wfKkUJUrtA6CbCyx//dHTc2iAtrhV04AKes9wOzYhI9sEia+5AivwT4O793OFuy
A+zkeGPkfeC+3WEQr32ia/CN08NbyrJmCv6UuxRiMKaLvGPtzwdHq9VvMFHUwL/O
QJXB+Bl4VldzovSrmJmjw1U8o8HKCaHcQMLo2sfEjVEASw38h3ZyXeGAWat+w1/K
nxnlsOnOpdC/YJ38Rry1eWTmsQ8kfgeDSFMzgNuw7jktxG4cIt/OsaQn3Ppuhp8f
J67W5ybc4dEPxBs+b6760ONrdS/DVCR8CrNzmbJwipW1vNCAAHhiRp/uZApWqcLR
Vyvgqd0wPQKef+zGRvEjy9Vww4cPY4le+mmUQTzOnM9qHJvWZkReAcbWZdmG2GPd
wXBlqdHZjh4/j2Edtc0t9IZXDpHYiz5m22XTCQP3LQ5o10AdKNedNta1A44bX/z6
yK3v/nXVyUVKDp0xJNKgVWm3lQMt+mx3syxfDk8lzziu/C0KOk+hv6YuBcbfcMtN
SFuu70tRxgAIAxSrD4VYdNDbCIZtT4Np687rguXP1x2TpMDG+C5nnqh6KV24LdXg
Sot3PbMV1g2Dpl+BnEyXiVS4hXEexYONLJhAwnXDC153z2WQmFPx+c9Q4RtyvRox
z0nmdajRqiEUabiWjCqqvArzW+AR30yDmddjWsGEgQ3B18BX32keCTNjcH9ZFZG4
/B7/+U90E3a4siMd1kgHTzQlNT0BL19pBd4y9oVG62h2lxEmSfrcy3QOCAAXKCXT
iziRUVh0A6nkgzew4MvWbH1/+hJoB3fO0wIU57K+FomVP4mkIzI9H1LhCnnXpn5P
DNr0YDHa1+BU1OC2/5k/XrGmyEFAwUTnE+mFuFNllPoDG/GGTwZjZJIhoSBNprXZ
fTuBhA7p5UJGjA/wusTomPrY+Gz8fgc49TaQbDgsOOhzaI2Uqm9j8pCBzeFf7/Qi
B+Yln8GWAUHfqZrLOiITAaRB2F5RqcMGKutyH3Yq0JPuoOvR0gP0XbPU/TqZ8dnS
hlwbqLI/OWnW1rvYE8rfkwZmQ08Bw3gq1+4dPKdCPCABhsEEH2NJxgcNttdNkUc2
3CURUnZfcQ/4cdRLU4x/BB/ToHqWnS9SH8pb67nqp18WlwAaTdn1B8yS5G2dTlTy
4WmaiCBATPYqAbNOZ+3D8UESsjjqPCT7SxMlQh9xYjjRBKrzwYqrSgYNJ2Jo0KGW
dJm5vD1225Awvx1pGzfV/fe1mSo2B3Gos3WzYOpGZxcX9W+oj6ko/8MMQYRMzDif
35rwQrxqZsVm6jxAx5mLA/1RwpCLE7WtTd1tRMD2Dqw6jjyxS52uN6rKLFmCb0lA
uVZXaSk2elsYSaKmXwJAEz60OrlWKWcHYPHVg1JDUKj86adwnMYow7hK3z3nWYva
0G0j+7UncHeBFB9U+Tm3Uc5TQzbUfIMIaPhfzV5TvGrPlpM+mz4n4IpyutAwe8bK
tOL7f4p7HfceKecSmpYBEu8wGZcUKxxD8i4DQEq/zlWEqpVCZCqpI5M1qtOU4ym+
J6S3dCIH7QvuweCp4+no0TZ0f7meyln3kSz70C56fmu4nPRXTo9JDGPk1nuVAafN
xBuKO3WUVMAk5HgokGekghp2WwRl/J8p5qVJw0fNBZdUJOktwtURalZdkvRgFron
ja8EWHrRUoI1A0I+RuT5uBfZzRWH9PEo0n/ugsHrSC0l2DyGM+vEI5zLX3zMnO0R
7IDbr2c/O8jc369h/O5cgs58x4RZbZX0nuJiIiYrhbQHpACAHFNlGr2BjJ4eWDRz
ooba61XuWJV/acWhfjTzKyrjgWRwY8AOdUsy77mTpxXoNkSYpEUqwJhlali8bBDC
SmvoIqEKqfqZaH3XvFq5S1Up27FOR1EtneI3hKvV3tiosddy/uuQealReQScFUww
NKX6SFwzq0vhUNlzjLTNzZriRSAY9cYMO/CyD5bnAhiAdGeVQJsylOxfZcygA9el
atiGps95SlaYIIQ0aL/0gL0q/7w8p6v/0EfYUj5PxtdADyxfbp9gSUXIB9EL+sox
J8Vdb01SJ+C6HnrkT8GYeafukCaJRAVFfraNtKOSAaREXgcdUMFQ+DppDnEvaCrw
8scaiK/12Q7MUtoF3xJayUzId6Svlv5ORpJfFbnRUD+M12MNmDoVmb9GXZv0GxSD
g9Hwh9vXJIrNvh0j4zZIOm5spyFXkfxvB7AYwtQFVVXb0FfgfEuI/gEtLkuce57L
IJX+nBeBPBy2uvn6X6QYv1UJnp/f9KZu/DGSAhjP8Vqtoj29tkuReMBNLqL/K3Gb
Pc1X0QnezXRyM04L1tKnKDCOIdqyy9yfwHG8pLR+7Q8WPAPC5IDqoPLCmvN4piOj
apDOcSxjqL0w//NKZy/WY1Sy68pxpm4eVDz0u6MDi6QNcmBweLHmjPTSGBWMoP4D
PvP+Zw3j+leO/M32z95kdmNMnLME3ixgjvMMwYhI7hOVytZVvd0fs6mKgZSUmDJn
CaMlWeUB29IrDbVm6vnmFO17E3FfTSDgcWL8mJgj13++3lzQvb6w6VI0WW1A8Gsj
7hmBMpZF8P7+BEqmzIX4Khz0vBjxr/bRYiQV2h2WWHpsFMKxpkk5PFIdpsCxmCUr
zrPerRhPw7//UUOWCMetbUM+mlxCjL4i47GNGOQ44xL5w6Jemff9AfwihtcXx2pd
zDpiuO+ZA7LwNdg1eMXU+hyyQR2HZa6nV4FPGbALHCLkiZbtjybACTiy5oYksc0L
ZYlOuFmI+kRTllULQ5UubcOTB/1aSP9nj03mcy2d0jXIblAOv3C1XYv2h7lyTkIB
0TDevminxQNvUjq3zAwDnzAFKiDHOOkLtoeXCLfqMaJYD72wtfavacBng4i3pGI1
Q0Z4eZb7Mh+U5QJ7JE2o7VO+c1WwvTorjCsSEabI2/QsJrnCcNRKpkgZeAN0Coub
60a8uS7s9phpXFlVkuKPJRafaU5txT1VsY+cmrAM+hbGO8JlHMpTKRh7CCRKN8o+
Pu78SUSyG9bDbh4EqjOcHpuJkkanYElvc10iw3BAb1xfsLiqVl/G7s9Jmn3O5mS1
1SQOfZYhhlOcgOnv1xVls6lA/1h1iTks9nNNkRciL4EePOVHvU7cvsdjzA6tz2MJ
H/9kyPdWRc78siu0Y72q7UYXysRGp54HA1XeOYnU57B775tvgtdz+Hpm5q4g01qp
e8LpqHQZOMZ2f3uXJaNVRpaY54K8JwsvDi8MO/8bR3gCuEcJgLr8QAw5fBhecX8V
iran1brJN7p8vuMz/9u7S4nijEticxx32pnWkESXn404fSwGYK+jAywOxCraGaw3
71nFTuLGzdp3Mf/2YP2n9Hbg3nohu+sReZR/CttufBHHxea07z318BmY/rF5O0Cy
KOfCTBpxQWtpFcnMcemNvjOotx4ujy5J9/dxh3TgYF5G/MGxPFNPiFFPG/iKMGt4
/OS0P2dPUdUWQJOB/4oW7n3Wmv+DUYqqS8Im9RfsUvKNyQqtOBG8hBAIdCMyeAQz
pdcSYwJjbv7GD6OPTcQ7AFiu8IDkh0MXupVho+9EMkUQKjd3vAgArLkW81wcG9Nv
6iguef9oDLWfAa46Pl2x11nM+yKc3Ejmq5+ZBamvfo+aY7CldofBD6JX7s03JHHc
US3Y3dD2g91Sl8V9gXGg/TR2F7QGUsxJzPA2rp1WmEhdSccbT+Q3to6wbbEdugCI
ogobS8CYBPvP7UMdcWysuYs/H41xtRzYVGvZ0Zjd5F/bNdLbBsju/iJidQmexB/u
vgBFcsWULcWw2WhYJ6uZOaSdwcwV3VEa/VrndByIkZ5qQeTEdLmVN5AuJ5SfiKH6
pYV2FYZ7UlYUFyhCvgc9NeutS9Q4oQhXSmP4oyJ2ZfZvxN0r0e4EZIbS9xGig2YE
g+2qBRgTbQttDzRFzvWGqA/OevIcx8URzr6BuvjPjb8utvR3AxA0qfUhFEgmvsIA
HwxHcUv8CqPnUzeqcjaY+OXvMes6neAWZ0QkxR19p0LWTxuSqk9bYsrXOsn6Eogt
OmaGuZ+7uHpMVcV4dr/P4J6iNdMobh+a56MpvY1zH0hDGqNHpIonLtLu5zGwz562
ZlzNr3lHeSURDZ1L/Slr6dpVytZO5Z8DbLdyQHdTsvikL3QJeZsPZmLFiNhJpKaX
dMcMs8nO0KsmWdX6BDpvEP2Um5yuvU9XXDeishMAnNM1bte4+K0N8uf3mRIjdaYS
Y6K7rmGAEwPhwf6E9Jy2O8LmGs3A+vS/vToEOGJbo0uSKKtXO5LonV6tL7Wd483z
w8PDnMxt95u1O32rMMtTygeILpBr1tPa14oaxLqBM2aRa3PwkXFEkdq6imf1VgLg
wn7cAhCoHGXoz9KuXbW1Y5xeLEBmw2twuIlaB6lnRnyVzNUUh8vz/OOp2MltHkgy
IK2jxPj5XpY/T3sI4MRuaigMGgcFJTwLR/7ljQlsoXA1MWCBi4el20kYIwQiJ52F
wlaccncspftuoLqlxG+ocGlZFZcHUKee/a4SfkdzSyDc9chZDqjkqu/JAo+nexDZ
WRAzTe3K0fqbDpIBnLOhj3QsJTCNAWzXumW8nhOcFWtlFV4B5DDEcOwNrzxbBWKY
oTtEonf5dguPGTgLS8WYFOWKX75Q1Q2w7OaBZTTUkEXFdhegaGYntniF+G1oB1t2
E4sCMLTvJCSTlhvm9d+U6lWJdqVPvM1SnfZWXVX+Cfv37cvTBIWb1lwUIndY6Pti
4QE09KS0ucziohadwdNWzLeKX6LJCBCQQj3bQQSfGD/XqCAPriBYrrKPowoqcenh
8yUCaUTSmDSWeoHUOJbn9phbzfDjR7Gh6uQ6EsC44ca5Yj2CQL4FvSER0hM/IcJd
8ATRMlR4z2mcCt1bHI1QVbdus2BSorwP6/NjMfW+tkPDo+WRhW0ts7VpYFMpVxjo
vFuLmcR5+2ab3y2ZOg/ob9dcELL5qFvDF20fYHHqj6edWUdYAkGdPeVJUEDkasMs
qWht1xCXyft/KKmGbeR8h4pR9Oa2rdsQDQ5I6hWoQw3bFm2GTmzQYt659EAEQNBd
1ldxfW5QHOwO7N7Ake+XDqN1DpOdGumCgbmdhP8PmSZk8zGXorRj0ARdNV7ZRFwZ
Oqp1OYfQAghZU9/vCYxHCIprrb1KZOZwhymTCtEeULdVI4PWtX1ZAyL6T21nKwWt
BY+tITc7iwHnC/TY+4JsLR6QrcSe4t2bit+nHHdP8i9I/oh3ZqNTDWu/fHjpDPvF
fqiUENDvNyqXQ81ehnvqcjTI51DJiRI4F4nE6kjOOkZBfNltER6mRAmqgE4fk2HI
68Er8e6enmoVIjcB2y6155UXqnn31VXY3wJP4l1y9BSGZee5WVbiarYB7dVkFtsz
XNuMa6Ps748FdfERp6xWx6NhOGiZGdHsRBJa4FpAmWYC55nDXUgKOmcEn8XEVXdP
invKzBLwMHABT+YaoszBfxoYAF/7EKDOeZH53pGAGJoCpok1Y45OTj58stsy1VbM
eJ1tulGTc2U34XrVa2LQE4lB/uXCaGPzjcsddtg/sqQoMIXYznHzwkrPCxMxJoT6
Eho1WiyVQZrv1Sn8CUytqWgklIZSrJ6dKLd2Gse5Df1LS3+E3A6OENM27VtIU9gO
ZXX0QS0g7IVzAADqQqF2Bq4F9VRJhx5N+TfPWk/ko2kgNJsyeHc8EZpZN0KlM4n7
70gsNMpSBKJlBE3ptodIXrZJsa/UzX3rL9SdMFj/qldYliNRCpokHRIg2RLb061k
1KZ38K9Jh8ci5oXCdL0xkXMTbnsXJsWPwIZ0V/lUaCBlS59E1YF705M1zgLQwj+N
BOILJhmpI+TZjb56eywNoh3VW3OovWbGQ3YGPHLiKAWfODtoakvgi31DleoP0ZD3
7OkBDIWrxFSZj2NSQxoVeJayO0ZwQOhNUkMz2i/57afQnbea8u6x2I2I2tObwOLm
TGJ2CCt2CPUgMxQZU2xtomiJKH/WzTioAyaxxusuk06XPN0HMq/rI52kIsnUgPwG
zqCsKptsXnhDeIFH1r+7hegz9dd3FJWKbkmdy+gNR/YnmDWodEoCcoUFYpzZsv5j
4AlXm+mnZjVtgevEemsQXOgSwQ6Ovu/qm/Uw4rZkqGpqkE8jdU7RHnLsAy186fze
4kvcZ8KITDYjc9vCXKZwQ93X7I/l1QQuhAwrXLRXIoM6v2V8GqW4nxEVaKRaGRrX
dEFrBrfc9GSI9CSmUsEMQ+VJ3VurUr/biKKbzFeTsuLkKHNagoIUsqw3V0Y7WY6+
GWk5OaLTNtZXKJXL0qSa3v2oD2jpoKCsre7QLvVM1+0lO+23J7xm0l4wHBp4Vhms
MxsHvjypaNT4ChN8jNyFto5WfU5RvZ3mrYHUymVO4Ui73HrJeCOdXbGB2gbpQSRN
Ll2FJiek4Qd4QszxTp9026Gd2wQsCjuZ7exqHTiPrCz49WUTN5dHj07ivC2WMWuX
F8eb+nwydxFTcXl/Qc+I2rWyxItz6Kx30h+Q9DIQxarDiMygkmYVJwkXqRNXkBoL
5ACepfmvjOjzwghEhJsYD0KRZPtEOwKEwfp2uF/Pg+YZXPQUhSzuBUnMA24nH3TY
al+XD1xErWWMsJWr3xobYSkZsg4VXwAhCKN+EKFXKNosKIBnY0xQ81cQWmY15ZSQ
OS33G1jYRO2L7IEcF7PjdeOUJGNhE7bNK1VG6+Ih/u0jxSYRXXrpDjxhW0mKA/AI
mupcahSwQ1YEqw7Ufuh2jXdXLx8oiTKBR8jHP+i7+bqGX2PlgypQrh8pQjRbLdSX
4VPgnlBdNdhY5FVfJJ5k4/S5FHloyqVfmQi7Oz+gr+FSke5fzxjth8zlW/ERCMbh
ENSQ4MYGoCOH0NVbYV7gmYvuxbtv65fglgATJgLqsgaLjPiDJTyH1/jC/cpZPhv1
Mc4vCPELD6efUUfTywzZNJZRI4w2SSkA5fs+EE8AS1v4Cudx8/Rlcfv7SSsWcMwj
mTSkkK5P0ps0Iyg+U/AJhDECLsUPIRq/yQ4e0Euh6lv236dXqiTgb3XKGrcBnteW
cQzLGxBSqNhcww8u3QwpW4yjiO8ewO2E4YJro+j2PQOOtou/pZaL6WtmEe75jFHk
q8FzDyz8YnGGpSBu+/ma30JfFYaOw75ywAzEmrmyc9nrhK/Qd1pFo2DElLTvvOk1
g3U2n7idOwpowNfUTEGPWUhfwm/Q3xz3G8jKcDV1Rd+5Yjeh0VtryzmM41ZuFTzN
HGHVYnq8Aq28jOYq0g+h9JmB8zPGvEtquedYtCwWkB81nr8RjP8wY6g/2G2n4rZk
X72bcWPIqOnPsVZ+qLYE+hbVgPI1N1Lyd3cyTAxDjDaqw9u2HIB5Xq/hZ613+bSq
79DTImqaWdWNT30XXgCWiuGJCEgvLawldt3BC6nTynKDiQIxqzWD7t9Vw+tTN7nj
A/GQBb6mxpCBz6ISeur63QTRAljW/nwdKeogDPTXHD1y4crAkGXWKSNoz03Rfnrc
MzP9E1Zw8JWwTYBB4336f2v1Qn8aOYCywIA3HluHvJWgdrnhlL8T8zY9m++PkWTq
hia27EaX+7IpgPoo/J50+nGQp+CmC7bVXyBQuEftqNP19a3Ezw+jSzKvGRJkoGBC
6Tt+Ll0etKgVds/feg+jf/LBV5YWshy/xT/uLeH8UTFFUno8P+8UUOaWSvyx8uPK
21EsmjioHvbQ+To0Vj/7jsSlQ1/eVM1JjE3VJbQvOjaRDdn9cU0OcohdWY17ZUnz
lXzAwjFZ5NxNxnXcgQQAMTCi2B+TTxBRkzT8wvIYk6HgNu53YwkyDJn3C89RpFWY
n/ahxvlvSRmJLYXKMJ6ylVjuaStVi9HOfqx36C8m18e6arQMTK/hLhpiSfcV5dIp
YtfLY06BQL/bxUAMN3qNRKkyYxaRnPT7ohCXxZ4VL8m0QMD5O6ytQtV/0zDo69hT
aMOaWxIUxdwMskqpMOQ0TX81J2YwfV+62sG9bC3eZt/meTe0V2fSwBorv+f0aC+C
16TBodMv6t6cy8WeQs/Zgw2pm9XNcgubgjEN+1TNwkHKIbdC+ezbwbShUMTOBvoG
hatlV4frqqE0fYtsT0SpukYlpeAW/yy73rL+S8VuakwMigXxpyVt/PEGKP+ZyuqS
BJri2h6lXwtiQWddEwn9YRwcQh+8F8s3nXB1sife9gXkc5nqCwM8srE6hmThMMJC
+zn5mG5IacuXjDwxP6dTi3YBcRfebftFJRTL2ClcRXdGh9MNuOMyUicLFAFNpkKr
ErrxBhCbeOw1+JiH31wBx4XaX3/ohOrwExw8FFjJSuo3IdMMLhKyoaOXe5cca9Yo
Ll94tje0wH/FxR6yjujvbi/aIvSgu/8HJWEwTvbFvpUB5XFLXs+hEgy6oj8Mh/cV
+6BbRnnmrD23rjlyfY3SNn5FAdITUrgUxVa0ooAOUgBVAjG1PTmYFQwZ18f4mvew
VjI6kpCCQZm8yVx4VyF3ZC3bacw9et44yna6X1toiJJQbJ+0fJfISGQwmBMwuMBg
rrYTeEF0sipIBmw4UHiIQJc5btaN+96nh0EO7VAmtibBYitOVL8h9LDUxkoiPYcI
lmca+qllnXq4VIOOJqzypQ7PPrR2GQQ6kSmaw57Hj20ckZZk+jiD6Gy2aLK4rekT
dzapAWa1ShWu8TJUe2QadPeyzhnTHDYApFGa1dY1Ysa07qOgtAWQVE+Ie8QkMYLe
rJh32Q9S2vQg1LQPIpfgWnH5NbcSlIuTcGxbD5+vu8DA4s6XgPSZkD6pAnhwcCI4
R91jZvwfD2Q0Z5cJXYGsf3hnM9Wtx82FkKJuIXTAyVhH4aY2hI0MxXqpamwdf48b
oXA0K8tuoR2Xck8yen+xOxzc3igjDDLxguIxavjvoFQ0IdMwk7R1BtqDwbVr4Mi1
T74Az7HbW7V1p1AisP0SMpXca0qrn0ykjhl7ecrmeiLH/R4kkeElemT1mcxTmytB
/tcLZpxtCZEOJ4oBEQ7c18ktZO0RUXJ8IcKnyika/72d5ale4pgjuJujS7RybMKq
eiqX6vu+xUzQH0LNrdAaxXF/j10uYojvxkJ6/HvSA1wH7ASv3y1/02WsAYQJ+m79
PY/dX2Lb4KX2OGKnD95KyGGDrEbvGnz2IOU9qMUPHBbKrm/tzp+OHsqUzkvh/et1
lJtTdAXnPS55fa0h3ZedbHwyWa3Cb0VmwzRkUhzTQUdu4RRdW1DJ/oMz5k9PFJDW
vM/Wne+vhUIiWVGmWgrXQcMTb1zQ8CbIW8qPm09ZxsZykhmkrewjWkrcmgzlccey
iPR78q07vWQ7/eOGyqn6Aappbdo7OwwAh0LOnyrjHNsOzbcQM7umWguJbC4/pTu1
ScbIc6K1Biy/+NzkD7XauYWYdQb7QskuAv10vNu+Bcj4YLqy+raDZq2RmzBGXJC0
2LT3mUw0grlIPE6HghbDAwAFhfRPREpQ3HwqZ8mxYbl1tsgxLudpgo4lZNCEAUsB
OqQUY4EzxWtbGv4658IQ4i46ww7YuKVTWWKMS4Z6IzAsDgNtoylieBSiel02JXIB
IgMIxCocqlzhgI5t3tSVyO97pc437OFucW5WYSyPhz99c3CVbwdG4gldVxYrF2Lb
tB3v2q9oq2w1g4eCLiVm0QWrcBOje6MoGWsiCUHvgl18wwlbEy+npKTefYGhY2+y
3wnmy65Ep9arqYexw8GRyj30DszxMiFf/wectzeKk1huFOgecIhmcNf+pDE5iZIS
Ekr3aBD4JlmAmSu1CEpqKYjSbMY0rR7webdEtabOjiNm5R/9zp/7O5T5QiTEPrsr
NFTPBnmziASYrYqtCWDa+8Z8R6tVNdY0twzoDActbYHAv+PZhFcsYQCAeaA+b795
F4vlm/xuhhVYtLSj7DzhFvbDf3T2M8Fk2hwLmJOQBkk1iBK1GEWJCr233LJYWunt
0KIdt0QmWYMhX3dEy3GW5+4YCLKPhYyAz3x0HWo9H7hAGJskLHnEnYXGZTdTb97M
aaDCjLN9DotwouOp/WxQq4NAeirWtOFjMpoHIYKi1OnMyeMSxPzhLuSdXfe56aXf
DwPLwv4RDC7l0vTjAFDtrNm9jf3hjX68lk1ka3zaRYBrWAfdYXXCJ+4yFNE85dN0
3hNKCb6qqFRvu11vuoTJ+8xDzD1ye4kTDJbv4phx4B0zulH+GcyS/CKqDsdRPtwK
aF+QwN9Wt+GLLNut7VOZcQ7cxl6HVHkggFpHETB8UlcrcG4IbRIG5VPyhSRje6uX
Da0KizmhjG/YI/cFOyB5tH+rP6odYmrFD85UXnM2cGyNCcrmoOEl/ZuvPsLsQkmV
6K7eI3SXNr/H8bI3N+Hrh0zsFTBxbvoWa/eYFClVioBOFajRJCJqGGH4ix9vefx3
9Qj46W+k8Ax2cc+tIRYPnhuIioJeKjj74FfLpgF+28SKsu+EUq1CjFsKUt2MlKyl
1cXjGdOFVjoz+4KSxCUCw1EnjHGS43TBXof74FX2woF1bg/hQ+dhde/MBiX6YyGI
5wd7fw/8lQ+w7saXD886sN+eWigcc7juKNeqiIykvoNuCwymHK3a4GaMKcv6mJKl
6Hz5kAIzns9cSQhQtA8sRx8NgpuhIHsY37bRtBW4yT6zTAg9uqNU3WJoVYBrKgzM
IVgA70iJxUlNUCUBYVBM40upzB7bJUxUbTidX7fMcihs3boBddOoJLwwnDlYfeIg
cXZNyFESFLG4nN9bRnu3pkOIH+nukr17pAwOWCd6a8OCtHk5a3hKCsW+5E6j80Kx
pVZshjRwO4LzLj/b9xoJo0/e3IINtyx3kYdhV3oJeNokgW7rWuKB3bhaHXOv9e4A
9BSCecqJbaD/S7SHAM/90ndU/IPhwHndfy+GpOAOpKdSXwDUiWVUvF85oWCSenFd
KxPiI/cfM7HNCE0N0o0k3rLJqI3dhIlHgF+nyJZKtj+sTOxTUzxNEhgwoposoBCL
6oSX7AOD8i+my/8wT62AOqZ1QQW0hsYUwjxZMVpeWZ3PS8zFplGDdXMJLU/hay5N
P7c9MR1ZdS2Lfkhj5yyHi2tzq+Y3GzGQuRSlhdB85BN3O9Eiqq6kqnXxSH4naLO1
dd3ZkULxf2gABKaqEpmh+iUREkeHD3r0Rb1CTMMwVLFHf8UIv13Piq1elW0e92hU
4EMRWliWp6E50m4IAoam1pVBx+aQ1iUcsaugJpienOeqraf64NxqKDWn3SMRLM8o
/fHlsdrqkFmjn5JbjYj/mHaNYEih/qhcT8LHE3yRJnc1cvmPBgEtjwK0jAPjzOmJ
xlyWi7agpcrkrm+Uso4FVuZU6ifQzyJhd0MJG6ci91xfaT5QCWxEXjOdLn/4ovVk
xflpEFiA75+B0tW5YVOl45q4HQxvzmX1bdkZnTzZ7/FS5PA6wF0aiE4uanSu8OiD
mIk9J+nSfddTmC+laq8DrhIcnHggpDXwjagOYAqo2CZr+VNSOEl3KR86T/aSvbX+
X9qxKHTEnXeN0Fh4wPDfpJBdDcRP4CBen80jxf+Pfd0aYwfYQnGPJeruKDTw1c2c
Im5R2aK5k3GTvb5nD3cdVIq2YgoPgJ81TdcSLUJ2DU2MS3AgZZDaOcZdodMi8MlM
Fmu57C3fqBP+aK2syQ68GhOPpNBGMzFV9yaYFFqsPwFdvQzrpD3yiXbDdO+l2aqv
pRuL9UQv8oAyMBKmq8TyJ6Fjf0BI0f0EoEjEIc0GGElm8sPhc9MIs+ZokTcrewr/
SzpGvJpCRUzT+7bcWpcRS6OcKZH/AaqKKHphRUogW2diooijastC3fDET7iHkYQ/
aVHK7Py20Cn+j7j8mhGRWu5hjl1AQQ163cwMBMBbWXpy0OAegD1pvd7g4ROOHKMR
klJtaDgcgnObJC6iN2qK2VbBIfEXQlWj1OBpCf6knDZemUue/ppsRkk6IWiRLN+0
0cowATQIzwJhvCp6nRgwKFvxBaGivqu9B4bPcLGpsxDmVzSTR9fgl9SxUC75ER2n
zBTiCrR9qYtnfgLnMJKidsh9xAinaYbEAla8Rabt+1N/gSZ41Rwq/S/VERr0CxiV
EW1w3ZaLX6WBcZKQKJSWvbtIUAnSIjAmXVcQ8yPZogLPF7pKybHj4k9IiRxpnqG+
N1RillKOcpsiAG4tC1Ejblop4/ph8t8H3NWW4TOrzk9t1DOT7KvESo2cKExrqC3D
T4CVzFyCat/0fGLG/o9RpTVy9epJ7JUns4Id47UUlYf6l0GbEq56t+SQR4VAp4KV
3WARqwYcS7lY6iWM/QecaiNydxgKb0TDmFut+1wne9vQtBpn+iNXjABYY3FR/DOT
fFcrMyLYNrSVW3ZEmgCNcdng6bZMUdBWYdiooKKEAlwrXMt1ZmxR4icovsQZD+g6
ThJNjk3AaggQdgv5pTq6DRnNpFA9Hrps1mv4csAJyreNlgfRnUVWvXLHd9hlphEk
ZhbjeZQzXRvWM3oJrTJSaQwgzgWAi2s/XzaTxNv1lNGr4fQ8Rq+j0gSfMC/OE0d1
tU3DfWEj6FcaV21MfNNpw/8KefagMgM6xqS8su0LttDUs0lOr4eD+Fs94rpA1Xha
RXOchAJNHrK59oh1z9Cwk920KjQS93yVUiPx4Z7eGp/6/1EcsZFFj8C3SIsmhT6F
t3z91c2T8URdJ6teqX2z4l9y3DiuQnl/6lQltiZWomH0LXgrHtJmN1WDBT1KoHVs
ECEa/s93++Xd1PabELG6uAy7V7b75P516tPLpK4XOUEZ3HxpezrKj6FUC1oH4Y+3
qLS7uuV+EcANTQcXRRfpzu9RMzCHqVXW8SKTXkAefNrqj16OrTsT+aHKENGVsrRk
ohdysIlH/jtzCkzX63pj0dDwidNyUTDohEMac420TUoKhMIYugo5VQfh1CAFDZjd
pbciwfNwb/kdoZ87K6zXTEXm4Hxf8grkcO9blRJTaZJP1iNTOsFlfGW5mHgt+gOj
AgQoxDi1xX5Dpes/KYzOcdrt8pUK/TVH99wJcrCaesxXAbvyzIQjX+g4PHPHEC9u
TuE8wDaVY/vRGVLQyOv97D/kfZwfuvtPHQc71sPWmQwGipKI87rqTPWvzW9EgOf+
S5di4NrkPO7DL9mqALGegkco3WFh++uCWSX4PuXK4SfejvlQEQZo4/Sp3vxn3zOU
SLkbDt0clhEBDqL0gyIdFobk1CAa6bmaU7J/GjGOaqHctbtvRIfyzZBrkp+HLUeA
46LaV38irKSz5cuizk0yreIquLN1VZ/5tfLnCS+UrWRRTRqnU0cb6sUojbHbg0PI
Qi8RTZGxvPZo/8qJpZdqCkBcwmfnJF02iRKif9kM/s4TTM5URWmqyPDKy+zZUhAL
ofiZY+KAMO3br3MfXBBBm/2NZZqDCdKoNJEP60i1jRhY+BoQDzlwt9mhG5O/1wMD
kmmytkHHZ8xml4ZVeVZMQOaMSqagsEUHEcya0nV/VHm+7xeV9eYKhuMcAI80Wt41
lDZ6HI75jtSewJ8yMpeUWcverNLRwhTU25HohXEj9uCcoEO8pOpQ8N5FMprWO+wC
7MbEIZ71FT8oIUffHk+a7d/CztYuYUQ1QIMvYNoeaX/Sb36rizWw71ajrvNCfo0M
NXzSUN6yAzL8OcmirZ3PUn20smXghULYXe9ij/AJWnyCsySaceVyCPDC2fI//1XL
djToOIvxZ5/mh5ErHd6WiTIPaw/TWWd2yIK9Ckq90CX/WKaFikaNwr+JgEU39T6z
TM6CgkoWlRVmOVRdLBW1XulyHQ/HKXYNaD1cJp7yyWmwOxuIxiZTfkIG1i7i3npo
kuUclJ5rQb3/0OCawgqhZZaySJyI1wv7ZTK8LEwnofOtKYeSE/CUD14xsHoWSQGj
iv+FeoOH0GEHMw/pFijws6ldGI420ISsrl0xducNZAivm2WgJhNrwbX2p26g8YY3
qfVxqHmdhtj+UNre7QzI/BN+V2TaQMSUe9lu6NJryafuTuPRu9dRtr/cZt2DztA0
kraI7GOHJy/aJJSrHVMJJsNz7WWc0U6XyZ0cAkNh+NJUaEPd3nmm2D30PowGdbjb
WRue/wK+sqStyrNYyldnZx7g60JolLMMbVSJ2eyO3/JmUlAHeVc5eeh8o3u+1ypT
F3wDpvxxecDGslT1jS+mME2mb/QKAt3eHBQooaUTuNPbyCidK6mPQcYW266tSWzb
3q2qcLJH45Yu3U0QEBLXQf4FSd1n+99JETqlZT88Ad/DxUM5+/n5L2GskGgVTiSu
aq4lohPjHVeyFGJ9xdLcwaEu7dKzgQVkQszW8ecmSu+uL6zrGTV7kNSxYBFqib/H
xCC4Dva+gYWc0RRLk+/j+u7KVm+XMuGRndPZZ1mEwm+//DHC8BcE0iTMO1Kac7PG
n+pOqzkSuxU905JJsDNGesI4norfPzcquv9bkLUUPDJgz0vF04OPivr/3RXRuYa6
80ANgMzrNwBknFidyEYwh4qp4Ctkbs5flfy4KCFHZOokfKv8BWjXSEHX/5PoxFZ8
52f893WxXTDp1oNiLSHalMYaNFpTPP9Pu4ghH+rO+G9zINGnIHjDhWJLnD9aJwIw
l9izpaivNP3IqfkO2vR6rlXLSi8neKQNytzb5QJ20jHArFpci4hAeeDLEXuRbcSz
nsVclk9U3/k+Zba/dZifTkS0o7DcgXq/zt7eHO8vsJqLNL15caRoddZBVlSCu7R8
gOaZ7LuO7zsYnwQ/8rjN5ZXXtJDByCfTYxXJuQmPwi7FEyCyQkk0+OBbmNw6/Zch
35xKvdYDKMI1jsvx5WecUi9EvUZcR3f3OYlp6i4I65kpbzE9UFTKhvnr19vzkYPL
mh5OBvnLcAPaftmXqK+3YryCenOQz6q1m5CbrrDFMzPxFPT+VOUzDz5jRaCdB0Hc
A5OTHsuB+ar6eR051w++xAHufeMpIyVom6i63euzL5hilX1FcTIveYtZuu9muEv8
AZ6WrT4EMwoZKUtUDR+S8XsNr9jUTNmDmI6JMCs7SZ19xY4jQS/00mIbRbKMHLVM
43yFeYO26an87xuDUA8oyQUNXdQkSIs+BGxWksiTNnS5sGSUc8m39aX30JvsFg0O
t3zdpnwWBeM3PRu/RJyfbp+ZwBOYLnqXukD2dUjTbJUUsEZ7vVUp7AXB14RCD1/8
oX2Brsm26IiPaug8xZWEhhD7aMOWlzX/AoR1lVlACBKqrw8lI/43YTgE703BOOkK
jS4HCxelU2cd1HvXvmmM+XbFzErDHNDaWSthUtnAvQNEAxY7n6Dgvxk8exqoHj17
Lqcp9cz379s+DcazTshGNhVzVf2N/XmbW+dx/Ex5eohJrbg7kErlCvpyihug1OVj
NOK2DxX5kcSYGbT486uCih529kqDq90gQ2jH8ZOoiZIgeA3VUJ3CzgwVRx4FGivZ
DN/lOu/7W6YERoxcYeYZ2mDJVduXsqe0s50zGaKjjOS5i0tc0igS8ZK4WOu/HWQr
1iF4aPWCSdu9EI4LK6DLUmsxIlNuIacUdZvD2lcWaWqED/ymCcBs9vhb9GSXv2tL
rOaig+pae10uocJm4ALviPGLfEBkFrPIkWJXRcVbMGe7YE0ws9Z2uTbSqOkE7nI3
3meWmyTLhOIRUyE/lGzjndc+srM7z4hDGC//MBFRMjllPs+fp+TZKwZAV0J+v4iD
M3tVHE7S8HV8+2qs7gVikXHPTAAYDCe0hbvOd8Ix2LDu/j76sLttRIQ6+R/9fDRO
5nmqnKFKxpuQ69O1see6kUIyVkNMC1nBsgMnam40ZrvqwHMKyv8um9dWqiw4pFe6
u0jQvxJg7doufkhzWIP3L1D7VnXiLZUuE5fVhDPz6HHbglYqpSE4Z8Gh5cIhXbnP
Y7cAhR6uzR6X4JFMXhwnOQLm6IKiuAhh7kqpYfhSiG+v2jlsS/30aXtCvrGQQkjl
mImQv0ZyAgPp6zoKoCDS3yzS2gUw4FBpOZFxWGFpRwSLvsEM/GBAAnzLfsAfCSPX
YnYMbJTOYaRYh0N5+6e0o7/+qLGycJtL0i/Yo5SrhJbPhPP3fTavo1QVfaBelpXe
ORWJ77AifNEWcUzRP3H6MDSeOP4bRAjxFdAOZ3JLUDpBIb62hRMQS4m7oplVmAzA
mlT0uHMEGUpP2LO1lV1k9jdPoHMmKCVPguXlyrGRGeqsrn6rxzMvUgGSlcxa+9iC
l1rMIer2QfKeyLHdKCeLdqlXerPv/hoIc4B1NtUaBu3u9rS46fWbuk7cZ6lEhS/z
+5iZliglYpecq6nhmtiCtIOTPaZasrPdJOh1M2pc4cC9p//s+V44i/HlE6kJrad3
DU7Whn1ywi0ptRJxr5hr/OIx9XPUb+nB6OS+vxqZSe3CzvoVwHYCFTNVImTl4i1r
SvhmIoHAVlS2Qdg5KLMczmfX0QgXrI50DJ27boveDUJzwwQc4AXpVcqLrBvb3OBB
UuDT5qGQuva/8ZMJp8SaOuCD1PGVvNLzHHlT8h4k9hUBRUL7TNFJOd2pK6mtCUuG
X7+Ne2Yp/JVYCM1C3qbqZCX747dP8UJmbgsqmxZE+StcarIo1JyhAb3DAuAYGTUM
Fc2aMNicr13wPG4RzX/pIzkDq3ecRbhomTxAnOMYB37LWbA2oAmLcfPSf8kU9KMr
382arQjlaN6V4nHGxCzmURx0Cs51tt4D6HxXGX8KGyocfxPQmThF/bOf5ROp4/Rf
OjhMTBkW6dJKKXnEdjIYCc+vy0a0eKarBDes1VXnsiiVwlwSfwtaFRb52pRH7e4u
k20aQjHcVPBqygDFDLtx3+LoqHwieChwa9Gc2efUgckIRe/b56xIm9f40xWSPYJa
OLm2TwU2wASQq9IzsNPHGaXy0GsDbHC56CdDQ+KMU5LojNDpD5+QIzrDZBy22Tub
j1M+i5+2u31sJfvQOq7OimTgLRwl2h0RhulxPhS4rR8anhqjVq/lsDgjqpdjORj6
V9Fa7Z+UmiNbC5siTkyQtSu7GuZpZ1jFkaaYI7LruHpvNQ7DcmJpNoQqw3lZkmhv
Oh/zfBJCJTOu6kgOwju6DWewLnxh4k13NLQGwU0C3HbWeS7wMuQ1/W7mGnwwrkKi
Z4T9LQ6vcI4T68YcnAy+dA0s5zG6ru/EbpQA5bjUJbfJ8FCq2oTHqgo4Cbp/OOde
AFf6DwcddHGbDohC+BdrvVnlZY5AIFSoeuf0WZ/PLda4pJuRqEQ6OBPUazUs1c5Q
Lp1BgcaWvnqBwCMa4l8U1nuFG8qLnmcJX7E93ak2XG4lpSSnENZ/mxwbGeb+zyda
XojVmXl14GlbuH0YJQxIRiQrcGPpgDjwbv3RS2PH/73sp87U/ON/TIJipKs83moY
byQDSmuNbV5nKqQ4NdTy2bF0MEg61YJHiPb/YOBMkMcfYq0Oad10jzgo/wWyyFGk
QlFoVNUgbHFX90EARUU9SyR/zl12N36dKMFywi9DNyIOOZt3Pauv42tlUSHnnsCV
d+lWPGhOJweDJy4AiPdvRef2ZULELNNqQXQcV10fPxk5JvH/u0aLb8iiZeBvpLLC
FqXSR3h+t+jzcoW6RPbHkhU+QLVaSmf1ZOwc64HhQvFvzkukyyqIM0jBmR6R1wil
N1fMOD2VdSmaquvX5ucaW+RwKCBOB0S6euYd4Ca/sKX6Wtt4M43GYQIGRXxUKDgG
HOqEM1uisUIK3ngmpQ9Q5bKO77ZS9QO3zzt2tXYqxRwT16T3uD2s1pR0dCVwUL0D
0cyNky/OLG5SZB9JWl0XpBpawATp3N3zmUCOyvjCz/kkd9jyCdATxGmWmVYADFzB
jCAw7lrupogUct+8ssW1vswU7PwQvn9oUZlljKYqhPxmkPPV5G6WsWqLbTFkJikk
IX4BcdakMErp/IUnc2RT+gt6o84FzZ4XcwP5bGIEAnGfQrzJ9fypwwhmyUjec8rX
vR+F14Emj9AakDvIOaN9PGtskbYXk6QjOku/+C/wr1YF68JBzS9qBx1+50zmnfRW
X/yoh2LygYzPm7+uzqtxjnnWWI9GeQdMAFLs214pVVOwQSrBj0+wC0FJGPKgpIQI
Wrh/d3qtjIgUNkPZM7Dp0JGTV34BfOeGl3QFA8VVJhoBMLDJdOnorWF7brsXbubd
VzQ7v84zjIYMhNDuURf1W1que8GfbFUbS1nAuDR5LmyZOd/tFJjgCVcvA/UNbOez
8nienQk6bxYFpBVfHXHAxvPXfmweMgs5JRTlpVc42934zM/sil7zEu1mx0gxhNQz
5mcJ1JN4B+PmfZj2X+PdcygOEMlsf1AGAURZ7GJz6VdyMfxP7eBlMm7L3F2waV+U
0pxupy6zfdiUu9tcit30uoDMJsHNHnipchmWPQi6XtNPv1TCWGDU/3uBWe9TOqd4
MwHM/Fw7IChcs6233wa7LAsTDSpdEP/hxQtFPQAQZ3yQ2agbrRc2aniiBbaNXONN
oTLJZaowMfU4ISlsmWKh92O4ePUGFMg3nl0gM7vIrXTufWRR4+U10ph6iiyxt3sX
wgGhAWkpFs2nlZ8asa7rEmYPLWeFFOUkPDTMoborQspbyTRKxOWbCwiGBxfkD1p2
Zn1V6P0vGEqWvTM87UOTIY3U3Ch2q4yIKKMAQBI7m3CWREjWbvmrNsNZOKlF8K3f
pAB3JEqaW8I7eU8Ia2gqKyqO248BqAWKkKtYSkuv4fQh/C9D3vBvmhQlkBLH59OT
3XTDxV34VCTG5YJkZepl+PWv11XMCYAZfPyTDOkVX4qxZUcPdYtFTSDRVuwFvqcZ
RWvbk5a8JutIvUMneBxZfzGrFAij+vGlxz87gmn8/3IketE1lB98dzXwmJZ5G/Lc
n6HbDyDsv/UvQ+zBJMn4szOTePR+wspBfXhADqQsF2d5AHLVfRRsHHlNP1k92HJ1
4X1zpNL9oh2ZRm+tvtQeovkzjrR5Llg3xIE6IjZ+X3BGkhN5/EpgqHau3x0yfE5o
Ht3ggXJr+MzeP7/+oTZb3QNvQHbaUinR5uCBbgezhAQdA29zdJf3/swKK+UqnbZZ
s8JHvnkLm+ee/2Pq28vFpBJ1FfyLRGYOFporoGE1DjI59VgGqkC61zEQIqCxW9gD
CFTr7u996Jn79sk0lK8QZHDWvatxHIz7cwihSPNqY04TBs2sE3dzejG2QRtYgnya
V+tYYA+kxnaoNsEQekcQ6uYDZ6Yyk+4F1pvf5OBoowiaumFKM/Aa7pcZ4O6g+D8Z
lDDKpydVyj3Y62Pq15uzEJb9GrT4oEo3G7KBmSHJrJQV4ipPCbtAzEE/9yFl04CI
6m4DJpAIbUA6MRz/Rvj/GQUZWvhjI7SBlqhFMcX0yEv9Xx6hz1qgAAffSzfdg0Bo
rNfP+eTwctHhOlZQpMboHI4QiWly1I2VIDDxK/2mle3plgOaBPJsnGS//JkgHD7D
U41Si31A5smh9bYrc2guMVs8nI+Ek0NjQqnDJf+7S770E1tpjreCHd2XDoqKAS77
hJl6kM6sOVZvJmOWa4kCfGoA//t1XfHRQkHojzW0dGdSCMyC3u5NgoIlP9HYbq4Y
d6t9cSCvR5x0vXalGh9s65kOcgEahJGCFLIUmGk/9R28It+LclP0zEp7C0OZeT1Q
Oa6jsx1mo4VArpP9MqWlTQUFGy4yNospVa39pZMXFo8dtyS56So7AI0wo6XUtVCZ
PoKSk6bsXPZi0z7s75X4g1RtHlrb5exIBpiswkvbmwpXIfkZXC4sA0jv6VjRG1vz
KSPqCcPqacfmr8s4Mng6iYahFViYdPQUz0wSYDwelcxnLyKxLhkemhjaDdls1cUl
vKlESaixlhsiL05bvVj/6SzuwtpYI7KUCvYRIZR65BbYCx/YoKCfAVwWKKemMm0H
hVdQpedd3/keuDw/VnYpJDRJ1ptLoilwr/67mw2qm8CiYrKHtsGhQXczBm6Tffgc
NoSF7z2nrb3biq8Yp8l8B8MMx+JP3KoqMAxkdG30rQ3D1gRSAe3nVR6Cl+HNTPpt
UUKERcJFXOft2ZuSqcPTnO7seCOA2BKk1ofFm+YeXK0Mf1x7Fw4Vn+8JbfUuQl1Q
K1zYESSuZTD4653fcYMwkId6jgdPVfOzmlE3cgx0r3mpyWnZuV4bhHCCcho3FD92
oxOYUm8B7ap+Jjbx1Et619pT1CwopjeBMd1h/xaD/NOpPT4sa3InSABncU63F2af
igNDCY9IBAn/xVDVYMhpAOO5wWR8Aw2s7P1MsqCekorHLDMp3G+NsUSwrc3TabBE
SLuK7oFTAFZq81gCNx/s6tSqlqg4jNYzf6WHR9rySiy0VDZRsakuXJHt1OvO/0IN
i7gUpOiXwcVznYU8ypz73PqoDotIvIWKY2eDl4cmve40wKoYf5vU8UalRBw5BXhq
wOmCix+JrADleLfui9sP2Tm4qCkKPOnDID6Ir5gvOjC1lqA+7ak0mObf9YQgDDq1
MIVC53XA55+kFuE40bsAV/H7wwmfxCC1DTTZV6vTXrpNKYYGHhm7LrjCoftKJ9fR
CkxJma8hDy4xszkXJJNWenDkJac/g/lWtsAa4O2moCjkmDrRcMpd8BmWaM13c71e
rkpv8kGcxbV4iEB0ygFF+HY6ky2+g/ceTPzl9NxKH3Nd4Rh8OmQvwEoIwaMNeLv1
per7yVNWLOgNWOQqoncE4ag1HPpYK+jw5TFQuPFLiDzvWBwtrO8NDVISEhWnwLkN
H0+RmaDok0KYUSnGuWtKg+ZdutLY4px1fNX16BFNrhb0hkpRDj4oK1I0bm+rDb6g
FOHrTo7XxaMXZng2y0RuRNuI9fSS89AYUEKyM9cxrG+pNur0iAFmpjcPN+k60jPD
G7lHagPnDUH3gGr+pxqYdkprPnRVUD0XaYtcPIxOJEqDeqX0VDud3mADL5U4dFql
JoPXZdgbWSzB5ZMCLvos+o7kuIXV/gvKz6vFXdZE/VyhTundpBWlwijV/FxIJANa
0ySB/xT9cBqDhjZ+bgRPlaVC5FUA8B7dmN9yOJoezpIl6Jxspd1FpgeiWT5jNh4D
8eKGxqgzSklMMUfGxc/1hOR5t2c/guMSin4/sLmQiKzdF1NwhGdML6yDLbjNz1V2
WLDhr6FBeDq5hDitYsizgOGJURa/PE074XAPExaYXvVKkHHJDyYBpd8NPlU3lJQq
zzXU1uMHSOaxYw7uL4TP0Mzdk4QpeG93o1F0OD33BmjXqB6Aq3MyOXt7DCuOONWz
u83EFg/RNSuZl658Y3rdfcz9rjsP1VYK/uXoxmYMjHJ9BFskep44/XVkrKnNf47w
FWK6S3tRG4CJGg8UbCGJ4tsSYzNxpmon7wRENKW11P1GDlW2wUq0RU2OswiLjrW4
VjMwFFuvdG0lqK6sBqm14RRxSPXrFVdJ9DhWdil/5/g/1QzWNqNf51DjRlpKqdZl
eq5p/n4MO59aOPNSezCluWb09MUA4ziSolkaUHoYcZ3sgQp1QaK4o7PLGqA3EctQ
GBh2yQ18kUagHt3mfi0z5bmgLH0jidx796YW+VYDMU61HOs0lJfD4yoXQFuqVKgA
hHHajF5Mf63iFlKvFU1SBAFNASij+MXSlAJhsC9fYfbTFqQ3IE2TobCwsxe4KrmV
lj7XDhp+pQzCEVR4bW34NJPOErwm7QEOveUCCqm6a9LLy4vDPXuRc73N/m+s+SAh
iR0MX1hQdsCI2zUfMkwmikUEVhWN9aCqPT2MoTltXR0bPzRifHsyl8ehNc9Dhhgz
7jLHqZC2vkf35y1j3sQwD6wOvKv5lEvqY7feXqQfX/ZFJXq9V1A389JADq12TJz3
jfjY+CGzQF9UfabJRLHf43A43A0Lc2OP9XyIhyFrKBQoLW0z65LkuRgy4JLDBz7Y
aSWrS++vGWug3rekS7NG8Hp20bb+PaH07ozcU7DQTngTAlsuWlFcE2baVkwp5tV7
si1fPoVpvhfd2tbRVf2pCDqHNRB9T0VYLNblgTXVtFRuXC6Ttg4/K27w3FagFLcy
k9S2Rql8HT5YSYQInALC33URYQgr5YgBJiyGBA2D60OXNwEG6mSbnBMXrokCl0CJ
sRgHkGITdF15sZ7n1b8NuBnTU2cbBAzLxX2cJ65wifqTuNrQe7dNEqCVBcBES6Sg
JJJZMlyAQuCR1Lcxtt4PE3giSM4tDD71zLk4zzdT1D1xaPLBsUE4R+C0+IgfJxeG
+/2xsHC51GOCLILWPxhtMTuAVJY0B7Jte+p1WrtLQCOT8PUB7v4MwIOfoqlIsWvh
+/IBIAbwASGqc52Ym1Vd+TOaFPS/SVY6S80xWd3LsSqQowLtXgai+t0sKNk3pPGh
aWqPXTWV919fXNg68dR3h6ZHTKdrxLFnqffZTwAojMPK24HMMLEMWNG3BY1e4grl
u/LCsmquS2Lluf9Lx15/XNJW9r2hOKJMzNIpo3hq+Xpr6cxvkBTFchaR6dAHbnI/
Fow9V8LSUs4FnCrDAIfS970ip3sxfPlp0sfSpVQh12ZzLiMh3walW7DQld7z7Qsm
FjU2TA3WLLBZj+2+aZcdOQ2WUdME8tup2sQZI+kw5gJY6tGjMxJy9BhM2x0nnijO
ya0jQS0SobHmJs8Br42IYj+0pD3YVAn8DtCYPAWNHkW6ZBcwiNa4kLRwQxaO9+3O
yHTDeICeaHVK/X6Ijh32NzGYMIFdFW4gklnVfk0FJMnJthmcppSKPRGnAl0BQZwQ
m1WiqVwvGLpCvH1Npo4oL5NmbsCL5a5r/Ouhxi8gl0aVmXHJE8X/sqjXuAYTflrb
FYrTggMYd1fG/REclK5SYr/ecODP0RYdSjrwpKuzGEPbDE8DdNR61Pw5d25RBd6D
oqHQY7uAdEDN7FPKniXwXrnZnK/2z0hWUk7k2dhcWPQC14+HV/JjOQDKOWz9n1ED
rH/1byM27TU88OcEmJWunwERXCmaMn+NyKzK0DbXjHlEJMWnvFOEt3YluVWcl+YV
fF7NpUuBset2htwZKlQRU5te353glfsMCHCMPGxNSLBnwSRY6S/5Xri97HRe7S1I
W+VWDE5hlxf7gjBA9n6uBO+VOcgKD69OaCYP0E3EDoCfSgC7uwYEpLXfiglIJGnF
0M89JFz3Iitq59G/nRwXR17j/UCq//VqjxJLeMu1wd95uX7W1Aoa+6wA+4npeX+R
KmttdKVuka/Z4IqKVJqXiH5/hresubEX045se1+X40+V1NKN38iN0gt1ALd7Vo3b
T1YxwaZwM56MMohYUPH7QnxnUzbp7EwzjIGxaDkT9+HC8yPnCPauZq5l6ry3rZ3S
ogLv5QDMQyf8pk7mWWLk4EcebO3ZLjTzNDXzPZgYUSJtUsadxfs2RZ7UmATbeZbZ
bCZySZNcwETUUZ6r9Dp7exRedu2/RLw48d2M64FvSLBgOLaL0eb/Ysg2HWZ+YuMk
c3jDcgT6Ktdxh6zMwGqvdMEQckwnen9FmMkdKDG3fgXvR5DKwllySXoJ113PEUHT
hwrgj6bSNEXNlUsBMHtkglA64jYXjVWjixNx01jubcR3lBQ99kmDyCReCGJkXqi9
L9efvlgLznux/7yuBKo1XDHlwb2pZZ1E8kvC3aAHiKbeCPg2jXc7xpp83/wtu8kD
Ke2MZiRTodON345P/w/H7+L/4JEP5OPsKpD7BHs53V8QBvxA8uMBFe6DFL/1h1dZ
hyBlNe+13CgxpgKUUpJ4SEvJIXVPBp+KH5ivteDo95U1CzBGnkkKZOL5h3IRQS7u
j5QyTcv6QA69O5YhJqy8M+dq+dIyjfu3Gf/r8O2dizRyvRCUTwvq217Yh8RLQtxW
NJ27F0WTWZgdg/3JDu1xf3ra6BXyTEyNy6aQARBQVt7PN4FVcRDUz2a/E8E99hVX
OUkyzNwGwsIbXyD4sLgNifxAnkuOcfpWZhYKrwAjWmcb3V75Wfvr8F2MVVCOqZrW
DH5eH0jSHgrHzncIGiGDXRAbmO6FI1zr05X+mIk974Q59a1YdmhvPcBj0hQzzA4e
rjG7fpHv5MFnKO9wyaxVrcTHS3hZIh7rl0vXWBvajm5fcG/anrYuH+4deFFBVefl
5/yhzpFRHK+YatpNCAbyfbIryQUQv/MHe5vL8wF9I4IoRnFgw/vaWEVgMQ9AukcX
OQsMnkTUrKFGgkoYZTGzrdb8FT8PXAmfifEjg+VFuQ1tpP/pcKyKQ5+sJo/yimT5
+EcJO+8+ileWnNl1ucmEJJzLyni3RTeMfPYtTt9hUW4K8eTjuKu8K9mg342dOkNO
hB8L49luuxzBKVHVZeZq+B245GiyucnexhQU1VpKtwA7ljywraTm3JEO4ZhxNJFs
9AJa8H1FmZNL13z7WjmYnCDnauriwmLIU4bncVdGND836oGN2IWE/zuOrgrz5fGc
+qScoO5eaE34V+Wl7+ApoDjfgF28BichN9vI6pjrIRefYNQTh3X3dU+ArbEsrLm0
GCobbjqdGvRHZ35NdAnnVjFZ5NNtHtvfgU3ZG/+ONCMFTgtve/EkgHR7NdwwP67s
zf8Pr8sjHtObGPnO5FbCBgNsaUygTtvsjuZGtHl0z/L+F6iRRtfZndmEv2EgjFHC
3uebPdeEBsdkq6jvN/TekJyk8exqyCgX6sx7VertMn2Kmg3AmfEyT1YAhD/KFZ58
GiN6utOYVJ7lx7+xYu5ED2FaDZO3es2ZgJnkXPr5/7P/Fu8eUSlbmxUHcIRUSpK7
wW9VjUvNp3YAlDoQHEDUcRAGwPLnrGTLpCGDAyaKQk2998hoIqBfscVGzYgGmpYK
Si2HIaJlgtfKCkuWQSXT/J0nJSNx8gQGXrOgVXWzMuH2cKPofj7IPa7YqCV1Aqgw
Y+xw3kpBF0ugCwAFDKq3Vu6iT2MrN1Jgv5aOf2Zfb7mEV1ZbKhT8asOjNLub1tI0
srUkesij/lf+Y/RXakIANyMXxUFnMAaUWei/GwrhE8FqRis3XEXZRh8/aRGAdHbc
YAGSYDmXAULK0DWqB45VG72T07U4/FjC9hirNFgqp+qNVyBX8jow8LlyD4ZqptNq
r65Lg20Zj3MDvveLnJZ47MJbjhilUsOqsjBAzRIza1CWu0O0MpoPgzod83nXqdcL
D8qQTRV18v1wtrBSHFEksMZURjqkUScWLT9iG6cEN108ASCvdnwVF6Z8Jftul5W2
OwmUa+2YflWBW1QA6A//LcW7kJsi1FkEjhP9d2k/Pk2Y2nopOnBN7wJSB19vLGLE
JXmHIAeOICmuwI0JXeO7V0n6d+ffmBQ0+hZ/27QkFfunSpeAMJkMOjK1RJJhRExL
KV9rhgPuUfH8RoEV8SKsCWNsPb4cYWkrubbKHHBWQ3ERJnV+M3vDJMjmhqa4DjkW
Yj31sm2Bh5xZH6IUsqAAPK1C5oyTIWp1tgHUfimNbTopnQq4RGNuJJzVgdroZ2eT
60b99kJ3HTG/X4uGLBi/eIslIzFiDMcaj7auwwpQ/eJEKNlW4Auw8AabgyJ+Oxa9
IpaC0kfie/wmUGV21Wg2dP1WVOyLH/ZjR4aUFp9awml+imiiwV0WlkGHEZS76LWg
+eLEBQrrT+MBGSLxOQZ/xIejQF+lvXaJ1NctHKv1s+Nw5RMVHMIO9L2o6GuF2+Y9
IsjcrmT1k8z+WqRYrr1XqhnI3NOKUVXPyuTWkiwThvCwqJHzsrrHkcqbH6KFlLBY
QWPl0fG65VU1uHy3kbT09B4nkCB8zuhactSK8+YMz0Hx/e6J/80INZwQoMLJ5Kop
OGJ0o0PSs4SaaDUpkTuN34PIBViKSt2+of5jQaAA0lVL0GGtpSRtXLW49QSRnn17
MA1FOPYyNIKdn/WYZZTvuKpNSCaCBbIxnzFZnZYCw6Xi754+t9z3+Djd3r+8+a6R
wTub0qaUGYbyrsURVOqZHWz0ocxs39bxHHRw2uSPFT8Sm5uOcVIo7/CywCilWrT8
P/8GmLcMQssk5tXGdtOhVNDy8Qv1itTu3f9bSGRKQiJW6+1EW0FsrjhuxKDJgVW4
WCqO1CB4/ha6Tz3aZ5Kw9WOZXlcvyZ2l/OYnwLpMwpzvaiUK+WudjliMmJvX39FG
Ck1d8p+4Z+valMXDmZ4FbOO4CoImAF+sB2uixQzveyERExd1RVTnDBMqhbEIcRl+
1Jlg3AgN2/0p0J1K+jIOuLWZYX/aGQL0OhqOd8cOT72zurOtP7xKZ1KOimiMjNhf
BSiUZfSQzMq88sIHimhLXDsUEI34IlKgkhCeq4pbNyTD4hCG1Fh1D4G+7Gd4Y2i1
7PKP+uOkjfFeqeYim8y9kCVL1mSkLETjuR6eRmCJ6AJe9ICZRiiysUMbRXlbgaA0
DxdGlbYmU2MKsIaWjbFgqTlUao0FiqgRjtmZjAiR3SrkjdHsa6QhAX5b4hgsKp3Y
qFdKyvHFjdJ04R4OU2KpSajRxIrcNeJJ+PHqB3gwLCnL8BebDBR9aQ/zoxcgNnGp
XjTlEpk4innHSdzwOJDPckd55+GCyaR8yeOmAQYMtiiWOobdwpI8Tn0AWO5HJAmm
9qW1roM3pXaKzdIczKtqW9yCwlXu+iO+sGeS5wU6Ucw8ut7CHhHQMhU9PNTU9Uq8
7XXmE8wC8BZjKKMzFRz1vneHGAyLwfAt+W5MBQD7OFEzVsynzXeNhPN61Qw5ktQQ
buScvQlces17T/tux7YzTpjIFnLItxVKbrtIkkvR/HcRx69EnfL6amjGNtQb78/5
UG7uSh7np9rzmZchoHbZ3cU5WDBXjiYlpL4L78wsbi8xtOyv+lgHGipuDpA9d6ZR
ShXum01njn/aCCqKtpU3N48/NSlFGO4TTJjTJwwSAjJLTPldGGmIefpkcFiKP0zT
v4DRtL2nQpgoAp5xiTUYRTeOE644wtAToVVdNBal1101Ai7YoBbTazzck38MYGGr
yNzltGPi6SyCLm/oowFBRUy7U5TE3WqQEuDLI9LDIvl8GJn87KgYqwx9t/jHtCKd
2COliCpJdavH2jOa853JEhmfKk+7IJeKEZlacsSXFjB0U/LQnC0+DOlRVneexFTj
Jc+xk1A8C3hSJuMuucoZ/dIxZaiNprPU2iDSHG2PPVIxL+V3Vrf5PvfgXvrTkHNq
xDeZNXMLg8RGvG9varftVgI221L3UXGhmQBlceDPyQngWg+I/OqHx8ypEEbL+NZc
mc874I6F9BBEm808E2U+b44Pp8z05zz/YPOAd0oZRuVhXayPUefjnVe6uBqy15wx
0e7WSqZLQLvJylMwgCBGtdwqZc8Zh2Alu8BXbvQmNmVRsruEa/8oln8gb2ODxlEj
8HWk3YWSVZwOneNLozTj/KXdV6B7W7e16vWGdD/T5JSM3YBMhh0lvQjtv9OM9BLF
JQqr9cfQBS0lAAZyxKd9ZZN7b4TUunFO0hJ2S1boTQorVNKYhK2hHyPGniNJ6kJV
S0YVg+X6ugdRl4i9PSNEVO7ve24XrajTrHxrXg/AFYSwNhys2bYURR70eW4KHD5P
Ode9OqwNPynYC62n3SKTt8rdQ6MgWRHxVNXb0cAkT6sbsEk7IGhyzXKM2pPz8UE5
+sBPkJJLqdz8zRoy+u1ujyBtaKBP9JGKwpGm1C/IdFMwAZ1MZpE4PEQ+jofKcz5p
S/cL2ELMnzLRcWpo97aCYjVN9SLlYPgKwsQP3QZJ7m4gykzu3wthsI84qjxXTfGZ
bWJ3qQtK+rCBrdMZVdYGGamWGB6KlIsijtR2a/lBCiFW8PdZUWoIBwOCWC1ModaU
wO9+xHvppKBAXegzdkGHlVU9qroqLyhYSXi75sRy4wHikNBrHI5voWyYuyfl3T4/
1Yo98pZ+o8k5A8pcc/JnpszEanmRXlqf87ve6vHKL5mCTcF4b98L9GOARjA1OTnv
wc/hUt5nCa9uoSwq2fcyzVndpMaN6gP/TKpl2K8KZGt5UV50CrqLnIDE4sFa4P6X
f7ldQmToCZJYFw/0qC0BUxF5cR1Ce3pwQEnDfR1uHLrgfT7ER0rbVGJxM83XAVZ/
rclpMNFDoAY93hbfDSvanEkLfW+yehKf2itHRrVFc4jHACBk8eoa/Eosd+8NvfkN
jamRiHlcqmYn4AngH46A7rGIgWu+/HlC42gNJAAiFZ5Cdzao5CF1n1GHt9a0bdO4
2uq86NT8FQLDeEzW645/PskqshlAgZsawle+8Lw9IVyHKXTsHTsEb3FA7HMSy+Ym
lmg05OckIeaWJli3GFv490TMfPRe+BtrKTa7AIPdkBCtN/WwGT8q6EJyjeOrIpCg
Qk4VwtEd0/Zq6+yYxcK2i9EV2ar/ArbupAnfHgFYsltDsujkFBoaLhR7JKOycZAC
AiNb1H3uXbeN5l8qUznyF3HmZeK3NJsLQ3xD/wke1P1QUv65jHPZst6VxTJsplF6
w2zOLUS82fQZOcsFZ8oCY+BJh90lL+yefb/RF9zmprhqEDAMhSqL9WJQIZlE1QiE
GYON/k0mxZBpVeT5Nh+k3FsJeAOx+y5ukJYjAEt6Q3WO51ZHG9YkU2LvHasOu0wo
kw2ZScmtY83m5fP3xnQTGLr4W+AO2l1uTqhXkGxxmbp0sC4r0qpfElvHNAtj4Bog
sFc2RDvcCOHn/YWaaupdJHDmGvj8dXWJDhVMcrVg4qyFon5dY6aNG4CQS9uXtQQa
ASpRoVvAQofZ3VDc8KJa+ERjx+rcEZvAxn2BqlIlA0bTLvNpFqfr3L0PKXwHf3wf
FXd44GdYIiPvLBu0+8rKvR+pjak4n9TD1UQc9b85mHFx/a2jLvmqjkOSKR4FlAd6
Y6VkKTeV/K/XVYzRb+J5bIXwgpitg9cHFMagqoKELFB3JoiH49FRTgEwrkzBEyo4
2y1qVZn7NXzzFz70FfM/buqCzyxtxVF4ymcloMi63oKGFnEwJnHtyaUD6FFMI+dr
1DkTaSsGbWOBsCu7sTjiypgjTkjYJN1Q4QvgvN8Z3q2vNDW8shQpC/Ci2MSh1iyX
5W2szFobvM8SKr94vupUAiYombPNNCXkFRusk0vmS/gqxAkpgGaBrw6QQZV+C9Ww
uchd3FSBaEa4lta9LOjqZr24Nh6RdWMVizn3ZZQqeot0+S3fYb1ro7ZtoLITiHX+
n22FU3uTUfxs4NBP7ml9OkuuOerj565LthrLqSIXKQytzdjy2aLdRANe1HY8rWdZ
GNLvJnIbpe/BCb98B6xhe182rUmvHCMMO6wj6QYdcciDCyYf1x1bb02yy7BzeNTc
XX6O+0/j1LLhIQSoEaF/HOEOzSi+qRTw+8oUbVqXeJ9idZveVXdcb4efWEicd3RS
t2Hna0SE2FzATW6nSYesR2m8BTfaII/lDbpVs2mcnpUfVNNnmik4uKtXkaptKcjp
EDwoooufOHFsRVCDVQWhaXzHlBHsmBTWPR8rYQARQF0VRZhkApfo9V1dJ1N+tUti
GlQ3LsMk3WIonI3d0JS5FBIiTa6qN6wcWnKL825EEF5HpZpfCkyGfVqxvhKGDgZF
L3UP2PcIKmgoUGvsanDRmVEB1Jf4luLUq5rtMOB8N2dTjDYihljIZbHIXyqzbpdx
ZBaePPelN95UFT+gSBF4UDawpOm/jUf2sn7lS34zzWcUbrI9oxUg3RtzOQXrNdyX
mwvxAT7E4e9vEzvrNiki8V1wenhBlZQY2dTCEIaHa2vDYM+UMMzaUqFiwpclrY9b
O2JcF0zL6yvTeJRya6eOuhcoP+giJ/xhEtDaGbttRMjJzHgEIwPuwh9k/yzXMRLZ
z+tWs/CHIQLS6gNiojO3BqBwYarT98oJ8D65Iu+j5CX2Jyg7jb1U2M/xD45J9E6h
zL8cwo7LbFmO2JkKsLlmec0OhQmgsq6YpbnyUL5Sb/nqpwsNDbszWBY5Ytowy6tF
boXuTDxGP+8vitzmUc67/CbG2Uhgl+Cgh8H5u0Rp+5tlIKCTVINPu1JjjiWdwGGF
klNhsyEkeoT8/ZiNTiXAMqgopTnRXyzSUtXDeul2HJOgWjlfIvl8p0kAVkoR6Ico
D3SSNWtDdImpysuBKBK8Xyxc0ZV8/zaWlHvgO71GiZsoFCaMEPk2JAUdwYFiBwXz
zyB6gXBYe/y6mbPU4mDbWZKpbIJ4lRP/dG7pxkoRBhEyvPoLxeZ8JbOu201LLFII
OQ3Is/+nszReVieiyVER4HMAdUmSd58BD8scHP5XIVmjmu6/VE+IwL6QxLbS6pSg
udVVi+ahc6FHnlUuvedZ2AotjjMZwTDDKSRgA5rbbAp8mAOvaH6kd8xL0oMeygm6
MeK/3BRcmp1IPijgp8oSlIAwXARoi8dFjfj5XDdWVD/rnSMDsRHDd1vmj+hh1L1O
UlBqtcimzy8u3cjQ1ezoS8gskbeyChWyTniVmkqK9Mdi5/bO7X5v8HOLTokFmdgn
j0QU/OhHvb16dund/pF+ha7FuUKvVqTyxJT0mrqieglKRBpz2BApcSK/RcMD4uNz
6yKN2RnJjklP5w+qkW9CgseVNfOC9v1NPo5zOn7MSsvUGmmR7pNM89z4/A/ij6HA
l3r4ciXjuNlpud4sJYabNKdGYVlrLYxGxb3RIlLiSOdT7GusOn1G7A+2xuzdi09m
HWqGCbKCSX2HZqbZlEzkYvsxOJPSKSwm+FdFRBXtKtCRUrofY0nGiC9GFr1shJ7e
KjtxbSgNKDKj2vS9zaagnv+aT4mzfgkui6MpUXMiG3G3xPogfWgaRCSqypR54FUs
BpNKHzugijR6/IkfZgmhZz0KXbFY9MOAWrW1J+O/2vAgwPw+mbvEd7B0tt6/PL97
7F8/kBRJOnfXx6NbZGC4AsbaAY+qJxdjfhMtJZd2rNQaaEd6M4OBXxSHOHFS5KS3
U3yof9hCuBa/e7ifh1rq95/72E2DEGOUuuWghq64lzH/R0+frX+EMW9iOfmbmWFP
qMKTkmTmLhshvdva2/YKyUj+XbTcXwycxcVBEYbqBJEiOkQB45sEmn74kl7yrTLx
o0VrtSBiXFBmdMCnLpV6QPgxejVwWKrp4x0wcJOh/ZbGvXylyYMSUAMcDF+JFtGW
kydYPCVRU+yZEJ2WmRbHOf/DpvRwdhE6tuXwACX2e6otK2nOF3kaGnGrto1cIWKk
kTE5coNbHjXE9Ic/I045+YpppOjAZ8R2Dq4Sd2D85JMLdU/OmscFuc82844VeChl
3gVpNuZmp2QLQXQyHFg42rXuGckM470u153QbPEYkrJVzFXYHFvXsWv9FXxobsnR
m8A/SsmYhIMUzZvR8PvaYvWU0pEJYQ4xIp03b0NuTB8uFH6xJQYI0SMEzfEzQgag
bddmVS1z3+kLvby7bPeizu8ITYBYkrATNJC1DEfmcgnJIdadGvOQlbgwkUaKzL3n
Bd5CWmHJ1HFdxrXWqazqapjNG6cY3dRzOWhBPpacaPbo9kazNvMuuUKZ5/+IwgsH
7SPapUhuZLgxTzXOoVFBRt/6FFfilIQgy148l7aqkZjHDG3XUU5+sh2Ak6xvD1Bl
HogKlw0D9YoKVuRQvKnHC4e/t5JJ8PC/A648zLY1DQNpL53ibFU936iGKssjNuTR
29+Uca+wg4+/BfJPkJEmNV5t6Sm+wpZg33WQXcNcb1IX6ZfS2c0q7tz6ft3HpkF4
SPBW+B6i/KyMX79jwuJxmSHt0sx/DEH7YSHndKK4qHpq6PXiwvYBePKENyaxUfFc
9uCsZBDEu0kGvS5cRqiFBTukE51WoPy6xKlaxsqFQiGI6DB9tQhF7S7sXlgFlyc4
9v3Nre9y2wgizPblkVA3w2g5ijXt5DxDdJ6V/2arbtXtn4fpoMYqIx5CkA9x9hMn
s5t/zq9kKekBGb2BGETxCNYdONxTB/hEEyrJlHNJvfxbzGKIGMf1HlL6ocm1TcCr
Wr7qxRdE+KFAs135RJtSHlRjnZnFim4e8hzjkOHCL+euVitqv3fv3Nl17kHQyjHf
fAZanUKydhs7Zp4cAyYPEUHj+Xw8yY1qLInCtiH/cjNmig2r6L7ENkE9iS4mZcHV
i0ryyy3SYGRGGb2jk0cP5MQaJ2LBencWBCrpLpqWSkijkrhP+XLkANpbMrxXvlrU
dreHvdKvYroxp9torV8rtuGfV+OpSJTPnHFlqVn5yol5q1q/pxj2gqxd0a+6iXlz
NpCice8vB/kHnSLZxbo1I/nSPFFTeSqa/ta7bL/a2Gln0lnZ+ftruay6oHsmhDKj
/D50CoDZpu1Cno5aDImxK29qPqply4qckVRE6BYFfuTBEW/yHAn9PCOK6LMmOTRl
2gMcwPLIjCxNPbxC36TyBBzxIt/q99Gs55njfoYXJO9ZrCO53C+AWTHJnACGdftV
wxA4XyOyBbwBxJ6VAatE5juhJkPhe8eA0KPQgYyLiluSrBPfyB6aaZrhBeKcpmbL
WXYWn3Q5NeXIdsrjRZe89ApxBO9T+snIeonTp25sXbEckrYcLORhumt/WnaqKZjx
BFItUFUZxkqmCRR+iXNOATM/Ko0ZQn8l2INZZ3GkwGPY/wO8Qg31nbibgahM6Qvx
IiguT3m873kgAfhYlRfJ/PELzJA1G+j7qQ0iyr0wjLj2FbqOAGXUT1sv3th8fLgV
etOUwVfli56WCRy1lEe5wiAsfryVuBvNml9G4vWd0KKvkgJkq/XZUIO6b19a8cdS
X3absvlbwDBMRqFBz14khtW85Tm627SUAVh2X8H9L2AzHiU/XyzXBs2uRtwabzWG
n1WHLf5jVIJ1GzLla/JsRa4T14gGIL95e2sDPMhAoflNh4RSGXdA1B0S/OZdvBHR
3OPIyMTONYSgYemxCCiBK6IWIDlRT/V1WBpAuIXxODdAahGcgGsc1ogc90VJ4L65
fRtpvOvwKBi6ervnsOjBXqe2XL9Nh2bFukFOQ8zWdYTv7bTtqyp/bR+yu3AIWoTl
kwIdYMJBEG0NjQWxZnBABGL/bXo8nv53dEIjiktaw5okSGab7ABuL6T+NncSSAcg
XBaa8xNICkWPMGq9v+8JnZXFDK8D26HYHarF+f30hGo0bz/ijMZTr4MeH7xHpf6K
jkj8bM3jQjlOCJ88Htt55fS2TBZFwhXKg7s1IdmoEvQ6Amj5CDgqDRosM3Gy5/Cn
wpH+Qqk0rNkzDS9q+qYUM3e5xAvYuUqhxqT69RXmD4pvpsJjcPL9j69QLCp2HMxE
kRtJwHNUfaf44CaPPEqRg81UXG0gs+KassKg3+K7759u16ULVjcuBweD7mxwbeM6
AIaDJy+RZ2Mjhub93kTGGdnb1HDG9zBBCAuoWr6eVpwN1AExeD8GUoE5C0/WrIcR
iZrd7Fu0tKeJxK9tPqsxxurn+Trd/uzFhfuGQZty3rnbCqFKWKrig21YPc8phzCP
fbeDtC5SrdLCZ4EcQWsnvlQAmdA9t/jhea7xFriqmfTz8azzGCDjn3alBq3vW2gU
8CRESp9Rv5jY1SFNea0KdOSjXlQz0xyBKT81ua+PN7gwTIcxoXiaJEbIOa2bnD9l
0aTTqI+/Nj5EY8TDb+o/nue8iHY7ggPBWCvUy6Dhr9xGLeI0CosIffgIBoDcvanl
iDml7ABuPnWrw7kmAJbivfLFN7kUjarIbiaD548ThqEpr7AplFywLoBF3nnqS2vt
OnetaCNkDp/e3BWsdj2PAcd3P3bePaj1259eyPg0Hwv73jO4Li9P4oZ0f313bwpE
G8rtzJk8eSeFrfiucLDG4OwHKaEbmGjOoPD+3OYsUNHOlfJOvuRZ9fz9XYUNAwi4
3RtdRcOhaU2NaYEdcBeRP6elsq4FsK7vGnFtl961Sj2zLu1qwg6WH5h3mZAKA296
NVDe5yZAz4pO2QMUml1yx+R18rZVL4BbVmdiBM4XwonJyDB4DCkha9QuKgU9XZG8
N+7k7iPXn6e2dJVeHIzR8pUaxwPl4FmepfTs1WadJykWQfYbWIj0YRTXO8PUvrfn
Efcq2bp+Z03rCTbXo3sklS+nDKzlgpzJFCDLEv19sYGhUaIExuCFm01hSAohi98S
Kfiht0nQ+H2eDEPGYolNpf/pDsptZaQjbIlAHBMpS7/bUNd+Diwbu8uqvQLT6N20
uAxHJVMJoh2NJIIcv2Y2KyUPRCPmB7vbHXTLwBKXnVZj+m/0db45INKHdzkF15SX
xpaJVSN6huRn6Mi35269z93M8eUvuyC3Fl1Vtgi0Iyf6ybbbTKYZNxnAno+3eaPt
6El90ZtvKa3x8a5cxAR/j2W6PKFBwDo+fBS9sZsp5GxYUZeiZXx5wREFurwB2f3T
mbcQnoI5e3TH2TJI7BkRfOyzDmzfmnbU2gVr4jJt1BxOF3P4RqnoGDJrxTP1TF7t
hHkBnwFf2omHqkC7930n+IjSnqrnxSBCjW6KI8sWLagVbS3ues0SsHRhdtLank0u
dqBPMD07iId+CiiG6Tg7ik4c7Wic2YV2PEct5qQj9rUjkLe+WH47O/jpeBHMvFDL
4LpDLDI8zAsr5gk/LIQ+Mz9OJB4TWwlh4ff9nbYbe/kpD3Qd35ssflXnhIVtXJvq
iH/89tvIL7D5iTv5uV2VQrHe6VVGmVxFM2Jz5DlNAfKCzo79iwAHr4eSVoaA7RTz
Lhwf8yrjtRqdhmiIhGW6x5wKSXATAe4OzNFiUvsQtZ7sCTEv+f1KPDvh/IARDvPd
meT9paSazhkNa67qAQ9fLoSlIn5QbxbMHCfB0Wv4cz6ykhPcGiC9agTqqOOOiRyB
k3f6m/SjwlN4ctEon2xUrwDurzBwZOEj+imZdMM63yYJ4rCBOVykeUbgbfTiozmV
YLrKuldh9MJdFUVdeZD1hKBeLMn2v/B7O9fc9nV7XuD786vt8/bE2Sw262GTJ3uV
prH5Jpss95R8iSBLKQDuFE4sdgh6hNArYME/cr9YqhWowt9OJ+Bldw5S39H5E1jD
LduSXr+Kmcjl94GtJs7tMOA/EdFvjS2XXRFRO9EZEqj+0GLzchZBBAxPxMKKvlZf
rt/J/Hagz7wXGxnxuaIqBONwA1eLkeNsSnuow15aEJhxLMXY1mXGXw7PY0NtPaWl
x/W9NaJqIUslPeMoFq+JQKkhfQOc2PNMkNIvv7tFHT+M8Xach9CfgvRbgY9kX7q+
n5JqcZFVu0s0Vvf70FbaBmObrS5Z209v8uP++P//iyd4xQ0rI3peb6ebwso86Uf6
nj7HNYev83tcaQS7PZcrxSfuLD8KqgBhvaNU5n13NPS/O6wXgEHpz3Pepdygr+rN
qrPCB8rG8bPSL6V4noV3exAyOXZiGoXGgYyLAIQcWwbASdHHvnQny9pUO827MHxD
ZQKOpkTpAzAu4yFMRf9ZIa/Y09kdf5yeNeMABkToPTf7IT+w22ba/hhNM1IMSSIT
r016pDXpupeIU0jPLdf9ZhTqBncbX0t5XaF4M44ZyT3I/RXZbcQybHXI2bXqmtb5
muL9+n1d3vJFmT7EhZw0r2Yt5GbcWP3uoPNuT3GLyEF8WWOyElYTS9efLh8tctQ/
/LP2XZQamqyYtGImOqJ+1kpyMkoaIkIDtb7H6wa6r/dwiYuSQOVxjcatr5Nv+Ybo
8udU1ypDHSg15ubiAejOmRoXV6/uIhRgo8q52Q+6rVqpnCvQGRX0rARMck+HrUed
P3Z2GZt15fQtBrdyYJTDFXbWGNoCsFztBCV7GwRuZt4/2DHu2cwcPdaFeCfkeoGx
ZZr/2z97s3E+JZlJ9n3/UapfC163rxvyukkUdFmin8CQhKErLcGBIZmech9ugDtg
gU8eb5MFelPzFoEVjT+gB84CEVnhLkiV9yj57okGtvmWT++/V0lFTlrnEABhgkkq
drEmY8atPaFsMPEL6BNS6/nyvSKuERJ3s4wKqQvcfuAzIr0lml1wAGqw91CpJoCH
f1XIaHKascy5zCwDvsx+QGH4dRGifiwwkizVi1k35Z1oP36QvaoHkxky1ybg+Jl0
l6mu1cKWc5m2fcCz4bweMtOrvw1EZOqodgKHYmp/eB++fQZUfSHjnge2BJKiafz7
RqY3hkBp1x1PkpLY41/rztpH80oHb39hu5rgbWtJRowhTfTeva5pti8k2fiWKo1i
GCv4gN4n+ZEqWQPOgmlsm9CfI/U+ZqZ5E5iBJuQXNFyhM7/6k4R+/Yv6uShKHd6x
6LgmP2tPDdZwZsWMzUDjlChdDU7RHl8vIRxCzk2ms6+vRuBQCwwCi9Dp4BDSg+ss
jTll7UOAWLSWW5sDrqVuSGga6xim/7EDGfzQShp4Jer7nFKgulRlt1DbWNadV+Er
hapG39CeGh2/fhyC5h64PNQGKRCNBo/9LLfLbmqSoYDW4l6ht2eWiZ7G3CjM2bIB
BT5tt+HDqvFJHPVQ2hy6UjF1KzPVmVra/oBI9GVLWyg9JmVF2YsxqWvMM+x4JLIM
POiE7Sp2MJW3ycS76F0ElI+zX38CHBv+G10CWp7PQ5Kk15vRcRLRIm3V7quqc/Q7
S1w4Kwr1TGqLJZvWKib82DdwTRV5EBrVf42LhePTa9TOcWXi9ASy47NH35+tJ+yU
V4Hiylh8ip+FT1JESLnyznjAu9AEhPHPJsU6SvLABOgZBxhxDwMmLX36xMVoPY1y
7WW3MnDioHngdxX7AV80k0VE2Ox7ZHu0z6UrouoLkBw7Ek03f7sJBLmvo4MfZge5
oAgcEyfnzGnjs6mA1wzFJju2OYAjVuCO7+BpQ8vHHa9sGVafIOW9RxMUK3H0ENCT
65aQNr0tRPP9rDoMtEOvGu1mVzaOY1kU0A5XIjpS1PvM0mKbnrY9mSOcmGMKaEjf
oVJAmKdFRVZJBCzAw2gtRWhMhK7RENRfmv29hFG8wItyXYfKmL6AvTu99YVxSfST
u5JbEHBuiHOFppj8rQV33NN/kDeTWeeiRVc4K8bcbStPUD2a2N/Mosv0azyCa0pb
CoU1E8d6hl+h7MtKmSBpXmMecBbEdLNAczSKphXkE5iKmlrJ9+KyPmBqQW8DK3aW
plepLEKKDcH3v1zC92TstroeK8th1TVrflb/+1PaOaw6zF2TCm3/5+h7h0uG5HU2
AtnARUbaEALY4z6vt8JgdMqHDkRHwQAmB8cmFS5albpbCDVQW07K6d+6k3SUuAhP
lMWYXmcHQxrOHp6sRE7znICRxFMGBInAAdXXkUSMojOQTjYfVNDS+3XTL5kQPtQv
Y3BrPqvD02uyQBJhXS6SblcX6Y7Re/Ez9gks4CIufjn6Qs6ha+rWjKQGlzYhvPEz
O7XZTeA0ac+xnUiXK80Nb7efmdght/V7sI7FUWayV999VoEewDXNE80euwaZkjrX
fY2euRytV70H5dOSuEVlyiEOtp7tVzUVF1qQj0mbAAD9jBVVPlzQHrVg6Xk1kabW
oigzYoj/gDBfew2/lvSgpvxh6BXrJTBFCw0Wv2AhD5ub1ojZp6n1L7vS7B/4a9e5
uUJbL+PO2J5XpQcLWfDGYSyAETZ1uwif/vSsrCMFvwXeF3zspBgzqwqvxryIbHsn
K2GfjrUBzLJV9KtvzQ/gsGpuqH1ltLGfFyJHMMouMctqqZYueAngNXGhtkXDrZ+3
rD26LA7QeYobt+s2uDfV56SKzBFXPFrSoNr8oSELTh4SvZx6ub5UUVniHaBSuEXA
758TMERjRykvjkbp/8NthrJmsYmpy+H/88RRploRBc2beduhsMgE1zAhW0iSF4PB
Xi07YS/KQHdWVNUCQ/mK/sQsjTnOlEjlv20snhoSJOqiP1PXkd1VOZTlxz3ErjBi
1UH+Bzg1UaFXIKNvS6ocMbQtvhOyGnzzGMnkWWNwIYpl+X4RfgE6vSxwfwA9oAZD
1Hjw+swkStwlREaxum4leUqWf/FMfyBrMN2OMqaOUtRO1E8eP3XI5rAgzkWpiYgg
3GHP+aBYG6mLjyyWw+aZJXTI9xC9llp8birOZ8OvDsGSSfaWBg0z6lGJexE+l1cv
qvbeDO0M4anQXeKjQRS03xdS6G9f3yH5n6oT2nzHWKVgZbXh1LSy5Hwcrg4G31GI
n20kITViq7TyvuLvYh9KJ3UgFBD3QMD+ax+9cHgBLz/Fd6Wb1JkcqRvIZpXOGWkW
Bml7Hpys5MuX7KDKDJIPE+1A+EJR7BaBkMIx1bd7euUccmvGko3ldDsGdOZ9Y/Mw
9Ap1vEYxVdRWeMp3w7+L3Zw7HVI4qqL0Jq9kmRh9u/Dn71nv+NLQHR6A6IKRy06N
lFdA2mbI7lc50sf2s11p0l4snTGNDVAijKx3yARWJyA1kYvRj+aHlZSjhw48kKj7
2c7S+jkz1VWxwpM/uDaKdnBJHYsKiu8Nq0B8R8PEUiTzPDeGVj4UbY+ST4AAsH13
X5uOuQ7CkyAjxVO9vqqggokD4Evj/Rn8TqnBGGfkKOT0od7iIPCrHfMYHUoYW5MA
p12hpkwKvOM8iax8OVUWEOEDVTxGj5hf9PHlVhzyZ/OlDlYCGhd6WwnO2+LJRhkm
Zh/8LTILbOS+ejT7LiW8g96heFlzECyj6S8OkcQDq20hbdavQWE27JHZk1hnBkse
8leU7fo54MA3MoOTpcm099z/bkLZN92RijjcBs443ENeZZRVw6ep06FkRnMXsrig
SlgdDsUQ0ovjHC5wQGGglaTg8AN3RG1XDAalhKJebeozNkrdPZ0Y9OPWtUsSOJmk
9q5CEXkSBhPGkoEUtAKBMprCfSc/yLSlS1qatgQGi1UX0dZQ2isS+L3jjgpGJHGY
4yLCgKFG5RobP8+YqI/pZ4N4wsI8rWdeFlwmyyBsRDKDCvxZuSJN912LoAt4EkKZ
H4lz6dPGLjhS3wrCx192Kc0BLm3i9S962EK8ladp1czQ0DnIq74PebFH2fJucRQM
ZE+PJAp5brkEbz0DoFMRQcVYzFWob8XmUJXuakuNbAvctb6lWKyZUIqDvcikK621
zEndKZdh+fk2iAFPzqoGBNGE7u730f6vWrHuOCVZljXNWzkR4IQrRqmepCWBySIL
PsbQRvbPt01S7DjWp9cmJeVHRAKSsYlGpzJI2xeWrQ+ChnF/x8XKlPxfWyUjZ4M9
+wkKJmFPMBVptAwvFt7qr/ME37Rbs5JqAfI+Jg2C9z6UZdFYJ5jg4XqXSDj89mh+
mJNk6DNLvoV13PAfaMgvUMO0YuHAs6zHdqI271T8EJN8Yxr8fbOVtBGslJtL7KA4
0Kxc/WSqJNiWiaNRTmZZwZFNXFTyEBxopJ3JE7BTghsaL/dwVhvrXM0UJGM31i6x
ATnARw6ZxIuslYwrOtsBHHTR+2rvwNpn51zBrBLE+cL/AKVTCaBHC3SR0fuvnZUc
DZGScZSbaY1ludfyLf2wyBZlHWN8IZjIuaeUzcQ3dvgkly5lx4mPrZ3Q4DDrNS8s
182afoXdab5uc5Q0ecq1Fma1Gc/IvfC/QUPQzPMsJ/67KMXLfxB6eEG5HHDGs88J
lINGr4wcWy5R0MQ9xBzjLxTjazYHr1gM+5wipk74wOSjQ0xNnnuXVluMGaIdbrEH
ItufyZlcKKOgyzwH1goG4HqHLghimCV8wZS8HruAJsEc0dIqLm6R0jyCDccXiefn
32hhLJAkUdTGVd0H+U8JWqAQK3552x1NfeF+iAvdBLUg7YTo6CTEGBnhtSiMoZJW
CtbyFW4Du7+w439txxL6AaIeDD19mQ9MjXEh54B1AHW+QGnQVoZpPGCfDQBKJfZz
lntQCHmvYvgEZPCogskwZLlb6DCmyxGFETM06ppKDak8CEEVyC5HNFRettwXYTVu
7JYEolgx7hGwUGeiaTRQwdUxqkueDTt1ZKAGWqGC4I0m3PXhHth86hld4jOtOq3Y
x2gu0dlkxvhkp1NN6fJ0WUcWYRntLFDCc4PazujCXWV/iGp504WP7kdDaWr+YIeL
+Ks8W9CXWtIhrrv5VQ4B/MUKm5J/S/YFvhDzjxsh1xJz68PMqN1AKSt/odcwdllu
UM9DleEabyz6KOneDfIDhEglUSJPFftxvKKKtMsUzwSzzx7Wf1sibSPGCZwRZI6y
X08GSbYiAzsfxslaPgrJP35MTsITaHispRPRZXUIsg/H+AFe9/cqxa5YExxrNj/2
E2wbwUgonvYz+SA2hpW9GjbwKll+kujmJO6J4RvkPgXZVrbGVYvfHSjFDcZdHrZT
4CzIocpQYiSXQOinjJCWk/u4+w5MCnutx7qknVDMYpdwFdmD8euSCyQv8Qm+hd4E
pFI4pFI0WulQC3GaQUjmksTbOnFORDCNui5mpUymX1HGh34wSOGDGfsyXnj+wU2b
FPy5s7g/k7D2o2Z4WGnJPPY4x9TQGPXAI+12NRXBopUJf6gsGJV07vDUFoXetJcN
yaubrXemPZkWU+PAfKVr8Iy9GtlXucjc6yt09JiwYrGWV+9/sL/32A8LqNt8pqqP
jx2aN96gKFq4MyfyanhteiYTa0cl/xs9o3XBQ7zVRrDwmoOJs9l5hgzMnWGyTvBM
qr1UUtMjLOPtY+jWYMM4Zr+4Ly+ORwyUwBE0QH9TyIbqSzy4MNBBAQBzOHNVk44P
L2J9M/b5ZHPEN/fXhab2b/C7MZ077ogs/StuFs4RX75xM5HFyp9FU+Epg+jgLMj2
FXPRcp1a8Y683earYJ4qXC+hVPFVmXjezBphMh+vHLb197/vgv+2zYaYQCIX7iR6
K+B0s/3Oid95d7HsWQHJbrxll7ls5oN0pGekpb9D14H0WxXqPekydXzqwLez+dYT
X59dbhktjkjRb0Q+l4zKcB0uq0OqzzgVF4p67mASX6o4MzTrip/w7zQ1Rcx1eFVa
zehNZuFTbef7q6dOyUbpF/nyql30lzupl3M96j9McTV3jIFCG6VRFnkTwAB2c2kz
lXpERq9GIbCgvbWBU9vGmI67xfkxwUlzNjPQZm/PAh0ppiusEZB/P6k08RbVlBjG
b52cgyn4SusVe7R5OSa0IaTbm42yqJnqT+0x9qZQrFR0GnV0xDQWJD9+cMHtMJhZ
5NXL2Ebo0HUSc/qrnx17kl2B7iA7L28CjXMR8H5ExGz21o1iNo/KtI/sCxotVKXR
Urd3PjV717GYHx82aHOhr6QnVxwNwobIXMjaJHSl07NnExwnJ/sqxGTOzih0D20C
X1A8NZV0SQyxdJY333LLYmwVDYQqLV/xUfJ8Z+o8cKJk6w2BSv8OCidEvs8OeJ7M
oZ61wlvYf6X0L9tyvrVNlBxoUwokeJd9WZGQQ7q9oeWsoJU96Ul7Vt+OETVMA2q7
WOiA8FNZOxUaCdQCJEY7vlsa9iiB/o0M2+Y9syrBon8f9MeU+fWZE1GpuNu09xRc
WLlbFlDRPRA0rdwuquseK34kLL3LR24xe0Jko+10ASbuZrGpPr4YXa/L/L/CYmBl
hTf99izUHiaeKjtQASfHF10mWm7a3jNV+q7+yhB8i09yOvHDPq+YWxsTv+b+zsKK
xYVroUUVsFtRMXwAKNZ7/Psbtxn8fczGJXjOI8IkwZ1LyZMqq/MSlMtXGrl383xo
U2Y4RTaYwyJ6GtUsgHseVa+KA16+LN947LQw1U9b5IdOXlhvh3IKMbeddtZF8oI8
g0R/edAAovElY/fIvbvTcTFbixIR4zrcnLEbS0SD6xll+bxmNngdWnG7KXUfpeob
NzRuQJDZfgpqKEUKX495BfpEBmOx9cyL3xfcnyj+UM4uAlez+vbC+yl6jhzAQEt8
vvGTOtmTXZJ0z9LmeaQvrPIUmYKM1bm4/2qU3wKPT9Zw87JFE06UVRl+J8aoFY1K
/JmORdkPl1w3LFb3beHQiFXLQXaz/GokpwD1m769CwBptsUzcp+jlmUx2tVOueWS
uHPiaQgdtXMOUpc7H2XsvepZzmWbuy3hEAgJphrbARPqGjzvzNkSqny+DBJIsFjL
mVpma42EkO6MzEon9Cxkz25LKxFTZucqDBG96ZmdTyElpiBioeleXMQYLmAa6nCs
uxOzPt7JxHJmpzgjRIhuwt4j0OKZimc/F1qv0136rr/uI4SumbWD+M2RKmL7YgHJ
iHABtexAJaW1vrpkL32U0haSDBuV5Icv8Ym/3/cjKCY16PWQncVNM+q1aD8LSQ+e
9BEL5nYIsFFAG/uFGGLpLRyko/w6purfz8wdJxQ3hP41rpmdBiKV6etDgbwfXfO4
TFayV967rUQEfWCXTOP68LGzhzaslk4ow3VPdaIzEMu+PVV7IAneZ/iV5SJvS1PF
Pq0Cx4WMw5PAkKCZyJtOXQe2sAulxQaYM8+SLVvLaI3y0I2FhkF2qJ9HMi0HY8Fv
/14H2HYA4aXOFJssOEK/nRHM8AkbZ6A//eF1BNO6VOqO/BmYE9CCFM/byAd/FH7W
/gaz9fF6a8iQnt9upb3bUWxIQTZW2Bdgi6eQ/ET7WTmi5JC1mDxvy58XDf8D54My
is6BYzIkAxfR4EpBh/n3FcE2Ie7Ko47ngdYqjxbri7O92EhGxrFYDZHZQgFAqayf
GL0hjFwC70351+gnk0M/6ivnYBJYY8OVY6KSCgOumcpaAGhqBWpt4p9dlDHN+xXb
pAyqxOHF9jkg9pVfDa482Y5q+CfrsA3Bcc4ZOjYvaSOy3hiZGltjI/SYt/Y0sBH2
T7NLTFp1m4MuR12PRekd4tq8RR7hD3UzqnSg0qYxC/4dfvqXyE02XfWGAGqWFoxM
EBCxLaKyiHTbfEB4TYBaLnXZhSxjysW4zu0OS3cdN5/UcNvCtgevqlunaeuqZU4J
cr6nP5Nf+z+6/kuhSn/mxujsS9teKxzxSCT621RzsJdSLcc8Ch+QsfAGZxnLWmAh
xSykKOSRwIZ5tZvYViuJRBrP+kaVx6aitwmdXl8uPIb6Qp63PrG0vajaYMjNHECI
CoH0fzbA6Dy7HrPmCVflGCs1LXBSIxGxYQaebmQ1x7LF1dkJxBjpXqgdphp/oThC
6EGKRjfZtvSL7yeXPuu3wFnHsXEev8PQ6XpdmmHt9H6BiBgyFpsYroGJ9QdE0ERT
yVV2ul+iHUg/jQWzjxsX+hy/tYTCIME++0f1Va4WegW8k1w9CSKR+3/N1cC7xZLD
7zn0rauPUWa+DELFVTR+SFnv+MipReK54RjYWoLWmrA+F57yV4VffbxD7Yct5x07
JwfE4p4bN5aQa/U/Kz/sRM+8yhahmPkqeNhKSryrUAMyMLQy6eq9GHG4IjmWibcI
rkCNTuJ6IznF4txyrTLCY+Y3wKV2N8rKYrwqJzMs/WpDu6q28HgQMlLA+pT5wnD1
/KQuz6sR6rYH9ziNHp9yxa0BEaDqQAG3WNaw0rJni0+5oMquBJM37T7Q+UOjMe07
9BFI3VWg9sgQlnEZT86E8WP3wIwyCH96bVv1xPFHO3zfV45xw7jq0CrThdCI/yhZ
hTbYxUswi19zF2dncsgmaBLxDVOyB/7TgPeGr2Xze4RVs/liUulLHhOmYpdj5sYS
9He6OSYL8ghQzguJixIdMmUeykvt0gfUBU2Qv3nb5cs1kphLFvgEPi7CD4NruYOg
9QSke3YwVdsrXkxrCJVbi7UvmlHMYiPdmB9l8ZsCd+gT05oqgJnW9dpDGAHA+uR+
aZMR48smznPuCHJgofAG3R3MRMTjnfYV+Fn2jwPyxJPKl8OY5NAiLnn+1IFXlBaw
hnhju+s3GyW7e9Q1lQjQDJO4jcyHDdSSligl6M2rcvl++W7Ne4U6K0roFn9ds6X7
wubOQkZnf4SpXazERkAJDm4+DOZ74DuH3dJ3vJmhgjH3M3jq+qop5lYzCMfi2usb
HXjPxTBsFffmPbPznpfz8c2I6AhjznExTAtAvqFsn1Ntq76YjCWlXGNm/6jnDeVm
gi0XCeoszIDikChX+NxLSBSN0o+rJhZNB39800OC9BCTIVRkDJQnMUFVPClco32F
ZFk2uhcYM/Bgx7ICol52UDqrVUqb25J3B6uzXtjt/TVeyQWAhxs5w17zlI44+UxE
bIzyD+NTmjtsFXsJrZLrDyPLUara+9NKvVyRktaTwE7ISqcNhu1II7LcTf7eysw/
jxgAvGJTaaGKp0tjhXd2uV4h4CUlFmPo/YiK8lmKmNX/l295TsCbs1ihshg3JXDg
wPzeWVjBYl0uQy51mgom9lCmioVJGDkOYXP+6UCgeYbsVVT1A9i0oKCNjDwji9t3
8SreppUqQvmxjOR4NEBhDLVk6GGx7AFXKHY1tP9WgVkS4NPlZSuSkoHkMDi3xgBZ
mLTxPbiDo1X0wXPmlcF3nFVJDMCcOIIWXPdlG3F5WRnIhH1M8bdd4TSTICvs7kWt
+9FzAPJ5fKoKNCuF99s3ZsyK+fSllGPkRaboZFmODe5tGWVLJlVxIDnfuod554tM
3txkIVezBhXgkCYcf1p80MJFtbdEVUiB/GLq45eufrW//r8dvf756hkGmEBVnCEJ
oEf1MjiMx/gC9dtbhVEWDgUY1E1cBFBZPMazAMfxfx41aGKDzoRWL3fJo0VynqW9
H3rj9nlXfWc6mcPVgtGZSXVmOV/2kHTWb913YBXhKfyfIcSpUHiD+biU+T8qkF/Z
ss0effNxlzdt+6QwQifyXNjMJJkMm52DcdXlbaW8+0YEIa3dZPcgzn1l5Sn/qbq8
gZAtirqjqi2BnaKB34MKgAv2QRRLrpRDWxEzm1vqt+xWUM5DnNQ+JQGyOTUktjAb
OQuIr6SoAU6bCuaCHz/+HkqV8YxNQ9RwCkm/R3iIhPUKhhN4pT+d+ijUFaP6Qyom
uPy0uV1XpnVcsYtPEtMO6gsxHiXEB7IcaiRkX9WoS+d5FbEVbkRrHqyU9WTFs2BI
xfk/WlxSquyPmzlo9aM9h+nAez6hJuv6cLjm+MZXgqnmviC10QPuWCG9GYCb777g
4k/wLVGCPL1oA/LrmmRgezdtTTw24i7/uEPjmSZRswCkir5p7e44auig9wCp3dzz
ty4BnK+N/HCNbcb5u62+ChhFjEOooiqHZmkSnB50aKPkvmtgpbyVx/0PotuVqY7t
Sl2t+vGiPDWYBlBfrV09m53lnFCGM9iNwreBTmP7YPlxEUmgLziXMlIJQPfdLN8m
5fpJkOI/frutRps+OBMayiqpMw8gtULGYap/U/JhIJLdfYMBziND5TpEqnN6SCLl
xBMtWkC0Ijb7/pBpLhl+vNj0Z3EGPBC5vfH01LSg50NhNgDIAhpJXKarAR6G6H+U
azP5ahfU8qWPG6nYTEqisJruVoXnlYeIMjsv1JIzowMOw7cSgNIY1zSbh6z/PEAV
fOucARaeFmeCJPL0xurgfwVxBgJyCMapszUtEMyUX8RcDOR1j8d6fZFyqZp8HrMi
gN3OLGTOYNGEUreoP0MX9FquPhqvp3IGiO5mgbi0Kc73eN3WtcDHqAqSvB1jWUO3
Pl0MdASkp/D4RcQgGXHWB50WMjE/wNnjTu3YSFdgB5kx3J4T9mb4lb4dGk+8f5L3
xkKhe3NogLJwmmvt+zWJlQNVFJfHO2sEg3EaKHJQttsFFyfimTgd7y0vG4YExaCR
Ue0dFIkqACG8cLyubyj2OkF1gL1siLkbZsPFn2ZiC8y8LKeE0U1WOjoSMNKwK+zM
ga+kI1d455myUE+fGclXpf3n4kUvuHfvOQHyzMae0IJoiSIvX23VYY9xrkj9IDcb
3DWGGlgkd4ZGVk5QeBLT+SvD8wS+yAG1krP2BeHcr5c6YhMsadZJxgMj1qgKw+bd
zwyAhkbytYApcD36IoiX9n3kN9K0vsyPAcmBDxbUxIw3w0ffYBU5wtZoHOxxnk5S
RoGOUYIPWFhzB3+RukAEuSL1R4O4x38aCCmkU7zvEwa0EPeT3dV1JciJE8E5Sg/M
epvBODjugk7GPt9+s3L+SjYTKa14SH3XVttz968zwKZuKvA4kb6Vn65QwPeZrKy2
1y1Lhu3tKlQDsX+r16Tqks8OZaWq8FSOQ/eus7hExJer3fnaU23I8ZuLl3WTrckI
91R6WCwZNWK2lgdgm3EeOY1wCZ74jmOgFjN/7uf4kNWsFKhS+sZ5MsSAaaaLcIXA
R+o0gp+gKOc0Xj7wZ5RgMTAs7l46bQrru+DMvIPV61QxSt/0XA1bB8PwwxNAeRVz
1hRIZ6ZIrjAYHa2ZrEEn5ptBRgpXAJKQmCL8RtTXiMYzwMDItIDD3DG16gTTi67M
xjmweXbKKAbXAhLHEvchbLTojB0ShBg1pO2anxo4XMxKvtOM6lfNitMUavNKTXdb
AzUtQxgYQYKiXXJHPAY2n7aXfvpNJaQOIHNcFAf38hcQixNHp2oVeY91+/0mGO/M
99ido2L6JSLoEzfwFT0QbdPckuvkEnTJYLgrOB589zq+9PrYnr2p5fJDFUuEdkS2
Uf4Q3WyXZPjvyB1/sBFT2ACjpQZannSTjwTaXa+QNJfXT7++MtgHgAX+bego9Zgz
W0MiDpfpP5NM/YRZcrZJal8SPYqHySkvAiRlwluxnu5nkdvANJRZDIOva+ohyqQX
OofT+EAG3F5G+jTIXRvikzn5oTLJzQpYwIMtnotsE8PRQ/NdsOHsjVqS6nKzghSv
NR8W/hIzhxIvGQkmXxEp+C71ZOXhBL9YmwsdHNPD3GzJtTgHMABOIfhvdiEFij9H
jbtN6N9rGh7do76n9oTs6ZqTQqmPkYuQE3ePzbUxRA4Sk/1sCejv1iB6E3PlfCCo
+QZIgDABFpUgxHFNoo5b3QAyXxfKNMrmebZpUPztelDIDZR03YyhMQUktIom71bx
Aul9zRTRRipOu5qRjzxnakNI3pNyv2Bgu0IpxUmke3LxPKKTn0gdwuSObxB/7uY5
5DTvMyJQq9Ubow+14EWAMOThJIBK6GqlqvxTa8Wr6mowsUSw4tMV4dBRl1VFJh63
30whBfSwB2JcO6RLksB7Te2Kx9uJTU1RfPYImpmb9nFeUCQ9yXUqMDW6cjYMAo5e
veAAXkUhLbSYwRSGAyZ22L3qN4zSTnpEERWWUs520dDHvdfMP/kmIqEPvsyWiVpj
twhw6Z+ZDObLDh4yErVESwr1+wHU5w5OtL3uQyzfAh5zy+xtmVmsw3/Y9ydJgauB
bqdSWGbTH1RkQ9L9yOWBkZlKiKVCB/IwnRqxYdxmYE7lprJob/q3o3LdCT2m+LpK
B/WOqPmii0XIDA1Jp8VKsZ45/XWN/S7/l53wG2DzfT9Klz7NSaxRQXe0DQVzR2wv
+JBYeaiqlxEmIqM3NwIv54SPYPTqYz8G9GZTxLdzLDeS0JZunhWayP/kgmHhJSQL
+R3kAfQjltpAaoE8hiSlld5mxM/H4MRjq3WP+ZFZThkalqAWYqgtTCA/RWDFi9VT
7ly7gNnmvYUIGLxNcydj5HEDoOf7rFcv/eRU/cEpwTnfx5WuA3UVIL44khuFvQ7G
YT3SX4w8XpUW7bd0szquAxWo0tmv8FoQhqwGh+Z3Y+cJyy1HE004IkPYEi5Y6+b/
XFOf3RrqdtpnQjrpCux0CN7mPm6Z63nhgwIJbIvsFFwnBk6FcpsfwzkoyN6cx55X
SXQoAgxG/kyefx8Asy8875YqwibedMfxoJxV/O62Hk5LsSowBJa7qQ/E42BuUyaM
cYfCRHd1uwi1mYi5sDS2kE/tKXnFI76AdwB32UpptSzQHO7CIei5LRFZnqfKfuOR
9HTEYWrHeGFtjJyMoypKZp0qxK1OdSSLXHAMIi1cJP5MlsRU4FvpcxpAppgc3wXH
vwSLsD6yl5rW8bj5R7mY4gwWvpmyY8kP4nacsKecVn+2y2l5InWcgTV0cINSALfp
KsQQQpxfOvlldMeqB//oojIn8Ukxv5jzLxT4Gm2C1CEcdpvRM+wf+Bcyhx1CvxEq
m6Ixhh7wXjNLPGPd6w90/Pha2ZzLmHXPnoVtlbUGpRWjkspq8yHaUeouP6CMH7Ow
h3XBBip0ziCURB2bxdswz6XAUWQ17yUdXgnieAW93n9heKiRgZpSs5Y4OgYmO2+p
PfRnAJRIyGqlpe4t6CmJuhubjjYhMSDRJjwpkO9GrBDcQ5ZxYErhN/IzhZS7Xm9b
uExRTa75/7pzXntzSArtMomhKx8fmamkWHLUv3ssWVRZvBall2OlEJkwd3GwRAvW
9uivpHcCXJH5AlpthGZomovIsaelO8lvn0rzZW4lWOciJ9hVdlw9XpQh5QJwYD1m
ehQBk7pU3AWd21COzQc2gxHcVf2CE9wF93jtrsLzUSbNEdriUeprxOW5DQDt2/kh
jTprrSNHecSVVJgMOE1mBx543scJWIuWyhO+q1TtZQDdD4i3CX57ywefokrzFpyN
kM3M0KJUDVOb/JcCn6NPzJMH5xIvX13q+nz3PxTHpUDNWLl92lyK6hNL6DtiTnzk
cLhRIlCOetHIRTLb+DsLOO+A8mmetSTWibof/j47+TXeZ5B1X/DhdUgaSKgHfV1R
xpJ0V3BhDwPkqOqaL6PXGOy0jDjOFWQPZr3iW+TxJ7SXRB86Sxoueu1QIDkm/QN1
DW/m/f9xxdsFNfMiRSqMHfYUp8BRGRo3DxRdxvU3ZySr/VZC9kRjc0gU+47HYX6C
Le3tgaBhK7Z3GVMYYcOzEd+UKrGqse32qbLy2GVBirq+YSIFnGS5yv1kiv1Wedfi
CoeTUgWYWFScVI4qfLK9+cZP3xQjTeAk//B1S3tn1uJoetIc7ie4F4Y/lVUYdmPE
3cXiEFhun5LSXuCdXrwfPuFsEOz+tI3DMUMPBSDeYdOZyeXn5tVxaANMeWK1eK1E
4I/6bf9EZjllv4/rxBI4iBUDlgRP4eHoqcZFtLfy+F2cLlXH6dJ/jIV4pkE/nkOW
V23mG079nQmcM9iJngNKOu8SxYK6ZZtZpd+Kd4zaf1UklifAkmkBKgVVh/O9qsjA
M1E5c5xZTJ7Gn3JtWZAKvQK2KpojZi1XlIRnGUBivMCtTtyF2eUr9arXhFQnWoKL
Gacd+oVGXdZH5uygnVbpqcyy5hZSnITfsxuvMZELYlV5neg5oWhYAyVwheXhVOLY
P0+Fp8Ry2omIUH6Y4mJIdj8XnwJxU1+mEsjeJA8q7vVMxDH+lzA+w1A92fsARjUH
6r0zVe9qaVVMTAhviLpMfyU6IJ1ZZUVvXeDHB+CN8ABMP0cgI4HToRaJw2MH1x9t
MRkilNSdqxuK5FWSCYlWBvxcC6MT01VZTaQm72NhhYGK6yfNtrO3SczDaI1Fpp39
U6/nAMKqildcV1Y/lsxZVwD3ZJbRoMtIhMMxDmoyphkNUWUduBrPzbzv8+mOn+mA
uBdoGhGtLz2z3yxDd79Fk1tmvyAjgfMFDWEENM35p7b/SkfOchW+T4TpSCmrLj5W
NSMk67VDNoVthx2epK+kP3+SBfhJYEEjjomwkrLyr8+Go6AUHm7z4h3nA79bmFp7
NMsZdaUAXL13tn2poDvimilZX9sU/Uxpv2wpflwqaF2gOzOxfPWx8+TL+3tYCwIa
qUVL0eoyl96CjzwpHliYwiO9fYr/VcPPo3C5dX+4cxESV53JY1pQb5pU7LIZRTQW
VgsifcPinbzQ9Z32qDNGU7A9I59D3YclpmsE4A3pusRT22DVJZA6oZiDaJMFFcqV
v9bjGtUGAiMXUDPomLOhLUrg4hzRgRtLSQyTp/GOTVNzCvek1kU1PKEW9dtOiCQk
04kGlQZAVsVAaP1og+v7tOtz8CQJdLTFVojivvra4BUbxWGTWW4O09DXlYmuX/bg
PjRWVa/yYmyEP1OXfUM/Iri/hkGSfJFOZWzGsVCvMcBWp80jY9EYp5th2eX77L00
ATmgpJI3mHxwTDS9aNO8hKazMpRFQZmjAWNeYxbzTNaLXCTuajO6Qlekcd6+R/7A
c/DwyTwkMfeTo1fsfsE4zja1Dwx2XytVDrX1kQiPo370TqgEM15h5A4kRriJDGGL
/0FJEE0s2lI4zyLhpxIfdKG6BUddfgsXQ17SY2p4hU5gzFIKVRjzehujjToWqGmA
q2P6lMz7Tc4MlJFgkbF39xc0Dv5ooESHMs8FoqguOboFs0X06ZVS1NF50EJMHbPK
EUQ1ex7nMisbdez3NPTUJB+KQGppHJxozST07cFvEkVurX5v+htY5N9mUHSBzAs9
khGwi6U39ozBogKTIXkk9voNjhgghGwCG40UD5v5CynYbSnPILb8Vgg9WxckZKwI
tPcppnWVHM0Xdvkml4+qL5h2MeP98tVKTZ8ZHN1Djjd27kOgZiCdWMXwYan3OWEc
VkYA6RuhIx/dXfTfYH+VFqcnoL/LK7Xnvt2WkQgVMD01UdFdXnVA/VGc3UmN/IVB
yyVd6c8A+K5+qhQwUrLIsdIbh0FHvKyHsNiOsIRoD8YyNUWeLwl45fdQCu5iTa85
fS+1fcT31DPaoFuvqmv7fZPjVSmsJki0ddwV8wslX3LMfsEPyGS1dHyTRIImoxjF
T/H8K6CdhlKUMf0Q2n4U7yLjDjRk5OuZLEC818BvUhdb8YmFTotiglzqHjO/ZHXo
xfs3iIshP0lYIKQdmSUs4oNl6y6y6GYJ5JI+mJwXMh2hY75zCrhM6nxVibBCyyaM
c3MI3Mc9B1UKmoFEGXhusdD7CKxagkDNRYODcLwzciu2qSsmgs7VfUpVXKlsFh0M
vFzdhCgPtosIfP20rqpgitSaAqwlcFBrMG79ONK2hpUKDZ+YW6li+6Dw493198vy
sqXJWtT/uYY6QHEwSkf7AxI77BSErU2de3xk1fhMivfRRJ9j57A5knYfQded2dpF
9lCLZehq2aCitnIByoKSlN+OzPo1D3jSynIZflSAKGFTlm39Srq/i43AfGlyPbKg
q33Qh5/WgaEqFjjJgKk7NABTzJfNX3V7hrmR9fjECebOjVZf8s3KSzZM6ewgeQtP
gPBBxAzX1Ws5Yh7MfU1AcYf1gJdAP9n5H95RwN7eY7Wvt+8q8+DuDjR+ZTN/Y6nM
ieueJcas+uYgur4neFmv3oJXSg+cpwHqhE50Jn7qFX+1LMl0mNH97uIkHwzJI8fm
gOygrDjvN8qEyqE51OpODRzyxeXeqCLKjhc/YPOA6N7WD7flQu5NTYy35F4VH3BD
hmRCJtKntGwn5coJyHCwSMiyxo/xJcikq0C75fJMykOAX2rvCz5zx6beORLY59WM
VspE/XaTJe8EluvEcMe2aMCXQzeLVg4s8kk6Sdp5vg07pq90WBhRI7hISt1d7B8C
KKUuKTnoEwI6L+AZkKMtWXTmqi0evbyh3hsuynNLxC19lX9q4QoyaqL/joLjmbnS
6qsprOQrQ6AaBZohFlb8GOWAZVmGs50lh70PdxeSWpwYwuCoErKeiv2fh+GUqXa8
z9NlMx93qQ0fHkVa4OjCztNobaq2Pg5zONHYumV2JWUG6lYeCGCn84HVa8s3e6zt
jmaervImoll/ikqVSLVvV9B7N4Ej/9nVAUV03RDoUTJQH1Dl1w8WtzZmnxKlqvUP
297HAz4K13+/07grmPqmAq/WbQVaV/Sm1m6MKy7I/Fpky2H7MNjeDzPiAt/0EHSr
sfMf5LvHe3xLL56NClNEBD8gx/pOKol9385HHNXpbmAIrolVDB29OwY2GpNCvHcS
GvuAdk7i2Kl5kgXSGro3X3Rs3gPbggdxQj30dNjdsLva3kIkchlfxnkMSv3ABHYC
NlucVIS0lylD+T/WoB5JEcJjZw3aEUk8vUyjQW5hbFioiZvM3Vgl2dBT06LUh8ra
mVlMyYj5WDeqm+0e63ULtubnENc76V6j6iBRGoI/2fhaZytCMKO1cN9tWaaQ6vph
7/i45qCLttrDT0t0Ta+9eYgQ69akv0WCj84+ELm+1iCxd1TfcLfh8PZN+L9WqOtz
EHnLPx950KdLV3Om6xyM1rJD+fOFfDhl7/bjOq+cx7v1hVK30gm0qEOIRlUWnwTb
QwTGYfp716F3LdLNNeX0Dh/6K7Pv/6xKccbeJd25/eR27AKiVFzAEJF6q0Rru9EC
CDr9VjGyh+ZDsAVaHXLuB/OKYWnDUHU/nWrGEzXnR3bnfMpmcIdJW3Y+O/jqfYRr
e59tD8WP6kYvIqHoUtCCRiW9e0X1t8UuwJXHTS2xKAsPkIw5KIIrnN7W30pKy1s9
pcO/KCKV2Tpc1FK6D4jb0VYmeL8WPg/18w1NhELeV35+3cO39zRk1nMFon7KomV1
HXLlqM5RuQvzekKo+S0cdstiVjBEgHIrHGnRGB4ObA2TawZTIKU63O9nYCmoJWaP
qkRp8zzWDDy1Y7JFiUPkEAFNkesRxHmfIjZ7WL8s4nBJMVsST/H82L22poRtjjcX
7TGvNUW30uTZ+x1swpiucIYp2M3yqu3Ncw2Y+LrnjxczQOCC4h1FxabjWHzlrVD3
hu8syzgz90Jtanla7QRruDZUR8IZVPGqGKTqzn/QXDedPtd6tIGYTKTLYU3/6ZZC
GY3saYuOziMTZ7nVfPQfniqUe42quHyk4gXy65v2SMaj6X2/P5cPydeuMz3khF1p
8O2v7GCFdMAJI6DkSVdn903Z0h1X5kl+3LJT3pH5r90HVDJjzpsXnQvt5K7W2H1u
DEqePkN4tepGGN62Adv4SMo8RmTH++lxzOJpxv7QqfgqZqIRPyT3YqAUgrX39LrH
d2axn7Aybdp8afcGeQdWTfwXzAphqtqBlrZwEtnw2wHXu3SZRJbD5SbqsuVTa//z
gh03Bgwaepue62LXoCgPyif4qqw8mTAsgtzrBmYArzBWWIPUSAO1U87+Es+JfxyB
wLnqHdXKI38VZBHrbk6WZeYQ3mjRVmZAQygd2YvWFsypfJPvIUkyKScYWaount+m
c7KF7GZuXmYIDKbsTf6DStl+cniK1frTnVqDBJEQVzk/t36YyYT+UigAW9864jwK
aD31v/wtYpd+c6CBSJI3p4uka5yUD5xmDVtTvvvWt0HVpYq3rMqVyrsEwcDdP3Tt
wCi9HR3l4cGxsbCnsDRuAuaSujOIZPex59eQpLkqI6PHJXlJdp7x/aHllk31T5nx
TsKkS+mBJQYNcv85wdRPsiXdBGiiZE5FYiQX4KKIgTarno6EFLyhNMsvKQvW5OMf
FVwTw2nx/QZnU+ctdZckvJWdTwOQdT+dW7yIGA9wNttQFxqs9vTLe7kDUq83fkYP
4B0NGd9l978WYpfFsN9wM/TgO96rhcLiCefVOFK3NgA8X1NS252cjs7gNePIxaUE
PfSqCDVlQ0AeO/+V5vJUW/rNUovsDCGiszZExiXZHWbFm9GFFjuC4T8g43R5/eIj
VFNDwaidQE1SQMU/EvP2Ze1+bdCISFc5b9Mt3hyke6ZSq7ppg4fpo3CF//8EeWHh
dYxDpUrh4fnO2WgiQr79g+ig5fI5bcaI/HDKSVNdX3U+K0bE2om0OXNsn4i1W1vm
jTmUl+30pvdaJBPu3kxV+tIZiDmnGtQsOYlXd+dvQEJFkfwUbLdfzFvQbuNJsb7e
xNGBzsqx2/WQy4gA5S/9bvIU/ggpVuNrhEjJCHf8jjC7GWZ4pEv4LzYh53ci4VM4
fPYsNgNztV64LeAhgF83Sba4tKsBIMihwlrnPKZlt753lApvsCrfDjwt/GtD2IgX
+6EOtX0zi6gtnlsjpisPDK/3jMqLoQlf1GT3j6CtGqjxKl+WhetdiCot7pn8BGoK
8iXChcO717Ldi5cd/Zk+jKpWCW3BNpdSarRk8LTEIYpwYUPqhCbcIuzz+BFf6RA8
daiSQM3Wi5IErS/syoV7MIcsMkns0axK4q182qYJqW8fKiIJzlJrsD7p+xut4OE2
sJ40npKHXiXeNCwQvGdO4UJw1Ei6uS3UJ8UMD2bZENy1tH6AbfvSFpApwXz/VSN8
4vlpNWxIayoJLk606KF5i/8z6awdBqmWeVn4J1WrU8XpXoJzLY0+peVwCvvwobPC
WUZzJSueNxA3IwPe9DNv+X/aFcHXodGMfoJHNKKlYd2Dm5VZpFzK/Dxqcv0+J0BC
2MHrBXdnjoCF7tMljYSZyxnKWVU35OPQLA/ehbNw8sKYViPczFULWts7vPK4UUNd
DH5Y62sy6CkRBMc62n3L0/tosj2CgiAVX9aZRYEBhRRCZZGHbzpnuuPh1NpCPGNQ
b2794ZveEBJFBRAEo/5U5nXWCdwv3e5wkzbeiUZWPVYZxfYj0j9GB1macwzPFTMi
YrQPn7sQxj2X1eMCdbggVPau0gM4lRoN6BeRbOoMPdIMiulqLedU2d7pcxvorLEm
XPbVozTwXBXTWdejHVE6JyvhBVzVIAnLnnVbjvDDMrNlHTqaNonKQV9ewzkfRTM/
GE78Q+DndKmbx84AdHxVaZiqAaPjO3Lb17Up9MmTvpUxRaIyAjn29hMZlGuz/Cxw
31V8bMp0dw/sAwDBPeTl/wexfX3Nm+udHSSmo6H4beNP1AHPSHdGKyDPgqzKzWdy
iWgsQXaZNABvVydvRzRs2uyAIn1Wu1YtgvFmN/QW0dKI0mU2NvAvgLx8mlY/kdKm
aQ7G1Pssiy18pVO+ql25rmvWbeog94O5A/VFiyWqYrWB0Lz+BWzFRARII3hry2MP
vSnZB3t4zugBp5wVbevlLwFChIsAzRSt8iWB2uaxDu8L933QMEJxn5WUq/t80IGy
EGm0TLKG77qLoaKQgCsfosWgOcKcAbC/T7dH22Yp8/Rm26JazSWjOJYHJimAIq5B
ZVDdm/tGWA5nSJ3pEypQSvrHH+KBJXRiy+LPBDz3378eTdwUkm6zj+srOROYjQF1
Od83dz+W8Jl/F6QAWGPv/ySGRYnA9tHt8FmUQj2P49FL3NZilRZGbRwpHvfiQIoL
KonE0bKdvZQRloLAeckE0ZYMFfvK8LlsmtNqpJGpQ2hBS7dGTBH/kJmgrAHQHgg7
tEiPfP//ZNoyfExXtls2jygMyhgu7mxYJ6ncu+1U04DMCJYPRhiZ0n5MicbJdAsI
ulEw06NC9hs17YEGj4aXXqN429KK7x/Zbq7GurDcUE4cz5GnWi1DF3mk+5iezNPr
46qJ+HXJdNzpwae1izK3qtxk+AYDegVfOITKzKqrvbi9w/L0+4pmp36v4hcKLmi4
L6BuvChwfQq9vMvevsp2ZI3h0nef2ok8hTzv2gNNwfw2RXk9JgaTceJSS/6S8/2x
sODVrSYKBLfVcrd/QLTj15Rd1X0cpjN0ZeFE9cdH6cLOemW9IJqh9EDjOeIjAnQm
h2loF2elL/ITGDqGehwwOHd1YZPJspkf7gJJvKle6xmc8m1VjWXFAY4oB/0O/xbx
xrxEbCThvresRAtRLvEHEnmkOaVPtnMxmeOwPZGffL2dSXTXMcVtXO9crtpcbfv7
dUynXHgpI656GIiBMEKV5N6qdZg3AriUhiH8ESZFtqp0QESwglNcs61bPdfMrkbk
C4rLmCjtVSl590zauPlW8Ws5Ebd4HNyqujCJUrzxeQ3ngZ3mS3lwNyX/RgAIm6fM
bZs0hbmB9wHLGT3f/nc6lpQFT6Lb8oq8/WTpTliClMC7sGVtzIxwBdwej7TPYh9B
CyC+jvnfRfEeWtJ5wH+mmVgYXwuz7BH4WFIpCLAzJNNxML0DhsWyxuvYFMtsla41
9QFjcvFU5NkB/MzetLPZFuZxlHCWQFSHlotbJmmGWqE0dfii99MbQgtO69m3TIk/
y4a1USu5CMmWvfC5zJTJRavdRfQ1O1ZTTL8tnIogdGjvHHvOFlSSRAYo0B+q4CWr
tu2pdG62wJNm/CVdZH4Gk5pTW4dtZshlGNouopiYm1g26NKy4q/XDMc1zDhMtfwA
y5cuG5wnUN+vVcwJ07c1XkVRLS8/avD7AUaSohfp7Eh+ZwfTycRv4/sgC2iHWFHi
vhalYzqKObtC+Hg0tpYT8Jbghg5b6cjTp8AOUfqPhkaFXjgk58/AlHnHxtPIlt1L
j84wjZWekYOsCMxXMjtmjoJwceOibFpzsqW5pMfDEbiZpOTzBTKPbr7sXAjLZYj+
O4FDuEZ4dHAVFpbAMfw0kEwcMdIxnBxCOQw+LHQP1px9SPzjJbg7JmLhIDbMCAhL
2TWkZMpCAW+88mfc17gzN8nJhRhdH0oc5y9+dRR+SLP9mnXn55G6Ykfzq8gKwSFa
HBNPLHd8PMfl6Zxk7ozqXN9cfI5/fcCUvhwgvuD2K+gnVDTXTOqtLc7KPnmAyPLS
g/Rxc33Qu70JTj7O5kKfDK2coAUg0BxvA4CqKeg/42XsF48mrayr9T+2z36/DIct
ZHArKg20Tky3rKHChw3Lo66DxhJ3faVa17ftnb6pUBJFyedimJRJtbX3IOoZ58KJ
EWqH0LGAHjDURNkd2DytXRL4bqS3pJVqkAkr8RjPJKO3+jZ3Z+Jr5z9DbCkhtM7x
Fe0AbD0/RkIpyt+/2UNiif7FuprmCiknH4Yhh5WJd03OXI9hzF0kmNQGSXEGsguz
n8BLWeiNuBoST5n2k6EnLMfGTg576t4RAE1/IpDgvWK0TNFzsjcdmhn6WAYUpquz
ARtzRsoV13pcFl+run0YFGARnZ20xCrvJLSvC5hDaF1oFCOXW5GoEsGxW8QJBgJO
3Q36Y6jygXyrzu3yvwD2CsvqPSo+p3acSmzli2g7iQ2Z5v7VmH+GswKOUi/i5nZ6
rcjD+S/k8nbuxqd5MuO6wcdrVShbNBjDSlSNXxu4DuB5zB58sjINTIIc6pvxS3tm
u4ljzU4icJTm6ckLXVLOXDsOOdTHzTNXqp8AP4xmAYcI0Ji7LoeCUjEfrF7nxkoc
pIHBaneFgJwXHkLZSOYsgh03ED/5gORPohUmoM74fgWrW6U7gFHotxSFMNqN1idZ
uIzESb/N5u8kU3IgHtPDXMnTCIdIG6I1PVraW+fII72kuB4FfRLWzj3msnseCFvG
MSp8B6KdPJ3C3NBssMo+lFIYRVzmyGCRCGgZ2pU0WoXYE7INKQfXm5vYw2vBHRFi
vcmLtjnFYHpEm0OXKOuLjPSFraOUexI4e1HI4Zx452ao8+lDElYqKEMAH3ysceAS
Ict9xW21fAmb+HAWmKEYJRiFgYvQCbFqNTMf2itl26y45IjUCsw7Tvn9HyDUVM+q
j7Zv3zM7C8H9meOdLQnqyiCY8Xi5ce4zNvG4jR3zHXrDI1m3mBdx7mmhFj1Pi5oD
7u4hDwBfR5CNbMXV+652nKQBSLu2Ky/uuLYudZkOai79ERq4T/BQgga+cCIeYz7s
ODYFpMW2oh+lrXWw+FVkGW9Y1m8zHQ8p5yWOPvqYBHu3MrQRDtmkTVxN80ttWoBP
i2g4w+bbZIh3zy3z9NGhY0OtCPFg2YN3ERyPLzimJXbLlu+i3mqILMdlbNhR7AFI
o8kIgCmYaanv691aigyETbqPcfHSvIRT9lqeQzvlNLZkmy96FoTY/EZft+ddPSiJ
/R4OS4oYm3udumiRU4OqgyyQwPSyxdyP5Tz3ebGlAGBLs1GDUineND+AoV353oWG
Mv07SBnx2n0/0pMn0+I410dMDH3YGtqe6we0yOl3LgFPdzQK+oKfduv+CWrLmKT7
Y4FkWpGrbZMdIFnk36cKPPilXPjAOlms21v9uuKVDSvFVOIcNfGRqPE9qaxMjWj7
TdGXZiO3U9LLdWQ5tVes7clqlm5RCmklOvjY3Nyj7DspZdGq1SPe2W3qVbXEANJQ
q8j7o4ea+qAmgK8C23BNLMK82gHvDNUjzexKi2Zzm1YFuWs6mlLgWu1AMPkclnEO
/9OH64D4r4nqSE0e8oC1+Ho94w/7YFqxudp0CEYF9Z/ulyEe99R+WI3qlAVGAUyt
5bRXNKiOJvpv0hz+LWP8vsjxVsHVltnIEPxzaQtaEsZdMKm1n/Pm17eR4zwa6KXE
HmpxtxsklPE0u392qZaTcerUfTtVfcSLDjgzPUyBaQgwlDCBAMo7YzzhZMcbkXbS
eoFq7wwUTcpXXq4fUJggx8MrRH/qhbKeDyGgtvNrUM0RCTyM+KsQgIj8YgeG7dfS
TFMSASoSbI+kR3nUBGJshTMFRzXY89QPs9TnYJnPb4rRJUdT1peFDYFLHqHLcC+i
bcQfhi8wygSK7pI5wL7ofK+NJr3XHDHymcKdir/JbC82Ss9Plj2XUbLLt9O/3hne
WZz5coPVF189sUIuEZDnyJdtP3yeCY8Ab23XXFo4O97WUmNzRgAEIuaI5hDFZztx
nK8byHVzoySmIn/SMKxzUchKUilMb+CkvXWQX4HLNxs62JJVjACeSFByk8WdLDIi
Mx/elU4J1nJQMOaRX5ua/ZzkHe8o6smL3xs8ALQaJqoRgEvMtoysyDc3PCfF36SZ
gWBXmGKtIgVoHAvqrKr7GGtYLFks3FPw6N3VBormdS37PCisxLtSJcAnYp1gO35U
rkvlbQqPnslfoRpgi5GFgnSF1Ky+UpJVkiNGshKleCd5fmEWlSPhajfCcFcPBtcr
ZlL7ofr5/RnP3dWlnaNrjI3s/1kNhWFZppWy4CU94JgD55Bzd68u/p2PyXHBAFAc
O8VlwDd0SNna4VjfudJr/55mZJYvuNv2/4jpuVA1frJyYupi+yzEfZz9XWHGRUA0
aqnpIzEkpcqNA2DOO2Fyo8mhXQdjBzCmdP2XKoImdq6iYQjNnufR+O/vtc68VdUY
tHhKszX/qslSUPT31CDbzxdrUzDgefcTDByecrMvRExRtfAljrrwTyuuVSBnsX1r
pj1AS65uQcWse9CZKYN52NfeD926LnnW+sXH8sjf2apvd26rKKH35yp/ZTQyhmOR
CO4y8sKgMuZ8bvzHbzyDtqAO2XXS80iOMbTxfvlYEZLD4OEQ6mI0X/PgnXZNKBRk
RXwQfmObUpjE7f0AoobiaoGEx0sZS6DTbiGhBanT8vkYQ/5zWc9tFOXtLnpzjint
k4aJzFqz0W9f+L7lpiWbnfHicv066BZr7IP9xQBRtq5RqV+JZMljFKEQlb1jVGaf
1BbVVytFNVSwfa+KgvqkCJMdObL0UHiL+SPDZnwkqHJNr+b4De0e1lR19hVImpBD
pqkpfm7twaptwzbfeusdyaYGTV51KBs/7q3VCJlOBVKjuHPxucDt03PuZE3qWt4a
Pt1vbO85Bm7IdtxUpw1paOUD6gptoNuadxCvcMtB6PT0ndrmc4ftsHIb9+90zoCo
+qe7x4XfROME+6HdWqNGQyhHe1pjoU31PBdYG3CcG12xNPH2PWoKjF+xBqhpI7Yr
d+zuwYQg46qC+lIT1hqI6QqcGWxpCWU4oc3jk8L4shaBoBuGYD7bGb21W9mwX80J
Da3qRfRcKTuumtQn2TXYs33XTj3KmmoWxLfHfNbAEQ+oOMHLb0AaI3MaNSji7e82
PTw4QGASNkf4c2AI9PmOOfkv0yXUQ+BTziFT8K3nllsPChMvijrOTdd+eUhFOeJg
Rp3KEq4FJGJteftTZktO4guiJPiDZAWIak9iOmssAq954ewCXzgc4A8lVEegcD1G
NHN6sC4yLT5qihKuNtUPYlDWeFfmDwsN/312PC/MSNnZqmhnVSl0UnWo4BfSq1DM
E11oqC4ea9Q21wrz4qLNrzwVOfJuUSSOYci4rGST8HmTVz8O8x3pI8tYfnKWU6DE
a0isoQRF8zZE3N3cYwc+o9BY7R3FWm2lltb5JpE4p0iCOjB1qtgFX1KXaUs2X9Rq
JXBPdwQaokguF8P8clN9tZUxUEd8UdS+d8o6h7Kp4/VOIkmuq6ieUPLwKA9rXOjE
VOivkwEhk3BGGckSGEutcyYCiXwnjto5NMEw/b/EVRf+kVNat/xs4q/tcb91CFnz
BvG1Lf2+ocQSX1hQLFgCDyjhe9NbZ8OAwWQfnvMwMS059LxvBEANLyEkC7Dl0sNL
6VlKE2Xlpj4dlC4z2KSxWb+8/yWc4cOfPCvKei67PoLRMxIznrfGwumFjiLp5XL4
FPNgOGLHIAhEoUgQ7sqPhcJMa/navm6VeU2uDiWv4D2QXmNScnq5DqTZ8Q1xPS4I
GKIpN4PZ8+gAdEFp8E+GZ16Q+CSueEfz/ern0jZPwCgWFGddlrSEXTWXB4o+5F+y
LGF5SufeFM3waudgH63r/xeUtrWtUBP6LxI7FLvmlExDmt+EZxmFX42llCrWfWei
RdXph70S0DL20JSR+0KaVsFp9Xn2sNJx/TAgE1sj78EiJm6OFZyufo6vMcsQJLx8
NKs1/ni+BJ3OlKBEwSVSikS6UFJ7nKYxcJRMT1aAGolguiDsWYwO3WAYsIoeGoTZ
BC8KPhp2ZW+I1+iYga8j1Bz3psEhFTwKa22dtCUmkn8kMLp6rcfQavXx2q1otArt
xsrx5UgMq2omtibSJbR7RIrnpnKqOtOro6hBZGbZvtg33bfGSzYNtERfT2bzmg1l
HLU7SbB+LqPd0Ecnj3HIigoTNb0HEhj93l1SQFx+btMSwa4CYcYv/ytU0TmorRit
A2X70MLS/4R+tyIuYFUSLycDh5wMc72XSGub68PGO5MO8jzrOX17hsqenqtHBYoY
NyDqPmIVwNwxUdcwpuuvlGC12VWIPle6ZYOhl+8gs1JxEFqXI6DXmbeeG9yc3x2P
c1PEQDAJiWbdW/w7a80eoIcpPqnpW3K1x6QEPmOyyucwKYbMD6ClJPylxxo29hhW
f4t1QIDj56gbgOkB4Qkyd1m/gpQK/Lp3WFAk8XQ9l3qjDYJPYM8o+oXbNXbDGwJV
wXnp1AyKDv+CWi0Sn3WeyC1cyCTdSDliTO45YNtO7hpxIF+1W9WCa0N+oDKBfW8m
DMPer1TaxOg9hu3GgnlGSGSZF7TWym4ezTa40E2XMIV60tC/Zj26BEeGmVTK42jZ
VKhr5GJLM3QmA/MMz6rNO1bbieMADCz0PKD9SR/wkWSMqZRBOyETqWv1DREOkPF4
bZmuvbSbbuSlscye9RPMWz4dbpuE3vfEotlPkChO2P1/dpOK/9lWuty7s/ocA9DV
hIBUclkGGvKDAqj8uNmFzsUOeKE3bdl5Y9zeu6W0rmsoheLe1HfEURLKcXlaXAlZ
FOHUEcvPgwAYoJn0TghuwNbjXRvgH3Xzf8IF6xJFVzDcUxXCCPcfTWT3ylnM5Y1S
2F4MYVfYy9Vywwj9zbFUdfSXTHoVeP9VfDgEKml6UVTVIE/ciHsGIy6IluG8kMfA
Ycqy8jbjL0eICzutGS1HGEwdrIi5JJ/Zhe6cJmNx7P9UjWXySCrFy0tMLPG73By8
KBfpaFWrEiQUMmYBGOLAj5FfN/jRt8V6p6OfsYgeFZTDODg+qLA+a0DshmWyp46q
ub1zoVPG1x7P+cDkmXuZsTsgcOil7jkPLewdXhNgBb6eLUs4dBugMlqQovoSGr6F
Ob8kG7dKfo9P7L3A1YbYDW6LMjo+hwmg9vTws3wzhm5tvk9WOhUyV/Gytmlao4Oo
WtH2oCBSOUKADGLbJQrmRGPTKtdGAzkhvWqmhOLwJHjPF41CaVwkRXN0iycPoydc
PSXRqxcQx8Hu1VZoGd6KLKgtdpz8WE2LOXJ7ZJBqBQ/0Zmc2MZvOc3HOPFlblewK
2OC/pdxRN42Kj7glKuwBNTNPLbKcPhH5BkOLhjBFCqAVgM9m7Vq85/Si/XuH25ck
F8A/hWPptRCs8hOK00lFEjrhGRA6FGWcrZmY5vu2VFYrWKLAxxOIHtiHzJCVOkWU
NkQa8CKOKl6yu7bDX+Ln0lTfSRpxSgXCLAz6Gjv/O3t0gjStPpT4mhuzUU8zaFTO
RjHJVPQDm7bkfURMCTatYu6OCpqqeSRUUuVzHoza5QViXI2kvtCIqHc2NDvWYjv/
HOWA47Z+QfsolsgpStl3VelRopXG85RqKk8zc4EPVwJ0b0ORPyDJY66q6yZb1KAA
g9akbHOeCm9LJNGJ5MuzyStKs9ADtyRr5Tt9O6UCKIadJ8YZbP0hPDTmomXJ+1se
I9YJVXLlQNgGGgAib/zr5iQNpHtdVTzQGBSRzRDmpNvOzVaSJSfwXsL6raHFZ4PD
yl8gEMqb3e9w+VGDVSQqB3iYTBAbG9jEqaz5uDUVLUEC4ByEuhmGXbueJHXSX3MY
FgwyDY54mrHrcuhKx7DTnzuVW7oT7e8TBP8IxYX7gjqqGZxCC53HCwRZkFhcgBt1
efeYsuNtrkK1xUmIwqsIbHkPil449yBgNLOqv4dP2bmkz7nfGKPrH9fyaMo5g4dR
MjG8Hz3Azp5MWWuFadS5p8HE6tjkmZqv/8b9WBJtG4j7oKjQJksfCCXOrJ/dVKWf
orwDHZ3HkTlWr371H1kl3lof2diOcZcG/h7t3Td2748mAXZwTvHT3F7Ev0+94xRl
8wzHfNm7ax2EuTtP+M74kGgwMpNm/zMythGdjyOhpqoLoDCUTtLAvwWTn5e8yhNO
Y8kyvX/+pLo168k8zYZB/ixyLN2TVdJwIVv5EJFPAotBuuB4HrwAIO3VB3Rnx/NA
wVwizssMANx9lbMMgbGykvdyDJwir0auLz+JB6td1JhRizea9hJpnrdB+pwp78hi
v8hf2yv0PkeVVBPbEk4crVFSyrlbY0rZKEoYTC3ekegnVh5CEnj5mM/x15U6ic/S
r+T6zzX0EL2rdD4M6iQWwUFsxyZgSPdOA+xuufTb0YcnYSoMNV1BqcmgVXFqEX/Z
QhNb3SZ3T7GXxAIZtjdRc7RikBb4Cb1bC72WlX9HUVNMAmPUs/EnkWzC6Jm05Wcr
UMLMIF0GuWzXNdNuWq6tFRmoht3Vl/fDEVOcekEzlVa8Sa0YjVdIt/jXDkYcXtjj
Mb5FpHSnBf3hp1Z8oCR58EQiS6usndyKKVqB6jfbWJkCa91FTsZ52sYooNVOA8nS
D05tCrHQPQvA/rgyKlVKx/K9i2oLlNvhWIxGXg9lXbr+AffXrgRMN9Q5qmK9wjYc
SFpLt4VBWPmv0UA8fAxw7yqAQlWrUueV2PjA1mm/M459Uhp2OG6ogSWQD9jz2Q+Y
zkH+NLSSf08blKqBszJrny8lRTx/rQfiEDqHKj31A6I9L65TneKQpadLym/sKO5O
jx3Y+jLrTJwIuvEfa6pHpiyP7A6GS9xWADGT0vWGv0Ki9LNPMfinj76LLdEz7Grs
sEY+i+/G1rmnQbU6awRjPHlrdb4rGH+WfJn8LLLfwSvrrYWvhVR9+PPx1TKtyHcM
DorFaK4HnUxjpAfQ0aa0Oc93w/4W2lLdaN4aNVpitRbEjmOTIHOvxOyAKbWbbNhN
AFYoXtWBCEBMs8j4qf/vvC4JzAm8zq1EyfAaklMPfX4AZc596OidMKxOR9qeQcV3
mIG5XZkoPxWQ1Ah4spTg0bWmcbJLCdvNfV5mDqEm/yYvzUrPADh28/h+FPrOVBV8
szJ3rNCrhz3VqnI70YlSgZn1nZ6oP/RHi4ns/0HRQjTV53uP2NqHOOxAdiUgWlrc
YE+bEEY/oDUYA/iNIf54ZeykHNRP1IluHxIw9R9GkrmBZo5mwkVR9XU8SYuoQFYj
RLovl1rO+fSYhtjhODUFRJJxMetuGTn5vOu/yobEEdfncIkx/Vzs5wI4myIVK6/i
0htaahLwI/fI8rDBzVnJf73TKPIwfB9eWgCKZRDFrBdlLNo6oA2Ug7etwoMdk4sF
wPcjJtxPgsLjXGvJkMINiSS3fyyb/yxmNRlnDeOFJa8MJYTvxLL/ckvzDhe1Gu+J
/+Jr0rrBh/xfblqDe6So7eZ2Vv8HHBq+zzTIXGcm0nQs0AC6487UvkHnEWii93Hv
J/3wYcb2XSg+7PwWrYNQEG2TF+s6HaOjNJbaqVl+stqltgUSyfu2JpB2Ou6Z0vVd
dnhyNFGSKiRJX6DJAK6eRZjopoKfI1pTehUSZuP/TjupKhT350Onx3Iwhuq8EuYG
KWTcmETHqrptCzccNSbIaTe1EfBKoz64ozsOo0weG/4A5fZiezGoV8Y/BI6y4Ttd
WZ3vr5fxQPwp3Rw+q4EAi6MqsTzf+NhfZC+QX4/DkngP68mdnsWEZ31uSaoL5YZM
fYy7TRICaCd+9jlccTrrl1FssUp1C5DmBHOcZM1WYFjht4BVx88gIJ/d+44FUpqy
xXKEqqgNFdgyG9o7hO4e313BuDWe03J7mHkS7CGW0kROaMLE56O79Mr3Hcl/nbb3
dxp+4mJh++LIfnReGSU20SQl8lVnYpFiR8OOvlV1hYUDc7L02RC9krlsS0S5T5R2
me121RJS19Bc3Ne+Por4OO+wdn7Pd0xlvgCe2vR2EMYVuQhL5CEyL8vvP8GT04R6
MICICDouTvDrCmPOusrAkFNKbjdDkB2xE8zeGzKiqyB2XjHNkSlhQ00BkIoryt53
gMd2iVm30XzCZZGf7KDMkrWMBEoULGHqjA2fBOXareOY8mRQUuJxxSJw3K5fFnFU
WNN7P1zdo4pC33U18fNrCC0dZzNZ/Cz20xevWYlJf1PHgdUPtk5PkEw/G26I4jfa
EdMlwmO0/PZu95CFqRZ6FEGdK1dhZow0cWQz4bz3g61BtMU9PFSF4gmLrC+koNYt
DFripvCAW5SsafE1kp20EzAjDNV3GpCa4V1PJb4i/XU9wX+Xg9dqC4v0L+1xIheY
Lz5Js3y6L4ch9NBbjZv7LwjIQW8WLoGIvepeMCKJlEsIX1uje/kzd3ajS0AC0Vvy
DqMtumwhZzjMkBvm9wMic0FUc8d6lqDhd1KvdntBs639U3rpHLMC9N2ZPqpy6XKz
A0qSfp3oXfcgIuswprlrmFZMfUgZeSHbqc0GZqlT8nScfc+9QL+D/XFPBArvwWvr
NGA8nntUxVC2Tn5PifBtm4GKMkx/Iltu0P77AoQtlLdjFGGHX7fkzsdc3lHOOElV
+BzzAAZN5IU8DJC7mUk4ex/vuqO+7xxNLl50Rlo6Qm6HexuM4MqRRB9cgfoxQ5CH
L+1r/sln5EOhqY2pz5Cayrd1yUUYISVMe/Xs4/zYBGea2Cz8tgEgf5boFP2UN3yr
EUTpNZkhQPu1D2O1W777K9oHunhj2zZP7L1ufY5wPMGM2XA9m2nmzKrrxGpnFkK3
W/dPeRG0/Zblk0ePHjwJRVV7TwKkYyo4djY5ULuEnqXeaiiDQPacF9cLh+oIUELO
MOheIshDMZXp9zXpm/3rL+zUo8thBHBi2/1ZpyUZtunyGCnWwPKaiU9j/VtuUcYd
0zvh2rlz+U1XJkLMfE5loHgd/V0O0+EvTICmBqH55+M46D1eAMv5yizFYmnZ+4AR
6tMjGTu8KRS6JzYxid/F6lNqIqHE3po+psDX5jTdvuVcYrC+zg9kKgD7c7ZZklO5
0K8Gttcfe97z15HiF2ieg8kit27cPPGguRupPWelPD1gqaAwd+tSb7MeWtmbMOoi
XNlg4caaS5BZI1gMjwTHjuTjUwTZyN49noFaITPyuEhXkZwfI/1Pjy7aA8TykjzJ
vgKdQXi1RV9b41ry/6sb4ciq0nRUzmNu26UEMZci+z25T8KfoGapHqnJgAZJlzds
kYbyKyWoSY6PYrkKcCWBry6I8QPt1SGOl8TEaJYRdy7MHcIWJezz7ft/Ga6yYEXl
N7QQwTLYcxfqvGNQb2i69xRnxul0nRe68GtgG19lbTLGQAeCKXehpBhnas1lcV5X
sadsBmP6kZSXWKr5fLRXSocaDpLv10bFncy66ZvUtcQms3ocOsW7Wt1sQ4/1BMBk
DsoUsC9STCJAmQzgathvNlZ14kTkhW7y8osPaL7SxWQ2w6MY3bsF2kNmHc2YKjtc
ZK49ImTv7rejvGG1Zbk+beuLjaByF++Y+BrQ+NKDozl1WOsjl1UwOjNPyQXVuN7P
Z1fL1+5ujodhSxkICaUdIerFR9P9jqsXs7oDycAbtSjrPXDFA6PUXCQcSZBgQq18
9PIN6Ztb64hgtHqz2meiWH5cPfKovxqzI75ut7cJGSXPZBQhew8A23aOO7uDxAqJ
FooTLVgS/drL8HXtsK598UzpTeGx087EYKoMFobPHYKyJA3RTWzs/4h2YS0d+Mct
s79REA5EIBsyABRj/RjWFPg78n/6bJDPURUgWE4K5JNMKPw22kPd7E8aA8Mrlf3U
lq3nmDYvhN1Ile/hef0n8CXEPDBBtpXFbD3eUPC+PxxRmtaQh2tuOywPGWBnQaXR
Wz8TU08IH9GzVli44thy2QDswRNbC4OQyAfwcizBlrW2i59abGXLdx+MHcIUptaJ
qUMEwTQmH735zxNwAto24LrBIJSsuYijw33Z2jQP5rLEW5C9Vii0z8LG2LQV/gMr
3DQfp8xw03r34OEMcORj1+cEKCk/qNJGlqSXIfDJVYareK9L4P1hxLq+NKUqu0nN
oC4L5vrgUw4WUcHVxdmHL8RKWU/iYvheSZLF8mHtAKmrCXiMNRh7a1d3M3LytTwB
wkFzIiOQPkbea4OkNNzQ7ExPCReEaUzEpdMQ858dMRnnBn73f3GlPzSYkLoA/g87
48S+ddDQPuL/bUEllbZnkeEJ7Lphwr7K5Iv3EuOjf/PwrZ9KzQUuD8tCIC0+5paJ
7sdKz4NhAONp89aeumDmynlGoq9x5/CpWEt0Psx4OH177R0zsPvtlWYojQg2ak4T
n965iBxcVsmakFp+4FJQ8pcy6JrmLa+u9XnkC1VO6Oj3eg1yMyezXfJaNLCy4dPs
0oHJzZUVnOmTYMcJ01sjSfyPwg4nn3gdlYfbhUcvvylzqq14mpAiUhliBWwQaeFu
3XW5DEoaAUnZXtiGgKy6AQFeJ5QLJ1eOylodoWXoxsVjdlxXS120jyoJK9m+nlFh
ta3snM/KL/rWDw4t8q7PpQ5mDGLWo1wWMwRiZjoW4JXN6pBghF4eoNlaDM5ak7ar
p2kNHkOH4+PwGEnw33Uga+tfD85b94mga1CT2jLXB8fMt/3lkIQ2C8LqrBVsAC2W
maeVUb9iF63yAasUK27L+Zb5pTtegdzQKYdVySHedTWRTXvQWWDzX+2pOIMjMOGH
ER6NLfsgnsu1zLyZ0Dfl4aXVJPhlL79tcvNiQ/JvygXr67WkYcAZsv02xAFQMtik
vdLvKx7SdgfMXNW+XBZ+mdd8clMo6mNEv9m2PII/nlro/5+RiBTZNf/RCO9KfRBf
OmxS+POdmBxYNnXIJC40cXhOpzgSm1nBuN/5DnbuP/TVT/j4+lAA5duBmyLp1fhL
tqiRQxbARx0B7DUIJePHCCmw01iJLfwVx0UC+JmOGmoxIzoPj3RUnLkFoYYDm8vt
FLRnArKOQ21ZcM/+zOkLtQ/D4VAEdtCODvyN9cwIlDNiTIR5wmU3LzlcolA+xYMl
7ef6+k0Qhr0Ob7OlmxqD2qWljVqUaN494iIq0kJaDqYxhtzJuVdictAgES0GP8uZ
Wq4Gm54hUnRHElmcQxflH3aZdGcAFcTpwYOJtArxlVWRUPlqsgJ7ND3lQCDKFYxW
qxBThYTzjGaAWIFUpj1ga+VNC4LHW+O93HETRDKHboWB5fAdrNh6VHKcPz8gjnWX
ki5NeF1MfR+qXUNdmIwPhEx0TiiGk5ARNdffZ5ZoFV5Vzn5bTXox0/Ob278x6k6R
q8Qqa0qtqIB9vDuuwmYlm1C59IHp79PtKrvursCQDrSc0I+3BcONHz35Yi5CmhPU
f8FO6iTv/MdFlKEgIpLFqqLGcNCESHw83iRR/y90YaP+bgJD9PBOCxaUsq6pQIiz
nTDtT85QO+DwIT/7NqtPb+sZPpcvj50xhiHNDuFMgllREQ4oEvb5myvoPRsTnHZO
aG2M2CluHy/YA7Rc9IkGB1xY0vdlRcEvqHOw9wHchkuzYQhDfPeME20Ig0KcmrOI
1bBIPE4SbQorHa40zuz/PfLYr3v0AeoCW8WzLDwtFj82F7mb8yfJViCR80f3wd7/
Z0mB6hA4RscRYIyd6m0nzdkRP+cLAgC1cEYFdFjlu6fPehhDkaUv/QktxZnGH5my
nHTw+iZmITtbAmYoZx35aL7xTwkNFEv9gC/oMVi5AFrFveakT6XBW1Af6bH8Dmt2
WYRDf4zs3xWU1kH6BgmckktYHPZDpP4mKqNGa+3gSkLdv8LDJFxbbT5+vUS6Zwe7
Q5nqbZUSS5eW++OS7p0eQWHXMLHQ1OEf8+n7+d999/Z3K9aIKOpnaIIXEKjrf5rV
gr9w6nbs2T1uOfkcDtouEOLc41ZpgFcxBZJVvLS0QawP2k9Sni9Vg/wCrPgYFyfF
E0qtl0piCeS8tZzOP/P8PCiKdy0Zw0KQLqmV53QvyDE5AiTAIXmvZZMj7yGoV3sv
3ElWjJVi4jH0+MFLI7UvMXy7OYLFHXlt8ONUw9Q/ZW0vL6veIbAOKIHTOCAbIIkx
+oZxN/9mUocT208uWigYR71TcjdhmoCvLIraqNHt4mEetzK6AMmCI7NXMNaqsA9i
sbBc+vKh6qp4mouzvvf7jZi0i6gR3CgjFSzn3Hduw801e7FjOb59DX5m4RafFZEa
jSfIvgn+S4UUzeUK0lRlpA8Eb0gZXj5NSfNbVAQhzaFYge/H7uuESTa2ET1+zuvP
3yySzi7MS8D9Y8s48dzmGSbzeGlhHUy2inKkSCMdEvSTay/y4oVyEf4akZTeJT4m
oRFtzbCWwByv5yk8cLbn1UiNv1bBZtJdJbCrRyHSY2ACSE34iRgyvmM8CSKRdTis
WnYHkTWiZwgygfmoh1uDf46Nt4dxJGRjK+xshp7DjWx/Eswt61vVIIa3SL3nz917
yZDzMVQq7xJEHTWGSVB+CrIpB49Erz4I4U/Us5gNibT9QLXkhkl3JweoBuzPvxGB
L1e+TRvRWLBF6N/iN+aEDHuPUHK0T1Qli2mHNxq5kVIz4jePWd76GVZIRo+MjieW
X9icbjA3k6OreoPEajlmcsWZFVADgdS1imjSoPYowVa5fTh+OSybW8cv7tXFbzMq
ymzvzkJnomObr1HRjjN89y9o1kfHrqneGxiSFzuT6OE7KuY8+Yk/inowLghP5n+V
9TnVoF81R3v0Bouvn/Z/j/lGRmO2tnzPKwuWrTzqkkARWMdpAyHPGK7+ztAMKRvN
JqlTVrmP1WfUpnrEiKh88QPmlLyf2IuA1uPSsHOjDfGonL/Y3Pqj6oY1n5gN56gs
fcmjRzRVBhB0ApcCOpZsVPmBS47+hAa3NOZYFRxiieW31qx+lSq380kqacW4EoGw
e0qFflnLLLRysyfQn6zfpAG7H5jXXSHY1scERYnrZor485vNOsaqFHhnMql7kw1T
ZrWoUTq+MMTEs/yq2GO4jpZfbQido3LjFM8zc1YcYy0CSujXkDSOHYT23Q1WeyLa
fXdYqP8yyh+xVbeftsPr95/7FhTvx/J6MzpM5MSFE1iMYOzHEKt1ClyNaoT3cW9J
hgob/BFD837mYGK7UAbsBTsqH+kzZiX8mEFsKPM+rbycY6FGihkezIjXIj9lC+CJ
dYtcHeSUDjePwSNT3iAj/+sExukn3zr6SCE3oDueOvFrObs0kjsWseqnGOIVsBk2
bjTMJ812OdOKmXInRWgs6S3dwkaQeDoQwki6KEc67ISa7Q+kbmskjRtt4EZa7iaZ
knvdy/3yhw/GOwa7eFjCjS8giTmc2vg8g/7Mb+o6FwWds5cop3jn1VwIG6QXl1Qp
vFmcwKN0NOXT6JyrnVHl1HWSgeb7aj+uF3X2iCiKQfGh2oIY1JlQZVHBt5FVGhEe
973r6/RoSDMwuH4GIO3jild2GYcwE85dlUUJp2aLuGtfkSJETwVqZWc2uJEZqpGo
QXWOgH3v7oy/ya5uyFuF8kD2PkCGdrt1Kn6FtRYdRHx6BoekDVpidtxXdmInekZM
pLfB9ojKaOzZV58i/zp3i3IIEv+oAZxJOPw1jKsCCmmH6YbsZ/ocB7/LQtYmS8Wo
FgQ8+ABrV2q34oZFennn2O70u1GogPhnNFX5xzT35DxJF6oMryUWK/ugNZAPRwoS
548G6FMjxQ8U8nzkY3LsZPRVWOBi/euPyUZs7kybqJ3oPMJ8+k9oVO2X9GeHkWz9
fvABbuKwSS6N5v+P20KA34e+PPi6j2oTV82sBOVqF/QYlnOaPvp0cOlhMamptKhj
+qWKXTEJlqE/CXHbBlrDnmb5ZDPfaIH7H9RKoDN5MdRnmbso3r+CNxXc4ivMPXFQ
V/m67jeVsxBX3hJfoETYy95lPwiK17lKuthZ8rQ6THhUjjIaHPILZWPMcnGTukMZ
Sd20jQmZBYjeUcCyom7UHOuDuGDMyGlXUJ4PewQ9IH8/MNidIgQZqhzaFc3h2pHF
trIksWkUCqoK2iUBPFyfhIdeUhZJ5N+nf6zhb5jegNy+AYsq02YDjIUYxfw01CjN
HoO6auWMpdat1X4dh1cx2QWOMfVUB/wwOGzJY540h7ivMo6BpS377Vi3bdRNNdSv
a5C13pIDTvsEVSVTBV5MsCbi43kWyG8iLXd7/3iHXO14B0J3XBPBna2Nn2cZQiNT
QhDu36Z/Cmwe6S+F7vSWs2CIFWIydKeqyMTPsroN2ioSbYNNnbuNPxSTnjbpIP9I
Nk/CsrCkSSMCXs5SpMrZ5sYhm5JrolL+8hosAUSatSkDagIGNYrLXbBgC2nTJ4hl
VfJ9s8TvZ7itf0TANQAH2WiLMf7voINQ57triOxznp3I8+puaUa6XtFqahkwo3WA
VsTK6N+r8dNgrwuSXFNTXHrPph+8uxk0mFYO17LWFGACqXikvmxwquRk/DQm2gbi
QAxg9dPBrW8qBMW7/WhIpSC+u2G9t1neFF7KoD480CwY4q9skm5rQofthpCGwUsC
7At51oPjYWAT7JcWAcN7FCs/zPyTcmXP32mu5NmsqlPglumS7HgRa4SGgLsQ4sHP
DgD3YHj4eKJ8Ur+hxt02+rFKzanOULL7jUBOOkPDvSzZANPxP1GWuUancw4CrooX
GDwpiVTvRelQvQsb92h2XNzikS8xTJn9ooBUqZ9TBp/k1zHWajEQwhwcQKXKwA84
ZITmcbGXBIO38e5cBs3rQrfpFK1t/7r7SRjKPLSaTqFsdRqSXCSudB7FBzlU+4Th
IgonKZVzxVQn0YDlxfoC2bCaJjFT2oJjYqx4NziCyxAGVbW7myo4h7/QVDNmVZLD
gDHZEyQaPn4GKt+kEtCVdW6/Uz758fy0jxnlPxHqLNhnNZMShDuLllIjPjw69XcS
xQposK99GAJbU5PIe4mqEm7kbGeaS+Aoc6JOKv1TEVGlPOA3/0HR51+2b10pkIsq
zFrb6idh4CDetxNy59EV3zO8QQVUUQ/9ufdLR3IkyQx5a10vm/7pY09p9RlkUOna
ePTM/Ae7MMCh+g8OGqcXYbb4UG62CLTnvtCe+Qcwb49IQmoNB9r7Tt1Wq2ekoMQX
RTXjd/v3ItQFIa4YiK79ZCrsdMMviwEuktmIy4V25cMEWtmYgsXOna9NQql4Jh2Z
/F0B3RQOmO0BdXzeClvi8NeTHTmgVhgAoeU1k2ZwkY/ReZCJxwYPWtzYGQLt4muG
UdBSEe1C1TlguKKYnStF7GOg437UtRtfa6qQhpkgXPrU78rseKS6+HADm6Mgtf43
O+w1JDHkEVNoeEzqnIb38/cQUouZw1Ebv+M5+TQPE7IBbNHEb7hBSCJl7Jgw/laU
H8bOBffp+7MYRwd56d0AM9N60p1kgblMO0RUeQ4yQzdgE2kEDeEDbQIspJeDP83d
WoaIU3TCK636VudpGdx3DLewYMHMDur5cndmSXZlGVxmD9Amt/gr+QlUMy51ZEWF
CYmErgrddnaqhx+dknBYuSMEN5Lf1Qz//SUNv80slv7hsRmJjHGI7KVCzXVsL3MV
ZAB4fY4SNqVLiIax/Tca0My/s9804g8RnV9mb2egMB1yi8wgmuKV36j5aCT5GXVR
YihbyV/MIAmiXEDTMjSQEozPuWK6RmDDuFPDICZOSFvtOs8a6o233cx3XvrNR8ov
0w+TCMIgvRwVrNfrToaLbUmS6Rwbk7yD1rwBwZ+4wgSdHRlrZfDLJ0LEXCgSs8tB
CZ8m5OxhcRC8JngDYLaO0lKCNnuPmKGuAITsbW2dW3aw141fisMLAEc+DEGPBHjo
AZ74kJ8QjVmInJYP5xSHKILBAcOFXD9QixpXNW3HWGpkGcKwVA8w0ykuOrPKRZ+4
hGyB9GmI7mLQUypLPgTjy0ZdmlXBeJOePMazsO/03Vi3v3BS5nPEzaYpoTD7Ggux
0wtWlsWyPUcdMQUTdGW1BRUw1Xmjb36sEmFMdfdiVtxiFaZ+ElV7dUoS+K7doQO2
LtIDfVqCU9ib3dzGC2RVavTfiVyHBNuAGP1OrYvUHnZsemD9hsZ1X+ZEyNSj4AKC
+xUlfr9+mKFOkcpsf0rRXC2jyNrDAWYvlNjpbX8fBzaEZjrJdEWxC/jIflClngEn
fWiwp3H+VIfv2L8LbqJbfNjuKYEhP7aaPSPxeVfYN1dMe3QQp4u8RW4lXxq0Ys6/
GU8fTZx1QbmJdrwAW6nfynif9qvtmLI48NNX0TzmDwcvZgFdNfbVFE3Tb8EDFlrG
W0oMp0qkI9TDdsc0pnsTSfKFzdlFtrfBvUwFQO/Ryq6jHL8MBGZ+MiJmqoSCWc4q
pN74nWgVyUIDUS6drlEDbSnlYNEYcBv+YKgPZSPu1SRrfkI8ArPHM7y1lpq0fU/+
ZR3zzrzdd1QjTo8hBjysF00g2wvILL4p3LXBQNkMh0s8pAuILyptaL97WLVwzR1C
Znvve4igcb15C51DBAjBGMnytjui5vbRRix7Y/fgyuha8G5e/0/vShYgfh+K89Me
illIgjyKjFhlkiJBda2hDPe6ERqNj5K564UdTY98piG4WvjHQPDylPMhqfDAk8l7
rq03Cio79kOsen+UR9JPGnH3as3FiZGCshvnAKGJ91TBW9gimBBogsWBDygzbZM/
Q8zf3J7mR621vDg7zVJ9i68qnXYsQbhc/doD9zdd1EwZQfWua3aZBJQ8K7w7PXms
h1m+FPlhcG2LQXjZ2FpYK2Rgnt9AvSvDpAiTkOUlo9erfqUCBERC2eLgpXO2FNA2
xI7UEe7+jvGdFiUS88frVDXUx0jVKHrxSqrPEaSJSXbtOA8s0yMxyapXY3b6lOcr
tk2ssvkrxDRuUBr2g1pphz29EJYnTxv4iCzo6U082k98SuUJpRe9M8kTxJV6stqy
6oDsnErr1j9bcdvNg8D1pV+/eJ9dkQd8ye41e98iVKyHJyO4x4vDSBYFA3GdnohW
0qyM8F/bElLiw8jL4S3yoORDfxvURJNGWJdCYB+IvLIvm+doFjMe36YAT1cUiENS
cM/Owysl6uWQCItWntsqLdfXSoy0sOPgSaAXx6/Jf5/e3Q0vx4ifBJ0z14b0c0p4
k6Nq2hPnZw9agDLQ58hY+X4H5stUsJ6KWkJ23qrIZxFeMuB0zz3UzUwMw8iR/EJI
h6pqOywSv0lNBO7ILq4XT1vbyI0DCwRF/UwMFmnTHBxRw1mRZ7UYvkqQLkhbYAlh
knB1ANYKBiG+NwXd/+tnqj7DWLc3QMHgO15UQlceVhVJCEadUClUE6ZPHYctVg3Q
rn6qDOa+260YV+CBBDoMPIm+9hYgj05k8FoUweLcLSoXnINZoj2BReFX/Q/z/vxq
Ho5koo53n8Wy8yn8FCppMV/THipZj1984wmaclb29dPOs8DoMLwt7k8iegaqEvVL
9nQ9DgpIMLDbdrW5ujURPMr/qnFGu/t58ud38FVjtqHZLbsm3jJhKk28cJHfKRiW
A6rUa0tdoHYTauZNibbdVPPkIWFeYs49yaRPhFg6yCPBsVCQtphYxLlx9/uilvIl
lXDl0gRn2v+ZN9cYt5xHG5IxbE3hBREHMG4tjCsV46UC78Qq2BZBmFpD8AhcpNab
9E9TS4W8z7zQmkhABeJoUUGhCS/rCWBpIKOyEdCeXWfBtNLdWczOBZDzkcwGc/+4
2bwyy6eSuilLkfAdI+WFW1ORjtETu/T33QNWUNc9ehEuqjsYQl8/OHO7c4HNIqnN
1jUhtwW59Cz0sz/wc0wW93Zqgl2goBC0Cus5gNMrOUJpDYUAUsjW04uey+Ze0MKv
LkHjckc7f4MduyKW93uV5/LhUEzUMm7PUQoTiluuWl8R4Kv3n2WvaNmlatExraqX
Dh2gkT7fJbolD6gu+DQpLGUauKIuFroQASX/OzZlF3xrEryh+hCOJG7u/wuT+7ES
ZrcGSZpHCZOkbTKAH0gZ8DUKZjNZ75/VJyPJ09MH0QAC8+KQJ7d/L3ro3/WhIhfe
WqUCqKmIRZYwih+DFFBybiTmirtQrVirYk9t23ZXmcdGj7aiHoMl1TyfJHuJyWx9
z8+6KBsXWqZcvisNTBaJGEvvnPQA0ZB6pJzqXx3Elt68aOW4igmuBGJyDZNTBbtm
Qmm7nUEZYdw1H11qnK7af0x2FuNiLSPtmK5IcBH1jXpLR0X29A2nt9S4tlmEcU0R
VxSKPiyMJGn0NMFvKXl/ruqYsRQx7vcAtshiUQnJeiwkxI5++a+LCuNWuaLxHup1
XLsbW4ff1pX3STvz59Am8RbDVMzoivQa8xtO4XSk4PURcTjItWCbwysI8Z4NSZot
xBl681foGTaftbnoMXIQoPh5dUBHfM6eQQbreZA0hZjG/P/oJfPWx02gDj95qXiy
1SkoTbBJM8CZVVqje5xSsLPq/G1D13zoNX619RvompDB4CpYLiTUKM4jJumUp/ov
SXkag6K/OSVZ+8NTshxXZHmBZkcaTwginQbOhKZr0mep6rY6voi8g8beFA7k5+hJ
hy83PEmoYHvlPoT+LmyW0yL/lj3nzKTxap1bHC816xPJCY9sw6ItQUY3/OolL4mz
x55onWPdiP3UL5F4xS1bLCdBKHCJkErLoHnSw4HhY9Fz9DSYkQpgs3bxLbpUF3pd
M2O4x4GHk8smSZ2WkndxizXVCbyM5ZGy3bOwE0Au5bho+dK2V3zWGJWGDJEbHSQY
k6wXTYSiQopRDCi9DQMEbcylSEhX3NHnvB991t2ZzhCxtYGTcLg3seiL3ExuxYfU
b27Snl2Dr1UAsDhDGJVp2DiS/fOxarKQyn+UIDUFEFdKG0Uj7tCEd45ZrS/XoBCM
wp7Yz7vz33farovn6d4L+cRATQqFrvCIwFVIAOwZNUM4JyI+iUIGmLRqzF7TDU/w
Tr10yOWnxaaQrXB25aLYu/ciiwILZeVkpcf5Wk4XOTJDaofWLF4H2XsFzg7qDHcR
esi/YwbVcVfN+7IYDe8/wrlRkAxC2JMkac560liCZOwFP9+BkwdPkMR8N2zyZ8b2
itJfj/mWGRMX5Rncnc8Mm3reKpeNTZjU3fBtyNOGzCUFZT5sGrQqlzCNmHs8SAx/
TFFAMu02vJ4uAFlw3YDy4MEOuY5B2YXBMnATltXZvgHWWO6ZeV2isSoO6EdjHRYh
LCIp0i8uvqvDtwoDrafOrIqc20IqdlO1vVYi4PxvmhrLY+6SjD0btTOspDkfh25t
Hjlo10VVCnZlBeUxEyBU3hF3eLZHkHLGZOcxoRTJkwwiGnPZcAIXQutIiO427ebA
36MI8vSEy9wuZkVJ+lmRXGZPMg/qtcNEmCgxJ4Ud9nNeFFankn/Kpw7mY5rhNf3H
71s1a002a63eO0QrGInVePd3TEvx6trwCOimaKTKmf1FYAFnERvG5q0FySpnLt7p
k5Y3QS2C4S/T779AAwiHAw7fTSgwXW16CCk4fdXTrDnl8mporYs7XYGJZb6oQLBW
027ptLgVLP6BSd/nzBCh1/FN7IDSDmgxqggCiVi4eMB1x6+ftNMuwAWrY9ceCp0F
D+yOyEKHIZso5YviLO1LJs12eKo4U7I5FCTtG/eKnmeLqf9lgL6GEhFrdgxQ9yS7
DLmZD+2PHiQbV+wXiRoG8kGE31aqNXGEK3pWIH2VIJQDjyCgjw7g07IaxISQIojE
K+Jwwa9p0EvT2uxD/Szk+D6Z0hm+QeONuAqqyeNC/qwPjDswoyifrItATU0ftLGR
+2xHMbc7SYUQUvsypBmf1q/aRIP2zVfBr/CBuypDkfWxXzRB7YkoIO3H8ArgPXKX
QtHs7EYZtXzyezl5vpbeoDQHSBdwbhwIMMSdJA/NlfeT3NZNTnDTLCrNvFNwM6/i
TAhgHZoJIet5FffZMZAOGN0YJHWt6RD96qF+84bgpo5Yj14qZ1c8MhN032m0a4vs
b9VLkb6KRwNw+ra1rxeL/vMLs/jVxB5hl9LeYMT/HeN9pupTP5U+lX1bnjH9If/l
O4HiRpJ3mN3mRR4qpWg0qV1St0g9kQjnFiZUQRA9QhGIqSMVxKpQ6WdaflzeSzCv
Nkg4Dh62iR64qlnwmzpmr72PkTnt/8wXcHtnmQRXHQCaW9M7QlYaADzsY5fdUAyX
wkbpL5D9KhempGHPCUyr4+UmTynb+Il9m1PyX4j6FWqx0OzcR76k4SP6kQZZwX3W
DMlJ6wWw4IHcpVD8CI25ZUv+x2KqoO1G0G/svbaCj6iqB6WCnzL0s7yzrmpQZ1k9
tSk0LoqtCGScxuduOOy/Z43IxCk8kOP4G22AeHyLbbCQbFRcCab4XQpBJPYQZc4a
qrSE31w/j/jtYEBaFNTeiBLp06iM84KzVd5ihGFmPJw4plPVYb+c3Jli2TNB7kAx
6L06RHtIZ0MRlmbn+NBcwY3/jVkBXFuTpfK0AhOinGFgAbrHDWhyA80vVPAyY0R0
xWjN38vyaSrPVPbQMF6WDk4/gm+z6pee1iZtmh/c+xWfNTPMSljMo2bF4y0xyk+G
6zDwqyCkbTSJANcw6s+9M+80KCItjDMbuA+7IpwG36zAcqZCB0OcS6mBpNnBkeVp
e+mvLRWpHZjugeN4JpBRCheF0VDwuEiUYivuiK5q04BYO6QBa+jr7VV5XKuaxaGY
5SDUgusqAbrnGjaCtRe+NS6NNzEfK8FuY1w61uu1MQcg17aut7p91teGYZGSv6cb
fLxyU10NEtwbYdi0YIWS/2D102LVXD4P2e9MeuUNRDiiovsFxo8fcxzW6cKqrTl+
GFjJiCaQdcaWrBtmJWOLp3QsmUyGD/a1tcxmjIjyWrBN8HZLY/qZAIOWN1ptKQuc
Sc8GosD7vXxr8CQbzKZPmZbSh5gFEj5pAkxG0E5kR9RN9nzDHkbe945mFKIyB6iE
YsKFs+xox56FfNf90sFKVGJ0Q3hAAyN9uXZzAghUOB1uZHtDDbO7MN9J/TndqxKH
EcT9ymZhrXOez9poO7+HlYwJmK04XctV/hw1BKwNNxmTUwcgQhiPBN+gUcjnuKPb
y9piVl+BUI0Dqvv7WFrDAHg0trX/NQ8cu+SU8BamEQqhG3pd/xaF/S5zzvAM+Opp
tltEcszbR39W1H/wN9SnIryixlUzAFQxP3OjJLLQBl0OaebCIuNbqikEOHj1oeGy
6xwOFUOtb/zWxdk9tgLEocsILixBqFnJz2/+WQuAGU9lu87zB0MbGSJHLxKDyt42
icNo1m1taaTPHfL2VPPiPPsoLsik5eznNW/YLsEy5BES4vauSUvMO3EoJPXFDyu7
hudTqIB2/RDxjSO9z9tCyWVmRpu10AN/FgqZOcitPyceVCozNc72YmySvxrwk2TV
mApsRbEbRG9onlMQ5zhsHwQKVnjbkqB2vBMFEnD9o5sVDnhGFsRobqRKLdWbmyit
npxx3Vtku4WQ7GhP0Xsg0A7IdzH4GFycGLcJY/nTCEIKunm0BxqI2uwBOJvR3fcH
OHlm3frH4DJqn3hnXHsKJ5+silEsIzY8TYddL7LJR5YV69o70Fhq1zmQ0C2S5ZNs
Kzw2ENjlzRb6bdaqNq9kMHqNIg5Kr4y/zizxIPTE2Bi4c4y4LEeyhu3vMi0duJcU
i47I3toa1rEOjuags7ijdaGCWyci9sN/wBOcR5oappTKPj7/xOF+mnW+PXMBux40
iqBhaf5yc5nWojN3gZVG+KV0B8C8RFn8CTdayDKjsiWoVJdDxfXGoxo6bOn3c8Jy
m/FxaoRmZ9PfC5hkLL+IqqV1snEnGzXYjJ7C1GceZjnpuLHefgE9javuCvHjlABW
pjCnJbMIJQJfX1cIIx7R5okskdBb4bfZ5ZcQ25DNG3wtwiWBwTPAhAiM+uw4F4YA
N7/J0Bq1iwBxNINutFNM0C7pIxDwmx/gxm58pyb3jbuhjS7aFU7AYM5VcDC4RekV
H+XVG/phfXymd/IK4Z4P3hKvwL6DZUN+aq0w0hvRqd8WwQczrNewDESfhlv9WkXy
RpVPuLOaava/PdY54//UPOv3hW5mecBCpb3dAQYqQvjFySaOvxTmoUAvqrSGykS5
eiaFIoiZviwcffpDEUB4D92l5dRIa0iLYkTGatzluV4VGm/z0193QZAnHzNzt50V
GEGJLR1pwJMZdBGuaZQ2x85AnJQ/BhTUaXszdZzzVKXlBIVOBLW7gg0fdXFt8Ts3
IZJYkv3r4fjBunpkJpUmBC8grCjnRB0zmtVGSCJoBflDDbyb90Z6O1qYSSwRX3CU
MWJwEop8RO1du0t7NOE1FwybNWJLBLsdzocei0Uvu6DIc0eWIDMPtV8sqazrIaZB
jXM4zbnywzVqKbMjq4GL9xP7HYXr/cMGwCYUcuQiszK8PKfBqDlQQokkm9GJ1mdj
b3iD+mcEci0VHjY3mDOBiUTw0h3vVG0P5rpRJJh6KSXMKEQR6AsD0PElHN2VMgq7
rXfc1Qjo+u4oQ6wyHeGXwWy0IY6gn6ZALbaTp7m514+eOHkkEx3C7NUMR4Bel/CY
ckH6R/o5uPeGZAzi3HCzfgsM2PkDc3Gfzr7V/TtJiuRGpIc2egE3QmvtoJy9xnJF
9l2mksGaQAoAQvL3t2tqzDCP5GMqg0QcmcacsIzdEG+yN5iB1/oGOv7/NeKMv9Dh
gheuHoEHM8YG5v7g+lmsh4jggp8Uq4WCLc2Qd+pbYWjN7Ud5LgRzQl/I8wt7rEtq
XfqYhDol+TYxZCTtcQEeBymvI1pLIxhszKOV03b/1QelYl+v2B8uwx4rtTTVHzPF
gzeEVmmCPYwZ06MkX61RypZ/A6reQB6J903sGL/Sfkb15tnZ2+Hyb7+GeSVN77yc
EYoisvDfoM4pDCA2KgGp8a8woymhTEm0XaasbpNiAUwZwwJv7xqcVoKfHUWMzsmr
3FIP7M1Ix2Lz5v8MmF7cjmiFY9VizhmoS7/oTw2wrGWggFHcEL8ZZ27RJPPLDeVd
tiLumNT86BLmUHylofi8AUaC3CcmqEdO/5gFcSdGmf9OzmXg2bGLDDCOa1EvJS5n
HzJaowlq0XjwDT9c8nAzh687awleNM3E6F9PcDJ+sNFIhriT+d3isfGqjA6OHmzj
YHDVpf2l52AaMK4TL7UFKNeM82v8J3aqLi9YHX8Ktz+iZmgU9f8LxVclonv4k2VH
2WJC3vsgjsnDhk1NWuAdj6K3kCbfg2rsifGRQnTeWNzO5awvLWoncCOopnwo/BLM
IO7KwT+aG4xMIybJCx8YngzqmqW+PHHKRjL0/8/zyQeHv3q8MoozOQQc8j6kau6U
IfbnSRBbHniwlUWKaEha9Z8GWaKcuDsc3Rk8cossdgWohDIwGebOEIUYkxLSS5w/
wuoeX0zOQ2Bhj/BnJMJQz8UgwzeW4TULxp90ZX0Zyz+2V0danczzQ4Gxp7AlFrND
hxivzybSN1tAl5EkG+gxskfEhXu1rZ06uRuA0Wdz1rS3yRczfabEnZwOi5/YLnLQ
UuWRaA/KK1WNvpNTdpOqUdP5NW38MlSmw0Nfuai3Jo84Srlkjonr1tbUAU5XN6Mk
HQoINItErt2efkViN1vzGcCA7TRpW1knKBH4WzCsDgfpJKalr2vu9lT0jKwbtrAZ
kg0Tejcc6rVCE+se56EoUuNPqbiwtXxO7v0w6qJ1MmJMAVn9nlqaIPbEnlhWxB4p
ckCFpYpBTuB43P9zF5JuYlUDIe668WMNcsyydIuV8j3nLMcUaN+pYheWy/LijNCb
kio7xoVdNIyxLr7onpgXs5NkOPDiFdGSepz1dme2ckwPuegPOy5ND2TzTSv1s5g7
SggeVRYlnakGv9BJjgKcPwMjo7GuXFFKuX9xOE+Z2ZFjP8hzk0zB/052mqRWpxyw
DqAFUOOAGlIbVmDsIC/Cfmlb0Y34JvWUWpS/KgFUxhL80+mipBUqaU9X97e+fhbX
iuP627jCWVV4VKGoSVLhi2KKbsWHuvgc1SrH10h12wiDRNAmUcoLGpog3dvoO8d6
npULd255oeI7h76W7Uhy7FvLJTOEd27/juWdkEbwSsQR4EVyz+G2D2LbTuyufdYU
RbjxqpBGPeqc4Wn0PJ0ukOKsKFKOQLD2mVTErB+uZdbCql4XXy2ksn3wJeEgTMrq
O01q5aPo2UKlqLvAQWGfr5h2lDJt2zivmyoW4UHIzRQHJHLphOCb4c5zEwzGzXsk
EfBF8SJ5Io8LVEHBInX2aQKKaeNRO4rpzr1/IoPJiaJ/QOiVXV/ZW2naxdijYX5I
QAqVfHlGinZ7Kj/k+dxHsWJeHVwZHIb9YYGuscNAxqe7fJMYVU+x1GjY3zKCrV+P
ZMpA1yNCkfoafzhoWa6FnuiuZPDRGfznkSHjxM+nPbnVFWC7BoxlTrZd9F/qPbsb
eKp6+AiisMHUuAvWK3yH/eNowNf6GFL5ISFKagv/2KIVp0/wAf9SuoKzpveZIrNB
kRDRYh9C9FiddqJk79c55jy6FsoUo94lpVnQrCdVKtL1zIJ4r3xrkzVMYIzw+wgr
ghwodiAhNQ4Ca87Dg/kx8kqpz5nu9y/C0EF8Nobv/pG1KRrStuROQEpnxH1y2PJ2
kk0eyaduTPJL+iAibYQ+V6a3XTZG0pWvtFnwBFxySK+yB3FWwHNxQdeV4w+3Jqm+
R59FYTfHaYYkpDyMy74+XpxFyEriUSnkRx361oNzM8qynsgNc+WoUySj+Ypvh2+u
8V9/P3+7aweHi5T5AcMabSmUWu7V7nxvjEmcEjBc/LvaYOeNgC2X76hPWoonpzng
t9tD8un1HZ6AM+oL5bNrS7vpTgda54YLnKU/C3B5JBapuCyzMM/AolCzi7AO2ATf
U/5vRfz+gtLrrgvgMy2Wvf6rDGqclA1A2MpuDEfbPf3atW4NCA0iMvJjpIa22J4O
ReC89MsCpP+a4CrhoteRTB8FraJt0Jt/j7cwB0Ul91cDkuRg33iB+ZpoCJCnGMw0
HdeiLyCgdWuKCuyox1pKxMnvuPf1smEfKvfwaUJcgfdIgWg2gSaWmqoe5XD1KShx
lkNyyYetbGNLTnHNzb/K6noNtO3/584mr4UGSXnELcP/i5HvMukGiatL8fiBEVO0
B01h67upWozSGOiRM/sR1V5Dybri4sdlu6cZi1zpUQ5mZnzf8Xm88Slot989+Ckm
fh+kvSZ1Pvrd5VdJJqYWt/gZzQc+QOhM8gu4Sjgbe4XsVqIrJrXBUlu1R6yV6DCt
5Lzm3rjsYFh+u+DlxA3gdKHv38Ven4gyjzTGn5heVaMw3YfHK6hXSvhcTItT5BfQ
RByhZ2p78N2Z/nnkgHxr6URa6miVnkzkI0E+n0dn8Rz7w9xDlsE5kyzwYWG43lz1
jXJ+zV3dbqKU48kVph4C5fvyVf9P5YmmVVt6YkedSvP1NvS83HDBe4TFPDcJ5iRk
DYi7+DeN/QhOoFjcnf3FWy0XSDnWVtS9+DAX4nVEt8TI026RbbdQr3Wk8ABH4w3t
ztwxVgpxx6+c+NA9R6bDrHw1byBOYDbXwJeTDKPWcMhVzkppUTdhdjLvOqLS7R/4
hLgeNLz6MTewxmLL5nNhWwr4Ola/D0Qepivs7xkBdT5n5tGDPJS5wOL1sRWuDCS6
s3NQq0p8606wc00rUfCIRe3ern9i/ptO6JALPSK4yMCgZK4I6o27lxenKnzanhqb
NyjiClrxfzH9cy9N/xJbbG7TOzHnq9ChYbfzbnQO1nplZ3P9WFPSMacR9Pg7AVtk
Oxzd3UnYtGF0IQofvQQ4bqlfXJauBJh1tjwFxMqgVPalz5Ilp1nzcUQEqVpPLfIB
QfXr1ajIB81eVINAuXBzvIN10izg/+MKYiN7v8zVo/06uANdTWrO472wIZFNpADp
3IYuh8FZStw3MdpwM3oB2WAl97InR5+q7t1AOyu9thRHJmaeoa1ZCl526u5bY3Fr
2XCqZfh3B6cTQjRnIVy+2G7kQHL7DwQWimiE+FoxIou4AzBOh/JZ/WXQDswl6mUz
+9DiIRKI93VeQgrumgjLgofeVurhu7O9kxo6WK382HfTwhrMkhJe1nmmhWfFPd/5
CaJfbqqWXETjNOOwnJOkm1ADVbSFsH79gz3FbrJlXZ+vjk3KDAnWIICwNdZ7gGC9
TXresXNIcbWpoU+qY9M1kKnTQprPSIlvDwRtCZM+6InTwpkHwOfwoRHzK5ONblqn
v1eKnX06wgqBFBPVAvW2gaYiOHivlMUcpgR1Fu2IluV5BsvcX2Memx7v89fb2KgD
YIGYBGIoMkl0nGtaII5/ioXCdzw2IGCDD6JhGcMKaaTHgCt+y6H8BxThNrktQAb+
lDOq0vnBWghI8EvuEzVPmraCL1z7c9bKYvO3kPpy3kWnDWNrKK05inapEBa01IQZ
0AV7BFNJmUQeJNRTIDrvrYASy5JqquDnP5h87LZ5sj0bQFNQto8rpmAB7Oy80qrC
lcA5b+xm4DVbJcK3ZhlnFhD14GEE+aFRI6HJkHazGj8sWgURga75MItxpdIGrAWD
jqQ0dUr6+5hFtfW9AQnTxodjqB1n0KvZeAPNyiL6V3AXx/ePZJS2cCn9cLHaJ4k1
2WBcC96l9TlTE+I+sUjUelj90F7Q9MEB6Y/FvqykLEL9+2x2bM5gL3j+b7qL53HA
jTPSo7GfioBCrxziPLI+t7SwnH2AEKXy8DhNaTyhmNLfwmmoNIDqqVdhG1c0U76y
pE0b52Mx5Q9R8a1i8NLYoPwyW+Z27c99N0Gfyqrjx/xnup0PqEI/3sM+nCaZEzio
WHhWYbj2dEAxBBMYm+ss7kITs0KqLRrlcYE6s5EDT1wYkgLX7vmMfAehzNvwJ3j5
QJcX/R1oGU9CDk1CZCAIARDZuj0bv4vJMkNqGQGc1VldIi9ZkGEjEKneNfUqy6JE
kPIla/bO65UTNC3G99lutYMoniBQYTtx8FZynDOWIQGIgEBNAPn08SEYA5Fc8hFW
jkDHZQF7yY55l5KNMPq8dhBSYvOA3ZV2e7lPdRc0zRQvYVxD2Qb7PkQMAncPQNG2
Oe9WVIJSj27oLlRBawE0Z6Cbp1YuwwTCcRo5dO2/rh2cIV92UmATIi5yDgJHRST0
+njKz352DHajIuEbhnnNjbdyUYuDRYbV9j201RHt4011HWv/m8e7IgTdBduVx+FX
p147/pfWcos799QR/snHjVCzvh8fsEkLUlq1qeBpTcwmboFtgUHOpR9Mq5yEpdzr
/2ZoVWzJXK6StJVHBbmBRxnyEYiLUYa2nu9KjGDAbaXMAVqN597Oah/Y30yxNpp2
wm4Ln6G3P22wptw6CnnlBm2e20NLeb7gInAo+M4PkeoH3ohHNn5U+RG9wlUbrPnH
Gf8ddPd1yoD3fUMXhWEi7Yt72jtL2xKtNPuItsCZeCiBA1I6wL9fk++pKq7QwS/c
jjwuJUgPqkBC8ft1993n2hxew0V/kjZ39/iIeeg0JPAC/7Hw0TifD6DZVontqDfw
8U/hLWzwdaDMP+UsFDkgLUhHHxubpmNc4qQwM6Huyom9dgOoloK2czOLzJZDMTsl
SRIlz+93+g+z7PLu5MLpzeYJMp5cPuyjlV9wVa4li4qWK0andLRfJ1JsIf4IMQFP
gVfqa+0vawaCyS96I2E/ywSvT/Rz07zGFwC1tbIusjzc+20WxwcdQmHyI6gGlyY2
CRsJPon4X1zGNA8FwkyKwqZnU369HDp4VGQH21ZI+5McjCvWBGCTGsKiqs9Wdn6J
/g4BnF+stek4HubmQFzBD65WF8Eqong0Qt1Bpdl54JE/H0EA6QqRJRHrzWZhCkUF
ILnYsI3l1fgP+jjpoM7TkdnEUREWdcvPlBsgMlLcaesf0GEVMqOU0X2bUIPagftJ
rRsHjjPzPrrpVS8HKRqh0KOCMSDlQ9SRKchvwdhkDiQIxzOWne7+QtexiH5MCT/a
ven0OM0aLNdeV0t1rlVSUR4YGJ0+B0anugF58OIRWSSqJefCYCk0hlMhCiZoV39k
To+Y8fVS0ChQLAVNEIjzVrvzf0OIGRFe4WT3TCruKNxuJ2s58fGPK3/u2s1sLCVW
Dwj2jvDWx2zLsNpZokAKhceoq/XJsJJ51dPF3pMY4Herotwi4D0+Xh+1moLs1AYT
CCveYRLP0BZKRpo4k+iRgzpbskEn5HnyNDNUzM7uUJphs4le+0Jv5H5bCmifBLKr
heIWBXBEAUrZ075V40l811QsYjCGz2ZXN8iRZ0bAYVhPIfrkQ4qg6RMpTqJxJPUg
ID2BxQ1wSz0FuudMkHrTgmSd6PCiOa3utT5AMx0m0UoJDWYtFeU1aW9+/UoVCXqR
nOXXAicJmtEBKrPsIsxYdxOKZxswTNDY6ows/dsYqx4Pc92GsnptMmmynrxeI/ib
6/gzGGRJveJjrYP8leZn+r9EfpcCQMjRMMp6moVOnw9IW1223hVDUB23Nj7Yzgre
HphpJePU9xOp2z/3RjVBgAmXvdhdiWc0mn/I1qmbY35RnyZ367kJpeYtc4quf8EF
QUjT/HIWcmkqHq+epp3/3xc505FC1Ll0yLqPB9CSmb36Qbt3edvK9WIpMoZyi+Am
gXd5FUC2eShJmkWfkOAZG2oDo5T4ruopg8byvf51bUc4fhrPEknMMO+rckqVW9zC
BY37dF+/8ut/yeh8BgD+4gnSiCrvLdGdwfKVDc62OHuwYicbI2jnTdrI/bcxxFAJ
a31nsZShMdRbtJCgVBf10w4G8Hk/vIvpc5UlFFmZ77lK27e1f8UAvRLIfqJQsFha
UKHOVbWQmAUd+yGCV+vwCbCu7dSdvsD7nkul7AnzFjhTVHr05hh08exrgw0CQfWS
Nq+DltR0yiyflGsez9MZy18mK8r/xlV9YJk6fUXwhq/3XVY12LXn3UsBSQWuoh0f
VRV06t2rTgJ2NVyBvzJ/waf4ILuel4d4dbk6Bu4U5+rmI4mKMMp+xvHuwk9XSBz9
Ibj3f+Xp04J982DvrECXG1m1Kz9QyibnuCJqS1ZR49uWLV1KE4B2pA/AbqwjoB83
AT5aX6iPzQLBEizaL/Z4hb0AL1XNXR099+m14rqLCyrvRZtyT4KZyzEDJHcp9brx
Wv8T00KEC7RsH6van1dS1CV2yWVK1YIRiFuSOHsGAjUibgPxox8s3HMDDLSvamK5
XM4hlYruChB74UXWfscLgip2Dv3CmS2VhKFodQ8o1v6XV5RtCcTIwvgjk6pRkpc6
dyaukQI6kVhYLH/fGYiLwpGgC69dkG4NzIIYCGXGfMZSQTm8zFzTHxVI9GvgIqOm
dz3Vb6STThComxOm6928sBPuJnL4bFAeNaObxFCg+v+HqQzgTQI3eTpYbyP/jl9L
JSkufjbCwOUoptQw3xC3BQKUNAZGgW6QF5TWJFrPDEqWX8P2ZjI0dbsdqEXqcQ7z
oZbUFKWYO2hJZFDi8bP/SSePeA75J2SNw5W0DM48oawtbXf/H6m7UDIErDF+KaA7
CjsM/2yk1waYaZkhqdm3f27+YkUOJLmGkNMJo3FRMWk1gIzbt1MRhZPNPa+2UpQS
brpDCsgPkAUYxsDxsHW3R+rGy45quN6bVbMLF2GZZGibA6/uNRe2ULDpbTuAl7NQ
041IvzWd+hn6Zxf3bPZPTsmU/ueue3gXmum5btZWaeb/6Gwo24E8ojsn2/8n51JG
zT5Dr2sDY1R5+jmUCRUR9nN7ZOc72FZEI1cuZGXo+Fl75remfIDiheqeabKEtP4O
phk7j8AL7sPiQ1IuTC6wzPaSgwxbfpmDNbgpzVRXY0DVHdMZvu5yR8ajzB0euK58
RPhXfiXQEIxBXDwLseDg8W9X1tlht9zf65LA4trJ/tKxl+FLEKoIKkLGLOtLufsA
LlFykOSPfvUKCISLnIPOpsB7VKbE+ZD6THGd/wUr5ms2bqCkDJqxdx74ZhC+8vG3
KnSx2asWu1CrlmcpI02rsUVXm/ejp+dBC1qTU4iGuFPjLUnDAmikMeouqPf+/oex
Lgb47T9xhVSccU1bJB1/62gnEMpH5OFup+Yk7pR47su06ukB1t6FU+hOM4V/appE
arJUac8N16e/cTqDXAJuL2NXnRWdkxUhQI6P4sVpFOzP8wxkXGtN6kRU+iCwc+gi
EtmdxlEMKrK9YuxTjzxBs/YvTAqKBQQwXjWPY+btjBUHKd9FajMXeeGqRQQ73ME6
/d3GV6tI4K6w1IJDgFXuhm1jB9qVm0XNzmr6XlKhaZaM5fGXTav1YEdplM0UUOTy
3B72kmOBM8XLSrqtgq7I0J+fcSJVLef22SPU1H49088ZuW+Z0hkkS5xUHlNfat/O
/6GQrg++9JnY1ntAHRUUTOnMBDDljTmXoi33Ix8kzJnQkNE8zamgjq2ANcbGR7a1
KFhFMyc1rD4VntmI/+AK4kC6yKKI/U/G4SYQgbWlPUI9QRLknrR6FWBOKgHWbzzj
9RkxNJ2rtXEyNSSq2qX6gBL544eFo+VGS735O10aTWh1Hh6eZwMu152+/zkVWsxs
MZ/KBwoVT+poGW1SEQEUBjbBUJLHH/7hm8pAI9y5+iKDkjmZgsyxOOEEfnXVfdFW
hMYapgbcc8zUV1rgq3PjMSJzk5Z2bT2dIIl39XLmt62he9eXGToht5Z2JjnAD5sa
e5FKQLSBWkNuadd2Kc4YOmSUabeZKjkNenzReoD5Oh+HvoFpuykCQX4Z50pcJ86E
k8FP7o4h8xg/34VVME4adnXOWMyz+fdpE6p1lHmJGOBazoRm1vmO38rhgzKTBuCw
Klgs27QylA5IAjjIiMIaiiRlFyfZa6xFTJtWuPhgxeUF2IPXBD5UDeWMmOjWZ3ms
W50YfqTViDYsazzeJ/XDtKIKVKAs2diJqcugJx8hVjkO0hTZHJyakT5DnLnLSOH5
fxwmdWjFrRXUPnRMWJUQOalNNW4/yILxDEFFVYxbY8hsezCLQWIl117Sa/IovWSB
GcvasT4nMNwjXaVo5WMpJlJScJ/VzbPXjRD3udO/lbCHV0h5hVXb+hmgdaqpgOA0
hOTTOIK+CAwx2q9JZDEKJa0IUbvHhyQWc6J4GMNYjvvGecwcNXgGv6SHjdlWeP3y
HDwLJqYG73lz3OiUPdDtRPJ83YKougP/fi433e77JX83T9+VXz3oxOcfD3XjvBnS
ewleyDoPbzUC3MmKuhJ8P37PUD/U8vDMfc0qZGZ9TOLaEECc8YLSVQJJdu7mtI45
FgG5CQYmd2/vI4AxAWjIYPNbB2mVECiF9ip+Hf2lCFz3u5jVytspS+NPO1fPTfLu
NOWjyRbt3MPMFwTeMm4FpO4cmkRH6zQySVSUQZPfhGw8uI4SydstrY+pv02b3o1p
UCDZsJmqpuzgmofPpYP0CILUNaxU/6ITw2e/0MiYMVVP1RgMvdm+iSTZNJafVZwX
JtC7bPQcHMuDE5u22HsyVS+1Jl3LHHTD0TJPmVNiGaQ7J5Gysb5J368T3/Z5vK6N
YJ51HFPIZBDEXdn9KZxF/Ei++XRM7SK2JqPu3DuEOPpf/Q4zhOLVE4riY3fLCxU8
CBNPh5euszzql8zVasmVO3TzwHhNn7Js4jpQf6Cg503E0LnHjjq1umOEvdTPlRGf
iDW61rWUSDDCT0dnC+tfCxkUjY3f6ipvdBM1jEV0M1bvko3HiFg7Kxvkthu9Oy2z
5z8QATSEHtfnoonARvqS3z3ZHYMRZ5lMkocNFtxZpumRp1oryCv4w9KMGoLYYiLF
rR9ZCuaIiMnh46DFsRU/ILYmKSqPniCNtlE0aSS4s6vULy7oyeHuBVSjt6PYlmSQ
O8Kkss5PsLNoSp6MRWgAStI2FOfQYQsBoTg0mIcUM7/5GBmO+VPcJh8tnsl/TPxd
GE8UhVUYimDJAO76BbC7SSijOU/vOuZFcsEh8+/KQcPK6lFDMgJvjuXufuvVCJpj
DM1LQCabzjNxvBIHixbsPBMmdiNqOCWqG7cO+E75ucVtUpre14cHMuRIIOaBlNTy
g4H6Fg5eM6ckmU99JgTf0zFGZUa9n2RWZSQ9F/FFdZZl05wkDgN2oZmceALqHQ1T
OCkOhs1uG9v6dNhaThwevBVm/1RTPt+eq0uaKOjJnETjG2q4w3k/X1uDMNlqrJYr
Dy5upNaofqagi6I4bM/AjHyyFS89G1L15oREGlwnOFvwuHdXzV8WXS6/emTd7D1b
GydAeULrbI+MUtq7gVqYuJaXWmlNalm9RKXYjDJ4ZQq6pmZl5UxAaIZbXsAS2rH6
ZIQvLJ16JfynyRosjJ3YCig3IElv+3J6iEDOlCkaiEbwRF1ton6N9BS9H2lM+F0n
o7wf3e9/e2IwGMcZb6qsgOrcdth4+rta/P4l8WVzL/Mrn66ZrWe4tg+ibq64sSFN
tzgp+eUaKNGgBVL2ZzZFkBU67jNNknfQCIpsPTmHL/bKVfEFvWffsXlH7T+un9+c
se8bI/NIVjV85ZJK79ynYHA89sRDtKjVTyxkGrVksxwlmnRGEW4ceFMRvtVdX43a
yMktWNH3oEaTs+DyricufvvuwcWISq9Xbj4PIlyE2E0KJHUgk08GJd2cN1Qhh2e6
ZBtBONS9eu1lHJCvSUZ37Ns3OsG/do06yIiiRViKuVfZso9J96UJiUuVHnh1NKTF
q3kJq2gmcJFqnZDyxyLysOk2w4ojp1pguRazpyB/nUekUDaGryuyJs9CeLoR19tX
4OrD49qk+KHAPax8TJo+p3zNBJPWMw0z9VHHEJUE1+1D9mFGO6uTi3/oHU2zr+AP
oMaanaOaeIkR9FyIlB3R+EAv/sRFoQpDxssyxdPPIusT9xyvDIA0S/jTVBoaIssk
0iBIxUXGuofueNsskdHb1DoVIOC13NpvIMerCfu6+lEgRCR+JiLckCn/PTwAhrVJ
aDmrJxqbxyxQyN3jW8c0/fGym22rzJK45yg2BLTGZHuDpcqub4BchKaKVoVq1JML
wjIBqHYlPDcRijXlPuaT+xlitSN3e40HUooqnRIvlZm5IKz/3vhmWDTkwSI1ICWI
rwNwdfXTUv0s51kbKJB9NJll1CwB29/ulTptkBEPvk5Yzn5iohex8NYMr27hR3p4
wSTubCw9+5x0xZzFf09Iza1/YoWUaxVvbX7mAm9jCwRkjEmCyn/Kc16DaadSzy28
CCESiiKx0foLOUBCVikc3+DdqFDI8oAWEM/Hac/aYKdNbWpnrWBtCBjcjh0GrgXi
f472Kb0tYEobHwu721OZG082Fp6srMqPx/62Ndvl3CKzYztPykjJhYe6n2lslz8k
Wpx9YSXTJ+TsYHpZmhcpeZ0THqr3Gr3p8LZzxeElZb33EKBCl6WrcGQU+FQtEBvJ
KmTId+Zf0RKc9SOuXPEjNysmAdppWUzvsSz4xIMUmjcJvmET58H0/EXeLq+BfUuX
o36RgEL6eRNc7HadeE9HMaHtGtSWalckUQWxdLqiNnUusLm5qMyvhqsBjRXVMCuX
RNVHtshqU1bZHCAlGk9ES28tDqbWW7mt1ZXK+JafViLaaHQwuL2uKP9H3YdSHCd3
scxuUsw/JwFVqmiTA/qRILUM7hB1pkoSx1b3jUZZxzwyp49XnU/B4iFzReTpeMVZ
T3b5kh+wvqMH5wezuaYLhNNvzhImBXVbgrKfZTJypumzSQFSGbqCfPG3WAXavgdL
WQqJB1NBW+4Oq1lcmYqZS0uceDIkauZ02zcm0VQ9xm741D3hAYJCSBm1yBcz/FOS
gX7Co01rSIoixVRU2H693EzMp6+aUKURL3mEhGsAqHyW17jrvB43tbWniPK1am0r
CgOuf5+J7QGP2zDcI6u3rlMAGN9CosyM5OMfRUtSQLcQQ80o1t4g2qEBLIhH3Gtk
+6DWba50kFoQ7mA5AV7wVrWJr68q/bTkiwNmlASPL/2zdTK40P8o18GHA91nXj6N
JPQMw79s4cfHN0GwX+HSvI3skgm2c2YbVskFAC6iZbi4y028cJN7vQlMJIxH5HF3
T1FAV0K77Ej4OXwNlt+qzT8w2mbaKbBfoYJY7lvoQsfRfFP+0dAtz69ImuxICVME
HNo0L3Y4ttSWmcoCKilI1VOW9cTP5+nJjZ68KYLlnJginTTAbp9MhYMP2SUez8Ct
/cH2k5a1Efwl4msJKDMk8hARwSju2U+dNmGWpgCts12TmSx7NUegQnaMlHwOcRg7
fQbbjSft/78f3mawpqlVnJRt+ZDGN6IpMKNYXadgIl9dF3yabr9e8YSVWZhTVWOC
ZlKv2cTcJNGN6AzZJ6OUlyM+7z0GtJmsoJROiIUy3znUHTDcN16mmc4nv7u0uni5
IdQI0/i01usYEToygEE2y1RwSP4PaRK3nv/yeVMIwTh9TpylDQF53apV+M/z47Qz
R1SK2oGTR01cZp20EPM/4D6iep8spbALWtMUzzX8JrLD+6m3OYF88ACFt5xMlp3J
rH6tIC4GTuTT/0VbrQrn82GmpcdVLlTqxnsCsClTAfV5Sdw6IH6v3U+FEKaWPVeV
PFNL9ob+4LIRzR0/23NJBJyQ+2ZKPqIBbHplMHxy+bjbqi9RTvGOIfIjuxHHGuoV
Rj1gdz96KEdwyTNUkhsHIvyuWoQI1z4Ske6cgzOzYeBVRoZel6/xsCbFNfmvTuUA
67FUcK9va6H6b3+DVPyqXse8CP+Q7B17fiDMRuNmWZNiEh5K5GQ2ctQselR5tS42
AfmVlpasD3mAjeBHl+yfG3IYHFxKOaq3HbBTiOXHZAnwGFtAxkJlcrfP+zMbSoYP
LWioJnNrdftXkpIgcH+EfVNsNfZJn2D7/d6V+XRpYYcgRvTF8jXAuY7t40RFsq2x
PEj1s5825vomO7y+r+OxdvXChbAXS5//+KpntmsAop/SuNNOMOKHjI2RVMBCJfrg
mF3cki73l4EouWXZcQX3COz7WPjQ216VK3M/JWE6du77MK5qvg7ehSBwKif4yD2B
3I0h2uQEpcuGCb1X1eW3BqTGvgaSub6XJoNQnYSkwejvtrIN2OSy3vTkZeK0mHaY
gUQO5N5betqlqo7Q6y/m1+SGu92eVcB2MgZEAlL651lwy8Ka+HYKDoPMZXRu+67F
6JR0sFlirWkgqLQx38wby2JwddDydeKQDDfCsQ8QAIXZQsiq2SoiVMmoh8d0IFWx
9eM4D2CCd/289UIU4qZquRXeiA2jTd9OGdWsc8zsmHBYW8vzPO8YUaXG+vQ6Sqos
Iki1shBbjvHfinOpfCKWI+GjLxiIOqG4ZF8NmwdOiqIK1feWRLjnantutcyjNUTJ
wCv2gLwSrYJKGI31gL4NlhvlsyzDt4PJIEoxzF9Z8KZmMO9gk6Rq58aUSIGmB3VJ
X3Zds8Scm9AHptsnsTI5LzmNtxfRe7pzxwln6gT5gaOMvXwZba+VmAvkQ8vJXEVn
EOmhSVkEm79WnxS/b315BDi8H4JSnWMf547Xnk8zMsYmVrv57RPVgOi7stiw4kyZ
tb8cUmZnmyJ7L3bmsSwF0vCOg8qVrLxqDgtOCu5T3pJJnwZgKMbeexaTj20pB2sh
p3Xf3ObNnaaEZ4+ALyL2f8nNF5/Yw31yHtNQlArhAQoJrHYCiNCp0T+r8aadZB6h
xdmawoSv48sc2dgkiRsRBHeErKncHFx75+An2tzrE9MC/9xhMaaajheNmwHuXfSR
oIKqRwoqsyeqd5omzObmDnNMRFBmeKHluQLphbp0cfh+rqoKil9dVPOnhVt03vN7
PGAYtCvd+fEpb0wApG6nLep2T0xv6mmiV7wfkB2PejHjiJZSQ2mu9oAP/2GIZXTI
DRKzlH5BxjerGD29kmiGZ7P9KguQG1lhci6wQzy2/5wsBGE4Anw9y0nnVThUJCIW
36LjcG4ED9iJcfMQOSqYB5G2G/dzRNUBiSD3vHITzoCoJ8Eljm2+VmNLXgWPaVnJ
FcNshfUFKehyvFnFUf3mMwnDrKt16YSXlV6FuMLKmo3uNQQ/69NBg336gJlTvxRL
MRUhs+ByED6h9bLeX5uAxub1fRy2R9QSdSUp+gZk197ikhOwpLvXjXt9KLVZ/GEI
kGhHvExCo83kMc5s6wEpJOjS+pJuzQ0P8qtmC3Kun6zoOAwB2iGstOQGmT7A8T9x
i6AijYiMQ8JDa28eQZiCl1jertgjWteqTJ1iA33H7uWR/xSxlo3vhKT5Pf7FbC7p
Kkjni4Utsvg6atWYQWE45FRQZRAIUUz7MmlWld/nJ6rt4xpBSuRB8Ue1tleyQuz6
zvhr6HTXKWk2G5YtSMXoLCaGYycIPE00koDk3U8iMPUeUz4+9iJq3eeJnbTRvZkC
PcxG0/Rhe2aJtoEUa9AtqcA/vGem7OubrwcKi3k9AkYQLUwEw1/xURFCHmsNtlNi
7sb3mVPWMhcu6t43iHdTxzLro1Lf+HrrY2DT+Jrial5L5tribGvfQZn24hj811qJ
bW04z8l9DL+9R0t1RgEVSbzwous0Hzp78cvpDs32bgtPEt7CyRrGd1E1Ozxc8cEx
5dU2AgD5e0MJMPpEFOBoFu6trQDrLk53ECsJW0+NKTAm+57QkMdvJKZEFxV+Yu1B
RBWuznH57ThfSzlLiMItZKF8HZJaasIfqz5vSx8vya2usp3UlLbGttapwsG0nmTE
7+PsTQQKtvaoJ0b+vaA97jRHNAK8E4Co7GMrP0HvR90S+YdXt6GYoHtlP8wvnU60
xkgGRNWJ0hHhzx1ugxC9qSMshX9tCBLVFYIfzXjdcU7sb/rp21kfMxBrI12jlpti
zVG6x74Id7yTNX6D7xJOrLr79IlX7gw8GTolyTmMhVAULG8MBpFv7VfpGsiNc1y5
DfIkVHr5trqIM177nMMPj9ETavXMfOt/LBqc6wgBnWjQXOLWnYAiOmbAH7PaCRxh
p2P/uW+1gKta4Sz2Oz9iYenIzQNpP8tLSsG04Ej/b63O71P05EM3L+GVieVN4XiE
4pvs8Ogn/nSLauuhX/fHm9Qs4o/p0zGx+a7Bxcrw6r9kUYNlXjdUFP0/xi9ieUV+
fLBizQhDOCxDSRfJHJQdPlVUtKWQvFsBdPwt7B/a3A5WguKHdEGzbsM90+M7hXGw
M7PXb2wQlefedg8yEllf1SWU7xmW0ZD9324xifCisy8zokUGUNkZMxwoSqymEwGO
sazEnwCjWrJ9Wg2aioeWJ/awwXgqQ1zaBKqJYgrI74G51Ff9SQi72XHl71WQS+D/
VY/Mw85zWP0dHyaFkwD6p2mrsW1EuW9ZYXlihBmjfuTK7U/qzB/fPAQsO1mMBwyO
ka7nUGW5BWlQgXefCW1XS75ujEHCj9KJ9NXufduepmMdAJRmuW04bwuqJCHzV2+q
vO3/hMz605Pb2JC1oeLfQHDRQ95+JdVe/6SfmuOi+5MVGhvjIUkVpTggjN3mbHvz
hsuDWkahviDMnJWPYDKxktF4nU516N3jMEna/HNCaObazXsAwsxP73AIRujh0wKF
yfU5nVaWPqn716IBAau5KPEeuNmUWjqxoHJzD1XGz2M1fjkiojo1k53A6p+ZG8zq
3pOL93TiXlcdesddsB4mq5oq8Oo1qsBecadcggymq3BJRaWTf48fDvptZWzpnv2D
fLihY3d5QaU+JDMR6YmVYWb1UVEaaxCwqUGYsz37HYcx4d1DUR6P33jvcv2lAy7Q
mFSyXHZofrO4AXGw0MQcbQ8hleuxVweIaI439+ayMJNi/FdgrMaSGfsJZP8iBp7A
mnF60TK4z/HyqvOdpvMT+KjcCxtfmB6/dLnijUGC5lYTGuyQ2Q26sp3HtMSQO/ig
q/90QnINwny5sNTgwfMGACO2bhihjl/2frZaf4Owwm94qKDg8iaXf5tRWX+jidhg
v79A8j4XyDs0K600coigzJvHwhTXNckuGFiUMD0exh8d/F3n0KPvZScj8SsOlP3s
15shYLqRbZ5XZWMK+GTQT9lLAQN4IdfNT5DOOiIEPeNrbTMglcadivdDUohdpQQJ
dPBMFL+lzRn6i3ytO09zYSW0TgTpcr8R3wLZoaXXVzYOpNA0wP5962WK0QOAxcYh
52XSoJpuYXBT4CzK0RAEuA3aUYZKkMHrk7SfO+mh1uynJDbwjYozYs/21+wfCAWO
0YFcJZz2gFEtO3TYhgBNdoYEuZnpD99uUmL7ofL0/aMkru5N/rfr1djEi5nRbHwb
QJkjpmhDpL6x36SqHsHZKayntDhiefhZDoR6i06HsfAyDVoLbFqio+pBiYYZOUbt
BoFiDARl8iceGf/p8pe1VtfImJybirnW5+apgJAEh8gru5dEQblsF/QP5LOAIOur
srYK+CiKrWasPhxxPBF5KHAhMN/3XmHhXwxhK/oOUlQb63FcQghdg4plTSXI2KaO
WMJz5nSWsmX2VWkArWdSpGfnVDFgG/Hlo1ic4eMlWHmSDvCA7O3LGSur8Bsl8VIi
0hpqran261hx+8uFbGGjVQ4eNBAa/FXFxJcfkPWh2mAwI1Is40NJGr/isBAbyvMv
Lqt2jq/KMTuu+j426D+2EBL4ScuTJHDTOWm6sWzXHqGnhN9NVLORD9iraB7Xwhox
XLV4L/1fIal/3d802AESAOmjWfka48nuKT9wUBtGNaUbWXbjlks6jwK0+ztmtQPJ
ME7ntkCdMsVuwhDuv9xikI8bCUmliuZQiLpuCxbYw2aqIn9kFL5yGeyZqZBk6u6Z
wO1qbk+75Ea2kf+9a8srJRXzOE5ON9sxtqIcUCW1JSU2BQmJ7nQzQrJ/MigusHiM
VpL2Uo/HH7cTKZyHC/1O+GP5VpxJhtwX+SwJhFBO1LjenvkpJwclJOgCoQMQNzY4
W6MU492ie2Zt664maGwgc9fJeePNh6W1a4/rzckjED+ZLh020+3MppytppyW6YJ7
BZj13B2YKDOseYXAbpzv5fNUl7YtDsqQDerbKCaH3ySe8TEW+zdUiFoTHarnBoEe
4KuGfVHfDMvbQNjXJRySuzgi/WIAth2Kek4oj4ZPMVrxzwnx8fNdtnfGoEuaUb4c
lMI4GmClm9nJGPfw46c8qNxBzL+SEG3koDWazJnA9AePRrKU52+8MsjFsqzOQ+o3
WLerdCj6jwMyionLNyxbrJxuasl+8Ise3CXlefgXubkI4STxXkTV2mmAE/CcYefr
Qi2Ymm0GIvcXArKLkGNivSip21/vIY9yTtRYZijb9TFmhsvq6EfO7B2omkjhQBW1
NfsLODDbbuLpOABZhS7ql8RXrKMgi+ylxsJ2015Bp9e1z//DD2R7LkYopT/kZ2Qk
f7CmGRVIlohZIQMXjVz/X5nuaeH2m+ZHTzoNtT/1Tl+pE0YNP+7RaaFFkjh0FLAD
LuES+kHoLWc7AhfQ23svYgsnYVCluMwf7qU7ZgZdZqa3EaRu5qA+tUYomosYEwg6
0eL9Kcs9EI8GDnZEk0qDvzItjDxmNQ4D8NaXBA1DyGOLxA74e97x8JbSsZVF+ZWS
RmUsvAkWzLNXkdiLse82ROqwoL9Xp6d/56p07PGAKAMOZy8/yQ0Fx1ttce6+TmqO
HcX2g6HQtgMLOi2VmbIXcHXkAmaOFx6/ZSZJajmjILZTKUkiibiPVNb31l7WFJ+t
R5YqwAdwJlqzjwY6N4E6/Ferwt13vXVLtSrUKWo1W7VTich5kFDH0RbEMJqix3cQ
SlfkTXOrttEHKGsU+SqLimio8vtN3Y4KSETXbpnGolnhWYXlckNoPI2Ms8Vp0Gv7
cxSmYQPgQAb1/IidcTowsMJHf4WCIL+gfsGFsZJriTta+/aqWXNbZPv5StJvhCYW
wlWUwcMXhB7xvQjPyWNAR/7HIu695bpY/j8TYoP15arXU4n6D1h0JOvT8/ddt2k5
/tfcJlciVorjt2km7ghbIDgssA3Nen4bLaxaxt3Rc7WvsH9B11pYgRdErN5ACSu3
M6ugr+Qn8UdIV9sNW+nbuRarGyTd74i5d9HSRTcsEgg3a6yu6tea7zSbiNpyjt4w
eQ7c1XVgdF16REn/Nwh6okoHmMKBIeYf46S+R/J2YfHvVBrBeVG32ZF19eK4hO1g
peF5d9bKKEa30IcZZ851Dezw0slDO0ie9Iib2yrlmXCNDawNVzJX6g4mrFFoOa+O
NSbt/apdPbwQk68taYRGPMZfeLabPe6fKBClBbwsUj3rIHtp7+mmsFZup4bHxmI4
uCc9wK6yG7NfZI6+7ctrAJgkBNknhMYhQPzyE/F6lKDHKp5qaq1ITLOLCk4kL0al
QG1CmEVJDj8nFwqB32UbF3Uwi0aLmuFut9yUIIEMgj8OOZ32ZmLeYuJCWBCSGD/s
zxPxgFBy/u9Pw1zs1psDfrRUDLs1Ta+cfeJyswk06UifWYNxG7Bsp+moUmuZxTpW
AqRNSFcip9xOBtXPWb2YZEeaBdttFffHWSaGsOBwPnNHZRLMa5xJqSNs45V9HVnk
4hd/LUfKgL7+Vq02+OilNZhqraWX9QMKelMQo0lYYERY4u4tqku1PvnviJu4WCw6
qcBBRAfZBZqxTNfdikJ1i+2mI5e7Pu9Uea9PmTIUcQRpCvUv77c5EhxmgEntLGov
yqRzR22ArbRUReGefeb0xEM7L3dVC6FxUCfX6qbwqBcRkvWXaYQDIE+z2PT50aSC
JHJ1ml1lvAastogoWs6WTwwYXIDw6ywhBJx1LXNmsKHr5ZqYyc938tMWqcwWizwz
CFeSc66YnQtopWfUwkidvnwBKDbPVWW6zTRVFmNe19tb0mCNtfBJh1XFjaD/ceid
Gj8sQmm0UtVmZQxesJ+oqSLZrExUMz+u7q/dhtoUzCHwiefb8BAhrlEATnFXi5Eo
CCJFQXEEIA3dGbScNS7B4JlyAcCZIdUaLj6T9b7B1MYaP4042E+WUxc3qUYg4UCW
r7qgShZ/hBUvfrd5LNf4cnfnt8Ff6IaEuY6nxTupWOgqYy5X+kUE5o6YpDOh5OO8
DzOpcZaJGPYu4paD1as/Wd99AP6cC6y92AlzhXIymo6gceaqClRRlHrerN7x0NKF
l/TyTxdYlKMT94YcFRLn872M+jdjeYbLa6u6RcO1EqdNtUaGnDWUKKaq4uVScLGo
kdEkFIatsBLSk0ejt7DP+ujEejw15XD4BUvtDDou0aiIcJ/xmQ6gbaMVD/6eaTzs
I3PyqOpPEyvrxIvOmHr/7jIgThc4GlEu+yFCBjktMruQN3QHbOm0JnF0XMXQy8Vt
868pkUgaDw+Qdo4gv4uctQvT1OpZhxFtRSSUG7uZMCCcDH73SdyKdD4qd050aJXb
tNAMAZo0oG7bQ/8d/yGwttHn47HTvo29Mx9TUG+KTI3o36Bud7Ukp7hYWO45MI93
5deh2y7Z1302C+23KIHCXnV6nlXXQebg0x1w0HhEr4J2WkeLTxgP8rhJ5WlEJuqJ
+iLzLFzXvqeorlfUWK22wnB2hWQMDh2n9LPP06NnTegU/h9aw5xTTnW1HZ5YYBWW
amjN/hYxv1cscOJKWEeZo+iBFDZvx331oGZ/TS2QOnmPardGyyRZm6vh4KoS/09m
UW4WVlwx3Krp0kLMT2C+Q5/f+ZOSvXy+K4ORQSYleN0hIH71a+pku4qllVtpKUnA
+IzFUZRwBdjaY20ybvkNaRPy+CWXnNHDFwHoPpPEkHJ3eyIK/d0pDdFmcoEJ30Gp
lF2Coe/ejLeeAFWouRVoRqDpNG6Q/2eKJqi7gSfHEqpITsoAyqMQnVnI4D0b9SLl
jiAGyuvVAj4JZCuVFLKyZCwbaU32VhTgjjcB+Z4lPInWszOM7/Gf5TyTyhV96a8P
6f3sYvA/xT6DJ1lODLlmlMCmRAIfQtG8nwbfTov1igbH44VuM5Zqpd+qGF4L+Syi
lDMJcvjI9omhUVJGQ0rlMZANkGUBbuwpx5LR1ZakbaaI9woYwqkRqvzY/JokG+KP
Koea4dS3Rd2PQWsBcXne0/ii9C3u/d3G/xyLRAk0wD3D/8FCYcN21s0C9Axny4Hj
2HkHm/NJGP99PmpilKQBXEG1LN3h/Vh+IirFVN4dO5HAhZkrGpyQ77Qc+cTErOnU
LbBcu+V8M0cHa1BA/skk1+PpYgpoyzNAi9dUmvTWfFNry4/CHu2zsx14YME/rq/F
Z3PhRRk+Ah7pVVd9Zm9hhspZ74LxMI0M1lOwLUBpGiT7kn5MK/vpTKdIrHMoIsH7
HUAgs61JcnI1wdMxYt3FYK8S/u/r4Efh4suQsczA25Wp2oO35pno/L1WKcwBke/s
bCfC3ynKf4rOlRGOCVxnFnGUpj414q0E3gB+WjmXJfs1TUJFJnj7XB7d4KeKGkg/
INMmyMlLW+9iHcHmNXyp3TeuVb4tP+dFRt7UYPVIu2/OTzlr1ehA2RzUCQGoNpdC
996/OFFDINx83X0rhKZTHbnkQyEo8rQkIaWxdufb/3EZ4cY3LQmYoh6uGv4urr1h
Q3hN5nRgACB2pjReDiZ+BVqnt3EGHEe/AvbNBpa0mlYVVwg2b9TzYiz2R9XrEkZ9
zDOOfyzUu9bdZnziS/WKbBcsIuP1BOuTNXX4w7lQxV++dgRdaIKom32yGvHAAIYt
SDaNpusT2wl+gCcAsLV6qnGFde0Dut2MRrajFwrNoZFJ2Uz8UthSUH/s46deBU+s
hU1GEBpElBc8WHaW3Q3bvO5y6unF8r7mQ4jP/UmbOhwYd/kcJGhuoOhVSTh9icMJ
ngknbYZXm+YGhYFCcD/QlxEvsn+ADh6l1tkXvLu8UD8P7/mMxqAFdRSsrKLMHoXD
e46CIzzpnAOdQcPd31ZeLpK6PXRBNi5x0qtaLYZP5W9QaECaXtzs5cBbeH4ag13T
WRhuhxGQ2m+4/SbbV0hpu54ZFIvhvZbEpmG9ouTlADxdvKNXd6SzOyHp1PWA9ESj
bj3A2iUndQ1jLT0h82wz5CfsYDxm6VUfzlf86vCD0OuSEY+30DbIcAiRjcXfpNTB
QiFblivYq6NRvXWsrey6MJyEL8RQNU4i0fGmBrwNmlpV7l+x3/XRY317VNsIxzaZ
fR8uUV9bZASFWALYfWRIktab0et4p8ISR0PGbi+KmGrNmeXBp667vx7RjEBtGNoj
5G80GV5tEN+fE0dCJjPeuH6g3+4nEI6euO0BldGFKrBnIq0JgYzqzbRNbLNPQImH
6KUgz46GTJIRvUrPitTqaQZTV9B67uvibGUQGNLoCc3dWhxY7aE1vZMXqfpKsUrI
WiM0kPxNKcgiA3CZ5/i2TE8fc6hnFI4nfI+x6fTAcAMziYPhgggpwHO5JONTbg3g
J82FW8jqEC0vwxONfhbeMuBMs/hUDVTrN2bfbZM07Wkle5OPotkDeDr5dYcsTg4n
xeVRAczhIy780ib3rdCnaB3Igyyhf1ccbfjBBO6IkK4T8hDkIhGQdeyTLa3KwnOo
aVIKcrxacCSlZPbREhtRa9F+2Bj28VEfjjAue1SieNKr7KXeYXHyX5bgijLjaCwF
IFhRh0y2KTQ6EhwjuaunwNPdGFy8mXR00rQlooL57wKlcVydrQzhYpR75FFFFV7W
E64tifEoHDAhuz4mnHNbAh2FpBeZW+CeWiovVeQvGCaKB5N49Z/F0k9PVlE5O9GB
kppTM83gmALRyRoXyQc7Y4UT9ESPCJtklaYR16cexfi0UfopeTXbS+ReRhDJEUbq
XSFBCbyZ8hvbo6MK9LnpHAw/NZLnCk5PP7pLuolz/P4dvRSaad0B6NN4Vxi46nnm
SAuQ4HnO2RoUYV7mDwaHBjVoKmw32NmQTH1yYRSiK/VPsrBOIPSYMr+/YekvgFMB
zFo5q7op/9KsS7aaPymHpgO8ea3gJCPwI1XOPproqD2gTzyVjomzV4OwHsicXm66
x1YDlAWsd2WuUJU//8Cq0iZkYGnO+Q2PnPm94cUGy05fbaz8QXpCxW9fBxbrZNMg
rLixnm11CWhmCUsZ00tVAIYTYZ9wbZAYUfuWH0xGwOkeTGrLnqk3KbKeH4hVJjpF
OumUD32Fslz3FCbgdd5aSjksORTw82GQUtkgSIazuadBbPT5kPbz0EDgWhIMPsbL
nm2QMDwE3B4U70giLBYHP7+WozcLJdedwZQqKVkyJVt9RCSEIbqlvoDVbgpenJJu
GpgnwtYKhiNMEgmhoymq1MRF0ahN2Ydf5/IQhiUDvjufHKBPXDzmT06hx9yZDBvY
1m3uyCf+30LnjtEXKwZbc8nkUSWTPsjk8v4bGnKDBXO540WO2pOZIDUHVAbEFfCW
/HMzqbv1wZVU06YuKLuNHIvYjNAbgRrUTjWo12RGKaQj236+RsMQOe0+zRyJjaql
qFJfvephXdUl5bkHoAkANmpy2psWqu+cDL7ojqTaj+37RygCIZU/WHfp59HQ1y8Q
5LcWWtnP1mZ2qM1ZiD6g0/FKyVtS5HDGRvQnH8mqg6Fwjr52RE2UwtGNyb1BqGJg
GZ+7u8K5chky4DQ1Hkr0HNI4e0gw86XpcyGTLIJz3J3AQ403f41HilnNVKaDZ3wG
IGbgmWno+kjzx3WAI0uR48qWsgBJNghhzQCE6JL/fh5ubqD0qeXLZrvn39ohYQJ+
v/7N6mvyWVTlniRoQPPomhVDLMp4t4fdUF8KhrZh6Wvootq5XwoHf9DNUMZ6MyR4
T7WQ+XbRBe6mMkw2c1tsm5G+tEcjLxxkKrg6+T2358zLUR/XQuBSMB7NW4VMC/n2
Q8jRvWvKp/rmmqscSZ2u4QVnaLQ0F5YQbDydhKmVMuNoDkuZQRMJiTWHxll3C5jN
W7rbZEtLcwoNDlNDAUZLGuqxF26VzqvRq5n7w+ZCxP3lqtsrdqZ2+tLnzLoAyRlF
/6sleTea/fsFMUYvlQ5VqClj9TSRVwr7Zs9+O0xOMEZlCV7vcYm7+/D9BFxEuliY
rVyWSAcjiPWdLofnhGv5DVGu89NXWWUjhuDmWFPik9TI6TEQD/54fHRE63HzgzwN
mowV1hjX6zfJ+47l1KijZhYrvJZHQh6/mSIC4VLlnVChANBadeRpzxnbli0eOGrU
FiGTvE1iDgfXvlKyd5Qlwjx8Is9f7McLpmDLGg2tjr9SPJNt2bASx/ofMVDn/hLO
86Rcj2ZR3bBr3d9TQjL3Vtwmi5NjgUTj9pgqyoaivt3PR1Z4+OHjMwBouiKewopa
to3FFcHu3enN9Eo6M07ltsvLtVXK1xOB2sSKISbX/9TrXfK3ED0ORWjshH5/cT9w
Eb79dvnca/2jM5l78CabMu2EKT4Egr2T372QFgSLn/oPqxedE3rMSPh1+7pNQtBA
HNwlWXt8fosk5Ud/Qn/ykBqgWuuCf/O3FP5ngfED6ZvGiJoZ7x9ReBV3E7w0G35y
Ym2ojKKa2EC7RJ1ss4jptOqnnwhYI5QHb2+dH1UpJQHsn0gTsAHoPOMas81m/hsf
eP3GkHGhESKxH0qaYdG5xyZ6lSkGyPQBPPjhooRJdHBnTxY+Ws8hcuxAaQqu/svL
0z5JufDXg8QLoFDMO3ZJoAuxPhf1Nx+mv9PW0lA4ptctPMDT3E/dpy0XaGZMcGpZ
3ljL0j7ydh8nmh5xsuxhtW/mAayQlQ02R6JuGJ9MZd02bC5NbErADPCbbdIzdrdl
UKaJj99GY7Utpy5ymnhAoWzdQcdCQf6bRl1FpVQV+/Zpm+JdmwoChdCNO6QuxOx1
uH0Vs7n4JXwKmdGbnt3sjpH66Ta2Y/VeAg/Ra58GjUKz2ZP7qoKAoHS+lZRRHOvK
QjrKaLyttAidSKoj64t5WXyjnH5Ethk6I207xIBQ0ZCTSdDr7VB2UWOf2HkOwuil
aqQpVtA+Ux5cw8+O56MCaOI9gQvcZZAq+Lcpy1Bx560IpcufzYTGvAdhnH3T6K/F
eibb3tsaSZ+Z+PP3WZ2xktNmptT7PwOPw8dAMYUjRHcxfhRCnV+mvIu16bfPIkEU
oL7c3J8wv1oIoSlACNthp8erdEn6bmpcSj5HryVLSEKEUYpCJkzAl8+JoQOdFYMC
aZD0dwXdFPRF9xzNDksGUl7fKt6Wl3Z7wFQ0GEmN7GYJE4JmLxgVckIh+ygEEMV7
GJBakzZeJLg+Fxu6DjF5P2HNEqnXp0ooHa0WxDHMnNZh1FWlReZuje67FdBQD8eF
Ou7z8YoOpeBKZn5+quiH/JeyLW2q/rNor179qnQlq0UcCT9/6pRGALMxsLLdt3L8
1rVVFSfRpl8SszahIyejVVqQVLm6A0NFRL2RUmGhlpdSPo9UMcN5KNIyF/Q+L28O
SEaUS9ZK1vw8tRzGFRinzGHkZGRLpAdGE+TcCXdZ7wJv+GBBqSr8mBYJx5XEz2pH
b4XJiFNBFFEokVD3xVRFLziaVX1rGv1/RyFHH0Swv5zLzSrsAi1dBXYfXlLh24h+
+5oOYbOe9eSLumB+ePO6qDi6UnO4O+a63yoA1KW/Lq/s1foHSGNHH99FJQtam5lz
PqE9B9xo+fokH0vgvBhrfgUyEFxvf4YYTvqVCNp7/Q3jEIOn57QH5r+UuKODXlU+
ItIG+PYggo9fDZWgB2FoQDBrmPTKGRtdpH/N4d5zo3x1ajP/ldeijfsWLV6hC3We
MwH6EifxwORO/4ruRa5nzHX5sbSxuSD40vJ4Z3+M10R9fllotpkFZcYC74ynFQoK
bCZFjhpWAhdzja6us6w3EpkOIFk6Ke1Tf9Ne/tA1nOMLcG5qGo3ZRWY3MFxliRd8
b0PnF7Zwu1jnqfOU4AWD9VeC7PUIvGgfK7m5usWj3XvFcYT2CTCk4P0gViupKiGf
IxmWs9UO97iD0VUrHW8iz8Bsxh53NOIdwCqN0E2c3ELrx3MQfGa00KKG8eq3Z/YM
oZzy8A1uTjBcVhP1lwqccsEmLhq9re46ViDqnzsn01Q3LL6UZFSdEBy95ZEE7nGH
VU014FPtPzoYuUqMRQ0SBxLZebZ0G5xxy4YZ+nBc4Y4iXmjgJ38o0/YyPPnOLg1L
JAH5q54JkS+//FrphKJM57Viv/v8dsoW0NYtVX1ddddGOHC/uzHa9NMl8dwMb3gz
bbVDR0jSsS7eoS3Ba52ZuWGtzFot14MG8og7U7pgAQe0W21t/lKBe4UTjBCrzKj1
8Dv+cvXr899lof/nV3+Za5/K6O+pqT7GtXIb05w/S2PM85Dw/FHUcCWbXja+69Nv
fOxAwK0T6fyLx+Y2rLvpJHvyFHzhwc+4xABY0eqy7yfGv9Z5OCD8TfXJ3cZcvHlk
CY8hUWw07ozc5RCfZSP9OJtcn9gLtTPRVqQ6eSn+htk98q3aNSzkRQBaxwMEGJRJ
1/DSoH/d4ulvMhOZwwEppJqrE8MRlgw6b0e4CsG41tX4keYtNiZxiOgVQMSMDmp7
LXL8B9TlKr+Y9vwz+rg/iwarXtW7XL3A32zikgVWrIfRG+5YPjG1CkH/Ffz3GqOb
PcF32orErF7hU9XoQcW4Dre++BYqjo9HrA9PBE7Hem/SxZyIGxYlAcBE2e5rYNHt
6tj0mcgZfXB32UOsibclacbR8oumcH5MMaO6RNX6W2Sr/EAUYwEUzwtO9k7naWPY
I+ZN/VBBcaWkT9nC3wPoy90jRZYCZfZTSl9N6Z7sNgK2zGzaTWOiiJT8F+maeLZE
ImfZ+E7JVL3RrvoUoWtCYAaN/HVbgaDTJXv/2l36HWVTQASTqTOu4EoSMSsmkkfv
uIkkHHvSd7Oj9usy4wU1oxI/3DYwbUTJKN3xzzVbrYp8E9sZNL7QOA3d+Kg/bMNp
SCFdnsoNeJGqaK1Tgd84toioNCqCQZ4v0ck4i1omC5SauopXBvjVt9j+wFDggNkp
TBC24ywkFKEksYcJkR5/gCqwARAv54aBxOxOxTJShr/j0k5kyucNLd605PBghQqe
gLSLMpQnNefcdm8sekfekNXiRUHQdhlKNBdkcwhaxN5BDlF9mwziygEdqtRfTx2n
qu/OnJZwin2Vm1tO5pr+M45Tzt/zb2m6/n+MjFyhUCD+D+e2AF6cBqJYNFVskZkA
jRojuJhZZUgH1H4PdQDN5FLSrOwXFOVLK8Ff6lCCFf08hxxRQu4L3JevoYBTZsYm
NckM1Yc8UdlT2iN7IBxJemPhxoDd2AiPhOr54Rhlf0rfyx4qzvD/0i2Uoyt7u9kb
IrGdFZhefBNl/J8k7bkzxlN9O2IhLxOM1sZBCwCgLtjWmZCvuFfFTJVWD9x05qiw
+IQosnbL70VOmkf+DTa2Chd3FZFENfyRyWezpTDh8jc92bYwnCwb4tcdLYbY+ZcE
nxLzoNJKIGQDMgdkhM/i+EX6aDuLBP77RuSmsKaxzxQoV/kh8ipwllrbJd/uoiOj
ksPV6fcrNydrWe4GGNsYk9On/+nw48twwzaUsrH4OO6N5WYmC+2qladoKzNOB98C
ueiMwLgiCGvyq5rn1PMmLqUzaeMgWZ2mUlhEjTWQJAIuHFDwOdO3y0TqEkCsC9EE
GbURyIKkG7XSrO/gqlN6GHINo6gI1+SXeGhRtS5JrnksYkP3CweOc6CnQ0rNXRI2
R/K8IYv9K82CdoTuoGH0jGVhKsymhZ+bR3Kx8u2BDKMk3Eb3+TR8F0JUb7hrS+N1
fk3gbelDJv2niavPa15H4ZkGjhW4Z499IThwK5lSztBH8FI5JFeBfevA8as4CkgE
q9dsK18xjXjxX+gYHAXQDeRMgPPxFEwx3VWz+K5D0ANaIooQSK8N3eJCsdLzosw8
utr6Rck23lRWgXKEFFttxRkM6umUP1xO3tTAdeK3d2sDK2uX3W3jTLmIroWoEDdH
5Nj3AbRXKjvLySl+NXEzIrqIT8ud3uI7zNt017GaPWL+1NN0SAyh6ryjIIHLMjM3
3s801FQ9DNvjhhFmyc4s/l1vKSpj4hIkxObKyOLmq6PQF5CSmqMJTleue/yfzsKp
xo2aK35T4CFXQ01vW3hQ3Miql/M1UqadfzbN4N3ZZzFCZCv9GSe5qMQLng0VmnCy
5pYg/SgW+EqG58d3hoICUL+9qU+9yyDtz4abNPPxucXNQE2d50d8xtOpDEAObaGS
0pGlA3EIq9VkDqDujqmIELOCiaNw9j23TXyunIjTR6hECMhJ+gRoGMwCqI/SwVjN
PbFJan7DfeAOvpm3FmtmYHF2nrxq8FBFFNmoovvrZ9AWVF9+LZ2ye4xSWpeb+P+u
QEG2x3LDHsHahL31Vt8fyGRaxuvs4hPmGJabwNsJTyXRK+IanWXCPM+kaVRXU8PP
eCGj19mCou0+y6WlCeu7yQoEnGMKuyPftzSNAxTfJqfpL0p9sGYU/qjwnHPsFLhU
SyRCVpMFZjeVmV6a1Aflkd3p74cvK2XXn/egelQ0waDAH1U5yYkHPsvOvootOfnh
rJcZ32zKfYWtVKAjtwfnGFo58b+XO2gFGSDpHxrsiasUDQiVf01Pf8ZBLSs+7RAR
RIVt9/FnbLVKlUFSZcgywSzdznp31h9J1vyrGl6UfDwIucXGEWEWD19i8xwtzlz5
6jAuNOsxV3VYFlaKoBxboHRkP7ZoVBIqoXSzfMgjTCE+YeeqZ5qj756yTUNl0mE0
buT8fh0VZHDxAE2yQ32Tn8nGpYSuQfHkUqpI3Sfp4x8zgzNgzL/AxVD71MLPfMM1
eYYduXrfSp8Il6G5eBd379bUGnqDWEMcS1ACXft1oJb2LrQhugT9g6RfRCjh2cmj
eTSeawNtcb8bu5ltDnSeZErp/45+9Qo6z19WAZUCY5y/UkZfhXDA68cPSlic6Ji0
vfbYHV65rd20y+uFNSwUkqfTJ9JwkV+tiftj6hXpJLhmZFOEMGXvaiS6dJQ7beLK
JXgxW3elAx9/H2XTG+dzsL+hY5DM12QYMIUfhQC6XLvhTCorIeHWeraV2uQqeq6T
9WL2pzaPq5wG4Jovmx/K62GOINWBpvTNprByZXYRFM8sqoxUIMXNvhMNCmGQOhZe
V8MZCO7l7JTc1pg7hOB3ftvcQPzJp+kKHeN01DTdQHyihhMucHimN03x0Y/qfEum
ZarHzUx+Qa7EOSBUGooFrF8QPQeatmvuYEVnaMaacJD5nFe7zktRxE1sm6iqCw2h
o+o+VqAlNySgl3NFcgCRuBAz3X9I/gzwQW0J0xZnxxOLfIcRgLF3toGtkE0oyZVK
egBJLBtDGjFeE8VQ2d1BqXpL1kqVZskgLS2mbbGOgLQC9pLEwaBHS0dPIRbxQrpb
z7fA0cB9Wk/n5WZqagD6KpbJiiYnSLKK0zaaTJGPpKsP7fl6FCyc6Yl5Kc/auG+5
dT3SkyP1SvxLR35epZxaKjH4br64ChOh+OQp4nshrqA++e42K/8L3bLWRJSOgf3P
qG7WyIH1XXGTsTblfXYoOLrJEheuW1VuDItcDHcVY0p50AXo2Eymf2s0D+nwdeum
G81KhuA17bVwT6rgpRvAFjBfCQqAQJ62sIPCPqntemFs5UHUVT8VCpaseiLabqvf
2942qJxVtu+vy/PmuUccBh0KwYguxbipJB4QcwH/m2Tdjwwz/rOnQyBm2b/Y/dBP
Nga4LHjPp+SULJ2Pb+zq9n26r5RuPuQogQa46usLzy5injxwK6oGbBLbBEmytPkL
I8IaqECz/Sr0OI/u6rkM3Luq8sDBwJ0Of7iJTdTyoGDa0MSH6BQOlQCRwDr4I5rn
+3r14s4uDOST+p8GnsvqSLC3YEuaZWNEmoPmB7BZ7hLwnQ8tTT7e4SPTwVCMwgVV
2igoX6447mW7X3blcyICTVhaYUcQRsrJzhk0Sh/593U2LrSwfnlFEDKCES1gfWvE
HlMAexyUFhVzUrRMPIyseXVr/ZfaaherujDbpDz15JP6qpKjxRxuGzWPhO62AARZ
8dry5jWc3y4fOAyxPEFE4Un7PdrZ8DECPH7tny/aw5OrivuhQ5xIxkSmZJvcOiDG
WIZZbklZNHpug1z2ZQOSdMZU6ilywUwDNWdJjWh+OTSWpoV6/V0lGFYAZiUbW7M9
FtfYc8svkXKKhYQeuXSlwZf0ZcSoekTY8gqOLHeXx3bA52buW29KVbrg0M+lmQ2X
HLBfr1s8nOSRZ16U/MJfBEfjMrA1X8O3pT2KMjUtF/0hihy3naaw4mc2Nntjqy/2
mWcncZhLz5T+UHukypwFw69j5oZ3Wtl+3C81Iz95k0ojo67I9iJgaWUMBOqvCGkD
VvYa2eQMN0PSKJOWr4wLYyEwZU/4mNGffZ/qQdxzS7hnMIqtXpfhEGMTZRbNQShX
l3J5KO0BMdSgp2qr0aALkXKFg73JmpUT7GtP4+AJwfcL/UCzYRMrNi5I3Thy5Cqe
pUQkEYg2AqDYH8tlDBNKpRVf2oRRGz0SukYDAQo2gxqvtuQzXgFMGBi5qiQn19+g
FTal+9GKgFYo+UZLxPI+6Nf1Sg532ebn+VS9f5RYjPfVEZa9/RjYZtmWmhTRr2PC
c99CSj3EyItT5tdExPbMSbdNkmEUMMvWIygUXgQGpun1llgTdv5zjMs/UP07ASut
mPV1TNXfIJ22nIKLh3LPT69Ufz4BivGEL+An1njVcb/lW8VfwbxFkQOYctiubYQn
mZx5ly9BDRBx2EDFMBcPvofT/EV7QiE+uJYmiiuofCO1J2QtJB7FmFu37HXWB+nD
lEtJOW+mIlAvp/WzIGhbeoqjfzigPpBpBJhE05W1lOkYNdi+zooXjT3iImCFYVpE
rMGdpdhPa68bE9Nk/Ano1h0YH2fsSdbmEO0OBzhKjoyhhJTteuKruIplOc2AOttR
tREqgIXFULOZfJXFFGh3cXVGhMo+b1Ccu9WLxS6qGPCPOTfyTZAvt2vUrhLyhIPy
5jm6rG6i/ct1Q+OknxMA98SDSV0C+y6a3VI1ER7lk7Pg5daLxPaqM21Q0A4awwtb
SMZFqaH2WR3OSH40X4Cgs/E7bbOEJU9IXn3KKjJDeL05r62jKaowPjS2XUM2kwvy
ufb0a8SKHDRbOjW3Tfr/hRHagIxxlvbSK1Iyy7+kW0BEpsnSSKkErM9J6r0IG+Lk
hl7csF72Z0YbIooOw3lHL5ANywkNjSNDp2HsIGPhj6mJ4Nop6XbcJz0nnxp6/3u1
uSudOThlpNgz3jDXmW/HGVyjeq4Rfv/xqI1vbPH4XAy49A8SsC/kfV7JtAnaqeVb
Ybm+hnBEu0wVVnn2OtR/08hhFau110KfB4ONTcj6O+MZ53vye/ijbhS8jDNeTNA0
zrfD0wFUhV4p9hZleguS5p6f8BcghGdZdxPKqmYE723XLO1tXFfFvt3lBPnQ0KCm
bC7GtS/X5bCTMsrWjpDC3JjdCrFvWGZ5u9VxokcLPORVSx74MU23E6e9JS7Lh487
zuv8/QHhGe85xKQkZbg9QcG67K/wEWUswiReI9duSIRjsF0L7hvtiDw5Q4zs3AMe
OHZhaf5jBt+pODRpTwQB1tIiYN7JdUC7SOH8lXVDWpGgtrpEFqliDtCQlbO3pby+
KnHvA5wmX8yPWhl68bCklc7G5XqkjHwBllQ26MeVMznq8TV0j2vl+u31h0T0lr/k
nF44NqxyffK+sT6Xcm7pyiRb8HLOFpxzF058lRl3MHcbGRpnp6nP/yIj5rSJrKDJ
q6UTOIvSJBeDfJ3mCCp13L806OSeeiYXP4cPADcSJNOMJY3J8vpqJfcG9GfMzq7D
g10aRJw80atIuodH8e+EJHmcGAt3ird6iJCRgWJyHdbEDY1UCHhmBPxWDoQph5RV
oKr5Dgv+BG1o62hbb4SBS4DCxPtXBz3G1W3O6zBSmQnQmMhLxTkCy1qojaO1ORTX
ilAqimgBxSOe1O3CmNtQXam7q+4TZk6pcnIKKimsY3lzbGDQQk/xvxa9ZyFOk/Cb
LEq3dTsolq/BxFa3wNVKS+1jkFe+f1XjY/OhTUhZ1zvA8S2a2m/LExkUYvypcbpB
tl46kpDv1J9UaqwBbXSs9ZmPBO2brLAPibgBOxgeV0l2gAS5hIIHKASDze7n3Jl3
qQ+58xUxWiMAZ7D2DaTVScntcYnBQMMKSK7WTExD48Gk30iJDkUvkxcEFD8trc4N
VycmgM1VNngKmsaan6KYOsGnhXfIrVXamOgdbKi7m/uDbhDKDpy193mmJN3c0/et
LpAB7L1TRNACv7/kekKJdIDxc4v6kt1LcyLV+CgeThWCk48BUMvkU5Ju4Xz1lPxL
W5+jFDFWly/hhA9njIFrQGwh2LWW6fGRyrd+u3EqhoBJmrAbNplffpMSnc6K/+9w
nXezafDdil8nDwcVpM6WUHBH35HhD7YaKBKf4ls0X/dtlxoxn3c1bgWi2w/hP7oh
gaHyaxGaRot8P0V9XZU7FkUj/4ObR/aQYo5+n/BbTvSyjdv6HwwyyRLFDh9YVt4V
B0jnEDxvi7wpGnhmD/dxF2borG7vjQ6RyBw94E7MttnoyUGb4+OOQ505z7RpheJc
DZTvNGOzjf6XzXz/xEAhwNoUnn620quf170W3dik7zN6MmGtdlcto2ugVa6PXshX
XzcZ68f2VAIiq79LCh4mtGwEai013c8j5yzuFnZ9Tj/DvNF6srcjUCDiYG56fdn2
xEB/so3PzdycSrvrbu85+YjYjc7BYmnx9s6ekEhCFcmTYzIfO4bye8Kea1KUJSGn
D7d358yo+26zLg0ykxse7Rl6DSmxWq0j3d+ms115ghq16kwm1Ww55tF4bheaDrUA
AnKW2ChJBXkiESEf0wBIcAVxOFXH7iPa5EedrNNsmIMLJ31vePHIL77yH7lgltcH
+nvX7UD18DE7lHy1YF82cSMzt0yKYKsY2GxprRe3Fi+Eepnd8f7AZMR/J4uXreXx
PiqwOLUNOHT1KwXovN0ZHj+nFsmRjl15Ea8fR/znddrIaw7mabyJskWV5AHwCtCJ
lC6Y0xio/ByBFCLW2HXY2QL9syNJlmaylmS1Kao6GJvH6Vkufh3HpEWyDlPGO3Um
JnlEvBzqTW3Sh57w6PYgMWQwMAfVrZZyn4GWX2w70LtB+U4rRoU2TaM94PPSaAof
zWthdoPcdmtTkhwjZT5TMZjKuz3JTGbNoypvBQz9Yt3OFyWlcDNbbyXNDpq6wtP7
sqb+F/XSg9X/+K+JP3Azb9m7rMpEf8d2uE4EqN76e87DrVIYtgpexqb7NV/fzWDW
CR44iRRmEGgtq+GOVYlWnhKuwvnWeR5FyXn4PtWFW6cxXM2RmK6Zgu9lDkM1TgJi
jN7W9XBoHpJKGfjV9TfUawKmrLMxLWzrDUglCaGwzy+x3QNcIpoI9aY2mzslKbdD
sdXIztnssvxe7xwk9KEbChk/nmEIxWj6sv7BEpk6s4N9b87RMnPJ1uZQDJH3TNv6
90djlEcgvZ3Pd1QGQ4GHE0hE7C0Ocpug3EsUe07JpT8Lu9tWjOhZNOblFLlynCwr
esy/2kmI0clob20ySLXfLH4Lem5hR7YaaJMMzyrEWeBU0/wLUYdcc0lf7ug71Q7P
13tK2ewcJhhhVg/9cmAjf9FJEinvjbcjt1CMZTBk9Yn8o5xTUXJEjCze++riTliX
SQ86G/efnmSLy6hISIDFxtcStzmRjlOtGrPff/A+LAuT59MHXKYxcH8JbpahZP8V
VM/PsH5SvwqtRH+RC6TLa8guCpU/YuhlEveCP6bdRUeiS+DGEP2MoUuIp/0YHUtk
IdsR9tIazxjAeSRxtwnMhq4N8U3gIlGDVZ7FIHQQOUh86bIMxwGyZVtJ7yguaRsA
x5CKxgcYuo4NLBQ7oOTNhfaBpkCMLNOUCguvsOuEMBZZN3JYdo4RAgLXBj3Is5HM
NbxmEKTh8X5mxd49MY8fi8VCs2GJ9Jlpmj+RNyZs8nhW4FgVZEwb9l3CYMdX4p5k
F982OB6ZxMQ0s74VD8G1yxVha+kuJJ4pODzXvxb+rjRtCQtbl3qFG8KVG5GHfxwr
8WjtC+hZBGBhmv0gpDAUIhew+JaOayR8sn9PCsZQnJnTYPSUKPF6iayO8EDuqAzY
vYz4GidbDrb6+aHbFvAqN1kUsiISnEMde74yGnkV3Kd/zPZcmOz/n/K7DqH4Vf0k
ZOu0LgxcZZZ6lRaICtPV8VOfiWiSwRihpYxOmZJqSeaS4asQDGAVhYaNqqbwKPpq
XHmAdj5PA/UxX74LouEAPzt28/H3T2Xp/6xFW6Rbzr7pUrAGH46XgfJuvGZF94Q8
o1Dwa2xls9jTgPF0GCHrgaLvJcZZjkkp94a/cZb+s9jSXisXsH81+Zk9tHwYRnFx
AxX7z6OL2iR8XEhDDr9L9D53zbBdAm2kyGU2FhoW+N+RMtbyLOuGQCJO9f8TnazG
yLZ650JS9e3UmbxzD31oOYeNOW5A9HNXWWVROpHGECuT9+ksT2laO6PsZ4rQ5fNm
AKt1qE3vQPmYVZj/ndwIVRuHevUXghV5TurECnhRY9YWJ+kEAJf2sQynl+PVaqSu
RwR5Gfg7pIfv+i0AjV99GpRjHospWWpxEpZvA14IlZI0/yx6onQGKKbUQAMuaw+X
nJ96dij6ks8f+/IvU8mUjXJo/rKyc/dORd+Sx8vKv7xjw9w2jY5XjPOQVZe0/7gD
aWAMQSou0Fg3+h1DSycH6vo5M0iBOnQbcyXNbCJprbzW6f1lobEZkRx55buTV/Ax
e/Cgz/3fpcsRsdQHXetdriOr/w0MsqBVjBKtRFwkdeRdBmpQZTMP1Tu9tEZ5ttRe
whqwnGF2ykuIXuQHPrl3oRzwzUDq1q7GADKxkQ/U6eF3UPE3LlKEpfsJxERXdGHQ
b+mXT8qmNOj8h+D1AfgK4WlaOW280MIxGEaGEKR7wfRKmqEKZavu7b5zAwz4K8XH
VPVizSApTlevvNO+qP8Jh1pQ6CgQJi4/ZVPxLhH0vaIDuH18BkrNjvkpDVC9uFrN
f6JYyOOJTnTgdZaxE3fQp9EmUVL8jZuDFaBC+i9Q5XPXvueVtwl0xfqWgvB1gtHm
a7LJJdVE6/1cBRS5JKu6vVWAQp0KduyFT9wEKd+kst0y4u8kqU/uWdgWwtvytHFG
L58ZoSXTyp2iKSSHmllaAsU5Kp2QCifbqM1HiSvAvCDVE/qbXD1t1r//31JAOgds
j+f59o8Rbpvec3R0cwpHsibj9f3KhbHnwvNX9XuU7sH11ns2RI3DZS+Cj9OQOJNc
mZVSiP4sl+qfWZz1iUXx5VAV2FUOJqF4EvmaiTrTfoiaca459ZUp0KJVqGXZJJrw
zyh77bPD3sOfYCnFeah7Fpi+Q5JPAt+dynmGHplfqvNMFtO3AIKYFCLPTIf07BK0
4IvfWUFN4Y1Q4cbcbdrJ5QWAscj5XtKKLGGiwBdsyG66xYZreUnGJCFOiFaduqCL
b3B3ZrHKpuk7YZJeHAPdgsgJuWoWPI0XQanjsZs3NWJSwqOtPXN6i+RsBHj2VW8+
2+EDMoeGakA9w4qFPpNvtWCLd/pO562zAQcNFyjIjfg14HuidPiybC7cWHj1kkxf
rKjevF1xft6VL1+8BI1+WJbn/dEQIwzmjF1Iw++BAWaqTdyqrNw9XaF9KZbL1YTA
/sXMDPvEbkxaMY/FG8goRSvAnrOc90/fvf7ubr5Drb8E0r//EJDCrMwEUWOnVc4E
vC8fiax+ejkvgQg3GGNZL4iXeoFJnXXtglogUfdyqReEkbk/NpksvAcaoWaNbrIO
04futDGohdYQOHjNV/btSu+l+BZ7YnWHrSB8ykzzJGMwHzXkgmQ+9k+FlL5rycp8
GeBA6An/V0h1rwJJw4vvj3esHrtjbvIOLSOOuIGP+Yw7ySpTAzZ+wQeXnmVKuUkp
iQ+oo/5vOY+LdhwRcT8JEyl83qISsB/jQH9UV/CGP44k5jAZurwsE8HhqWjjT/hC
bAeo4llk6BcCnHExMRG75lhAYiVi4+fJcaZr67pMpApuad2lA5TXjDfLiYnJOp/C
+FRdT9s9VqI/IoarUT149JeaNHaSoQ2vtXs8NZ6rFrVPfuYQUOHJUoxRz0LY248J
R8cDdy9aRH1iRwrycdLYN7nWTk2fqCHd8aWa8516UuKG26kL9d3B0zHbEcB93oBR
cJAvvin67YKORq++hDtP5q3ZhATYujd20NbQHbfODimE6gOrRDLxKRxbNI6eeWyo
X7Mcfuhfn/C6TKemOSbyvwclfaL6wxirgsJyEGHDzRr4iYUKhqIriAX+AjG9ckgD
hg6FNllQTOTL/U4oFwB7sgu4E9SsfSMEYt3kE69THBD5+Ye+EPknoX/LK5wiEvYR
qmOPDa/r4wFgBv5l0tTm+08ikr8mD8IXhJP9pg+/hYj0uJEbuC3OeU6/LctsBXh0
rVJhvn/JEL7O5p/gK9vbrvT28JGjkEN83avO7eBx0J/6kh01QORLEMHq9CAi2w1L
EG3U0/EeM6gPT4+Guy76Tca0WnoPxCAiFsSYqOVlJKkt8Ayh/t00Q8t3g1GM2r2l
ZRJ6m50mvNwqC6oiXIEgooAJfbxSe3faGP/8QyK7GW5hok9E9T10iHKoN/vVMzOB
H2C9CAHrg42kIoVfzOqb9L0q9JdJuf5vdovixR++ymoRy8mlkwicqCYQ7sBnjDVs
RnL/A972g7ygiic7lTr6V77JRc44PALr6hPCM6FAuiwm5hJvvL8eHAUHVUjfH8oE
fh6Z9zisgVILWn4tDkcAObTnzpUQYPVsNH6XjZgZROrBwylBxbamXFvxsT8CjqZU
tP2v7bxJ90tn0HWVzQ6SWbR3XDKd9l054wG8ODxn3Pslh53w7F8CDS4ZiYTGJ3+K
5DrKoFAgL9wEItp2TsShj1SghdQ0VIuWq4qBf2z2alr8DSQtlOogSdzOKXeao0jT
nozuavJ87E3C3rBDXInvu++mW59e6XJ8RkVUejESEETtNxCN3Uyn+whMgY2obzuV
s0nt1T4mAm3PY+cLnUaZBJdQ/ulRCiT0aaPXAaGqNAwq7M5M3iVYVI80msa2apbu
ltsC8xqWiVUzcPy834M+DcTLPODz7jv4PF69aieLfpsJVxQ0EOIoR1nXIY85n7r6
KuQamwj2zR0SUK+BFr2LtQEZ25pMfbNu83zATbusF0rzCen09r7COk9+mDX8/Epe
iei4rGVj63X8Glkz7I8CsZmQgAhHj36qz5akKSznOXXajUK166hqm83dc0sMsqZv
xbHA7NaQu7yLSWnvydYUTKncAt12zxFUQH6wWh8x7YzlLfz81kYYwyH1IlYGyMqf
cEIAFt7ZbR2Urjn3D2r0ke4vi1Pg4gHQKfSt2Q61h/tbzjYvXhle9VZxXyuMjy4J
O7Ac/uTOXTPzLmu15CigRLgHjbcu4KbZmpzygz6L1QgG4GtPA891BzSjMMzVPAes
9lNJ+K86sleqNepJgHDh+po0JQxNnvhflpbdKvpVWc9gWIpzscybdrERaLLYaqaU
Pf8hhxAqWWi/kYm0Jh1/GkW7Etdw9y3FDh08h6R8NfKMsCq/m7RURvx7/bXrMMzW
ogD0qZQ+6s0YOtorDhm5QW/zD1DHwAqTKVbxdHK+d0zQ/E+GHSWFmTbqi7ycYNVt
aK7ij/sPWeuafSHpVN/iM/Zb23Yd/1bMRFsqXzVqq/sT0u/Rtd3KcW25GLg12Z1e
22ZMd4ALbH/gPP7hV7QI5Rzbz4gTJja0DayIr6HP2U9S+adVzKoFnmVzI4Cacbxh
Md/M1lrbFkM6MvuZmBEkoJLObXu5wjq2auFW1vYSr+fBS4IVnjrAKNdlKKeCgzkf
/UmHuXPhzLS3cYOgrkjbz23EWqobw6vp46FjcyUFWdlWtX0xYl66lREbuxgWAt2S
1/HzTP2SDsTGTJJlcbg7dPxHXho9GEdzf5wgaw1fEXr6vt02hhHvrolNSXPvosrV
RMqN5dWYOi27YJzElMPRns1e6YMrHYKhu5IyLJJqUc6BRZUDjy/Z3F6doVewPiPT
oEjBrIc0mEDKsNKXRuZX9/3oAoY1IGJBWryd77YyZJcZwneACouw3mB2BESv6DRK
VF+7tCxVzsOemPrdpgvPKeOYhWzPvhOcBwgxRhOF+YZyY0/7mub7wJDGAgCGCDDa
ACYMRmzYLsNqkXy96sgv1Zh5ohlp2MbYzdMFlLwjv2a1R6spXy/sJUZ6GK2avxhr
kWWYSWE9s/3UFr442eiYGYd12gsNG0xcTA+XSvuEXceq+tKsa7W7yXtCGhRR2U+M
z3CyUxeUTOtdpYDttqyPJOHWAYL4J5AcyFhFJtLi2MilYaSmD/Afg2olQw2j5zLN
XuWebThbuV91cl4ggwq6ZC7OjvN92lj8Gs9p5MxQe4ofr6z2Sew2YCpbYNVxggWR
bvURZdItO7d+NN3atVZmBD6QVAOavR7m4BBkGn+9SE+5wMrN4wAscmHJHZyVX5vZ
QIg4Ls89u6KvEkIk3wmvQc1oKR8aJYJDic84KrCLAUrZdCx5KzWyBhilvxpNg9cK
s1nWHRHyr+S/qB7uQYqSw+84n3C3jsjHsHrynxX/hycwxamZR82V95s7kEIt//ze
vyenJq2E0TEcMuCU3qM0Zsfv8MzbrOBLJugjyeGFLn6yDY4ZwIkuRIRMuZ7yP03g
GK/WmDah/zXopFtF+Uu7yJ9knURD9UIvC8918sPA6WHA1p8xhEsby/c9xnQNWIjD
wwALCfjQscmOcTqFLY1Vs4nVdiRWTI3iW/W/bpZE+kgPEbQlhADrOfhkfzhar+qf
bhasoWJsKHTelOVLNJ/KGgnx+RBzrxoXSLbxrmJjeJa4P5RGaazmSWgu74ILgrMY
w5PjjRQEP0kWgCDB16JVMlt1E0I6rIEPA8fzIRT/iab6XthbOrB6f9z08IW3rwzA
PjhwmvH36OHvlWdcJDZPD6QrBXIVVKkuTZPcjXDEDYFTmyktp1dxy/DkCm1pgO5s
Orge+Oi+VRzozRsOdBFUVzsPjmkzFZYkuMZ7B6GT4hVSL888dURnWzyQcXlVe/vT
uQ/xhOPfT48aPGw7CNMlB6qMZhLwoWIrXj5NffuC/jerJAHlQ4ZkYSpi6bdb8VEs
2luwkJmQgLDltQhkZ3RKahVdTwa1QFMeYoflCcYpj6QSvhCcc6/6jKN3Gbj3iZ/b
+3OKUTKePUVAV3I3mbkDwKCHpD9D8eP5LtecypRlmFPMGJvOSSllgJs1QA8Jpts7
L8wnt6CxCw3WIUmBhdsioo8xV0L8eWjBOL0pahQ4UScSgDeBXQHYYvxs7NwScZVB
2biBUFdBGY6sYVbrRXELqg9sbndSraJLU87rR6ILe3YJpOgEl1XglO3N3MsCjiDI
WY1UaxX2v28xcqdkRpjmMjFwxlUh61DNOjec0EiQuDleFwphkGMm1EocejfpGz/x
jDYCexbK8YQwkn/DwfZVHv9eR2stnmTxdHp7ODu0vWTOIN6yjGEqXu2E1967sEJ3
oGs7BQ8t1odSqjmxqrsIapBWIRsRHDlxKBjbiymJ/gwCyK0/RkTsVEWPDpoTQNdh
oXoT1F3tJV+lyI6dJ/fOf7b0Z6vxV4zaKlaHnG8rp2V6wkEh8d8I8UeBWXD785GH
lZsXNBA8OWY+2LCcXnXVG5ZEy3fFcYycz/lWmkafsj9A8G8zLtaur8qDMRI23mXS
BkTWzEoC1xvykCBCz9PNZIDMXfm0PIcxk6ilUMSCaA0bdXFin20gqhXtzBqtX7mz
p+1t2pYxclQJxZK69/JSIIvNRVXlCwoCnRgkL0GU0U17F+wMrmnBCBCbmkJ9SnQR
UvQwQeGSTAKFBzcdv2Cpjzzx/vqRiPk7OtDd/YUf29sPQIk4nx4GuyQatPWDLcpi
/MxVtvUyIBD5MwYlVai/4T7AUwPGSQbw+RegySaj3ogS/JQ6EKmNuEwKIc1purBL
bQm7ZSn+9FQ2xxCb7wJfZaNJqUJ2u3unkdbHz9iMrpggd+VDW4pZZoniBmVH2SWE
uvvwPonN4EZhwZcaL+BleNSciWvh5mxZM/MQixEEn/lJHhLZuXlodDboO+eAX7f4
IUDVLtM6NnRQBJENh2sm7EpHhH2THDOx9FePF3KJXJA3CvWzB1kbb8+c3tcj5sHL
3dFATZQz7/s3qFgphZnd21s2JOAWQa/oGtAnqkkVUponVaOLMRLZZjeu30lzUloh
HNnerbO/r8qMtTyFM7ISQhdIgtYm3GGVOgRxUWYk5nGj3amRIKqIOoLiiS0gQ81c
M/fVfgG6BQv8/h8XEWFmJwfdIKrL6pVATi+Neqo/5tIxdRiwNPepwzSoL1HT2+m8
Bx78B+OhMU4ffYPAuC9LACEe5OK5S6LuVu415m/++RuHTU+4oPUNCi0TiL9j7PbG
mnTgqVG5N3RHRwM1zCrgYg08s4aZSOyxxFNSfpRQILSNDziC/FXWKI6a4KCR/syl
uG7/Hfve8AoL1Q6C5d0Vu9EC99DeQMxkkyF85ef2yWGKUuupWm8dPkAlk/wbryhU
TkUT4ROGouSAOpqP7ROoYg6i1xtl9DMTiHFWMKlii35SMTI8SqkxsL+Ss4p41CIZ
bleJ1QJU0hVUoQLCwUPNgNPGH/S6Zlw0gBAe6ZwOWyMusRiFsaXN4xGk1locVeTk
ctBTFkna92rSCRghkXrRumDpl4NQywNIRxqouPlFFglteDQOaKZfcLeRKGyiahRo
l7aFppdUQNGiE2Cwo3+u5PGmIJb6ddyMdQB+3rVE28dKhjKZBekLdC89ujTeZqu1
i+g7+cm7hBioAWXZ4IQSnMZ3U24ggkTjL7VqqDkbgsh98cth8nMHNilaIb7QGiWS
vmw7/jQJepRgC+JkpWSelpexUw39cXsPLEsVbomt+C6wLeGdpU2qwcj+LDInOYLz
6rFmFP2mfiwiZR4xkf/ps6oNrFyFOMB8fQfIVHVaK2AgQ0xXrSdpr/r2F2OEDONd
6uMwn682iAPAYUR/HMvEop1pq32Oetl3m+vnsy2LbhyLlUOI0RoQuKyn087wxmDj
EfC/UTt/GPTxKMbsPq75pMTXnkiU4StGjlOGAa+EBZpSQ3cCPzsjSSoG2H+RnIRF
hYQaH2C7QXYTm3SfYEcw8uhMjpU4DYGi0OHJ+a6FD9utXuVcAe2NOYYcbcP8iCtq
41bywlEgbgFqiQA8Hm/CN05brStXsTAMz9EC+YLm+xJHKL20t+bj8NtZtw2u36Ox
B+peEXM/044c4QmNZk0roTR+rK05joSTwXdq5wK4+4ETto8JFj/EzVWpSRtxv0SN
t8psb9/2cPTin0kLuNJwbbMK4E6fDb8OFCINqYFNGgTF6LcuqK4DSeoj2RGqfsZl
5M0VVDLIMOVe8MpZrEsN+WAEASRLOaJff9TqBfenpAYXOkxBTAECWa5wDU9lZLnF
/i3QA8cwbG/nyVms8OdmuYrWOkHpNWSRcVtZAaBWsG/BjjElUV82og4NP8hvvtTY
0987m0SREI0Cx/Wv+KaDNjUMukt3dlhFJDGbJ0g3ZMVetTSyJmbhqIRwKnJaWZ3o
xrndt8AdguWlm+Elp+ttA8czJtjzOp3iontIXVqAXZnM2fB5rwQJGyPLJtXZ0o6Q
83WAc8wGqlbbhCrcmF1+5aTymsKAqBVIhemC+aWd7NjmKF73dz6ljLYkeYbzYODV
yLZLhkmJByz3WrVedro6iSOHzrcK2zLD2/BlHbGcBvELKz3bKHtf6giX9X/ybQbC
f0rnDfIpcDlsXVth/TO+dUvH4LSB3JBuPdp71qyjJUqIsIAG/fKtPGSYDpkevlWS
DjNZd2NlPrkhhW2JkgW9dzT26EvboEtRNcGmkYrMdZaFpHkb44EwkIpKQ58LZ+cN
v9XhYHNJS2c6vbiai9q3gnTt9NTTpe5qMjbbLEMfjTvP4iNtCGoe3z7kzNoAZJpI
6wLLLCshbbIqFuED8+4In2TbpVPfg3KmNo5AFukVFlYO4WfLiK8IaCjbBAJEdDpw
xwVkgnVrmOTzNZzmeRh2f98must/enZLia/0w5jElsOhTvGBKaOM92/SDR/rUVJt
YpUo5BSluI9NDt3yxHvGA42+88RKOOiAiaVrxsTSYHvS8A1cDvGpwa7nkEGcTWdn
IgKmv5KZyi8wlsxoCg1nBpwaxPzXrRj4CBaWE7jVqES7SwgdWl5dVWKKO0EVemSA
g1+tOw5WrjAA83+yaoiAvtpJJWfg267vImknXMLgBNC4MojLykY0WWbJm3iKyC4Q
AFHDMbbmkMOhP9LeacAhMv5BzAASzy9AaWJvQkXZ1gE1XBCSTFpsMxcCjC4r7C1p
d18604eRBmch7dpmVdAqSoHyVgidARmsrtIdPwHt98QgHbYE8lOMs1Wla+mIJcCX
H+IjKEqf5m+WzVgYpdCF3INCsFRH3mbsfLIhid/ZRt4pcR36pjCRMgDp9HFPGcoO
UJQq520nXGsuiUV5ytp59XbivBNIUPOHvVcggB1o3GJcavqP2oKu6zTJwO9fYVst
QlvOO6HMj3JIDRVI0h9mHgLuCz0IoaskfUx5cSc3gQPgfJfwBnxUtoOxcgr9LiBg
W4XSaqbnYa0buAsF5t4eGQXF5FyTyZDyF1aPORA1wLIspyP1Adif3O/eDPsecV48
sngT3JK/ZSajxc/FKpmUARcrsZ8a0J0em8HN0YxYIVsZlzaMAtnUykDI6zuUXjJA
9cIgX9uEG5EIS5cRYcnKkIJBVuEXsVqk5GuTdxQQkaIhDn9qdrYgCUCXj2EC868e
uxg16WkiVNBzVHs3qhNQdMx4opN4ue3HeZvaH51zULvf7bEnkdmFpyGu1F6sTd0+
AfQmu+R+YqVBiKHi7qNXAo99TTqxHyAFXJJGFiV7UBT2X1Lp66Z2HBQilYTE9BJF
R+Q3yc57JN4/EME2ADAgKqLxRcvO+EQoUBITdTr5UQ1uQkH208uRh16CrhZGAGsF
+J1Wc6W1xEsIL9k0vtp2XU00IbB1wq4rHskte7SqBRyGdVqWz0IiiUib7ptF0wHy
RgHEmRJrxT/DQ9eHoma3X1VWXs/cGLs4SiwMDikzOPXVIiqtTVgTBaAiB5TmFart
0zV50w1AD1wjbALzg6AqFbWCtL5KLGMDPvx37Kl5EOAXBRmnC1sUW0w+uhV4KuyB
M5v7Jk55Ikq+JS97tTRVXChd6ijUywFuj2hpe1czZlxtD2IOlsh28bRYv9FUoNAv
LRi7OAqKrlrRwWMw7shhDfXZn3aFlyoR4NxPD744TljKCrD/cQtS8c/pdj6m2tY/
l9/cyTXpiQxstsckIFZALQob+37wMhwnq6ZSkpa8rx1zI8X0YeRBFPQNo8CjpIeU
6Uqqsyxu5ovD7lz9Qlv0hg0iC4zIpS2F7PdxuDY1+4HdQ0tHr/vfGpjwqLdomjv5
86CZdWxD/iH7cvd28HfIJHqoI+jLONmGzY8Jybeo7qr4uTdU0M4ps1sxA3BdEu8W
hWCqfaidfX3j/TSPq5gxaad6mNJ6fkFxPU3eQbihe3q3uYrcEtBUFDQu7g4+J6Va
TJfC7dK3SP177p/sghSESwyH+25lwL+DWv5R1lr3pogZ6ravVRaqn1bb1cEVW/T7
MhQR868DoWjaPVwZIn7IfzmyH9JpoP544K2HYrlv6P+ViPO1Hww+io3qWjdOSQ0+
R+bUhKXSWON4Z/njRm0I53ykz7NmT3/BIs97iOxRXm30pCBoSyBtsHpG4r22mqBv
5g82ZxK7GP9Gn/6iIF3/8ovY9fLh+l3iJcBJG0YJIlt9TfBmQM9vBvp05nxQgroS
RdpSdcqFhpBn4zGCaJCEFz7RyibxcXYJNwrvv51Ssy4X1Dnp/LsQRGMwNM0gW+pW
dEnEnGPG3oKNX8/CLWgvUxVhjXLBO0h3nkIA4WobGNuhkbIUjPWK2OBivvzB7ffG
6M/1/acgVcwJevL8njb+fzOIfSpmVQEFYtW0fUO8bGXiKGDyPdRDjXXgZZa4hbuT
f8zO96G64LOt9fzfS3Kg1VyOube5T4s3A0I4D0oJ6V6S9eqEUmn+F6CfgKy2h9ZG
rFaI/xR6gwP5HuqJynFNZx1jFZ/gwCHQKkHYamElxhL4/vuOqUzzUxiADmLbgh1B
SagccYf3KlU3p8X5ZFrIZq7whM4gbSwSkWKtU8oLnmsF0V3lhoROx9W/wW4pHAHb
Ilu9VT3iocQGrfxsj6EtUrwEwwoxi6q4KsbPDQ8ZW53tDgrJXb6svzgd2sfz/EpO
TuIMxtRgulJPBYNsQ/tdFjo7hhFyfIJ/ob8wxzHwckW0DCi7dFpu4H3gutpF5QTQ
Dr2umRQOgA+glqy0GH1VuUi5jlkP4YKfSia5q2+0pmfW1YXsp+Zlnli/Ym0H8of9
PcBQeoHMQ0E3a/lx/3SwiUerpNrWOciZ3RinrpKhf3q1U0cwwxDFRivUsdteFDcu
eo3Hrn9s0Ky9kdt+BfxEaZuVspViaua5CZ6AICRyP0EVFE+7I6Mivuiu5ouqnZIN
v2YBbrk/47FeSrAdlfCNho8oqE6R0a8LkxEnixsde7M8KVIQny4GJcUmWRCH5d11
oZaQXmCYN57Fa/VNkFZ/a0QEPTCngUqQoYogmRbJ4EXac9MFD3GISxB8XRLhB7em
4s5P43tkDcjoqSrtHdh5x/z5VeygcCSN+WyoMjO94wThiSlWexEgBfoZIL0WpYsw
KmlVX+1sgMG0EktXzX6kG8YYZsamLQi0Fdts6GKJW0QBUbB5rsbwTnCtYSpXII96
4C230uEtzNE61OmpfoWh15JnTpuvPFDZ4MiP1bND2BD7w8m2X+l0pYghDUJZ5aw6
RpnGiwV+ribSNyaCdGwnw6IrFWCngWYLRqgraKdgpItfTvv6qa5uhB7yBpXo0ExU
15IElvXXiK4R4XIOjEhiYCNDKwK32ba5VK+sDcj27ja/BWcQ7ILDmljKBX10zXM3
09Im0RPJJXA3+a6iJuMWBma8pnTIZZnaQvtY3rIeAjs1xrCvj98sudJ+XJ1YEqLU
KAoLxc+++oXk9iLuRPhRbY62fylYWYpbHyTKKEvrZ36sWTLQBQu2ujVU1JTd9cy8
l7yvyxcRs1XKIeZyIFu0qaUMkN3jZxohkcVzRPu/1JDn42r12eFgf80wFrze9ZSD
AcSnujCGoObDcM4bSLkqdYtQR7thD5UynfosYViy7Fs+UxFVS4LiHNiD76JPozmt
TtzM4LTE9YtG6QfTFCPBCXbGZkhvdzG9aYPn8JUFY8/N1vbUQHsi/TpSJ+SaDh2E
K1sOBMa8DvLXBj0uZnyKUnbcqrjWNdVvBlFaoVqrsRiA7jWpes91LfH4D5FHVt6b
flO2WP/+ZIWXIGReM2QBSfZoUbAZ4jHt9SjmCENoQ7tIftYCKAlOY6KBy0Robxod
VYa+Mz7Exc/soAz6rTxcOT1gz/V5cRaCQShS7O5tQbya506COIUtvsM/RPwphHoI
DVxWfx+DXw7I3MbAUet1MRl92xxbK8IXNfsG8guquXsK4K0+GD9vEvyeI/GyQtQB
6YkvfEqWsrDrQPIDOYBiu5Zo6a1xANM3bHEd7xp7uTWlNiHq+VpE0Fc31G2GwNH3
4+AcKGUA0n+aqkIG0OeC5kqIrhnVIsWH9iHK5+2AKh9ygPXaGuKE3Tzv7kkkiR8I
qlL0PEzDvDYrLrqTDzQWK/KXKOqC+ZcLMWbDNvNEqoqsOP2N6ZXCCnzaxmUCwrOz
w1/g55Sfmx3yYHyJYgwmBr7sYAHgHvjXznkT1hbfoR+y+1IxOYzpGdgIRVH8lBFb
vGCiPfCBp+MgP9tL6iMhkO3gWf5soZjoJk6N3/J1DXDemL7C1q3XujHmjcqTJy1F
DMJD3WHkGjAHuOnDpvFmOVCLC5aQZiVPEKXKAbVSm2xyRfEJS+FOGGNT+j5u0njZ
WjSYr4pLo4lXnUBsn9QM0l3sUF55E4r3DAQhfQLykXOgjqh1S19ph7GgmdSDDEnA
fh8kdWsBrfBcKieHBS0+KjZUbizMk0lg/qMocL44VQ0JRebRR/tgZ/LTs/ombKzp
Porf5rt4e7DU0BfsBPxgwAfySiDvqY7pwFCjdMTsQQOqCz0Abp9B4jw1rFdoxd8s
w+Y7o9xAMpHpzC8wqeIOofFtUn7UyBfmyc4vl6WDqnQPPvPLXlqlnOU4szTSx3qg
2UzB3UkOCU+Nvx6Ft/lJ785pp4YGNHevf6fcyxEA3VI3bzIpOWcBUDEwBJQs9DLl
g2kSVls4p4iTjESSk6LN5j3TVax+bDOgkkGnk9TSntaJ1Hy+FnoTbk/0oQMTke8k
iTQmWCnLEK/e6Lmu+K0MVD0fkF8KewkVx6xlHnghzE7zQigNFV1WlOQkczb75IBU
qRcqnJVUeLrt/GS2C3pg+1hShbnfrc6U+K2gvIXDTdqJPTCnEBoGOdN96+eEi5mA
Z8+S7xUXSMKfeC9G4K/W7T9hNPkLV44oLsBuGiF5Kk8nPUgwYdaSV+5RP+GlQiCW
C4GEYiF2UmjEnOPaCnvo1yj3vDl4ou41SvvWMFo3Q53S+1wBrwDRolyvBTLbAUyZ
qOWLlCD0G8irkmPYfu1xL3W1DCk+hIJ55NUrCvGT+HptpSpU4VVXXU6mnXdNNv4P
W6MpRV2dFjjsdSs1QtqOBvtftLFY1Rg+4H4VBl3WZRvOPwu6jhMTIpLUSI07re1c
SplfNLzCoyMTBgeetzfejG1SEV4qpMAZR/YZJ928FTdw9vXlfXwukGOhLaubmTqI
hd7QULhR3wKBF7KeO6Oo02cwadE9PqKO/o/xHPazCN4m5bVoqdBVEEDQ/X2lE3iR
GwAkOLk/HVL7/BASLaMm3WjQ5eAXIVeJc3mO2rKUGUMxwXeqDfMZm0sU+EoC5B/6
RUjvFC62+FSQexbrZz7gzhde0kVKUvB0NsZPW5s/D9OXice9mE2KfPn/7PtrXH4x
+GJS8+Z3Uke3ocGSvP/vt5Hw+vqHNlIuPjmQAFt736RnYwz6fuF4RIF7XunRfPPZ
XlEQfApMcgF9IkJdEL5tyyZArknVrRU4szlLYF8EiStuLzKiX7c1ebZUa0ccagaE
nF9zXHkuTRfu3Nh8WzUMB/x7/mNYsSu+8zYLJcKa6r3Venht1jJ2hW6aR0YApn6b
LPvpgKkYXBs/xQ2GoJFqFCTPRYcvo4iRDRhnFufSy/qkRWGHlShE6eHNGjeEKC//
NW2gD/0oc67muBcIR+CERVvjV7JwkOO4pzpRRvc1cf4UBod2T/NwrpxHeUswiGOR
yOSREZ+ngzfq31PY12grAQ8Mq38Gq0fEBZoWfvHtwa3aRONLbps3FKK/2mkesmnk
HhlMTFEpT4iUrse3BglDG35gxUHFHM3z+7sFww6mdZZ0AnxWCEB5Omo8Hd0KCszG
suy7Q7oDzqTcw6ZXypk0wenKQ7q2kzbxUBhH8QVtr0ca5fkUUc1oOpoPkbz0eC9x
YYwSVcJq1BaERmqpIVmyIZ8p47jDWYVTywTuSUPGXRe2qzlYrCmh6nDlGWUD+ozB
sHQxaW4mHGEL9eKDiokZ4LMjtYXrREveJkpZRD1gmCAgJz0OvgiVTuNiQD5BD/2z
yzuozHP/9uMKixCpd7AZUl7TIES7tnPkmx5mQgQGb+sTSWI4/HJ20vfYLsCvqLMF
nlHPok3ePTn8IK9uvFc8lbLV7KVZnabChFKYCVcjET+VH5Z4OsjWikoslMBliBJY
iSfLEB1KzsvNmozBbT/OUSRGHG2v3ROXiIr0tMgq/+SlqBhswF87DR7Qrw0+yG13
0oXS79xlOdmG0kO2d7ecWfSWghEArmdaXTvlVrD1pHACFi5LKafZdwL6RA273KSm
Ix0L+HFJUVZfHjYI54fkat0cGeXUGeLSfhji1v+pY234GsZiBaxGUjsZH/NhJa7C
vTn0E7Oo6kqD/yG7/fSgb6muM2Elk7BYGw5+YhAMTtOoT7NzmlDHC7NbXNL4mAaA
qRWcUrevO5cTJU5WY3fBdvkBPqsfbOx2Fsnq4rvPq7OtB/dEyvS8cEZMxUTjNg05
ro6FKRUg0KMJo7LapmE5sJUV9RvY/DWjsee8N/9C8lpeNWjqpaZqYMDasTzFp3ga
T/V4j7ajo2sx7cDuS5ZvTyhAL2dK0H8zIMB3985VHcJQRl/Ky1CTd2R/GAXBxwbl
5V4nzELIKlhsR5JuyklYCGDEiO1RWwuBcRvj6yU6s+hqB9UURjVSmqqUQaYt9UJF
7isOxDzu3S0K1KGMxbcIG2i7rVf4XnZ22Y8H9Wg8qaTFlGIzOhHaw4cUnVwcUJds
bH6p1K8j1wsok1F23QywRRkkWnm61xSNhtZ26ugu3pxrZENFl4+JwbqrES13UNuA
KY4Da4PSereeaIpIDFWuyAzBjK3kfd3p9VTFCKi2GMvLEc3GONZI/mXP1/9GwqPX
tER5BzgqvqiuMrqtu/u1ZqfTj8FbabKqfe417jg63h/Q5VmkRg5I70YuJSOE1QFw
ISfnVpzSzMXStsqEQCpRDg3Wz/17LPcYavWobemYBHSnIrY6ns3HUgCupzbTA+qT
AabtTkt4Vddt46EeExGJ6JLay+adhF427HEuaakxej2wcPcEzF1x4j0uAXVEWn6N
AiQNGV6pDfEDz3bRRsx+9FT56c6QxHY1p4iZcBLz5bVKg//CGlJ942Bmp3Z3EI2B
sJR28M2ou5pPDwC+V3lBBgR61G61C9Wd5SoWwxypRM9TcLPzCnOqjD858IuLRoXf
PnUID5Ddt8lI8O0GU/GXc6DIY3/F9EsgW46jqPGSwDOyifbpn/sO0bmPj/IbeWrs
a7BDGuSMOJZbhx3RnIf3S4bN9cX0bAxzPmZ6ot+/HocRtQgl1aKefGXXC5XVARrN
SmQl93cjFBaHSL8e3a4J9pjwPgkXH45FOz3yuWDF650bXhHlq4ECFC9IXCeGu3qz
Wtw2d8TyFeOQFy/PGqTUDF0bPtlaDl/3vsBydIcQ2VWrG1XKxfYBdTWHTqZmxPcC
vgxig+akK3m8VJ0boWHOHXzKAP9AALWgZ4hQQLshsActfzp2/flFha6uDpnaw/D8
R/tCxPR39VBL7bHW0lmoHD46UNULBHLbj+eP23gO2hGihjk5orOT4/37q0NSWeqt
190oD0g/XJBiu1eAM22hF168fEGe7ZArhds/J/izmM1d3YttLSLQfdwIGLnTK7Sp
0sSakrIT8vaLyRhPkonzHMyG4PznfrID0a4pRPm6sMezpl2kx6BKaNCXDIv6S1JQ
izAb02GmJJMTI+SeBupbx1j6iI1+KjwqPcKTBvcNHCSyHLO2x6B7igjlyW6hpQpe
hSZs46hg70NY1go0N44SX8HuSdOe5YfZMRjLv9acRT999wyeNFjOe3xExOsDlVrd
2LfTIuxiDd9tNnogNQoZVDeb5oeKlf3N+j4TuDoWOayiaksyyh6PTadYSPBUA1Yj
I1J9s1sZOgVgiJx5fUEIr89eNY+Esvt9pT0E67YfRTmliV3urrSn+o4BnZfcOsdY
pAkBf5mkC2ZeE3/LeoaFO65ZDDCzjQkt3ym9BMXGRuB8HL5c230uG1rlrwp9y29g
U9LDp53OtX/GP34JD/MMYuiZch3NddaO1lRVrUD4tZLz6xyx+6AmDel8YpH1DAwC
Rw3sufJ8bXwj1QPXVRW+XQvKKs/FuDgNVx8WAhhCzr43E8kev0nBiiD79YwaISze
vF0UHxzy+oPZCNloHb2XLJWU9HVGiNjQnnPzXyf/n40dZMuKBfiL7lD9hl3mKIyP
skRRLfdJ7tyhD6IxgBhGePSi+Sr4Z3yintLwaNQF9vA7gndhT1sghTBp8lsgisUb
oYNParAT7/LCA7GwPsCw3J8Ph6o4dWw4FfoPWcNvF9hwNbXlKW0yGwDkySLexWOI
z2jL1A9xo3HDcal4773m9Gvz4D34IxzMb5jkreNpdRt2uus+n1G6pCI6x0HqYZ8M
k7haz07oWXASOCEIN8zPB7z9hha2Az5+MjPqgbY9wXQns3hc7vglglgJHJWMhng5
yxVjQ7x+7LxMXDrUWnqmegkbjFRc+nJJ0qVNX4E+Uc8V169s4y3f/Rmins2Uolu8
DEDAiif953fs1NC7arix0ZllbGa0je4bC5IBdz8JE8p1DrKvGzvblJDGBSTch3Jz
kWOJJJpWcptDJTd6HalwDR/3VFl35e+2HbZxGYKQLZhDXDobe+Pk6My0LZgEO294
waq6PMO5OSc+Tw+UNZhaLavE8O85mlmPnfNdbqq2m1rydkxmYolHNZr3TmLbAMMd
SQb+8WNeZeflFxetaR1fFdTQvYzy9kxz6OkayhSrEr/WjLWQMe+YnD2ECKgc9MHw
f8nF277BXi1YQQY567EWdDrOAYwgVhmX3F6I6PZlP2hmjWPwlAn7tIK3QBWi8bfM
MUSv2ypFqKvL64J+UIB4WyXtLNwkX2fj9ZWdK3v4MlHbI/h4TO8f5oW4m6piJ4iW
3rBTtWygNnpRqIM4M4a8q9swpDvF9Dtxwy5TqLbzmuzAw1sItpPpPgvoVO+11StH
lin1e8PAY6BmStsQWcMkVopPjTPvFquESLBgDFyp5saCqhYzHZ2TWqJNNGAo1TgC
8LG6epiNEpt0yrRgMiqfjaIqbT6jcVdenkJq0IefrNp8K95TopOgIIOWsSmnm9Go
pUAoEyW0Wa34Shu6bFE3Vm92AraPd+PPZ0lrKc0rtI/CccBbMnojcExAugeecM72
LqQsgip/GquHWwRB5gg7SWLO77lkAkuwX0MvLETeh/QWMFwGdHRAVHyOc+QsKkP8
F9Mr5vtcUTa41YRlcDvjb1kSlhr6m3KFZFsH/6JdHzaTVpBbmnVogKnhZIYnUoQ/
BBYnXYNNuSpoE9zwp5L9bOlGYPiQXo5IdT3wMxi96rdIx1mmZ1smzXX0sBqSSeHE
yjAEOf0VfWtbYEwxAYqwl6FhEmX4+xG1c4uwHTLwYOtZcR45qeTvUdLRGnkVrBxk
XfQpMwY5i0yHvl0BiB3MCl0hQvPIQcaKOcM5ZG4J5sRl0HLBgqEOVzbRslH7lT7o
/GwXVZ0VnH0WKMnMsfOmRgaNTtVyjqVvdqBYjbKPUbrUBI5Ioq9DXs1jk5OQSp1e
nFijJTKEMz6nsDYIW8yIAA8mzmlK7ZWWysqWj54p6e8GVYqQuomh88j7fGea8jyo
quqbziqYbCT2FnE+xjDppBKCjncem7nzSWGI0OURwVRh7jDh1yoNIqoNynFZEtxg
taCvSh4Cf0IxcVeTMUeOuggVnxgqwh+/bFs9Dxfjgu3AhiRh8vMZXZUcD77ezKZk
IqC6cfFx11kcl55lES/Qae0RwW8z9xnjRfLzlLuUShHV4jP3c+1g1FKvFFM0uF/9
peeKjMmFNT5k5K7U24Zbirt0CkVI716w29/nLXYghiYe0bbcpF3wb0RfO3IowDpQ
TAxw01lSot312fRosjtZNX0devtT6k4eoYY9aJXXAWC1zbRqgbwJuOpCDytnH3v2
iC7VvovRK6E/Lwrc2g9VI46B0oqHXUlzI2r3NIWDnyVb+djvVhsigd282mdstt2o
JldKDGql/27lSvO2/RpOgWMSFOr8fYT2gmf9JdB7JpfJc1FxMFdtOgQABs9dnoM2
yYtVxXe62JQqJD/rI5DidQnzQVtyHlzoU1bWRhDUV18sOsoCgvA5Lq4UuYdojdn+
TDsZgruV8OIMqfG7rkxFwFhaA0AHZb0K7QgK4qSE0jDYjVdBsbLTMGcTxSLnhFBi
yXKRydsGBleyZ46HMYEg46zZ1fqgAq1iBclV5ESEplczLeIlBPV9F86YmUQS0EDx
BWq+if/UhXCvmL3BWE9j5/4uw1OjHNnkudHM0KxAycAdf4Hx/sV2dFx82A0u2LsT
/oH2s4Y7rneolwsOJxphgWHv+DjWVnxYXRBoYlmbdbCKzyAj0LjLUW148BYL5Ocp
Njc8S6IydVEV1S+O2/cM87m3QvY5OYp7qR44+dYsrIK7pVV+6Dp9rhky4RFapCEq
G1HXoWa0HM/bxwvimH0Egq2c8S50/PthmxfOpqP9W5bnLmnoZ6kXUWxmxq/8YAZa
SdNuF6X+Ogyo8G8cF5t4yesDga0khyBudSqjGusu2gMQ3oU0KdpTjaE9nU7zs2zn
O3K7skVNanZjsu6uO1gWmtjs3nDM6Bwc6W5GQmBk1smPBHEnmKrshQlFumMvYjWx
343NuvX23kZEZeO/1nWjJLJo4G8PrGWObS1tNH/7MGEPqq4zkqeqku71O+PYT4PD
2EgowbbFwNUhmXQeeIOi2bU3WkHivSkHU1yAD3l6ZDYq4MOY+3FuyHENujtK6nrs
6daKakXFDm4OKbQ87lnqoDwPKielCyOGaBiqg4aguJc9JmmYq216wx9Olz9Wbuq+
e6jwWQ2V1Vg1T3h0RfNsf9ncgDnzct58H/gBN5ZZz1PJ6ugdIUiYq0jTMYzqCVKz
N4nPTXROa+s2HzNIiiBH70zU7BOxNA3ZeXMmj7Mfra1kXqMXyNORelfopBzacM/q
CC5ZR6lSh9XCdJ6b9Cx5WlhFFhCKbwYot9Qvq+fFWphVmghqhxhQVOsdypzDxtaT
QYFQNPTo68jlv47Lv4J1GtsqitPb2exmzpUTUeNrrgZqworYSWm81gnpKEVDP+LE
/uVtwn+4vzMMcdPi172068C7TVtKNHNnoi6/U5BMU8jy+Xu2PUzNLR2dRK/tTEiu
BfEsTWQpX5REY32Gn4ACyORRVMSSTPreHexLlxut2c4rLY9vzGFd2oJrQhla+LE0
thVIZSsSW1grhpBkvfVJnNem0OBmlvCqj5Tur2u2pUrPa0Uw0aJ0ZRX/i5V8pToS
6p0z5zB2UI9aZaJYmW0k4QXogQp2Mq9TlnyQ5ogLmLuNaY6UchTzDdg8tSD49lfR
dCi78174e1OwH+9IW+rZ3tQHJ1PS4BxR5UaRYp/6qBRkSiXx0pCra+udKhkEYZvr
+7dHmO+B24dy90LHFFkCckdQ/wZSaueQ7gH0V4QiuCmv2GZbaidpQl53Xtbz64F0
4cUQagNWsmdJz0BB3rzeYlFgf9njUzerzuqpO/ZPjFToVx2hxWEJwm94w0PdQxxJ
1FcDxzx6HvvnJK9KXwxT7uIKrgj6b8z/R4O/ohIjWKKaWGptxWXNxalphsoTrgCY
9UM/v4S5mUG3iz6syEy2WMf+nr0jv5ZvehLO/nx46ln97UNuuL6RB4sE+G6J0VxA
RvFI7VJKVKOgL837p4JawHPQYEviOEWBs9yXV2lQ2BvDok5ffAduiIF+Z1lf0lD8
Cv3cK8An0tmiE0Xr7VRxZrvbYziYcW5x60Me3bvQwpKshqhlT6oh/+VDVlqYdBZ2
jogPXeSAIjkAHiqqeCRrDvH1LLdRmOaReLlBBN/rrw4i++W+cA/qYVTloxSZqbyA
qsxotY66IToTd/fPLR6ubcet+R8vR5eVmCPLTi0kC0+xBwm5gMIkJExHOnPoDUUt
Hq4WsHX6EQmDXKCaoN8AmKi+vOkwC3HRvSZEO9bYsrwf1YToJmjWuP1gk90GCvfT
ECdRdVG1gcJw3WbOlY2dQTODcHwzqr6KSjq99xVha2zIJAuKLb5sbh7srupniZBx
GLiKD7AdTJSpirhEzXodSHPU/4phC0Cy7vh7jNdP9LD9gVvERZWVXiWIDWfXOVyC
JfL39BjJAOPyWw/SyHiJPzRAL+XOt4nsA34AvbyNFXrHfKYHY2Yc0SM3Wspzk3Pz
X2V8QMz3+j7K7UqJBUCZEpZ4mM6u8sDyIZ9WvFT6um/eBtxQv8MYQWVg0Jk7vRZC
Xqp+ZqDapAo8cYNRHHpiMPsvM+/9MFMSNMM8ZbauHbmj9Mm6bgE0QO9NVk1wdPkU
lE+V7dnughhHqlPrc7DbjAp9Kk81bTTVw6lz3mS4yHDHKvsCsLr4T04fgEV6NOnk
Fem6WzbagIT0S2kH7OAWXXC5shZdkzgZvSRKxWkNOYOCUuoblMj9xlRxauKCj+x/
u1xcB3oRj1xYvE3CbG6vSP9smPVH/eypI3TPDMRr/zIc3hQ2ZT7jwmRaWXdR3J4v
2cTVrx0TRH+o6b/GF/3Uu1QlmYSfPxPhOYliKFSijfWRtSd94npTshJFGwAZOXmg
PjoU0QjhWI4N3hzwKvM6ODYUYEXZ7rBG9XJmGr8MiIbl1BlE5m74GN1LQrfsMxMz
8wH6HyjAFeyS98TH8ku/zIXQ0YS/x2vNC4bLJDIRceKej0qcvvOCOZjp3ggDkICn
sICbZEuhXmKkN6VSQoAHYfMn7Xex616JNsb9RX60e6cHP/YiMv766bZ/2pd5PgD/
2+Q2iux0VyqwtBNLlf0tkXQ2/+BsTx2OBVQ12lSpej9lZQVkbIlDawt2ppkRneIN
MMcqiJ0HrOXqw9tKpN1lLiEuWQawkqRVmORoFA6KggS/P0OoQikLRfHIJMJXnAEW
1RxB+o6MNqWf+hE2OAF9i5fbidmwUocMDbEDZw57NQu92WCQq1CIaHaUe8Z0Frgm
ParTBdd6p5kBlXGWcvUXm+R+KiK/e0u3+uAVpWo+4siyJ4npLs47skUhazcBeO1z
dYsHr71xVxgLYZJQea3xC8wBcSaSZIXWzoWISH6TapItAbnDaEI2GAjXX2FWvKG2
vZTJ23l4FXge3OqKaFm32mK29a+kPWj4usSqPXuIhfcd0q90RjCcxm0BIJqDN9bb
4tRCgQ3mRwYnTRlamCGNQm0A9A2IPjVqW+lri5mY4M3H2Pf2FFmHLFZgQDvinEp2
/JpMmov1YCtz7XGM2fDgzo8buc+AwUcPLRTd7fvtfgq9GrUkyWPG/Ym+hgCocVG5
GqQuZKUvGwdK4U2RketUYbH8BmN9jIqw7hscfQkNSRyGipgTkXb29D8bi12ld+9O
GKfPAkG7wM5WTkgHldqvvtgfHeeWfooqfqEpcqLaMFG0uZeOLF09fgFHTF90oArd
8iZzGBxstF0PTdObp/GyPqZ1Rsr09QlQCFDrFv1Tza9whra3flMH2/aeh39SrcHl
BahDDyNT0TqDrfudI9wsvSRe9Qg6zYQwuB2YEMN9ISgxciovnXxAEDpnLmH0PcQH
vCX66yHyt703kEul5KKQiPQ616rHHS6SiRwTQiEJpsRA/4OfX1tld9yANm02IBTv
QmP78JiCKhFbquEII/6PY/OBxbN1O+TSZjZ+BTVdWzl5eBjMcQtY8ai2qREurSRq
6XX4U1P4ZcwOzAnhcGBrKmyLMHml4LgP55LMyJihbG+TRcdKeoWP0zMTG1BbXGVw
dm14ac4nNEFzRkSKJCFurJ7p3aRRhAuPI0GaqH7EcVRAmc51l0Wm2Is5QUbaIzCx
OBEOyewaDO+wabJqgnkQlB0ih3L2IzfhJmhBqOoORKSDkn4kWI3YznOTY/RyeKTM
AiZ7P9h6JyS13oDxA2KH5k3SL+BUfHSpre/0tsvawYjj3hI+vCLoVT3+AFya48Kh
/Mu6tYt65ODxquY3yGVHTM4G95DWMFI+8iR5T7ne7vhnsvDbMbIc5bqnsn/vVS5p
mDj0pIPHzZb43jpyGwxG4WLmbL3btXi3UWtinUzyGnzzappnf3MzVZ/alLb6REFK
Fmr+GM2P0/Q0tevxoUEK7KqFL12vVYZmk1Q4CbeCq0wexJ/q1g4H8MqTA374QjMG
zoeKXatulUNQ3yBwUmgUKsKzcee+WxB21jwTV6+f+L598FzD+N4JDqLSX52sOEye
c1knLQQ9K9MedNMV37FncWL5po/FNxOLIc7oG+YCFxgHEhoiQoHBpcwPjQ9O8XIt
ES1lzCom0eGWmpNtd9Zw0moVjFhvV1qk9qAls6MAgA8VcWGc5RoIOhT6Vt5Tf8uY
8WlyBngBf2uTHkA+w+knFKcsnDae9YaXtPzad2tGHfRpw5+Ip5wT6aKPN235/664
x/l8B/J8iq6qbK2fAgjeyHbwCd53BF+PZrA7oPW8JTQYpFR95gNRYf0Af4iaVW4G
sLu05+UZD6Yau/3LktubuI1XG15UNwpDJllXP4VCmQyvewYS9DjcostmbDLVqwlO
ehzGc/sFpvi2NFpwYfcJ8tePu3+WdT4WwjNY4Xc2/UGeyj7PaAVlp0MUnCPJNQh4
6SkjtiID/LWEa9srTmlKHjWd/7tBCxv50f+IxWG0+pULc4vBqO3GxhTr1tgOFwBV
DODi3NAp2YMW3e68BlYBK6s2dxcYU1Sfn0U/RgP4f94z62AC4QMqyKlWs/XwKt+R
qDSe1XCRIUnFalXKSO4SuQp7twCxmvBUSW4M9XoX1u7PNGOdlPSm6c6tGJJEs5WD
asdmZdyoaB4g8IKtwgYAuKJz6XWInNgKXEdkxN4OoyYKdUgnZSvPBy3P0annhNaj
Gn5Io2x3AopopKMnz5h3yNJaQ7Z6eGyVBd7dIwJ1McQXeas8xwVq+G0FQc52K/4+
5Es6g8sgdRwoHMlEwtSG12ZoNF4bXNBDwQffR2RhvjO62yGL0uIt/Vo6SVErHpEp
c6gH4vxWypvBScPAk/uwoCf3RZIBNrGai+ye1+mCE6gGhGxzgDDs/1mKEB2U1dKY
604OoAKM/WxZjJWsC9QFAv9iJxz8IV6Ew+XznXRJAKh9MJq8edhdHbawk9L4T+0o
XYxu3IZQhH5MMKM+2dVnVTURh4VAJcGjt+TkJfOHAzAKpkKr8ak+OqKJMhiPYlKI
A1tz15ALPm73LRH7WHZaIM+UXAE1DgauVJLkj7BoPg/Ljc1oSqxdcTH/9KCwCiut
6jJ3VozlsIX0PwAQyEtNeQs6k2vKWmJ6JaAh9ik2SIjQBclQE8ZtIzFQF7DVFqD8
5hIL1xnroD8h9XGtntfrfyfoX8bhcNAN4LRV7gJFH66YupqURQjpWafEf4PC9wEN
w6IFT2BmbukXHhI6XAw1MGIi5YLygF7opZHlZnjtdd3P4RQAVl/+gwc08puG2uKj
xSUmlVXx62MrXdVWhOmd6k29UMaYVuIdJwDbudD9DSdklKcFNf12MWgbykDJda44
s4czTkaJtR+PnF7Gm3DjSzsmB2QkeMvgpAireGMWP87rcG3rC3+FBa3MbuRgfeC8
ACm2c1cYTjLflP7KqsfOUfWawnNNi/U7pVwU36UH0g5cfqcbAM7DX0qtVe55W/Q9
/e32yYok42Mshh7jhrzxFyNZ158XN0Ims/JVjmUr5bQNFhmfQgrhcQnP5c6vLDq0
JrElnJwlag5QorJ20oOef5iTBk55B/enwh6E4A2nyG/vpER9YYigjvVm5s+Z3dhA
prnu326QtYuNgY8FUebnceJYuAyS3GX+8HYeJuoR9Ad5dCiVGlbazopffmyxCUd8
x4Im4jjH2A/jmv+/BsIcWcViXUBEzPqzi3z8qYIEsJIk+30kejL6oceEP/f6mlE8
ztbofocp6trzVHMdIKHnf4ru2TtRcFc5iO4oPwlRx9deVI4LdE9NgApg2moXDvvM
zogr55fvNvJBfnjC/czaVfXcOQcnnBAJdk4m+GjrgFyPrg4X2MqKdP3bJGOIHKMg
A1kGRYYXt5QFgaARW9jzGPdfZ2QpDxd+W0o2O1+sax633KU2c7UH0p1sOIk4cg0r
4fgOV+vrx4MpHwfWELZtuX86bWPjn8+ykUXexpeZRV/YbonMYkEv8tzaQeow5UrJ
MGH1cS4yoYctptxdprcCRzU70XAnC+DbE4UZdyvEuLfTt16npr7IFkmbBd7sjy0e
C5S5CB5L0RQnTVCCOLigSXtv4ZAPANTbALBwtq/lhuFnhpgtk+7eIO1bwcigsyv/
eQ7rzpe0GO+DnHpUUoTmEkkr/wzCUDLUa52u8Td78rFxnavQ1DqkjG1iz90O1Kmz
j35FbNKaRjjlyK7Vqu0j4ri4OThwcrEHrAuBLzmvGd8e2nY/WhVgkA1BEEl/ukt3
2IT31C/OYj80s+6qaS5CCEiWvfS/PijG1/pUB5Gp6Omc8HIcOOW1hND6+ccW2BtN
BIslxR5j+J3klzO/qxRKQUZihgPUtsC3bkLTTVupiQGrVdZLOEJxdkuiBgrkwEUn
jGiqxxrp4kvOeX3Efg+c85F0uNZtAMiNNW+vDQYxSOhYwhb5vpp4P1samijezGqm
VcoPS3vKHlKQsfxEFtRK7XrnQER4ENcoajGTciscujFojtC/0cqHKmfbiASVdh7m
mj05dKZx/m5Rx3jGfYG1/cIwsuNCBAUZlrMv+mwHD9gCYy/4+kpDp4krEPMPWwP2
iTnLmlOAlsfJokXM0Ny6oPzXG645/V3ltxOh395HjuJMDsR0slsG/pMFYyKrPMXk
3yy0PIqEIzEd93A3kbdpV9ncpulX26slXpvC7BorMShA9yf9HI32Ou/DY9UNcoVY
6aUQCbMF0g0WSJK//L3RYVBPgOW4DvcLpiPYRRw5096zRHpce+0Y50W5xTQUmfRB
lyvyPZbLrwlsFtwkCCyC425UVpbR8CaqDjmQk40B36Q02U6lfmTNCPyK1mkxRz4q
e3iFkN50/bUo7HYEwUhlmTa3S8QbmuZFPtsKuu9IHvHCosp5KrjGe99iFtKDzFI9
zIG751ckTwE2DpjSW8MsUFaZiNbybooWVSIR6FSDqarU0142UzqFMivz5YvzpiHW
wssyn9zo+GXxlhEGMF49cr78wZzBsVKIi+JwxnwNeSv8lOoRwabkOgApboAKTwTI
zTbjoluzlpKqBi1yHS+nqFE/hBXg7yaLDxZ+9dxus86d6qRWvVCnzYeC7IKopBdt
VAt+UdN/h98k8M7EqtMU9HBtARyREBADOM/uOug7O5XoGAQxu8rrSp2STqW2kpAA
oZt3MqGYDsklc444JpsUGm2kLtdx6YtJ8dbbB8GyJUofIrpP7We1fU1PMn8+JK3O
ymEqN1GLC1yNe+fQvn6kNjlEc9f6IABKS6F9QZZz9i18/utr/KFdRBp3qMcOVDB/
gj9t81Pw4An9ZYwsuhriICLdeDGTTvHt+vLG6sU+Wr0w+cbDbFpOg3yYiy7VNqHt
rWlEoYUkMXagVu9DAGSGcez+XuoSxSPixa2IthTBNkD08rTuku15Fh2tySJsPD3Z
mSPRNwKFgoy0R7f1y8AL5mOySvGbnCeixGqTmBkAVHZJYL+sHz0OokHW1oARaUsa
V/H1Ap88kae/ixnKeEt9LkoxXyFthu1RkIRcGgZLOE2Ul7QnrAbgXT/SrLPZfK5c
6xGa14qg2qY4fbAgQdyEKp5BCZ8yGesGi+gKwKRNitHRjMCwGihle3FkhT1APnxG
DrtUSyTBhjHabsQJkjHY8lopmrNrxiTXRFRdhXK/Me3BLAdB6VdC6r4lnelUC9Dn
1XBnUlp04uZOHGoMSIw9NwVHKfv+DsApAruJ52v3iLR+/UIizRo59oRgYTiYJW6I
nsdTcISlq0JWhmoUGTOxOZITtqDMiNm6mdHEYBAuwg4Css+vMwqOnzWUHoVPcecK
/AzIAQkA/dPgsGrs3hWTQEhFYMmcDsjfiWaRWU1b45fEr322JoTMPPxOO53OXWOS
sNT4xmxu3ZAAzu3KEcigVg4iGpD2Y6sy7ihwW3K3SzgwJjv4GvgMixn9gWKTssIm
bIYZjFeskxn+Nby76/5XlZmG3wg7l6OKU4igEot+LmJY/gHhapR5PJm+0eELTuYc
r1wVm5QSuTO0iAVgQhdPP2k5DK6ckEoo+gZdrHpbN9TX9xBO/hXPBh2NZdjHd/j9
DaFAzGfZvXUXM5j9aNzQY5fH+6WQg6rhb004JqRJ458voPXrnn9Als8oTSVs0lyz
ukXfXwAbd4IwnH6MYMkvUN3iUTGifiTeD2Kbq2lX2qJg3oWJDO6TcGx7aldLTWUm
pXh+IW+1PEk3xhIuHaiwFezPhs+YilF0mdfrOgmtA4eOsX16vZpYcJJ5q4XNKle5
yPRdmoj9VakfS9ZWSApzLWi4gY+e3Du68uiTA/yHb6h0Sj6C7299/70QDqDk0agH
O31aJCbY464wLg7R26HK78mvT2QubnPbh7I45is3WXtf6o34E8kNtPSRBfwGY9Oq
dTSSBmC5Ukir19FBrUOloYB1s6Iwz+BHl/u2GtmEdQGEtA2xEMXShj5hKkFHC1Sf
UWAuj7TBXvqmiaQMqU+2Obd+nT0hOn1Bn0oUEJVrKqjr5cCju3Fy2VXiw7R3go3+
6U0FwM6snL7nSZKYd5ztAGDqMEBLXVLipqd1NThKCqpKPVGNPlWiXMvg4A59T9KO
5K093PudkD+NdWku4JDZkz90v0HWhH5Id8qOwLoXqLIJzm2hR/ArQC5S4WT2NB9T
cQS5A8CUy2GAYLOwOd33v6FatLRaGWipnItAdQGdDYYYe1GgQtQJoqzh+TOy4WaF
766MaKwIP2DdJ30zBFCj2WgzVh8o0RRqLFe3teDwVdOLd3tr2C0Oi61n+YbI4n1W
qHYV0g50NisBem+3hfl14RuwbyNXbeGj0I/G5BIN+X0OLHiNYKvVtMU1bTvSWw4f
nlgMQ+6mHfOsalDU7xxF1nacHVDX/cUVDKqU/PK2gXxELCEvWe4tZL3tFnqtqTa/
nGp/OupjRj+p5UXNPoylXvDTGBnyDCBhhhQ2BaMxoTBVAa9duOmSiDj/aiqe+T4Y
U7KAoyyYxZL0E4L98FDw7cRtSE0nM+CZGJX+CnC7BYhIxdnTSVJFThUMESJvJ76x
LA6ZMHb0qQA/JIUrsvxuQf7hPWqksq29ACglFo0TAs+GtLE61WSK75A+o+/YiIvc
vJwz+25n/YZT/0+iE3kfZ8lUNMpm7lrfZlnMl7ildjQGlmcBwtfLxljpLeGFPcvz
Q2oQQBMoYQDzYchlm/xE+EJuvI5VUNNrdLWosxTK89HQbC1tljpwOS1fmqfBkuEy
uv5BnUblCSRBkXG4h8DtPKRIjmnXU5SCHDBHZ1K4uqjo0wi1fYHtoDji6PONEOq5
QeD31jiq/dUEIg3wFtTigPDY/1zqeL8zY9Zr17zLKznqXlS64WAE3dP9q5cbw5s/
vL9etbv2ZKfy0xEGG/Zh07weNhnUw0ZpwMhhdIk40zM53CzPC78MDVQ/1RXpA6p/
+ICV6YntSjNIRQvt5PCiPg+fngBNp2K49G4HC1l5rtRPwvqWlwD1c4iP6mt7Y6hq
UDx/UgEsetNRWaHyb5MKd+IlCV4QP9yVb1Wh40C8f4tCkB+b4TWYvXLgaK/Baw7N
qWga7fdA9fyFXK6h8Po8CDpk8BCTnJEkpmsJLV1kwzgtGL5Vk+w5D034mp5Vck+7
zYPlfLxe5aTQ5Zh2fQJ8/8frzoIj8OeED+H5CPUSEL6TZ7ZdNlK2lu4HD29pFDwU
+W2YRdqeH9tELHxDQbnvJqG1BNvSGk1Y7TrK4MNMweSWSpmZfyWqv+OlLrggGN3H
49hrgO5cVVXf+ZXCV1kI+5pqXMJrfN/Hlvkt+2OkpnMGC9U72WH9TqA+B3sIC9K8
s30ZHjjsBXUKNZOjXgVydK9+vaEy9IcY0M5anO8YwfND3owEneiTR0Pt20KS7LXf
tyELzPPWM9NkR2TSeZYEz+2/gl/ndHvl7REqqBG75ThSsjaBFGlZHcUsqbyIrQ+w
LWhvSl48EHfOd5u3JKas4rvsZawu/y5Iozasy7okOubgq75XyeCWHnDkoVv36GUs
7NwQhuKslbUk0cwYhFbOVRPxRbq0hFCRfjfscPTn1WX9kTkMQVa46eiCrDnDuuHS
qXk3xltW7W7LUozPxIhp3INI0bf2W9t+EqYjp6XXpV9dTDJvOOYrxXZzccE2hmhT
nvxGJIWEHmpRfkGlYA3c+Wd2et28ix/OOwNsCTeHe4M/2l2jw/pEktAlNAUPTFBI
XNJaPaZjD5WabIGChcyqZ8XtCMcXUqAxEj6jASWtvT3VLVuvb+uvojVoUHXlf2fH
5vPwLtwJVFT4PCkDE9SfzEBIWRx7QrDqBvnctMMjstFrwTxx3aYO8VaJan1SIJRB
7d/7lYu+2Ul4oxtHmRI/4r/iamjhGUcwJMxxhmdmcwsYpO/mZEe2mXef9o6wyiik
ZmUMU5QR1ja6kThEc575IJnZUcBiKGwUJXnH7mRJxyD8mmaVTIOjF24PmT8ZhKVx
i12mOAJMKEKKHWiPUkeD+qaPRi6hKIWXiVwsf9YAzcOJYKPB9itZKQtu5LhzwqSd
ZsTP/do4oUNQ6lwKPGoYm/SoXgz1NgUAE7FBY9qSVMlqX8/XJEpD/d79ygPzj3C8
nwjngBV9jLO+CrEzsRkQJEaHbN3WKROVZ8NlC6ovIu5gPqIkTNzeaHzceJONpMay
lpVY980M/pUy/oo54+S8zYOBH0NUBMniJOdEGfg2PiNTGo7w+jQuIM2egFrvwKzZ
TczHA+GOOFzl2yTSqIXs491BBrRYfaNTJJn/XIxfEitiWt4SXSvo7Ie5itdCwSeM
GRfyyJgx+b2EQoUxa6UBnbQG+gbmmvxim9jtXl422rlohYZTFGIOip0f7Bxw4ywa
lWsvx7XggkENu+akSqdhhFEkZ6/ZsEn5TeOW/MKnaF5fNb4fziUhYC1k/OCoN1nV
Q+amc867jizWc1v6IE3ngk6eEPXRpwxk/MQvUO4HXGJFJUEd+VJlwzOUBFfVIb3N
jqBo2csRBp/jLw+0KRpcJHVC8T/s0t5XrsDe69I4lpi8NLJt2d9nEsPi1kEfpKhT
Yakkju94yB3/TMtP3+pD4OQLM2HSwsMLaEkYg3dSiobUhmG9PnA/S6M8B+tm6Dhg
PRdqx63gMnzpXglDQqCqrJO7UJ6FCoGM8uA+3kLk8MZ7zK8TERHdd3Lobhazc+18
0QElIEjFHONgsZMFfIbzxw3gZKajvh2WYEym8r9RyysrNbntcf3rxlqfSwGrtJww
3zqkelStRQj83U1LOewnZTGK8CuBvYbr39YtznRxMNrcMKVmhrzwQ9dSSbCL/87o
VL7yC3k6Nv9Y6YQ4ugqWF/7QKKwjBpT3EGBxngzrgZ/kTbhbuM8Sb1+lqIKBcdI0
/SGpJPElZnF1ocjQus8eBM9ta+lnkec5CluK5NewD/bruGbDafY+06SYuRSetmho
RzuGB3zq6BitGVSJ7M4xiFfwm9rdB0+/4ZG3NMFvCaXiwTGcJ9u5P4UUuDExXsjm
4LKj6zKif8Zp2YG4PVvHcd2xOuD9ffy9vrBCjb6afwcPZsU52okazQqcu2qYxsJJ
lh4iEjLD5+UyEdMZfe+jbORsTS6SWRT6RC7d0yyUmvDfeREyJyD3Hwhbzolihq/u
+Bc9y2HpKhE+WVojxAr7Vj9nemnbc9JJDF1bLecIJ/giVMiNQgCSRq6BtWg/P6JK
Ky/WgsP270QLhDftNsKLL0vP/LOVzswOwLesQQlK1Op5oo2O64S6Ah1OGUwEidch
IPCRQ5bZ85fjAZyezOZ86CYlAxUz9MbXn29xLUB+6oyhfy9z97dVNOQxzQKCmPNA
2ax9iYxolpOa5+7FVy+WeJhmmhzSpbLr+cxNxn+5G1WX6ELNPXnRd1qJlH7s53r4
e1UN7kepb54aru0mTStQPqBhtgFWivLVIzNw0RSUb+UOJIijbVusa2c3/WJDbZ1/
G9mOlRqORFZfUtzkTV5tGxIg5X7VjIkqUtPZNw8v13km1Fkqw+bWxEnGezt5mj22
IUftLaGnS3AgURUsAHWcNWP85AW9W+JHXC7S+IOtUxmva2Ar9CRXA+JdJHTH8dOd
Etyf9dNTve6FR5/w+azVx6JlQGcg0+U5PENn055NdIjXlmO+tqDqz+SVGw3lhERC
iImYxGBNBGjpyzWlNDJKZOUDmidXVIhdJHD7dvzdWrHUeEXI0cYaYPo455CawF8+
8IOwTpmRfI+Hk4Z1IDCyJh7EJge4WexzsJfywiRKPK4xfbVZf8u25y1g45DPQFRu
HEEDW7k4yAN8AGgU//Goj27tJ6BUNQJWUYRbO9JecjsfkyzgwAbARg/tdDUZpDpG
yaI6cc3vOQj5ZguWrCOKea+srJfoEfowAu5IbqIrx+Fs6GB2dKAwHof63Lex0VWF
xt3mqcPoDg7hjlyNEQHHbUngBG8T58XRO71HuKv+Ymb0dFOEFMVvHnrCG3Sm9ksD
VD6crSg3hOFcmp6P6YSIBlfPaLlXqnyk/nE7t1zGYXuDTFm3NfX2SNWgVvtmMfXO
KbeEXuWaqW0yWbNEpDs9fIeWQyEIUbS3vujyxdxE3W1paFqhS3houIia70eCRTNo
gXneYSJomJ4NvJXbZqOn/WMzUdn4uLhiPeYoJcIs4ttEU4M3seoTsAv3zQyXQ3UV
WbZEOnhUWSkIb4p1//aGSTOp/ZBJ9VNttNc9DHXtXDdSgNyWx45spKXHrcIV+BmZ
IHu4XeOxvqpNb4NPopOPOb0oBXTWfoFDMjovtEwhPKa0fXeVBC8NhZjmMKJL+NJa
w9RjQ+T/2z+vMiNkXyxy85hh2O2iLN3qL1CF9N9Js13knFu5S5UDzYkq/vKVJ3Ku
ehYj5pMYNkC/8/wjXKzYmCQYHLvlg6WRYrHt+QfQ9KdK2XwevKbsL+0LRMeGP39k
k/GrJH71ivss8bkkdal8JeSbry6obRyJ0S4OIvXytvE17v9Iqfpqu6OYPpZyK9z8
P5UQfmODdpC7rWNgZkBOCyVhzrhorLtuC1N4IZifb2NXG9JjuCR6QEzkZ9CL2KTX
nwhcsAdsW4ikAg+0HIPb0wXH4Ky6pbboTk3iEG/9AQWRNz9mxE2ODAcBPpP9cgPL
0fS3OO7LgNVCAsKJCRGMAonZ2F5yxKa6tyO5mJxVHNXXojxqGVRpkkFEiZte3XiR
pRoB8UIORxZ+OzoZgN50BwmL/aboVOYFM6xKsmF4kj+Jkf2BmQk9Ww9pSUYzswO0
ihEBF6VkD3WmbMha7cBKpFx+U1eY8ZbTm9rIHdwzpqv1qIOP7BnJZbBb9YVVyIaf
oi9aTD8U6lIFRNtMNL8zUgqLoPbBIXSekM7MosLuLUfbYVm+1gHHzSbnFTICQuRK
phLkZp8LRqZm1hjYkV3bLDI/OVCHc9TPDGe3UJjAyFQiJ7OywCR565LPSzpu992m
R84nzvEZ/etjOxHIy6yVAGW69+mq3aLlbhsZ25/pkMQWdPLKqjOs4TwEW0uIcwHx
qp9IXVzUHUiopnthE+oTVd1HlLyN1Q8BAORG8baSgVzs/BSpiEQ9DDor6aO4tEjj
TYq3IcaD6lROK05vQtcADTxt2J8vsUYO7waYVkp/z4SgxrLuO/Fcvm23Ndt1FoUk
sZpDgSMip2XA/zCBMm94pGz6eVXq0FAXiDiKB4NmYTAlfz6wb+byM4TMfjegMh5r
vepRxhXPRplP+cLUV/PJdPGxlU2PrTKBsylXjpkHcxlSZzWRaWE0Yc3VqU0CYXOG
Bj5j0ULopZwRGCZ0DuID4fzXtz2dIfW1j3qUWXuqFI96pUBo/RiXtGmnwRgKgff9
u5/BHgp1/g+GoHJHGREtWxlBF7YyIlinjLoO0Pcvxj/sKIZZrnLE+uWya7xjBd2F
sgaAOPw/pdGtx/AEh9VwdNfBn5TlhO05GNgpn3cvYLNUoGXW0iFak4LYdxzb/6dj
EAqFoEPZoHw87WhnDAop+CKHh8TExHbt8k2Pfixue2CZdtbcFlU/c26o8HZPocSq
UF0NE8KDai/q1aNPNY0pYK8EpWygBGhAo7IxeMQfMrXDjEIdcWwQO8o0PH9PVoKy
DcutJGMYOdQpg8toGRWszybr8XtZxCFFvFyhLKfQgFy1DZnoMoUSIIskRX0pZfGl
AOWuCDUXGhva6Bos5nuFoQWcVjdHchhRRy2mG8WZeTo8OTeIR8YI9i9C2V2axFmu
YgP1Iq3zdNQEUuZisYOFmM5cTI3jPP4vVd0StmEozyVPUTm6Y9tvCPRN/ElGWaRD
30UwEvh6VO6PpzKjwR1gzeIxRDOtBWge68ocoNII8d1X1ecGkFalMnrug31aK5GM
rinN2M1T7tPx24WE3LiAeHnRm1+9csjkM8kpTe6a60sucsaYP+j9RYjQFU7wkv4+
XchVZFGJUHF1n+yJo75ztP0aQsLxNX1Exygc1TGd89oEBOyv5/5IBqyGdxUk6bYD
Fwssek5yJ5ZNa0Gwm6E4RwRTP63upFJ8PYSRXMi606BG3v2oAxuhIxAwx6hvCYMJ
r61lRO9QMOpBPwghltaAdg36LYdDCo5aexZAAql9cwmXkcOvm7SqEv5bWF3T7/L1
uwf7cSVH+JRCXaCKJTtOVIvgPfwdVWC9EzUesJvqLa3oukr91gAsmYMQRmZpjFMY
mpfry1RDGhFHh/i0QaAkOEA+C4gcqzfA/WMszvZE/qz43hoqkttfZ79kWgAtz9lb
2A29qtFoMQC/Yzy+eQShkA9IWJjtEpWM4bO0V9OZ31PWLPHR3Kb0d7vOhNNRfLDz
z9yU75JSqLHcoqTPOxRKIt2QhSicyRcpEVMtUR0JTmm+5ybQJ1V+4wh/v8ZGyX90
vlHEQ4cO2GHXaM3v+zOtUTa6jC9/BBkwH8PWj+O1LYPBWvWbLzt5r8uqnAQh10m+
g7dAgLhq6w1+gWXhySHQ+X30WPDMvMdVB/PQTKjuy+MthdHi+NnbUVuh4TF4ov8Z
xM/PxdeOhRDrsnBnd4kxHNAJ+NjE4cOKLHn13wghQuU64ijJXfTjTQjd5UvcC0OU
SQoX+dqL87SAbUHsz7Vrl95Lv/+QcwShhfhxyhr0eA5FgD2s/eCN4UqWmGvoKJL+
7kSdgzPh23SawBxd0lEwkh0L1AOy+yttsuAYlzm6JGZ6iujiyRgc84fpBtJGWmrt
EgZ7PniGfyR2kh6VOKj3ZbcCNfgqTIlKXN6WbDTV9hKHGF9y0x0ekYoCPa5iEPjD
XAPV/XGShpzyzZxrnTPoGsc6C++oJlLOR00wsIYQYDqgjy+ssCUETD0L7w5MJr3o
9sBfAcwzi1VGSVkxFddEQhB6u5QxN4ga8Wv1y7WS/LSQL0srN0Cvh6V1kaI971fE
QfZgEC2xtdhkTIuj1tyxMwJ0gN8FU+OkhD9IN2HlYtK3/QEoPxVoq3M3pQ44vkUk
jjnSIACD5D5H8vRtuBBHrdEOcL8JCr7sBdW0QE0UdVdQ9hOO1UBj15sko01AXlkc
XZg9qVCaIX2bi1KBOiT8O5my5bKJZ3G4McC8vKA2QCsIFqrHbV5ahKfHNJ+SFz0x
xBa1o/CWDvcx3Zdv5P86cv3S83x8MKoAfMQrB8YhDv3YMbWqXFIpzjoHNER+2SqS
LZZEZ8f9dueZ/eF7b+lQ+gK1SQIQVgEcN6hRMo/7AZtoap7i+IqyL3A1HGl5t+Gs
pkF2NTSchzOhDaR5z6GJQ50SZQEyLQxEzJoC4rwn8ryFUI/fHc+4H1vHv3RZxdvo
tGGQm0J4X1SVTDBu0Zp8rfSegW2Y3Bv630pUgRPCLNmPb/ywseEj2UX2iHHBJrTs
w+y0BiMWstqMJKR1/JqH7ZVIiv6SPlXsDLGI1/QSivpIZEr4JCWQ3uVdIbh6VY6Y
83ojRC5CQzrLd6gXIGBqxqREB9Z2p65oM9Po4ev80qIzcHEYIp3vfgab5UjOaI81
2zTN/YF2o9dwUY8NTOP+EKL5cJAq94g9IezqKIhRCQBOFRwMEguohpoN7r2JCvIJ
kJgdKaetzPUJt7MLUmSRV9MC1vVwoaDSyN4VQNNFXmVceUr8RECmqHqwI6HxskI8
U3Rq26MQWT0Z8ALmcI/IRNyp8mEwjRHLzBaxPz3mDN8Omu2kN+rphdEMrFFaNbkv
p1V6FfhC8JcdMdmyRopi8IO2mMMf5teqnznzJDH+1g7LJL4sTbWBM14mXJQtg7Uh
53qpp0foaaa6w+zt6Bdk72058IejyjGJhdNsFoB0WUqK62MXJvzYfIDxZz5NfgUV
aFUJLGCDiO0+BF8xiwTQLVhpCPCQtx3hGn+G/uGOffzIyHa/QU6oWY6G5tqJR29j
cJTX/2Iq1drcudxxadUyOqGNWEJkzcdl40pD2GfjuS4kuZcUV5yHahCo+djErvJW
7TNNHRZ7y55I5K55Ktx/W6H6rxZczr22hE8NTl7H1pkTomKbdhSBkvfdcfYxhbCd
U8m1GHI0B4eD3CCG0ASsor1J7AEYHU7MmAh62ui+yLxu51roVnhmv1sgFTPnYntG
u9/tEF/6KKbNJ5q77VO7NkMqZVI40BocR8bLuqv9RC4CYT/DnDx6NCkJEErCcHhd
qLDJX67aJ94N69McgU/aQ1vhyKdQGgwrAunnU7TMPdI8CxDxpKbICojGg5mNJ1xG
tKg61FqPJHlN09N5nnf6caRe5ohW+XiToDQq4uUDYz4x6C1V9o+jsDE2DJnErGUR
FhwpmoYCF+yezGvpEQ2eCax6QP2MvL1T6fwQjzC7V8Rt8fJhkYPO9/vXKNXfuVLB
/NdcUSkkabnL+bfYNvsFiKQ9VUjdWJFpRx/Ikliqtkiw7CSCE/HUXH3H5iLMZAJ6
uGfP1SPjCR32q/FX4Zt5U/DOk3SeP8UHgpyp3MCEt3BUNZT4JpSNxZqB8nF+ahJG
gwgoSbADOHLAhM5ub4fQQlCg7m2V9kzs+bpqhCaBH7ulRYZJBDLBDyWG+YNb7YpA
NLoY6Rw6U3ehfKcrJ4j4W7iLKGF+kgM1zhP6mDcGBtvP4LJD14DA2mJWNoQVblwQ
p6w/vzTCkIKwe49e3QY4ltoPHKq2isaKeg1/Mx9GpT/0uH9ZfzNj4oUv64HHBD6K
ceJnfQ5L8EOPN64zzH/E/C6r6RVHU4Hq0vqed9kcoPKj5w7FihaIyfzUM7R4PC8z
9TCfrp1ZDL6W9WJLeZDkYTx5rd+M5OnjWE5NYaeJ8+YyXH1ixBWBHxPGo8mRaVvB
S7ysBjZE+otQ5n0ZfWLAdD/7gTwocPMh/DdRtqp2X2Mff1UrgOGXcCwt2FBUyHIx
RBD1NDBNrPMtejWsi/5/N1YY0VXBGapaW8N3+BQr7TkOpZ4qhsR0zbrnpZx3wFup
zuJEgmtY3GriaZ7bFGNv4994bJfgiaJS1kNSPSU284p2nLxDOH4lsduQ8ZgnK29r
oyEetu3VjE4+VkaEgrODztlcVnikcQxb+8q/9s2H3h8jw+gNk3ZMqXvzDKTQFedi
UGaEiPQL1pFR6i3tLBshFdgw0hKdlgNzW3TPDCfP3Tz96iK40MTzdVtnH+8gvnU9
JM59HxfzHTZD/XuC6+cVA+1eXq5v4up7ELSF0Af4uKXJChZqPzEr3jcS0dhOuNeP
HQRUrsNbixyelHOG3RDm98QIwNnhz6VwQag9Wfyr8D1AHK8jkLcfs3A3fSZf2t2K
2RQG7b5YOK3Bh+fXAjSJtDFNBrN+2JYKCTWxNz1i4IlVgHqbWwIWKgR6g4C2K5sd
I64GT5MWIP2f4OzqjROkFnrnWQn1dIly6RxVA95Ab+s/VLuJDj41cH3stuWKAfK9
ZRoeWIOavga6NdvVGq74N87KXMp2LJE+4LJ+HGZq+B7q4XJ0IaTjHlXetdyKWTCa
OcGnllvMpIT5CcqpinAdopXmx9VmGGzqHqCK/EjiYDnwS05Y9R3W3gLHJAQV028q
6W+1xhWCN06YxSal5kIMRjQE2DqQC74oV4fcAeyZxAVLfNlCglm9OL0GvYrfFGNc
NGtxme+6n1DNpCAKjdJxYUlPCZaDIuFRJFf0JBNJ2C48wcIRGNfMR/WrdWtFxhXa
7SXouJi55vo/xI4jnlaUCG70hiJW+1HyCCCDvd7+Z4hiSl62o2enHMROMmVsfdlm
AjUOfIOc6KMA2aLRzuJPY4C3nk2gbuf4m680p2dyXbp3QW+5m/4o52dSnlHaaXS4
6yaGKZnAAWzHW/G3vB1FhyY04uC+d4wIaKhwHxyOLXFn6s9XxcXMvjURk/2eadaZ
jg88Dgm7+fxkTmNx3ZqhLTj7mmYSoM9m7hyLcYRUgcZ1RBRcVoTABnUe13E5kYJE
ovav2k/dsOznXqiytgFJ4nqmpBjlJHqQXvRyDBl/8mCV9kM6CmpJVRfg4+em9K22
I5ITyYTf+5hcBlkFmQJNxRDu+CQWRkAFeavlIaMe9IwEEG3OCn9M49YCqbQLds39
auefa1fKPUuo+zH/oeAY2ml/ef8PaTlsdyLy80QA8UyILBkuYzOpATeZrYvAmIxj
syVvYeRYCRaBp3XszPKHQRlLnYknuLlCLXGj7w/7J1jsHLuTMB4Ibw9HeFv4CfwU
HAZIijLusjLlzkD+KYUJ3NP4aormkVDs5GSmQJDng04i6FJEhZkSWb6Hpo6Ml2rC
ppPxxKAa6p4yf9Cnv1cmjkt78mpp6+8N4DDDzu3RHnaIgto7UjoGiQHdQ9K0lNr9
8iluwJzCshvX0LFPR783kRpN3ZjF4iEPKlEhK7UicJ7gkS/KCHsdTwzi7xH2/bS4
XTmxYcfXEbmnW12+in7MMqBs6nck6Rz5Vv8sMk6/4st0Js84NWbtBr6BmASi5KwT
X3u/QUQdd2lDJMpRF9bs4UxeRQBXGj3cK1zFO5tw0euTmHdhdBgkcjmNqp2vI12p
k2A/J5BA/1nRKHoCczaeXkbglez2FApOEM8MYu+AksPIJA6iiZWV7+bIuAbks8Q8
VD2YVP4UDgUmM8VDkZbTUsTy/MnUJ/QYNgi3cLFMAhRQTxoaHQ0ad2sp2xTFtRSG
K4cQvDDvSKRyJwT7nwteGfsiOiq8DUZseOlLYZrjeNfOdRYVnIPx4yN31Caf6VvL
AWh73daNBUPuwyyd7PPbvXFVSW64sZZFQEH6TKEpdFcDDKVqcq+Cjj16iBDoEz1v
yOX169xygsP29wExYgE8ZXHC65X3VgBsx4PAkNj0MenVNmeoKvq2atu3rHgx+one
z/4mbq/XRl1k3OjBQ+KFf06SohSScd2d1b3FRCf9Ech8JJi33fBvXzb12IqPbY+L
MzTACyKpyNM3auYVMSxQo6FQX8bcGznfiW9yQtxrMCLUt3sDCmCsDXVXeyyX2fXb
jgIquGPt+nAaxEVNrtzDJIrxWgi//PPHYkzy8Qq5y5niuhC6UW6FUkV+5HqGaB5g
6DzTuLjROb4irHvxuq7/Vittlfo/wEy5TAo9j7d6I4Qmr+On8DfTHRiDrnEzcbVr
J70NwX2qCSnHykwUoaDr/L3XFPIFCsnBlPymxQf+oIZOHCbhm/Dw6XmEWcf2unOv
Od1Cbvtvn+DwV77GKCviyKsBk2liu3y4ulm4HPSN2HigPuFzLylAOM3b+jXQQN57
0ddZiQyHc7D8oLlSY0aaIqSnt0V1CGvPuMDJJBRNmzEZnTdWSER+NmCQuptQ8DHl
YNDVsh9klinDF+Uy+MwUH0SVzpREEUMoHod+b+MOCnKLF0+Z8PN4PSHMpbLcV3NW
26Y5vDSngOBKgeTAvgA5lrDoZl4zWKGpyQ9+8j+37H5RYhLUzn7WV2yCI2Ofh6b0
hXkA12nmZivtNE0SIbOn2gOx/q5SYXQFgtPuefen217tuO+TjHjoM8Qfc+qBOIzJ
OY/BFVQxZNjnff0/TUK4ZmOhRm0ki6EHgUJYmbB5rPiQ0V3LCK6ywyn51BdPKYZL
nxaD7erHtwF8iEge2Bbh3s9GTn4Yq+8SXSU+xKKe+DZZE/ZD5myRnk2EpdDwpSrT
KF1+3kp5VnGEWdLXVUQcEJFw9ve2y0MvpqRvhGYE1X/fII4YbdVSr3SnaJpSC4Ym
jgIz6Y4Bcvd0sGrs8Ax8a2anesfF82etU3Hb3NH1qW+dTnxSm/r2jxYnHae//73f
553ktz1rQx+cxOEBq4xsRjL6tyh8zKemG1TWg9/yt5fcLrZnDanJRQSU/3KBG+So
r7wFarWQ37QgT+WssWkUhlfvQX7SXofJmMWlIBfRxCK0GrmQp+GKu/6mOsu5+Fv2
7RQ/R//0IztPaHhMYvt7AFEueKV0orN/nPNvrhjSqzj7/vemtK6DXBImsRpwIwq/
1ObjnXzAU3Vj7dUvFABvbkv0oA+6/QKoPdllGoa3mLu5TfA3PS1Umn6WuHCpi9pS
otDF/1gkrzBYusUN6eGch2hgISwCmGB++0MvUcA2GvXQIkbCxtNP3YgPvRklv9iH
H7/WjBJvQvTU0tb6NprZHURRFSc4d4S07aMw/uHSL6y4yfeIyxEZgw5NbpbpbVBB
jLvTFbZNEZkI31RFZ8E19oAsd+9WHkAmzp7r49sFQo4jFUS8JMEhxDqtg85fLXoo
eqF1hNq+FL9F6FUCfDsNDr4bxIRRzMWeTig4/Jq1QNqwC5hKggoKCqjZO9pL7lkV
jy7YbGeXeu6sfElPXsPJgr3ATx6AvkLfew55vn3ynjh8+yzdURZVpuvtl2tzI9cj
SpXuCpHj1kMNLjuLSOVMCe6zR7S3FBZ1sjrRKrIea4HcY4ecGC07yMwVUBm6PCmF
Aw8JEWPq+Vt5JBSwVKuuxKaPdQa17FpwiveLXDLHTutCevwkverwg2N43hIyFE/s
8AiDPLQIiR+BT/yb11H0xzej4LdlRgDm/U5HQU3dh1jKFzEvkPbYbLQIfnmmc5Lq
lYPftOXZmk3eAllZQL770zEriIsxA58y3wfnaUQ27Zdm3/IH+chHtbpRtwpcobdp
oSq23gf8cKA/qhmra5CP5+Hn0e41JCmb0s+gYMY+HW96YDtVSEmsZa/+XNePrxm3
fhiJunovuYYDLiD9SeJS1A/3cxeSc8t3pg5wDwI00DKV5QousfVxO8by0ejp0hJe
1kd5W3757P2nCroM29HZz/MB8xcjETJeLnXBsM+6k6HRbLCVrrAMqUKjORM9piEg
AObSvZ/nG26FTWvg+uNBFdVrwd965PJItvkbwbMcQnkNodSjJ439F5Cbap91VAB9
SxjvjsOXdctymecF9T6uyERO931h8sGccOZ7dvexwRgno1BXBqgNmmUVte8LFh2l
xoMhzJL9FVu/D6ZAfNoqAKJ66tmxmATD6eWEFV5Oy0aSzV2VRBebqPSvg+2umhgc
srpmxSND3WIJ8r62SM3IiuttPoiSMoFqJWOmkCguc+TpVWeLbAbIWbMT7omNf1/H
PdD+g8aMC80tmJ6K0Gkzx2k3jG4b1c/O9P/WM1CXBRqwIB9+Jtw5JCLWAgZQp1JD
vUkWTw2detrWoGTW5EdTel8FL7D1gagRqNDY9oN/JPnynmqPQfEm9Wdb0zMik4zp
J8DwZoA2bRjSStiFV/BzUqHbv0heS71MD8cesxzke6yqUT1Mb3dop9tzPh4XRcTN
YoDQmO66CGLGyUjZ/ZXw6zRw5on+LQKITCDBjT/SVQghCrslwcFHkNAfkdbJbi32
SWLRS9Qyr/g73FJLavsYT5//TjGQnjOqg24sFDbjrlyujbAyTFltQlRDAROG5r3W
Wt/OD6gYf+0rZx2PjLirFbmUnGzVatm2TC5eLagmwjQpld/ILkv1GAVpIVomI2U2
2cfQCiyg8iDtF5m9gBTKmLje7a6tsxMQQu9l2bpLRfQPMiUhXA5ll1koA9KsTgGq
+NXGOA1YMxTwOhaex2gPkp5LTK3MYuCi0x6x2pKZ3zEneDYdPSY8TJxyqCYwvsLR
m82Siop6cPcLvLo6dPNLMc7SoVnIFC5IgWr2tQmlHqjA0f/RyagSsIcHWmIpGVth
dYCsl9RG9d71LfIK9gh8l4MX/riyJ2bYH1s+FMRtnBayCwXmkNRMRpjyIkRsV7hi
H3xCOOMub3Z4I2kwukS7OKSgIeCXfzo3lpggBec3j4bOCq+3EM9K55FyRoS3i7qO
b5JzKspYU6K5kaRelU0Px1gco63nSLUJeB0Qa3mEyH1KiF96y9q55cOp2qYZ8sVv
qzyqFu0RBUXuga/vJgRO3jn9jAfwiSUBA26AqU0XwuKoaXpNmy04mvBC78pMxqzv
OaGn7iR9SYp8nvoeTu9xyB/OCXFuRFFgAhmDnmdAd7GOECzgpKts4/wDE8SteC9b
gwWwr1BvVVaAm13hzrofQtVVBzS9nX9hcxYQHmIWtwS7q2SNy2YpchBEsdqdKDBe
Tq3MzcOOh0vZOqKNzUvIRnMtIc2s1V08JfFb3JiSP5UEQpuFq53OXTLbV4yeXQA0
i0ku6G3wm9b6Biwog5Wzl2vNHTjMR9zS1Eh8Rf1L/LALAJMPUCx3mdjQSaDp1FsZ
O1L88UXEfdAQM0ajcvp54Bh+tnvRSkPu1jlTClcenmhPd1kr6o+Ks/NFTKfq6XEI
2ppvIqPGAxcSetxtqN5h/MwEgRZluzTPsegLeNDmp8h7XGIASaon0PBJRnv8ulp+
BkAh/I0/sgEpG7+6J/YV2rIjK0NhU99ipGYwnqwCDDKS9YjcHV8aOzqcuMCtgrFb
3AMg6WpYUbQyzcIhidu2pmSUpPe4i+qP34PKzPDCkxrYzqBQUckxFZiYYPnSR9SQ
ve7ZuXICLsGSwvQDpgI8/HEdrlVHdG0VJ9ZfAqIQygjpR81Iao8l+65543/komyQ
pPTDq5pdfQQM82QWeYGR1l1hab9TvwFSJZ8lmtPjljcCe0uuIMYYW4fftzIyKixT
ryIqv24uguYZ9usWitUB8X7plCPL/3gBrguLh8VcdImjlrpK1xhr1P5jhAuxYzFU
OAZ+cDhlz0ZEXD/IHf1kNEUNgkWVwqYIZQ7Sa4DSa2Hk3zDWEFqEXLuI0VUKN3T7
U407MlkuJ+LsQ2vDhpMgpdGzqeP1NIvShuTOxCeXoZoXsyq7ig0p9GgmBO45O/tR
Du5CaOq8vrj8sLSRTPF2nf2Oj5tjAbsKeUaTn2hgj3FBQM+SlKTbUcNxZ7blU3Z3
3LyfBrNodeAG56luAnNDD32GlRuik/ih91VWHf/ZRZMeoSWFRaD6Pb1bhte6jSau
Q8cxp8TbzNH09cU2i/Avrkup3A0gdLH0jygmsYsS/+kdbnGR5e3XbUu/4g3mIKA5
GNKCsMxHIQN9LI2Om13vek5D6ld2XvDXP+hQjYVkeQGKXuld+xUH4e706sNrXKuw
qiUMXjLtunQMe/ba+gAkLrvsPlAAWL3be9rkE8DfK/LOkk1PVTbXjLhiX14c9QBG
bkC0s9GMFoRP0RYDr5sFGhh8TcVHC5CSE64Uig0O+j9hKZdoO14RvWB5obmcKJKi
rQjaltdQNeBFE6hbiTnTYHQX9vJmf2c2Xrpco4XATyvq8mm5Vpo/z2+CDyJkotF8
0fmCBsZVzWPGDbABr5PDOFSkH874JkJTo3c6+QMZgzHV2n6ol67ALe5GYL2fOdHg
/QoaolRx8iqXeguPXIaPUKNmbqpCpWL9eUkeMcyDXJcg/0qRcG9+OfAuM/85cdMO
GABkxNwbR9Es0nV4EmRIy5Kzq2TxJyjCvQdRio7yOYsPdHOcG8tbHbPmdHjBp69c
Pu92zK8SP9inUBzRtYtBZxLOG1Zy7Mn1EPJ5469jT1CgkJQouC1WnaTdc01DQjwS
FyW9NJMFTiZOi6CGEX6T/MDRVnd9iFHhh2qKjvIprxepjGMCy0XW60M1LEKKIp6r
yG2QycG6n9ud0iIJTD5F0Nxq89RYp3DPnQSU5rFbwMETZsrFZx74rbZ0kx5lAl0W
xSnMHteTu8NaBFIkoQRGm4dD6V/ul6+jXy0AWHgq046JdL8h4UqHEa1fWpUVvlAr
6kdvOlGdt3bq1P92J8ycT8+YSEAwZElaDn9f5u8Eol5idT0HciYts5ojN3Cbnwou
iLrCiVQnrtX8hB1fBWj5cOXB6MpMzuLP9YTY9UNEoz06yYTFxmKvAWk6B1R0xQ2I
b9T+JH6BmfgXBvZSYLHEFlkUJzM45eOOikUgJKd4f0I0BNfVl9KmuAmI3S1RFslt
v491RcnYf2M+xxjZYYJSjIY0CQvH7Nro9NwQt4IPOx1O9FYidFxXbQX1x14m24nn
25JmZEvsxfjLiRXYNIVobLVw4FfB3qO1y25S2Iiu8ZHih9dIEcVWk59lzZOl9k6z
dFpYF60w+9jdFqGXdnugbU5056ACTZif6SOlcxKrlYRS+nHaHqGETbgaOraCAfH2
3bFgavJ6EKrmQplo0QX/qC3IWONYP8DZAjUxbvdbESoa7h3PTF4Yt1A2HWIDEcF1
P2U6dksheGcVdJAJzeiQX7aKMP2Z119mCz6SH+Cyjhz+YTJhHOnXUztP+tikDnZQ
uq8nsuBFh3rmrEzShztSTEvZIZKwHtdUDzJpx0dDQR4Jixwa0m30AIB390+g9Ryl
G8S0jwteJXtK0o9GS1I3hc9CDinkWP4148WwRL1BFT4iPKkEEhrvstLMUlC+QyQX
g3HeWf/cEvMvVPNYCEXXRb1SN3s8dpu7uJiOLntyMXpmjmOlSXJ9bQeaC60bnDRg
85qP2/lVewZjC5ubaS2QQGsVwrRBKGXPYbXWLptIYhhnbnp55/cxojt6bZBGObad
ATb3ZqLAQCewjpfWzyLDRQUXkJDTg+zchGIF5G4XEICdLLrQlHfFotH83o289l21
cNu/WnNC/IWdBir+Du8rSkMPTzsLIMWHYBMazVdoS20Ao7eHXu+8X6BIYIoc/kEd
qFA7lQJNQ+7EujZ6xl1qxJj6relYcOiSX2uUc+Jg8H6d0vVfhXy2vPyD6gZxS2Kl
BVXNetwyEDKcNy2V6DCqU715Nrmc2tAgvcBd8asIpS4p1ZZPjfWYxTxjYexKrMDE
58P3PtP+qoMYLLXDocRUcWZLuOtrVkopbqk3kb1eGvZ2TRfjWqxYXb3ta4JZuOnQ
/U7C1pd93IsrAK/FxHgKnP0lkttoFtdAuwzxAj8fmBeLI9C2zbnPSUvMJ2ATH7B0
g+xcm0o4kKydQWwXDRj6OdsQ3G8w5/ndD6+GI7HNJx+DZQhcTzz7SVPKG1NmUyOR
N5VwGyjiiLDGWe5Z07W3qOxadHd8+0NXB5ulR1LbjWDFTnB3tlf+/MTfErhjC3oN
oY/1OFd2lGZHm62Hgww896O4f1I67KwcD8O39wMw2pHeg4F5dDoLYNWL46IE2jqp
Urc8nV9JKG88SYR9XRcpbL53YsTigkQgVNVSs6vp4bmQ9XU/0pI8IF1VrjnIaprb
9JJaHlMBiKRD3+qfstCwllNUIUJSaI2P9Ct4io3dtbxTn+ttaEGKpm0tPd0iPlHc
EF5StEUKmmTN2Fn9suJHE3LxGVfgmPs2Z9gQqXwHhDHGnX0PpynnAgoE15OdV1v0
ZiG/7wJUf2jB2fzOuk5pSOJqRC57DZRYewl8jMYbvIFFlV5N7kpkxWDJ6yWbYNT6
IjDfPIrPUEukEBYwew/pdW7Lw03KxCy6JO8x3lGpF5oXooFZ9HoQK3Ic/+o9Q2gt
zK46/38oYyoj2I9meAsg+y1819Vxillpx7SWWZIpTQr5pmJk+3/XeYdOogehB7ec
wzMNAgh9k5mETBQzGccOuA+kcYbk/VDp3asCu3po5/kToC43dTAxHsXSZPS/A1RK
ALVbcFkbbEybjRVT/Mnlj6KLkFutLOmuE8z3l80J3HhfWkyU1HEXbJnySfWduB3X
/yv0kgP70zML3FterFlGYcnBfto1TSvGq2zaCeBSKWciFbNL2cjnJZLOP5M3Vgqv
92BBZcO52+gdkjtbuR5X4ZXZ3luyo4UR0fE5KerFKnNMl0UZgnrOJwVJliDFjheg
vLIx5I6IVUoQaEopqY81oWcKfBwNru2Z5jUbH7THad8Lq9oMbFehl9j9HcugAY2k
0w43DtTRAoBj7woyNsdjjoGsPHHkj0O43VxvodSiPeKSoozQ5W8/aVQ1za319jJf
qWBswotsbPuTSnaxJSONpqw6+30uXYI7nrRkH60Abc3KImKtRaOpZf1WBU7aRoJ4
XDeuSWRxAN8kUn+xbOU2pcd8BNH6Fiz2aBl+Jctx+KA2f+gyxOzoto5iYeG/lhqN
Lgf8X+Iocsuyuj15wfCkMjb3wSQKi71drQJeDwL3MB54sKog8hrDaC5XZeFfyIp8
gEHXASpRubzmUIoNq01YL9oeeu752TQoj/6cyKqBoCp+RKsa3hUiXlGXA6kHQHiw
mXlammdPiHj63rwWhTS5MhRJNT1p4H9WMk2GIr7BaCsOHggzV3y2D5bhZmNrm4/q
AkfHP2s8CUPH6sQC6v2CCMVvyArXMFz0iwUn4C6wA88ERnk11kJkKKoKv5lnV06u
bWcT2vZupiSV7i/okz/rfnjILT3p2CIzDcxbcH516slFR2VH/Rg+Yykc4hIFrzCB
JQBBemC+DgsQ/FQxBDiXKMG85kMMzWeMIkLuS+3BoELplVCfJvKOfTWJka8V6KcV
4dL0IoiCQdRfMze1j8zZNjZzhyRvWxziCJPiq8Mp3xdcKeZJCf08CN2mpQ9FJMny
N+4DO09W93qzi8XhQjiq2817tTUo8x1ohA4vzepfRioqkb4X2mKpU17LG5EXJGvq
alWzQ/wlkxedZb8hZPtQiJjsHLiUma9xtZ2D1HPkO+KXW9BuSh5GMX++WMkItt0Q
0Uh3ANqCfkPF+l2QWe1a9HdrEyd/hgWoDIBuvmoWCAKTt3P91PFRGfgRC7duwQU1
l8uiVa08jXIc4J4J5T558TjfqafxPlj38k4RMKTaxVtRrr4zkJvPkIuyh8FQehaH
ry2Gg9tVblQXCtyyoZga/ZyO71FoUPm7aIOTYBosjIL861f3XejOHC0wgFqAmTgc
rimQSTxqjlvI9CpEtdB+F3hd47wDZDNGTfJ2rHm0Idh/uQTAHWgox2nEXHNQUndU
kI+cc8iqr+l8Dei4bGFHYTTrPWTfNA/lTzwy3HYgBjqKC2g/MVsJzxWWt4YKpIHd
+0AGl60TXLp6RAphzT8HH5tAQFMxwyHz9AQwoH9X7CArpjl6yfBwELYb8EWJNIu+
V41DCkG6BIdnqh5b2xxe773Y8TyJyc1D4XxRmjurmWBsCDbfk42SuJCv0svdiO8J
IDhb4wIH6pAxoT/zH2L6wbHL84nTRS6zTvk3ZZfLOYAigXFMxzDlNlNVdITmC3o6
SEL8VCsYoswBHEvIeHrQ2Fn+1GgBzC6Q+os8scAIBZRTUoxd2bZLXvgL8nqSaiE2
sMpeDnPprNVIyA+87LLfhQjMT4vwrpc6iHRmgREmhmJVWM026Kp1adr1TbTozLUX
yBid9u4MYsEl610llqxBtJu1K/JoYAryXtr226WMT9k+JaJqBKUsBBuQjQgXJ6bW
X1sApDq5dnMSZMCpMoY58LJtv3ogKK1E70/bpJnmcaBAFkRNDsSnd0BQ2J8tfIO8
gtJD0Kd2huv4uIQ8ZWhAPwjN71bEDtw6STyruzborJ4eHDKFxIvxjOt7OCa0prXo
vMFyDJA7fFTbOeC1GKtUhRis/tU9rkYJ5mKAVV0dVLyK9wkc02L7UNM7/OZUri3R
rY/VmJ+Wc4bn4NaLN9w1StZNgNu7NvzcAVcbIzd57qjH35Vmncgh54WrKlSRjVe7
QcyhKMZ2B8S+xexY78gbqLkNfv7aexjxjRnoLXn2xylT+/uwpu0qROhZgBn5QLge
lA9lJNy4UkmhcZPIgPNWN8hcEDWmc0w5wjIJPdIcoWQ09UbjgkTD5WMwz1Mu6vTw
dCItkpNQLYOSKI3e2HbtycnyL8ZUMxFYClNLqsWDojIJOGs5JrE/hiitvgTfCiDA
p6TF6eHRqg3ytBXIBMkUF61q+NbKLs2/o+pqSPgI/yw59PMtlVsVYjo46+NIEWCO
/JGaJjiz1+XGG3uz/J6iQscz7pYvD7Fs/LbZOtDQGVN5r2Ot4u8NDKtfJ8tCfFGy
bbQvXFNKokemsPZ6F6VXFi8loCBeW3cAFNJ34QuGMx7yq9kxtJ+ie0LunAZOcLMq
qEnckBBA9DM2+SUTdx2gtriBmoGIk25Gs29zMg1B4Za8TqjVi85ZMj0N8P9pbfKP
lK/fET4taCVqAn8WgXBqPYJx1ZV/2JPIGavktUnZZRn/a12Wi7qh0YHY/lUYKxSx
obsuX1IpY6tNAWc3xWJTzCtrAgizOmrvNyzjJlqqy4heNes/NNJUHH6zWbovDr/o
J8dlommD3YQ+U+7FwJvNyyXP9V+iXdGZlOX9Sd5GvKy2SAv5abmqCzQ4pKS+o0Ci
JMQ+qmifed6QFIGEjQjoqKzb4QVEtfecwIRgquMJAjjF/Tch+P+0IUrLsrfDghwv
xOMWJa5JGNHFAXYvY8Sua1QV4+xVKMvTIAeXqKTswtMxFAwL2WvjrCE/zJFqeZM0
XCc/ouRuJfzi1JvRwuRWs0l78xQs6eRsWhYaDTBVlYfdToVvI3FPZPeJPflddMRA
ES1uZRnjpZwtzMsm2kRUTpQ/e4k0sNHEkNKZLmtVqkEJYBXeCiJtOiW8EKQouqdd
UpnI0HD/fsk+7hq9m9m1ZRB2hy5PkzJrB0VbP+UU6aDbow4JjNnVWItAbvvwY+zn
GMxOzGS4n+McXAvfJczwpIV19PFAPcA9ddVmMUkxfJDTRn8oIbA2rtQRp/QqOYeu
eJ481dF73ur6JDJxj5gbK68kktBkl9OPlqcgOE3AJhwOKvlpi89YZHORVX9G8+tl
BPvIJ00do/y1QULebXQ5eTYJTzDRKqCyzseF89201H67+Vmw/3Dyi8wwXmjs2muM
R3ZOuk6NMxbqtPdufH4xOt3QOIAH1rfiCs6z1GR5I9RelmMWi2PL9HUdXJVr5y1b
DNW7lO523tBgP+YUSOqcD7pD2M1XI6kQ+G9cX0jVeBbuYRz4xUVqLZ2FsduX0ZP4
5d8XONd6CLFB3CTHKf6iuK1OpO69gYJVPiIYiEnsjUAZp1J8dEPxxwHFbc6XQSyp
2xRpMpIUQLURronOxFa8Hgi1u/cfowRf6v2yWRtlSbDTVqh3mlg880a69fqxiI0m
3bPrgJ5iYlz422DDgpzvcdsBF9tM4ACp50wuLO+Q0Z67QTDbMhVnS1n9W5knlqQt
5D8pEtAcBM+KXiSJS2WSpK+A3CtwcgYiTw9ucyR3tVFiTenr94tw8E/1zPiChMYX
zEZ3AHUK4m61r7B2LhM5Txh3qg5hATIdaQCp5wqjY+04YmWpEje16eV0RjDxDV6H
lTag9i5o9cGgInDV/EI68h/auf0Lay8gaejtbuvMmrtWFoRuK82uzYxTwb0esm/L
z2ctvJj8CM5WhwtfIf9dsuT3Wg0l+4uTNafUvkzVeSOfvca70kJiigIPWxc6JwtB
CmSnrlbH26OdrCLLCRQ7jVcawwwzyOZE2mAomb8sv/X0BzYRYANqfbSsWxrvdgxO
zWe2JVD8KskcO7yd3a0uy6IryQcJHUJ52lr2/GrIHm4t3MdcTDuLok1iB6BOLNJm
W/5GZIWTHHwj77TdjiUdB9qdVTyKr2JSr8L3QO5oC4oyuUQCDl5iD6OCJm4Swcy8
Q7h4bg2EmxQLYqGdZDRAPZuwEhlntOgqEclhxyUHfG2EmZbjbvf5V9S8LPqCNh2C
5cK26XfA/krEdqrwC80CP5pmbUcG8TM4p+U4MNFnVBzNnwGQcG1O6Rm+rytcti5k
0TZk9e+Xitv39PP4Upk590p892GBzEluepqBssSkvceURSClqUNZz9tE64h/HoUU
NF2Do8vf6N2vkuo/o9OEfVPVn1LCboZOJmtI6yMu2zy1TIkdqClMLY8tlgYMWqqs
m7mo2m3BotvKbcvs8MKy1fxX5C6EZV3GQRGtMyPlV5DziL1wIcunRrMOx6CEX+ja
Wr3LP4+OdZ3kJUgK/81i19/QLfIm+lmmuJ+UC+PiKhQ46BYNAM7FLjO96RTHrrvy
PYI8xrxcfAuVZmYZpZja9mjlssVv6inFMijYDuSu/UXXmFOKwQ7q3s0ML7sq6jJJ
7rnrgLoNQ3PVGiYf5V67LRA3wb4GZXhB6gxBpJGhU9FrjUL4GR2L7SYyF08bVXkh
GVB6br/lAbHJXNnbymcARwgt0oLGrIvGCtPKOyOxULh54UWw9fQ1LC/kANj5jCka
m7EOONKjJaq9sEFaip8cjWJLNYbr9DrfDSD4dK7958smf+iMTxnzJvA2feQ0/03y
76LvPfvSGgExxobohoc92yo23iI3w+NcrT8ZhKPWK3oaCueBcBPkZfzc9zWvEwqs
ErkifAMJXWdoQODXbsb/77FB9whmqEqXNr4BSHb/iMjxjGw6D8JqOpH3e0k94vot
Io71kGMv+W0dedsQt8uPWZksYCBIHEY6qWQHsQh5PsX+IHLSHLT/Is1XBQuy5rBv
zf8BpHFFVZLMvvcshwWpyAUxo1WcrAZG/9Y74SaVwG5dw37ji3VbITNLbtw/+L+W
hQO8yv0WS8WBwEx8wKAibLdKfzyoV10LIgDEZVRRDsRF8nhJ4NhEqXdja9iCJiSQ
WAks9OcKFTk8fcUxCDGyrf/qbTZIbvUb4qBJuklE2oO5EBDgieoN3ewsDcl2fjOC
M2g8t+g/GmE9RURw5DQLo+eDrukhGmWb1GfVrfC4CsbuBHWtZq+QcehnzRNs0pu5
37PZ1xvfFLfOAf03n8YcbnnTKOlPvBxtu0fl6rbmiLzPPVT/21KK4v2w1s0YJ98X
VsrOwFafxfIfdRsODMc78sM89ZZKdSOXVvTYHxEx2P53xvVttyXKxqu6Vr3NWisg
ctP87/45JTjED2kj82CPTTTQBc3BvS82iDyCjFOTC143cuOUdJ+jEG7gUJeG8yfO
ZhMvwxH51NzPm70ZiUPgHPoNV3D3pk17k2HSGIxUvz0OFIWn5fG8kVeWm1MlCXg4
8AoYvp4bmifiEoHH+i4yiRoF+ni4pBjXxYvuvAv4rhJTODQ0jg0bni4hpX9hrJ6N
fyDRZTcBgqImqiR7AK87oqZNbUVfphq+wuPOlpRoUbq/UgCmWvfFH8AFJvRSlAhV
HScRUlU2JdYOW7bJ1C+0s1/89CGmnIlAh/IH7hIUfsdRj/PUnOdJxFJIPURkO8fG
uDuvkv0flJUfnky0jbL2kcnpCF4Vb5NRkuxssZ6o1ROa99E5WDTtXF1pHUqKj8sz
DhKVx4qoBiaa3OOqZhUwil9mTRmhHQIlIZvYa7RppOsx1ceU/laaOSmuWOwpQty+
wb0ehAddCYbghffQviT7FU8Srlzsr43LiRqyoh2x6ErbHA0CtNC5KStO2FiAY9Jh
ZcyAp2MhAgmv3Tk965d2Vq/lngA87MIJUeouy5zMWlxe3fDZ3pIVKHy5r9PyN07R
JEKi/6LuJftu53634mc4TRQd53Mcjcy/nZCMXRcaf+zWS4Tt9KefHvMXaz7C91BY
P8Bf6kliNYQZ7Uc/iXRc8m3kIBy1ZUiZsyAQEcIgi6F3uoOID1ObIIs1ZIF4Aisr
PrB+rDRN5HN0TF3D6R/LHdmK+a14R3/DG1feQr8NrHkSTHChusnyMyy8uJG2i+Zl
GxsNX1cVE5dibqWah3eVdKv7BDggW2WEnxf+yUd1L5XLrMrkThS0Ak1+LxV5Wir1
sUi7cuLj67tFTYS29t9sU5WRKaHQhtwSKlh5ckNhFeMssjsqxwLerua4T3j7uojI
+3o7JrknhRTYV74+1tA08ocO+u0TrrgJO/x8LU+9gzIf17TioWgkc2HjDQySkhoJ
CY3Y5psKcYEeqKoHCEcTven5ll7p6+jwJ9JeuXquVAQzN0bd1U2/zknIsAJ1ZseA
ce88xVc3Mby+PlYsrDZ9yWI6c2CxnugKd5A0lMOqsAKTQwYVlTXlj9nQuiu813eQ
oibp3iOD++QIeZzNcwmZH5/6LIC+vHNPKnPU/mR+9LV0OT28Hx9Qlt5RrhvSRc+I
ytqK3XNQ6gPtStPNA5neajCLktswLGKqWapNYV551IOkejly5pJRRamg9EWtuMHJ
nJtCC9lbWC4CAk77JwQ/wMa5b6wxM4+N2t34MfAKrNMsgmZaa7cfuUBqtQzLVMLs
HVmhBFCQ5WSbU2kmOjQk1GNFPIrDVRWOtfJLetxA95u6eCDqGecODIqEnGLXaJk5
/BQHhmNk1XmMRS3JCs/MFDK44W8tJO7iTVQmbSHoyyUf2dDHkko3gt4YigjPpEPz
FmueRKKfhcFAKjoiKpxJeMou+7FG/VSeSJRHkwS1uRSGbKc5nvEC6c2e+sTKHQMe
s39HaGN/ZqmTstnoq+LUI4o3XrgsNfqCnPim/N7urhAB4KyqiWazV+7KC7HfXKE9
xbc/y72+jrCvQUrrOTtydlMBsaHy9xJpL/jOJXy5rJRin/UFOQdr6d9eWXjAUqQn
OqxFApSnrJkZtG/hS5/DZdppHHQpbkdrZA93AQESV87QxaqHK9rgDL6aeS97yDFS
H/mcJhQlATl5GYme0NlI9Lxldk3PrWBuKI8kl8QqUAHylhkHwE/fCZSTPq4h14L4
uBhZu6wMyuGS6LWw9wDLoUn6YE3eM7+uBwJfPx82L9IF4H5gov1VYGifKoCBW9PU
SFbzGe04/yhtRnS1EYe2miaxOOir7t2bxJL9UVCtSn6PcuGTZfM+Vxn9UUxwEFao
JGW2U9aFk+8pRPbC0BUjdRqtGVPsLfTPF8MekgE12yYkM6+U5tyZokAyIuWgp3Hm
hptOlWx2yFj9IPqCsedUhUhUbDplqGVOikXaxt6uzbcRciB56EYEezl4+irJjxNi
4E6qstJbOnvE0yfYUxBEgIvJr0FqEJ8g7X8gtQnHViR1YeR4QSeH9VeoLuavYgas
FmTGAulvmjaJAKBsKDYOZAsPnN2pN3mkTosiuqegRWrhtaixvFagMmEQ9Vc3vuxu
nl2iejrZ7iSex+PDU/Bl2TFxi8p1QyDInOcSjIWUrepQuIuFuE26Py/UuxS8sqO4
PKJnnbU+s6PXo4peP27N0Nty82WMS3c4HZjnIBeCinSCu8cYEQmPFpH2Di3CtN1w
rIpNAxk7CJh+5WxNQR+jEzlqFrhOA2r1R8Stk9MzWQiXyM2RPauTxLq+t7qkecDn
NS/RZYfkCFyeNylYwTo//C+NtRJhugytB40cKEcNz9SljHOIKV/7EzTzQ82lRMWV
BfJbOh2uLQl3DstfD3WvZMhksAESDQHdUktCeOa8LUqPnaVjvxLlEft1ZU3DxQq+
Y1468ccirbNvqAuYbbH4f0XV+qSnD+uPoZDVJro+lC4tq9AgdViUKtw30gnd+dDc
qr8JbJFDk/ZUCnpaQkIRAlHmokxq3RwyyzGEX43kGhJHQ9SQuNp0QKcGGPX0Tq/q
i0KL1hLLxoPU6dcz8In3RRMJD+ktS9QjFV5eEAsq4JCeIx03MVIMjcld2VCyQVBx
qYHchXIh9oH++yhybo+fQtpN3kBIMbD2fw36yIB6Pu2aBQItu3Uy61MCm0bRx+XQ
LQEJxSoywUKwoRB8yS4yOycOjEwWhUkzie6qxabOJSDvRoNhlHAyyQ1RgdZJIyKY
wDVSzRydOrEce7rB/kKlBluDkW3GB20j5Q3+qOZ0Z1GcBIFbvcE12+iioZkICfS4
u0d3YRfUGONDSZ1+jYEGAWpC5eRItboKsNC9N/t/oypfQEKymJLFInHAFiDA1uRp
gIhCwbWCK+uPJzabt7o30nRQ8GuAYprUxW5BGo9LlEfig+SNayp1qz2DPH9NSNzn
4FniId2SBYllBOOeHq8DkfVJGvlH3BnK1cBIAqrRQYOQUYWpzCpGUrn5sPs6c3J0
brc3rmoycEwvmWxcJkshLIwMABTZ49AymGO94jjJSM8heuXzO7DC3fbHlV2xSTtZ
3CgR/ArbkUSvi31itWrJqphKZhDqvNqNJe8T/qGAvE5SdfMzlaaq2YDqtrklxeDO
X6S6i5eQLezdvQe2MJFRQswjKBt3Mfcuc7oXmogre1ye8FGWs2keNM3xOMWd1kkV
69ZBnNStjxIwqMjes02o8bIUhaqQ7CAY2x3VM+gavgZS5lHaYuBpzff5+J4S8QZJ
zh4Q0/t247rF9u4mWfSOU1jOlnB1AHLi1ysuwqK0TRpiq5hCdEyQpBniTKm33E7L
qAvIUYYKXjzYTOUx2XF1Is3tTqGH9DI4y/gQ9eU/DZ+F9CsseGRlg4QlfpxeN6Cf
0sJRcX40AqBTSqwId+ECGjIGm/7kUjkN7ir1uwqiib3XJ8Z3XAkvElod2F44EPxO
uxgiRSyhwM+USTLEgWKeHsHBPEZUAUogr5aSe3TbuGcPptCZi+8g+rua3vXg5cJk
SNQEG0cUzK0DLiiXNMIkk4ThmbSat4UdT+7c6/5CT5MdLbRjt3Lt5LjJJ0r+U20b
LNQNi64Pa4QzPyCzdchXKx8ntgjtF+/ibhDCbtISryx1/kY2vdeQXAQISY9/HTDf
knybAncAvM+T27I1a90uQop/JaR7uKzSwQjlwXM2ooO8/avhWU8n7F6FVuXxPgVA
Bx+ZzLcIBVrUxN2cC84oSVsK9bj5IE3a9YTwJLk8USsQilQF+Q1zqkcXxzeONUpm
N1AL3F7NTKKEfO6ORBo8QULul7yhKjen7VETmzUynjEhruQWmiuut1pnjHAvOVeT
FS5+WbwRHItj6oP0aOZcQT6SnmzpWkf14UbsSrewfib3ayu5OOqNhmCWh5GwKiDD
ofy3LYlLMqJFloK8opNPWyyRWcXcPX5HXz6740ikEbCIFXDuSfYz0JN5mpi+samq
Lk2fzl2Lj3JOw2n/fWFOv13YTBEl5mPpTHU5vE+ibcYHYKNmUvXCUdukI8WTuwWt
rB79H4YG0KyKL88DPJD/r0Wfx6MYjifcJ2rbteqo2egWQWFy0W5FygYetdnfnnus
IzpfGtOiqUYSOSCj73RjZBT1Cg9IPTc+EJMUCzcYlW5U3oCJhyeGpnqI1bt8GZrT
HtnDQyc6BSQTVxgNay9ci8etMA22h+G6Xs/vT10nlHy6Ok9MBhBfWzTvxrskh8mZ
/XxJxLms0xfPuXCL4teoO/HQ9CkjNT0RQeGlSxnNBaimomHiWAj0p3SpWQEqJ6hW
uwbQJS1VomyW7XJfQ04aSnj3t3aC2/jgbhe8MSozloN2WhFTkGU3tUFIm/PxISWJ
n57DQFx0qfoOmrBjOODuNNV/HbSHJi4m4eWRH2DK6Zl8i+1nCOCm8mg/VlIWzv4O
94ugp+GacrLpEjXZJmTaxz8nFp9oGgTA1TgCz3DekXTCH6THlfH8uvZv2lEkLvpF
WhPTITpzQvhCeclu+mrnYKt3Mlv8XsEKDfbweB5XQrunDDVqH52QCsQWbYQExwIE
8on9jEbqQqKsK5Y9iQjqfs4MScvDN/4XSPQBPLS3/F/xYFq+RYlYDKIor+bYmN8+
IeKok/JIfO8BTyybFD3sT8C8mJyQPhELO9Kj8+3ja8w8jr/Oyfy0LpU6GtAb4v9K
IF+Odd1ayoD+PLLXyOu9aojRKeF3m15IlC6ecZcbAmj8XGZwilPdTwXPKyoX2wy8
Q12LiyozzUcB3Hy153kHQwamtKjAwWCz66QOiwElxZBT3fuqefjTdpgQBxBmuQGJ
mnonnkdxv8nelPMx+T7Ad9i13cF5n5I7ga4L8B1UpNI0GZOvDL8ItvenFyWDUo0T
qfI2y+df6VQ5rYmuP2M41Ml8yUV5plflmWhcD49H3UO2W8BhXiY/U39/dGFjPie0
jdV6NAtW7EncdkzAS/0u6u3Hq6MNHEZgQBpGIAtrOWNB2oFzdu+nqCSEMD0UCnnX
qfdgpNsMcFdmtYhjYvhgPzxkZIs7xgxtLAUxfG4pCCWMBd8vlyhjVom6RYnKsYDT
tfChLl77bb/ud8p7SCPF6Ws81csrRtKm3LELcGlvYG14Rxs5QnI2HArxYIMRJVt9
vULQx8ovzyF5iaawcO7HNu4DW6naR69LxFpgKAgfFK/pN48VZ7z3Z5wSAGGKu79n
XXBmOzJnl2ds2oKSE4MEkVyEKHRejG+jO31PIx+1erdPB5ptAIGahR2vriJmgmUf
bZI+/mEPysDsQTsjE3KKY8ncsiUvhqcprAmv0jKsfCYI1dQQoe+69WYP4QtddUO5
8G2G8p4aUcil4q9u9SNIM1lgOjA3gHuDVz9oIzlAD9QOQn0CFHmXDCwA09zr/ooI
AEg40DLGED6ktmCtUN/vtIfSoL+ejZx5f4ELz7Nwqwfx6QJ+oefBn+32RNqz/DJU
MBlLF5nc+vGf0m/iWrckvxxg1xGK4UCnMyOmxULmmSY5fVK0jXvU3Dn1lzgZ8LNq
XjZmDd4MVAv5E8bzFAVOF6D/G0zk8PwLv5eNObidwcKewrmCxWfDL+INZvUUDkir
48XYzSZpchLPbdiD5p2WfZW497WtgW8NJwaGM8IDGuc58Lg2LBI922b9ysk5dmgz
F12Pub/VVgSXEVpTzzVi0V926LrKcs7peJ7EWQMtZHe1sAUhVLDD3U3gPog2sZYx
ZpeTS53SHWgsORZXPJECLoUJvIabXHrDmlBzvTcst//may6SF2FRAnnsKOlHe/48
4ez0prG97NnBoRuFfbrVj9dKMbig37JUavgyTefmgMIryBa9WCh5BfumXaQ8jPqG
+MAhiIoIDKxZFj6gDpoai50arKZ+iyiAhmkCqH+wZzfaRjsTG69qCJOMEKYM4Ssr
WJcoKx4107AFmsFKF1Ccpn6KyIuO9qhg426Y8wemHLQn1pmG2z9eT2Rr7K0Bt3wg
cGYYEqvJ8emoVwH55VjydqMb2B4JYKb6TI8l8AFLdk8pZA6pYLIl6qEz3nXQPKc9
m77tkHwEDxs5hJDSme2hCOlFm6evMFWvyQ6jDiZPLAM10dP1OfaWcyVunyZUJZS1
JeQQJzxLtPBie/k95JTqWJaovbYhFqFIo9F2/rX/Q7bAk9KcbZmacz6QSLqmZNGr
el32hOnqMKzxAa2iJZV/3GlPDz2dtcK6XRqm6mOqNDHZQhFo/egP19z5PB1OjpmX
QFp9+CNzMxEhpGeGqVDfApuI8lD1X2XWKXYtQlPgHy02oSKawUDESMWo5GMyfY4l
LtZ4Cw3XEl1aNgLcS9Jhnvs0venY+Rh2YBF9L2EUNfABbDOQwGAZBlawvUHvUTkC
VfIE3mm5FbMDcQaaT7pb+tN/qk4L5U/ddqM7IbnoL30bO3Tnqs8C1aCQ4pBpcx7c
K7K8TgtMTXaxWKzfEsWNn69+gcYbxZV+e13tyHB3rsfjSIBVZJ7eV5Ncz0b6ZurY
Njwvyymyh9j9vwugqeDtcBeattBKqXa3+f/3UUaeGMEtHZWzezZhQAJNpH0yX6EV
hyrbv4MvX+S8Pud+Mkcti9ObqTdKfg2vHUueuzQYFkkfQ7eXl3jdjR+rVNshUhdn
baRyPNeowXHfWbXALso+iIoP4JIVcNBX90Fc1H2A3OKo5cF8ehfytutgSVnjkMn/
ZDREP0oaNEYbYuOT7D8d0IrsGycYsqQ3Ud1xKIMCthAbWHXWsA6rU1aiX2WiBWQ4
aMWfFY1pys8jwjjO31a87E3ETwyUZknKzjIaOlxAniW4Vi3F0UXRJCUhIlVCN5YA
NGcV9PJ0Tdlt4ER8q4gxVaC1D8rFvx+YhjqMaqd/zVx169jkGzDW1BZi/u6+3FOV
zU2TtOsbE2tkylOtfWr2DtsePOwNE5I4VzKBEwhvaz1Y6JBQ2qdg66NIDc6OhrrE
QS6UhPuabTgYPsh5LNP7P2aBCk7Fs/h7qLp3UZjm4mizwlhQhWC/IrvPRr8vvF2n
dmtFY6B+MioASPwz8BdLAwBznClZ0Juf9sUbQIdYuZuGF2OFa/22maYglaNum4A5
iXD3dpPmeYFrP1Bh0WrC9akBSDq9yf8Y6OaVylikjumd/k9a09RdLiMEvQU0vcHR
GChO6AriJN6/j4cRP7WMdenAgrRVS8vx4JWII8O0EzF3yUsv63YcR5P0+pB62xqT
O5piPdFRoUs9OfpGaJseZuA6V8jY0as/woU4oznTS7MqQCpPaNW40IKXE6gpR5NX
Up1YptUXaz1j6dvoAk2UxQ7YvbhoHxNOJeC4WAiQKP3G/9aiTXB+iXCg7FrpX8JX
fQ+LMnM28OF0V7kNhHGT81rmaXzGK9+djyKJVG/TSiXKwdwPO2lL1wsEeVbLE6a2
L7mP6EUxGHG1/JZfsYJbN93+6y3QEK/r7kl9ly0Yxhm9vK1GuNRzQblPjenKszmu
sj8btdzcoi3yWeL5PZzDf5svB/Oe73grpUzQbMXnydBKLyqcpiuyYOsMJIYKK/Yv
XxuzoHCcpD32SDJYZrDNenB6q+LOvED7jZpkGtdoaRb1TzqDdnz+tIPpuIhxZRK4
YNtJZ6a/v5YvgDhQeNXzsLopolNNPRfu5dttkRmMOWDfrp7H/QN7U/xuh4O99TZl
avfl3FgI1SXubSgJhz55Z58RLc+LJ/YyQnvgjdiQbcKiXrogx9rQo9NeOxNaCy6c
wYs+ffoiclHkEMS3RnpUvO/TjETwMhlnBcqJK4oLlWnhP6w75b7DOSIdwOETXyi0
aRE08PmMYjR71+1veklg4yGd2MzMSK1Kf+8O+KyO7iU+oUxsBLC0Ljta3VgPo3TH
p2O2bwy1HHQ+Vui+oZoxScFCt9ZpfhDeZb2sgRagwauwMM32uDAKyOvx0iBIeryo
LBXDF/LhhJ9btxAYLSMCnHkl4iMtThlrlpgA8e+aPlbhT7Jy6uVSG3kLlOLQqWKv
cz6FgWndmaWHGPho38s1wpfZ2qu/N7E90FZ7IjB/agYe97lDUihWOv6jg98GVJsW
9uksohKVUhuejAXoEzUcCgl4F6KNLt0FktrLmPb5QEL7OneMhqxCnNB1OShztpJ9
PL3OFs0386pwYnYG2/qoXkxtsLXFgV+v2FlCWPylVfgrn9KVBwrEcVS8+2e0BtC6
kiMRkDJ5RZVmH7/V4E0b8p7V0SvjCUqJ0JHBU9562rJfF9G+PkUb1mCUmA8dfN1+
YGl4PbGqwAwmuCq7gVsOhzWutCYcYI2DBTqQl8vJrlyXZgUVsg2m/HJgHNm39SJe
iiKI/Q0+6870n9j8xQOY/Z/uOhKcdiEG45Yv35H0ZNtj+53jtAVqrrdH5KAHRG8K
31pyXDsne+f0KaEmjGMA4OQNGf4rJuTeSBKpdlxoiX3OBMbTx9MuAWey/y/V5QVn
afgj+BmC2PNr0pcd+snWHUqXkznDqQr20qIN7ChX8n/0OSjkiCSAJzi5oixqKAWr
C/8mBdYeX8m/tKUVT4hhx1ZfT4HFc2KcbsyygE/FK8Murw+6Dn0jWaXdKgZM3xXd
eDIW6zP4Rt8Dl97NHv2hOgRMJWeOtpu/CphJhswfAcamTHKb+BqPRoEXeFW90Sfi
W1GZYgVs+n8QctwOYp/s9VrierLjuZ8I0V+Ao+DoyyGghQZzK33LKThwv9pO41EN
Xco0jW/0LhvnaZgRyBNhgp6JT48BPFYtUjwaDqD7+2iPch6Hx5hYvb1oYEoqvLPd
qIzJJ+3j97CHB8guFOxdhBEUzni/rLgBIk5YUrsOP60Ni3WnrQ7otKAebHBZYNKe
ArVHyferSB5lygvbGaB+rfQ2b25EJU0Z33dhzrlnJaa6fUYCETG4aw66EHcp4kwi
Z8UqNOsLsjAEvcrJm//hr03LWGBF18TzHB+T1Rj+e77bu4bK0SFKt7+ePjZsZuV+
q3HeSxL6EBBmxUmdz8WtAdQp0QnDJwBYvcCybZ3g6NjI81Vw7/cVUoUzp32/Rkov
tu3i9td6Ph6HY8MGBfNTPjsJNVbEIl3rRICB7Ts4TvuMl7kSggE4TF3Gzdq1XKbh
MBrIZ0ngEXKegmwQqcdJLfA4V2UrEVHfmTmnxXFZx/kVge1ZVhYIhWDAVSNHtBF5
nQKFD5rCGSpjfKwosi3KpK/hVXrhe7W0nlLcYcw7hv0tyuxZATwhdVpzmVe0Ta4g
ew+ravfhPtmnOzcf56fuhRvXN05UQOND0vjNQWMG9qCo+GZpob9ZbssEE7St/wzA
T64TYwNWFxt5mGjJ89PuM6ExrpV2ldQ3pDcxATYKwDkxJNGKnE7L/dZq441N2Mz6
B8jLQjmdqgiplB0Q4/c7lz/A8amB/EYHC7fOawenwsxa49f1BDMmJQ/qvbbU4Yj0
j+jAHzK4H7tFH/6VlSyr/axtYLx+e28ik3uILWYT/WdJ6t86X/nLEzQGlzWysw34
d3WawgEZ/2D3Lnowj7YYVebFtFMySW9vWPqXF1FN7Nf7yIaunHGeBXDSI9Hio6+R
Lu6xyS787qoRS7NkL9P2l9BllxicLvZh9ESgw8ieeQ+AdU/D3QlMyAF30SPXYNLZ
d6MgH6xf0ULnjqh3dAi/IhkSK2hNweFCRD+6vIHrU6LtnHoy8CouQLdygrTrYrP2
RzxUEKOT4JvHwmbx5d4LqN9X8Ecatkou9aG54H63Xy6tefV/EbxTHph+MM5SfIKn
ec7jp35yzJ1V+oeEGIIm7LRjKag7uOluulpcPtZqulnuDZFihNNs5agqQVHS36E0
XNAj5aimGFLAMEzijBFwKKgnEz4xvtTimktoqn9FQOOgRONCq5hKDKR3Di1OlRe7
9dhwMH9WCSLe3A6YyRutYmaD4pgIh9yiMy/0QVCsxeH/bAygpHbbvF2T/qhFrEsO
aUjCS+CVuupKPuM994pXBMwHwD4fMjJ8qFZqxlqofLbwQrRX7QuwhuV5oO1Jgp8H
/1aVTW6tbfUJO088u+QcHRBppKDXo0qfjUEEYX7feUgHqGyMsJkk22HlP5ZzkgRr
aXM45L/84mvwqHl8+vmWAy8IRqVxq00SK9Mf5JpnnJu1km+4Uo3CkNXmbqi3eY4j
oJAGAWaTu6YvckJPoAyMsE8DFs7J69pvXx3XRPgTAO5xpdCQNY1usc9XL9NBJ7GB
rjoh9R0r4sOjgbs0RNCsQe5Bw5VB0j9SkCAVraG7bwLEGaFxa+MtCWxdKThcDgAS
IiKXTEStC/GGK0r6dgAMy3xqg0CQ9/5iI0ij/5wdbT3eVnagyxREeYT1tdKRSxaz
FodhxhxOf+LjqYtQB2AokaG5E2hN200vSyE1lIsUWuL/hsB3d33H1e16VqtEQ5Fd
PRbnAsFdBYNa8JJn4Km2DS88Vls9tntCEN16me6ccMmIvfEbhn8iVW2CUnysUPP6
vVHcKDha1oMTF2MrA7yzezNcEmIL0rlbzCsod5a53jqpgyGRaxzZ79/CGIkYx96E
JCXhftRJBpixT/HL86vOIblN8uqhJFTza12kfJukCVUn1xGMKjq+lKjT1ve7K2b+
hgTCauubWX6J9vxcEGqYet8ZCQ9GOdF4ueQWzz7gbYrCKyFjUb8XvZJJ2GeIHXO8
wZjBlXDvnQVv/1WqYw5nVWRujZZkzK6xw3Nkz5ruXFEP9V+SavHDdQQFQQvgy4HK
aqUD8kMWc41qz2QLJL5Qzq4HWFdmMCYJtpSNS3+yDACXCNOh9Hp06Qxg6a3nka+f
Uc4itCQYVKi96lkxdHY/TuGLUUAfHWGseYXh/jj5CZezSWD4WP8s7IreQbzuVjUr
V1YoYGdL2ODaTP81dVe782wtKprlEbFIpu7dWdibtY+cQRfEmGCUajtJjmzyEV4L
1l4DGRnRQXSxLKnDYGXxHC9P7ZfK8kB6jnmd4EIawyrB37Y8oJrGjERuwTAMEu/C
KXg4c8EM+xbzU6LFofJB1QTDH6wOWF5quunK8czTvAG2P34tImkobKIyJT8YcORt
0G9x2T36XDqXpR+iC5sfom3kfE5WdLylFyISbzybkv2ANn+LUhMdbdruh8Wo6RbT
MEqOEEANLTpYbLBvISOi5IbGNLezMMxp91gh65HrcI9yXVOkOQvGt+dpC36pvhUC
x3QJEioPKJFt6Sz8LpHWFwfItxgji6LLaWQb9nqWxbOP2X+xOnQkJYHdkXM2lDGO
/5wAfXaIvmiNfdluA85oSjFha8NtfctZvgMTc++DKHbj541tqkiB8y9RwGs6OUFC
UN69d/aNZ2a+Vmm9cwpbc8lk0CCBq2W2qM1Vo/12jjO5qlHwRrhuVIq9pUk/C1Nr
EJfBuyKtCN4TA/xhN4loOXC0tDWXsbjrd6WedWoaADaehgLKcaEzXPxAyNa6ZDqu
dXh9BYbEsJxew1HFIps1CpCtDOHuifRltJy+uxQaGYKpdfuRtHL37hBUbNNj0eHw
NW1I7B7FMH5lP7FqzvuB7yrbJb9x0OBCpJP5bv3iydl5k8f5vrC27UVRMynfOHrs
B+i8LQZ8LTGle+gWrTP1g+wEc8wpd2IUemPbJE22e7S9DUJYBnjGk3n9Nbv42GpB
97ieENc7l1FzSO47Rm9IheoBIjNbLsjSgMMTt9EVZkLfznG+i2gEOzy33g7H4BIL
Vkpp83eZQKXheYpIAmbTfzUbx4/0Q8wB2DyBFSa71h0qCP8SS610OZkL9zJiII9C
r45AMu5iZndae7PRlgRoBv4EvzxL4xR9FMK6N991dWNS3sXPN7ZeO+3FXV6viHA5
NETETLp8ISKTj5+ybxzO7LUEiVC366LGB1XKpLEDioDObeDBpJDXiT22AQFVLedz
Erm3FDUiiHqieSvJYy7681Teg5IX+pevjbxSQwTU93Y1zaZrOdhWRgy7KTIZ+pmU
JgcZCe63OVGE17CxT5mRaGy8Yqi1mUbEhtyPQlj4HT6J4dLGZQG3AtexNe4bhsfW
Hcnq+2KhxOaFU89GWN+oOWBaYg6KDd3g2lESffQdlXRM2D0ARLyoAcJJ7i/uWZGA
qlicjqtQGSooZhFecamb/lfCup74/mIWZXwrA4trCKrx/SuoMPbwyKlEHcyhg7zE
dB0ZkZiWpYCBmmrEEgvkutL2wShpEfvItwqBWRtlatxRzv2w6xIY/PbyXoQ5RI4j
ChOnBecj9vpb+gCJyt5gCvf+b25zlDI7i3OCIm852cWANm1FlbpajnhEpOfqToqu
9KxgC/XRVOpqveDZ2Ef2xQwVqNLQqvLBDkhZGxcuG5Co8/+uhQzaQWxOWFSVhku1
nD/R20taRGRX1pfSSF5nGG9fFuvdN0WcDpau8qCZdyLv8xsnJrH3jOt6NYG50vMY
j6jZIEzgUfhMQAyE5Gu4lEGc+eVnkaKDOMwLfqEOmZA5yzJTubf75iza81hrIxUY
nJwowLCVknaalgTxwR/nYbLmH8ogUmZTqOQ8hqbMQYl97KnLe55wEF9AfGBTWMH9
RIUqiVyG1esxQfmkUqXahRJRgHtWUJ3VVBsa8lNvXsh3rwOp8/OU044UBk6h1OEe
2mtd4C56OWAyx5gS3r6CbMiBhZzDR6Tn33FTUeJHht773pqF9/XhaeHf2Gt/v+EV
40qUfKfIY3KlESwza9eMC14FAGRLaV1mx9NdX25Y3yQfXIA3rKjynt1JLu0RfVfL
BJ/G6jOmbWr4bouLNXp9HoKoRqAEa1WweLrh8l3F0CgnR79Ek9P6I7lVlyM4P9rQ
zdisj1PSHn8U/xzo6UlLwwmy8uxLPlBXfok2Luz+73Mk6jbj+RR2ZfrN1Dylgy2h
EgGo+eI7PlA+GP8j7Or6hgMKrPC/XasrzZnwYzQoRBb4UZNxICeF+5cwcOhPsRS7
2t1PnbFonqATqvrVhRmxjawrxlXY89IxFnXVelHc+syJC+mGl/Lz7m50DuTN/wGU
MD7dLH22m6dtwdeFnyU9LCYQ9O/Wwxh4mbOeEuqPPHkxlrpPbgxQX7ZwxxMIJArW
oGginGXv4b4f7pws+Wtw1hNWe+ipREesSQTX1ydMcQB8EMJ0wgHFP/kmljvjsPj1
T2jWhOKzqzwUApcHwGchxR0ZB5LaSbNNHde+x19Q+M29urlKh0VHcYx+1zSM0WaX
TX0Gs7AkTwg7h1KrRiqsJwd0t6b5TtNu6xx/W9I/BV9xqqel5KOCMu7Y8ZLze1DK
M5Wd8ndQj6xqH7QEKtBAmUiFyuITYG03XUm9SXVGjUZVt06OjWVdTDFjTPwzpbLe
rESIKcB0DAFewrjFxyp3yJeAOuYIr4IqsGAWk41w7WRh6ii9H4UMkh/GRbSaO9Mc
NgM0Tm+AMbuoH6ftSAK6A+rGiY/JYWMgQsqrRp3fPFMMY59Qjlcd1GuSHDiO69/7
gLKlb7m1Eobh3kcN3jpSGzBO2SoOUgWqPwbQTDfCwsXqLBs2tly21wLjAWB6wR1I
zC8dpTdyvLl0Ab7RAKzQ/tghvm8CzX9FFdvHuV55NOBLNgwGmAmMQnT7pXT0XpSd
yBwv2tE8IBIZwD1+m70LtCnixdZWLFIwHFlw0wTaCrFSPwtxUNznFXJmZhE5xlLz
+1W32WjQhxOuNB4UWM+S7cPu21qLePBdffK5I3H6wbhG4ja/bcaY8/unSvaWMlLm
sNiX9AjLLg9mxioYpqPDIvNvBJJlgImok3i6LLCg1BEhyM0JDN1JUb+vXHX5lxM2
SzyYdHydsvIHVZ8GVX9XGojzm+N7g29JX3gCnXQuaIsPvD+Rb+VhVmbiwZQctnO6
tbE7utwb4P5jQEUUZZJqCDmlTwvHmd3VtYPpgcjsD1GgREfm7jZ2Zs5cPVjRfOQl
PwypxwMUgL0Gleh70dAo+9dj9Cdxb4Cz8nWyQnOJlQaFAwYry+8qZuKbaPli32Ga
XjA59E+onUkmHaCYhWjpgExejZVP/F6qlCvLYttD6GMAA0xhDsiJ5beLqnURWqco
LXjGf3F2kYwpBGSUixYA78vld176s0G5OBr6ICb/2rk9bciAckK5i2p0MbuDUcNj
SHFegYD1RhyVX1JaTgytzmIIU/RlQ4snkInJWzF0b/OyXuZnPU5uaYqniNX/cCqO
Dg4uLJ0wRO9QdB4HZNS8KQWau4Bhac8VZNqPPgPnEFt20JsDbK/JrMtG9c26IHvp
GItJnXDd/YLM/spegRtaWbc0b11qiD2g1p9BUq1rpsLR4M+TUHj4yEtyW9OOmBAv
Jf0x8YLmbBUOM1TJnGPNy/n3pKmPVabpsqoPTVY6x5APbTNjrRRrRd+Q4CC9C8Ie
4uTWr0jXd4UTQwqZFxCvSoryL06M+cZUahSEtuFprNmvLRDCBIlBhQOE+cinlqJm
qkoTmSqYnDozVlhviMXcwdkIFJiH5A9OMAZYqy2/7hX8aW22EuCtubTnDCMjBBHv
LGOu0+8u2wtUmhUzIn5ROdY8RboyXeAHuIwOgmso1PRDgY/9tCDdhbsclyXRJVRY
xRVuuQaagVvSDcEdkrO8gsoAGYGjUdGcdSxAL19cg6IFOJEdyxGZfQxvRde9DqYJ
udvkEDbr2a+GheabGdcw/IA+hRFoHergObsu5GpQdgbFMXTedv9VewBVkghLuKSz
YtitS95p7Z1mR4jWY4m5gBHytjlEBO9xYUlFeRG4qpYWwMez4jUIER/dn1CtQQXR
Ex3LGTd5C1lug2QHjBMPW4PrMmR8RPe2xCPEhoz6kwzqcy1sBLxXFbCOlXNUME8/
i775F+sdU3XcIoIrFGIZHKqNdLktQYwXXU55+8vl2JeZw/aJPcrGE5kyoJS83pyi
GePsMHDPk3l9Q0R/XchlVpt+SxK1CsA7hZug78lvyigdA4mFud1L8EWNBlCPQeDU
y4oIKxT9mET8Lwkt3Qd9JENQXu5E4bwY/Swve2am9rgSmSMBylyIf035NTtIOM/C
Pwj94uukNU40LKmrkEIuBX1gVvg5kZArIYsKu5mJDxzPfuYRRPG9z+4k1ULrCwu5
YV5Rddg4dYYe0yU43jMRdho0man1wyLXUJXYeM3s+oi+oNEW36h4MkWdoHBlX49N
5Pu8tOmCIpkI/pxpjEnd08Atfa3KStYOywCg5ggCyX1i7hn5L677dbfqesksmxKr
dwo1fatBTMQHEGS2+aaQd/v/LAokmLXHWPoa0ijtHMagE8o9SsGgeEQLt6d7AlFs
AMVh6sAdAXj40intjcPG1YF88O5aewPs7yK5FErkbI7RgnUEjD2uPOGTcdTLoUeJ
KeTxDD+d2yXdFki2CJBtDwYeUUjeVsn5kbMj3+m/EI76bw6PmlsyfIdxhZTDoKKN
eC0wKb/7o9m0jT6SSBSMIa2nY3euO88MZgPhYwYGG07H1MdarCaPu8MhbrZXuz7j
ZVTc/RZxqXNlcsbTz02eptJsQjJyajHuA0U3xVKbB6E1pmAdc8xLGCwRLQ9R8vR9
b/AYbB5EnlAhheRZaSc5xIzUhDYJIjk9PYWlwfcpfC62DraJJi0nRe3fZ+PqazSi
a94azWm7kH+6TAEUShLoez+EPR+pChgw8OfSrVPBe7752Gskb8QZww9dDeMzg9gS
kD06EPgLS2GMwWSBa43chz2Tj93KX1bL3zUntrSXc+KjNFg/INxfUwjFWXhfAbJY
yFyeM1IwzivxlQW2VAP+q9YhBRYAp4oLAKj7lSPvV2v380p3iqa494WdYgr59Vuk
82cttJcM2NAT5D+yJHCK2x17TqcqDEShy6VOkCbz0cKYTeMTu0x3t6pvkcCe/Ou+
tcaYsZjSVLa38fUYE/TrUkx5B4rU7OYrOOoK+qXww2jXOIaRTRu/aMafWgkiZeP2
hU1Se7fuA7yzAKve3Ud3dzbY1qbPYTCiHI8uY697p4X0bJOrjRfxwSyJMPJMAmeX
ffBTeduqvfk9M7N7usohR42nM8cGUloxZCjpNGYUBqJr/A9sWJpako7X/7qKBAZG
cRvtreck12wnCv189JBN+bG/NZ91B17OxullXH5bTqmijgP6QgirYRdByn/BEV/W
pSn1XkmJxouDKjr6MoZ2rfu8ZdxIB8ga3zZEV1tfpvKKD4RUTvvDRIscctCAYE3o
CwjbjfmLfUBCfi+kjJxbOMtqPV9BZjNhs7nAKPKEvLXbgn+AuuC79dCZtlD4ZdBT
ZUNFI1o29Fl2pf93k93pQvhNKIdTQmWrIXyxL3PGy8faTp1d9wgfJYWKf1nnwzZ2
uvSuj1VCSMtvY6Hq/2ygpUgAoRvAuT+oajHDViF2MGc+0M9MdPYXZBW8p0bE8rex
2mRxNW66AlRdIN8K4RFSxNDohFuVLc5ElvjvwkffeubmV73mSsq3tXEZ3fkIix89
rjjGUyhJzh1/ssztP0BdJDVWTJl/6gjlhwwtyr1n2qu/c9Cvnj4C4rs9ftX+o3uS
MLm3ySRktDCyxRmoQYFYFFi9It44sTSd276JFIoEv/e2c72sgxxWib+KL6rSY98z
/dacf4PNE/ObERrf9iiHNuoic0HckaqbppQOGhvLWP/oihpgwkZ1jHl/AEUs1oUv
tSXSgMWbIJOCIM0lJlJARHm7FmbfmBhWNinNJn9sU3DpwVh6EX7tGnEapMWTV37o
WKUBCjhsTzzIxjNPGM+/VLQiUWtM55mgngFAn95Ou3dQRn3wU4r/9I8wQ1607kHv
AnAPeZQTgChbnh2e5KDXEMztPkoT46sjyk6G7I9dHFzuYYl6I4lUvNNB3UfSYMrc
90VZ+aJcQ2Txcucw/E0R0k/HsAs20wl2rs9oOZ6eaFCrGeKhwJ6aBHlMWurDiL1h
hrnjj9MaCWW1HZDpUwS3rIeEkr+8kpYwkgVCpYwCzJg/cXdis0i0QqZsHlEJERjH
Hy0ibuozh0J8FNm95p+3ROc2mpVvPU1ry7LJ14OHCpLGj4G0DJBfEAMcm4nNBLV2
iP1ZsUoHkaFJgG4qlcLDqej4Wu7bgELYRtPTICvwJ16DWSBfVz128tgmIB46UcaJ
EZFE91SfMLlqL79191P4iJLYsb6+rDjzoNaV0I/I2OVnKb8XPIrOMPomuKagam4X
7xHCxbVhTUZrXQ6c3FXaPAF5s8i2Cr3ykAJnheayiIWAwaQuLm7KWhB0845njQ5t
aTy0D9jYwbZg9uzlY9q6ZaakYmvdNMQd2h/boP1uZr2dk3F86YN/kfuI142KUWl0
cXy4OEVu2/df2op3imG5fAhtItf8EN+paBI/oBVYQuYV8v8xAugYWH5kvP+Xvuyy
jk2P8sgA7FZy9XN69SKqn/asugKvjgjtG95K6sbzxJxFdpeVy1hF3pNVsLl5j96d
+eZp+d8SibeJmfWuIKu6IDoiV2jptRh+StX3eUJZnG8sfCyxbrl41YbSeGaknwfr
1akl3Ck+5vJVnO4/1CEaD1iqKk7fNkvJq1bpBV7X1XLQzbSZMl2yvVyoROgW9kOq
cBM1gNZoOECr5IQU2dI9EKsIUkI5xhXOqAQae9uDqICyYgwtFfDXp6jnWJsehU6r
yIA3wkvNldJEE3bbIE99eWombmwC7kGdStH7i+rxyK/eVr20MZBQ62Tas6OnX9jK
9L3tq7L0TX4wND9E+PpvX0I/FgW5/T5audleYE/ecOZwZiHcU7FtkJNsablJ4fZp
ByCxQwndS20LeLgkwtu5TaSZbNVgPcbDpnuYgWlH1S55CT4h+6U8/6jSKStWQChc
ox7xhz3UZGYOd6ZKPH7P1Bc0sHVqazdFTDklLD9laadpsXZc9dRL6ng2Q/nQ/Fx4
CnVvUVOQV5AnvocF/b1n+4viwIvldJ14y7GfRvzY2eeyh6k6DHoq5ueXtiJEla+o
Slinxgz/uvutFWVsnRyk1k+t34/S2ASe/U+FEVTVbhyGL5wKFrDXPqWVR9qhtU7o
JkS0JsEaVCL330AmkLunmPULvwuEbFOucbyOrp134SdKpQl9glvH7KbfiGS+TiFo
lNG7qEFqn663dK04x3nIBanl0VnrJ1onEhEVGwH6uaIgUpaLVRPCmT4KDV/dE+Oo
oI1hnPlWH91O1N09LR3fSWVzuRG0I8ounqDWYUMo+O1E/Xgh4oFHl6HA751Bl5kW
KwfyxIT5He9+1j2nGq6RqUj4ZpwWPxAeZEd3USigZnCAFPfvymfrUcE2q6pZcmY7
sko9iEm6LLtMQPGaN6XlYzteNps3BJ8RPAUImdk2yvNo77h5GTYPNUTexHo9CkAd
2LUQy0/XYnTkfm+D1zRRgXQu7TH1UqcrAnR9Ld9EKwiIRmixSLeEusYH52gHBjiD
ORsF7RUsFhGQ1MSKaPyUI+3KBCtsZubTsE+iHlDeZICIiyRDHPvDHWJF4l4vfnHI
cPKgq5+OF3X5M4PQM3IdKPx6cGbIm7f8vu2QHk904LBVkg0bEd9Lkb314Coyf8KN
vrbbIINHM6gJ2WtaEgbIXnxxIQwkjcDSX41v5ZQsDdc+BxxDCBv+mxnTglI87DFT
IXilhIkSFi9rD+7g2x5SPQd+eqOigxWwiKop3A5Biuo+gmBCpCgNGHlvz3tRTMqD
hCD5McYoWV4VZbd3R8N5PeOgZ81Dap7NTB7XI8L5cGfg3P2raC5NJIV0735SRNTS
fVQ2sYyIGaot+XNDgY3lD38jJFI+4V6BNll/7p/eQHtQ70c39j7Pij8s4tNHfmlm
BGOrSlOK/mn/kyT0xF+1q4inmhLVESDjkIaoi5L1OqVkP8eccmMLqulz7mcWGTsP
ayXBzD2bBVxUaYamma/V/28zdIC82Kr4IedSTNKdCQO0ucmtiLReSUjo4M//u7RI
HmvhcbUoOWoaZ+b4fT9rGjdgHSsTcgcOD1x5IRA8lgqhVyGuE8uyT22XMYxSyEyM
GGhLwa6wlHW8n8qptO/xq1URt6EtV9EPgeNE4a18o+G3nY2pdDTXHMOL4Eh7TCAP
3sAhQHfrmzxV/b5lhgl92vShG81C19wlofYLC/YyxYyCc/agpJWrv/q6nHdhE4dw
I8+LYEeeacholeZhw8Mh7senrm2R9i/fLoi3HhA6IjcPiZXRUNMRgHL/YYP9C4zR
x90xdnxnjAYfkTpAiS/L3oZo20FbbJT10pNTaEVXdf+6zUUsWQCrU6MKnPtWPDh/
iVHGPQaODaXJotM9AFiM1Zgvc30OEHx8akjKRCDo1kpFA6LQNYZBqx0OWEUfQP2Z
mlLyGwYHKellb536nb6WHglCq11KXxt05oxCIG/WtbHwU3z3up/IOnG4v/7Aux3j
ww7rwI5+OSFfLmT8Cg1K6vBnGcT1KZFixib1dGbm9yNZs4bw1f4SXoMytxLg14WS
kqpX13DmQNVg9vVi92IeCtxmFPL5rlk3N2h4wAS+b1oM/LQdPrD5fAo14AfWmu/Y
HSTfQGYXA+AYEWHHzykjjW2tu9IIrdIxck1hNaY1uMjttmDW2HVUKV6MDbg3mSW9
ACf5YIPhmLwa65dV3s0dbGbd94KQ2TyuhMv4xDhB28HnyZ98pjVeYlrU5u7EAD3v
T4v3ejC5Xe9FlBhVQkmE53SudP0byswa4uhjCM3MK77r5ikiPrIhh7BRhqfdvl1I
y9oHIqX26BG22OH3s1rDsA8DHxMPi7iUeTOOwLTEnTPV0qEX6tMOlFRAee53MfJJ
UM4V5yS8wnhS3y/Yhxj8uYjJkVTANrG2sfmroi30EdpuSLG9AN7Od0r4HeEPsPMn
TR92dXeVNkZYXr+Bvpd3CKph8ZpuUdy6kMPHougnQgeJGalpJy8XBzrwtsWq+owY
yYBSXYIT0V5TugHxXeT10PnBP9lsTPFKLna60/PUzg5uXpAqlP1Y6QN/nCK37JVY
FGXrGDhB1UCE0fQGi+jCdRjXKfSbIpDC4d2U0FGcdZJuHfxw6pjUe+Kbat774Igb
AIN/fzDCQT47C9luWMJlkpuL1DbNhFrW4ZIcXj+8xvgBqhurbQITAkkP4mJ7lflF
pH3BvXtIydlzbtWT8j2VBU2RNdrrS5zAYKHCYOg0apZUNq747gLIaXNyQVaO24Jz
OQ0n54mBf5AeYF6xd2PVxgR56Qj7Hj/PrwaOebyOPIzdLm9luE9MmdytoGEKLHYE
GqjYZrqACpFwouuSLQuheEhan+v1wNrNxAQgA+z9vq8TKfKEchqVRAi4D9gyeMue
3hFWzeCjyCf077Q6V4NgHn17BGW+WyC3z73Bgx4Vq2LfwkFPk9VNikAWiYnQkRyp
c2OvW5TNqdh4+MDKrseVisYaFdbxhz6rDq8FAddph4ctRvyJkcql0QeBdU+ezvMG
qs1cQWsbf0IABsYrfSdiEvavAUsqXuzR/xviw10Z0Gz+wSZrLO9q9NiYNmOTL1ow
j0wtGmSHptDrZ4W0qKB5xFT24pNGoP1zOyLNFV8w5SWhUCA+sR+wR65wmFRLd0gm
8EWGljrEbRplq3m8ILm8NiGlSKXeCSS3l1ChKZ1XbHenGfvg0ekpcx+A5L6E9AhE
jWsEYyMqoi6HhnfSNGpknyniUEzFWWpM9GXktRyFw5hyn/aH2z2LaTDOpMT739+C
dP/m9k6Y7oc6R78gq/QRJTTWdd82RdzHIVw0vYbcqkW1OOmBEX+ST34lIFrWU3p1
4PXRYMEXlivlFJEhHmUDpeTml19amX/peqnhbiiK3CbLbhN51Ghth8NpHB6p69a9
xfrs5k+kGQcOyIpXcdAuxHRB10GzFzJUZyRkLwBPGPEoMfzXDg1N/67P6IlQSeoD
AQ3uNlwIrY0wqtK/t6kSC8JoKxI80dUnugu1G99Hw0t3Wpj/TkdYzYVszgOs6P4F
AxHERrHWsD4fe6SXsNkrSS7sFpV9mfTT8kTUUQpBerjMvVmzwWznpMGo5160I5/Q
GpJy2LHwcadlQff2VOJhwN9bdJZk7vMK4mcaqGS3lP4MF2ztVgEE9ktfI4/eImkx
wr8HUqoNTxybrWVZ0A3dtQivR7F3TV1GQr2EkPOiTDGF4U9EAwRh9X+NKsFhOSFS
fTdEOYASITeRWoJv4HDgx+GWX8n79a4So0ZcpKyDi3X/Yh25iIRNctxKt2gmDikt
35A+KFWQkD5HHgYMXsFSOczPSu7hhTCIWhbwaGSmM8xTXKZK7vuvoktH8SI4wIYI
5lKU3ryoAEsXmtELINIkvGTLIhSxx4CZInVzhImyYeTSAHqqSzeL4dTB8U3z90PH
f33NNWrJZBMRV2y4ruwpeX+sKvPuVy/OhfNZD80NUxKKWLJ4oib3s+vrIcxAsXFo
GizJzwPWeiCXsuwJ/goBJT9fk4pc0CeG0IrGKvNt3ckYuq5BWqI2O2lccS5RFIuN
kOPdqJiy5xW0OVB0+w7kPutRcZfObgs3xwNUN0Clw9heJ2lIL8t+ozhpzNDnglw5
E1yD3bg19koQ8wjwkQooMf6aWQ4GCpSbpKFcUIojsenoiEIMFI/8KFgSBMoXTqqO
ST6Cg+Feab53VLVxr7zcJFbjZ1WjsD4tBE72otQq8QIo9lAis0WCvXS2GIZ7Oxjs
+kNMbbQYeYAZnpoPPMGvNEEIXSU3OkEFid6I3yQwegzVhNj1BTmtT9U08GSDXQvL
XyPBApv/uiKn2Dv6o8MyZ7JuDzjA0no/UeCFZ7h4mlYONwDllBNZtjVGS9hz6HKe
O8akAeXMEyBDqQ/m+9F6KkzK1YlVcqJKJQE4Xrps4ceUJDJVgt+8eNg8b4thlSmH
XWQAzS/4dgx/s4gcpLJzYSiGG381LGOdYMUyqaJMrkiyYuEitUNNLe+qhgfw7k9Y
tghrrULvUib2DcVyBqg/o1N7d1Hq1svBxnzxWC6S3xQ4+TdnXOqk4xN0A1Rwn6pP
6fKuQHBRbC9BU0E+eueBF33LpuuHR4+7vARtSWT7L0mdVKNxfetTzTRdg/lreiRX
ggiB3kJTFRWcKLArseIlicix0s5rmtqi6sF6mUAtnJdMw3ur/bev+n8SlN/QDDMO
vcLKEOl1XlGaIMvSOu/AkSPIVDwXvrV2mCDmUK0PcyvgQNWfWczPE4htzZA9U4Ft
CGYS2q3BK8w8G5y6JQMvSbLgFJ3OX5liFuf3TmsW7wExlM9P6T9pGR2hceZQuQ1Y
oNBiWcYaZflt1O9aZvx02mvEvIdJKZymE8o/QS5rDvqKPQLtDou8Ic+dDvd5U5Ar
ZSYfovlCgRu6L+wkJLQrtzAxDo9IVB31daii+sma7A7n0BXuIERUtE0kJusf2xk6
367mjLsTuCv9imEzq0ceqoBaokjyNqmJdjhHz0FKJ6ecfPWzx7YUbLLDfVWnniAy
eaQ4g03TwrHjTRu3IGwtCOc4NKOKgnR6urHMUReGXJLTNKW7MNobUHebXiXPSSoK
FDKfjD7tWftBzKRUtrnRxtpt5f9VnmzDLgx+yDLPDoNS1+OuIqj2tiNY7p3YfFZN
Eq34tOYrPaztluN0ZCGvZOdx7HtvnJ9gIbZvuWQGh5udzeGMcxfOpt7w27LdoYva
k3MMcm6OcTGCec9BEVuLqhn7s+Ew/AzyplPaWOOXObH6a+qKJJj9X0zXOLv6ulIu
uKD2cgyej1F93c96jTSyk96QOuAC59JGp1sWJVlsrBtVKwX4DcloL+rYsjZmMk2q
3sTW7wg0y1ubDcQwnLj1iYt4ZF3IgwzcXv1cVolDOQiUmtMOoN6HxlcwvBVhPUwI
/EO7+RgqSZ2iYlkQSyMazo84addJ4b9qiBju4Z+/H5X+ZnUWqSHQ5iEoXj3kDshy
2ZDCHegHy/jXxiqNE5AEpKABvGTFoza1lslGxfGRNfJjhGUX0UbxFa94lKFth0x9
aVFHuKN7AZxjxrm/xh7/NQfy6dYRwqU3/oBP62+DV8obwSl5YrGPaM6SnSVRkztr
dNHvQstJxgoBrEd9FV/+X5P5Wf3QgO1gsl2I0W7VNL9CcatkiDuhvZjQYBxVIRfM
xbVxZTblLGgraqWA7RXAUqWHbY8cJ/x5lYxqWzP6qrEz88x2LUqjr1xZpFL7mZZE
XOOotc2VXTekCvV26A0+n4qci5+PVEyNl+Rv/j0v3hOkeX6The+9fw7FyfieI+bc
y5latejSllFp89iMHl5f+e9rGlNKmuiK7gsodliN2KJOVa05jPcWMRZY58sKqp7S
sj98iX1DQPqqPgIOaWUAn+sSwwFREuWMVxBSk2F8RQpzXeJOFN2WNvrG1X5MoTCH
7cPNgOt18c5sknuOIBMH7h/0TYAFvleo6sqSiCys3qsfPiuUbKRhBU6Nz10JmDVv
/66mDFvXsEC6t1WIpQPXBtpWFA7iktOVcWX/GgSoggXG4n2bEz+DUHLt7hBwqS+S
K/uhTS0ASwaaOcAN9WDbw5ua0uJbS94FwHwDtSAQBOdMRnWanlrMsNK2AooURoCT
Y/bMVJA6boCt27zFvppvPqsXFOx8j2y8uROqsAO265ZgPKAnScWqDwmoUXCwgCNX
U3Hx7ECEfHOHcpvcMhNt9Z8dDgI4HFLAURdjHGIzzgQQ+UAUc+mLE5mmNPsvfko1
USTu1bRPBQxkkvXKYuxfcbV9pCBmCcbrI8rdcxYUkQM25eZnITUWFRDssl9Rz0BY
vV4q4MpDQM9nK8DNBk6PS6KAu6/lmsLSBuQ74rcYkigs9QPbZQ5grDov+L2wca+h
Fbmpczn+Z0dBYX2zaNHxi9nJ6zGxCY3IFGhlMLsiVKIu81uy9B+2A/Xh1JoT1vj2
CUtGF3VSD6cHkjJAJEAdJiWuU+Zd5PynzMk/uJQnv2jVv42VK6GBEPvS1ZFCjml2
ykQF8AemZTrN7ELBrzgzuNrvRosH2Mbf1Qr5YujKiY0OLq1Nh2kDSUx57B6q/UAt
4xk83ROzWajXZJ0sdpuZSH1qo47D4A1VUlPXJMZVe1ehBPmuE0Vy6obcwqKR80Fl
AY9LqHnWhYTeO+o0A9wfQ4GkwB8/603qN8dN/MNruUaVBXS3BH8B1Xbb4s9lRL5C
9lr4jxx53G9JmUzEi9ppD5SBfdCDVd4gsFMNuyqWPB7VhvxwHO/UtSe6nRsyv8bD
YRclfFF+EXuxyYC4xvKE5bh/DM5fVgcmMqT8ngc9I95creJhaJYdiwbv8vqdyq74
yWFNNNnqFxUl5BYREUxKPVRPe8d9k+Vixmbw8Q09wyk96CtCmQYC0/5q6+SPNWc/
gDPM5oLBrrUyCnDudjjUVcF85KbcPXnloFRcIqCfhNTwgfWTjRyeCuFtnGeG27hn
99jaBDDqtB808Y1nEpmUWRetFc8Zkj/IW6XnIT2WYr02PGS5M2N7QYUQ7ni53Egk
WfASgtfBhQWl3L/J5LMGYt2UIYJmQBbSIDkmTntWOTeAv0B1ij2YSyKjINGv/ZPA
rmLvcRrmeGM4WiSParDGB2bAAeVjKa3bzboIk0APmdNI3wVacPhQ6dJnQsVoHtr1
IXsxvt/zVc8vUWVXj/2ito2B2Ncac0rVQuSV+T94nMazgLKfS/Vu9UmgYpSBwvfu
uITnVV+n7GGitEmJa0M6L/9nIws7u2HJ/CHtT7uEevKPBWjG7PHsUyWBNPxBeDK4
qZvxTANhWkxJCudHEiUvPrFVPHq52MjCiBL8smCeeK8r3dB0GkcCrq/xUoMG3o49
UyX1mPT50AWzoXvdDaxo1UmfJqDft6E9hukXU2TADO/LTOcM4Bdmpo822IxylSjh
3C/aiUX9h9XwpaXeHwp+MNZKryeg2ig7FFO2YCvhZNs1aQHy3ho6xT0c0XvVws+6
U7z6v+u0xse1Xa668H7Dxfyx/HrUCBRgcQKYiK3ETU+N1R6Ec4+WShJH69zpzD34
e6DxDLrtBGLIxdq2JDUPC8E+1kv506+IM6h32vplJIVwQs2ua173kPXb9hppKBAh
6W4N4lAhmAxBoEEHCFAcEuxA6+k3EKTYkEr5c4EW7ll7VT8GzHbWpMYOi9MZWLDQ
lb1kP0BxfXqdenfdOhYdoQZqjkAoJTkWIW9lJ044dkQqEPFE+9kI+Z6KEQvRWg1O
SwerZjRQ/PakjNGyzwCHO59mS1l7JO2YXHAQtIeMFYN+CZJujRpNE3Q7JuRB/j0F
iQKwccA6FjQFdIDHElA2hMJ9saUFqqKc70XK2XTJ8HwP/vf/mbkQaOwVI51Qa7LT
iYTgR+B6IFarzxKgA+Ubg2Tsrm2PUxfCDeWLFy6KOWoiX+Rn+z6GlshUeXstyszy
P4kQ/8/JQ1UWoLz0YtAkq1qJZcP7kc6TsAOczQcEH6PcdLaHXpKNFKk0w6kcXiTk
B9W4Clq4z1T2SdsT7v0kVJL1o1pV5fScz7vBA95GDkhcG+GKEbYkBy38eXIaHOSo
O1IbKklsPSS+dtw1UxJEdkWRzx4MjZ71dNjoWErmEEwDodhSD2MlnAo9eUeudcvW
rFRUnH+ojTyITw0Njtr/Mt49ugGtwwi4lRlZcuT+dGQAh0YfknzWFZ/2ANBjyprk
yyehTTGgFbOLdlpYcHr0keKgjI3yrGtD6dg3MZUSd3n3b9q06NgtaiM/E+l5UqYk
Movet+OxA3xArh16PDKPLESyKMCUf2Inek3lbmX1aZBpJ7M7m8aV7/T3PR1in6Dy
Ns4vLsVd6YPoOUBYJf6+0rTS8ERbki0dXIyuOV7coqS87HMh0QF+dIUJBcIiqcIT
vn34iOh1i1UoBTCkLnrFgfDtWLqMR9+q9uC8pGsnrLCrzmpRRTO7MYnagZT1+Jye
mgh62JF45kNmdOSTEV5pQvWYv5YmJLuRpBFJ9p74vn/T51Ac6aj7lCZMaVh+ymOP
zXCCrOt9SdU35v4/xo1PPP+srL5XYgoS18jhjuKI5i0Wbmap/PsUG2+0rKRIVdTz
LJ5WiabSB/+qoFfjpaO/YmWJsMig8AHL3CMZNgWQj4W/F/zn/dtloWRLE1AJXvOR
/+LCnXtDXI6114jwQoIK9vr/iOwNXGbCWnXjujiG79oBOJMJVi3TPZ/7GDdH0YB8
H5nMhzrLTTmtOvOn/lWfAjVMol8F+VZP1Ge+2EUNN89K59H1GzslwGRmazijguxu
XUX79hWOOdvhWsbQU0omjLwDW+D/bPBq3QnP6jMunn6USuMbLhJCX47gFJl+NxCD
UYxCQExrxzEoZloE1wT29osB1ZLW88dBaXQ7qGFPyhxwmCDfNv5V8tMJ7BwUGh71
bs0Ejn6dDNW9cR0+khqO/yIMs/Wbyq/Ckx2SDfe7IN23b1rvAwu0y4SpYWVeGKZO
MFg7+nC0EXCEdkIJiNGNa5k1qvmGDHkUhQBixSGMIngwouvLuNu2eSofL4WsjPbQ
mRZtuX8+iOt3u+OO/epu8GDxmh93YEKY7LgeMnUq0oV32C38MDWphg7TIZz6FvdH
26qbBD7UnOS+IyL6AdEKS09x0D/Cuz3gyxklydbM8xXEdjy4HzOcR3A4gebthsHC
MKT2nNEms4bE223BDVWP9Ic+pkLUI0v9HrGAVXmE6uKStO1yfBX+bgo6JYzxOAnx
KtkJuppk1JisAkgyvFcc4yfOBYWxWb/XoI4fNCyhhsA1TOCcyZZjHJPYM6HRH8Wp
sapWxY1mnnXyGXQMc04gbLLH4mq+OHetSDNOi0F71imHeuq4BHiClG99WnA6l+rP
J2d2dHc1db1huj7R8/PiLj152jyDiz9aMZMMkTAOp40dtOS5kNpWQc+DhaSXR/zN
EwuUreXUkgFp8bhcOpnxBa67tED+q+v6WfFg7wF648tcbw6OorLU41mqiJ3Xihgo
R0I3hVqezAXuHo7urGu+OMMoVI7diNd1a6y8sgoejMZZ79t0a0IK7TMY31i8IrjM
pY8Jl3x8YzMSM6cpeVjEtF0A8aBd/oT/tlPfwjIT/c2gAwjMuB6PWbtUXv1LiXkH
lowPuaqUubwWUFecbdMyq2nFaRLh7XkO0txv/pvDH4vdbbk8CYATLorWm43rV/QG
5OOlhTVllGP8vp6gpbAi/ncfMWkzEOOTFvQMyXWDgbF5W1QSrlDE63XlT9n9pya7
l5b/IMIdrugkTkB36OfHXgl6+BQqCYHG482QWybA6IcOY0uM8Jac4DT5I71pZNaJ
C6xdjx7btFYpl24hTDGTSzlQ7NoQbNPPilHdB567dgOsP/CcBRtlDfZagBou23O9
0vDKAzy/7xWRqVUN3igG7wDptvJeMFOJ7rHkQpv2w4ySk834nRi3wdFmOLb+N5PA
FtJARj3BbOTHf8BqxkTR59kiG4UaCSqgHjln/HkHSIR7KKuuz9zhdqIZREfxiJb4
KRJOVSCR37NmD4bMNr+/NtKwMsWThY574uVZv/KwGJOF9zlAVVyFxr9tVifW6W1O
g9M0ulq6RQhOYWw7PL8gcb50+142wBby4c/DTSjVU/4EOEkManVucZEatLq+DX9S
qEEKBlE+3DZ88iepxHa31UFc79t7lF9wC2qmlC8A/bv/JV+0SfBMhR+rRBd+I0CP
ZjBUiF5xWIp7x0JoH1iLJiNXXfapfPJ/7Sl5gsfE2sPqzkHYLTjsb2tkWYGEMBEZ
fkCqiMSUS8bBd5V/qcoS1ez+zQEyu8XPINm5tYut6hloTqC6T+KDRV3MuYZPdcS0
wcI5hmpoAHoBkM7r06ZYKjjGWvsC/qsB17ReWXIj4wDJT585HFXTItyhzvPVai4h
ziJFAOiSCLF5UYHkQXdf1dHe4EpRF4SkwB1u3/Mp6/sU1ZDMBGoN4E8d2AqjcOkq
FozVSQzwdTKVT1EPREmoZPgzA/9ZghBfkuNS2YmEtB5neel2j9E032URJP1e814X
T4QBk6xj0L7H58cNWvn0tRrko942NTnuaiYSQWPyUG9BWba/10/rfoPUaPYXqIjB
bq4tLVNOWDBkuK2AfiajkvzmS4B0kmtlXc/w7MnXm3Zbu2tONnx5VB5GelmcLWgO
nd5pf3Vjj9EiT/Q/9eqHdy49izvnx8RwB254v3A6RWvu4oWWtP9abKvPBZIMcTwI
zdZQgQRHZWRX0pB/EAvfgROfVvsPzuXW2aKlAtScVUmHgub0D/yY12ssJSpqDEO2
KWbppFyNE55GXFG6GPzz7MPsRyWDGs84xA9C5tYkU+vMgO8EN5lopZThn3mD7H9I
Fil8P4yj2Omj2j67d3IpbHxfcCqw/kaHYRxsS/d+jIDMm74R/JNRSllUP/0UvCF4
FX1jrKGSJofoZujvqOmdYkRkz6UwhuHKTi23Icbam3wjGUdS+puCPJHPAaSWcWVr
ZSrwMiOMiWvEZ+5ohzoVRNW8/oMkl8rBL9lTsl92JUqGcJtjiWyAg2ZuSGlRJl1f
Hzx5uj2A3PxUXotwucd1ofb+gHHnJRXcOn2X2qdKU+65fO8+hEgEh072FXhNjsWb
rKG2O6PK5ZumFrNUoJxkdiKTtOAJkm2Qv2pZ7W3NXwo6Uo/1RSIgUEs2JwWicL/m
2rTYsgjxTJcFIOQVpr6yqtVM4STyQenWvTalLO4XWVEEnLMUXvZQ3VGMmKYrIlR/
bhBgQkDk+78mkbTMWQ4GHF6h6xJvzSLgMoKnokSxhK/XOZfFeIb1hKg4KNhY7ukP
UHyMabXJn5XrHqRAYRZMaYYML5WkkHzxeLhl6C2qFoLc4XQjFvzW6bRNkSqtvKSV
XrZv1NDUSIBZONNB99sy8xkx6IirF73ojlToFJsGLXgfCKI6vQX8wpeZ0pTAk6yC
6c7XztqqN+sHwC0ohahFxZ32U8Wifj3z9xcZ2iP26mNS+GWO3J+BYvdAVspEXkLj
KvfYaGeJtI/HBthWROwCXim+4JbneB1EeOYHp4KiPH5n/Z/ctUUGXkcG7qDaxhoP
+966XxtqvnQJiSmrTxPUSKpTDaHRvccVgEAm+AkIa6tPY6n+kxpe6euQ6cLxNpdC
k6EuGpf21eJdx3GAl4pPe8wAiyspZvbgXseGhZA+cRh6YRk7Ylfs/0jIMlrUbBCq
UQRX0+0hxym8cAS4dfmLBarAODWsfrDXzDINpBX0qHxsl99DMv2Tvur1EyMu0eLZ
5xQLOAjcZ/A8txSPn7Lxxtm6gMQ/qLEOIonuLOMjgCkSNNmy/N1CmgnGN08nCPll
ndr2Tp6TkiIc1fDpffjNsJmWW1wo/c5ZXZcIgaor7Hn4O2bfq2ZJ6FdsThym6zPB
qBtLWPRoEVlINAnDMKltaaZ7jTG77agPOOjvydcdi/NAI6jjjJd+A1gDCg4DTSFj
uO1YU890vNj4Dwq/Qmqvul4oscVpGXaMOUnaCRux61WCh/rKh37VlruwIvGvCNEu
FboGiF1CB6xroKZLdBwdz/84d6WyLh1NYEH/WN4SEfgpFL2o+v+E2eq9y/SkqqSx
4yP6foSGbvD4U62I1ZHoLuZJZs+ox+a+nPEPPIzdZWiwHC1t5BxnC/dHGQZBMBC/
wZtYOHaN6Ps/P4sRd/FICJrsI4Clfo7otOvcxbqkFdxm2EKrlrZEl56gJJpft0KX
rBiOuL0T8N5IEomHOvolIz5P1wWyQNJZD/4iBa7Y5iU6VvAFVSHOMnsReGM7996C
w8KOwjLkm1DK0OmijXe+U6Wd562HRKCAjhjxZbGI5g/XN1tyYs7wxYkzzNIUSL4t
nB6RpHvn8kbqq2g/X/p4nwDc1b65ZWkGVoLsKbHJLgfx1uukijI1UAW6aaxd7+CJ
auji34IPMu2tQcVE21OS2jTqFaWo2OlLMzQexmpm+DKITJ9XKQIfA0JWO57Ggf/+
KE+LYb37AP8ra8n09RSLLcBvWpd3T+zrAhs7qkKVifiQiNwYWoW1787D5zRHHS9M
Pq6YxAW26f7+czJ/G5GaU19iU7kySePRc3DsF7iJKq6mE159o7ncT21uVqjUxJQ+
9EQ138TH9xS+XoAQ4EC6tGZKXb01yR36fLq7TgLun6waBffk4bP918YChH2W+TGG
S7bkmt5/5OslDJY+Tfne3IC4ePsTLEEflzI5sGY84Mx1g/xOGZy9arQqnHm63WPm
9aBa5ccwKwcGSHFRyoUVMt5MNpDkChRZxxtNUWhaVjJaFwMxAFMA8k5rj6fRlAIV
TgMwI5qSthGwVD0+cs+xx4O/9MBBsA6P28LEd8ks2XEfJDnDJs2vHUyn3AD4q5a5
fQmGm3xxSR6xAoWe9sOyc5yGGdwkWJKtoK7RiZA+RXccL+DuJNSQoLb+/bLWyE2L
dzaRn7/7I1+LSnxJRQPeuZDPGYUvIJsKz5Oz58RZklIvN+/HP302ofqB7fQDZIHU
eln+8Mhu2YNL7GctSMgUhs8j1oSXp6lc7LQhc9m5pV1VUiiUGEZDo/fXcCFfupCL
yhYUPhtzjOqcQJaz/7/yc+MglbYRM+MwHY42ktKqtJiREexySK3Gp5PYKVxrW+mz
L+S2nRwfI+XZcEYtQkJD+i9PFLNB1Wg3AttrRds5oy/8mBWye8ZOWf5kko9jeMwJ
cJUXmVk1uLGGBryUghTckFJnZqFObxBhwRWlqBcEzl0l0FVz+P7qJ9sT4xbCcGan
40Ubu9W6JoURceip7ntB3lHMeuoqoab2Bif2q1+CaNlb1/MxXlaXIkyOCB7bCNOF
laDvycG6ZIiCT8uD0UNOeIKny7g+ZRIX5emiZa4aonIGWYafnWSyO2K5V8AOVYuE
Ku2PGNRYDhTyRdUQxxEwZQThfibpGzy5WMicXAh2dq8s+Pc8vrTomXgF8RAFyFwn
vaP2CRozpAoE+/AMhotzyDgbq9QvWvGTsKL7glSQTgkYsJwY74vzTsCYYa2iQQm/
VDmK2glu+XY9CL8HFsILpzAgVSo6ZPSpV0MIvs0BI63oFHxKI9bdeXZBYCVlnqqL
yojYm3yQfc63UEeHPxjV0lQQolPP1moo+YRfUyndY5zGlf7DnAj9CICjPNWOZNY9
+KKd6pebsnuyj4pKc6pVvkdNQ0NHJLkWubrWVvkSDpwnlOM1gEqcddJ/l0O9X8fY
P+fcs6cIT4Kg0Ktn6mDdVoQHrJ5B3dGe7PnYaigKWRSD+A5PV+zxPT8YVzpXCDmW
DsyZtIZPMOqkjP/6XK39mTPhLXAuiekF07/v8+tI1AiGy+sajPlueLWxiMW2wjqC
hx8HdVaZrlzob389CsS3ReeVTE//249I2Vbo8UVosVIaCaOXVBGPNxkWe2lOCI3i
Oj2mfzR7KM397I9wDBS2QjZ5t7TT6Vh8Wn2Ya8cLHGgfczWaE9I95pg08Xl8989n
+HmJ+awV/fhHFwEoSY1UoD0b1q2bP93Apb/zGq3246QvPC0Lv+9NtnmSKsvSVBxU
kYsCTWdbsdTFrDL2PTsZXwg2zhHM5ufH3XUWbgy8xwqViibtt8tIFZ7uZW3U1zt4
ZKXd60F9AAUS7gIjxTMyzeBstcd/z5hY/0q0orIDyktr9XW+1U0rvLSwLW8EfCBn
yX3EWWreWV6ZJtHx9Nd0tC7CmjqXAhy9REoZvKH3lrzerNme+4RRLlmaQ2w2MwIl
Vi2PLtzsj1VR/QrV3nkj1nLRkm8i+VXsS1bCltVem7/XKKEnTSQtkJeu0GHfAe1p
8l3yX1/2WVco5leDqJNMUWD/wmHo21RKxuBuDsMXIA2bMkkOuB8uaOhcezbWNMzF
KGfHRWVeoMZHiH+xhD6NPWRUDumMnhVOYTbR/T1mFognPhrEq0yt+EQQ7Rsahz6G
BUeruOcZERbkyxhMistIvNIHyQOpR7MKddkXAYBSgcpRv0XF95XpIxb/U78DgFVe
0ZydfnEFQDaGv29uR0ikl3GavUUUrbvsSbz9RjrC1QZ0kVhfZCY7tjYddkg/nQ1L
uQHfV8WL1WPYXDtgBJJpbJHopSEPIFXe3beB1xDM9H4rVN5//B3+85/iYM40iJts
fCd86YzJH7GF26VyMFhp6UeaB6pjh8KOTcmZloewaYITRb+eIGefRhzMLZ88JhoK
IM3Gw7edlOZluZw3THc/YzRW5HKqq3lcg4GsQSp05MKcFUuuFByNJwcuAj7F6+OX
zA1G6CuVDOvl5zMOihEtyubu3LrWQ3Hff+JMpGswV6zL0YvacSfsjtEQdbnHptx5
8NnBhQj+MdlyeGiuscOGtdSOFXUx0tCoNHFzaUc65V/FF/q0K9GZIWoznXDh8Nfi
WbXD5xCRWKVp/z0UnxF92EiNCtngjdXYneULuOoUUe1ZsCC7dl9L44dx2DFwasMJ
sYviqNZWAuorjL+EesAw/Cso5pGIzO7AV0ONDdN9ndcJ5snUNwL9Hone3NoAt/iI
TUGt94Br5bd/3nkinHzBiQ29SmK66GAhUf0xtzG0v0mRDPKT6PCpkCpVd7jJkYG1
e3/VttfoOokh80+G3Q5NlXJz2s/KW/LDR7oR+uOKsRtlf1TZ6cy9gCd8ZVebgFjT
Yk5tKcjCBoX4ZX/a4VHR8BCLN2JfFpiQ/r2xyQH6i9ajmg7k3P4NjCgZZQjcqGnX
9tPWASqG9fX3uetz/dX45RP2VS/YVBScbEiaO9i59fSIOwih3CZCXr+5xbgLYRM9
f4cJg8McpQBuoA4MeQKUCtACLGJgoz46YCZFiezpqcpcv4tfwsURJ5q86hajQLfv
3LTbf98WUlhEgLudx6AEgsTIutNLe7LTy6rdbLl9R6LYcBgf3i7iI7N5vr/+tHdx
QtoF1qR4/uKZCOjMzYmuQPwipQOf9c4EzJ82zpSST+4V8l/m137daTLg2jEYVmXB
AuGmYosk681VL7Mzsl5DKEa+cRwIJV9OVri42smLwit7Ikzc6IgsTk0WghEWznkf
L6f4AGGjk5d5x/TYa2UY4Lu8gWkYziENPbWKTg9fx8YCOnrXTO607oItcceShlh0
LOIQkN5BYmtK1hlakpYmdZM8dpqcpWIngx0dRaQGyAmEbkwDgqPvh3R77OicyCrx
fp6S/1CUH2XNo4S/406f8U1sh+w1ylTtOYOrhF+dvzvXmiuCW0g81mC1ytFrW1oB
HIHJnw7QGU/RdlZNnPdQbsWbgchIJO0sZ6nqDyt5+LRYS2uH1rMZi6SUsbVU0VLl
LUndgVZPdmvpF5r6FgQqEb2y+qWzjP3py06Vq+rVu86sQ3I/L0YAbbBqGtUEIRLl
v5bvOM5ShftjZKom3qb9oA03cebj5sUguy8TuhQnVxU/L1ZojF7KasWVzAqUIFaq
ZdIzrMfYfXsq6mjOnqhxq6bM0t+u6KygkRZz698wMBciHzb9SMclJTGv7iZjeyam
D8ZnroUZGIaN71fuCE2DJnDVtRSuNeeXOaLJ2odffGx+qstgdGkpC4jWHIi/2lAs
nErEdsmttljJWc71LlnpjnhSlEdJYL4vFjg9962AKqoiA0fbuHMno3R+vzwgFi2Q
Oj4c8+2M3tq+hjGgG/JD/2anmzPhSu+Wz+M4OKl/0OakyudWPvRF85ess3j4IP5F
wdLCeyWWMYYj+5CalFORHlKffxd+l5fS9iPSkr9M5EjSISNgX4y3KCKVbfyEjL/T
SrfQuiemmYClW6qWWanCXE9VG8WdvWcv8FA1QJWAt8mxvNrojnuFlrx7wRY2uJ40
CQ+xEtZjTWB1yFRemz8ziA5YenYb8rGrHhbR1nBzE9x+cmic2fwgeL1QYJe3U/uG
9EJJmKMiWW/EuGAVx4hi9BzPwRnAemSZ+Xh44DjRWU8/axZHnC0eUOvpZ5jhzZ8n
NhL1T5CYxFlBZUoMnjrWmcNTbuYvDes2XxrWgzW4znI5uczHIxBeb4K6I1NXNlZ6
EmeovJjyeChBQk00M9Q7Yz1bpokRUtIpZfdytCYXypQcscKCU0xnP+ulQVqFP32s
cpG9bXl4ZtfCIHeWPv6lILD0UmB+GU9F2AaZcTgYtOgPher7oTtepWqPiAobNtgc
Awh12WiFjBcWS5Q4TlNWKJMiYt4hDF/0sYHZkYvzl0z0XV0e69ayCc2Da5kM5rMI
ar0A4v++t07Hk2qrmmIBy7hpTDBcc/jgXPHs+sfc3uly8ttXLwsEx0uzaPCQzD7q
awrWcjHGFH0r2UfRpQueW/yZtZcfF4uTMrDX46LV66USgr6V/rpQiWuRnet3yemC
cvZty/TtienHB7qOiqW01ncuSeff8ls/AEsmO/RFzHbKLtQEUX3KHdp5ZAsUzU0M
/5yyKlMfMBgXKHMloySAfj4G0aY9EGR5MzGFDo2laJKYIA1OoDvaRyXvO6unoHBK
AbXltu8bMOvWEFo5hCkt6RF8qKPpBAxerfX8zU3+4ldOhRVg05QEXKo+SrtrWG8E
WEEhar+C5JpGKytsy/PYLt4878KXOwZA7JaAZMYiof2o8fdSJMLyRJcab+Yn3WgI
jv9fg5pfeoIoNQOtvpaVajMjdicPnmSQe0UGBJv4F0OIbuaI8sz7XsIJoUnsFTx+
JAa90RrPUwjuEa4AuScqabzy6kIPOYcpGOPH0RUMxIBJPqVvKSy5eQDu8WRYo0Zm
by9HbWr/8Z+j9fZssUTki6sEJcBa8Qh0YPzJ8/Z1OOKbxnOIeyH5P+v6UjuhtSKj
9KMXtxyI7EVxHZut4UdHqwMOoj3sMGrDjY6von+METqewsIF6RdO335/r9kyyvVD
ST1PCzW/skoNtbvgC5MRUuoHm8/bqSFjnqheZAvB0YvWIFABxu6bOXph26aLmg1y
/vOjogjz5Qd86ymcJBGyQf0+m10SmNEH8zp5E7CfOxAhSftqhZgoNO8vMvoS5PIs
jDiy6dDdYrgCTUaHY4ZacgdHMXFvYYn6zEn4UUrtRAtjFKjfv6DO+xrfQ3bFMXGQ
Lny0fE5zTtFqVCsljsch0daicup12YAGqKdk/3YA1t4gutJlWDOPh07rgxeZJn7D
LLDJfSrBjmhXx3wqIXUCWXr7av7PO7GkLllU0a5YRKPd5BMbZpkXpViXLQecvzWW
EgAkPvB1WdRItnCA96UdL2O0JNAQVB6dfVBJbQphOSSkSirgHwAJiMScvPIMFBGd
XHPlTVjdCCSluNmgPmZNmknCGL0gpPDzsxNS5SJeARvDiuJZKsPAuV9K35Novxv2
64lzcLIa4wHVkAMcHasJ7pC8fgsroPxAcCV1CoBoUBXT9/okJkuo6CS7NOCkMYqC
s4CTl6juIt1nR5ml1sPY9T5WGrcaToDiCWA1YLvdvx2BwwnByoB5P2WCWUVU7lfH
Q/bJbd1mU250CI9jgMY5LY6O/PHix1XuUq/au49leepvqXP3O0rH7+msr8sB6ZkY
XF+FL3TA7bVSCzKloJ0SQB2BEojHt/psTwehQ00TMoLh2a+7CtJhWnAFRjKfQfE6
bpACygvl1fcmSkoLxf5l4/aI2PY4cJAGapBAG7lk9H3qwcL+g3GVfQv1f/JiAcCC
ByYCgccrQ81zK5rgdaU+2ds0WwbMCY0EnIhC7lVYHpKZK1XgN7Wa/SDwkR+gV+Dr
uI5tELkbibQYs87d9C+ilJUZUa8p0hqo4DwzOBROkO0WlHp+fxYI+SalFrbnB3Pr
l03bLiU6WUMsqFcHE6vqlsIOYcsts6DoNqxBynQjMxxvKQeMH5UOgGQVAlTvnB+Q
wQOOB+PILLsnCVh3+RuRY7tHRC6N39s6PB2TFzGu0r95StyjuUnlXUdsjiZ9nEyy
PEhPIyzyBSCLcraRgnneBH9WD1BIPG2BtSfmvS7E8vLx3Mj+gpRHnkQpQfUwvxpc
7uKYp8KPy2KQIJtHR9gqt1gkFWENHbNPhJgT6ew7HakSOdxS9kJzr6ghgRaFU23Y
m4PW+IL69/mMhVOsDhdQ/Vgdwh2vgnB8vnZTMYUAw4bqrX6LLm0wDi7Kqc0WyrvO
dsnwT03pcVJyueE9IckL1a7S+Y2UxvNU0eqMjVBBIGtrCGsw5fn4TOjetTmakaMy
AXcZGEzX9JYohUzDfW3oeTN0DT2fzRpaX+lCskScJtqbiB1KyROUi0XqgECnBkmc
yaAVzhbbFb2/QtQ8qAFTKx/47Bt69Y8ntmKLw7B4xUWKSDgOxlNC9EOts+t/KDW/
4jXGc22KWbExfBvaY7TNvGS77iOLpO8kws32MSnlajpRGquKMrhCj27tgQOC+r/o
5/OLbx8daNaR5BChK916JTYNrOEHRFmB1+gRMMRT9QXHXVFbsAY67WqIpHwW2pi9
fBMZatan9MyO7+1NFxYO+FWJRDHZEKpkVM2mOelzkGU7uBi6csRUemUxQYP15cDN
su3x3Inx9IsWr3lgAMmFiCegLvelX7m2QlOjr7RcHnfxwiw3/wgMKC3Cg0XQguDk
onNQkZJdKYFC5AAPKUbkbS4RL63S25Q6r6CXfeCWkvOmf4h3MFYgrxPbfH8n7Xv5
j2iemsQr12CtU4uD5K1kzZbzt3ltPTBKKVkN/yoRit2Ol903HpqUNSfC9TBjiKTW
wQsUcq/slFAYdB5OSfE7tbVjK5QzY7DZPjjGYLC668Led8/BOJdw1bggfIe9v5Hh
vmcT0N30Xuu/3JxdBRaeQCIcg0PHGq4rGOe45OxWW/a5Pa2O8lnQ1gP5WsFfd0vK
P/wQxf+4ZVcoKCOkl5KtalCBmzAVEjGPis93wCrNBwDSrlSAXfhkOr7ePJutGul3
KIyy/0FPwqV8+atpQO2vNf93dG215eW2nRAYzQSbchLRvJ4KuiR77ffAY/5mVkGQ
YqtapASMI4kvX/bD94oGxMq3BXySmPwouvOYMox2Iar/2xX+EDNJ8zXxKdsuINr4
bsXyr6D0VlYIdbRLi+zgOkHvf/E6YTLeOTlv38g9TaXdnBlSJtgt6GK7kOjjKazx
XeZgj19coYRf15ejZZNufMpZZEQQcXBf4Mb5h8k47hDOubJEKHd6qU+gn8TN5Fo1
yqtE0aOBAcXzLnCC3oJoiQ6y4DXywvfgFlukXopxU4gO1LN+AA0wwDtymsiVdAyo
R44EyVHFdzEPOjxKgvQxteBIUF8ArM0jVUqE3r4ar/LAwSBSXPAUpwQBCp042wF0
f8xmc80QLENn6ldN2RgKl1264pmql1rtNd3eO7RzjzPNeyhraVcW2fMbeSysTSVy
1CqZs9GpG1tlOZ6Kal7q31wvWqBQclqC2dm8NSI/8yJ0tAcqi+8F0UavvAcsgH4v
JhAY2NSDMuw5/kq0UfWsc1aogP9WFqjRT6S7KC9n+aCXN2Ps0cvQ2Z/YNd1Zy1Hv
N08d1qB60B4M6x6RkR0ubgCfN8K+6cVdyEIZTX+uQqozOJPCw3YJ3eSSr2Mj6IDv
u4y035FWivoMXCu04ferUR66nyOsp/xdGcRoh1mal+5YrH4jRdHa+E6Edhff/OyK
xVYk+HHanGMIhFQXuFplRIRU8XP5F2/eFBUu1mN9l8oVQH7BNhlUcUPhZbgr533i
dzP3s9Yj5srZyUOjCsaTsuYxmPCQGMGruXM+4k8piHUm5z8MKGgaj4FUSxHEkZYc
EXXBFJgO2Tb5csy54hB/M9R4zPxa5KQkVgyMEVzhA55cqy0M3pyf1OhyuBzKpf0G
e+Hx/tfYvC1AdbojCLU1hjoFBNq4lr9KAD0pIBNJ4Q2CoGIcTjBl37fylc7N1NHk
I4eJDXgTJ5Y5D3NrDy3ABWj98h27LoWKNutNiRlS816XcvFq/jznPKg/PjiBxDPS
c/aOXGV0HIEBdhdWgWAvACXJAJsP0B9iHbnv0XkmPvFUY11c6CCyjNDg/Esz8Mal
PpSculvO3lxkvF5VICK+W1Do5dC2Ejk0fZkCAUe/dzE3FXGCSF089uIyFHg3tl9V
R7e2h7DoueB0d/nMRUJ1lXP6TrjX9qNRawMCvxAT8h8Uwa5Ohlh0snxJ+1ZvroFt
6eHZ9xONhcXhR1m+k+fXSJFHQMWgpRd+8qvKW8ZaAKJIS+FU9tJqjUCfQ20vp04h
LHr8ByT27boO5KrHrhDtk4U/TqAN/QV09XmqmE4W0JIZMOvvaSoTJHmVegvgy8Ht
fMZ9qbUQC2qr2ny9nEWef9CeVH2QWaNZI49oFvw4rVx74u8jb6fWIvchrcET+RIP
I7ZM5dM6Mo0RjTJNQciQzi2uG350MCcziQsaG1aS0z8INc3pUs154eSupwP5NYzO
EpKtzdHNhCXEt7/BypKpqwKFMR55N0jnI/txbnTfag16G7iLx5XA4u5upd3agbGo
fQqJdcMBYQcJDju6w2CL7Mz+bcoXp/w9rGUZ3uCmkNLXxW4mxHTUO6nQFWEww8T0
SLIwVGomL9T04le9V5Fa6VhsyLcBxf+lS9/tzMdPDctVnPACiKa8D53hHULfNLIK
62t98aEJTgcvCFlAQByW342J31lA7mBgwtZpMNC18iP7jvvO6CBlfY7QvDk/8/FM
LBlso6u2pLiWnY3+fgxWzjAN8Zf74tOr5m4Cwf8PGztLuLIWhFks0BV9m0smrjBE
/NE95Yk5VgsdH8xTMVYb3EXQHoIaPF4fFCOo+Tx2OgG2j6Zstc/ZMLf9EcFlXprt
UNeoNE8LpPlmKOmhxlNTHY6+SLH+IrACW0gWgu2N+faaoT5BukABKW8pCskhNV6a
rT4yZt42TQ6BKg4OD6fbfgEVmZxMobCsRJiIQHygXbNZlJYQEVClW4hqgzIG3iRU
AOrop2JBeShX4uNMyV7EE02Ux4FklAGQhsxf9gDZB7BaMTw9B1cWCOp0I4kPkqHZ
GPn5jzxbyaK23NPCPnzGJ6RUpVNhCtKEV01VXtD4tBhN8KuSsl6p41PPJrmmAtXF
Rvworyovicp6u2SWHJp9vVw8uyo0USmznZRJENYUNDUk9rNj1kKvVjxA+o1+hsyh
oprEDY/YrgeO0NcI2e5ZMaqhAQy/JNA/G38FVscPVv2HUkjB97SWBUqq5y1g+YP5
aF5CX01k/O9ELEBEv/9wCdpsEPvsKmQg7dqp+nzEDgIT5OlArdbkEeEG7C64miZQ
vJoO6hL7oVPlM8Q547s/zIqxx1+7G4gS1tYHNvvGocEh9QAKa3xrWoIlMCqBAeYs
Vk0W+JlHl6ousLpVutz1pekDPYYi4NCNgkA6EMNkPWBdnVqT/vNF5Qh63FhKuMzr
vQbeDD76bn7BeyWQUcpjn91yNHOl3KAlxzFmADnzhRSa0hL2XZn1XbAuc6ITG/Mt
47P7JZ90/PlGtdxbQPS9hUZzA4jXELwx6P4kC6QYg1heB8ZyjVjc6rA3cNIGWEa7
jCezBV+L9sPQRi00FPzlM9rov0KdP7mS+fayC07rrFzputB4EiQypPkeKtVNC8tX
47XEn4Z448Ud0YRfV//biVFcdRV5ySLxMudLkX81zJaAfAm3i+cGMvdHFQJppJzo
pOW3JnWjZphMZdpScx1oGfUdidJn+54xmeO4cEtcngQyBOtYKdc71Wz1Yi2j8Lwr
pvMXoKjDoQHuzjqN68hnaELf/N+/uJCWUWTFWtTGeQksFDoCecGqf5nXislmk5O4
fEDdiaHC+C1cB0Vf73aqplymGLkJ0g+gY+ulJ+frNn2hXDVbWzArH8QWqtWTJFij
SyV2QPIU4uyxAGCZgbouA11mhfIAaM9i/YaQhqILg4qxYFok7YsD5eiDfNP9yXRb
ow3XkN/vZJjLSYjqn5NPt6CQsiy1OYI/QkCbSR+vT+vXueyUZ+1l3Sbe3T9V3a1k
Cl+ldDChAvobHkDeTJIOrOgPISFRdZsHH9zmmutgLplBpgquuNmZznUPslL50Nya
kFvGir7ZgSZCYnlaClshkBr1XvCgtDeD+XbQax/k4QNc3w2dPQ9SYtAfnj85W1Ps
txTcyiCImSchm9QWDzbLxE1+tZvGif98ogFDJ9wqrH6wliEW4WdwZr95r66JKNQi
7k2aQ2HqNu7Wq8d4XJ/cuEWthYTdmZZSB4N3dfkStT/JZ5Br6IK01QnkMzxsJz8l
zbuaMm664/yWCSI1NcpTOCD+kjILwjuKrNWhXBd+f5Q3bR1QZdCL6IgOQhtNUeVq
1+h6XZ+tD59m9lOS8s+PUtNsE1hH+Hw3xqQBZ2JZ+RQZvEYqSDSPjkQcoamPPI8b
6wnja449A7jMv4tThTliXJnTCmiu0kNo69wX2OTGodOS1Xz0p/wOkRp1h8pW3TGZ
J1nqNkIbtNGZy2t5hrO9+AMg2rivaeGyXWrELIwQonVjmr19z1zPQTh73KXTBJqT
02ZXbK5JtqT/NrlL1QCTyeEo+nmwO6RDBkLL1mI2/g1jEOM0TGNF1z3TPCD9r45S
bRMcrO2xNM4M8EZozG2KL7FG8o26SscqFqQeMbYjWCHynAIRJAi0V5wBIQTrGNh8
cipxCmweyrasrJUe+IUs4KyZnpT+VKQOg2OEwz5ZwexaI/29MtblaAMtoczMtKd6
9VzY0BqtLytPFDgjplFcXaVhqvpH7NcaLVrHuyouPi7hWtUGmMj1MgAkVn87+VLu
a493sgD009dXFJoJjPJCnMbLAZSHgyZCYrHRrSgv51ijbFcX4/AhbVNPZbooZ96+
PLjyUnvpcvt3HZ+hj+YjjkD1FQTWT1AeoenZdioDhkNdo0Nv+WTvtyJ1HbiScBqm
38JIAzu3o5krL7od5wcq9zpiXDBNcfPADL1uSYeomaYmOLTROE0SJ+i9bgNSeB/j
xxtnCJ8ok0WPAahCtoIYQa1m83QAeUX6mSc+ZkceT9q5yHKOX59U9+d8faVzqrfn
B+1N3P4awOreCws7uUaHxu67uI92S9yNgm3j+uAEdI/qdDJYIaet9Kigmob/wmHV
PxxDUcvulvcmWYS7TDz4uc6xCTcf30RPrIQtama644NYwK0wggQ4v5JstjTJEeib
Qj1/9LaSu9lQIkCTF0CdPWoLKojvZzsU8aFW0GwJvv6TwkRIE7G9t40XHuRVLLD+
HQJF2AWnyVb/mNa0Dg1HPiUrKRviBU19rsMr/7wBvZDrDt+PqcwmYBcyhXF/8aiS
CU4MJsZw6FnucZ71tlLBUZC1C7Pe+8suMjGyFJZUEWTxljO3O4s8+BOJPcV+VmOY
9uw/bUCnWvLOKu6n27Lrz8hIG2FwTDuaqVAmWjN55/fIoZFii2cGSW5LKxXS3FFp
h7sJpDgh7oWXTgQGsGHoxJH4WZlkjsoJv7JaWN7SrijJvE3/+a8sXAHgqA7TWxiA
uQQXTvrMf6jQMTZoMP2ZxK8mYTjm3powMTulinZMdVispxhtfnwznjqYfe+gtlwo
Z6vvbEdGia1HD2AoqrXY7JWnsGbm1pmUUbWnagfcgOoQNkKZYm02UxEIXuPxVVZq
e7xSlG5z0x68fZjFCn1MdZwsEVp8U32YST1OxLxNJP3NiGnSpF/5tGCYpYFHunR2
k9uyN6mgHHWQ70BjD0o14SyHN8RBmZkTPOSBT5uz78bLioLSRqGGhn3JuH1NhSra
8otXGO1I01P1KAbc8psKEtaF29J9VqARUSQqpH07PAUrFOduqT0zAN3gcP+2T7LO
BhToAzI1QoPv6bbFtopkoDzu5Rgy9voDUfXtPsfsb7DuMacxl4RfbzsluFMubWxk
W4hNFRPg09wNOhHAHRGkHFS12XjZPSPQadPCWO6xF9UGOpxYT5WSZBLMx5SXDI49
hNXKq3YojnBCQDt2LxSjR0jURYkVC3izUREEUjy8Sx7ZxVK9leoaK9GwUOxnae55
8uMTVH0BOxG7gk6YpbQ5BXSB7/mVWr/a2+EQ5bPmnCUEAb9gZGFOzJiE2sSN+txw
A0QetjbmnYGtvp6uu2HqW3qykXw89u93+yYWNVXERH9a7wiWt8iU/HvsKnHQ+bag
B68Q7x9STFGz1hFv1mv9mB9Yji8bkBqU4Hzv9vJeYRz/fVOh6/Ll/tveISdC2d3Q
n/taZA1uu98vXLCrd8xEMPAB4x/nwfP1nVRQrz3OSCHUcNMBRWZixehisggruu9s
vWC9wSUnSmopPqQ5Rh7+bpLHXkdGrT++xdtaXXTjNCTmcIbhudkAeDd2sY2DBIFt
PAKBMeo/0CpDiL/zFBD34Y16gXtPsYXmZrnivodswm8yz90wsMPpWuftH6/z5r2L
TkImd1SOR44u8UcSGnTOkMe86R5d/5llDbqH8idDheYzlpT+gtuo+evrydL5FLlK
YA3sd36FAzW7G5zoEm4AhrBGiEkGDn4S2lamPksXBlq1UaBIu5GbYmW1MVBY7tUm
Z29iDKuGBkTvYiGR+nqHtzc67iNjAabyEXVLj9aXTnoyl1lL8sMXAM6zBlxVMTn4
1B+mtBPLPgzQUSi7i1+gU/Lgp9s/pHh1gw5sy0Km66uKfQsgh7QDZKBQ77Q/ir1Z
TTBYX6SjF6ZHc8P5r5Oz++rgj/6cnZQ9x1N0K0vrT/kWZOAEu5qw/Twaeckblc10
FukKKdJNlvRg674zqrIF7tehkGn6HhsE497AdBYOKmUGDuaQlHkpUnETDG3yBRTl
71ijYR3DrzEYqlh0gMu5DVycT4JIb7KYnzFzuT0yfRyHzFoBXkFLwkGkhQuo86NK
skGaDpQnCZqFdu9l8R3LOA+0enJ8AA3F9P1w6/8y7sgoYJUvzKieb28FFF0+eogA
9cwnL+skpVPziCjF30vS8VWjTLLHYBxoa0HVhx1HbpyWL6BSO4RAbof0ogvwhW2g
VGTjQ+snXuYzj0nTWfDbrTQCiqSpER33AR7nzlEHVjTxw/zDqrY1E34B476tMqLj
GU+u5CeJ3PrTW6LQXBTD0ftSrmH9n07omji76K392dVPdGmzn29bEl5khxTD36Ym
8iOjp0U1l/syagUD4w9iGPq/2vZHeMyEuYZdovOkyC9qwv8QVDZ6tJKtVIPSCEpn
RwPGvLuxAMtSw3j+P37QzQD1s0/zbfIH0i5pUW7Yd6f5rvHLAtvQaIeCWblWjat0
h+dkXxvhz2N6+DHrME1J8ERzDfeI6WZyHh0zr0+YU2bRciRa2xEXN/bXws3wYvcx
V9c+UO8f004XxZjcaslnKmF0xLY+0ptdTKwRO0QJOnFpBrLBGxh67w1A21KAucYH
yGGTBfYrv1KFrhd5A4fZ1RXuEdWEKK1KXINxf2zk3WzOKnmGmDBmwuoiRJ48XyP7
KuunWFMLgs06CDOGlpLDlMu7wMvn9OZYbf/ZZsvN1H1mlsNr8e0mcjeSnopBZB7J
stNfKqHK8x2T385nXf6LKbzKothTSO/RUb56XW4T5uRsoqCBgSJV75KuIZIdw09N
pFbEAd99azuj8M66V2+E4mSYJe+eIbSmaX3HVm7yStNunp0SO/ibNvqJpWGl0TuJ
GbR6sDehqFhdHWxnev6CIQOKkiKg3BtOkcbofNTdhA4tLslm8SrojG9rXguLcgs+
9oFj0CdHy1KcIlkh6Bb4uJw0nUIxtabjVdG5FRgEt0/qiRuqtgaamiV3vTtL1wGV
EQbhPk7xyhBmGTjxcXlBvkevlubnaJHrL7Z6gWZXE7S5ljf566OTPAfxHhn71vVA
+WF01Jed1Ssbzx+mBZ4q9MX4mIfzHYDfoO+xP0mIc4BdIoYei77n7S/Z9X0v4cCX
JQ02Y3VN0V5hONE3zQQHK0HvUv39UlgsKG3R8Em+TJziJP63C3P4J7Msw7RDZRFa
P7MtymOPvQ1V4hTj7pOtjO6vPWu6R3sxeGlIZmq4wsJOr8LtvY4L3v6sXM6card8
mlnejl7INopj3jwGOOa5awY7l7yhbHc9aNmH6w8vvYgQtvl1I1YayjIzB3RDBXni
HFI27rDm1OLT/rB7ccj/0G+fWJHVJgPiRuEXZiK7jCu5pmQLSPtsN+0wl2bOOmQM
783dpeBDYSnOYalWifK5XIzUyw9CZOxjVAj0D4S41rMM5YyPWhj3ULl5xuhTEEkw
A2R4hPSlGSGZ6i9fir64GxqdQ22Hj9DQ3Bma5BDfc3EJbKDIVYn3C0cSWFNu02YF
1Zb4dXxcsnpPKTwVTebmIACCzMrHCpJYm4K84Zk2bfC3NBCwn61l1LGhkT7fUGd3
yJfkkkqIZRHpOm7QvJMYyOczcrhVeX6szLpW/ugGlRc/tnqsuuujQzepzClE3OuC
HMv/eKy7yL4hVid07dDiaqQtT0+vrwFjH1bcRl1snbUv5tpJbqbNhde7RvcWCFxe
n2P7zx1Op6+OSidfQgHhIEv6ifk4soJWR8eKJ1piBpUDhgK/mr6m4WXzg9IrmluP
V5c85DayAJeLP7ydosfs+d/ha3bI3pQoawdSbjaQIVna+bkwKi12eUeGRMXARAhi
ptpnVw6w/zJh99FLRISNHxp7YzqnB+STp2NKTRQBnGW1GD9HNFCboafBQ0bXClXv
KHni7e7W+LHucSiNW7gS6S7UdCYo693gLgnhBIIYij7dc8CwyBIf2F0AsCTEvRse
To71EFXErs+sJ2UsbGl/tQy8tL3MUu73/1TTg7H32S8sT65AR6Bl3EYVkq5ck1D2
5kRoQTdGrFvJ50CKlEM4kaBYbnoLaAFbYL9EWdxoEC5Am1EhW/s3xNu9uPAxp4qr
5a7u1KDviMVSuccpB739dIV/LdaD3pM8OBAqvplYgZXbXs/4vqStSUyY6h6lJBNK
Z1Odl0DrTCLqghD/VLIk6KRIJZem1qwxG5CY/c/gpk+gdNFzt2dIl4bVb7R1lLDZ
hTIBABe0rUcga1VGt10E4+YEFBjCLqqE832bWwx7az1mqzSNH7ZD0VLHmD2W14v7
Qgs56R4DZjHEuiVJSJu1sbC+t09WoN98DrSFr3nWcZvtjqIBMXEjcYiNNCs1/1cW
UJ0BLKoVwh7dfG6cCUmKZx7sM3/WEaoOeMFHA5sPb6KJxUSulKRvFb69KhQtoKoI
ZGxB5OqNeDs97e6KbMuXwFMfSf3Dm82+OnQ8qYg2Mt4Ptsv3Vtz1VCz4qjKyUFvM
LhH7XfevDh/oS8+/bzP4btwQiEVY/vtg0IKo19bvF1jQkdlurJ/GrC+rVYLXFq/i
EzJXDIjcRlvlGdjqTdIn9JUSERTHcie3Bx+1JPqcsNAhNFRz+bJSg88WaG6zLN4d
rvi8nRUhprIn/T0pEgXjAXFFg6xIGJmzg+ob1ZLDPSPUUAjz0EYkbHauBm5FFW79
vD7gpcqKByh31Dg4eBRWSR2ON41Wu8azChwoADA9aoVp8CubMGSja8IA12ZCgX1I
rSjrJAl5kaArI/P3Dk4qmCUEcMiHmgPCZ092ts4wnY4xDTbW1p3NO5PwqsoYJA2u
mRv0bQs4aV8OdoVpNLJi9HhTfVAAHLbF2AEaxqVwxNZhCuYgrmTvbucv6FpiZo11
Q+6EcYBMxE+bMUPRGwoyURw9hv9b42xc7AkSPv5bWBScIsODPPrV4MfMV57ggPPf
EbJuhzoMCmWES5s/oxAyJjODPr4VgQ46rEIkKLlrTKJxPtweH6/WPnobwX8flge2
9eSsCNIlsqfvGfmRIDzdYGQJX3+mJCnURtGR5U+s8X9SXc67+FidCqt0aagELd2u
dSMTcHWBmpXPG3CQo7KqvXrdlJTSbipCM/E7nZsC3TyXmgU3SCTgPOJBK1I4HolA
D45LT7GtPvDQpqOgpSS9clhNDW4BjlXwGoPZiObuQGB3hMf/olPMquWDVz0GhLtw
9dosEJIBh25tvpUfyzpLqKKBhiMgD/s+HIF+T4MBu2LV6ocRUHHhBhmlBPhrrlti
nG+r2sQu5EuzjIpgko7mfeUzt5q5YfYK+JZbgHUSWeWgkGdnXkDKMV3e0eN4U5Kg
rWQ/8fIoEi4hydlGf0oDDaFtFJ1gf44+W9dT5049O2l9qfQKeM73MmCIAzSq95Qm
sAwdnR3T1B9E8Aezzt740XrOP4rvgNftBhi/0gh5kw4RicVcWwx2JwAAlJkEWImc
j0V8w7IK7lNU0wxXjEItcE0N8xiuRme6jzoo2hbsHyG7bgDrUTyx62PoJhelT6bv
K25RBoKv3B4ToE6EDv1vQn3ezY9+EaDemPckkFCz0BwkLlxGHxwErrHyC9ga16IP
rCrDshP14d4QDEjBYqkKSyETM6cal/kLl9XGEdp5c+UT2b8291xA0NBS2V18Yo6L
x+u22Lxz46EbIyIJXEtlLx0LOl8hyfPiNkN5VSDt44S/dori9mucyk5gJBozUgtW
9eg3wkVQ4YxJbYoGgEXJgeuNqypgoKqUhPnJ1hKiGMCS3rTWiKZereBqZM6u4561
wu63Xd0+Adc1+ofwQAmnSSNkrVjQ+GSrCsby80o9PgJN1a1w96Yp8p4rQBeCHn7r
50qHrIJu0f6EmJnNTvZLgwZweM+ZaGJCyAlEAdw723fqyxpf45OWeHUs0WcWk1Jn
6DVotEvLSyqQc6IODayoRsun1EiXHszyc2FU7udsaX8ciyg+JrFggLdUWh/NYxJy
qPCmAmOIyNekPEwbYXYs3xx5C0zpQEuIfa1O9fzCHOfZ09Nx7wn67yPcG7M0SZtV
yQTAG4+Iag2jxCBzyBoJP4EsgOQ0Yr1zBQTABIK4G82xK2St4QLUEXdrOuvQI07+
e4jqKwoheetNPeWD2UA8K/nX8TskLcv4TgE/OCTywQGRaJ8/qMhSLYuH5viPNVUb
6uQdF3QFa/aubEEazGT67guvwS9PIVXRD/UzEH9Z5n4sewhpFxiCpiMV+2+8WG1B
cWc77kDrrfvRccKML0N3B9/0oGUxRLHe2OWcoEmSJfFp8QrE4jCCvlEu4HuFwFEZ
/pOj3htzpacwaIxWk/3PlWC1S52bFkqQu5c9vvgLmWlBtA2DS+LVpfp87MkQMxXo
iQdhcdQZXF3ju8Q80nGsWeeVyjSqEsj6Sjg+EbnVATdZfM1+ihTpuncuKsW/xMn5
54G/kdhisRYuiJt8fkTqhTINDPuf405PqFM1muo6YShV3WysHdk8mGpNZPjEfIG1
e2aSvxisnHWRCTJEURxu+FQx/4IKQuLXX97CVtnm/oFIJXK8rMt2IvQSJXKzpvLm
ZKLGcMbugImQLgbSJtautPsUztBiaB+yf9MaiZO3cHERHrckInYGASLEWDbzgPp1
MlNiGWiYJlmkwXaI4twAAOq9XDN0i1WA/QQC0JiOIGDlMJLa0H58n0HbiFZTzJUI
iEPSgng4STEPEFyCizMUZUo2/f9nrFP8DEcM3vNUnGs2NgxOIa2JhbaoEUlUJ3L/
dtMTJMJpwG+iMG4Kmh7EOPabB3uBrCpN0KDutmGOcKU78Ap3l7wX4xYJ/YEdUA/x
rBxFM04SOZy23+dG9/k1Fi2G/IaNJ0ZMIRqcAJTvEpT9vG3kvniYhUmvI9l5GQ3y
anrrdScoJq2TDZt0hMYshH5vCTe7+IlheKfOYEneWZt3Vt6DfJWac8bWTM/qk2g9
JbUwpxJq3SoDFJuSOZFPOMpfTfQ0VRWkCrj9EVtaRELaMvrX83dyBc0bFmyHScqQ
ioExYYSfJjaHauH2cObQi3G0Lam0sitX6BkAc+YWXHi+aYI9JFRvDQTFC8nb10O3
UT/HFLq6wI0t4pXS32UN5ALU0NDowrPcXa2zliCONwRVP4zTnHBEhfC5OQGF4PN6
Jik5xxZaQcqLdJgJBaPReT4GEEc/kcPGsos6B0BV7zWitB1iZPhfQmnYR8gV4NHI
MfngVrdyB5VYB6exFIAwGthlEspiiSfRreGd4CtXDwtjedg3WiyzhAucnWjBgWJ5
Ianggto9FMOzgXHQNmy1DCmdQyfoE9pMSKYL+ajj5pavj24HbS/CC+m3zJ6CCQaY
85dkwTmETAP1n92pgenIr1Sv9eh4rL09eJzGeCeN27cN9adpyJjaokNy5gsdCUM8
hRfrC/QMBCRd5fQsPbLY5/iALxNGY8W13hLYMMgLFHG2BNHdpyWVv8lUJ8hh8Slw
YPFOSqeEe292wuvwqiZ4dvghEuzvsGsQNejlkqIffVnXYeO+WXucu7XmkX9tVfDu
xzq3bnacP6X1ktrfkqZdFobMt8LXi6k2snKQE2bPec9m1SURdwVgTXojUOBToRMs
rvA3il4w45rAuEoMskzkx8TupPhTuVoT7YxBYnAhcnggxLhCcD0XNaYjzNQ0zqQH
dp9E3lDMyb35ahO/zx5ZlE6AjpOL7S6kfDmfwv/ofPLvvlUnZ+J3Tx8mNH9s/nnF
x0n7cc0soa4ZwlkPKxjYoj/mTlgb0tqXx2iHMOTwKw2qUZ5jtCramFj32Ne1TmYe
wBQacsgpZY1gu+tPFTXtTaKIERB9kv6leKwreBz2HczP0qoWL5RzLmy2lxXgAOdZ
+VWb8YVFo8HhfohqWzlGUwc+HjXbw+F+xjKIVOX9b0V5PF+YOc8Nc63ccYqp1FyA
Yw0+imy2WXr+AMt2iO62tlVrwGOIRfAsvJdP99dDeC94+bYVxFS6c5sTgXXkc/My
OkismSrF29MBoURbaaY1/R1erKlluIzD+Z1216up+SQzFxeiLcEoyeR3rtqeFjxs
IQFBXVrtpmg3u3TUwVggYIX82oCYeYXXWhl1BqtzrRz60dXI4wuQml4tdPBg7ZmR
LU/SUfXVBob6f91J1RVM6w3LLQapdWoqVLaNT/dciKlN8lpeCmxrLS25IKFWXAuK
HhHT6j9DhFZ7mjaFDfnyinlC54mDey2mWv/vvj7KmHsYV9Cufa+YDpPt4xabEDPJ
qjvGzEqW53Zi+5XAzxOy4IMlTFxv7W4Tjk33WfJ1mV744qubm+/Q9YUfEHctx5Tc
czUCLUkgM/awncJK+3mKDMvUKdMTthK/DpG4K0GQKaV819Ud5MkLmVy908uRIADq
/uujvUpGa8yv+orIxEW5OOYQy0zKRKhKZPhpNAd8fWyNDvluX8zq5vRvzzrTY0gf
CbeO7Uv6oBt1sZ/Ypy+2CFCizuqpceyWIO7YdqrP6qVQkI7iQ37/IOweeFf23Xvw
mZAZ3xWWBpROOjwtoLWOdcJizUdgAOjIkuTQg/OnLz8c7UdUxMgpNPxL2xOPWyZj
RWWS9n2/UvGFt/Ogr6VjofZnAGQiGapxH1jsbhcqPtty6OuUUkDC5EqLddg1Qymx
Qr8iavjIH582jjnW+N4Fkc4A3Wlv56DDyeC/dClgXD05Vx0K6n4EvyBcTS6ZUm/m
zSYvuLNwQo3ewQuQA8GKUHOGUjIUAG8t0BOMRnEzDHrLtnuOy2gq3uE9FCcfevgx
79r3m+iB6oWrtb5TunE7anfnhQRgE8HLbjOl7vDeQ+NT3zVDZ7zKZQ5rVc6L++td
pzKseWHJUREgkReD+/D9Nk94emq303K9c39lXlU896Qj3d4qwBIvHHycHMfQ/mSj
yqNoiABPYQVidBTcc1wMmr7gaL7fvoRti03PIf5tKlfdOajJf9SqXok/U1gxMPXF
UBuhpG1Snu9yRPt0YeVjrjV+1LJMKkPYzJv6RHhqIBrEgApEMiwpBX+0oJl5pc05
Z2J76UuOKb7eb+ZeuB2ik6xy0ICnLOuIKGHSEJCj8VrafPCf5XvFBHvcufJFp6PD
kUhWWdGjBmG8q/6kOe8UMpxKtzuhMxqn3L1tZUaJP63iuxhnu8tpRp3n5BzRc4QB
0SD33ZvZjJkxT4F3lU4cd39dPTZljl0q+iG+WJybHbhX2nfzAc2ljqTO5oj1lOcD
ac1wyyw87wO7kdAdH60Qjs1VTKkg92QEhZy3+kqGkjjdZlU3MQMblz3Zc0FO5mD8
w65IRDNKc2V/JkvwCFxwk3oYgshVPula0cSR+X6tPouBb8iM/RAwt5n56lVskyCB
lAbI8JdTrw4P682PaokniZP0msT4TgqZ80xa07xar0PCyEtdGKp04YsHDjyoiZXu
IoZrl6Cp/u6QLOd7hwzto7sws2jSWNSfwlem8ru3vgKxTFXqsLIvXb5WZoz3ac4O
49FtFcNZO4CggoO7zR3wAQlcVkfIwQ05BFGmI7WA88eyWcDAE1fUxS35pWUWzn6x
8YfqdjPbLnUgkftEZ2jgWNvHuPMiGToxafuHAJ8CfAq79cGd0zd+AT9/kQ05ekF6
waqiXNkgPiEuhgrITE648nlD4llXY/x08QHNHNovkvK3f2NXeVH8hlfks+ydWbZd
G7KI8x3rodGyHHVOC4LqC2486FWZFYLzD9mW+CbhelGYzZl/anu7HUjoauE0aa+l
1w2LCs03Qb2N32cKZeDQvdApq3bFFAGuNp6OCZVSdARTpZahLs2/Tl4Qq9z8MMPo
qUM3Gp/GMVh0BSrZj1jOyowIOPFTroGPQBhdQYVP0m4r23OShXoEP0qKRlLJoxPf
L0C4DcKlFR/q95TnAQcA/nPFiMo/xbHto0sOrvkph6g23URcsTiMdi9ghQJIFlQ2
fzSIF5a6c0wBXvUuZf+1TKsfwcrokm/SLWcw5sqmxpUEh6hWoNxVoy5Yd3VoTCIc
20gK37JFqDrpWKEs1FWn50LSKBwPziSQGR8eWdtX9tM0T+GJuDImlZihGLmfVoZG
RRQQ28MQU80RacYtPc3DaYdo9jEgEEZOtTwguaiNQPUN3jifNGihQsPZLT0tBpfS
r193e1qem6+yN9lwJ409/IhogH1F539rfJ4Y97DbBSmvIYTR+s++i1jts905DA5I
nPUj8n8mqlypfqAMqBJ779VWkeiM9pZ8ZaAt6fY9tHcqmd5AovB8uhsFF84d6A/A
QJcPdGpSKx6Cy8I4eIE24Ic4vyWNGIg+hLI2jc9JcvE/DhUkwEn8O+LKqhgYp7O3
JApFWA7rTcDXdzI9tpzWCXtp4mmpO896h75xA8nYnNHe3grunDWqGUTFOthFvVlv
0W8+yTFc3VzHOZeFkWSVkTGUqFLJaccPNkzPU9fuw2Ikf/M9DDv7wKk0Shtruyze
nRmYRlqANpJ68t2PvHDPWROov6vhCEsLcQvrgtWDw9JRyGVdNfvXr59/jtCy8Gc4
3mlMaGOe7OQriyXUW5kyipF+cAWB5OFhDROwnlocFVozNMRY/XrEv2lQvXI3A+F2
57PwzrbtfY5mmcjP+jFeATszOpO2eU4XumOqF8g9PCLYJzq9mEhZMdnQuQXfsnFF
E8VXZpbHb8skQksL0NcjJOuAYkiFo9DduMD8/0s79u9j23uxs5rdVwkx8/+btwQy
my13cZhojFkdmkKKR8vrGK6QxrP/USNasLL8uSZ/DXykPypnra1Q89UdU0nDchGB
yWySpffBuwJjRGwqzqn+Gg0/nLng9kPB9gPHFxAj/nkAnlPHxwVkSgnlwqQXZQpk
izbPVTYgaYtQgY3pkdL8ATUO1YEn2jVEbgXtvZzysveXHw3TketscBnRLYpe/Riv
CVkHSBhTQ19Z4qxkh0cpzwQ7Xo1cy0YCAJtbgm7qmUEfae7+I42AXi991VIHv0zZ
T+YvqqSLMqHCBVfT7VEss8iaQZdO1PuXWTpmRaIDrYwMdyKGkhzO2aqQDPN/3hTg
l83n2eER0j9GskWlrHHSV9Kk+zgkT/fNaZFdtTqizfz7SJiYegpOYTf9jhqVckrC
rqeY9BkMd1IIaHfNg/EnOU6Rlnac5HfsPTJor7heDWhfoN5R7hePSes14lVV4yHK
tF4pXUXul6XLp8PFdWpe7cL1LadfrqWxGySzQTZaIZREmJNyZKyx4SFdD9pxlV9B
XWlqOrT0OOWhxtsjDbeMIp5jfJzpBnw2uIv6E7L4UNbatVRwyLBWzjhoDZ8psNvh
pTvtBJ2QISa88+1thabotFoA4wVGloR08U5aDOalXNPtakETdc47s1x/91P1vgYC
PwnqU3U8lTLahP3AN/0o/wVvsvq+0OpdNwtR+2zrXecnPVYPij1pPTE4Vef+U+ji
YItN3+H0/pJtOgeONx4poT55hmCf1KSd4zLiJXzR7uWr4VtNn17gUifkYkC0ptam
gbDTYI5jEVPDky5OSm+ZaW/hHK3upS5V+QkzBYDsYtiE4rlpX55CcrtEeFedWBtd
eoXKZSoV0DGExL9CIBqYpeY12D3wKR8k8Vd2R0WRKBd7U1cvnisS6DfMGKMOlHlT
jxxwawzqjBR+Mypzw1AtVVYBKy+2eon0+oEsX52Q6Qq2BgLVXpj8JkadEq7e/0EF
mn8QynQwKF+lzEDvXg3AmAb/R/cwza42Ytxa0X1rj5KoWvOFa6ZtnC1pvqp4wtE3
g2tZJO5XMAB+IWSwgm0Gx6r89HSI2NiJY2bxk+pcy8rWI+KCjwaDrYGPN9tpc2W0
YMHpXlAlnETdeGEFqpD0KtQJXkG+N8AMosXJzVlWoskjCVTv81OpFjHulRrNo4u1
uyaBIGrbgnAI1DIc6pZ4Hho9sPahRePvpsMSByp/nnWxoG92hCIHgFYfZJQ4s3++
+/rK9GOpe+Pm/d73tUIRsA/Q1uqKc3vUu3z/0OXzGUvvQoG6niBlAeV9BovkiH0f
Co8BBrDQZGGFqievO0bLmW2aGYOslrQAXRYZv4mwqm4SXj4+2KXGuSVhfyc91UUQ
RSY9m+VwqhQ0oebjM/CRNRRJpmkyosWwB2ezmeRo54hErCeNBh6bGFh4WZMRB/BA
HK1QpmkSSQRUF3S5F9hb9hjqVeB8gRNgrbTfwKPZNlcDOCiW1nKmOaDBmYC8VehX
LiiYxDLf5BIVIAH415oAO2ZXo3GJAtpU7AB2StQdOKsMkK9dCsJBR51JpP29j4OM
+PYeFo9hcMb5caA6QpFRlSOje0gJlp4e4LTi6wbvKisqLPs4GLpqN7AnHkgLnIUN
2gKKfANtCdfFA+6L8dfpDpYLWYZQXx8Kk8L/U3rFpbyraXPt37h3SiZF0SUR5kRa
wh2/noJbx5iUoAZflFlN9sKF1rXIgIQuF33h6CxacRdGNO+vv/HfMZ1b6tTqY1eX
ty7zoX5uw27hs14r/Iv6jNqqQ2mjilpRNk0PoLnj1RJ87QT4AjgnS9E8iq8pKYO/
tYmjLmvh0Ek3V4w0y6oxIrd28ogRJzkrPpSRt6GXjHStdi06/Xutxxw9+Itbh7Bn
OtEtvRJzrZ2hL1mxgeRMOsZlh/CmMnDU1g1MyGFY+SvdC8oy+j+Qd2Fj25548B/l
et8dnMMj3lhf73FXV59qFgzvr72M+Kr2UlQTsIz0tAr8p4D7Hjm+8mIkqw9c2dFH
4TT+TAHFr5ni8wcnKKIHJg5wj8QtRSn6u2w+MtyWH9hhQB2aK/93++S8VmoYpom4
FM0EN66HhUFDtWFJbMudLD9gzAmKkZTqzQUtKi3W1l2FRrWIEHbhF5rrCgh462Ey
Jg00r/ZL2zPpJ68DvLkSw1I10H2o7TgjXFCMu4J53TL9cYFqaoxlE98oOYQgvdYC
YpUQsPVxfzlyaZBQJEYrbjk4WHBCASvv50U3UQdMRkX94L0S9wYeERLZxBhqvG7m
0J5QcCnpK0BujQt+crz03/gf1Ogp6jsuy1xkFZmfSOlBJhPNYTC+OtxIyZZ+cGzy
wQxy1MTO3Ha0DDF4NDPqRHQYBqOGEDlf2otdsv65B+fruwm7r84hwqU6m7008SXf
EKqDuOKibNYp6FmmWR9OXBdQpcgf0+I5KbEuQh/s/VzxvzPYIKjoQAb4KUrzZxyf
Em2m4FmVIgbJDSJg/OiQKfI5la/WspxNF1xgyCgY3+ael7e0e1EeACBy7FrBBPOI
0KGW/dUVUnvXHC3TRRcSgHAlPCna6+6dr1+GABjIiPvcYEGrXqRlmMHrzg9L8h0J
s7LvDWOMPVFgAGpUitDrR1uRQpEwIA61t8Y07rViWVA/g3svhG7x47nFwCsHjfxi
CoZjGPNL9HEM5OIMQKhJ2v9OwgdlABxyPjI3Qt8lUKDyEAO4s9+Lp3IuE7iVnDiy
f1fYULlO3EV8ipSs+0b+zsMgId5W6YqcOc0QG7Bc1a7HcwyUXRYgx/b7/KCOMdno
XuQFuKx4f60bf+/R/HIVzk8VmEA8uh6oU/fExbTFUOWPHb8Zg/2jkq2IYd6AfESF
f110UkNU17sn8HbYS+RDW7XvWJhWcgQ7FVXLEiQNDcuPbN96QSdF1w35zO1IZFFD
pnmbcome4wTQP1WdTINgnN5ndxZ1ql+MXNFbjMm+mUZRsXXaCGNBNfILmaPW619n
w5cT/SiHSNXnYJrAdMmk2+/mNnX9Do57z777dwN3/7kfRiSsQkCOng57mQiI2NId
w5YCMvEVprj8d3GzualiezE7RlPO9HE/+nXm7UB5c+RmziF1MuJeryxpGOKozgMf
AAJhUpNnPQitOCzAD/aKwE78l5qwGbg1RCvR/zxIEWCQT8AjtRChljEIw3BxXBrN
J79pVSUiHCeZfvRPoCYe34EJPrv7DTKsZpD/lxwktBYTSm3Y7XrPF0JvJ/t8zhIr
v6k+IyNmrALIyGz7Uv/1u/JXquoYdy+qyDtBy+BxMkeL7UJZSMYZN6SrQBafpWPz
+D6fyT2JojgqcgvrXa7RfjdldVE+bHid7JQdi0ZiZ4yFj0f5Lx+AQzJIYoqwdAzq
FZpDDlmc56BML0LOeTYYpogEYMhY88SvnDVIOz+4ghO+jbIQqYdayK+Ipjv/wT50
+sJ/VuwdZRZ4Jd6MA5ZhLls9wtghKpMQQO/5FPjdW15YsrU1Y8+l3tv77zs2kVTd
7e/Dt4VvRuEh8hR0KZ4NWCloLM3rn+cvMF27ND9brC55Mp0FBUXD9S4d9+0HKEfY
V7T0ihCbbNkQZovgh4MbjrTya+TGMw0y5mg0zYBOMjqOKUjgLI4b5M3GYX/LQNPk
G58OshRZH6KMTCMPrYogEADIUFrAfvPLtQRVmw+Aq98ODdAFwu8C09Y55wfRvfXS
W+Sfmpi2x8RrkSD+68s1Qs9CSvjwboTtzh8ETQtuoEjD7IkqUarrUK/UoM3Cf5UX
y/3japlzjcz2TRPyCT0y5G74grt9x8siPsnvP9OHawaXRPFzs1uwMPqCSO2eoRyN
MmgcGvoDl7igujblKns7mR4aWBGhjleV3N5L4xWxEe9UacJnBKCN8BuLVjvmELZh
iqbnyhbBomlT+BItQd/tvCZ81c6l7290O3RqvER9VaZdMJKZzXuAnqBPHuDhguyf
jFCekrvMjhNUWrtj/i/Kp3NC8dUw/RXOqEPCErKZhP+KjheyK/DribEj0aXaXAgQ
Wr7VLb339NruIU+WR3tRTqKvpWNlY/fRPv0NYc49YNKEtJ/W7oONrHhOaW08Vo80
4TfhmzHSdgC6gYoTN79dzOHo9oQCwH05owQXpwURINyDdesPmMfyCo8nsEbYp/3T
Fcp0a8WGmppfPYknDo7pzndhBFbev2Dtc+dl+bZ5sjP3oxmFWHoWSnWeGLn0DiaN
Jmn4tRpbkrCml5zf5eZtXedeXM7c8tcDpUZphpnixSMGEvSIGPhnv+5N1HppliEv
SH0GV/QOPVj2rF1Fn2ow9G4Z9hOnTLyQUXg5a/tL4oFbi241LAqdoUsrEsplsJFI
7Ye2IsINv0+yxuTdamQkT4dexCCsRcR5K3MUY9vZosPyInn5ahiJNgqH4dEqp/NJ
1dmybw9egtCRizWIBFDaKSv6pe19t0HEXbdnfLtu/qOMJzHiQvgxFIQGw7Xj/FNm
lxABir4f0WW7IZP39s1OVeHF7soFhQBca7MOBGz9lD8z7TUwUhefxekx7zcn2p1Q
w6qkWUx2iYkvwaAMHaKlZfCHKYM7JXmpO6efWzo70C3b6/z3IzLquKURAjgEyZte
S+ns585HWsHyzWcr5KmBUe8hGlpzV9vKcf6YqjfF0wmbQxFeVbiSAZ8VbCOZgW6g
Q/Fa0w6jg/ktQLgvDeyOWfK9jLsVWVo99hbxoOv4bVFEqf4/ZDltqNhHHWWG6Mfe
24yIadrHNSddpvejl4mVovF9hQjhUL7BTFWXnNVjUmr5XBL+YlawAXEbJqzeRL2j
NVuUrYsY88htAqyMlmaaNLm/Jndgqmm3umK7oXgsPrWhpwv0CwbqBSo2hg50pGvX
C8CrHvYuAweihy0TmVzMv9TRwaijrJl9IAqS2Uy0KzMnP8zmcs0wYAIFKNgvc+4A
ARO0D/DIFx3rEedny8xmGWMi6tJ0nsISpScmwQ/xA4qCMvso2ZNc46knypZsuEfe
mxO2uxtIzFJVE6lXJGMIggZPUWqwJRD25+U26nW7IbJrIo6Th+ZehO3ks3Mv2FqU
eu9+TY2cJNsjfHd4T8f1rCS2OYrrLe47/hsQg8ljp1h7nbYUKI4JmhVAR4iVTxXI
Ks56sAhbOXg77+6fxDwzxGezY8LMHvPRvekduf4/beuRRk2IwC0zUaMWsp45RJjK
h587mWEK3rlQk6vRY9X1i5UFVJhYFwF4bDEL4j6uuARW5gBqZ6yjCZi5ULk6+z5C
dszSK0MBRSwFJnLQGYoVaOqYWe4d6D3UwMM/usxqkIckqmjvIQz0CgF98N+P0kxQ
KATtI6Pq4tIzKLtjDvhGOIRMlGN9WfHYuWl5zzGkuwlYpwHRFKQzDQ0Bu13hhGKA
Z7sMY6yT5jxC3Bk9K72KuXlajxZ4yxqnKVkRvlyi1BD0grnc/rWAmzoBOEcq8frW
O8WzLHkJxdE+IKgfotP4nmy4XRcqGEtPRc9ylMkikQz6hp8xdeekJzJssliEfafc
jgiMiXadIFCuXocbZxetbRuqbXMEpiaXC14kQ9SET7+KC1WnqHwXUJXHBBmui76c
gKvHvuliYfHR3tHLtDMwrqXpw6K+vx5uFM+OGUVOjz4F3dN6ZuuOBfAbn2MX5PM6
JBhqsH3eCKLAxQ84QHyEik00GwR76al5wqAikOmv8mzcz7fCb/eAwlRY1SIZwxOD
rGHFYvcGLRiyDyRwErgDcLc0i7LkVvHxuzToCb3cU3aQ50D+Fk72duQxHmO7Szm6
ARpVK+z95ewrTtV/x0+BGmoOr27fisFmvOwt8uMsCLGoHCgr4Djb9YOpPNh6eKtW
rTCDs48lAS3rPlEnCXeehfdj0/HSF2FofXBAoC8HvCVff0wQ8U7W7NlthloVuS0M
B21vOInoKKlXkDYFKEMpQ6+piEhmqLOTRfPWEklV+7zAjUYTNTyXDfYeIqDj1Rpb
0n6ZKLSHvQil7ax1N8N1Ems7/77TVt47P9ElbJ2RJjSCFY7fRuCuwJJBmYU577S5
3pMSuCLPh9j4H9gT20laxf+1LOZPOzbWMK5dBj8Xw85uCTc0IGFwJQyue5PmRiUB
e9vBellG5Hfi21uwEX5jggascrw2gp75MSaF4T/Dwprjb0gmkEoP/j+6yJ+VAGmZ
DeOzVKNnMJv89FPxObDLkF6d+CeSi9Lv4TBDW8SH0Kgb35xyzrF6RxYfrScTISsz
reN3boHgtImEUl2mRMA2zjWpUH45iCu34a70ndxOTBC57xOg9mkxcSb9P0XlPzEW
dYOVgt/MQIDJawBIPNn+mtMqGETnmcAKsJvgzW2Km/AlHeysi+Un3MbxObieuGvZ
W02/Dw8jn2lMb+KGrAvF6OOX/zcfWWy7LpfAU9kSwOKjdCqD7/w+VPJ69PU0gXqZ
+CucqQUgi283gmL9AzXQW+98PwE26hION1VWbXYfmIKpzk5lO4ojYaCbDTX76Lay
zasiJKvptlwPVewZe9jINREK2UUjg0125GXaLACsZr5+0k3g60SdiwTWMRVHuggB
Xz8JLlz1s8pv1x19YC1Ndx5I+YFkVqCD99ssC00G1CNX2zUz98oiFTVVqjwQNIAj
GFBsmcAqinwjgAoQCt8+Z7b463PXS91jzBPgwrtK9R8Wowi8RvQxXNEDe9fn/b7D
jGSy2IXF8T+VDYiMkfjgUm1uzdScX/jlwKUhkK1Xl0aRUj4pxPStgl9ujJk2ovLH
sM1xBh3b2i+rwgvMKrSiIVwxTMxcO2RpbXzEIR8mU7Mt0jLvmu8xvypdT7Mn3tsC
Yv7+hl8lZl0I4aURkK4SYGLOBgU324dIodZrsgfnCCNtEbgXb46PLg4WgZdVRi1b
RRitBM9fB9Jl1d1DAKX/6L1Wq4GTT6q9eBflW72sDvq+zPFu8zICBSSLu0Zyh2T2
yvFqB/Ma0Q5vfuQxxx05Pfo73t2yWtpbU+SJM4cx8sePHd3sidEi+6byQLscvUhL
EEAQ1KF0+5Y+dq2xVnD9U7qLdsB1BD5XH+NQwTXH2LInEvGJa5rulWUyWRxjQxh2
fcIdOqavVT1et21ZQtTGL8B8wlM0WgVSiR+MWaxVpZKd8keN4j+BHw1N12OYuXe+
yZJfr9GTUhjRlSZ5yKN4Crqq4T6xokFKftnoHkldXPZhFccX7+o1hW4qYDasEHhD
2M4xShp80bA5aeMqjB2jvCOO0jFK1AC0HL73U+2VgwkZkez6pGbyUZmREIW9MOBE
Rjeg/FBEIJxbpEThFXVNMp9vmRw3UHuY45RVD9yCBh62CwTPqpjrQy3Rsvmjxok1
G76tXlhMA+XjwyV5BSFzkGI/1JlmOFrZUpE3OJ0/ZqjlMnQa3hDccvJbYL1qD4DJ
CPn3/Z1qMC8lV/t51FVSqQZQwVZoLrtkrdyevxobdgAiU7cMlbzFOyK7C7GtbjfL
1GcslPyPSW47DXRysQTnGG2NU7DY4NzbLyYWSb4gxSu1xPTJTmdep+SP37TKsUY5
XENRgon7drx4UhQkVklAGEoPWVSeCpQ8WbAn0cP3yLgTgHbVCf6r9S5jOENTemeF
IGo081VZyU5SqDUHL6eGRh4TQZVcYdDBBA1GvQJWwRAMWxnZAOOo5qWDHOCYL16Q
war0N5FbcmF/acfC8KDi7xJkgPjEy0+eQfjlFCmVRPEcEdZC2Jkgt+xMX8g21iPq
FYrszInqyNJsUZ5m8SSJhD+WgnFrHzHi5MPlY7WnkKpxUrc4zFrp0sskieYOzBCO
oRrdjuEr/8DlphPMEb2ie9e8+bB96dt9KeIyGBq+SicKWYUHG43HiQTslIpMLix6
Z8jTV7HLxyEDaVRFZ45hKETI8IRuwLMhD5HmYW6oVuHN0LkQY0IuRUA5qRRex0Fn
vdtNnvVKyd4dUjlw+7KMHbw3miiihylPqm06l3psCGaxtgj5b/KQExMgX44KT37+
iAqnrfmyhh37H1ghV2uuQwtMK/MRM3YN/mEZCo9gIyEIZdObw1I/KEfhGpW6Ydxj
QPXO5TsCKghO61rUfQdTgt8uJVKpcPJQDkZo/y2Ubklhwl4y+gB/BO5ppufCtlUl
e8QJT/X0ZOAEro8DuVm8R67l9emkHsWmvJUvMVOgfsFKZVRKLFd8ue8lxqcgVKkY
C58vW+tivEJ72KVg/Li/hSEeOdqI8iZ7gBLRIh/SZRFeSWiWicdLHYxZtjELMbd1
Ik3IzewUGZqd2M2TNe2DzKgP/fsoGqXDnY4xob7V70UNo3pyA8eUzEnuMOPqba5U
mibjAWwZpBI+0RYve1CQehQtK/k8kgz7aNhjBuH8kK/QUYfdnROXU09/qgc5lIfy
gdYkWuwkx7p4i29lEiakQdDYSqFmnMVOP09wMBXXdibvdYX60TDjz2OcyTxh2FYa
cvGRya8nmjXW848aCSzta9h3kBNKof7DTRJ8mGQVsglYQFrBTCVAMkzjLwXhI4tT
shYSLXcKwlsbKI4d/vY8DIVFv8lyifiKOb3hq5ytlRZKVZn5erX9IkH4divR21pv
9dRYbaK5biS/mmj+LxJzLrDq5b5/uPdZ2Odbp7EF1DYuOPssLO5lu2fEo6GR1Lsz
oY13LYO2FiRnFIic+wgKSOnuHNH3omTScECQuziflGkKSsx9feUq0ar5CjIFVM1e
oOfDkRdJtqo7SpUrSNAJro3nj6QgRprOVxGnr3U8tpcYK9FJXyBVFazkpUCayeCJ
gv6L8RfisbdMIeLJMtOp2RBnbDa7lFKaQdLKWRPhu4SA8iz+g+yXgqH1ovkWINLZ
yHeGxw4dPwwNnWvKWy2KHSiv1SDMmy3UvPVSBB1Fi5byDELhY9x9+zEz68kn3m7L
xdFnKV70hRbcv4elqAQ/k9BEaf67xPb01jgmBbapf0mWZ6oeuzXcfArpY9H06Wld
Un2hvTm/S+++EwFfH3wuVkPFDWNFDDoFvplgxC+gvpi1GPo+SWwL9c21doHLZofi
x/AdA5URff4qvA7KcQuH5Aodi0yoTW/LZ69F0u41XHqhTZbdpjh8DZxxlBP4qq9D
EDt7mDrVPFJv4Z9g+VzBIOlbEUkijuibDDCmK/Jqa5QEy0Kqu/9TwGrtGidsTV4j
esPuS8kvjhCw7bFLAZVJhNFBSr/0DVmZVJyOy6IMZBZNZ1SnVFt22hwFLnHj5t66
Ytt3lMosWt9j84zdeAZuHEBp0VMFhxqQcB5olS/X6rbKDlOqSTqKo7euJb2URXxi
49UWh62dBagiQvxWCaWo+Z0LkDumM4ceOJi1ICJ6xTRp1QJzCj3Pwof4OcpiH1Uq
0jgb92h6W9m/uKn5V7g23ioC09E7VP0uvv5p1z2fALyDRtvJ3j+1XRbbx0Yvs2xp
ZAAPsU9ictDOdnt/4//uDbaGhZcGO43EOTsU9vWU0lBrPU4A6YspBMKaWNe+2Wib
Dki9WkgaAJSrTwWwPPUOVK0ftFvFdde9VP9DhELNG5dUgE8qIA7ICcGOQ+iTp9TQ
1fZiCACjijhsEY2k//j5acRj1XSxg+a5CiiCOMxKe45rz/SUIJC4CHYl2DGBDD1f
fqy2ho6QFDNN7df3xFWCI7+TH613Hf7LWrsDsBmIGXY8I0+x/Pqmw/F+3BSfBiHB
8yKl4sg+s0WtggKDQMkUn7Hh7vOQBIseZPTOilxaWE19HYdgn5G1CAw+cQQhi/2H
2UZ+oqC+ZDx//VzulWX5RTtfRlKua1U7tP/mbLuHxQsREfXR3momNwRFdvplKSRr
if0DR5cmKpH7SvWl3+dXeu8AYG+2dGB3YY4SoBQ67hnzxXvUdP/yY66quOwrPT9e
I+cHKVkFrRM1bvXNKEGGfzgAqrOmKBmAqQgo4nxh/erL19qeRY9813GbBYqK77Jv
C3fgwx0cZOrMne5NvrjohQ0m0EdRuIz1O/s0gNNkNQB8htIv3w1zHjLa2CXT3QTx
VPB3eJQapqxCbkgwMGCLswGLFCCPCk1ZliAPGuQh/Xtu5zBXvvwcVbnNIpKcEASD
qFmNHkwuRg2R5mtT+HAhPD4t9xArdhCuqP9YVvT9BsFc1rnhUE007FzGuEl9OoMn
ssjDSjViiuRw7huRAytlJKS1r2L504fCob/H0ds8SH4H/J1Btbnsg7Qbl6nP3QMP
W+GKK+AVJabAHSJfLPiratbo55TqQSVoccWeyg3cFgMpVuM1Dxq8SQPPJ16zd6QK
uQEAqAjNGKicUlfTPPKhSeLQLKa++492gtRSQoRDoAxnHrGBv3n5+uJkrF3G56R0
y+PN2G2/o7na6ZuFANbaLObYQ1KT1xtsMNBAZNwHk+qWv55+nLw6aIpuoObdhyhl
xkaB7asjaAEAjdyPiY7ky+f9v82aJlWJ5eizfVUCmxcCtHh+fH7lxja4RBh9JxGw
23Ji6wYEiQfOGBTCiKcEe6jp2jxLyxYX9i1+Yi1W5QFI6TEmmrkMscL0VFrAAYIU
SFXAqekgi4eRMsPkne+kC4r5s7TxvDoyFe3mnLBFf1yesCYzO3v8W5GgRB3dQK9E
QtscbsEjKsbY5qm8BH9n034U202XB6hp2KaUkTjvKRGobQ47VFHoFaxvdjC5SNqe
JM5YY06MLVdFvH1+uFf83OKT/KuWT51CoU6eHM4Bi4dE821tJONjEx/mAK3JP4l8
SQNJNTftRklZgkqyYSbdusu6YFXExmK4XjXQerhVE9Y39roZU981IXeTlfBprkc0
iAPZx5/DhPBfehoLLVvx5OmmoJmJ8d0FT6XXLRbGPJ4OMAC20tHvP+h4TMYP8IyS
uHPn6qqtVuevnew6Ia5H+r+EvGASDzlUjM+WjTqNSuctuszytHkB1iAb7J0+8mu3
fJFXAlnKh5ltZMXCV+yV9gMIQMpVHEdXYj3o60atOJ29tvQ9oFM1nNg+1vhF/DPn
lmo/8YigxwHUNq+/gUxhhdK3gKyJLJHHd3ZRJHnxJ6XMh6Yh2KH+ih9jDeKFx6Oc
kKmcKhZTQ2VZII0qj2VSDItAjITqfz0d3yOVEoX18RCudzORTADNdVsgfkuCcS9z
iC9o4vet+xVBrqrssHkg0+niNyXlQgjTLYvmaafGYY6XVRqfXYVjWFlH9JC63z7I
2OH4j++bmtodK/k03zFo8fZIanFjkDxDbaPhkSlvUiGdEGIe9JEtw5xKgjHGZ/fb
5zTQvwm+qKJzjh4QNxpDiQ6dSzkaOZjCNWVMev8XIM+YAHp38mIBsI5EPV8Jmzol
li6lbsH9WVzpb/XldI8hrFVsNc0AIw0dTumnH3HIVi9A0uZ4uhzHt9/gKrSsWEaM
EvsfcxqNmUfWTXL8/VIm2qf6jlLUMdLTk4rASTCw7PQ9lt0x/IEmpshmLOycrQ2f
/Un+Bcn1I07Pn+7bhupMNU7cQYa3MueOg68+kxGtZLjl3eX7ioJxS4CHuXPgkfBq
WvmHOexGHQE4WmyhlgvvzAOhBI5/CNMjZ0FGsmbh2dV9LwVHt5wIcqKhW7sYdpCp
lTwPQR+ClX6Vnhz/k2xiVQyOexKpUuWjSixeQu0MYzpzYcFmpjzv0b1lhnrNtpGZ
qt1yfc2XIU4cmtfyAcP/UPlY0d9UUheW405EVaK49qYvp62m33tWwtYouiVc26Ko
X2TUeeB07FED6DVMVNEMRKC2eAXaQf2btjBz1eZ6ZiTagSK9dNrofdk9q8k0zv0L
xK8wpZahmioHu9lBcKAAvRmWXO1bCD2H3HExflxhetHdGsW5kzTrQJ9eab5q9oPL
Drb+uejXWJvwtoqc5u1/2LyJfCA8R67HrbbELapEHdxM1QARwfXH9ITelMorxizL
sXQEhtNqWYCZvseLHkFDJXXqVBsQxLBW+PtNMBBVlM7a7iXXKpkrK4SGak2EFvG+
K16h1MAzWv4Q6HTsotEIOv8uvlA/f4oqepfWJhdzliA3XdIx/UHoqeziVMFeyDP3
u58JV/tl/d8iB7tGumC8erQM0rFGNQBpZVwQf1UHoQnh3vnbdtPREikS0DST5LhT
3nA3hppzfSj3ISFo8SulVfK13kY2FeJeZLMV+qZqsWc9FZT++unV8CurCVWXcns/
trOXilL8WN24aa75Zyf4/TNsPgij6g9DYukg6Fc7zQ3s8VUVx4NWcJxhBj+LlHUq
qiEn1TJW18JJwZwPkKEv7H/tBc3JZI361ChxB69VOkmCYpcSqNk+fig0issww/E2
bsU3MponQdTobHZCRjPtqqzNBcHaVbybrgOzeupIatU/aAfbat9mc8ftTsP+7BqD
snR8uteMLNKFrvocIuxZ+qFgE7thWqynxAD9dvbzirJXe5LdZgfgjnsmyrkabys7
BZdOcBCDZ7EMOnBcvqx/kBW4dVeQ0paJr30a12OnRxai+Em9f8g5f6fswF1Hbc0/
0yzRv5wntVlQUU93eyEuPl/W0P6KWQgthw8LibcTAdDUH+NgaGZ1JUvtxyUC32T1
UX3CQtLCOsr+UJ/sBmIYxIWN1fgtmEOqs31v2mKr5GCq+070ppZ8r1iv0F6LS38l
AGX1VnuOH6C7/yY7mgAlvNF7LAPeX7EOBNpj1TFTPz4jigYyuocsy1zJ0F6DCOKL
ezL6nDjaEysZ+kFB3Jp3FD4QXJ5q9vCm/6m7dvK6iVthpnYVr2NWXzlqlXfLXPVD
MVI0J+TlSTvCRuuf7NrPgTzvd+jrFuTm0pKpaXk+tYncofNqiczBRMsvpLnoon42
WBTQUPCeKPSR0zFLgeHlTErbiw4mmSl/c33wONlk3P8hnoe0d1gbO84UNkF9NtpI
w9FVjm7smZXMWjhkCxh8XqCWWuywrzfWExcsZTBS3zYPGuT78A6behssb9CLyD6I
bX4DwNzX8lo0AiXdTlttaOjVhi6GzJL4yqSbi4R4ogaIKSzXN8l1CcIZdGoZDxln
wVRVZqf+j4/yuMVCgRMBKYyPuOSAlqSbpIXOm5i+iSX0g89JpfF9k3nw14jyl3qz
c5nFpvLZwJqbVT5MzySqbM2OMWuIVgUnPdv2OMUN/rTI1JhOXbiFgtWKnyzzl8Lq
a1R6BP8EY4SVK559jCn3MZbrUugc2g4N8AlA92QEoMwTXe/5r5n/WjLgrA2MS/mq
YYaDOJBlfKitPNs07Grvod/H0rhCaCSF4upP3xxju7MkrXLeRf0bqIQz1lAWQODC
bqmdEF/2yoeYw87fWfgPGpKT7bHZdk6TF/rnwbxjuG+6oHZvXnCWNYOGpgODs2ns
SNnZFpFlXwCJH0XRPgd+2VlpSccOqSESrHUJNm2z2gMFjkfvlH0yqLKPkNjO1aex
d7omIxLMeVFVEnxWVTPvGYw3JQoovTNbDVm+YhmbFHgq1vcxuMOQylwbISKmvoSV
6D4HZ5dmdTL2+qBMAmb8C4j8VinWLZWVYpAgsEyJjzcnUtYjG7H8l1WYpGNo5JLP
PKJ13gInveDOmQAtR2pvF41rkDhbVSAS+pAhzjr9FzB2Ju0zmz7qCyWRjYHF8Og/
nzLgajjpPo0MwXfeGUn7qolyyZBWl2i4svQEHI6thY7eEytXkzX4xoIg3uPYZFpl
zcRltRmkT5Heu+Uy04eX9HEz2QQ0bSIDzdG9Vw5A4XqKn30cIZBupDENBpBWHUwM
CrXRjN6SrcA3cQaFv3rq7nsCkpKSJZPGcNQedv0md9GE2t3Gheutd0winT/rrCvI
fZzgS7E/pdiltyaNna5+wvh3l/udhMOh2zksuqQEZ/GODLAdEsLoyrJnlFuzVBxp
OPjpWC08P7VzsiT94pwDgLe9j1HZ2gIEIzHDFQxM/t3S0sJ5G+3ZAXZOOvilxm72
XimqSC/5EvlDy/g4Sys+xrX5/muWQj0tjA4b2NOihyl5XzEV31g2UCwaCU/6zRPT
lyX+0FC6zosIw0hqBE+KEExfKidDAnm9drtk9mKueaOEXI7cgjjcQtlLP3tkri0t
Bbik+DqFYHZbxTcflg6/4RHkN+sXA1mE3PqLd9nge6HVtYODb85Jwhj90A1Kbm5X
1bWJ29bPUoDZdGUOLNDeJjaplX10Oy0WXyTTArZ02WjF9NoSWYzyA3jpD2dnHV7G
XGgdaws3GxdmXS553i8Qqosjhx7KlnsIoBM0WGc2YbggydRn8gdpfCwbX9i5jSc7
/DerohYCFpTN1wcPiekAFUPfPqnwhIVeWrnwsCpsW0Kl/He3man5IG64BLwz75E8
uuhO7usDPq9QuJY3UGmrYWANq/sSrbdm0kFXn2vmo9EY6ZoxwCZvvXYwUeteYElL
HXHZzFbK/yQrHOg3E4mj3bV2mjGDCJeHPm5kFRzny9IIOSk2bU7WkCQqsOYXKmKl
eY9p/gWowB5tPxVN4YV349I8hAwj16mRkXsJ27M04zf4YAn1TFC/iyRZF7jZsbsX
rOKvTZknzxsrt2s+VDKxFWbSEZ0VrX6S8piWh3c/pesAQLUjfw4QbmSuSxrXIe5T
MUui4Us0hHStaFkXP7Udu6Y+KPoRdJH79OQZPcAaN15oW4UMxJjjdT3ZCAxSbuoP
/HTv2nA6FpOI3l88QzsI7mlNvAcBMAWghWdB/cY7l7CId/Nt8ksP9ZAczKigm1dr
s3nmDykiZAUNOcl2/3NlFhH9mh24c8koe209CrzRH4YhJqOYhGcmY4Yi1nuPVlRM
Hq/X0LPKuHysYnF/u8urevQctLWnJhxGQGRWQZCMBKgETTAQ7Jcg1jLCQEg1nYzc
WGEbEz1jxmo3hfQArvryoPJuD3z8mGQ4kFm8riouwOW8AWa5eIKVzVAJ0LmJNKFd
ir2WMpwrYX4I4HF4GhNCyAmCRcoUT07FI0M9g3DhhNS+2TaPp/cLtIiTs+HR7869
yK+FYEwi+18wtRQtGoU93qUGUYaNw9gwi1191x9Lp+/ffNSrBL7mDsDVTSb9xoGj
MpdBgghQ9awVNRt3aqjugRT8ucMsoElaSR0b7tn4yzhqFRbRUpB14RrBv7hgZPKn
b1ZYFBFneT+yTZkjZr7suYzhOHICrI80UxqVQrX9gDQGdUYiGutpmCJw+AjFZeMV
V7aB6dajpYnoacV3sbnNoHQlfImKPsucZlzwXyIiV8xidFqtRX3x0uFwS3MP8/1U
C7ZCT2epYqfuEiTmgonoyEkUL9FZG+z/lx1FuTNq1EzYJKpkKW7vCZS2Xgvdj7uG
9SBWIbiyQXNxDXrUeaXRx0MVTN72Nk7k0QuYQJ15brmeI1TT8/9lDvKxXcDEtuLP
IORgpMEwPInTqkbctztcYilDK8JLgCJaDqZZH6K/jo30FYznIPW+NypgLFYT1VBG
M2t4wPzg1QiqG+fQqgQxZlXQc9EaH5YBNEX+1EANH0FDTT2N8VqfLnYjeyfeVuHF
JMXq49kgk5GE7S+VAWIHLBr2z+x1Vr/4HiXICxS9HlyrCnJtoHuorWKitKZUu1KX
OttKHWpN1Aj1Pnh7832crQ12sp4L7QZLm+T28ZqDrdT4EdQ9dRYbfOg4/M7XQyDQ
mLKPcxKb1zt0EYybS5BwOkRijy0YoLzkWoUYolxfW1/g0RWi+VpXN9vTZxHyib6L
Dq1q+2Ou5znRuwGDxf0U2iT/8Nc2cHG6ftqaEZujWjs53l2B4omU2vXNifrm42SZ
eceUIz+fCqC2SxIyD8DwMnaCIkPj6zaiVnFxUTuNSuOoi0YUiHrDQmXED+dae8yB
5J4/J/ua6tKYLHHC2gZRkG2s0uJIND8JSrdd9UxQtq7y2DI1Hl6Qidj6uI2ERd1k
Sm0VQKF7EbIWgdPKuiwwmqKMl4Kqm1+hnrfUQ8+u5VI0ZDuAxDq9RSFrfLqDFBSl
l5G8ibTG9N6BrYytsjH4VdCn/3GOM11gFW3DwIDSA0U9gzVxr00sd8qfe6kU4AUX
epCSyIxIFAjxHrmo1JkvUpPvaIq+9Kl4HFyCTLkU+WlNdDVMkIHL61FBj1omhgLX
1qy93ZZW2lF2Q+QVZAWIU/JKGUdaw6DhnnL4OQS6J7ID7JSu1h2lKCuLdNsRDL43
ZBv0a62rwdtLtcjgtEhKQBgzIqDDm5kRsH86oXZQ+RnA7kspinH+5o72vv3dFaMc
RmJLm9GUuvI8Qxq8Hqa2KUASPBNKqEoKNY7DeJxFWlig9uljw7gNjvG3IJN6hEnZ
sBBWuGYs0fHI5b33tBulScxFiSrfVO3ReRE/gqqnc6l1oAJgusjNu5elMjzubKnO
DVUD5vaXVjUVI25DrB/QUPs20ugnIvH5HVux7dfQk9CDM0C9aWCz31n/fBnwjPKb
rq2rlzgcS9c5dJeDhhpb0gDsBGfpXw0G8uVY8fXdXZYAK3d7Dg4+4Q0KMqYMa00B
q+uNKhP6+Y16inU3yEcSJBQ6onqRfi2lJ6MQX7gyhcTYx1qGWO7JNSdRRsz2GZ87
oZi3iytMRJ0hRoenO0Vffs6hV/MpPocQy8LL1dDO89XeQT+rb02LqtqCcIoUB6vb
P/j6VPPyVKfZa50YgHnBtPLJh/x6AQc2WEGFOAPOyYm56kzzJgDBxqMNQV7zyj3i
8q/D80jbYKiBB916LH1BNo5xnTbjAmwyd1vU585SJoyyxPrpTU1xMaiMISrmuLvi
nBHQRm9dvVM94BovbIyu7+KVEhHmfqppbd8LbxgeZbfyLw0dsS8UyNvQKOdQf465
0EUPaRjB+7WDeNO7dPbYgnJG9usz47HJiVz8wxlev6J3RQMhzn971nmBBsU5/9EN
gIPBBDdzFOE5mOOAfkbFMg5WnnKEBWcBfd/pxuRu9LiJFaAUwz87aQeDr3Y5siA+
ozdZX9BZ4PSWeoaBtd8zl+ZLZYxWQnXRvZJNXQpqgcSATtC5Cwk3jHvjf+rb54MI
dEuDFETB5z1WQBno9lg7WiW5/80p96SyVU2WNgqQU+rc7POm5e05CrHzMjT+J+Sk
nqK8UWo42Syk4umh0Y8trotXHdvNPD5k2anDb3VmUheXzDGq4ytXV57sLYZRQVHX
Jw1q9MU5Lp2Cas6FJxAe9fhLt0YOSQRuc5XHEw+bg8CyhRHu4XXQRasx0zrub6xp
QPxHHz0v8HHmUsBNPqRLX1ufRWrf4WqQQnq1DMlHCHBG2Tn5c4hjoYuxxWZWpSpn
cfNZV8uOKuD8UPFhNjVSbpEeRlOspVCvLOou3/i2ClgWd7bzyOgXvfCbJeBWBBm4
ycpa4EpS3exozwT701YwZJVCBIZBmT+Xlnyj7Pr/lL2KIJysY3BpkkBT6P6BYCek
AZFPEJNKdLiAXHmo/7xMpwSxrpglEvJbasAuSTKAj3pkWeA5hx9xQHzDdSe3s/XR
kaRRcUWHzj4edrXBJrWpOeunsu565lAW23AUeeECyFZMvmFDQMuSndpbvG8zVxaR
E3isX8VxnghERa2AG8NKw8HIF3c9+3EE1YI6wA7Lflk/+u07SVuZTBt/VWGaNvys
O7RKPcih6q6PCbnhAhw7xY9h2j8O9TcabCLXzzPAqGcxo9SJMHw2avEstgcc5wWk
TIomGhjmIl4+mU9EqS97Y9TV32mqJDnVUcuXYWor+/OKennOKoS7LmU5q2RKRlBb
V0KtZy/asFF77F9/6NO2Bl1Sqx2J84Dot//6wPFYeNOxLhSycl0tV8yrLu48LjrB
yqucrQvCUZBifb5Tjaj4xsN2H0JT/rChVzCn/2jEXNeobEFlUZDyIpqycdbBw955
4zIsURnSu5bStYaareH0lIiokP54wi3NArMcEeRaDMv60QJ7/janW+0u/O6gqOdM
8Hy5Y285F1FpZtIL2rZ+QKRkLjMi4QfAMSDS+DHJ3CyYTDIjo1o88nTfxy1AhVTN
rj8pd031kvL6rSU1J2GNleoFwZxcphNidxcHkL0sJQNs48BxB0VmQBlmgQP1hH4t
SrnCvsMLnVkz3Gco2t7jONj271uQxtyah2rMyVJHIeJi8rO5Bw4pO+ftMWvFfSIC
OmdJFhMQRXJQeRdTbMRpV8av1iu+coe9JEizkOWKimBUUZ8qf/EKHV+k7bpmNXTW
PuED23q3plqF0Qb5TPM7fOm26vwjrIaLdSY478ozWx1XDCZALRwiGTgs7fT7OxlF
sxySfnMP3oLRiYxLqVVYzjikC8p19zeNzRRZcpVEum7nSQwkA7mgvmX59AkSXaG1
AklIBcHRzRwUx4s1eMCk47YCSNoTak7UvTQDSreGZtxkSo7ZlgTuBFOcA/HF0BeS
RvbnFuLksbfh7biayYqLxaUP3n4hs5/DfNg0l2IJhPVhFMUWbnzaa0EtaMze01Vg
rE97i/6l4boah/QSA4XmUfDnhkBZUGADvTiC7VzA+lzs1SO5u6axOv7E0G3LU1cv
Iup5IKK3TJuEL/glBy8rTpFuRLzflfBrUGtu3glQhzZOismAYIbnpqzj40i/AwrQ
g+tZDilSMyFY7m8z/oR+frxDOKBcjBjm2EKEWMS3ITB52EJfxN5OPlzOcR0qSpiK
5AsyHN64hmg9/wot+RjXmiyhqzty0R0J70XZ8NDLJznhfx1oybtMMaab9MUMyGA0
qjCBfKDlKhKFGpy5zZYainelpSmGiTkLLFC3z1ksykqz5lCWsz1tTTLlOE4+COCh
TEz9Kci3zLGJbJGWua9Vy4mtmOTjy67MkzKx7OArbfEX1sQGhE5warEPMf8xVICW
bxUpJxOOoH8qyEDgfQzB2W/IZo4wggOTtRGMcr8kVYjDZYCPkCGUeVTNs32BMgzG
QuKiTb0NmktcjfigDHx1/UndE09jxZVhaFNNruvPueeF8K7gXH1DW/TuUpyz7gc+
ff+3J4JvfPU/EIhx+dK7VLWNc6VmSj9BIMoHEqVIfy8a9+jVJlLZeYSw5DO2NVmx
FquHzGqU/8isNVyldTFq4qkBuhqs2I85FxinmzIVYa1lXBBvKZCGd6GYxPoltI20
XHVN411nwzgQKlaSi2ncgE3bWhJKGach7+uF01425Zg7etGhLY9DPmH27mXAFAAG
sJ9FYUmWAFfBSpMBWhoveQYYD7GjCHoWACi+w5WWAR95iFNKJUliZcl3y4+RNB8q
5H6MboWY55xw5dMGwE1S0DLlqdmsG7+pXF80iz7uVf5Ad05Z/Q6A+H0UxwcmzgCM
XGDXv/ucmwTe2GOgbyQ3Upf0XKkwghwFolGFsOPArq1UOp0Z5N1o1ag/vOpbMr3E
CUXs8WN4FtZdTOiDJ0QdJouM9nw2BEqN6l+4OrEhBIQ8kEmR0KLjD9jgnv/cpnAL
V/SYb1K5aA4znK/afWdgp6VW+8A6nF0CSkesKN36xZ7lMlEsevoPcDq2uSB4/up+
ScdyqP8Bb4hap0QHTQ/5Qo3/Jsp9VavqHKFMzLfjbsH1i1w/+sHq7dtWyfDrJ/Qh
bHGRjOS9IbEQ1Knr8DfQ6mcwhW9VIwBi54sO2nBbSONM/Dh8pp9s5G6qT7PdfBMq
uGhaIuLcJL/4gQfTWJek4ccmO9J6wc3mVTFtS+sE/jssOJ7AOZrpcFGZokC9HGRZ
PQKx4btJ8y6JWFhxhKt4oxroAeh939I2ZejLukxEtT5J4eLJgtZ5EWqHpcJCeUVb
FpyCCOsubEkvizjN4n+fYJz+ap9lzKOHleuYrz4oz27+1RQqsMyL6/lkTSRLyu4h
zt4P+/yivMXXicwmOSweI7vTrWvAc0ZccqiH8GL9wCmtYgA9lDhNCZj8G1mHCIKb
MpYowpuFUBpDSSTllKc2XamdYicy4km9Fv1+lleU/ig46Nbm84fTXneo+WERQ5NL
p/R/8mocquV8kVcaJHKxQzqFbxWjKet4QCGRAT7N9MR+MM1j+JgDxTx1TnYG3okG
e3r3Ky47FxsblAm2DwfHwMpkL8rg8Joalde2DOFm9iLJrhDzxmxhXMZtaRGIm/kU
TBR/ApaHHiN4klekoTXFGd7onzoSBuHpyoFfITiP2yCKtTSvFKwyyngfl+d+Phsq
TvbCOer77xNQuujI47Q7WeVM5Cd7Q6UJUS3wdNmYVKOZ5ORkCOI/n3kRX2fYu5uG
rF4Lw5nxv20mVJx2Jba3FSVujjGESVau3hcYkEtWUDqZ16nS2IXVijPp5cEtmxgZ
683l7PW3x8r8q1Q7gW98AGF93RPpN3u/EcjAyYWjNYU/C4+rcZwLZKisR7xHJAFB
CKr/SjhCgmp8i19BIEg7YI6qPj5YNTIBzJSAyhwzygH22J3ScfcCJVl9rDsXV8tx
vGQ5FajsgurTdtAF1TUMoXiv9esoz5mNN1wfFiyvm78ZoR2WSPYE4tJG3DuQhzJh
eTo80/4lNb5sT88vg+EYlGWvJVbpiwEhb4kze0cdF2xeUtlAG8+u7IexMrmwYFlJ
I1iaJMvj81hE5sH+FkYRpLjUgKuFOKpS3LFUX7qF3JhGCr2Yh1SOYE7dtRNqsrfL
xCiYuzdI+TSvXxmefeoLlYrASEYRMkkci7nNG4kB8Sg+wMKKVizTzjV+HvMr/mUV
K+TXsjTub632heCKP6pHaQeKOzuP+LupckF44GxhOzMlzAtvxlc5BN8RBCTovXis
ZTHHybstnZAodwFBLSXMsQnT1habfgngXuToWNJKYfzug3IunyXCqY+vLzeXSoSN
3Xq9qEeYA5w4Of+SFU5l/YqkwASLaBY9/lYVtR6BsDfUD1wcUyZUfTG54XAdKbOj
5Dq7uCz7tdo2PDTX6iyc40uBTPFrtk3IbzmXZZEhJ5jJcvwjDFHgowTapti57B25
8YqNIKsyLBLM8GSbEcKGsFDYr6Gi8yR1SFP1Cu2cyL56OrWrqBukpoKg5bS//2/F
bLCLGxgcgoiG5poISsgLB8nupFFC/9pMIr9MJYHIPfUZ4npzgtNJcrwnGTGVf+aT
ExA8uFWBkdPMh5yUfsQJBrsWOKnPMQTpupcHYNE3z9MmbWa5ypKesSflfnAGVQEG
TVk2d2Z886b3rQARDmFXU6hfvW54+IHmaUsEZaWNXQL5qZ4Zpae2GOXaJ+M2ol1n
NrGtVszZU042E+geViYUS0JXlOIMfGdObWiWH963oPcxXtUWSbkqJ2vkO+jm7H0O
RFy3e91yfE0LHyjdbDEoTF8eNaA3q/fBPUBvsmO9Ddvpqj+3K1nfLs6RGSACS7vV
ft/jkotyb20s0398kgBKh2G1PMqClvuC4QR8XfZDfS3pHxvrtEU9r/tCyxNPRfly
hw6JlE73wixxg0pVq8FI/MsA9C8s+rThyXHakkQf/zKZLDhwlVmTqCW0R43lqxXQ
JN69sjl1ho3SPA7apDKTRasVWuClqqzyrBY/qdCJ7pTsc3boEZImBzEPFgJBKnTO
GvtB7aQxy7jJ1J+3/wjgoAJin3Sh7qsl2rhhiZdfyYJQHBZ1k49HES70ojl7qCNS
Eh1G6ZmpJU35w4CJ7U7QLAvgmFAGe5RvshLM31vHP+1h3edd8HxUf20deTXW9h1o
GS4gv8I/+cHlbzi7FxKaFHtL9K1rgJh2xs70qV4PsHthLnQs0aLvFYSvhHYu5pIc
FcIT6/Qho+o3pakjJIaX2F5ICCuf7Iy0u5ve2Nvd4L7sv6bn5eWb27+shubeGSiL
5iJ5O3GKkRM0M9nR1rNbEXH6FTZgljEcoaet7Sn11HZnQ2gJb5DqD9Fs3yvLtV+l
uEdkR8bYOWjl68BUJ6zOvi2QVBzPvIlEyW1KTcfGx74e1+M/LdH+uiiOjTqbeNqF
xf3E24UIEPr14C8mQQERnZSb2FSkXh/r4wqDC4gsowDohNIGt2Iy8dm3WWIa826d
GrAv9Hgk308OnCWsBhsgU9Hx+6tub3JGA2OKiFPEkNXa/bTID7zoiD/5HliYwT21
0Oyi1+MfPDAruHe6DThHM34XkULILbppV09Aw6a4Fd4RBh1FvqBnbOq7bBnQIlG/
Bc6vY8S6oyFUd2+8nQlCEV9MHE1Ghu6YLkTSU8u0u+U1X6vp47rIfy8PjJ+Zjuiy
Wsq85jxJoAjB9Yev5Sbzr3zWt+xZQxeE7MOONrZ7phDcpgJ23dApsjjxJnwDG2o2
b31jKb7KHoH5GcCEHlc0gvwJRx7dlLrkl24dZmRzyS0VX7Ki9hEMcUGy1gVzk0bb
rZhrWWEMGbR4kesuCVfWF0g74nOvJBLD/OGSkApjenEaVaGwbEm49oq1fu2yH/Mm
SiNkDrbCPFTqeuUzxl7F0qZadc/YoIfyK3YwrVPiNksXqeJ8zdW49delsTgxyqTL
8MNSTJKG3N6LHQQnbPTyp9fz9mf5cbm0zaLA7lqDptdFev/3JdfLWPzo1RikISHd
0ED6A7AST3HcaZxP4Qdgx5usZXksk43hQedeoqJKHMK+0dEgiwfkXOPWEjS80zh2
GfhYtfvkE4rmg5tJDepF6uZiKS6cGaF5Ee7kpvSHBB5WgQaMOQ+WKj4sUdXiJ0uk
FEzJcCJwwhVo5ZBIY1AjG4FeCf1qtkrRtQiA2GXLw7xIDQyjMzo+AR047ISftYqV
D/LIedmw0qtx+/tO0SgUCbWXD7mAnXEScrwvSRrqxTWMI4XBGdNiELfBgAoOgiiI
AAD+e7JpJhmoglTfVvzHzIu26BkwrRBoPaNhDWvQ1XCFPs2Exf8ts0E5efytiQ6t
3FxtL8HNCtKAiEkjby2i1wZF9nWLl6uolOx0ss8LnmGKFZRCrUYMvMRwBKAl4quF
Y2zDi38ZQVqxhY7IVH0na4KO8TNPq95TmN5Uy0YnKw4/3sVuXMOBR4FhNib038U3
f4x3YnNsc8JTxlZ/KR11tsAo6XIYwMTG/sFVguEbw6/bIc/Km6zC7pvDYL6UUWUe
jY1rHDafj6JUDuV4v73muFIw6e24/bFdWiuAV7ZPlEfEkAHB86hgxHftTPSNQY/Q
zUr1ygwz3a3cX7UqQVsXnHYYVsufTfYGp2c8naBRe29vLKsyEj6YwJA97QLg/Hm2
hBETV3ivyUBbCSPuM5IeWWg2qqjF0+tQ2tBmXoLUZahzob+rZAbGfuFHGRBFB3vT
D5uI6DAngI7OGL6uiCAVJdBIyeooj7/wi5H5hE7dfmPpbhxX55A4GKSaGHx83iz7
zH3iimClorMWHC8Pds5eVsPcuipUBaAPAYD+3AKBzjz79JW209v1BC2xEpw0cq+x
qjsbV5VQ7I7JbuFwHRc6CweXD7mjZHp3+1ecsXA9AR+LXsME2hwHDkcCHoWzC4f0
nzsVIULRxuNf9hY2ivAi3ONN01TbpG4D3ZFGPsQSkuWzC0XSk3baPLVDjK8RXvx4
nmERHLmyp7HNgLuDxc6WvnnwIiGiCmF+PjKTORROsjSSHwvByYO8ANcR+roDWq8G
Vhnj1B59T11qMY94xEStsvDvMQiAN7XQ6sDYHwIPjipcyyWCkc5oNntgqD6/MciN
TbTVyKG5CV7YKUdc2icPIpIdX6B+yaJgMjwQFhEA13Yp101+0LgrWmdXpPyxGwA+
B6k+t4+Skqvv94qQx9D3lm03LGWiFQ5Au0f7nCt2Ao6CgLFsQ+1ca2SHU+Xi1bjY
sT8Sl25TwANbVw12Zk0SlM9O4uqWQ0DBrazMBXpVAw5lENDTUkUfitAFVEZyY/H3
hQR49rsBYxPTNeLhepXp8rhvm0cybyMxHQR6PO6pVb9EyqVMfBYa3/eOoCXbK8p+
kq+Hrqlp+TDWs8EgsTJj8c7PEB3zFPYA+UGEo0p5SoF5HN31YNW0i8ekDF08Jg18
EWoQigCT4EP/b7cjjM2GQ/RhHUQyFRsNFKZHnS5ynZGfXuKmcd5OP62TWlFPPHbQ
zGxKQI+vhxdo16FsgfL8ATNRGPyl1pZJXG4NMDxmUKndjwvgAydn+PqfwSIyJnT8
HnN90sugsdf+ZVFDLrh7xoyDx7lZlyq7DXCk+hvNhvAqkeeDdMszxMJDLSNwLHWV
AeMy3TD+b+lVuP+FHmnwHYf6IXALq3jxlne4KHm0CI1hEidOekUCGnMEh9iL/d+i
5pVXxGBhKGjorm3wc1QaaxadZRPivkWdYg3HxvZKgIykpAnLi168gtsgDhLuYmAX
SVVm823RFoHDUdL+hsN0Z72mu81ejQ0vgVmRM7AY2OsWKeM8O2GWB62FtJ/S1mGT
TGs7oF29WhP3OOaVvUkE5VoXk35kUEpfKOt/ilTAGNEP9w03HAc7+xXAuHzXBP0x
wcXzVrPUw4VJf8FU0zrFhps8+Bt8WqC6HeEqvehJBMAq9c2YH53STmmik8p6NOJ+
PY0I7bEBZLXzOU62S8p015VoasRgUU8c301NwBQrmbAnI2TuQzDETIBiLLxjWnyv
zQnzAD2JKy4Tnq9K+TLX47hSGWc0SUayO7YMo6kpMhoB7Vn/7szY5jojsRb6fOE6
vw5ubEAEMUCiTKVxhiYDsvkAoJE0gT9XRA7G2VxnqTQpW6LAzalvkDpoZR+rbbNV
nuEjUInCte9Ig7JrdKh2tw605B2tzovH9prmqOoTDJ/kXXzKAzQd5kUuRIxIdVkv
hDK2npIAX7epo+ySuvhxGAcZtRzk8n5OtOMzVyrZdVPRVR7D092MbGyAJI8RfNjQ
h8tNWOvUtZgUsCHGYlX8kCs00UJ1+f9g8bTfFJN++BgCxf0XviWVVa8t4ce4kTJE
tpQca2w0PYHTgQpHRkFUdL1LkhPe8WDmK0O0WjkDo9QP3po6VM4VB0hWR8KL/jyR
E6EPpgVaEEbz5BbBrIMIaLBiuw2iuNXDSpbeLG55DIfM+G3f9UyKY1r0a6F0Kt91
yk/pS9Y8Z8TyhQPEpobaH+gPxF9WB+PkxbT6ScyMlX9kGq3+C8kszLGtyc+eXNpk
1EpQ9DBOzsKrdBSrgSZ+wQ9zRBdXD1c9enlgx2577IMd9yta2ZBSnxxPrwcRudUC
u1SHBFHtxVJio/QC/e7Ey9jZs7tdC+lt+kaUA4eMwtSezecSMZgAzqdZDT2Xkd4M
a3Mv4XHfxzK4V2N9diM5z7jdzlALrESgQANF9YTuZTSFSelIDi9AoD4BXQN86h2e
e209e+jzcqMvNrp0K8TiWNB6c4GKJMAj8VYlA9H/JI/nsgfsYkuqFzFZ2TKTOeGt
h3ApcTPIr3TMbOpE8IGH+GAwn85Q9A6FCfexV8lDYgHKM2uBmZgxtkuyWAH9utla
7I8FqXjrASAlczHa/WHzJozJBnapntF3Wy23zgNNw6f2HZ2Mcsk7QDGswffpIMZD
315+4uPeVWadU4gSYOjhUw5YBW+olmaArY1HjJuq3pu8Aez/WTPBzb7II5lCYjJi
i9wxxAsWPAFSct4de32vI/sWSSWXvMDwmrEVHIOYIMyA0bxv54SKu3k+GVjHt8cL
1ZGxiK8wmWrWhbgYsS5QMc0+4k8bbozdV3WmRyov+tanDkXgZ4aA1ZnwJQpCnkKv
8GDls2tTkJ7GTjE4pB5iea/1BGvYBOyVj+OGxM2KNIBJKRuTyS9RT0s1fqHWOGCO
GXi1lizTFR1mCgBuhgZ1yCT4vC2QmLMWjR+vanQpTwK7AtcL+7DA1yymak85svWX
JPA5Ye0eilj+pDPIUE6bY8eIO6SEijx37IZ9wHO9SVlTYpWNCOPKC2zVG9l314qj
US2ytJ3GI76PFaAEIIPAidVcJdosTu0PFxM0GWkSbZRUpLl7zK9msW4GWrZz8cpt
sJJ6lWbk6Wfzmi3ZwuzZu1/pyoxs7xvbUY6OKLKjL9SjJyyKmNw4sH8GwIT53DyQ
NoD7XBfAjnkE3uKukpFU6a9HeAR4o1lHa6otm/AzhKAkOpuHzgOQk9UNKCrTtRvM
XUMcNIZNUJIgveeopf2C3R0V3ESB8XY4Gf6atN8k5cyeNhlapgpoVgxzzDGAvWs4
tLNdMSB6ukXlZHAFZm7hzbasNv92GOgO0S4Lo8t8Er86wgOHJ6l36Afn6P661m4L
BOib3yqnCBycKojgLz2gCMBoOWr1Xfk6O9mrWpVc0LUiC8cnvvMvfrD2IA0gyhad
odpDaqgGyu3Fi4OJnwuCH1OD8fW2lcqtwn2bcgO3vkqxfClYwBbRzpO6pi5RXWL5
9SizdK7ltYv+U3kJG1BBpC29eZgWkVhS8c44cPLlEURTEF8XrooaS3uInxRZ5xpS
2Gaos2Kt6HNwCxlPZokxNWOj8Kx7L16VlTpdBswFQXykOXjgzgl2E77zbs2cSUZj
+0C/4hCJiIOs4wbyZo+6iSh2mE2230G1JB1DkwyeQx9b2VpHK6vMakocKQ/f22BX
GpSDkK7pSnCK12nhBpaOOSRFGg+yNMOhiYbku8twfuEfckozVW6wstPAb9qy9hBY
DAI5/bjpY/vOvNfWFoquu76V8eH+Nj37Elbcy7CXvfeVITQbcsYBZX7jPjwIdvQg
9ueu602kHippRBt5/pEUMKYdOgRczcIraoFEpaEE24AFbGj8bgWDqafc0pRAcAbv
/vHMLzXdz01wIMHL6mCz59gG55ZFazuQyK2VsWUOrjQ6TF5BBZ+DqBj1/RrfX7D6
oj05HjilAA4BXkiCGmIc9Cxt7XIuIn01H+9oPPXpv3iH+vydvnHfNOpchE72cTPs
REKedjcSBYggp/hXwkG5D0hPuOJURt8/cfzII8KKaNgRyarOSspRSEu+nA2P3z/f
3ELsXgyc+lrFtpo3dYJTrfL8YMP/D+xcBj5FkEZ1ZrJta+vAwyorwZNBpJE7U7z7
blXQLKWCq2Odyfda+zqEOSjEc+ZtAAyFx/mKFE+nDu+93zfuc48D9tbMycRIEvC8
8d7z9AhkxJfT7zb9brt4yrX8XS0okH5z7DRDYDfiTsNetkXtVJQBnij1l0wpw2is
PEecsxMVb77j9ZyJDXHzDasRury8Npblmpqdrsx4U7BMbqWTGHp+U+OQrnHcSdAp
LGUNJ5NOHkxbzB9bhI5/nGhmD2HSH0wKWUtiRTrEtuv5Y8W4Jjwd1JcHQZtaYkAo
o1qLgBfzSNEAxaUQZV0b0Ykd1IUZgapWcwBQm9iow7RteD6T6wygDLa5g8VfLrMg
KkgusrRMq44XhE3BCQ54h45JHE+HLW7J/Q1UzMUEWKTcsUCcGKdXcqtrYiZxemkj
oc9ZGAj98Ih/q4AAEd6W1AsUC/Cy622J0r3G8XYG7qrsk93UOW8aXOFz/titUc94
1jkTKtiphiOeiftV8Fk+WO9npusxFwTrsEeV/Ilz42zMM2ht4SfZSkFgmBuKlDD/
4mT4WKePhER6YB/hq10lCFeNzG8CFeTO6KAi35ZBRm36YdnFGzGbyJBHyYhwAaHe
hiFLTFm5ZwnsBwwTlr+Zhd4MsODjEeL/lmPWUq7BGiQgXePc5Eng+oE7/9V05nWZ
WlKQdu57QSSOvnNJh+xaEXvb6kNGM0r4w7cvDq6HxliwTkaGEn40entgETpUhtoF
JkhPacL2LK2+pSRl2bFntZuzlGNHH9lVyURnpcXJha4MDC8eOHGpbRZcIavsumGk
/kfNyOJuqdEYu5xlNU93gvfGzyM/nSPByJsy84GVhHDCVrQAHCSVkfCx4Q3GbE80
pBmqL+0VqSWM9/LsSWf30dJPq5FSf0/mKYZEURGEIzuX1XS55tYeZaRFE0vdW+Zj
yQ2X0V/V/pOSb9dACv5K4SlqkP07Er2OFgj1F8TzIoKKJI+fvqBx0sh91pksh3Ym
3YLmofbaoI+joDOy5utGGRIm089Ij1fsHiGH8SnqsSx2th/p3wi+DH1S63dUmI0O
5XHHbZNNEEaIc8oJ9WWmKgItYRhH1oeQgBQZ5CUWL3/OkrwZblHz2pzbMIxb5hAY
MKwBm30wp4bjamVww4QGwsYDoNNNn0DrNsVLwcnuoES7BFW2RjleCSLyJba+Gk4N
KdpCeP5Z1VGJ7T4Ldt7kznx4PKQlBqkAnM8Bk0jNQxtcCm8BNxApMf64V3iAUUUl
oYzs9RTMHv0b/YUxDHvMlZOaDiqMrjYC6JIK9f/HlURKzGe/E31Y7VC6293yAr6Q
XZHQpZNN9CVe6Hjmr2BjCu62hLP6Cx13JX2iXcXiBJnkn+NS80r2i+m9t6GOpk5u
NY3Dh9FT3GTLof4qHRinwGHmGJfloV4YHLBdghCCxHSimNwjVXhyHq6jZ2/tG+HK
2J8X1osJK1ZnS8PYrsQurt8BkBlnOEfCCYrUYaISUCoUNjz3zduRT8NV4h50sGkp
QirkQGUbiGVH2ggKgHKAyX3OoJrNgLc7oNp47+F9rbIEavhadJ7NT3KH0DFP5Q8b
QR1JGLWvATUHQ2VgkMNASWuPkNBKYPfIP1Cwrf2ystpqECAST2xmylggJ1WwQlxT
Uc1AL89WLByeLc+dG/+gs0EnJm4xuhaCk0wnQEONm7TDH5rUHFd4f3FJKnRYDeUz
e4aOfn2COz1xe6CXgv2f3lSKc1wZootIWALneXb4SBgeFcOA8CcMDFftKaTnePSi
tvEWtIx5XwV84F7tHfpgQqk/k2ozGoH6JDzR7E/lVP2R4LOjkngLwhICJ/23cJVZ
JPqJFOVw/UwKT4ybh2LVAMKv+EduBNLCzLWfOfXazAoutAFlqG048/DilsIYjJbS
RwjFiNXgPHNaGmyjD+fu/CVtdRTkeUDlWcoLFE8OTz7rd+Nfx9edLsRmQYrj+SMS
1fzCJrZ57puGrIh0h8MSFM+9AzZnVhBvH7hBjO51y9wIliGLiUd0OWRZJ3Or8yG3
39chi3cH1KmQLZsLBhV7Y0ky9UD0f2WUX4WNaI0eo5ga6vgK/CtTDZlhpW/lEH+s
o8DdfRxDd6w3y0gwuXSlQIgDFtqqlUMgCtuY42sXi7TG2BPo3ZAMIIt7DjcUryZ2
Nhd5r9Tq1YENswsog7v+DTSRpoE1atqRWnH8OncArCfF7is++zQUk66mhHu0sZeA
eyBRngm/n1WwSJEgd6bzjWw+RwLmFkeXGPGRV675nVJfFQy6l3CZiyItuXVpIDlu
sVvCtc/9qfS4yiTmLkUwlN0dMwdC600iJMiYCdhy8kVwzxxWGomkY3qsBP9nAynF
ktTFQJEnLIxkJ0qFRFx6x2F18LqNRHowjygD7kpV/8q42T1XctjU5JavYuWRgRPw
j6VqjsM4sRhh/CHVbYMPgd7N5TK62zioS02EY+0StbVZHnEWsz6toVft//PYUjcH
EjJP1ysSKHBTI175UNJwI7MfU4BMapGzAhCXpMvCKZgSR8rHz1iUz1SZn0hfXtFg
P6x8yorY6BW5jwbhacd/4YwNb0ITHeotgf69v9HXkUyvMv7kiE6FeMAzvX1dhZBD
BETOfEZvu6busaRxJ80UAP7uRf24o1hK7PrlR02w6EC+W+9uW2PdI11UuHc9O+45
bx0ikZG9XpnFCYnolXiLFIzilwB3xGk95nbZKY66cDzUxyD7kEM01pkIE4a2Yljy
13QbNn66Zbh+1UXUQYQsvM4/GOBAC+snNUUeWUZrObVDxhE+5q0bV4W7es5d3Rad
E6TgXdQEeCiCjy5QP++EItFRteHiSLFu1+4q/gvLVjwAL/6wTapvHnV81wnrB11A
mZbp4Nz6sivTdNm1hXQvrV624PR1Vu2OXH3mbySPbl0oRj1WQT2w+g0gBsYa8kyD
MA6aNfDK2G9QJ4G/LzyUz7lJJxw6Idg69drvDtJqC5fwgkVlUJ017oGG7y2N2lSL
BINK7US+Z4EkDumBLxwMWgWsmZlJbGp99rB3w4b17K5TsQUqdeD3wEEgl8dxsjh3
UdQb6533ZreT+37zu8bzivW69ADY1OcH6+W0MYraI4GEtIA3uDkK/D1Ws0idFT10
KfrAyKQtIiEn9UpoqunWK6PgZ7hu2qX565fs0c5xEKAJtI+BBY9X5/arEQkkU07J
797Y0OG64xU4RyhSa7dKe7R6wt23I1wER8CG10nubswpy9/W+pPhb1xp80D/kWmF
JTzElxU+6N3rHHCEVhjv6EcvqxPX4VNp4nJg2rrLiQdddiGH0cErUUKW5eNK5NtS
rLAeQg+zcM0l4nggHa3Tu7WAcTkGu4eCOLy/HpNzY/Sas22rvmukmbfaJaxJxeO1
2ULCiyM7mNAk+eV+ZWmWIAIbsr+LIb/U2Mrl4QSJE3UZLfEjSAofJTlw7bQ459D7
lIuFupoh2EVdcibMtQiTIxLfsTSbPC/B5BW7nT5k7USF/PKEFASY9fdFEjUCuLwK
rbCcGA4mvixZXteNp+dKROQP+tnmdAOqqiC6QK1trVcV4gjJnV59aSBhbPMcLJbM
7YTkKclefmZnBesx3NxPQprJvW0qgGFP6Q5sFc1e0RVNg4Bwu9FY8iCxYsiSoceK
HA/tI2hQ/2qx+Um5dNArXO7VHtPLIi9DRaIP/+uxQy0G489fgjIgRMkWGKD14OHf
bJ7Em2oq2ndVcbA2Qu/iORO+LMX/eEjSu86KNO5n1sjZvaR3IxZ2i/RZORqv12md
/TJh8pedtHsB9V7zFfu8guX/ZtoXz/m+6F/pdnR92l/ti2edejcYfDst5vw3VI7q
CQDy6duXf+ac5YuHGAgEtRUiTr16jOzDtDrYDQzkxICE393asAMlGr7oqWVnkv4G
th+9Nja84gLI8xgCYRDciKlf2nHLkv2tx6+2eXnAGtvd5tGlNl44Wx+c/J3Iv4s9
8UuCLFe6h+MxjVZaYe047QF6c4J8soRhGewsDy0Rpbo1e25rJgIHxmX2mYKmV9Gc
9JXRJezUhBXmViS0HJtSrP19uGK9YDxWJSfsKNqiYfPwTtW0yOoMBkkbiStqZp6C
SdAxU7M2PXAhdyCJEtDD9kcMaRLJUBgYyDgOWUy/n/K8Lhy1Lq2AKwTIB3nRqd8w
vVATWU9qf5mrHRg43xlLJWFUlVJmRapqYF89yEaJBsY5hRUFNEDSCNQhnoodbmJc
mXfs0FCSRBbpLk4NL9KnnxibFRlC7zkXvkw9w3eJ5PxcoLghcdH1GNJ9IXx6UNh4
Ypyx0cIDm12xZLTb/iHU7Ad7gkCaj+WOZ57SGXUr/hZWpXr9fhBkceEVWOueVyrc
fDPh5OU3jHV1QIgQkvhMcSh3r3p2qZb23bNzGE4GIPK73hG/IGmGQukLZuBXKW+w
8pvWDiucfVb0k/CNkcj/0g37hhcp+xVbMSrJyo3cd9at648EMtfL6AqbTatGbh1a
XZh0+FAz+knFYc4CDnINVK0RBdPdUD4UsnhaOJJ0fzn0Whw9ytghClvsb8933c/m
/z7LlFNLuOWRaERQ6b+5pkR/CkoFfw6y74j+2qOzWo6qg4b0zqMSbG4GNF0zgT8c
KdnqEC7BQ5ndHjO+Bx3CZ8+JUwfL7SHMjO29b4QR5D0edQQ1L4478AE/uXQixS3d
m8NzHVcZ8zC0Rs2Pk/L0tCOpNiKE7BlS3Yky0+R84Ugp7KZA4y4NLFGXhcx1nigi
hKU4o+C38Tz7JZucEtWM1hOr5jVz+v6YgW8Q21XDmBKdBp1gLmhp1DSspjRM56JG
GSECoWKiPmViD9QaAhVKdfZenONNwsj1VuwvxXlgZcVNPS+XopoWKyZCME0aKsK2
LJDEwxDaE3nn5AjoLfpP5NKJE6VTs6I7AcjJ94soPwXTsOIAS4dOloDxaX6LItoG
J105v3JbA3nA7GXM1CwpUxliG+HShkhmNzsZqD0DOtSpjEzl34nfv7qQeFmRFolq
keeL8J0+uOw+RLY4scKKHE9C6VKRHQ0RR86auzSeRQA4Y2C8jc9A8Q7hpmaEOpwn
aDRuqZQ9hJQCIxiX/pUQTu5tpnNDLsqRoq7H/+8j5TkmksdRGM6Durdidt6ttDZb
KMj1IGUdfJzmlDVEvUdVUvjZgpriB2vpBS3ncdSNF6Mc1+dpvyVFF+zkCh0sAXIM
aAvd3I9SDiVz9aBu6HFPVNv89L7SDhX2hW4bphNOqVJ1Dsvh90BDJsyWf76XFVZF
c09l5a1CrR9uMr+gWRNLgB552xpxgMrAeSV5wUzSwiq+YE25nd3vDY3NUgePpvjE
fSRY/McUvSfuiXr1GTrW5Z0bJzAa9hE17K58MmVrDIHPH+AFNJNpr4NcK4y6qlq5
TvSRtIQGGO/0GEBZyuc4Y+5lE59ZfWB/oayVIPu6HnMwFptreUf9vcklQNp58bmk
QKLwRuXZm/X6XaXJLGoN16Fzbjp3WCyK492VPvI0EGkvrOLjn4uv8gGmAHV84HZf
xblaW4/3zd7dovqE75ogft88UYjV+zHU1KyUB8JfR0hCBFfw574/bPnJW2mkWqxK
7BT/HIgRu9qNxcs+shGbLniI53KjYkKSOe72YY3CkvuiGKlju5qn6RL3EoBxmwwx
0MgqIexGnSxPIsHe+t7NznB3KpyVdEGzsJqFjklnFLmw9rsDEikbiCM30Vlb8JfZ
VL8mV9i9gdak6OVtgjnUWruloig70Xf6UUhPDLRKU1Q4w3pRnnnlQzTjLxnmMn87
NqLSJ7b4/oixorbokLutRhSgacMpOZIDSvX5TisoNiQngVgOwl57C5TUbYYcFWUb
Id3Ew6cRIpnD2+3qWKLU5Y0oMd0wFl+ItDIWziSZfoxzh+Rjib+KfeQJORfE1OJF
MW46s87Hw7tm+Mlwcbvr9Mc4HMdvBaDYnHn2aXagmCzwIY4tfB10peVRJz+l5XtW
egDXoYUhEYO6b//GCQwKFiOF2ctmZYWm3AaUkGjPlFAaakfN7jYHKbz06VeIyF7Q
I49PEBTONt2B/30Y9Hj1HHTbz/XSanBvgzAItHSTUkYsPas6hk8bGKBcaB3GR3Y7
N0YZiTLgkkaQn18ZU82a2Q5VzzzOjRKz1eJK16OehTDjGwAhClA2cikb08IIeh2x
znzZnyZl/ovmCsQ1HWyBynx4aisVyLjRyxAavW6hIeh7u3KVRlGzwDgkjNPgs/Yl
zTOCNLqsaaDD9Kt1sin1ZIvJz0BNyRwwvKfJ6HOtTDWBGox0GI9zzwN2tZyiP2tp
xMa9hIeKyYChKgu2Yn6zptxuwzUlt2AIrpbwW77+DNnO1AzVr0mh2qP2Y1vqt52f
tOgKZ1lArpq0fIx62gP7gYOcJHsIM8TcrJT3QFN359u6KIqOp7+5nYkVdXDyuNXT
AwCdqZfVWoKw6ZL7Yc9t5BmEnEGbw31CAH+uCwjRr8zNQfeyWDY8sNxyQJgWu65T
gLeHmUsKlWggom6Qt5qHwMdOvbn1/cEVmsUV2iGkIXAqpIZ9SAYv6lYIRxz2of2T
AZINLN+DrnstOsUA5lp+Bmhj/Hr9//mSeELR//HuVFpC/C+WcmnXE2vEf1Cz7vRG
MCbBU+WXpM2skiSsPJGhuF25SnvDyq+H+FiFZCgTPNCDxhN1sAfCjmNKRQN1qTji
hmbuimoN57O8+3cR/kOX96BqEDYfHef0iow2RXPBaafs76upFX5k4f8/EfZ7hKdA
t5VxhpEDcoqv2QsuPcUmOyHgtA42MGY9SFexT6/mpYhmE+ZADBfmdm7L6JqyIsot
1nuquOea+i63hb42QIYJDx6szoiWfGIBpEXOCzOUp1AwMd8jSHpiSGnoWz4j/wmL
CFQSjXkutItZM/2QdmZB2EW6WaxFP+36Ufk5qGrFuEuBwDet9/CvR+nnbo6WSK31
7P1RIUqanbDaGTyWxycwnid1K3beb6Af833zKAaTQt51mXxY3wHmwZuYus4boeHf
DUWuhk/Ufb++8h7MjElUZNH91FnqPD9cYG57xEv/ePxwXSijNqdb9PYBxwih7dVY
/7nJyGkznGKt8dlccVd3Tz/BZmykb+rOOKFwmaDjwy+jeYS1qTRrhXcbfxmoB5+0
mkZMJBbHYphh6ukaIuDD8I8noxE7u0p9holBTJQbzjLoKnX5w9++JYRxXHziNDwD
roTzz6ft/uVj1b3RnkzzZHfIB3CBBuUY2twYuJ0/Vc7kSutg1dPie5qKTiYrtvSc
T6UkdJo02dcnjJ7YTR7h1jf5MlwKnQxFM3jujZqNucrPKMMFSlJk2Wz1dGziViAo
++5gJhD5btm7FjZ5E/FFYm18lnwHuFUSaL5RvbmScxxJgjSsY0YYsYALpph72g+H
f5MLJFD4gqr22KTtsH/FFnDf31WK4ut0OA+Ef2/GtXgGXozjw0Yzf5fyFPlMo/Rp
21b87LC8yRFB6Gb7P+S9gLWYBH21vPLmA2d316KKoJAdq74/kyQNpkwxMBq76097
NsbeU5Ztnq9vqTR4mHZGgESKY1NACTDW6yocsI1TPkzC3PaWQKLLJIYoEC3IE+ei
AEVggs5cIAvZPEPBJysGcgGSp7L3e5FvUUXBJgXOXhK2BaEg0QU1WLqrb14suNN3
GgOoiqeHtqveaCrz1JmZXW2kcAfJKccHbfbXfxm4KYAWjryxgWm5CqkgYFjRLiH9
Y7GW94+EirZM8pMH/Z5EJIPs0V8Wk00s2CFKPeC2ktlKkqppQMEYBY/FHoFOR3Wz
BMxurTcWZCVVGdBHDS4TdKXf5jgDg/iLJnvKu2zDOTh/RFpQ/chYhy3KiT4XVaLV
/aozB0jvM2kYJUHH2NOrNFo6bqkzYaUGTZcJhMyqK+ynXZhOmaCa/lSqaX8cD6iN
23ie/YrfYXsA+DS9JvROQLnAuegK+1GTc0zVcLKcPMNnpTrcuU8Z5U4z/t935KNo
Xw9zIj76AEQvehOA510z4MSct8gswwb2Fg1E4m+vKT3KKcDnzzJAtj8h1eN4zm+a
pwiFbM/D/GN+dhGQmp9bIHbyXyd23EN9q1NsrvbJDk176fjMw+ftq5rm+tQ9xsN3
Dl9xt1gfDKsT/EUdm/vH6y78PsrcfIkrOL5ig8Cusv7+FE9V3vk9xNs1WBTziQ2F
IyZyXqZuMfIJa92FvMJvEPLnlsXE/y5BMm9zX3I2VgmUz9AF5cty74XBlZwYNa9Q
aXmgI+PfqRUd2voxZyNscfdos533u7AD6c6n8sv4ut6QzpYsmsGGuHlyQUDmyySW
KqiIoAIhLMAuuNg6S7/mOsFl8jC5okblTItT1rtl5jFt0VX5ozPb7pxyijfB7ozu
Ma/X+Qa2WKqqdaMkKSdCTUEFpzj+WQ60fWAm1g4c8abyID+58htl/KymB5lM83Y9
Iv7D9j2PBx2oVHpXQNCWCTwr51PWuhlr277Z7UzGhvWQl13DS8kGfTnyEzh52P5l
QuXIEvUenbrJARMERh+BZIGZos93T0eFezEc6br/awCTTW31l6UhEm0lJSWtHfoL
47OQsnoOvGnZECykhAoHNDgAKnmEXKgc2wNOvAkVDD2h1XxYC9cIaY5jmYxyVTgA
RhIqC1MIWtKRLt6gMmE76GDehYi5FuISI5jT4+REhFnCRexm+7qH6g3tDrImeQxf
AhI1maDNW+Tn15V88RBMHulmquQtn7EExzlmWqrteJEZpZRLZufIe/d9MrDDXD8K
zaVU+nzCHTXQAbwT+Rb6tgsnm8QLvbhBtKDYCXbY/2xzEhe/qLE6jWWAzmsPI/4U
SQ6nO3epTqBMCfV0mXz/frqpDq29tYoDv24ge7V5vHRZRAmGKvFwfbojJoej9b5b
gQOIPU7yv7LevJXD9Ix1UVdWD1sigCP27GxCzAA7tgquPyCqoKlY6GgzxeQ389wT
XrlOIMqYhYMM3HAf5nPms7WeFQlUcbuY0SK5t2iXvF/CUOS9oM5Sl2xOjUXKZ/eg
hZOB0lMDdTX1qkgaG19llSjZzKTsgBdfW8qRnSlR24udzVeuB0tpNYZlDzm8sjj6
PAl9vysofIqus0ucfENaqCAhBQGak+i2D67yYfKPzElHI897gLV2Kjb7s2YCPG21
Mgse0nf5JKAGlXE8Mo8Cxq/ZyOwr52xTaHKo32K747fX8EsYM+mmgmbSGfVEPoFr
3IF7hsn+Sgeu6aiyNJ6FLqEieJO+fdJvNuJLQ0pudoBvX/GDjDME7VZG29TuxS+k
69VjisrNF6kvmD1Cvt18AIe1Jbdj+6CJTM0l/Mn4w6+T1awo0a3AqW5wPrFp43Gg
EX3Vu0RnXv+/rz7RQwBlpSCVvNQhIGc7DkFakUz2KneJhTpNsGBhzbDYzPuqF/Ib
T/NTyvhYCBpEZx4XW6OwWEaH5sz1EvaziMGxDy2RlsAxshMotPQMUDmrAL6PpSaB
Whk8Nr3IUGNVdJ0QNkfVCy33hbNYYAw3x9sczTFExsw17fvMhTU2leO4xd5RS8ae
r5hT+w3Nc68DFSFTO4QPs2FmEtsTeIt9xTupwAE1a1TwGTggROC1BnzT2w2Bz2A0
aurxwS3NbO3Zpl++ECwOEy60MkI17D76Np0jfCD9XbD6qGc73dDjFR9ew3d4W4AY
CrBt/3Ke8jhiNHuuZly7x1yKt37WfFyi81fKfvfXV6iQiIrGcx3IINVyM63ff+zM
pVWWoYLKUFsES7bCEgrkFUas1U0a24rVArvkxZD7Y6htWm8N3/pyt/u/y1otv5fR
AQiRDOGzLpPtso/Yu/0SUf5KLh0KEVz7i48eoYimZqvjSF1W54xRCP4Pn/3AhkRF
HmmoeL5MLK49f6hUPgV4Zam3/aXqb3M0q77VXKxoJ0S1U3wtx/I5i/XEKXFIWVFM
F+UmF3N9GHqzrQdL/op/s2Hi5LwuGXcUklkz+KOw6SS+UImmx/134IjajFKpDkes
lgE5l4rCJpTZ9uX+bV5XSdc98sV6KoFgMnJ0gOt216M12DanACzYZwb5V49tkqxB
s9mtRSoNWZbd5udERYo5yly5obKLcr9sh7EE4y4A6vSWqMEkByEb89qpqci6ytrb
XBKsxu6htiwb9Fg3pIMk/7uz1V1Qw0NIv16oL3rxdig3kn3d11E6oRNo+Z5Ughzj
Bf6qwNeaNARgK/MPZptFmAJiH80NZfXaRMxMOemhPJfERfVOx5iOf4ou7G+viYMF
Iy1NpFrdnKnsPPc1lIKuD0/DG6q3CRnZM97fgA+vaeKjMg6Q7Ad1fRdoEuudxC98
m4MclIl5uDTzi4M2EKu91ZvG3kqT4tr8GQ1HWCDmdVU/UfR0TgOPQQrur+c3YsSV
M7Dc7LfFSyU/nXK9wHTcJMbt29nGYi5YfyAy4OGnbOhtmMIeRtjVwUsjkzTYulHN
ZJsowtqPgNekneWZgI2yS6He5Nha0vE83drn8VSTCtFYgUmkYhtnhUsh74FmYfae
pvMpPc6pisUksqAJd6E4BO8gWhqkRkCBsgCVd0uHnrLHEUOSS8nmVYID+VSUVHup
7EWpIXBcE86BQHEjqp+ICbRtAcQUWQ3XAr41+amq+/CiJyPF13d9sgK5aO8c7SUw
ZLPOP0weoPyGCDfDrc1BHYRNaqHn7QDj2hfT52Wh9O+EIjWt8ma75Sv23Tfk72+0
uE2hXINGjKX/cdeMSUAFkJ2TwT1/HlEVV9Njzk40XlIDv4+7vPq3TC7+VUdvXAjP
jzYqWBfuIGhaSc8YuC/86vVc9nco5tXy0kNkD1kVrZ23e4arL0+Tb5slDWTfKXde
0QBM+5mVy0MMQzWWAKF7p8QJN5qu+AQk8NIgpAHxtDe6aRwLbtDdossyHwCXz57v
99gKZ/M5kwT3f/O66YLv1U959vwRogho41WGjiqv76ImHj+hTsn5bnf6qar/INn6
ew7Fj9rgkh2QAh+V61fZaj4Pi0UTTB2+yVWYKc+t+2t4TATOgHOxsxN0vnJGfIGd
FgGZFdAnNmylVFK2E+7PyV6qQXoG+5DXc6GVj3j7xpK3zA+3vFFYZSaI1AoHraAK
gVeS9fx4w9KYfKpi6TaATqQpl87ykigjhImEsfmYh4MKqKs8R7V8DokS9oCDpdAZ
IiXDo2p19Z+2RQHFuvQ1eQvhpAS6g0T+lZAhN6mGYZfJ+MC3mDiR6tVv0JOqZ5x5
K3vBhI7qztFnMJzxt+zyn93CqLPYFbtSIXY07EDO+ojnLBVHZKMJHL8194kO6qH/
pYoAgTTPHVogY21UcCSE4KRD3ggZJ34zqPlIwduMaGIblfniUCghISr7nW5NMR1Y
Dc86nFEU8YozJsg8a7FymjhuPCvWWiVRs0WOV4uDE7JKSyNgOJVCoFV6GuuWVEAU
4/IsU2g7ztxkXblxAmT2ek2jFxbjeHQj+6l3jJLmFS/wp4+bZG89nG7d5lUOwAJI
JmpVGbLl7++LIQVl7rP+4sKiDeXvyb1rC4q7hay0accr3a2irvWkAINsV1XOxivj
HDIGoDEdxfh1cBr6jlXe0/qJFjcJbSlQQK8bgLA4rAYCrP8dfRqH8InE2dVJqeRZ
9NW3r5qn0ByJThvYW1uEr3+VG3TR4DNOscUXq/F3Uyl5glTfHiuzXYLwLXqQJoa8
xZqRUA8dL847nYiNVQhpvhTxlFDEKmHGPqR8K44i4Fa0CXE5vimSYLR/UWjFjUVC
33dpLViuip/t+hYoEo9L6WYwTuMa+I/EqSi1OgFNIWRfo+7XAsYwLnbxlJHAPMjO
hC48qHeGlar/l0YJXV2k+ds8NctxfC2Ej3+cePengGqdxtf5M94HUV6Iq6iCJbc2
4ps3ECyjBJGXYZvzVqLz7pYM5kku01+sB+KWJNMwZ/wEi5sWnm1/zXlgLVZW1tCs
ralyrdMmW5JmngDdAyPwIhAQXHO1vIvCUIT4VCwh8Em33jmi71iniCxHFpytJ2Jo
TIZJqr4DvHmz4NQVX2+XxqPpDnbTuEevcZnfKtWE/2trOqmcuN15eR/SLLWt+xGD
57rT3FGznGVPsPcNg+9cgmNS5tSrBsL1/rCnZvvWznqKFXj3cBv2h7mCOwel8e6T
bNLF9lZVMN5aZeWyvzDm2mV80M86EC4e48EE4t33F2GzShS2jZ6QnP6B74y9hULO
liQKvMvcqvvUJ7emKFw2iTPBm6F7swugFb7JD+oK2+du07DyiVAFxnfpDDP2WycZ
4eFm7FTrurgWBg+iVgaKAW8CMrF1vMfR9DPsXLRdiwcj5YKwn93Q1u9Mvc+8DB3W
xFnhXA9/pO6tNXModIZvdDBZNkMarr+azIpeN6BTh7B0WdRnsZyTapy0eOBawsRG
JWfoEHX/iHuRIf7RCiIstceVvB16kxmE2KsVK5M2TGLzQYauAcjHR0DRXaOmOPig
QVqN8z49axu1jtjb9oY+0qkK5duNz+CCcnfKR1fIa+CEOw3FTfjBnd3KqdeQL4HY
SKxXv0r901H0j1DkZ/goEx0xliuQlgK+oS2cDvvKAgeXIQ6c7I09SMzmdwYWFtq1
Msxs5Xa7LDk1bLY6ja+waz6HHhpq1tdB1EOvU2EhfvigzPyHVC8olC4huGkioQHi
gDbo2u21qEkBGiF3XMwFMJerq83UaZhJOE3G0bL3r2K3zFJnE7N9vjUhIcUFmkTo
WRh/+x3Oy9AQbKVC4PmxRaH5va17MefXkclSk1OS6TxqexwtVylmdcQkdtvvaDiT
GzZRX79rwonuFMY0Wy+YJQ0mAxGDJqitktq7AWyYjfGzPPrtl11UHml5xctkJFuk
Xc5C36vLN0TLyfNXW4yg4FaQXEJGNVDE4dl9WxM5X21ranXom/2I21ppieaZ5hZK
Qd5rpsESTHP7z6baS4ZdFgYmQxam0V1lF38zFoUAiRe3Gbdpx2dwkADo0o/ar6n3
/vYOj76AQJEV5aUfu/R8P24AVb/Dju2m+uyvuTx0pUabLCBKWPOOSfd0o1YXKlMF
cWMs7e3c4y27aZAM2Pt+ito0f5l5UGW1uw3F6ugO1kmp7HTHVQhvc5zcBT1ZMibt
Rx+NmI3qpK8DAFmLi2zAOQTI1USHuKx+s2QdD5pRBMRq7urk1amo9ZcKgleo/wei
ovOcuFRgBZ88YPlNR1JpkNlMZYRufWS0uYzwt2WDDxtdXqtNR/KEaIP2r0OXHbv7
wQpKp1STMXEa7rD7l3Ms/OvZlQ7zRz1x135QGV2Vu/qN28VrlCKx8s1lbhnxxH+D
BP/mWMnRYaBasMB/iFK2fbHGaLuy5uV4/SgcNFoZkH0ga4fWvN8odbXJUBBZfUFD
fhpQc+WwkCLpkU2BCLdGl9qCWenMQtVo9Q8PDzgBLl8MvytZaep/bT21a/5PyiZo
oYMll1Ew59pwTdOwSkS3I1dlyy5e4wlq2OkOmqC95WLtTb04XJr5LHJ8KzwrlAXw
C2ZbXIlwOb1W4c5iHtVTnXi0q/8piVK2QbU36dO1fX56/hnh//CAKE6XaoGnke81
iPtZVJIaUhc4V7Xpoj6oZzb17IhFtfg1W0ba4gUs8YKWlIClWz52oytuUg56BSvH
1OuCY4IohM28XdYMlOxtEdlvp05P5AhweQU7s4lqT0qR+mRdzs9dRflSS99s9IMF
PZeZFGmK2OeGMVXZ2WQhx/DQlUdq6ID6ggBujy6K76yOK64ArkCfQ3BztivO0xIP
f10+Xm1x6aU7BuQP8ufKuNoCngmkidZLrBS3rjBGBkg53haVryYyuDiJWFDdTM69
UH6538t7D7hP1nTZ/p2gRR4sAfk8KCaYgacR7KdKaYzmvGMBVdEpXQu0scVm4Inb
E3SNqBk+/S6tuKUY0ByAdQE9nGGVZkERgbvFkXEogMH9m2iBDXGD/yfKVHsfsQRn
65y0gLjQgBlRIr//F3KVVwmAMC7NCddPt2lzOnsvwjV5XawoArDeRgzqzGKgzihA
jenxGM9wcojaCA+YUMjOhPQwpunYOJ+m/PxgDye90wh5rwqMhAwVRfxGf3iFHuWA
5GGb4twIzSLVDMAUMbKucMCK3e1yxyGCN5DcfVDjq6FZXigQuB2CbljAEjeV+n9X
6/V3rJq2lap/tFL/PWh/dC4WjlN2AEbAGZZJ4qqxOby+FR1Gwub4vYDPoFjj7hw6
eMMtY1aQC+rqmREDB6prxNXKGW4hXv2UpmA4tmPhrNADcMwzVx7Rnb+XCo/JtkES
KU66x/NEQLVglNBBrkK4usa5oVnID+lmI0sLoTN7j3sBvuvdH+L1zPJALpxIY/Jt
PIZexiwJZK34U3fhR8qlFKS6rV0H0VG7YBn+YAkZehXO7qOVezrNVu0k2AKCX9c4
7hQlpzPxkqcsk/heLWIsYq0GjBhYZJbyieQ7z9vLInSW+EazBj3MzUtbBn6itjYG
D6oOzFq4SjRMTVNVPZhU+2EVgfKLcnfbRbBrpIqYssgTs6CFZLq78wb5dX5jdt4b
lJ4oGaMUrGjMLzE5Pn87RCJWLon2TKKb4P1pmzVrZ1AbNQ50Zsy0NEKqrHVAtbe4
DuNeV+6czbN2BzkBoi2pHFfmwXLGbgfiWIr6gvwTOkg6fnuL/bEmy9+eat/JPIHc
DqYg8eObSa/mFJ15b4bagySyxIuL0b0oVD7a63XtfqtzvWe0CFbuL9LS6+CfJcPQ
5qT+vsU4E+Q6AnqaItzj9fGK11N+0xjzJNnPbFJymRMVp9n3BNfW9IJOogUI4I8y
yPk/0P3KjKKmvjagiyQDy2CKC71LRrHTW+pN9WCRlgTuKilarpPJVXyMfO9jdva9
xxrL6QY7+7VMNPihoBNICHQKH0GrXnB8o4fgmXfEtTS+EP8JcCkb1F3OMZj/DiH1
u12hR+TXs9cUOeqcKYNz68sDrvQqVoeMyVIc/66fH2FhnjNmKBHA5yx9ZFBvPu4y
UNF2Ym7aLm1ldurxXhfVPutUBfXTsGgymJre42PiOuRVsM3LWOTrrLXr2YKbSqrZ
tAdkQlgkKWe3nRDhHXzVWT3u2Yf+u5NL5WhE5dvpZb20+TZoUrS3zV0QTtLBsYE+
k5Hux+eAFPkGYd0C11qCNMulzV3jNX4MxvMAuu7vAzajZa7iBpb+3SaloExAUg98
MRzKY2EHIQvpGmiSdX3xXxzWFJ+EOMKJEMieg0bV7lMz+wppft+N7z3kMM+7phLG
Rwot1HY3zkRX+ipNMCcMAKm4kJUdH1keP86S2dy/dOCUV4uJIqPwkpy/AxrxMAGf
RI5mMe8mNC5aCi5efQHiiXpzwhUuKmv52H88ZrrouZSTD+8YN2GNe3sfRrD+E+jr
p3WPI626m2Tefq3H10U+xn81rHYZEgWRMiUpuiiHb2pwtFVrTynXI+Y5nvuvGqF+
Ny3de2+PyVx9eEfyWcDTeCbrdYUY1ilH0XDDThVRaM+/aWTcXVxXcE5gaq8BBbZ+
UTcj01hhSF92J/4Z0vNDLyt9XhBM2XMncdde8rVddrvKCwkn6g1QfRhn9eW6kviG
oxN/yKEeMA6zKEv+glgjqHLoirfTlhUXPRZs32zcF6LVl7p6Ao1egdu4axn5L4NC
A7UTaqPRlbp1w5oapHsJ/gNZGFPv9JF0/jD/3kjHkzt/QdTSIA+Aw9ZzCiFCRDk2
UOKhTUYo6sFxgiA+MOEsdmYHbTuDnp1g1OCOW+GcZQBxSkoOdeGsj7lIx9JNrEBz
pwDA4qraz3Xq66RwmmZRIh7n35A1E2+HqsHhYl/XmrW6b5aDOpfxiCYwXemGSkJA
W/2pJcbK6mJYYMvpCz/dTc50mIHyzE1HHSKHN3nLMH7JLecpxipbqqL2ts5BlVh1
JnV2ruzVa0WX09STuwqPfC3A+U8uENfEcTOXbD+ATGEEQ1IEKmQKguyEFRO7yFSj
Q9EWHT0nYSWLpiW4jVANJJ6/cEKywgOvXx4frE9KzCgc0WbPs7pKKexco13jr2sb
oFC9uuCPSFEtkviNraLzCKGhZdfbJAPCKyxmISFufQy9x4czpAIIzbDlLi/HvJch
AlSi4ORoIG14MQe+389/kcuO1mSudpw7eh/PoQut4yx+r2IlusvsiR3LVPh2OQKC
yu++iwFEUIufGFFueKpU0yJ2eZhe/mb24zU4nV+WOUQRYtdTdSxHg+YaQf2ifVdY
4rXKpO9ujAAheGuYzmdSEw/XCYTOh29m/N0T86yrM+seJd4tv3v3f/N+9nv+k+Tr
i2Gbt6GWsvuoBOtDvg9OgK+EJOsjUTGS5JXdQ30/nuz2ieHq9uqq74LLhsXRquBE
ZU5+ZNTnPXyPNYloebmTptmaeoxg/Ki2X32pqxv2fp1UM1JRrRPpJah3SeRmEDpq
rJVecefzsn6sgD+gT/EQ0v8V2ZMZIGwkH6n7IJWQXeHmZegAZaWUrEVUA9CTowwO
+b67khYI9lsH+1jKVee8c2mdQKWqsefucc424SUekMPNhyq50aJdk+olf1wA3yAE
3JiX1V28rhwP50dJM1PE0/xZ1XmQ8uV80CtCF1YN532AsmeATg3f44EAPsUDv0/O
MsVvPnpRNRWzC3/fIv8hF9nwcK3DqeUG8jQlxmXSFm197UGWfkMbXk81i2jOpIbl
KXUCNzeTfQeGf4IMm1tfV/SjM83duK60Hef2oPqIy/0aD0otj7JGy3FbGhCN/jjA
Q+oBNjGGadKsFeEioqZggkZlTvcfDIvaoKgNcjYTBZSZifA/PPV15/FHYN4Vkkh2
+KQz8GY6/Qe+M5UfHxonEqxdGM3iryAhtz7bvi3Yk4FrkIjuhsCrSzE+D0isVnv9
ZLGZjp7eTU5JqcmKPRG4JAeeReAgze41VfcggvF/7ZgO/k8DzLd1mBcup4ieQKwV
01g8YEmLfBPYnmsIF1n5D/OZwaPC91/bFUQ+frlogUb1Egb9IMmoaiP/bmEPSQE7
RhB0kZRUSJgmLnYozV1L4rl5tYXYfkcI7Nb5HBHhpptgNggZKF9LvB4Ot5Tcl8LJ
jc+C7zp6F9sCVPkC3a089wgAJEgPjwciDHiWWaUd/qqIbkoHNwQBYzZyAS7G7Uof
kJHu3PkVlX54Xgbv8+W5AowpPxDyYIjll0jvP39MLrXvID94istrgG/kclk54lKg
7SeF2YOE5CGpX8gRno2+diubEsoUwd775zenrefwn85kWRPNbbvAmMMDiGYjUatb
DS8Cd4+71eZZjlOrj9zM2Yaqk/11C/kzZv6Ynw7U6dqS9vfuxKx8Dh7MiSex8JYQ
Iqw+Q+C54VpL58Bu2zckeerY2oIA/xgqpvkj0Byj/n1SJKp1hSsGPkkX9UqBC69Q
7UlYKF7P7zrV8klPLz6YGxca1rZq1rbgWjtV6265JhrLcZait0JQ75OO2HGPkiMK
XC7pVc+VseXVMFfScUUmC9/5YEM+Omy7Xez/I3QpIoMOB6QBw3n/Bu1rcAlaw6gn
1/10zUUwsYN8Cbg5EsroRKTn03KgKP2hd6RIcaQ1Hr/5X6qVuMW6ZgweBkS4KJ0l
uGVJyvD3aD+twn5TCKA3WIZeobvIjI+edW/0bx9CMcaundBNv0eP4T0c6eNoZRF9
S03/ABUSXVzZ+M6Z9AIGN1Ce2U3BLPpYh1jwgqyOeV10wD7TNue3nwHkOfsuFwde
H//STRxVmROyGB5zJ4AtLVTbPZR2czr3P0l1kSKxqvw4Wo6JrHGBAc7+IHoaEKiN
J3HK/EBo6MKmobIx3t6VA0/sERb6hlwZFzV1TKyhvF5vI62kpV/ZQQTvR0U/QrlX
128cfEjfrd4fVZgI4nquaYKQLziQNvbdJEtzQhDf6/lINyL4E6uks/MIKcPbhKSj
Ea6e20A4GpGd9hUlP+seHqsdMNFLCTgeculvliQSzVzN/pqQOtto3EGeinCOvu8V
/BiHtFuz3zK8Sr9m3nZeeEee/fvTg9WwFE5gPM4VPpFp/Atx1YMpidtMBKwb496o
UqeHxtUOtuN1yID22aYdrmjrVV9YX6+9v9s+3KlMKpsa8Ibq0ETyFJ1Ab98hrfVv
UXZ5C9w/KPRla1hpaUFrwgNY7R5eAp9Rj1+tihGK1XgCzENMfBfgBIKYTvpitCHA
EOlt9HwdCr0MKGmaYNlZTYSDZGz+tFQ3ZKzwZEYqPYvvB1BOCk2hjiKh8gwPB0+K
wPILAbOapmB8cyXQrBj5QkOxmXoBHdGi2i8wAudOL0+8GS+t69v9/PKMRTOO4VG6
t5tCcB/DUGcXKiyaopiZ5paTuqYzBUqoj1u94STx7yvMH+L2AOD9WsZM9NuSZA5x
v62RvjLpXMp8zPLuHu83xV9DaxsuvO+RmfnlUmvsqXpCUiYxVrXW2faVEeoQqA2E
l7U8W7l5TnBA/3McEo91YQ7gavdoY/dbWPu9PEiTSxPCd6XTi2XGejb0xQ+ybq5l
xhGxSuwddWdZYdUxcA1oLtH3+TBUJzUAFt+OqENoMqaGCpgkWeed1r5/jo6zks+O
qvWTap9CcsO620eaMXXR82hF0RszU4WI9JvV9FOGx/qwtyeJPUrDSLu4GIfkugZf
LD651jXMsj3LF3yOaFpjLbsk9G8VwqgRX/BfLRH068OjBOJG6mXNp/3Nh027o8bD
FP8XaH06bsKEJYLI6sIInaoWhgO/ea5MOKH2r+CpZhTSaQWfXXf2VlZ3hDQ6Phk/
F9L68wBAryIaWx69iXO4g6elcWl6PH96iEeDnLklMdLjKQugvn2ryMbWrD4K9P4G
AMgXD6e9p8qqWjaXs0ZtcggOyff9gHBaR2QgMEHPDFk/k/gCPKYP+r5ISDdFNqoW
eBoEE/yxFpuN+zIkjLWFaVi2J2H08lAux59VPONXDz6as54760x+Z3Id8NJhJWkU
c0HDVr6womR9qgOJkPKynB1GQ4HArlO60zPfetMdsncuM6bcNG/PlWQMJUjNHEXP
f4C2j2xRyqcEkFuOvpghq4YbTVgeMn1D9PHzDX7+pQDNFhQHTEnAef4WWPo+lHWN
jOLj6o5QjI5euZzLEPg+E5E+3qXSZvoLwEPLQGM+2dCNhNh1rBdC4GexyPrA8iGg
N0hmyHUTx6GyFuRErHAb7wvgTo37MAGm0bzPOGLmtu7oP4k6w7Gc/WK634lDb7e+
Bj9jbdnl8W+GlUlk2D66LwHcpI8RhYn5gdM1aLVrnv1Tfd24n7HFE33SAponNmGP
1EAY9HbzfBzVQeH6gMy4e1SO+Yfzhr8M3VhjQxMnKkbKiGoIy6GGdqJnFMpKykF2
ePngEcoBsByLvzWa5qEgSDeXCs8/atIaMxQpXOW21QFZKSTZsgrtb7gKZvVPG6mI
IdHSQRYJ9pqgIMAe13pb0hZXNXVuaa8D3sodtiXuBr2rbrLDcCN8vhEZueNi1w/E
e6pdrvovtF1DfMQNNWyqQdbyj0wFSHJCVuMO2sf/n0ROyH9W8zJYih9fDpuCUYvc
ZYL5+4EWI1eHc3SeHuO4xWTB8keDXCU7Bpfp7LFGVQEkTY7v3h0k83m3wH0OEsPv
6v/JdnztdRzzPsUuPmp9HUuRk2oHEArBdkDHGEqCzYAlT5NA5thvx/PPw2c/AfJq
VsMTt51gO02KzGyZ+81u7j9RqsP/z7xogW3q2u1XkxzPPdnw/eAyLSrqs7u90/Bx
JoKTRZdG+gMD+GCx4i0X24jiHn9O/BnsHEbVCBgEoryhc3g6LnMFg/ij6uUXiMAS
7PPdvg7BkMGva4K4nYXv6qGibOp+hxfRQgNJGIw1GNhnAlI0yvKNrAzxqkbwzEuQ
8QN29GJCJoYFQ8wb6m6rvFHoT8OAGY0KavwnM4eiKycADRqt9RVYDiAAvJMCov/M
IwBgeRMqK5T2eEdwcGFtqAASfI0zWvHynitW76BcW5JG5dFFRHE6h/ZDYzVo0Nqx
ecY9UHRRKoIT8P2H1Cq1tfhd25hM+b7OVln89fvPVvC4Sn+0XyLLoOwEaiK4Mv6D
Fm5AybUOiF+/L99gio891ey8djPqyaUmVUxdWjQNaK9yGWMqvfkuEeSW1GBaSJVq
6vryI4cFEJcC2yUmgc0LJZSGveZqMd/VF8RbRXEGl2Gy3wKe5K1SAprtrGtQwfJX
E3gLSeXexwsV29F8Zk3ejWlDdX3w1Kya06RGpkvE+8YBfl0QVlGyZYCICNN4E8dZ
3uj+oyMxnyxEz1j+UVo4JihUpu1lqTS4SCjaxiQHU8zlL/OT3Bz5qLG08TRYqi80
bAZNwK5xXqs4E//Pqi7IFnkb7bIoqb/ysy4Y+oVMv4thEhd8MzrCM9hgD6pNjMN+
Mmi7iOhpomD+Fh+HvgkKR9b9lEQVGrpCE8VDfbawONZawIXKi0Dfij9PyAy5x4cD
YeZ9kkpTpAhRWWW1P7YF4Eokyd1J4Iu6GjMq0qSHFvhMnkTTacw1NAikjcQxE6Bd
V7B95MlNrbTOk+Dtne1wRxULTCPF0Zs+j1FcEn9DMdQeksstgSv8IjF7LueXWr1u
YNoRIm8EqS3XZe7VmxfxPxqVDH3XFxdfq3eev2773u/+N0hcWFoTptS+eLzDobrQ
M5j2A4oOWph/RhyxmguQ0HEEgX/U03LHs4pn3m+SyimZMty38UoNzxvVxh9jVVOj
y48DvGlUezC8KAf6zt5f2EsmWLpRPWRW2scnRam942HD/cukaXFzTrWKkRgM0J77
iupDNX9s234xhxKkcULVo4E1sp3NACJ7p25jjoQylV1EnqQRbMKcUakWQrUOKqMF
g9yC1an8DYuAVC4W4A9v/STTX+nZ3r4V6B4PuJfYjnL/ZiXtfxYTcAYlYs9L45d5
O1bTYRoDAJjNLFC+y7yGD22pmE/NYTIkoyk1X4O9nW+50r550JdNQAkM9totv8Sw
6SKAadvOgMkmzGBpZgw/Tzx9T/pPrOoXzJMFgg60uGZq4b7zEfaVsTFLq/0l3jBK
Ps9HyCLVKgyc2lVPks86tzRc9oF7Z7nz/zkjTEzs0LHeZYA6Lg8CNMz7NMJbSH/y
CAj2UltZ7Ey/DbobBizIAVt7Zbm+JvMCavRw84L+/kDcNStwfsbWGU1fGs6pHS15
Pwv+fkfq6kBDuaV9ce0IFV3LY0nIVeNE+v7FS0IEMrxvNzfjzJKhGYPjhXnF66+x
11EAbT3JxEJFncUCu2rZJF08+DN8N6/65RYaTLVLO+JU42SZw4BiWiAs1XBMwMaU
2YE+1ugymQT4GaIEFdTAzwBZGDwDzVFIXM6Yij2/a34mOWovsTXkGX+B7SogiNvG
e5pCgI16n6/xV4SNhxx+NF4NctekBXFcoFCgRQmVmXWyiecTHb+AngIOmN/zXR+E
3TSdlvDbZpPTF+Wb9IKHDecHuCx1aF/GkCYc/zvan6wKginMBCZmXHDC+qoVlv7j
GZKDHHds9vu74v1dFzVVpgfDfuonreRWHRk/C22Af554uek/LPV38bdF3jiAEpHw
f484FYjjU31cdyE82bkZFrqLz9f3ty2XpTHE/C3Qzk/Iqw8F/wtkBCYP15ukueVm
cp0/qbT3W3t9zuc+9x5vylJKkJuyiq9GiTUcW09rbSWaHr7cXSsVjsri5xZBrgWk
xqOtZt5gYoENLkip2iBopbeopjN3fWw2lVkeShhrf/Hdpsm3ce5oeuufcPVsVTdq
oh+snErJFhyf2KSIsXAwq7eC6+cJeim4Ha5DZ7JbP4G4vWnDZQi57urVRnEt+90J
C6IA/gNWQXyiDJ8wlUWSv2pdVv1D8zHNTX97XXi/leTkxRTtu9oL4uQ8aGp2c892
03A9Fbs04hnQE/lRL+gsEQ5b9exbrjDb5lGXy/LZALWbghNYWdxpn/yZ0da08SSU
aY0oLlGhlRWPxYArYyIguFR6P6i+9WkaNRH7kXsM9AoUhRd8vdQEmA5Ss18xNS6o
xKtFwtCoirOxG2lnLWNzjsD0kP+K+CCQnvSnGTwzPZZtj8z48wGfONT5cjtQLg58
5wbhKjMSLl21FNNiHSgwoMp75xx9PgrFlibUZFEyPUVVMMGxktcRRKzfSHFQ0/xD
QlP1yNAiUGB6MYITQYgkZOnkDBVQkA802PB2zEfeYzPqV9wwFsxHF1IMV4Qth5sf
9UFsrX4/4CRj2zY2UHPX7gVNCUC6K+bENIOhV+LbaiiNnYIBnzzzm/JThs0vwnKJ
VXqXSTI20gZBHihRqo0/ZMTnFrUiNtLjzFH4vw/dIZD+3+lBslwFqT7PfuAL26jS
+tt3kv2PjuKtDTVD92yDpkvDgXAm5/QEyGz4QmVMiD1e33WrU5u74R1aGs3orUeh
mg8PCXee/U2CZWgnC4WpOESFfblPBMM4cAkd6zlItjFR0LzFlFk4XqUij5gLE0W4
wH+0lw2sKVVuyrXWON0H7q7CijabE2Vv1QMbQRco4b1o8ZRolP6iGXEdOqreBDoW
wf953QmhetuM/AA8cWYe27Bp+d8b8QwicUAxMqfzEzeBfeyOMf8G+5Jg5Q9zlOqX
9pJzXXMItgHDKZ6u0JG1ZJktBDA9+V0hc0VCups56knGAA0fHB/+ugmUbVwbqp1+
sv8CCIzKVjb4IjW0WcMCUUoXYX+OdCs+JncLZWfu5iCq1L7Pez95GnyUZ1ql7/Pn
2Tflfu5rQHgSldXwBBxco/359b6JE+GMUxAjJewr3XJNZtzT0wXuFBfqXaDT1rHO
0arpekHYr/IeVY4f6omsDlniNaNfKaMoqk4Ead9JT+GWCw/9+OMZvVOZ5OMj6I+L
JBv3oChtp2qFSew/JSQPFeHsUpKhg0OYMsjt/Zj5XrSpwP2zNldKiDjgXBmmL87y
8qQo/kYLneEGElfHHRa0rxhJSeBy0HlvXCO+5wDLySD36+oUup4Fcvh4y0LBydsA
H+Ve1NmSCBv/qlSLMM7ugn8YylK7cXB/COTwI9nBXrMkZwEUlq753jiRhJCWOH9d
5rBqTOl6eQys3tmtCEyJHmEjyNLx7C3ow3U6HCVrPx3XgoDaYw78rJxm4W9AZj28
b1WXcRLwlA/eZqKVaHXe88qCTWP/WZ0hTORvsjqI+B3bv4a1sQrxnvFc5VblBdoU
y/YaputAei8paJpS3AzKqkTG81mph/bHw5Lk1enuHvU5aPWjoEDi09Px310d+vfc
FezHqpjhpxcJOyE4qSsGaQVXvsE0c0t5uROLbPOT71gijUJLfAQ2Ju8eyIfWtA0y
zcnlgiKqfr4z5BY3GM93XMa1hFegciYlLt8rw21WDmkhovb6r5MWTW5EufPq0D/B
ZbDP0IkFP2hzFVaFn1ecO0Fu9Um3FwKRrNwPLhd6BiHQgOVi8Pv2Toch4pDFP6wG
bo+VxeIKqBZvzjJWa0yBPCumWHpJm82TCjAlHASzY6u1cMLH/JIdMNgJYFVBeX1Z
mIm84X30JLKudDDc/jALqr4ivSa8klo85iFR3zKxYJa3muN01CZGmKdTYEd0bD3j
8PBqkP/S7CEBdGUtiQaHtRDpVH/BMt9UOjsXsF4ZJ+DA+LQmqUIvr5+rDLU4H7rj
Twj98elCHJRdRDqLg3sXi82aktNJMarPJD/5qhXSzFAp81d9eaKfh+agavpjXCeT
JtxHDkUxV4wPGWWz0aoTweU1ijSFkRqlM2saBREQdmosVzOJEtCvsX1Z0zsgUF7d
8dFDTz9EtxiGhXT6UFiYsE4sC9YX/gCZVhNCXWx70hwkOGxK9hFTnkGqy2AbG1a+
+WA4RQEH0fO/j7TonkvIb1Z58lGZXen6fH5BajSRsvXLo8hqahO5HgBQkd57gKlr
dfwojT3zd4zToNMXZXaif7aJtQHVbQpM/lwI40yQoAUKpWEZ8WipjJdd8G67AbIQ
+WykG9LAfpDxaSHE0fIcVs+i3D7L7ayoUv8kJHjjCUin7j9JWmOon2YZ5xN7tpFC
B5io+0KNdHbk/+vzrC3kYXtdztO2dBYPz8dswYcPVNU52gJH9Iy5a5u5bzvnfXL+
B8NN+yt2rNLQxc9C+flIGxcc8Dotam3tsYgKFOTg48GQHbTSgI89w6Mz/9uyp5as
AcqvXRgGHnQ9fjd0YeuIUu28CmJaumRt/j3nuYsS0M71BSAcgVxPI+Pgo2LlVj4G
SF/lQNAEz8ln485ujBBJTcPM/+g8lazQ9yS5EMSvQIdnNLza3SiHIbxDc7bk9rwz
IiN+Cr8e0XsAvikpWpivctAiVMtUxRqRLa/ulDaFYmB/05xtbJoNsqqmBmQ1sM0D
60J6I2+fj5MK+tZJJkpEA/wpw82/762nMePbWY4uyMDL7Zd8sWconunzaDcj01n2
b2eikHQXzgHm7Xn0j3+msACUWX6gwy8Fw5DyzuFL0rSnfUsM6f1Gnl4ZXuggmliL
B/OTD7A0nODiH9LFTBK7+YZ4mjuUT//f2j+ilUgEi21Ld1/+KiKrwTRBOowgOpqS
QBx4DOYshH9Ji3KqApdEXKGNNg8dW9UrCq3xZ5BEIPUlH9tSAgWW+BsotOXsne49
Pn/4yingZD/XsPvf/YmKZae7Vm+CpsQxQp3IRzFFB9Bn6cO3S5n23FRcjUuGvz3y
RySIvp1QKqIgDonbTvmaEUQXEfjQ+x0kAfw+KqdFlKOBvfsfc8XZiTmIFaeV2WLM
Paudn9CZ4g5RuDZkRmhPSnf660EMUJYKC1n1xLi/sCMEm0dMwlkwh7mZCb/OfHNx
FfM4vd5HhZ/yQyghZmA4hVKcv3DF8B+EeCps3DPNRDcAXM+5T0WZ4klKr7K0SqmA
GWigPEb0vmnnDfsigXwrn+l39fH4t6Ooo3zoW9l+g6CIpm8s+hFYHnxATmEpbaE6
yxnrWsFVvzGol8nE8zNkjzCNJekavwbsGjR6pvr+9DrigL0t4Q44Mj8ytRgOB0ze
2bMSThLavk2b4nV1AJgGSKyJYL9qvZ8X9dzi20PotcS2vM/A79re+CsNnsi2yjve
BcHn/zlEWtRzGHG0l+Xm6akrzGPq3GHbawJJ9TKzm6guB6OxEPKMKYCoXSZMqyz9
l0nrwUvCZigpQg2rfh685wOfhC8o+oc07uyhOuTuV+B1W7jDNfNbVqR4Pw6cnhLx
4Oot9WNHd2h6zmj+VuNqO60cFhFW3gENYqhXAQVld7WBY8T79JMENF9xPvfKIwZU
i4u7mGxWtNzC/TuqXinBU7dFY4kFImI5y6GUb4Luaq3eYWNB8iEtnQIFcqRXXt9u
idZBhEB1DiBj93717Kev1FCk6l1QI/oTul5UibUSTtgRJhQNMnio26LfbjzSiBf9
1DDk6+0iL7zxwbc1eX9VqZlqsW/fSxR/xS6LTL0TTGIORyd+06HmH6+lqYHRjMNw
AhUvpdJIKGXdDrvGysRj/NnbyVxAOorb/hmLF9Y3A9/FyxAhbwU8L8uh0Vz0eJfa
h0wiwZ0JACK5vrdYQ4jXtHIf1UFQ0D3He3CntabcTb81K5est22AwJoAIJW6n+GZ
25dOFU+/PLHN+K0z04HjOfs7SV5UX5UZ4w2+mwjXmRy9KKgpHqe70rMsZJbYhIg+
cWf1IaMt7UyDpBRA+h5Vyjz2pbI3UBNbwXq1o2VXq1vi9mrj5C9JybjGblb0uPg+
vPs9vCl9XL9VmNzCBQgtRJxqdBF0a0819v0zznT1CGNqdtwFYV7jkzFyDLDmLfYg
Hqz3iq6dFlU4ZHuGiZzOb2zZfJ+Q8w7dYNEV/P/0Ee53smuFrzNOtcltjfPAb6Iw
df7c8MNis4Ptkf9q61hsawx6hnxaV8PSbKmkktW5XChEgbxp+NNlZxHbRjEfGGid
5mRmnGPQm12n8QjHL2uC+q02eGXcdRWmFqpBFBvaTiPLX++3uUm5Wmz1JK0uy/La
nCuPhIZ+7JXg0FtCG7IZ2/uykD7yeMg0Xl+lSGn62XD4R/qVoaZiZrN/bUULcbAb
QCLVVEp39FlkGWOhCdBauaT/M8cms6ecBB74ySTgo5ivAYtevXdKGSQqk6K6f0Gr
88rReuQs4T/GByvRKbniUw9CWxQVNLVfm2tfV98kU7xdZrvoJiuN+jTzAc6Xjdhd
jft9GX1mRsPADsJrXqGShDJuOXXcH9L30NmlSYuEMeXTvRHut8Hr1QzTPsz/TXc1
4HYTA7PK3ciF2TXW3xH5hsOvsrIjmw29N0k6WN0m6N9TZdAL1YUUOafX6YmPH0xn
dvG2llJYxw1ofswrpNcLwGjUDIakqLyNnarnN2NB4PP/l5txT7+YnFtcONSD461t
J+JZYSdXV76ET7fiZwfIwzfFzZ0ERcva53UIEOc+oS1UzuwQmV/ltYwb5pcZD04T
zMKYHowVqxjzwfTshYSTY/9v4QS/58AmjgXmJYLLYYLpAhrKsUfqEkngjJJoPCJT
zk0UJtGg8HxKUYM1izhGf53Vh2i1Gk2Q+v/pDg6xwHThRD2eSjtQa3cc52R/YH6F
chY5qk0fRxmkdbSjVv8bZS0utwgkHWHaFh83HNiRkJEJwV6JwjxXCEWfCc8caeHN
99fbOPRTfV/lNcSj9h8StngL4ZZW+r1nKDlEUWPecQccaVgBA2zVTHU5UFVofXm9
UocD/SCJ+cWQKA4LHgqaXiidGHX3/+Hr41J8c3Ns3fZMsyuc1gBhsWKOGj5WPEL2
0KvgK1kdno5ldSecW1AA2FRaCXHU82uYmPuOsX3pIOvyJ9OWZ/9n1TMCyvRjSejA
K/tgtToc0bvvOSWcxXPJ1lxEyExGnFlSL9esK/RpMdhUO2cE8Ov4ST+ASPyzxTNT
uxFuT819PONOu+yrEcxnSDvaywDSREJd8zW5rKV4tekl6AXI2jL6ZtZE39q95bxX
BBW0/A6gy4WzGis9OYhB3JiwAbjFHKrTtd3NPtSxQ3ZDkfi26SG7dfJbPyzxX/ue
RYf68KqBJabkARo+vFlEb1dIKFiN5b64zC9L7kQ0aXyHF7mW1/ia72XfA1L2OYgS
uIldqUgavfsV5XwE3QQFLiBaVRVERVDgV+zmXduk1Pzj8Zqcrw7hyO7ydAJwY0hK
DTHZatHcKzh1r7mlty9wAufAmI7avCJ9RgIoQDszC4FDM3cgdVLfP/kfcWAw4vS4
CFdEMPB6MhLPmwCZHB93ut+WNiK78jOx7eA/lu9LNrnauBgJOZRzGtBVmhGqua7e
/eG2TdLwrSSONoOPGrNkShwfSvKP5V0vORR+isrOdt5bm+LjejT6xd5ROW38XReA
sILAL88NBiMT18qT6FtDfU0XhR9e18+u14VhWRhq7+cvp7p9YLH3epoz0VZrUshN
TrfunOhGQdFQNEpFCRYrEEOp0hksQcO/EY/N9ZlS8c78yTgniMNaQiJF8eoy4syR
y0VPOvflzZ4Ap0STwpjWosWvPSDxBTxEtbZ6g/lLUepF7rk4ca1B9tNPsubBR+eG
YrG1fJDvjDPSA0n5t9e43kYyycVI6/5nOXwqv0L3D09cSg3dGySnRADj9ugRLhrm
4O3eRczt/GLZ0ED0jcaDBrDhMzrhSehgAMpUlXwH8RuSSJOOKg/8kflmsREkvxaS
ApoOXA2RevcQ1+fJV9u/XqwYq9u8PmsU8ziC0eWkC72exTyEMZ3sr/mMXYlatVQC
VoTXwopkyOzs2MS+DGXje9roGjwZ6285i5woWSvZTTSgX0N/pEZrd71yXbeNfvxg
3tDcJfyfSLjFiHIEiOirFCXKFZa2ui9cBF+zSs0VSCWFZ1oyAYiIhiUzFLkAzNy5
rKzcLvLRc1jN8CsT3OUU7DrOBeIFdIrvwDxLD/UIGH1vPTg9QZM7P/eoOhXcUdG4
B/X+1LwEJ02P2J26R5QSEIgQHmBCEym6UinNBwh3kF1VQ+iHgbBKiTy2zBITS4ek
AcApeoO2Pg6x5neJJg5LTq9Cmc6wwQGLYYNeCXCAB0Xc39pY7Phsuc0kkITtnNzU
fDXlW45yFiKyrnlwGFBj+MRk/3aeD0Hx/wpdedEwD2SwAnQr2b2grI3VNd2ZkyHo
4f76cgdhlMDdVYjeI2+kTEYLqf26bDBOrmXZshiQUZz7MiLSVf9kNebKCBumAKju
VnHf8CNdK2ztKRb/UzkZR54GhJw29e95H6+5kKFoF7UZBnl3dRU84fOkUJQIfZdu
Nq3XPUXlN5eEmV0SuiTtvcjQ3UUiZrVtKyoLKVLBaH8t8CcMcIKVriUTaYPDEqF9
Y5HhAOAKm0RjZP/VA0cPwKH6INeAwTZUOYHtQdsWVcI+iUlrh8xEqXxppGVLIXu7
XjdaVC/hWr6LVSzcCLfmtxEECNAvY2zaQNzH5VkvKeYRjaGR36oVOPJ2yFSX4Gvv
sBT8SOMAM5K7jpmIg9yPqgm8qunPdupu6H9YIy4Nkkc1/bKurkEs1IhNGr1ZGHYG
953i0Ya5o4X3T+YfrqL1ZNevcszAbe9NDDFPtri1Y6ZlQ68QYsFGPS5OSzyUwp+W
RVFni1gv1KiY1Cu/MXIjvXctAeVp9UGazGb7MT6W1XqFkg/0F+z7UzeXkmSD0CiM
Ao61tTX7Ulrfl/sbqRlCwdYme6u4rDBsZvc4N6tjNp6CRyCtf4W5bDB9U4D7m0bE
6n5oKZZuVRBb5LFyhJ7bzZWXxgATop3m1sIgIBSBcv6n1USmP2T83rp8Y4LGpLgv
pKuNoJzM7abINpZisHEo+7KAXAMIsZGWJLaIvFd+9/gZi4Ng7xkCS+UMVZTMd1iJ
pRZvvI+pSCyXpw83ep60uK0Jkaf/DYPWbbXqiY93y6TbK5k9KJrzNa/8BbDAe1pA
wWa4JJm2NJNTMOvOslbVgfTxa4Bar5EdNEpdfedn8JCJnkNQaHNwmLy1AtwcRTgk
iJX0Kbv+3WkXpfsyUK2aWnvbKS7uVgphqI/jERA+xMRtpvjX1krSOm1MofCmK3Cc
s+OFAtfAkvP9LaULPpRsrhbq2gU9+rfLs50M722iTAYKalOCqfIHtAxENifY/2pE
j4rllohwMIrO7r2NbqkSZtRqqAtySJ1PTW9Ic+PO+5xrKlTSTcwj0l61Q1EH0I5k
vFhXGRVb0gmWFO/NvXOApiHBv8OnnhVA0NVMM82K3dU4Eefd4xooszK5TYlyKOBg
jWWGDe3T4sPma/bHg0dlO5h579WyyKEZPifd9YTffrajlMMAEPztKWKUTKqd2Aik
OmcwJy+pR07McVgIonDK2FNe+BZ2qG3eKxXfXNyUIedd4MkElxvSk4iAtS4SR9iC
sbyHVILs+egTlTj89wIP1Yk5bNPaKW4H39TFwyK/GLrv38g8MeS1mlKS7j0COgF3
z4iNQNdDHZ6WSrLflsJJfHDoojFS1FV54m9QW33mVZMgrVVh/USw2dMCWusI+AiO
XdWp869gua+liJDvNEXLTaoNQgYnF8ax3DjnFONWDIY7y1m8TiDMaixuWzgVfyhA
d0saM+o/qhBCa6zQStwI0p1xMVserZrjE246d+rU3m2LwidN3nEYdqTYLB6sU0Ob
VJcPjTn/Po51WJWPaETFxmtZv64zLLNqOFUIGvzdAF1UWB6hjF/IdOSkWPTHU+49
0ftzd5OVwcQUkwyOXSdsMzkyx+6HDNqlFFS7NGai93OEPnKMpXedAUTURxg4LmK9
idrWUi0zmDNKNumA8a9zgwP+EKoP717WkUw3Yp6oVRZyBo1Rr/jk54e2C44WyY/B
xyOpWSf+cjeB4NXyGEym8gO87dt99ejM4l8RNRh1+BCYsTaMC3C3h5j0Q0zKnrcc
auv5aTMcjtVPThBthGG+qB1w8THE7yWbaakHEx5d+6Lr2e5978m4UCeKihxcttGA
T5ayF3eeR68bKL0fC6o7uJC5mIrHlRLyuAR/KD2mC45XOwzik/khijBp7U81FggE
t2Jdfz6oMDE6HnScW0gbLfR4fweDPo0h8VPk5tR0OowY155WXRs6dhChPQpxskPD
ygwNCPPupaYSMYHsCJPz/vRmCNMjN0ZmvNL9FyajtqaISzSA0XAjmFD2iIGHnxtp
vCUIjRJKrx18/iROlj+XC5dLa2j9ZmRV6CcEY+S6h0n1xellJLkWCbEovrkXKvt/
OtwE3AoTu+RNJLI8wH4UcZul5nraG+iPIJc7g/c1pi4zZCmDC49KMJcqzZPx6+Kr
yzBQAOPqKToH6lefQaadOF3MgarJht/QN9sAZd4+CiNQe2UjkATxiSsBeTPvuckA
Bp5GmjTgvBTTTuDBx9kbiNuK5sl/084pNfzIstCWeM+gJj6QXivklRpY8R2J3MNk
EhVO1arZM6IoBHbTf9SsxXuCrltZspVmMnBHvk71ldmbbpnjG/yMVaFjOUPbCYYT
L/O5ddrJc1NoWEf2k7ZJkejtlTmY48bXQ2sQngmwexN67ibdaoN6FrbSvz76nisk
XZL+zoUqHvstIaDU8E/znXZHRtwBcOrzb1aLmjUIx0+u2mkO0SkA58PctNsmpNSy
ik4X5Sob6j6wVtj/TD2PadzJIZac8VrRVv0c5j1Se2K96YgTVLgOQWVbWANZ1jbv
DNpJwIlbQCamBUz2VFEo0LT2d2z3K0tn2OWcImCiZ1VOj44gJKMX0jWZaKoYR3HI
KSLx3y8pjNqiFYG6HgA3I7LIG/e8y3fg73VWsL9tLdchk9hIyG99POIlyKB5TcFg
0U3H+NU/WqRClDquzz+fyfwrmv46RbakP+bSlDq7n8DxPW8SXCTrlFoQB7qY++Rm
/0vuvy/q8ETQhcdI++jZVBaS++K60Nx/+mKagtL0ivJWtZ9F5kNBQ+rp30WevLvk
umdzLyYrqX7o6DfR2NE78av0e9iQGINCRJlnhjPWocGTPUmc6IgTL9Y6TGxhBYdu
0VphvTVZ7bhUsb68qNprFEGkNPX7lvdHGXNKfAOExx7H7DIJCyYDtG62w9vdeO4D
bsM3pLOPIftiU9LAUpfKxbQAKqj9Ii6riUbhycnzB5BP8A5TX9Q9WudG0ESP7jYb
Jnp2r7SG4ZTN+Z72pg/qrPqLyPzOp9jYsKkq/qYZHRzf/keaDzzlO1KIvOcuFlM8
+nvAfAXfz7Gwb5Q8M/n9kCB8+W/HC0LraAT7diO7jrmmflXXarqIr4VauaMbsWyy
O2aUqC2h6BN0JCr/d4AvRlPEO25U5uM5NOdsD33ScPC9RosRshDD8CIy2mn2BdaB
6W2kCetkMwIHUngGaoYXXWzObB1JPnLFyQL9KoBdE+b90OUQ5/lKmu+nJVuWAJSo
oJQBx5wXqKFaAeY0515HsLtGea+Ts9ikyvOyXtaQGwDw2ymgv/mgPEg5xFjWmGJ5
aDRf8Wd0IfnQqrzUQDL0dxsr/M7APS6IQvJ5tcYyy3O5evEwlQM+O1WQH8FWaZ1E
XN1uRT+akoG1zCWTer9p8e87k9y1lGdIPktczp/1AHRuKBvG/4fggRzmRK+2sHJM
VZ6z8sczLJZR7W3ybFqIdVUyzfg19wNfIb3QsW9VV2JeC9zqVMk2qoh/sq3ndm3N
4IdrTiuXPf91HNLFTqLoFXoPrn6BBwlf9jpWfKWYuCi4JJQLTLwGVFtwJMOuO2Pw
VcIY8+vxaGx6c10eQpNPUx69Dr0j1zxlok4/FXcfbbInZcGG2HzTegJdEE5sEylR
z9YW75YecivxzeAFozHdVBay38emouiABCYMpeHpbgtHuLZWBgeUiaM/h7Op9Zj1
30xiZJdnSOWl9MbDA8R5XRekg6aEguj3CVEdHMcuwKpiJOxQqFjqFTx/sl/eMrud
alNuxrWeGYPmv9LzsHlmWSerZyNP9ZIms7BbtYWM2Ipm/XXWncHtVadkpcXGJ0Mu
X35fSiJ6UXZQ6H7SaLNm86Q1PB4d9agZ1zRIQCNTfF9WPbRwUIqVM+r5/+7hMqIx
texMyVzVxt3adytY2QK6BusLWEGjWbMyDycFfO4Q4IEqORM1w0xjAIb7Fm8UAMRz
fwuCNc0SScD66WgDJwPOTACvGTOJsBZJPxv2LL76J0SRmdCyGIgCKuB6AOm2i3iZ
6Zqn/fGSGhA4h0m/6eeZOeSkFWkmdpTfPVAKDYgPKybVyQWuFeKxrjJ6EbGIsq69
Oarhp4QFWTUJqGWz95csmEnRCcrP2XHaonQPpqq8V80FQToNsWYnb1+tLYYHuxDL
71ixLlQjDoSH50ccQzygDl6KdRxaxtRzhO7p2C2e76hlD6tFhz7Kn0oEcxvcJze9
XKtoo0GPv7gzdQyN1mkgtF+E4jjgkxs8tFEu6A3JjdNPWgMnvhIJebB+Ur91C18j
VhdKJPzbXIWHWqCT95e09BnRxXZmtvp5SMCwSssF8+CSthf6Ft8ph0yZ7QHvm9rV
mIBL6Smic4p5aioe+YCUKZ2Ap3uZtxuHGxlg/OSo8F1VJnx6MLYBabhqvoyP+7jm
yGctwtMlOnsr3J68XM8ysmhDS4014z2BKbsCg5SEvpNUhGLQVLhD5bcCYF8qdQBT
Di0OZW94SB78GCzYcp9vBBkciW7lZEsRS+9lqdoQd6yciH78L+nK+0lRmzyAA0tx
FCs+vkcLVC54E/C3wUbAFHC0vQ5dukJqOhFXmC3zWsw4dGhBQE/3f0f8QT/Z9LaE
gTI7lbHxGLDYtfdl7wC8GC/7jVc5wDdnj1LYt4qTmnOiICSa/TVb1/lNp5g90AD+
dO2cUk6BJbrf8oIN5iJbSHUUXLcdVA06wK23sSbF0LA0PsfIEBdrOPbP1qs+t72A
ob3HXV3YhoVCiQzuvIgDpRWGj55mvpmJ4phnGOFS17LH3Hlw7OiQd5mIiB28cUHT
GTKL0xxgHkqJ7lfa8SfhytTE6be/wc7g5EFkMr3GHtRJ+thWenKZJJTQY2qkZHiW
26DDKbpsfo2CI5YpMCdg0wLznVeVoJwNWcp0q4NN1NrvFjapmg6PmYUMVHY6lp5Z
Xwe4XLPxNHccZZ7sFVasaEvumMLHWYM4DVsZkot/AVGR1RFwQxCXKjTGMYJAD/iU
YkGJBQWISVhdBj/gJOvkyw1eyCBmWUOoZy4Xyu4yb2xjFnJ4/n4VqL3yLRPcfi11
B0oM3vba7FWwzlijPTTJw8xeA63BipQCkTX1EjFUggDKNkC0ZQbT/JfDNtjDcNa/
stm69oe5qeHZmOscGa3mllz6QepmDMWwM/HilsO3uKIhb08ApIs+bmOwEJvCpT/c
xZ+kj74Vr1aCIUQUKbyXqqMbiTGy5/A/hhH/WqHP6HvRvOOKL56QtrrkxW4ZPWzl
6SkV/InpLzx5AYA7IgWK+VgfvYwhOB9jRx5WU7jpO1UM+iXJJOVzPall9FDYftg4
E5C2lOg6N7lIIVfBN85FCxTGo8ZWpax/cW1CovrCIfYQGdspL6I2bJNMNW3uvL8C
GTPzKDt65cnBp/pek5LuR0KFQ9qilLLpB5jYjBrMe+dzaC4urV2RMAty/IU0E3s0
ayNobbOijTvgVXyBHx4+CUuC1Z+T68NoH4QOjK+lEfWPPu/ny2IBIggvy2ErADbV
9HUeW81BZ75Komom+4QqifbaBLe0qGbmY9ULTy1oVnhVoePf8ExE2KBmsdLfO14J
BmUg4VZ7BezCjJ6F0pNC8rSyMfJjO2nsPSneHbG8vLz8vU43u016OnK1Wxkf3yqW
61GXwbP21BV2RSacRIRVc+Iay72PTa5/nHTDs9kqvEZ14b8PgvoIkkr2hXDRGALk
rsO/TQkaDOYNIcRHtSMfV6/9zMMvmVP3VyGVuRiO/PC7T6wQScWLZHsqC2DittD7
QMLfdJHcLbABmNSQoC5as34ekp60j10jaQQOAa9MLHGxAZCxav4wmS4NLp+3YJ5Y
un1M3GtJE5mGT0sXnlfkj/sqfo7JZwNQDmVvqchjyXItQ9/2SxCBibOtRM4OsbQT
ogbIkkmBiNjVmtFCldJl+Wlt0eAHq9Ceeb9E61N+erxY/CLRa2MoS6dPfAT4/nSu
dVDfdef8jaqrN1VYsV7TIK+3N12IG+MyV9mV0Rk+eIesROrJDNDit90AuHWld8F+
1uRDR7EIzRo2pYE/jhZivaClxVPKhhU0b8NZgS7FPO9rkjLB5wMnNBZLRaS71T00
BX3rpqzGPXnbzox9uE4W5h5/2SpIt7VNcIEFzE9YbnEmnLGQVE2QJRYkzB+noa1i
u9aKWevRqnFp5o4aEnco7QFApba2iI6uVwD1TYhmUNk128rtD8RTDq04Z4rVH4ti
EoKtvdbc+x50jdfg1Qoix/T1v6Gm0iE+qOmunELwpQYsGIFodDDgVcvE6Vd/fBfp
bIXDDdO+IiNFcYCl9lcb1cZPbfT53cMHjtH/pVkzYpzNOVvSV69CYEYCX/Z46CFx
EgY1v+PG0Lew4YCK51vJJbsSv9+lqNG3AGT/FdxIzs+46tIPjCXpmDEf2XfGwmQ9
Dhl9eOpVQSqKgBUueityT+bLYxGFMC8cnvJoyMJfdxJefp4eo2/qx6JDiMb21FGB
+Q8F1l2b8iG/5WhLmfaniDKcPjSTebEj01XcYtXy45d5HkQbJTFslssU9Fyi8bjZ
gwVFgzhmJ/s8jqQejoap6GA55nHk8zQeQ7E7HWp4QtpEAdKT28s4GSX03VAOKg44
njzmkHVCZUjV/RacCg3AmtP1WCqtdjTJzTbwGi9YppWQIW3+nyd6V4Sagdko/Drw
NkcZaryMMH51ouZX3tmsSWEX+nhNYkyvGqrVFr9AqyTFkNr2A/J9izOrM7GsVntJ
wwH3kgs/r4FYAhbkW9piZhdLdooKMNsVFDoUItvsJCxv+QnVciMEBGHaoNKCC6XO
iOHP1dUuCUBCQcfe6XY7khuInhybgF4uaO8FgedGGAb3ztkhd73jy/ZUTc0/ljaS
NVK+JcFojdnyqPfz3z0Aw7UqA3WaNp3oAY0qPYSC/uxV5t+lVDrvCYBOz887vquG
bgExN4pwVlXUMnEwDCvYmV91TErV0qCAowg3jY75JRETCnlLgNe56cdGiHGjkJ5f
ygZBPjgjBTqO41fFYb47Gvi8UJ4Ax8mZLSBYa8b8o2IxJdW4FwXwnadxwmRHYQee
urg/Kh5mhQgvK5triV0s6Vdt6HCCmNJ/HQs/LMETogy3xsI3SRlU7SQt7sbn+OvV
hv0BEdpO432Py1DfoAOGfWrE8M7PC1sPHSi3yl5spa059DOmYiq6Nt+eHkEEA68B
+DOcRCtQ+QOvJTA7KUvE/1BafPLxB++jish4EbAolXB5e+odCMVdAAm0/MK84DSm
jlyRTXBgChcbdNrmZYXBpZ0Ly4GOowC0qOl2PkBvIV1PlOP0IPn2rAQ3AmW0eOQE
gJykmdTp2bB/XnTKuDrROFY2Ftmhl95bv3s80wz90u0kmAOdHQHMy7vKf87Kyowi
GyeS866HBrR2yJK/KDcDQNjUzdb4XhNYoxM9ODtQ98J6zHZtiSywVvrFEg9FwhWI
1/1TuUJy/bOqWGGPBjtW8A8E9ulnhl5bDQxRMvUhowr6HhqukeqCaR88HMxVH7cH
TgYYyhds1AiX9EEaDwihV0fRlgl7Xh6/Z3UnDqgDNvkijslW6UocOzzRp4ZAMaTO
ZYkMPBgETFs6tuWuyJFDsP6E5oK4g8qtwRnmr/dZt3VL3y+sl8tQ0mDvYDdAJM1W
50bKECARzOR1niVzykJOEL2rGarW7geb4EhOMcZq/a7ZfddjS3RsOvlsYFQ6E4BL
vp2kziHB4xnxoEnQ6N+Ab+2YyuC3X5rQzcC8a4iV6cMQ8A2V6RJ5UAm++O1MaQQz
1lc31pMNTG9055mQoF8YLIu3yBUh8CjY+L3guGEleHkLCohWgxj8gIItMCUougKx
onWcnvxochGkXhDg/0JGc+6Xvgam48CUkviNRIxoSU8412D409Knxfpp11wxzgPl
cI6k0dbdmP7axVzIWUqq+HnCU26iF0ST0lc0r/pvZMC4+40TqKfcYJhcTvNRKMJV
1/6gl6tJ6gCNSgqHGzLrTQZqHhe1hucB9KQ0c28NfTPg4B/e00HZjjj5c4dtoVI0
Dq7rL4+kujQDxdP0Mor6e/iluTYpPExVX+i3jFIcgIvr4xQBmqUfP2rUB1gR3zjK
/9BmVlcaFzZYxor3xHQR3KBxsRSW5nPNWInhKFBUldn0twDwuMQFY3xDXm0+L2nk
nH5nYJEWLetpGp8RSQ9hLS7i/caZoiAszxo3W6k5/j7KiKnz4pDr11ZZ5XMxtQz2
WBTu6SVD5x9mktngnLawC5kBKHUHdRfqWCyuFmUZDO0dK7uDrG5vWBfD7fJH2knp
OZYDNCZhZZ7Fq1IOs9T9ruOvH7xwbfdxgXN2f2/o72Wv4fvykcs8J1fNK4WvPTkw
MT49rkIji23fOyzf9AYVCSeCgJJ/418IsibJaj7kGLwHuSqpFA9CAX5wiVCuOWla
6FSzqEQon62nrM3dn9zPLdaUyIaHZyiR8Pu12Lz3izQ34YB6Z1rJEYRZTqJPgaJG
zwLw4GoSnwZz3pBtt4oTseM591WR1VnRbAE2p33wcUHiZBqRAUzFOJEd0OFI7wpV
Fq93VDGIJlDPi4rWk9n4r/sYIWS/fwfwbXOTxjsKyjmzzMRMdHHNZMuwmnzbwQ2Q
XxX+yCZZGFN1IQGmFnfEQHoPXFlN+ubldBuXZw3iy3V06IvOU3sLrdK0lt8ZEQ9A
xtmijLe1/Nz9kx03QYvmaMJ6QcYWJmFKGAVDrKSsoYBOSiycCIhbdY9dgIHDgC4S
xUkVCGlg8xthfmDkX4c3J+M4Scb3sdoQPryGbDdSSsQ/ksIYMSuX4fJk+kAs2Upp
AwKZDIw5nsEm+deXjYzQPuVzZk5an9X1NZeAt73+fmRicY8q7SHZjF/G/bzKMNsy
bzMjED9EMzb9RYrQ2aqcwWort6yXDlEDSCKfTmkTyjG06i0WDvuo00vQrYmRPSG8
rJHTq9bF5MsTgLX4YKBXJyb1DyOeWJwmAQJ80bv1npcOoXgTpmGbsKi5EviFp4Yn
0IIL+ye3bSm3t+i0P5+c4HJIjxv6zVcYnfhpQAy89yl5GTlmKnUkVDXd8iEENO6r
7fb/hNm4CVXpbiZp7h+so2gY5IHu6pLvHbfM/dMnmA2c6/BVq8KqiUelOcinSs/9
TkeSYsteheYXC9bK51HaxroX8OQfsGgEmbLUo3TJDFmQF29lLAvY7z3ujdlvnu/N
sRJl9Sfql2jt0q2HvUnZo4+cYzqBRClN5BGDUWJfqHMJTZnzK5dm2B7MrII93U+g
z++abBvTYghEapEGntLgMy1Lywg4+nl4UokkLHQLMcMSJ0FLLq/BrN88MomHSrce
xKhIQgxAEKRGXQHRDxUoSRylR+uxaToCrk43otopYP4BGxJbUOu97SOO3CTbmoa2
nFMxSay82pztbgYaJx3hp0rnWFZYmssUJl0CM+PnMOjX252WAipSfSMycmFx6RsN
PddltyFZS6QsM/siLg3O4WV8FyA+bcBGB3+w8o5luHWcA9NKNoWqMLnXMxTo3ETM
YivgFChl/vMHlCC2amihsujK5NDLwC0M4G69zDlBdOqNhaZS7ZO6bHejLygfI3F/
D/XvJ84JC2phvs7SPMzKV94YoQlduHnvOW5cxcUOJcVZAIte5VMNCDHuJ0I0JLpp
+g7ccFL7bNJ7D44f26ZA/ZMx+cYytXI7B6TtHLRNaLDUUCejXtteuZWfSC8oztI0
mgldppZfdbLwj+Cnb55OU5Tpv/XGFsAQGvNDC08Q87yIm5m5bFW+iD/v472CI07l
wBggQK+4W2+Nq9wMkCzNF8nx02Uk8fNL+Cu7qnS8RdAn5J2tNtoMwDxrvQ2E0//B
dex6iL5BYeHTTV5sAHKHoH1Eqc/xTgcVYUCvSsVvzMUKOn7CEmbyXujVAkzOthbR
EZchx/VgKMe1IcZNwPHK7KKiKt//aEZbvXLO1Bqd+QQbunfylzzQv1DlfDqQDMcj
xcYZVBjE5LxGH7Y8nup/faCvh8TuT2nQN1rxQ5MBDsI83OodckbFKat1t4zxBw5f
C0YhSQz3VRHsuZg+W4ry1nKA0vjCxJZSBN6ACet056kuLDKdZSgIt5yR276K7gDs
QC1fVAGvKhFC+MR6yhHxyhMB5MGSogWCNzBZUsrxo8K7IeOI6xbpfo/xsyNgFu/k
uHzAVlzfC+uXMJNekpMf9bZYE2x3cxFA/FiO7dD4zPTuConNhVid6zkweXitqYYA
BBnZorZ3kMlDrXb8S6uy3bSI5tbFCxj7VNLXORofnukOwDkC7kao9k1lUHSfiuPM
Tcrbxj6CPazMFmSGoKZVGfxkCGM/OZM1o5BVVZt08OQOtq3O8NhNbUb7ePJZViRA
GfenuBgGRaICmwsO9nwxCKon+7ai5QDSZE/eNVXMkBIjaE5f6rqsMaYiCjoPBiCh
r36BWOhE5BdBJPhwxA4s1vJEU6+NNNm1N/fQGpFahD+yv8Yvj1GV/7DLns0ouc8L
DzqpZlwkAF1SYRVk5F4hj0mQHHNXNEVfP8fqth8JW/8RdKcB3oy5PohEj2mbH2Sf
/j0a2Pk+mBg9tyeXXV+jOcJD3SqpAmzFNoP68mbpCash4514B1U/bHEhQlh1f7n3
TOadn5SDBtFTtD5TWaQ1/0rIkWZRzCcfatlz0RQZQG0j17e5UIs22cfFKel0GZzq
QDfc+NaKchLVJSiP2XTNOXN+6PWarW/xljmXQ+Kp65Dy7CDQ0Dt2PJ1RQUkTszvZ
popaSR1N1BRjq7xkhoJ9H4tvy5HD1ZiIBn/3n7dMBpBb2I2EPFZ67CnEmsu9JNVo
z7AklSPfpX6uT9ttB2beoGPirJlXRL1RvIeXA0DCXk0BW1m1X8e7bg8IRBx75UkU
/1ctF/aK/TpPgabpqLyrMlAsR1oc3yFXehZZoGrikUWAKQWf9PIX+r/hbDM74wD3
Tljc/l19S3Hyec8wz0Nq895a1XKdmeKMDM8Mfc8Mro2Bsg1+rgd87O2P9JP7Id3R
DF1MGgfPlyAOYJiKbTipPFx8J6UnmpCFUVlAMZK55/YmIsJyEpirYRLVVefKPxyi
fTenlTHKhzHp8LytgmJ9ILKzVfhwXyxpYS09DD0wZ9VELN2zexNL/wsgJRHv287s
2BMTAZHbX3H1V3hLklzU6uOrHsi/CjUrZW3DBtxLoqn9Vixo8R530h3bU+4+eICO
quVElQAm/Ef0FSiKoCOr/GDyxZYtIqyfl6DQNsoWYhdBDkeGLXv+/kNHM2kOm9LH
DAiDm8KG0iqNn2juc8ryRxnVIJ/Xm4wNOeobURFyqhwvJt3/IqLyGS//tQ61hL7o
H1Qbu25m47ghLqu/xr++5CjLoNHEQumFlaDkXsyq4azIV0f1Qs0UNmFbR9U/jj8m
wZQxxgQBKkvljJLUbpQkkJhFQGBO060wSyNlS5R+AFxrzvgkWJQbSL6g8TWYR61r
L3kbSbwtVSIMyCe+9tcoWxQhRtF+qKYnc07BwnjUjr7TCehw2YA7uTmDgdXTCB4l
PcnT7o8X6HlI8fIMvlrGzSNklLVjNhhmSlayrkBKgAb0WeS58/MIqF9R9AJFOtaz
3ElVqxdrvqb9ShOslTBOGPWSqJlvrVTI6GLRj7CRuPolkhRCG6CMCvBIFCctVKDa
yBtW9aLOB7r63IgCGHUGGLR6sqbzTAxPy8nKwCyy7Lt2Qepzu0d6vvCEdknm0pcB
kYQwv0Cc3xZyNLa4WQan8OMVQeGEHw8lCWPUcMRxlqHWhfh2j7Ht2hY8uflyVAux
kJRdW5/zOF5vqjZZqytij6A6Xk3OjZST/fxMaeGFUK94cmzAknacgZp5ysPYI/j2
wqeWyQkqDLpUtQGgoy21BvxI6SrxQcxj8nsGm7Pvn9um3XdZ6XTjUTpmPlvjcS+W
sz9K3AEPmPhC4i5Wf6WBn7Crm5Q8rU9ZzZXCQcnNThBR50FE3q3puv/bFqqn/rgp
o6IvDAYahFBUt0GXT8eAjNFB/HXxF4lqR7Isqs6ztdp5qyloO7/Jt4y4tS8UA+/l
klESJuWb8NYf3hH+f2v/fS17iUcNnz2SS5/+65EeHaXOwzQ3epr0+7QSgDHOwhhh
oO8L3oq6vdfWHu1PRhiWWoV1XgZEblaVtFwyBzo1rrJ91KuKVXNRROwBxKOKyAgN
Mi6K3tZPn8/PBtObwZI455k0B7uIBZh5FyLntx4XJZEVL5TyISrvkuolOr54UMbI
UBxqMHOBJrqktFTwR2GwRnsIwKUcS/WrtgLz5EKzmpaTEZAtzXUz809A6lo6OhdS
aYDSTBKs1YCqwDrJRJAQJKH2agSrR/yU+gx3PHnHGj3KcRrA2wEAO/HomlfeNB/x
ZIWR5mD9bQ6KMJbHCTpXfXJfqgpNuo1p933aldzAVxeP7dn3pSH83ZmNTzSbJM1h
HBEL+17rjqFNjQhTRs/6VIj8tJcPl8ntaLzCYeTu2d0fvSUaSrH+kXYThL+tK+GA
+w2yTs9EF1Ti3YJD/P1BjSnzZcdynQnEt49PVcYqz2dFi9SGHlLemZQWKgjj+Nge
XzSgR/pv8l8XI5Io8QgVg5H62Nv4rTxxaTi/81YyS4FD/lx3DMaOl+Y2KyvHW7+8
vPKeVTVUtEtChcWwPtJGawDuStZ6jhcqdeDa+AlDyZC/YLesFuICGaesQNr75hxd
27fT25l9vaCL4sDu2LV7iV85g6Lfl41B7B8EO10yjSfT8iGMnIMUV8t2PeW4xkSf
C5QCz1MXydbTOgSZ0J1orq4tKzUPK9RBxoiaFcP0d6MwFs58H7D03kcLOYay6r7v
QteIfaOs75Tz/gUmmhU6OPCxVkHoyJg0skE1V3TlPwfViMcXEs/x2c8f0pIFyTyM
DddQP2CJmkyuzOHW5gJ83r8eBMBi35rpbSr+qvyrKOl10O7PXlgzLBtTkf+j0Lx0
SRVlBAzm1X+Z4Ns/J4wYdoePbK7JPotRtLHRIrC8CQDNMiFQ/Tbu5WTGzrLw6fX7
E135o6mqdaO/9XiEt8kW4Pjq6+N9sZvD0xsHqWZZRSnv9SG0razBou/+/mMtwAnr
UKrs4LJFhHuysw+pmI24BezSIGw5434KrpthTO13vLf7PjA8bNXQwCmiOerLTeFF
FMP5clqJHjunou6hMnyI/qDZkefZ6Uft8iW1KUCmFbD/kwQBf8IBIRc37ODESOT1
LyCL1MDDUdpk8uJ6gK2xkjbLvgAnNSIMhgmlMK1vkdpTw1ufxs4Mkd9uT0adNdNI
KeX99iV7/rA+x+R+lcqqLWdBKMJj+0lvrO46uDodruZ0XWiIqypejg3tp6fzV1SL
bLX+sJ+PZPQU1CZ3h5vdXye2FW6at/YnB0oD//VyQokSxBbBS/DhYP/Wt/wB2Bqo
AQOke5PuE/tsVb6KLLkdTx91fRYjkghfUpMsyLYT4wzZz7mCsP0gHE+laHK0r+XB
XJLXaReK1WuXiUXJ+xSSUK5yxBJZFMA8lrXfTJY15dyWBsus3N6LBJaLo7OOknOX
XNBqTPpq87mSIKX1RG0XimnmNA3tr46EwvocEQmpwSCwGjbuPul86aoWkxaQO0Bo
+cqbm0/7/4k0Dfil5Ucty6fBgmXbaWRFL+A7hdcH2b6XPb6wvzQA7Y6LWCqsQMiJ
8TwDXFh7ZYhxXK6A7h9Rr3gdcQhgp5ka0sEZcBP73pPRan2IRWRGaxzjw7xcLID4
JlPo4D6B1TQ3Y7xgTi8KEgfGY134Kxyp6PLznNzig0iMH7rX3cuLl+t9pjAI89LP
qayD2p1xohajJfSL8BTTyF6wxNy9wVkg+PV+2RLVDb4BEn11ay7+rJCg7mFRw1/9
J84aa9texhI1+Zm6NkeVhIyJH9LLdPiT0jRKCVw7SzI9zkfrOYxbkG/6LIUYI9D1
ujIfJvECnbx8n78RnMHQKy2wj2oTsOWMFlI+vpmHK/Q/pGgPz6WGW2arrFDCCmj8
Yp6yM0DXXJ09Hs6LAlCRuGXkE6t5HLmyC84KlD+ALnGSGoZpJ5BhF60zjtcKdpD+
gN6zyjQBJFfLwAMkIfKDvnr+h2KMkw2QpruX6Zfcdo8dQTipT2feARmir8cxHMxc
JPMihtUIHX5WAoefNWPlP6HrWGurxBp0JhhNctCQ7Wuw5SXKVrjsOhJbDIdaqQ7e
U04eWufvLMcVZnSGGuuppQgE0+mB06zl279+uWY3kpTjuR5EjMLYPxTu2aInklNI
3MdGF5cdSKitvyKmBJ2vfZDMvxpY2fF4Fs1T4ybuhaJJrTl3iUWe9p4rx2WFAHEF
E9/p1b02E2SPth6JmNovSQcVOrY0WTDVoWNIwpdRFkeRLsinK9ZEJ4xEAu9DGOZw
w5JH+N0njGEgCaA2vvRT0G4NsWkVcXmGS2Pin7FuEPaHRzeB9I8JSuF0dMmjegPm
A+ttKYMmdPPGabZqbESGmw/IIGagRKzrfmB4Z88x2ZdM0bAOpIlMYIUs6HFFATcw
nV3jSaO/s4kFpX3wnjAfyM94CiJOIlyhyeMEvx+rnkbprXvI85HJ5tvlYXl0QZuX
j2NuZnCpQ5pE4xuA6Y9YHhSDnVtiy08CSQBAi671Y6jV+yI9R9KwqwQ6Alf0Bo7o
PAZEvCQDogqPVxbiBkmZ2QfVhL06bBDNXNgD2Kvcojg/00yaPrKfoNBYygCI1D60
3CjpfcNhG4BJrwTL7bKydaD3TcxGgoT0J6HPJXgBEmrFIqZOx0DiSRo5wjgnfd2t
4hkWR9YrlcqsrDe9m0eXCvCBr7M14kf6uWePPPtM3OVJknuhvAhz/T61+XZjDxV6
4L+qekboqCLJIYM6uf2TwielCDZfTH/Ij3oZw9f/SqBeq9nWbjL6HaNY/+1oplIv
25PLZLywaD5gEZcYTFkQ6nqbxbayZGgr/RWUhU7XCGFPt8p5Xdpj1gz138Rc48gc
1niRaWATd6YXDT4Tfrijj/9IbEA5RDh82+TB+cyq57BCVmDajH3Ogj2fG+xgA9BX
sbK7H6KJ5veDfZhibPVtKwZvSf17RRDKRwoLKfKrNWipyy0E7PULyKWbVj5wmfSp
pQ8JJB6EAfCRlpKDqVyeNi45knJLvVngUC8IgGcCFlAfpCQh9OscrnN8drDM0MLg
hLrMy7mrz7+QnE9RrC/HWko5Q/ER7lvZb6POAy+y2BHCJfTBRbtj9990vxZAf1Tf
0ggqvdz+V7xgX29qIF6OlcmJVxJ3B5URvLqLm87EROdX7DXntxpQSI7z+RHx4oyv
l3vt7aRFivCwbDAmgWVuFB6vNTyngGuy26kYOmCKdFBeCAdX+9wSK6vVNr4fCNZg
IN0fO1Mz4DxPcDQX3Tcw7IZcxXTk7VpMnBraP5W291HfzGB41su5T1dRwG4vu85c
ue4yJe3n0dqHpWK67/jZfrTIflizDLfOVzHTqQKxhkvR55qbHT6culyij55lxR2k
rvY89EDnjvuL+2VvaQf5254JP30BvNP7papiDJY2QbPbLfKs2MSDRTCsBrnm2+Xy
g8FAXawOVp9EsjR7lpTSCEO7ggexYO/W/CsHWm4/RS8DG0NvMMB1xQOeT8AvniQu
NCtl9+Xw/Gu+YB0/eS0SgMNE1dnbMp+u3bFpYPY3l8d1kMunTzqjBrXHNV6Nuvq7
Kc6ceAapku5f1nDU+smw2g7IMH3VMSfLUt5sc1W8/iDOMyCmQtZz//W7b+ZqkjZG
uhpvNwEMSaYRxyYc9AgcvyUJdXMAaUtOFzJi+BWecZUD+Ltbej/cNYksVG694L7i
SmiddbPU865RaiUFcLoyGklGJrdV/onHsO8JZBwvi/YfNVhC7IIjHG75h/YLviYW
J4tu/B1l/ltn/awYQUyTVoR5ERmmrvS4Zzbp+yAxhR9TBuWXewzTDlMRuI22SVmw
O7XHvZuc52zqt2cHlYU48OWuyhc1jZTN/3KsoZGLPLoWCEoPd/ssTdV6L5suqn1P
KQCnpiRUFPggyapVptVEBmrLdEIddrd5ACuIbXiF0JQUXdRl+0kv9+vaBpWfNEQ/
BWXkPxYrWDJ9nQGaX/EkjysEcPE56KCQKdlguxwRGTaTzWoDOfVcVaZg4s78vHcE
bowQ1QKLsLXeoWOOfh9b5nplulPOl5nrjENR0L1AsG04ReyzWOv93yhV6DztVNm9
WiwItBKTMyvH8I8gzAMYe+Mp8T6iiA8CQlPlEdm6p6MxcOjxC0OqR7BioMSptUqW
Ko5og16kaDqohzVGBntLKOOMrrBP5eopXowm12TmwvQL5kUNo15TuRL/kB00t1/5
wSjGFh1DE3gEhDWqRhSvRvi07L1JzeooArDhTi9DRHFRY472xSPnHusln26mLWyA
X3xoul/EpaYXSH9DEwjU6du6w8bbodVjadAXCb3wtBx6ooIhO2h4Iphpx8mzPKbB
OzfM1QyqCjjRV61da8FpOX7/gUOB7Dm2GbGJgzc+eJFKlcLjupUGVYGjh2zOFeIB
yDpkunBY/3ugI1+X/vkfw+Vlva/ttRqCRQN6iEx9e9VRydGV07BcjB/sg0Apk6v1
0heZ5lKGmJXKQ2Q15cWR6dwI80ib+R6WLdagopISCRcQV1lhxFHRHS4vgv5r59Ym
E23a8Kvf2c/fdVJhm6A1I8IxuQHEYCyyK/7p7tVjqRAxFqOqjWmTCWuCMam5Nrx9
yiNpKNcRhdj6Yi5kNfhuE6mJiEN84HKOoVrP9pEn7Fd9lg7dsVjV/H8QixWkGkZP
+tyrf8ZfgcZJoFDovq7t+eGyHlXxLhJgezKP/IzkJdACrSceEJgHYmJFu7kdK7ao
+PIyCwKF9grz+ppvKRhllSMuXHt6kEkVPv+ikXNN1kbP+2enxD67aZoi4yYcjnL/
yUHuPk2Bp5Hh7TMnOpjCUP72UHg3ZKm9hzaZGXDm2DXZKKacUBhCwX8I6Ub46eYn
QTS/DIAyxxg2kn4FydA6gYahK0YZemCBEC2Pkxd7SQXtUsacarcS6oY6hzrRXW95
zjTq0dCGyJrRrdAs5QQbXBvCBx05WZkrmxzWkNMhFBxZgn5/RVMIbIoTF8Hs7StH
cqtethD8vtCYua2/8/UMYRcDtsm6PBLxs9RQSkihpTc65YrshAdOLxk0L3iOmu+I
oAW2E6ZLdPydayF4FJhZ6J+mI5CRHUxVIQpR8ZHnQ9yCQ55gP7JAmAl1QVM5k58W
HltrQl/teLH7ACjGhwvfV2Tkywc5cA2Aq7hC4oSYxjU0TvJU3EoIEIKtvVMTjiZR
mvkfPmUMl/l60wJHJsXLgghaV5XlMHwxtdbZT0XZCguTD9gifXSASDrHqTwL1kPU
M3rPbPaEllVwApvJeaplo4Va4/e7be4mY9v+7A8Hj3kWn/bDWTQjqsbPnk2r5TMD
pdv9tCBqgF0o6l/yAaJRtyfVTfk/YAHkuj0oixT3VntMGWCBVdnEA+x3J/snfqEo
z4AayVfyz9WBS2P7gD4iqtIvT1RciIHdazhGxJ+mXI8tpofLr3caF1mdHgsiBzvh
vY8yd+rbnt9mTOTJv9ZSaf+5m5+yvVUBPNGBQamuG1FuNwWOj/s9B9Nf43oHYusN
g7v0l00Zo2gglczbO/A5ncXJi9olRr6A8NFIfKrhEUsXZxM+mdPrbECQCx6ghSMM
hQY4gyb9gxMnjr2HtEPxXgsjnSpV3Z9oIFMDvLUNLmMOm1rGg5l6t8PjCUd7ykQD
9Xf3mWczvUSOA0goOsZqpATUGUag3oAlY7kq4sc+zC159MxWjecxZkSjzHybX2eq
fELmO+3flpk9iLvTKEx5Wad6DhMe1Jd94B/8iQcZB9v9JoE1fmZ9XW43OWYeKClD
1SF6ah/khHxacMmxqmJqtfV12/nuKCDQ9vt62KPho2l3zJSG5cOWy7bB/nlZIp1i
u+JYYrcV2fVEKoSjrtElAUFTGhXG2Ga+yqaPsC1XKPc8Xs7UFOW1DmaUrgj1JAT1
hvcYFov4uczyoAXrc0q4UGendb05cDyFc2pbPj2JYFMwQf3OutJjGYGTRxnfgEBq
waIoz5C5J0oh1ABq9M5sapcVX+RnIQX/wlY4d6+wmZsq48GyifZg1Y0s+6dn4b+Q
DgXoDpOY0GGM97snDmyVDtI5T424pQKojm2xxEyaGQdUo9Q+/vXdtWW/08kBc6R4
wM6XS9whq/TBbhu++9FMhihKuY47MKmJmm7tnaVJGiBwlv10l3tj9dxKvz46mZlk
SVajsu+aaHa2fT/79VTORNROYdZG4F9E/Ree61v0VxuISAmjA5/T8RcSaA9BjYmf
DKKkojKNf9kaND8OIsuNUN2xmg37gV3k+jcp1jauplhMWOYfe6qZC3D8lpdRXP+u
2vEUBGLH5PRDbmx5jFkQqGijkUqY6Jv8TBIpyiCathxWa/89kJFTCz4QuT7dE6K9
5+AEOFY9fSq+OKVX5rZWwJEbY9utWsBES2ppMQLdD5OcZvwpapVq6WDsyNxIVDnQ
quqhrpmBF7gtjqV8pFvNKOc5jp33fljuqDia/SJqFG3GAaL5mOps5mE2viv27mJI
YmqRoiMhrIkAq8cJD7QIwEgWy6jRwohSp/OSbOwrLDYChW1GPCq3zfHqOTiDsiIb
5INSpJxIZaH+6R1NjI9/fO/ho1n7BPr8WGR+vrEdLkqDcLuokWqXsxZHheLRFxBl
IA4v3/J5AkdafncecNQNwI8WAQ0JW1QfMYCkuvZwR/oLQMU1MszPMN8aZWXgWjeG
8cK/GGKscVCJ+yTDEc4zdzyhn48etTBIEEi5KiOGU0RxCX0ftwKRFYEkGobo2th0
SmBDrfopH1ks1S4A+ontBun9sHxqbhslKi3zaGtl+3G0K7vL2eeZ6uUwVYBaEWui
xgqNJuTQlS/B+LKNODklqigLXm6c1ZM+1Pu5XyE6BheSkboP6r6vZ5GPIm+I57cq
onUQ7ewMiiQK4Xhr8asF95sYw+Mo7Q3ayGt5q1x1vWWPXlzV+HIcfippGI2SfIrd
QZhj/zZxXZWbJuciWcfjrpZMoK7bIX2RV8r8bVVKC22L7E1jBayz1EewJxdCW3Dl
RAh2BT+ePNCc+IE4+YegbqqCEaLsIq1lzkojy1MSAolMA3mxFwWpcpMPHd9J+vfe
D6WNmV3Ikc1oGLy6dHI9awetQafSKsfYCfxRPtuU1/a7s9r/ojnJwiewRhOjrz3z
Mggc3WvFeDNcUSwPyXzdjneT/ulg4V/GDuKycaAbn6FkNvwEMcOyi7yFeAkKmyEh
j8ihFkbpMJwGyzOeCI4PMj8hmyOO76TiEfd+Xk1JVfCzs3RK6jTovlit971dqmW7
NKgPJgeq2tao0w7bRH+XfoegUTVFvPOOYoD88V/D7SU9XsA0RtPSNcpCwUTNK7z8
avXAq/cbiwFtokMdA7GYDxoHNtBWKVjAkMKW+f8PDSvh0FqQjaHJ20qca+xCImCH
BKCoq2r5MnMsCthLSYmp9wMDeECkdrPQwJi3VfvDqNTHIWc56dO8XZsEOvmO9kdg
bovQUH4QNMzmpLSXu7+bVPplYrALM0grc2qIuksCFQGotnrIEhZMajJihERToRvB
lSX3Bh8ftV3SZDaFUD42+0FpnxHB+NZ+ASL59YzE/m8DLWlR7SHyzdsHFeXeHjlQ
xxCUFGEJArW/t22uwj9Nszq9H8u6EOhmwNe7HlOa7oALms8K6zVjjbwO2nyknEVU
148o9MzH+DmbfGUTq9/QLeaU2ipMOVsgLTE5HemOth1rCfkWv0Jb7UjGFPnhwJ/e
inDu78o++tECj1+eBB7dFUPxii+nGt7z65DUVwlwodB2vim5IJt37fwgdCgwT7aG
r8YPMJ3YITraJFap8ekhUJrmmj63dvnkjI5rrVtP57Tbg9RyWDjUmhyjKV+eR8ju
JZZpun2g+6t72ISv2yYYHwE7rQWXusTd9a1xWMPuYc84ZSiO5D67p4unTsgjgAQr
e5HRFfvzrEwJbmA9z0ZmmcpIAbLzs369IntEywRKFCnguNEgIJLmvnjTmKey3khs
yaMtPHdjoAyZyCQm9utsuFdHRA3mkGZ0YJ4echodXTCRCNO5nFm3APl8t3YVhaNd
oIQJQX2gRAdynMQErp6Uk0gWtzzC7oYc2E1F5Kz94/hKPaSBEplTEsBaKgTHE5Rr
eJ1G1RbpBANodrrm3asgUGNmlvF3e0OV8/MD3R6mVjfNar+PtgMzGAfmOlDfM0zo
OL4Jk3tkgdze8MV85UswFkhYep5lWNlpjxjf3isrBRph3t+EURQ2a1nCtN+OcTLR
ceDXaHoK6ShIWRYFfB6QCVvjP7bmccCCF7XHky/xu1D9udikS9YHlKDJK6EEDiM3
QxtCsevL/kKjBHpcUEI/UnMHqtLuDpKGzXAdZ9ZgI4/dgJgnBJlq9yjHanNjNSno
rWdKveEbfT/swnWagoGrHHBovbcLNx5CMqyM/8fQoogd7kpsOnKujeM1Xq22x5ct
wq02BITPb43HxRECa/iIQPU+dsQ8Eho0jMGCmNg9e7C2nwJ9swBNVxOO5P9ZP/94
KITlpG30l+YDPrerQmlxOnaW7lJro3ofGcX2Gxa8I5XfWv8GEOYhvr2FliMyEfyK
LmNDswrTcebcYWb1ubqQGiAwFZegIg/DSy84Ty4Huix0FhGFcvdYHh9+BovvLvQW
mNtZMZM3B9gbeHecGlWV6+1qkcNAtprrP8jExjUb2CqfamFAtMkER8R2d1XmIie0
qEfSVQlwGr3HRICGRHn+tiWuunF2cCxyGYZwCZ+bCmC6u5RTHblDTAkubKY3Pekb
msj6vl3GdU6a3Cjd7qd2MO9TzLClMS2eKasl7p2E0tjOQwfc8fEJOHme4orxC2Ly
c2bGgNYAPzVqJMLMB1lm49bFU2gsspImz0bqqYfxtYyNBwgMO+H+AaYDW8P59XRg
EGSSs/wnafCVmWdTYs3MbNPXf2NoqfUVKAPpu+wDsrVic8N+na/ZtxsCFDYcxRcX
MFBMgpZdNs89FxoMPRx3NYlf2c68x5YiFhUAZH5exxM2DmNtDOpV6EEI/cIaskjM
HkO+T5iIE0c8qjLdmvTRyiR+IuPBLoOGmtp9HEey5VH3Tb4jgwx8shYR/q/Qdu1q
MHXdO99sAvMaocyHvVYx4I9OlmZkjOfcQH8hkx3ruFHfReBqX/ePcurKqyAhbA9Z
A/SGUeqh+FYqiafAmha/4YQ6WRj60FwZBMkcHxcOeAZH4K09NyhSPU6ui/o0HAvb
0MPR+C9J7bFwwfxGDPMP9QBopiRJEUfaizZEUbT2RMktrhwub7F9D+0w2BEXAoiV
/8ebIRYWa2KSDA86+vvoUwbtZLmE5CLBClLX51banWXuMhfhj5yl9nlmtgm+XzRt
bGrATOmepy6Whv1eQaZdxJVyrb7MoF4Tb5C3TOD+AU6OlEB1BhJT1d7BIHtXHWp2
qNKiyBQICWYZvLUAcBE9Vv6pLUfLLxQUwpT+lSX/P3UlDqg8A1UgrWSmquBejE7K
ngJMGVeSJeBzf1+eTdOs218OYSN20sQsj4rl3TtqDfc/T/Bit4pYSv4Ng1hAGaSN
E6YoTGwDJ0pJ8ndp7OfkaBu6Q4AHK3OQlhHuVmG9EEIhSO1UcGywu5G/c6XPJGVG
0w3k7XzMvMiVjluv0FZzhGycbot+BY4CHQANmnnLq5T5gzjEbpVHIb2RVWlY9oKA
EN3NNpX+5+o01QIGWVkLbDneld/SVLUt+QvfN90iBv8l5pQMZz0ilT1UdtMX3DJP
TtTmkmapMvV16wweOHhKexp1uoDX/HItFb9Mwjh/CKrN/CaP2n4TEQ/BFh5eR/qE
pAT/gdw1ymxM7CRqD67mwmFQmmxDLx/uGMI+BHPWxyT5z700DkEFCALQRRH/RMyT
BKpfisldOIYpRaElJKvRFDz1O1uv1HSEhFqLywWbQseOTJT7CPc+2ca5loCMAeg4
/Dh6gTzykUCfkHq0zc61gjuRiUXkileHH9xeC1+YrKFIWq2FSGHG1tuGY6vxQ5lg
oOw7Ct+jfeLaPgLazgEV63AT+g7S2LK1R9lmPjGenT0ul5VbMdaqPs+bDcnmOD5U
xMaWhKeoiKDSEmrqkB6Atbfl6XtZ0ssoYDIM2UKVhe8sNlXflv1Mb+KiufDcj6A3
gwgY0Z9WcFTaerl1LiWdITlGZtuXJ4gSMPYdORyBLRY1d6U1vRD2+E2BET+heiho
uKbpgMNSrV3WD/GBrCbXwP/Qnb4R7QSScyCpcHXkTsOcc68bS9HjoALn+b1RSxZT
Y1SGuYq+On8HSQ0R/W0yd0A7H3VXAFSkU+VGTSJnbxwwUCZyaYFXcIJ5AsfntJ+5
e9pXULGvidjV6pwgQbIKVN6AvJW9EBgxpQ5rYtuxFMqn0AkqlSEeq/o4QDgGotGH
a3U0VZVgumJ+F1KPGzsEl1N6WSmE6OgmUT3JFlX+2ZAanUTqSIY44CDpXXGXJgl0
oRIumvM7Tb3jqKuPSUmcl0u5HsNtlgrSasXR8ZjnKNOaoC/tXeMKwCRj0ANynbsK
aaG4SDAfGvvH8VNoqA0rRVZU3NCRIzREVt9h7FpDunslDJDY++hxyKhCpGWotqLU
MlmgdhXThLXBSZgGlz+r3WkeSrs7MrJFrz4T/bzpdmyPOo2oaMol3r+oK3i+mRKP
HM0cSHMR+wCJxELtLOt49aC9idSlaIDkY7m8FNlW+OmU57/s0IMlSXMi986iiPpK
uFZRdiFMdG9xqqNoi3DLy3NhaUCWn6i5YtrzInCSsZc23puuV41pzFbWDKOCIUfZ
MWo5tpBNWa79vrPGcfkBm2TFihV4CPvbFx+9Wp+i+3WVnsqKuMWxhthsCI9fHfdq
sGtbbBdr5qbECU0mM+RbA3eOtKIuykGx/C8k6EUvSX0d79FLZ6Wozt6kbwtpWUKU
Iwre1Y5JR6WyuiNVgCAFGFycxKuZ/XXRRW9ypXVmAFao9UIlLwWDMlMkpuRk/nZV
LoDVcMl2zoFpeXlVpsMe0f5yqxCft1Res0UfZXJVATFKj3noaurtOpWwmz8IxTdY
yV0pUT7iExtcNWMi8EOKEbx2jVBKZq/3R+GGdG5w91NesUOTQND54A3+8R2TzbW9
6kjAktOmXJja6OUAW5wFLvm0qXVFci6IIdLUHjOT6l5X6BQZvtQB6SR0eAwRQuVb
iSh0d7Un8skeaCu5xFCI9L6JukPeb7dNc45WLX9o443KOEP+BcbcZiBZWyHU0j4S
KhL7gU5DwyR8Ohcd3p2Ncpfgpw8Edfl336mgMgnJrmOrceKlxlyCwlTOI8qTbwz1
500KO3/RS6YDoRc1DHWQvlezh741zKE/CNYWlZxdIMJbNHvay65kzeEG93uWoVOJ
E2JqWCAKFW3ZTAJOvvg70SOtBRv3ESuDDpYmSKxcxwnxWEY0SsQL85HbC9iQVgTm
NC7UGq8srEXVg8KQSvXYK+jWT4NUUcfRjcQzkhd3j9EHnx1T0j6wbQIFu9YX3aCN
OdA1irYOyuIiMEQ3WctNfD0vis/fRNENdIjkDSRp1EjunuGryaLK0AEBWx+LWIAJ
lCYT6yP5iyuvgwymndfO79Uyd2q+AonUy+q67hIovIJyrmv5Md/tJSJqPmi1y8Hp
tzdnV1/gooMrKXfI9yVA01es7jLe5GhuNfThrKqUHxwvXS+OAbUxMLy4FNuNaBI1
IGwNQSZoQBjXOaGl3btcYLLGz7iZ7mGFQWDw2McAVf6wqgEFkLl7VZ2tC9lgr7Ed
+uGjfq98gjMOqHh8Ug68+Ka0YT90krT/Bq1KvLaRXrJW3UcJg68Ip1GjMZjH/C5+
JCsJBHTTZHnLaNWSd1w8GXFrXmbpxFESy03EuJXq92objgFfjtUTV6rk9gDKY8me
aSr+meSV2yNCs/kSJu1PnykmSSkwcjm3DEhoN8dflqHjLE97fWNUkKvWxnjQdEw0
Blt9n4PkX4uHvgfBOEli28oxhSqkDEcPp+zoXv4bVrdkhDXGbWs+nyawHSeGEMI2
dulKOwPTAnSR+pc15nUtkElcDtNVi3XcHttub4gpE9aR7nin4P2rfIk0APyDFVMg
al/5nDjvJaIR7QRpBEXaMyK8SS3qNE4DFIM1u+n4Lsfs0RVmFUggGdTmDC3rl+Pw
LRS/6+V4LdCZhZnVE3Q3ZvBm5qRaULpnYG0zRikWWOrcC3nDZtNso3+POMTgpr6o
qzDWKpXLP9BaabL9YcqtbzWry8UCX6Jpp3pG92XGqCbOGHq7X452mOIk07nnM/UZ
NzEakl69R0plN8OM1BM0X2GxmN1NyFI3M7bmWps04ZYnp000tJVI0o6HattZm6wv
x/2JPySa22Lj6uVa4TIthDNirFe8i7asEM3wx7uMEfyTCu10f9ikA3iGgxUID2Ku
lYS4j99IPjjp64EoJ/Je1hhgLUR+hAPzZwYnHx/b1JPpcO57Tf2689TVou68CK6t
SRY2Wp7JU/X9hHtYc8+ikvZfX+XCc4rJul3mwroRf6qHwzsDoVDkeIhiLTONut0q
1yM8OqMsFFtd4q7QS4lCJTas6tXPTgX30TlM+jeQWdrtYXGzB+0OHgrnApnAg4Zw
vLxmaGVg4GPQ1mUvOhsX0ZIg8k0WhXotvdPUeSCwLqKUOvTBpsUkBKxEV0vmJg3b
luF8tHl2R9RwGO5XgGXny++eOO40NJzM7ZX9zIw9YW1VFonlcfFu8Bjy+i3i3CMk
4ewTK2PjSGCVg148ZLKXcLAFsYaW44w4ea3OgHwOnvAvrrDDYbb+8VNCiAdLtUNz
mP10Xj0adgguRve0pB1r1LU3nx+J5HzZiCada6m/X+g84EUvczpfBTwhhnaSzUFm
ZpHGkoN0w0svsm7GGtgkhfUiB3oFqmItGzLJjze1ZG+tOSMjkCinPKrMXfPPeN4y
7pBW+E6EtEPrwOSfSyvAVb1rtqLaYA6uWKRRgiSEr9KpcpVJOVUZFFKpgc6WqopF
u+cpbugTHJKSZY9CX8FqYbpAL8QtAzk6iIxv3MecYFMeyVHyqqLNE1G1XTSt/g1Q
m/k6HKB1MGSe62sAr+hbRmVzIoDvNoMjdfgZh9yfsPzqoTzxhtveiPU4cZZV1IxZ
MHlfRHnWJkA9NEBSOXkEd2WzxbHRPLhnQNswQaATd1IUX2v5OJCSN4HpoqvHukFE
gpZWMrKRIGiRPhlGpwJLfYvLoGRrmo/mBEVEEaN62VyuEig0/GePgDXaXA7a/pqp
nxtrsPmSqySd1eDMS4a+GsniySJzrLWhIIzpMwLLoyNPTB8grEOOO0vafUsNwdZR
mpyxXwO010Ezyi450qDZmhYe4PPR++aAmfyqXi1i/T9SvzYV23zRCwHVe4udZoG+
0Biv3C9wWIY7m7njqIY17dIWEj6wACGqXRPMHkzF0McNWMeTYMxeYrhi+CUtZ1Hd
7jZV1IulR4dvXrSQGGAzYpBwC/KhB5/8Jrvpfjt5FTuCkzkHcgGtbaw803ux19kp
7dgAsB5FLGpAkarV4/4DUB0+OzYLqzHaKQU2JyoDELDCp5/yPCJAQnEPvlWwUOW3
4sL4QKbEGmiIYLEsj6B4fvDoIGuoP7tdq+1jXz+6pvwP9dL9KOxbWUkbSeYTDYod
2kXv/ojHk972FzIzBpv3hhmSoeQQriLEXr4POKvSp/AnM71VYwLwiTdBqADqQa7o
szCOxWxgex8R50mUzkPyORZR2N/rs2lwWneIixE7SKHfX7ExtOi1Mzj0sBak/vUH
nI5C9UKGeHeKjE5yAao/Pmcmn3tyVONMBgwWdGvu1PzioPdS/WEl7JQ7S/Rcy9zc
9+ALxk4cBov2wH886vCs/8h3ECGUHLimOCxzYfiBzgRMgzKDdGwg/NRLbf/5de9C
wRbxVold8vNWU2OVrRpeAKcv5CxPjziEbzuIE+tRDdzYNFU4756BjGWX2m/l7whA
nWNbuun8S8SMzZ120PQUdAybAVlHqBe779R1Mkx8w6JHdq7YfyiQlTCaLXZcyevi
kLxxV4AkyR7yrzMvRvpMm9LCy/XXLwPbGXZVJ4s3iOPNcxgZLi58h1YZD9y6KgSS
K8sX+u8uJQKlaturJvkg9aZ6wv+nIfYMl3VygnmrzFG9brZ8VvSXvCYwSe1HhZLN
cW1pyx1n4ou+zEmSdgkm7AVPUt9ixuziKMJ7CDNlZXjlT55XXB4NglrboUupeOB8
JWdSzUuSPN9sTLWWxHrkdxT/nT8HhGkykief2+aQdDC9X+9Q5IAxa1jY/IywmDHc
ksBZosPi3tRE3S3uIGANtGZR1b5mk8JiuTaoRNfyvS4WyAoWYGj7U8Qr39RTV5LC
b4fQQ74VErNtXOlvkSgk0622kYyqsKyEqKlj4DLAbizxtKufNwwA3KSr6wEOk8or
yqITv7+TlB+mFCHP7JQAtPrEtaCE01P+pYD5a/HBP8SRZvvcIcBO/LTOrCm7bV1c
jfHZz9dH40+4crkyRs5j2PcFasWGSqgvV5suI1paFrJP2qUnBeSCvU92MU6y+2zT
/kToGbKGJ4DDNYSckLEo6l3asVNWNwE9l4Rbf0KfigBCH9yKLvcOOHujVDNt/xq1
eG5HPdjaBcZ7ZI6+Wbl1coGlAguOY4R3Sz8eSKdvZNA558XDc6XmBcqd5Os5qhFz
ogcCxypleBZuvPqzyO95A5rtvk7+i7unM54/WY292NdxBb5FrDtm6L2KX9IPZGoV
Di7YNpOgDm5z3LN8c0Dup7lNAqAR/JjQSrJ9NhrrTLfh7R0Ycbd1yjZ8XfHKuwmR
8WovOfcoBG4vHzHuGu4IkfixIAkS+0j6CDEzERk2uP5TInbMKBCIYeUi43OZN8Gk
Iu0eu19pjYsyvnQvGcfSDhQpDO9JqH9jFEt6BKB+J4Fq+8XUt0ti7Vp9tkVkKLff
NZweJmHEIqoDdKw5xlLODMRBT6VuuEmHfrEcbrOyJl8Lf9rX0hN7rJ9fi3OX6KKq
TVeaxuviejlEQp0s25P0S6qMdgdnBWrWiZ/rUp1JWqPm8q+zofZnFyhKoeuqnzBm
uWEL135mJ0ErADf5zZRi8RYjWglda6swkRLaoHs/rZFl+rAptv9NPW/pmRIoxzt+
SikOUhztrWyOAtnY7KRJPNy3MuYtzOjqyNnXbXgxDyOzMw7gQSj1mfCkkKnqwZRK
MHG3l83WonQPxMtsDt4aAZV+ATHqkdlz5El43NPbtDZ8lJ0YqZPYb+qa3mMOhPfw
msw9BVRKrioGOGmSiBWUhSWkJFFrf6gvDTPi451BCsM60G7i+zp6uRcI3Gey19c1
fKKvUyDWXG00PI5IRHIxXW0umc+r5kleUbFGP6oSXdw/nqCdk2lMknoSyPjtBRdD
GLJXvExUFbwwAP7J5+jVm235ltdeSkfP8ZEVkJUTBJknCKVBUAjo7Q9cWxCxFcsx
KXyQGE3VykbZY9HzpzTW2++xlGj+ddgSqCmZ4BaMfPzcWNT7ugccfafUrAhsHu0T
S0W2ZtVyndNnL3R0dY23faqiCAAwYoje5krEw/pS/PYARL4MBni+OZweKTmpLARp
EZzmLTDPMuuJR1KupANmJa+WxqIUvl1tQgCDTuYFZNKknLo/tjr5fUltkOFqNl8b
nrEuGGe9jK517Nu/ggNvG5WnoVWo4mDWPcb7ur5baZpL1e2t6Tr1vdTiVL+GeJqc
lJWH2QsbNI9jl9Gu11jp1JrdBsC1OueeyJp0oehL6bHgDQy0m2EXDvfv7r3oBUvV
vf9x2sxgrRStvwZhq18NabTvPvMStM0Q6e+qcgcCHn2FoAc9Tv+1B4FhRBx6gJUu
JQ/fdnAi75dCbr8CgbuFUgBhqtnSJNn0dJjQzqX9ZLUqUuNK6zzsWLobFEHBUK69
rxKR/6M5zCyAnG5Rf9CSs63i8DVvJx3WByeb1c8fN8FPcd9OHUve7xQBGXu6FhH1
pFLKhXdEjbP0f7e614RizkcXFqLTl/j5k+5zzJX93WL50jhIFRUhrhtDZryHmRuj
vjnuxylBUy6MAz/RJ9Dk2FCNND3ZofKF4GstBD8Mp0MlcmWc4q7UZklEwTx+JSsF
CyyQcIwFEZlvhI4r13QEYnWAUU84KQ6we4ufKD4On+cHlBuIEEPeWeBFfkE1Dsk9
blZFXzvsw8O2wyvSOirvKzUGUUtVTfP2XA+Q5jLKvOjz+FIjf9afTfJcft46EtsT
y4I2+pZdtQiZe4fypTycCXMfGEymPfxUOCgPPGIglha8JuK9f4PGb35mltcza68t
fjuvdLTWjVJyfiZ4+D0P+fNMfcJWmnMMJjGACWH7t1HxC+/SWvdW3RnRFtmLPQMU
gg9cfPi2ZyA4VIfFiSmvkH+0O1sGtjLampPMN2jtw9PATfEX/tgBliHrkCKhC07I
TU6peiWA4qSbAMruwzgv/5PGdr23aDecSFCIx0JMf7+NChmxPJJn254QRpKCusDQ
LeyJBANlKXx1HzAkSRE8Hz8xL5r4Tmkem6ZtzTybBfedmiruvb0XhkITp4I/gWcf
dEKlzmCDXOzFBLI4o0OzBTjN4qR0++FRDJQ3QgrzWM9hztaFb+JWXqPHZjNoG9hO
4j8JADbgu5pzxjHYIIMxdhgm+7EV6FXu3aNb5i1OuYzgm7bFxF4WB/6XWVEjVUaJ
cV7i+xZokRXkrv6ir/LjFD5H6zTRVAGBTlrMT70gjQKSHZ8Azfp5xEi1UiFyGE13
VoY0GYYDNA53Zh2FB1vkDCwkakpocp2t+JrGif3vPJnN6K/4CIZwsQoF0NBviVlg
SXkr2IGyx8xukh9thcPcQeKPha3G9qNtWqvblcuOFXVfKbKWk8DQnfs/jRgfz1UA
ALemKV4gChz9bAkaAVmZUvKuFStY6/PfVDhYAHeVF2TDqmyPs+1fhdI6BqUpLHxc
OkrITwr+E0Qz3jyWBx3J4L8oGxT1Kq/S5d0NcBL8BPjvZzgl1im7iOG6av7LEnz7
W8v66u/FQjh4egsUUGhO4l6fh+aX0rYLb+QtCWNeWXdg+EAqmgq+gG8frTLXqsNf
/TCk9WTuqhyCjDGpLPGWmFyR7fmnSg4mzp69zcLiw13m6ykBG5N70NpBwBnwPQRW
7oBqs2B4IOxzeTZNWFXXz1pDvEHexKMNKAoMXtOcVoyUEBXwsuQDRBLtdcQN5xuv
xWzpBo87YSAFHTk6Thciu/I3TLgDaX+mc7VIfIyPd0RIE3RrwhkO/LlKGqoc8oi6
Bndblfteg6vEZg6JGD5SG6KTejA+c7Hplw+sEcK/qGYkDtq+oH6L8q8f2IGtO61r
rB2fugcEYDlOiW7GGclBhxiWFPNPrFhFt/qhRQaeq6dF5qmR1RL5SGpz+S0L04Ae
FkcpMNXWDShpDbE0TyLJFmJomr9ZVngEYvxN1zdTISCH13dYQ9cRsnO69WvLY0dS
1x66mhhazE+ylANW/8f7O/OVn0Kn+AZxAutNcmx4RrQIKgcObwQ4cNPEgr/oWUXL
BVi7T3UyyAk701mB9ek4KHtlbHwHg1uOrGNlchrTsP3CR+Gm+BpmVL1sSw8SYZtR
yNIzPymR2Q2RulFg0Pi5vwId1XlpSQK2QqHR+Wrllhd/HzWvLN/PE5Ei1BzgbAp0
+J2B+lwyHL0rcKHpml/txBD52lpufYNuZt/qlBmwiY8CLsknw95BkbqAW6a/2rPO
UTiXLpMB4npkUM9RQmij4nUlmSDUmj5Rk4E55KOjnopcqztgp5SbLJwmYB6R6hL/
DYoDFm8g/vWCTcV/cHNejmQGoUo66abDF36c7XtlozgM66ii9P7/A5G4SVe3HgNI
NJ36DrxVEbWCXWH1z+Vn6WzEVdrqKjD3OG8rNau3wCCX/PCL0+L6D2EZgEMZrMAr
5NVBjtjjmmI5J0kt+GG7SeD1LfkZjNfN3a7QQkM90MhPs+vSGLyH1XYsz0ri3HLt
Ie5+BYIiw9UaM3Kwc6LUeaDGd8sLIbpyjup2EZ7cTm7x8lW94V6QPeNSyWHcrO0m
bcrhLk7CFNHIC/xq0ScrrNLZxvqoVM7EpxT02ronmpPkkQ5zJvCOLj0L2JMKHQ+n
DetZ61TtJ/w27QqKfs1KNi3eDZ51bnC3NXG9Hgz5cCElhSS9UuCYX+wHBbgA4b7J
oOk4Us2LQ1Sv0aC90n4yAX3X+M19ZkAS6hRY/mY5wSoY73MhOtrq+yUWe0XczdvG
sB3PCrMXpnWEr7NbnU9y5wmelg6kOi1W7E+3xih0ZVXECpm7+333SlH4+gEltBA4
Uu2Q/CXfxlm8ZHDWP8s/ittWJrIpgIpT1AqnnTD8xDsDbLoH9JeK15qnLiV04uvg
dr9QOgxoeTpmUN6rXQwuPrpWfsw86xFBBK+4WxPzIbQofxJrg2p1K0KEUpQ7J8Es
sdwUaQC5NV2MVIEg4IsxKU2Jj3bRdxW+/jChe4HaN0aasO5U3LMU/HCy8u809g6+
yd7z0zymvoK8rqWEiKaJPTtM6+rtvKPpTcKY+uPeAlSy0nAKFRxylGZVzJAqtrfN
Vf0B1T/CplwL6HJ5ZXUUmcri7yN7roJGvmMozqtXr0kml7+W0d6NeubXZboy/fws
bsz3VrWp9UVntDj7EiWLPi/8D/I7jy9r+Ct894MlvwwnqTcTgE532v+8QlvWYcF/
FZgD6D7PCJApM9FvERCbLMeWOg8PxvTz6+4FsHAph51KlXeZl4Qa0pJfJoK2UvuT
INXoR1rHIn0NYHxXKPsvSgr4KX/bgQoqg0v0wZ/l7djo185IqxKDqQprz3a1LFjk
xj7V2pJ36IQ+ETpb0ZYFi0/Vt+Qq4Y1QGH/w6hqZsu54PUXJy36984BWE0nXH+oC
AYiAeR+nlh09UNlmuF3aJk0EXlMMpRg8G2/2TF9r2CQxGDWY6vkngA4yJV+dO7Kw
UMk8tEmWM1nws0ZyFNZ70ArRYfMK/Kv0r/j9hPwCTSQ3EVqP2MWVhskhwA20hxuX
nqd1GZ6IG40VQi4kBEoAXPpYj5qM990ZVFbaplpRIuqp6sWLVsR/iqSG76R/1+zt
iTUS1/Bcip8jjsnFA1qc8xOs/Uon7K07rbJSAQWAr3AX5JZg6DmxgegldVDC0npS
ZgyD9APl7tKbxDkW93Z7heL2LlRNrK4upsTCEGLAJzkXWuG9Csl7X1pQ4xzQjMPJ
56DLIasSIzcco61nl9TzXa5RUUzjJ4W0FeXmoCKZQYJamFAMLcfnIa2VkyfW1xqg
5+ch5bqAf2cc22dyO8LMVXf5+FjbJKz6GvvTLbxyQj4odhpREOtwcC3d9mWm/j5U
gsfgLogWKfLXuQwNriJidxjb+OdvTxxcqwifElXvsqYIBG4rGVQymqgDDGXg0LFL
usVxYTq6DSzpcXRgyo03vpXgRnNbsQykd+E2mhV1Ho7yNCf4ml0el+13XSYDD9ba
WAvpP0X+zyTHu+x5SN19LljnpYaoMtLvrPHTaLwjz9GOThEgxGIZx64eS/1N7PaY
2/WPFhrYQETkEthIyMwvkNa5fC0LDM1gEWETxAgy8l5dbOYiaKMaGNp1ZLIVRWZ6
MBexcFOMAG8ompx/BNXA16jTRj4VdhR06IwfpJivZbykKAhkUmrXXVTloIvlih6W
mmM8Rav6Bfm5Lsm2p0HYvheB4f/dDxv/90mR5s0IdL6PIX46a43uHfQlOtHJ+Gh0
rhhuF6YkIbiZX1rz7MtdMrHHpqR3gA/VbXZ0xrqn1eP7wf9Yf8yVyaUl9AW9dkNE
IQZfZcf8SCTD+zwZeFh8PbBOTFeR8k8wuRPSJPfCDbQXlYEuUgRGN2PnMyLdW01E
FcSPJp9Hm9LHyx92KE5oVqid6lxCvCoVcsBWSgY9yHhOXfNTcgzTSB5uUDI7UDYF
/ld9JpdvZjSRo3O4LBrKpFf4Y5qQsneuhiv3cK4V+D5hmrQn/tI6zxfLEfEBRxZu
2RAMS/RzmbW8kIdH2ReKc9XMN5J03TTgRGTTKFMsNnZCnpFtuk/YUEWLD8kQD3Gc
Ul/behX6ldygaL/tyww5mi62nh4zbp0Ndz2vi1HdJI83w1jU0CCxs5NBv3IuVjA2
3odxK7UWIpm6AQayCwlq8IxTQyOe59I8KZIudLM53v3eiuEii1N5cG7OOLV4znqs
A4iZL9x8JJYiJnkFYZLxw6ypb7izV87sXSk4K6EaLLTPaxJMUI/OmcaF6g/weVJT
S6Szxew4aLylxgmNWtE2p48ZCH+lXByuCAYySpf9NPFBQ8m9BVQzhbm1DdzF6tnh
BdmSiIB4sv+5lsqA0RtK1jHbAcLtYGCH2KPBgStwrqt7YF1KAb6LEwBFDPdaz7S2
k/u8EGcBUuaa0ejk6nITGF2H+lA1sU7j3P1F3Pr8lM6H04JfOevSrLWt/IICZFPz
mj0BMn9RsthXOtsiEH7sTPKPvrowgAUUjqcghQ3RV7mIK4CapLl4TWMHQ3SkbuM/
RPmcuEuO16t0rD+zQlJ1V50QvMvd6ovwSRwxnRNaj5RbxwYrEr8G+yyKE1qhRNIk
1Zmci9c92rLqnid/qrDMn9q5a6CZGJPzt1s3FUZu1yO4AJOIfXdgr3TJrjz01Xb/
xAFGcVsvIwGovmZDJEk2eiVekhNrpIpq0pJqAyIfA7eDa1O9iVCUlXPeWnKt/bXK
yWYdliWclOzCfAKmmTfx4weigLzwds51a495sd2Cc/mDwbAfN4B/q2JIfrLBGmD6
dLvT9hbQTMo+oEiE1+UTKhgv5trI5Bxs7IahiZqkAIdRUWe7hq/J+Iuj+pyngT+N
Hf7H0jT+Dbh8Z5uPrsZ+otNwEPoR2S1ZgQQ6wLYNp7Ody4OfUTlYJ1/l0S6qeSe9
vSV1bRNWlLCuTVXP1+4eCqoIfm/oD9VlzHCfJptDFo2vMOpV8sFrcr/Q+a/XA0Z2
eAwRgRuD5U+OlZMsXeVFOlF0sjTTTmTOeHRRLb1Nkx3x0UEVUVXXpaogtzunN2x5
S2Ye/+JchsHDZHPvT4F76IThsOLfiHlp6PARMSjjNcNUO5ztS6/vAOnA/Jftogwy
zcErMEcJEPhJZUJN3Mxzedi80R4QGw8Y51gdkVhOPV4yc1GwQltlVirXjkUqJ0w7
E5rjHXJ+wr48XJLvNkGEr2bZhUDobuvxWWfogiiGzJQ1r52ihr3zDhyWW+71gGUo
tqGgmlUsX6QTcybKlmwGyrDGHgvRS2MC3wdxUKIbI+NCYGizUf6Ixa3ArzhyW0W+
MgrlcEU3ql2v090lXj9oz/Dk43TVKH3o7nVkZUuvkEYfxrcGQvigNq84AnqahSTN
USilBra94a9IggKbPZubNSHC6aXHxthp0oukSu8CHGUc03XdROK5W5FCyG1Nz9wE
MfLU7nlQtaGfYmHsEOk57gYShU8rMWu46h9ToFthWdN9pHdCBTWwDDvBVFTcRrGz
iSNmuLunlfSBtvExGKIeoYT5ThlEEMEyLHc6t0fT//9byut6tZsDDl5Pmzite75f
nyVv05TL2Mm7FMWuHce8L68zunzCVcCEl3wUQRtmGQkMeZwGLHZkStRjaR53jRJd
nRdrvUVPBSowbAMmrQWdj5roqCDw1iKPGQ1LzvV2WTAiplabnhh2G+Q17KtkJieW
iGARbEGb7QQaOe1srfx6DG2hcy4fUPOC+ZqwfTFc7OahN5HCZLnqRs3v4n7BkiPU
l3tMI5eWHjI5x/i5w00qy7txAz/mIeWPx6XPQHspDN5E33tJe8wbhUnS5U2h+4gj
aF3j0EcdCUg8Cf2SZdUYitFUVrrar7pCctdswJieGsp16iD3+o6q3svYBR37mtZC
5YGchDViYzwFVdyXMhWjHUaeT3QJRgQut7lNu8xq9W65O1bEilksh+lrh5X5kzCh
5w+Xsljgjud+ci4Mqn35jYfFSyZQa7lW3RIEtAmSRdT6MB0gSM1qGp2wWEDQ2EXb
uBCN3Ei3yLZJQ/YxFlruUG4+lnVBtsT4wktB5dCShfXRwFvjS/hhRF3F4sPXKEYV
Q77ay3s4N/XcQJvBfAwQUM7aCjAzldPkG8OOAIm9KH2ker7mUWJA57ZcwbNSrDr0
u0QvvHyzF5IhBlwVo47qmK9HhTdxvaPLfIZbxi0jt09W9OPD5DStZ0sa7akuM46x
DQaLf0IJY+mPIUPEtQnUESLqcFWQ96ndhk1CwNQ9IDTD+UIBaIuu5oxK+s2S25eR
5Fn7Fajy7ohINH7FkH0jwiH6yS3vcea4wstIlW3z/u06QpaCnd3jE4Kb8d4ENBft
lX94OW4FK5UFA8YR3R0doeamSJZ71XDxdTXxtY4aI1fRkaTYmtEiBY2jWHeL6EXL
OMtvmBlAepASoBAn7KE97n2TeGNKR3VFmovW5CVC8sjXD95ZIr0GDcXtvYzo39+T
ziAmmNzJqu8CK+m68HQboE39Xu9IfzVm6CuR07ii9bOCw4cnS1gi4aVPDAd85FFt
lF8sf8OQMLDxy0EO5FDXa/VsA7OnneLE2oyj5Bt91OB0WpbZtDsXGCpbIJdU0Aiz
xV1uAwX7wUbWJuDdC2iAuckLGcd815AD6sOJ+uAOrT6UBNIEZbhr67lrx5567wY5
CK9uly4HC+xoJ0mj92tuh6g8RiEEpj8ZJchEcUeyPznaOErIis4vlDf8SiEBzvQG
E6a1Bi9TFxcRyaFiQDBdkBb9R9bfdDLyd+aeeW/qTPQVM21udd3KjiYHxvu3908v
oPRrH+R0XRrnoT/o/0eguzW4vccYV6L2X5dA7ni/vqM1rgnYsFrM1dQbDvVFex2O
eMEwp+TQRWCxna3SRjf4aIz2vWdIcMrFLz1THrUBIPnYeyCnFl6l49NEowI+IjUe
6C6eEx8UNBFTp7AY8je37MrHfpuMAXQyI8HsisLIEbL9QD55RKTNJtLAiN0GFyJP
J85OjmOeP86IXXgfwHnAcXOozx9aUTYDx+mxFUeR+otPvBnkqh2D7cxCRwHOF6L8
GR90eztw/mLATqhINyLRSwqOtCKTEtO47Z/3LObeihuatFdFD7dvydgSyXA3dlYP
qltoZqmFpIoWfhTscDFPSWAdNmj48Jz9IbDGMHZauWIrwSQ8xxCt1v1K4YF+RSo6
Drk8Gy2TmVPouqJmNhVaUeeOuSoL9kFyWhWInS6F3tnvi7bAKQH1a2pgF+QgGNYC
1Wl1A3O//50ks6MEBjg2gZj7qV7I8P9FBvfPHvASMD4SCd5Y1zxDlB8pEi8TlyWE
sPxnRf20+/Aaj9v5qmLqFZ+MMoFsxu/mgtsPttmXGdIQdmkmc5ghsVrhVCfZRqUV
Vv/WxCNNHOc+6//hsu22N3mdHzwaVXQLf0wHrJRYT2oqILuvxj/isF66Ra5wGpOR
FdljPkar8OpxaWLCnbFmkxz9Pv1rz+3CgRLfJ1GD2zsXPd7sdBEUsx3thd4zYMZo
97gQBbwZOf0xCsVBVVkCjo0TDjhTnixhzPZhr75GywnSIKPWY0lC1FA4IJrHJPqi
fTelGYoNIQV4WXdizsFsqkcRCP7zEg5HS7shgmTyLUfEMWfKB1FnN45F1Y93xMes
/Dq9faQCvzGjmnn8xwNBDSO/OlF/TiCuMoDblCEYLVguaLOB9Q2JWEbRXrVKg5ny
x/pOZC1rP7RaQpO/vBE3fNbdzJfjz9gZF0PedFRA0e+Riq+bmnKOf25SZOPJPHPg
RQsS7x+gJMbgyFBu1Pg26v+NzVmw1w+LmEw2psYBSM4ryAsOGcOc4SjCkLBU99LM
elLCHljByDouVsZp897s+sfLvjMuMeKo1Gex0ief3tA9sf65OjLO1OMdIU330pNW
gWwns7R2WXMkCDPGphDxupZf2Z+NwgFvpYDnNy0cejYsKNdgvl8PB0t4peV+ql5h
7CE4/ZRczkdSgE+DK4jZNAzldIJnAWo8xt/ORJbwq3cOTbaOqOqeuskn0l/7VMrL
2McfDcoGOeTDYkj10WQHXmbnYk4ElnNonGbb0zQioiAjocHludKsw+46RHYBnsiu
DpUVSmnniKM/E375Ci6UMCrH7BfEz92yWSiPw7XE/oOctD0p4+WMAaNxFR7nVZh2
wy7VwktdKI7nuYEa+uCvQy1eBNx+M6xbmV1ofubhoCioZcJKSvZXSD7VMB6IRbPT
cXzzH+WueqyO7D12mU3xuOFP0Exc84FvYQekuZS3Keip9mNYmp4rJNQWydSKV6RZ
UYmGHAyMkxe3ECbpg+jHwDlUrbTHkz8GYJS5ZLbZtfjdttcm0NMVQgBRVFWlsHKD
nLB5/eV8HbHIO6MrUIqjkH0mgL2fsmeCmhccEkenBZEsriPt9AxmG2hnx2cbG0aH
DZA5Z8WjhXfyMK/YlSXvuzixh9d4QspgZtFYywSy3Qha9CJT/XqPB5RqifQtfJEh
5HZr+kBfyPDEVz4rNt0QxXmGw1puo5151HdVyqJD0kC4OBZxzztgaA9LSCSKJg3m
kTZFkWZrNqfyLQCW5eb4UtZIerZreCIgweZxHqY0caaMsEqK+ZUdheegKfnyLStx
9CaYCIKJG+SNe9PNPE6zf1xGTJ0jkLQla3LxYWTbmYd5ZlcCstSkNf2wLfv5eK3S
6oSWb+UW2bAJoaMEB6BcQIRa/HYg/SiWgT31YZnQsGg+TIpati7SdFF1ic7dKWEp
3UImOiUUIO3OqKwlLmY+WiFV2opQbO+LPi3ar32U7cEYGmFF7TIBy2IiqIkTOFJ+
pOQvoD7HGtMsglREP5LFgfSmolpb81F3ENq8VV/oPjYEC9lWKMuzVBHqp4Wsc4Rp
ukSD/J8e1059ReDSDMP7Z+exXAviJLVLSGJn7ONY/JosO1NdMZ1YLR7yK9q/MtdR
8v6Ji7ED7FNjXLHnBqDUf/3keu6tC4sTxFrO24OM0L5jslbST1a9OyPoTiQn10er
JBWQo/eo6y2Bj3KhlFNRILTg7uJNPhClkKhERdRXKwS16klRf2LkS534oFZxeG0H
DdjZhQM3eB8SxX/8XMplVKEb9OwgT3YNqTsFjBh4b00NiDbPuJJej/b/DQ6yvYj8
CbbpWfpsae25p0OaIbweykqmb565dUEKzE3cC5MNDkoKHv7VV8G1UIoVy+FliMX4
yqgL3X1V9jqYU1SHGWOn4rknTKv1irM6CcQPdu+3SPvGBq20G/ABgoa+aHGP/7S2
VD6moMhPuZ0q43u+InAaWRwBuZuARgfxgEzjzb5oguuJqodKpGDVxAxQcLRaPPZK
DMqW0/gCNcXO1jLJJ3ofUICQXMm1AdakGvJHpQlbbtv21irDNwPuyNq/AW0aEt9s
h7skv4jg1X80hqdbt5TUTYOeSJ9wUpPSQkFv21bVEeZ/1pgzFbVudhFif782tasR
L9ocWMC+H9h6BIqanuvw2Z5uoDqJWocVPhc+m1kwi3C87UxhvoJ/BtK+A6l7LxMh
kaqhhg9gXJAgE+vCa45AZHWElDSBlrACo6pC07qHJVYHr92eLmbcX+Z3BpMddjwo
bFvqNRk+kE5rM/o1CdozQHs6R2vB+bm4gsyXxY1vZm1f6dUjle/sPYXxOG/jUAyJ
YFdEX8KCmAn0v5M+ufW8N1/Wpiwb4ctbGW579kno6zSUlf54ocTwZC0W4XOEoiDx
MN1hh4g4fJyKh8J4IssupqSr18WwGyILARCJPmcHpvK1QMNvUEbQSYy5EdYuBc3S
6ZbS4SKj9CScnhPTLWLu0H9w4IlgezHYAERHyTx3ucsTn4CAH3fBReXIMHNDII8m
fdDgAMkXjXs00sg9jDANYtJc+L9iwvEmbUYMfHzxQsVvPCK8Mdli7W6GKB7QdUTi
IKRV7E8hpTuxgLt/9VX5RDMNjwFoeEMA8wuf6YNDrUN7wus52FOcPcm/1blho7t1
1NWMV0xJHzD9UPi/5SGYThJl4i1Tkrx8TfP5c6XjZhJQWMt0Yx/P4TCRHJ0aW4e3
9XOgGQ5UApIlQZoZ1W2atdesApCybHGxQ73VNzIIEb0/g01SGLctJ7RsYmk6dJ8N
KsHs9wem3ei12mvm7hm/3KGNFJ6wx60KjaS7/fbR54FTwNzM3vkjcBJUPHBNqeO/
d2djzbNpe2bY3Xv8rYhY8aoOOtRse0AnLr239Krx42z8U8kfQHxYfCrD5T4OD36V
75o5Zj9tKCr9x2Ml+ZjuykiCASyxUsnP8WLZAVfhNoTZ8ss4KAr20N/jd3kWx/w4
meenRA5uPxMyGm12lUwokpTtRjaG29krgzKsvESRdN7UtvDucZsl48kGdsMKh8B+
yKHYNAfQKENivWz17W0oASrF3hg0tyRWaUrb22r2Ake91o5PBw3bl7ObMuHYwb3q
UCkqytqgWvLBb4N/Frg4SQ2c+RLAauJ7ZklrIxlakGNr6YjOQbfSvwLoVvm41KdE
NB02bSy9g/DURk1HMZZn5riuFLmiPy0sbu+IP2tSyU7wgtbXKZ4RmxvCtXnK8UMe
ccxEPbYKe0QJq+xPwhHP3cQEQ4lHylIljQkq9MlET5SMs5V+8lb8sGovORgEQ+aD
bKykviJ6j0qMWXXWpltT6a6Ei8DIUAuUUA7PZrKE9Jr36oowXCekmxZ6wFxKN96s
Ao4djPNWpX/NLgi1lcVNsZFmYUImOACWAkUG4TXZTF0K8GKv2Qh5KN4xsy1BzZ3z
Wd+dw1WFenePV8UFftOrMSrhbIRtVd6R31ZkPoBUMXytUvwdFOK6vLpiOXPnVlG+
K8z/zLRf/VjvnxoiXBdky9i+4F68nR5Tnc028BxkLyqA2XVPkx7QYfWmrNms4sSf
OMQEZNkuIO5/f9DQ/DQHYnUkyJj27hq3+9IEXIy+WUWT1ucUTIWPBYWTcln+r9F2
U+1NRcbwzmk3InihDiu+QymdQmfRIrQ15iGQZqQcWW/Ce3nKI/GrgV5szn1VUF+t
a1GaGxNzHd7RTqICMKTGKE7pO5xfwmcFjLz9i2wz+B1+6u6x2B87unzW1V0Qp8PN
xVLLnI2DX+djcwscku8m4l3EwR1qanIEWm8nvQYxcIOpTGgPGiSdm8HSR/MC2JS6
j29PT+Q72JxOTO66cC5xmlG/R2yQqJbJniZKHBDuQ07fXEMPMJOApjhBpRkRXmcg
E9m9gozwtbC7cBlneR8rLuQJedp19wJOFMBGJGSgcGSMiEo/OuUNU4rSK82GTlqO
uGk1qwUKLIRqAqxJ9S35MP3yzH/KqIp9v+bPeztBOFUEo9wRyq6SPvO/QSTnToNh
RMDdT6/WGuZM+/jIY2IoRQBe8TYXaJLTCi2Tq+p1Stf6FN6wf4+NRJq0H6sKDVvD
ZmcTWK4+WAfr1Hso3NTOKYh4BuO5618t6wZgRy+QXqNtDPSHX3MwbJs9ZwykoYQH
iePGGwiMqGO4Oq1ZeakJhVBGSU6hjLddWhm/L0VxuQ+kRzpb0hSzQRN9CbPYDFjy
78x95Q/cPp9d7R+htsI84p9LDlxSBBbDPDgn4/jOHIRTJyPJWoWyFwXjYMwEDDEk
exGS5eqUztP5zT0VtEdRbh83bO+sYKhCvbmUT9jw8BaEHjpj9w35gNlGQJPpUqVU
SpsROE44Q27JrpJUYjtHV2vGVodkwUqGBMDR4Bh55qXP6FfUfAX4jPx9MHR8LudS
WKBy8mdAI/TSKVLRP89vDIZnOEQiULbwR2YQ6wNlY6vDfP6/E+47rfpxpqgDOFB1
VZS5CDeBAA0ct2Vx9FMXAdp4CXrB+pG8hn4NGyy10O7xdhoxvzduJ9eaLafxii0T
/Yvho5gtClpmStbb+fVE+5g6wfeDPjGsCu86yGDDweO4ijX9wGdvVk4uWiGWg5Xy
WjR/sEF88hvimoaCtjHeOuLs3/fxZWVrXf0U4b/bX81o66v/rFNLBcBlu5csF4Zu
JgCdpiE4MWxP6jp/E3X3GuIPSfX7wQyXOVAwbR+H/mKnGzjUi1hsse0JjnJCzdte
BsaXeu0Nqc9wdbwXYcsKE4oCfDad4VIlH+5NDRIfSzWCcWzvI6gMi/RJ4GcqeWBf
fzRzCqGtPAFxO0BmWGf4fFY6iCt9OgrSZja7q6+jgqUfm9P6PZaU9BkUl4U3d8IR
yDtWVTX82bHv48mddiofzEH241NQIEPS5EZu9QtG7Fcpaw9/K2QuKb+uncaOUuDR
BZ9yw39R9AoqVF0BJRXMl07eQX6wnPIGggaHBJp2Pk0Z8Oi7F3vEFvYNGcQQbTh4
rCWC4Bnv2vigUQpAd+tzW0wBD1WTcXLVxpI5tBK5QKG3SpSJjZSL4VlnYVddT2Ce
HGnDarGxYnvhmXIspM+OC9gExlLgY3KB6z7eCVyhI4uFzM1fXyHYjZ5cGW0o83qY
HaEHJnosVkLfUKM8sPc9ViafdjBRcQPMy2abLK1sFPMCTuf2EPlInqip71wUFqIq
spf5MTtOISYI/w0T0fEpLRZlCfwc/YP+4UV1jovh0ovUw/TjMt10Tf4KIKNVy1S1
74Vni6MDrl7Z2x1/V5hL26COmmpKSNWI1BmED0dFlwfWyZhxqhSYvo95/is5c4b3
UKZ00/OLwjjzK4127ihsRB3KeV3/yAUs8MoJJQU78A6HgkTWHCo0UpmtkFIG7/2j
g5l+/HMtBkKn1TxJ09dXByKVTfi9Bkgy1U2bnHXf2wXkjk/wHjcLl15MfihwT2XW
M0VNPBki236qZ8IaPCN2OrE1oxHEjbcd/zfg8dHUguzj+jnd0a09oB3n503krwNk
/R/LxrE8Zce/QPcp2gI/V3bqsuCJkMjfS51axMZwT6Xla6tHghc5vuOAaVDcyc2O
4SbamyN6M9nXCSmrFQFvRjtgVQbJdJfdP+XJT/95jnSpa1iftxGypzFnjMIQlo6T
J5rLIsEWHkEGhPwXCr+NXFeVa1scN6AbOz47tPy6YAK7/U50dkJ0H0z8fymAG9uw
jcy+BfPjW/yF+0eL8cdkjoNTu8UN8KTQGluRJTKbL9ciPew4bKdi0yQcCvGenqRP
Z0zArDuFQH1Dcdmyq3ncIfM0rePn8m8/5pHzFL6nhQEu7regq9sat2sYNoMx8WC1
SaqOc6ai6tRB7BafdfoveeBXW54A2Agy7xL3H4byJYmUv6AzJWnNfe6fR27+nUDL
4N5VCpZ/F3quS9RiBktIsQIhtP6cEvWz6xhvMYZCwtp1dl/USyFpwaXHsRYUfLhb
KwXHTg4T2Q7Bg8f0B6Ycar1sYuZgeKjMXelkrDeA3/2kdPosUi2trFfzoKAScf9T
N35vcOfshPaeqoDyVyWroUNG6TFW2rVsLQkt89Ra1JSNsWQ026e7kxX2MWVsp0+o
cuyc6YZYzO/6SvJxVa/F81I2UR+/sNBIK8mggM6KsN1dGjPZNbnODmatbZERpoUG
6oUKla2PkzpGeb80TbPyo4nWiueYorjm4WiFl7G5Ns9fl2iI7VQHFzm6QSkGJbBm
nz17mlMe8sEVwTr3OlEc16PAMaz9FV6dNkEF/BNmMt8hGv154JkDyab45ASquiku
urF8qwCIbS7ImLUtYxu4JzBK7c4o20pYHsHLa3VbFO3usym3CB8z++KpvLclOxxD
XR1TgJ3S429/z/kHl4PsBfyizExijsGjnnfZR/yhv7jE/3dX6d28vV44WKvsLU4q
iZhYBf4pczD+bdGCerfkjmFSl43SSeehzwOuBnx3RpiEDGys50VzRqpMTydBA8b5
PPRXjOCV2K33If6PNNQmwmmVqv20N0I5KhqM1f8TAwYbZAHBz7JkXtDirmZZyHLY
4mrGC7adVaxjG6Zk43npORM4ooXVAzFw5Gw06m5424NkgQ7wn+ZpCeUMUWt0TA9k
8fMLjH7eVzUCLZxyvNjya3gh9vFkL34Ihv4ROeZCjtbYmBRjjjSzOXZ8KFIl/WLf
/MMErS8r4y1Pk/gPZ2RE1RVlYnnmwA4MFvf3mcWhatS4otF9PJM0a/MIF35XLs3k
GUIioDh6j+2wvNPmzurlVUGxQmngFuFQ91toHU1VK/TXtpL81zZ/ExuTSqRjJBZ0
Q3yj6Hb4ABRp7pdk5N8RYvTUrn6IUPpH30x4m9Tx5cJL6Zw+pZ9cvmz4DBfnfhTU
5EOe+921F0Ctr7EJeIQ4BwenBpcYMomB7iCO+GwjfT2CW8RsdgWutR/fl4ae0XpH
CqIj/W+UESppzMPBuKvnoGjPIyEyANNuUwzheBsEKp42FgSSmpsQ2zu5zBZz4LKB
coqzL8SVq4iQJJJxdGr/EFl1TTjXfzt6Dr8ZmYQzgt/evJxJfktA8ryMI3/RVstg
GyeT1VGRajo0P03osZ5tgFwP6zwJGM/LFCFfXKijCLWjSmei6YNGyjtmNfpH9EHN
PboqIFJRKlbhullaT78nKl3jMWopJphD/D042fURZ5qwcerr1gdnP27WrkMmJp16
WEttndEmLJ3d0vllMMmwmX0A7z6FJbHAuVGmzLGUM4a9n0HUHW9GIF5vwxefhgq5
Rfp9ebtMdx5eU7vQrfZA9nmmHvAn0p5fq43kpfK+gN/SqrJpO7BHg649gMO5xRSl
OARRaDqGy12NW+CmjulLo/3N6qZrYY0NylSDBnaUoNaspTKhooQSWZQnfdPh6lnH
TwcPPAhby8JiayZqPifIu+qtzXP8mubt0xMh7vZW7lx0M+fb6JzAyaRvxx5dH+xh
c0i/Lqauu4zRNlbYqaXEsqpKt/g304m5/3oufU4IW0na6eZgH/64Gwu9NXTBsnv8
4ugjV/1vFPZ7+lZpXd83JmxRpEMXz17M0UVzdIA4pX9OQSnu6xQ2U92ggZfz7ei4
Jbc9xfnORT9IJRi6z6WjOBqiZn7NiG5yPSDH7viQ2UZX2i6Qgr6+4XqWhUbx4BPZ
zavfAy5hQsiASPeR1l8dVGblxrkS0f92cdNOPv5d1f1TCVLPw3JXLspoE+AYqRI7
zwLjHCEHA5im3Cj4lROEjYfdmkTT9HQz891jURCfsGnlWiVIe1eIZf/kBU8YX47z
ef5hTwCFt8nN8e6hJNmpgZk479CTdVowIrO8M2Lxgqx/oZq3lUnN/GOC53cCjK/6
4MUQQ+EJ0lsdpKExrC02IjlqJQ47BwYsI8xmd3GRhGoQ9Ji5vaYMZaiQHDQsAnFc
KwKi/GIDTwKCsQYimApCRYKydQYLp4kSIdfxpfEEYs5kOKc8CvxXPsLGPLgDkh+z
LMv6/fVM9awy3/RvQAY3HcCkf0gnsokOaVlanFECq1qfl3v0Xm74595tMjXwDlXj
ag3KS5fow2XCTHNLtbCbnyjkvunF8EgK0WM6/XXfudYaEEkNihQonX6AJdHiU3Yl
7IDxxHjyiQuEUjavHjPz39LBlqlMLpN8Vzqllx3hZ24nhVBtqDlDhFeG8RfAVyBX
Qb8meAxXm9gkVTzFwYQuLEGvRuH2cAjoo1Z/88lKrJL/BWBX1DvcuKUACmIOIgA7
JJ8VtdKUYDKJGVyxP56ccaR/m5jsx+sCCsA6HS5TwvKEXr73DNyU5CG932FkeX4l
2rsVO857c9BOK/SbkJQzBTtfAr1x7RQjxhkpZ70RRSv6av78QWv95JWEgM+DcatS
0P49niUc6C2AGHESoR8Xic5UhRh7FXkpPLoDEvqf09olllqvHBclt4P73WHyNhGA
Ew52U7lOhbCVwlSAa805T4kpemKtDA9OowqmTQINttKK0mSGnWa7fp7H4BLRYG6q
DM/caZZ0vlh7vBFaTDaXIbqonrmF9WR41jJSsCYDodY3Epk96HcpVAoQrlVxSuRl
3r1vYR1io+Vk77m6w4sV3cRdIQtTVfwL56k6LHDOiISAnyarLskIYI3uAmSgv7rI
BrKtAUNXOtiPb7ZflLxAnaRxTVEi4sHTeilIgnajd5i831lSvgfJzqSBZVdNStGK
7/OGzATdKmrXS4xtQEP7soJtHB11EgMkZVWH4976qeJN1OaW50y+Xpw9HVcthBw0
NtwAeIRbuTE0ku2Ga30vu08VZ+/V9eH4rot++B+f4FvrkUyj0bBklFJWHyPNo72z
Qzy8XoAhV66sMnmJTinjEMxDAnxeiM1JgKc4k96V3JAEHR6whz+o72TSoBr81WlL
fiAXhyasFsGG6HfRCgWHSJCA56MIbtSJGksk0Jz+60zZopDv2MEuk4NK7TtjVK0F
7hKFPnvYTDW977bBVHJVaJywJj0P+kSyUFdZjk/GNBhPceprimlCJBRl8KPG2HYb
KIMvMYtG49oTi/hDzMBP1iQyGmiL+h8JUGTm4MTmkiZ7MYdI78LxhOcFXeoUZqFj
RroyqAvLjJ9KtrEuU9jNpJ6B8aFFlUBE2TeMI+BQEY45551/S4xDznWBb4Q53RET
P1x4qgevJIgm7QsfIz2S7pTA8v5XVn2MFjQcQOQRZ1eZQZkjXDwO7eadU6c2htl6
WaJoycN87dGQ9obZc2VApxW2yFhJNG0ctAGh8F8jsXK+KLTbxfWmuo6U57Du5DvK
kevROIrKdop6N7SVc6BPwc/RJspHrlXwfsSII9djWMr++xQf18Og6RM7PEBPq+QS
Xa9x7f5nzJLmYBqr444wy+/ml7t/WG+6taIUylhEsTIfPMttAvtCOJ/9hIQn7f6l
/42XccBaKrGtpGw8duGmplP8ZQUvO2zy0N8yvWCSqHnY/+0fJOh95pZf0tAGoSlc
k0wfluJowpV495CoM0EGeX5F7QPKQQFGTQGWMAwmC3wi4YWx2b3D824udsBqGUH5
BFGE/IGBg8um2d00yyxyHM7AMgQ2OZ/cw5nBUKGw9YwfLx1XR6uUDisJSj8Ps9O6
yyz97hmruXnWkf4QSWQhrVDG/pvJICO/vcbKuXbrKUSrD8hpObA9Id4Tz+p5k4q2
R4DDrNiDvRVN570GSO0NBvtws1nCHydhrm28HcSxmBdGfEuoAKgjoDbH7dqNyCVK
sdt/oKuM/HzotaDPLKTDIaVaA7eXJAwBk3a75OlfBsdpVoo4ta3JaYP5KSzku8Gl
X5dFjftc84v8hv8tK2zlxX32c3clpfE4IjRPYWNaWhflOh9EozGlLanlbcA7l826
LZ/WLE2FScwrWjmjBGgbsVcw090QLKWcu4RkbW6ucVnP1sOM62zfQE/p6MPW376y
dSs7aXz3AKxGniqv1DvJj24uywnXK4II654XyxJVyKuGyYpbt+UUzAkqQAlG7jwx
twklqtNo2VX2VoB8Q+2iM9USzmVUDCYhKDkGYlKIfgVcXxpetOEWgjNaJ4DY8Xgk
bLq9oMvRS9xSTHbo3Jo1Uo0cjfkkRIjk4JbvzRupwQJFGhKJibio0pTK9dorsDvC
AIu6rSNQEBtLMk3wSe7hleDMe23IW/ik3v7ocJt5C97gr/eu13r5tzigvSNwnuFJ
iTpntaFtH4G5EuEZDhtUEpBuXEbapHAglLCWwCASfrVS1Yoz4wzx4JxagLAlC2Ok
9sdIVetBep/E6RdsVDBwjUMVsrK6rt4A3aRB6wSTkVhOvpNC+8Uq7uowjgj+mvkP
A88+ZsRQpGJ3WrIJ6XtHybV2fIh1eHoIbVDu0pHSuvu7D8qbLdoQwI9UBjUbCCXA
V4aWH8pXgmAkQlOUKUcZB3Ca6rkr+dtKbHkYkgRH6oqGBSaiUEz3RpzhEGW1gewT
Q53K4Ulmkfa7B5yfCKQIRO1tbbl4hm03XoCgDX9xT5pXgU3EW8TbrCySZZKezrgV
TAKNFUX+KWVwrAS9vzUSIsLrlJyLk99LoyZfiLW8W/CvYZbJL2Qwdu1Ie7fxnpzi
gglhrstIbgobNqUOazz5TFSuxx+aeX/y9VX7siqAtutAciQj+JTpDm+4lpM8lLbA
kDXIiV7Y2m+KzxWfOQV8hrpSPG5YJwSOixUkMhV4zJCvI7EZaDpEqbjcQg17tVf2
gDMBfJvU1c4obKx064rdu0ZZMCws81oe5+SLOH8lKJZTJNb3dzniFkV+cy8g0hSk
B59bakGObxWhP/1usIwRhw9VwnyEc+qbF9Q6OFYmj8LimjFLo+Cp4LLLsSnMndWk
wCHC9dq64xeN3O2M7cip0YMT9YC90j60fuTACWxEI9Rffwd2qMyxTCT+TWfHKi0t
SV8JToT/RT+mA/ZWLHvURPbD7mtTADMtR7XAPu3MeW3hMUjhkYVA63M1Qmw223jU
a5yo/+zQt8eYdQFMkMIkJYXVGHyyM+vNZXh+4FzA9//bsQeTn9T6bfiBSMpJUKmW
DdZqLxeoP5yeYxsDQN3ehOuBvMBOeLID7AdSNyaIDGg6zrTq2p757wqLpTd5AMnF
IEBDYRpqdvQ+MmhRKOCTsnnbPWycQwhwYBQ7gV2TdCPPRMZvqOS8x8aibCTPdFmp
EZ9f2eFUgfmiH0VdIyx3CmukExZ8XNxlFXYWqlK7oJtjRGZDA3avxV2zrHJSIWIQ
fAzi9ucKaTogivNEu31jJUs/AUM5CDOFEm+/63Wjy+styApsxxf61P60llJFJ7b7
SV67Bl/meU4tuZMPR36F6Uyt8y1zre4PKfolfYIZRbJZA1C+oYyhAiceKRtKKvwi
jNfLVH8xxiGL7GcmIGPWtXGAnL6C4E42MGj5RXRZ18b4uRAPPK/TEqtNYKRNlVnE
Et058tYwJ1RjBzYQ/SbQfFutYXtImutHPS1i/TofRWTW2nkW8opkAehFTaA+w9IT
9JUcpEafbTXTUzReTwOHTdAJJFS1aWx9Vv3xh+s0PtRYOoekGq9hcquZOXpZR1Hj
ZgiEY5IlZG35rG+vMqn2PcMbOP1rrQSSMI6Y5jYx5h3HxzLVdaMfM4kcIucKHFiD
aIdXO5J7Y80yd/UZLhSpwCED9SvEo4AFS+RSOFjh7ygO1BvlKO6OotA/v6fpI2TB
hlMuIwc8l44QaA6MuOxXJCDN62gxDomQvjASQZvMH5/wVwEoKRS0SvlI2iXDhukl
OW+duTzBjt38orTyn6010b4snRQ/+Ymay0N3PSv8JnMrvS+QIvZHX7ufsmQPWz/K
V3qTauV09zKpnGSdGI4ojPQEI0y2xFqMuMwtVBFxY8QoxXXxpUxzwng3hhdRWgkk
FV29q58z0t4eXwUWFzoW/ldTGSixOQH5g2PPSmUI68pZ2tvD0hBMJEZDeI11OpjM
7LbhJzmcml1M2UKddpzCpHva2xnUxxI7ur/eIBbULArYLobA69cPXAgCPdhg6S5q
id+qe0jHe5xACWxKbhos0uy2wTB7ypzde4yw9zqCnrJNdPrDDCPLxeoOuSTfBAMg
oLNyUrEni5IYI8zmW0jb0cuJiWFwGBEXYFbdv05DU9HF34LgY0baaD5jTRQaJmPu
Z45ZCcCorHlpcaMnWnjbWbObm6iWDwrbWBR1gHXC2KIx05kkz0/WSJgWIvCyoc/6
ua4XG4B0X12e+GoGw0xO+WgwxSZxNcg9XG5Ojb6qcLGxAB+m4z5AAFyMsC5TMk+S
wbtOe03lZ4wGvKko3AHxRTgUA/j/mo0XZufZsoWtF6KlpMnn8aQiH2+B/sM8hVxY
OkNlCgkE+8Ja8dr5s1e1f7j2g5Tgl0BZ3JF4PNPBPvHt05BJKuS5CNvxmArGYnqJ
zXOaOtO2S989h9dS9+KtsbcDwSgLu9P8xMZ5KilhGGCRGpj4e/H2DRUl6WIWe/It
qlElyt0+SRkDnqKrZRhRrHtC/ldGSnzRs6o3yC5AmLNFhxhwKqBkkNlgie7Zo+n7
jpS0laIDMkYuDIh4as51ojiNVqLG6bmf275f2ZqfyRdjLUunt5PN8lYOthF2O3ce
HTlUPRCOr0Hm5Fnaz275AlrVK2eEJOETMWVzAqZdCepay+SvA4EYLcTgawxjnR7/
0Iui6dzl9icOkndTRGZDzcGmkGRxfgPyWIYXqwiP+kfOmaVb536iul+3+xAVSPV1
96wK7GsxJxlTZedjU+klIEMyS3qX/QY+bMrIKBGiXnIf0ICgUzo67a1P9RYDAE//
6SXyp+E9e2Zmt3Sfdhl99epml1s6t1hcsnyq/VXIBPPBoTE/VAueqUc+IZSpRmHb
bPPQQC2W4Xm8QlG1GYkNXUZRxLikNuH8eYWDO+63Y64VHw/CyRJCE/7P0TmGZBrx
6ic5jeGI/GBw0QOFcziUkxXvEVCP2ae2TkoEHaSLNb3Bo8dn3LBS573baPtAxbG3
TKFn1jzYLFTOD5YzmYygGV+CiyteBhXAuWDlZ4r60wQOyvNyhA0rsIDxB/byUfxN
gSuMDFqEyiZYAwM0dLuvMifRohIqPfcq5k6T1+2tpgGB6EVaTsROrviZBKG13Stq
Y7D+q+NDz1wi/H7nFK346Pb2vZDOC+daRMy4YBBRpG+mwtgOL5qAMUMeb54qMzm2
YRLeTf0pTV4RxcNL/zMwRtu+7WYaFuW8TTOjTcrUtszClLnAAnXzwW0koaa23TzL
HRXydnp2qcAsA4ZF9bAePxWRFx11Q80Fu/h86Be3qyWeNdUq2DY/bWbjob5Bl8HC
7B2EUjI9/hqJBR/H8hprLoraKW5+SjqQEr68qtimpmIIRKWvU0IDNjHeJmyX7lAL
3sLnPj6Ylw3+DpYGCYsMiyi3MnmeRlQnOMGvU6Ipc+sojFMt+K6saVDTz7iiPHgi
stJP26uNHA0Zi9fDH/ZVC5h2z9NRByjwtDmUyPUObUwRGQnKEQ+At4vLmb09oKxB
s3ggHA0QDBhxSx/f8q/P29I5Gbbmk62sfS0F8UwcJJWoikME6NgeNQ8Qydsh2cDK
haGel4hCLMky9FVSuVRhuUV+i5W15KOeTU4v0+kEVE3w96lSqQ29Hxr86JipyCDn
OTzEI3Ot2AzOjVSwaJHPvd269REO91Wz/WHCrnTye53d649As7ZBaQDzsTBC+2Rs
yQP2H2QUJRtpfrQGt6Q918Ro85fAcpLWc7x/7dN7WyzotW+DcPdVMECQuw+yUp4b
EJaEh3zMrY1NasjoCFUSw+ndoufxLLbhSVUAmPv4uTiWiEbAsK0UnNNEHQzWPbZu
Sg5ZhXD78G8pRYTja386BfQKD1NDcxEvZ4NPSGBYVW9SyqlXIJZoapxSdxz0R7Fx
KOoNiuzieu51vuDagNve0Wl/nVCF+6ZDxSG/QSA0yQgbJEBAj2+BQxNGZRibQOnI
TZ2spVleLmgVufCB9s0Z285Ud35VqLZW057UPI79TBNDUh69leIdPEfwm1/Y3wQH
h5dQjDTgSN1VvPlnZRqT68AKqX2bA2ISa1Bm6j+8nYCyu7+oGbOxQl5D6MRdjQkm
EF0S6RRcIPLBbwAQnpGyQKvuxu9OoPPq3AIoZyEyp0feRfACvXBCiOLfi3PD3GXk
PYShCT4acQdU8WFvydj1KQ1RZ+YncFd4rPOk5qrSDgbPLnAdw/0rcOoH/FJYA7UH
rSqpOxhn+mFxu+WhzR2GHhs06prYrF+bg77m8g1gfi1ZqrvjSTxOXLlAhnMuBo1W
TcwVRkNMqZqY6GQWTg/7feYPXQDfzsVD9W5mVbWZCA5iR25EKa5rU8ghSw4WYI5A
RCwAUavYAdJy4EOzH7EDY4BosfGo0BsxvZjR6oR2ivEKJBh1Mfv83cspEvgq791R
cFmopR7bgoZ/ZJsCWzPfANmWXyxt7HooB2roIrditwsE8M6HIsDMz4mwglzH7NzG
xIZW46YfOTFfkbBaUeSd+Qc3kuG3yHtYBJxyCacyN81l+g4ZvIbNXNlRtmCMKLKq
ZsARsdZPOyLsSutp2WgjfVyTkC3RiEt5JddE95TWDarJF4qnUz6ccCAN4/KjsDN6
pV9ff9VSv67Y9a/r4ZUNe/bCW8eMFEtyzVseCAuKiFjqBxM4fkJb1SvbyeX0sK+m
bV939U6F4anMgYPhgwhL/rHiSYl/lv4I7lSkz/XNJYztQ1ddjJO9hmYsS3W0NHWx
4LMRqomAqG9QU76FInflI63TyA4VIz5m7DbGIC7YJ3QB7jnvuxQPlGlU/FM6s0W6
mcVEb9yatYNLTYFGv2T/vTwXYApjlNHop7XNTGpHISBNjeF6PNQaGiUWYBTGITtK
DEQGhmlEgMYIsGcIcwD0twhwCMUWumITIjO/33U6feq26FhattYL8vLbOoRkjOl/
wbqtObdqBimw0RkvoZl/nVqWrhmHfM9YNViS78E6lZFsC6QKZcNBi9G4pdKzEnmJ
AjAXj2IxW2sd8CdpX0XMBLBWYY08x6uWxiNvWsLEmN1UHWbAKq8lAIJJFl+LY53S
bklkHJpeGB+th6VzjaA20ZIu0IzNGRsVBSy8E/X6w0D3NMSP6vmJYh5t/idDG5QE
wVyOd/RHyiz7TcM0wSmbzo6vHngHd6keZ9bgDOmjrLUEVM3KNlI2EyMkI/hhCW1G
ewJmbfTVFUMQ+15WQYTiRodMCQblaZGwgaBrXQ4+r6VoDW1hR1UTeVe4xCtvn9nm
MuNrB8t34HysP7kdWlykEXov1MZehceijkdeuYDZG588WOgKKKDSShEJQS5IIgxB
bslBIJvQppQgKB9DOUIWL8Eg/eaonY7PV5AXikc+BGD20yBNhzcuzVbleNxVCkFL
IWkQi6sD53Cy+d8Sw7nMsphBTF8PV6afDPDm+5XZAwOhBPjGZawxJC8W3NVfsdOQ
kio3CuOJwtdgiQVcbZAlCm44+RmbLhDv4PuOPk6rMCP8MroDWN/ZfSq5E4ffAFlX
E/Gi2CVoia2kOkrAbwThFwURjQpweWswGaVU2S0lC6g+XZv81F2Eh5Dq9o8xC86e
iRfYBnDGtj3jNsKoxkCHRyU4F8MpJJiRcCPIDndCFx+Eo0OTdac9qfAmDQVC0OIy
KgQn/UZ+uqjPoNmScB/2P0bVezO+j1k1jwg5dLzcBYxy2Mj4X5RuYXF6DgKDGOuu
hzMmKCCi6r9w6iBP/BLleFJXgAD7CiC4J+A+Mc4eBRQFUGcjgjVp8JYTL43+1EDR
PNE5m+NrxzGlF8SgQ+2GImLcrzTGu/BNip+nBo/w83kusTyXU8QlIpOg+bJ9noKL
rqmBMAdfviDxLuyd7fjQGqx+7PtPtS8xqTBIGGfUYpLjZqcQ68H5XO3euisgNff4
bFgS606HQ9q6d8gdIOun2i0TrTQ0/cVesdlU/w/x6PHFOWj7W0oF23xeYsauzb8+
SEIyU/t/4dm237fpdUniYU5WlV3zfNKzOvzdxjLZOb7xYOQ6PS8Mt9LtkhSKSvpE
PrRoEzLFLRXZQUH1FqU3+waEqSrTvxnCLjIe5Qe+aoYPen8QUOVTYRS3le6Hmmf5
urr8hrGUf4XYAwwZWzp4wMpkHGUHvJAWyY577VoXxgbIJua8gWNhcavy1ZtldjEc
OPi2d8xjW/LtqLRmYcRkCo79e6EERN/daTIyjqSxlWgWUJD0kOdyutOsj/TSlXek
kGR4HSAclbV7hh2loPb8RMj3D4koqCf2t7R/CPKkmu44nxSqjFykAl/aUbL8ioxQ
u1L5bsVTPoWfVGei+mTXATvclXjhtMjKECqMAPVCn1aGMF+7JaUGP+otjdosl0bP
ok7ZBnPMvOGyfzVQgwXzzc7CUCeGmvrMp2rp+dP54485Wi3XBPfwGSyfyXdMVonj
O4IH+2v8p9wnODx2AIka9tQxtrCz/EdkqMnH5tfRwLg1UJv6vnR51wsEbKMVnFtU
3EXSIr/g1uT1plMW/kcCnqocEVRUtajzlv7OyzgR1LaSHEg2zwUd+OisRZyNm6BY
gHN3+O0Ede0Dcq8PmSw3i9V6bX87+fU1uAzmSxHF4YlTwu06doVtkR8pawxNVrJo
XTYGElVtnyXoWYMT4q9LgLsGBVoQHgax2vfqbnpS5tjvVrVzYhcIhZdlGSGNMQhz
fqY5FjGPVjKWk8TPP9a9jSOp2zAVNrm+1qwZRss7ix2pj7nQTc79AUQNkaN7juLl
lsddRnuKupDrvrCihAtO3LLZ8DFCEF5+2joc/B5q7PA2JKxQEDtqUtfZoehvpOin
oX5g9C6Vizrr9uY+I/QlqcbjZ2TWgtE6cFSn2eN4kv8cNUy40ePaw1b22msNQEHC
SC+D+9hWV/XubwYH7/E3FnIFJjoZv+AdJzqT86win7OWByUGXr4Bl/ibXUK/llQe
Usc+bk7KolxPndd8FswjdtrGEaig0aguSpr5wvbh2XaMwBHsWPD7qykPW0NkznSP
78cNOCXVeth+EYntYlef79E1Z1K9G2jMzYLP091xF/cG9vdpXrDqLdHWR6v8DLEx
UDA9SXRbQ8CJdOcbV1Q8weFZC3zywYW9+faeNwWvvueZ6jc8qS7dkorIbajT7GxT
++1Ws4pIAqBQSQZLh87P5fpb15RC+tWhX/nUD1A/wpG/6c5SPU1MgZ9owo5jRjHr
vbBd8+JyoOotwNEOoUcYPZAQ6NuLzZGqI0hu8uhmhbWUb+AusM4ZvNwz/NHNcM7p
hWIRo8p1B/h1ypLBTLLXBQ3fKgejC2HrZGvVHhMvZ1Fo3jtJIYPhO85vmJAhIS+y
gmCGqgLN++vRYhZI9QzKMT81fF/1W489qAMAb1wubar0XWDvAYhAwdXMs9Cm9Saa
Cfc20XEJWw0fXfD1UBXL4Zf0R5g3zPbtTh/etjMMqP5zHDkD5YL9UlLnsRqNoMm0
9pcTigL83DJ53rm9R9VYsUw6aSAPXq2KkNfwZeYWhqVbPxfO07FabX04wo/6LTTl
ca7BuWLaqsZTOXN2ZxEa9CYvF2Mn5GMIxH4JjF6B7VnVdeA2YkJaLK646+J3PrzY
0j2o6DGwQaP+ZMAFv2p8YuLGsKm4eZEsEWf5Pxmpg4gDL7wdl09QldFDM1alFCAk
XIBw8U+A7To16XujKYL3LJJ9AKu3wDn2aN0wPwEgU4EHxQSHfOveftncEiRE/4GJ
40Izf3YDqaUbfJc/UtMrOPUShKkyEin4Jb25rnOt3QGr9nw5cQnvmmsMKYYw/AGz
X7xdc3PDYYZtI1Tsswsdg8Q6y1kHKJaMyI5Jwb/2gqmSWTa3UwmIVKLt8/MKqcGv
pwTiVMbgsZgJcrkJ5ZWfIYIBNV4UojlJoaOjdOTsjLEomy/71m41dyRhpIJdxsgO
gfW74SntWp+MCqJKnznCYqbEzapG4Yd5UDXHMwyM+QdQ5xb5F0f4lloMMLNxgIsr
VdRWweH7Iv1cuyXPELlZYsUtejFX8hCC/amEqqzuMFnl54uNjLIZ66/+AI91EHQL
npYVLU164VsVBWfgYYKo7L16tjV84jz0IwipeQAYLb818atkaa5NvRlwiPwCDlQK
/Z+JRyfvyZGjJQPe7TvLr40YgSMZttwoV3N9+iyPa2yoTjvuWCpSXECSQM4kt/9i
kMu8UwLoE1KTzdCySsaFGUlSReNKtqY9mR2K6Bd+nki3kK9kU5L5CFu3W2D35g1k
b7yMk2E+IsoGxJxRrUZZlr7QJDM7BocKEabEPcexOEeex6oErpKETwQa64XwFrrM
rG4hefskEkW07mHWIt+izUNHbgSqGKlmWCtZCzMVKTYD1b741/3D/EntlVejCLYz
sYH/Z3X5iU3fGjWx7sA9t1QS9eGNAGn6MJUjX80yklAkBb2hf5IkbYbyRqxqkg7A
2bfEC0tYikGBX4ZIGweVmljoRudcvT6Z6xnVVVVLWBPsvO1BCvH/OrzinCfrt6nD
65sNadOv03eZs8FJaHVIIPiVTdpIaDQMH0lFwagqfDSd5GsPPc0OZ1ojzT5w7sL4
eJvLtZqpZqoy6ds9waVAi/h3bCxmqqeThAubdDJyqnynGB8JRcskrRXIb6ggxQyh
k3+pDBVL8LuE2x4vFoFD2ZLI72SZkLTOGYvzjQ9lpoKXeg1qRo3yBxI3cDcEVhp0
+Ba5VWAE3c+nvkufE7uymhBZr1DU/Dfitwvzw3XTndx12ji2NnMMTRcrM8vr3eZm
OhA5d/aXmuu5dRIs9pBzAGBNF1H3WokhLT9TKbCoCwt5IBKOm1Ytvg5clIpTlTH3
8a4J69H7WTBFu6k/FTmJoF+jTxm0+vSHTzWOunW2hB55fuPpcA1usNsZc/zcmFjx
4nk/zS38BQk11dwxlNeP1FNINKuDnk6PSzJceJiofcCM0ZYdLgEJrCehcIW3q4aV
szppjv5fiVFlLLSGK+M7uxDsdaf1nOMikdeBeainVxlwLEBZKGcORdplX/dlU5aa
tIS7kCru18WbZ/jl1KMGXNKFfWZH11D+1UzrEMNsQue+wDbgVlzD6DVhuMIk5KV+
8o4mREuXmpLlOuLljGkI8oPY+bK99Rz4JZtypSpDkNwbod21hvk3rqZ0+aJc6lFB
wcfgCtXpku6o8y/lmXCbgfW/Y/pmVUVTg0QZo2aFdtSmFe4dVgi5ykDVkMOo4Jc9
rGxNmDwZiu7TNV+9QAmZwd6M/c87Y/E8G0hKFrBTBupnmS2pfmalUzZNjDpf+eEx
XMEsIjRQDyzgXu/Yfs01pc+BpqgV1ttUhms441Odi1crVCFBDpfFWLmXp2hnLDZZ
THVEE125BYrxy+x6VPo74DG9xbTa1U4O/xt6EiXCbabxRrIwlByNY8VYU9JS72KW
GGCC4dL3bcmffV5IfTWcVS8W5zq1MhberSRaT+F4047z502fJsE4pR8guiEIfXGV
M1MEliIvpN6w9aEPEm9dX1TInZQLvpubZqw7syCao4Fq4S/1jwCC/gzdKa3GiMmg
HpyqABISwBt6kUH6RW/QWNKGm3c+1NT1+XAlvcDNBm4S4FqOAVGJ6XHB+ISmHR3n
B57OLnU/k6R7ekAGN8Cu6SxTKBXJMpCyDdYsHwJhMxpoYcqWm5kC8QGqSvGttH8j
pgCmWKDQ/Ff5RgHsIq7+pVQ+jScejyAGdW7VDPpkSs5b4DHet+YN1EXtrB1a1wWP
h50sZsMRqP5RGunrYaSbF7kpNVUF1R4Jv6RgOx8jw1+Ba1Cf065Ik+xKP3uK/7iG
suh3ddaWUQi86k6BZT8OFWDscJOnAHaWrg4NYtMe9IrOeQ/OhVYsQojhl2Fi2RZy
q2tR3FmPxlQKjenn0DB/Y/Piw7h43ebKmygE92hs8QEkWSAqlFvglXjp97YO1VIj
hu7Q2syl78eFCYN1h/J5bMgKByVtdUK/sHd1oQ8TkqggSVfuX0x2aIfp6dTwiZi7
qiPkiTjF0uowas49FGCfUqPLi2Mc/KG7iRxSmQfYGpjeozYud/KiyKpC42KEX7Mx
vXvVpNct0ZvIJUkK3TUSk/euTpJ4hPx3ww/9m9Y+8sTgS/u6LAwQ19D8Mcv3t0jF
htXF/eK6DpGTwK6I1YokcO0UnZe04z6F65UBux4XsBQbBWYyRYOGd4UvaA42bt2X
Uhwsq00cbXyafK1mvGiG4gQ+b4gEnFlMhh62I9YMJQ/eb3IGKO3R8NEtcOp45IX8
7uHQsdmCQoJ8GdUB1qB/2oQBk8X8oCE3ZiMSRyyNmK4EDBWM/Jl2fLTiG/gS/EDN
qLR7kEVDu39JolFVNaZeCSErs9rnUhh+PeIQ8rPAv8RBtvVsrRKNVNg7ZLDz5Nux
UtQQRIc73QSnEDWg0y68V/pf0bpWSZkB4RKNdRUNRjWr363AkAq3ccqzl4NyadNF
EKzSpXfrZkmDiXdjzwIihKY1bgy4Py9ev9OruHizFxRCRRFMuezxrqs1nG6vdl5d
I3mETiiWdessSr+547B2jHzIm2DR9jqIswG1/HyE7p3Ng1QzJ+zQ18eG3pqeqPDB
vva8r+9q7Bl7omnroFk7LqfmbV6InVO8tp96Lcl4/BYO7PsErlsBrFxcS/jJqdE2
RPwFzj5B6BWPx+utEt9Ksby8mQz/LxI63HL7UsxtFkcFMEjrK+QF4BRMF9lQP3iG
YucLBC1HK582Aq9GnZyOwyzIe3iotV+ZliqsjFvo3P5VSY75fzyFkYGysyIo0QUN
EmttsIUp6rvhZJVpGLIsE2S1X7OYVkTc+Yb+Ac1wmacodO2/wT6IJbVAl/oUOnf1
JsMXtLR/N3X/GjqPZCOWooZ9fsSlHe6+5aesBqClUvazzX+ObxJxulIOTLk1qOwy
07/ARkgml89cBeqCn4VDn8GXwI/bJ5G42UAswhfUApQx811xJdKHLPLnCfD3cioX
UUjDg3bNhI/yh/rUpM3yF4NTLJdV/WeZZNS7wR5RNpYEAur8Cnh5DJ2txh/gD0fn
/yLgmhey0yM8yZ7tEHj3P2FHMRy0a1saJhJxr/HvCp/tGxLeiW1+KjmSOO3hTam9
ivmi/Ub7jwMw9yDVQQnK5YvdN5tf6/Pr4D4iTFb8McRPyKLCRtj7soUm4+NhGY0T
K0LjXnfj84syseEta+DD+FlyIDFKLPiCa+3zuhs9LJ4tNfzDNsTJv68xyT+7EuD5
6jM86jzimgTTDRePqH2A4jpEu6u2oB7H423WXC8Uf0inVGZGYmMwxknacxLntd6e
2kMvj9iLmsa0yXqviwW59ODGV2jeJv9tdpF/QM3vqZpFiSpMARBlKEGWw8Yw0nfZ
ziVi9nePhhlJiPCNBs4iby0mdd3j6DSokn3XMkkIYRSOmRGKqsDHb+2g8OapyDi9
GkkxXuo3RjRXNM/w8DVv+7FlxxOVM1iLW7dxqSsodLc+v9HyKz77HC8aoEOqDcsI
w/nj7goU/ZzDOAjGKAmDa3l39zOtFrnbQuv7YCcYl0BvLiYUT9MAWxxhhkS45ZBv
uPYvRZTd22sgVv1Q5Enpu5JoPQjBKuEKkNFgf+5zAWuG6ntdK/PJiB9pTabx6fz1
gSptp0lxpH4KOHQ0UCfKPbL3ZFOpMu5Gz85ioxo486eAzKjDc1GuqXed0YraiB4d
goW9KZIDxDgbmjmnJXiQltKHY0Wi5ZK2/so6mXgZjdrrSnlTkwhdr6t/HVePZl7M
MdtfNc4mkfOjoaionYnHjqtGGtmC/fD6XvHXRmqYnduksYA3Z/rn5BMw+SaJ1Yck
H7PdYC8d09DcrmOc+c/fbxc8pKTnHOvPBmc0hsH2SkJStFLSMp1PxVuGqSOe0Jri
i2eJopEgyARMrfWBh8AylA3bs2iGiydHgpGk85Nro1W3t+iB8tpj2BrNleOONDv5
K52Of1MWkHpkjjfl6l2fS0RtiO7cX3MQTcTwJNN48aq1y5QI3yeOL7PaiGvG7+Wu
mYjfFLGiW8bMTvdiR5kwI9Dih5afbGyN3mL4yHN00lzgmkN9Rlg+KFoaiDk9UkjU
nYx4WLMsKboo2MNwbxV+jRYjT6CCExpV1R0QIF6N6q6W9aIw8H3kxqLY/oAafrRu
VvyqqNj7gwl7Z++5W2swq/uozyWr+uC3E7ApUPgYR8r/YBGGcs5QhB62XfBbEjoW
t0jkL8j1p7FHRBo/CWZewMAZYGyJ0b2TBSzEeApgE6apKO1PcEy1xsO9q/nllFP/
S5dlFh8lskulsf0F1MjFEahUFB0dmgZrsjMWbf1KkTKtZQpNQQuBqEfzwfEKXS78
Wr+IHskDJHRCrM9pDU63+JU7W+ox8sV7KBwcBA4Jzv//vTQUaP/+n+68Ugjq6H3s
jU8+JnFLT1uxrXdw54lCNj27j6zE3VDwQKSfaQPhy4TD68z6L+t+MBJKsdMi23Aa
cI4gYanmXqUsVqlc89B06fv30a496vmN6aKeayonJKxvm40Xh9z0tfVGhSW5c9tN
L8JYIwITWqcA8skkmSGpYcF0MlcJf4O4yKRXnF2ixi4K9oH7zQGxYMCoE6LOWSEU
tRI8Es9Ax1cOUllYdQluIkjzvV7GZQJkPEUIkcdKEglZn0sSEsFjDkskJI6eXbBp
jUyQoCzN2eQF/VuadYGMpfR195k7CZNFF/WjTpUaJFoHPLb4GOHTda6vN4/M2PCb
U1VRfuWZj+cnzzkp1ZZQAXIQLonYVLRO4Fg7AWhhkXPNG73UWtfMsz4FfAqvONHn
eiXBuGhszHUuazWMLWWrE/QF/9IyBE+8/YA9fWATcK0STCTDt/N3hTxx3mJ9sAib
XvSXlV1ORLnTTIzzfAfmJb1US0+tp26y7N5ROsl/SAbCOO4cnCBaIdKKuDJXjpzE
xIMNflNKnU+Y8ZRhiT53KRNNKd4NRq/1HFMrk15viGwaLFC1If9RAlK4L/fnGDgT
+LjscvZrPOPRmEBmIkvay3JkrpFMHC0uc6rsUJPFWmOcgFDaAnkUXZ/S9p9781sD
xLhF81JVQVGZn3L3WsouPHvpjjhyHOoFL+z8SIz8h5FnoXRQ6XXFAA8m0oIrnAMU
ZDZ6YI4bPr4O6zyl2Jr9UgtGEOshyFRWa6DzGnleEnBq0c1GWewHp2CKi/jKwqPx
STOe0sbjHKQtlcCN5/C78y+qqVzqFBcR1dY56O5eTIzVyvuoYMC9ngc6pN6DZZqL
ESY0XHwbx5VBnzIuAaNIE3GvZ7qXYiofZ7rmn9cVZY8KB4gaO6v6aepwXnm+L0yX
5MnBKi7p2RSXjdjkYdYqe5IJdVXYmv89S/YZGduf+mc2/PTw2HPhXqkV8rrf11y0
lv8YGKw7fbDHkZAwDFVrsbqQpznpv0IUa17LCn8Kt7jKNkOM/54kLx930XkAgErB
z1HxMhq5GGdSLQL/SnLsyvNqBvOcpX8MjZ+IxPpoo6XIG7/CxDXl6lkUufnB0XiK
SHWcs2I/uidd60oPsZsniBv49M9ExzzaFABNfg2rhffWgRSaiKn6RkPYfsf5me3z
MWJrGCPnEVi3yAwQg4oSosZswk6wu90yK8bihv3S7mZsTZXcQ11CH9mMwYIFIIfp
r/lv7CRWqJlGybY3P+jRXhxGtmR+D8aAq6yQlLAxQjNUg2HI5ttAiZErV3LMApYH
xFtemKH06nvpw/hHAnL4R4dbCLMEHJXqLuIxo89Zp41teRa96K3ScY5vXKIbjZjl
n9LZlnI+/PPgNuZr1uaeVZc2chRQAPuruAf3FYHLZvAsokKWdescqVYXzBi1mCo0
kNz/eBe/Kh01uQ8Rb2Z4IgxvMozNSyeiRx1frFUwbeHH12a5FEC0hlYmmUB5LtE5
WsdjRsfV2juJHrX2TEzyPhA3H13CC4WE/jT1yFJePOnMgbNXroNwf7o1988RqlzR
GB19ZU4KzBLkTsrd8r0kPgDxCKlSZ+x+Tatw+2trgYauXxmOJtAbcl+/xRw7Iep9
27KN/VbJAfFKq3+8wjqZ/yGG3gSs7Sowq5XWIRE0TPzLjwVKLNb7CSHFDyCw7YJq
GZS51mKPL1ZJ3CvqihZCuCztwqOCeak4Crl0XMwqxkmA0TOKE848KoHLcYBx1rm6
UxMpQKjZtbS55oN0ocdvsJuIJoqjbTXOsCAp32oxd2iinYo4qar/C4ZX18nZgMiI
H8NdFgNjmZL6kUADszJnSZJUAvDCvbQ/zl9v7LL/GD536hyIwJ03S31Y85oJD4yE
q2lgJheSim8ZGqJAdtNwXqO8yBJ/GBHtoGJ6WPJGpfJQe8HQeiuCqiZF8WOXg0FV
r05RvP+kz88lCoZbynRSCzlJjiY+kO4thVJrQDXRSooGlCrFEWPH3wHfwrHv4Zbw
vtonOaO/U7o64FILRy2iSzJAE7C2c7TKGvzd0I/9ZW0Zx+hzVOsRHDshdD24DL4k
lCt9bFnt6Voz0Rzhr/UMFvak+R9GB2MO8hlo8ZMFwE3WXKYIdvOL3iqKuafTgEoW
WH5MdfZ8g3W6xSgEwxeVE9R5d6WaiKbTvihz9Iev3IA6XSaujVVw1sbDOv/mBGH6
o3JPNxWyWRj0X1MGJZPuhtao8R/7BuBmz0JZNA2fo/WC1kqCecXmR6lpNvt4WrL0
RPUNaW6Rb2wC8aeJk+e5ImfEC3ADpk4PMnSkk3PthTVRFK7xkm8l01vvof3y6t9b
ut9ye0frC1JmkX6ytVEjWUaW1q9CQx5/a7kAETk8QXw7Lda5g33fFSbwWPI0OoBw
zW6JCpuNg4XA3QRk9tQgnYobq1wI8WaSMdywl/vwH8do3XE3CSV5oAiOETXuO67k
c30TuJ8c8txMtcmsotlUNli5PsQi67Kxct0X1HLtSHsBpLYrPDua6k/MvzpPiMA9
vuiThQTUsoFkSlcl+FupCmw8Pa2/G3vgZDjXkqr0Zm0zNYVv5y3m+Ysuh9AbDR++
XAp41kNbLm9FjcKKNp6/BY8cQ0oQysdjULubREEbAacWA3jeRPWHLtZECYjVVNbP
6GnWsz0G8auUUYJ0WvkQAvWGu0T7jNsgtrRKu4C5sZb5nbvBRBRnlJXbsxnmPxdF
SMvIIqWgGallO+uUj11LxRUmf/vCbyyDi6RXYFNezgTWk0EuVYN2ywZNik3j/0ig
ZxfAQqwteG+SG68jINPixlJGeJCklw4BvqZUSnlcyoqKgr//Tjq5Vt+pMsov/rdx
PHBs4gmSUc5zq2x90IPQEdNv4RgyAuIedNCq5202g7IVAwp4bNKrq72nkpNj/586
pMA8mwgA0OpelTyf2xQQjqtxgRE9UZ8PzVqYXNhtG9CdMvyBKT81MO8rHVWbjLoF
IIH6gXtiey7ZiJLbJop+61LqEJZFQPz3pgpH4zxcawlOd3liGZIHcUTvzCY0rDew
xsN/unuRYC5MNLeA7oRt6jPGv0VBF53NwVv1/9dQoXoqCpu8gRjVNWtOweXbIGQI
sXmBPeYjLkR4pCR7F3u5YvdUn2GnH/G8g6Zvk8fq00BG42PMoZS44s0rmE9yGfuB
lxWv/R4gf8cHRtFTHuwDX8TzeDNsW3mYKuLdXjA3X4mNUhDhP7fmKRXMUbH7UgEZ
Tm+3eiw2bsPG0QnlrZv1Lg9LN4+hH1bmflCGmym9pgJ2+AnRsETvTbrPyCcdkWwd
y+vP4krt0PELpOo3UB7PGKvzHx31bByVejQ7qGZBRQyV5lnO+pMI6douYn2kUYCV
45ZCxUD3rtgq1lThb2LQ0cK56Ww2C9VEvUK0qvm7xUpRmV9p5E1KBAcjRYdx2BFp
7iC3Rn9Yf8e9wnF4ABrF/Iju6TSeh0ooW/tRWN+mX1fw0/v4wsmrPFJKCoPhYMhM
rTIpJYYAxxxXXZAJJXePUEhH7wkQZnctVbjW0CktfVQF0JKlEWlGthBU51iimifR
c7Jzf/8shWQVW5LE5XqmJ7HkgqVAPyRupKI3BQYk4OyYDv/bJ3Mvz3GUvmg0lcUf
RK4v2vMoCf/y+/uUPJacRWoOok5tqdOM7JokpZRpjv5+FQzW6D2ZFzTOXPvV5rLz
x6jJRaNXEA06bpDJ3PmlUhqAK05pGEtop2qzkwlEE2K/RTgyGqNl53JFV8KlbIBt
gZAPOX1yUlkglBsBXMnJ9R+ID2WXpWtd9zUwabHk5nloedOiBf89Vng9rZ05B2HW
ViJlXvWGE5MZxX4OKFS5a8y8Qw/OXXeTyo/3zrpocU7h47JSnh9SU2t6gL4OBeBU
yYVyhXK6VGp0VORcfHWrZEl0ia9hONK0YBLaaB0kTSij1cgCple8UGix3Nr6hfAN
4+7swlasKM/Jvho8tx6RaIiFDN+UFuPerAUUR3QMxqzRqXAzdV+UTg7WbpbSflc3
NN58rgAT/2fMGBd1VhW14Ovj35tXETStOX3d4L3cfdNDSXRFasVV4c6CoYnGYRxV
5EjK9L1/gvx3VejIXJhcbTuZcuXmQzRdZTOHW3jNGF5IM9FGDonFhe5Te2DJFul3
/SJhy3TWdOhYGmQwHvqRFrSCC5/gnqMmn99cw4Gu11m8qkX2e8UVKOmZpEOVtJ6N
xIToLfxC37Mxvszomk0An7/bziBzr/Mp7vGIQQu6r4vbvIIqoqJvuZYkosnspnjl
A3NOsbEOV8XzQztEAxVV+uqyCFKh9nWXFFutxkU7qzsvCWsJqWrcwH9wlOYNlVM0
jp/tBArCIwIf6roq/IcugUlxcXbfAQw7xpTXzbNihjjNejotzwIPxxGHlsEBbMCr
AgMnZnzeUw5P6UoYwqvroLWV9SVYDmJZuMSXDisPgOQLhgD+LDiNlngVRsQP4em3
u9SIBjrw6IRJG4THokWSwrOpFCEn/X5Fskr4LCmb9/2Q6J36JIGI38I7/+h81xYw
WjzSwjREkOeiLltkzvZ33v0HZyOdALdQ/CXdQaynUHDnt8cPam6CL45XJFbnHQX7
kGoSaQcNyEiOdHDNOsMVozuldj67kA867iAiHXYhfOF+KZaLDa6qu1r16Kzd2bxa
Jj+TauO6pmBeiZNnbZt3k6BDz07Blcv4Jcxi5hoVWFtSItJQEsG24+56S9wKYEqd
iPQhoD1rfD7ZEBheWoaBmus1rc3MPHHa6+tdL05cigSDXRmP/aJMRIIYTbOZt9gj
o4l2krLLGowntzoWwQapNTTMLUFmrTfDsJGpUsIMgSAFELkyqYi8Ff4SQvn8N7T3
3zb9Cez+/cckMkBWBd8puFusmi1fH6GcZoy6Q+L0gfztkQOllbXTXME+EyR0c++A
Pa2Ep+ZVkmpRZfUocQgOnKth5PCBnURWboNVj2E8Yr9VhavDmltqdpgnN/MndxC1
GhaP77zqiqTlibFroC3fB9avgGHo8+Zj1D21Wqu2d0LY64OTVQu8uiIjUgF2GDPz
dh++SJ3wxbOiariXI7y2RzrsWZY5Ptb/sJwgli0bSlg5w5TNW2gyYR5ev2C7YDeA
/5p8uxYj8Io9sCiDErlx3vSLLfGcipX4QGI5oMca7ZHEvIhXHb/EEqbSdJ95R5o7
IAYFT/9bkOBV1CDWRKTDZHYos3ngaKynwfAYQwrWJdse1AQpR2Ed9p6lqnFdYL7C
6NGrLb7f195utLzld4wKesbBh6X/hIYHknOkGoV7V0HqCllqJ+8FuxA7QAl+23gg
T4US8IFhaIFdmHwZLFmA3hmYPGSDlUDWSz4cah/RtI3ZBmkkZZhZZe9IDXkNLELA
dQOQ9mwX5OB+4W8LrowNa5I07DlcN+YsC2mQZudTXSWkGX+ejMxvpxY7kPhsLrsp
32Smid/EDxnHPJmpYr3Wf5N7RgkoLiQZAYZ7XKZCJwuoAWOfa8emyFjmBTEotWto
a/4ezZzbHDdq1RJP3kfqatRLxrbtfNYnM+5+LLLzyBIpfzgZ+wpG/CBfNSuoNyAM
Lz4HsJBlwWX/Hkt7SZgs4Wz5jxPibsx2JXyXtCsigmQgNTSXJz1T33GOrNnrfG8y
D6FjVx4y41FJpKaFdHCMvsZO/xZdXGElbNJ43FXrGEuNsUc1A03dVljdJsM24Wio
aNn2JwFN4gh1hf3ia46deWqEkUGUIECXtHVEPJ/ygfplqirWGXI3IiZ3maoNLY7l
SKi+BuW3Vt+KV+tNF1kES0P5+9WVP0T+w9OAphl6wM8BYMNt/ipjE6Ty+iciSFH2
n3e7FWB6WKQsXLy480cIeTrxk3VyZiCJIwOY2Wv6LhcAcF4HB8vPRo6vv0LKEpVS
uEaVCIxunQsS3fkAi4XS56VDAHtmpEiENZ7F29OhUUFvRz2XImiFwZtpR/s7B8Jz
p/U1QeaVNCLt8+GzAK2xjBB32bL/JuGiFvWmUkb+ZnhjzEWVZVPEhx3wSJVEPWab
U9z+XTHPp5CwZ2niyh+ZbeqCVfOODO4YqkgwEsAhYl6CtOq6PP3WH2DvK8fz1FA5
v4zyVKJ+bLtBdmIGCbZeMyYS1XSfCjg6uMy6E9bHsbdw2cW3CaVUwF8TtM38C580
WxUvbQmTvc7Cz16e/GFg/OujkCKDPMca+wBKI921onDcbhq3yolXES10K/0ud9LK
7YWY4u9+pSp32ON28RvJFfvwK4mH/tcbVaPAtn+k4etSsEy8tyhEpb5c0ADPtpoL
ZcDyheyFHzK6Y0SlnmhSIKMlC33FxOb63zj2rvtw7RhcSa2uMnAXNo/QvuBkdy4I
3X2wS6YziBHh17vdLCEHV3XvLGk8s4S6YH36z/91rKmTLixaeVOkXclwQRJNwxLp
f6C42ZhXpy19QoFmffkh+rIE+d1V44MUMuzfs2UBbj8MOttSQbv0bCtVaKyUPL2z
BvT0VXIYHZ/HePaDSwIcOKWyBNdlaTRstebQuJzdLtJ+XOkCirDOW4jc2vghk3vK
k2pcUaPUhpMAiXEQcRu01pLe7oybZ75UQD1nRgUhUKjD3oGqSJI5YdgmUB/xKkXe
sv0YtDJoL+3Zxlj79v05xsZFRAZFW4rZyAy/Tpt0ZYI2EJKsenCFnHUoKzT2Ux1x
xolk/tYcWXGenfXTGqDR8dX7G803WTNTM+R2hjsG+e5BBPlz8AVXKz4Tqtzykhl4
F3dtR/p71Eda+yssuLYZ09gMeSeI8uvWExFl7Gxl8BJj32Q/zdPF8GHomGPIvPr6
WGbosH6RfDpGHRAnEpWMZwUx08mWu8x3DoUDAa0xsXUa9YVXmPpAilw4Rb6pGaZq
gdTaR/OhHF1oL8uO/YxmMxeOF7v2UJ8mhrCBMMlIuJhYWKcYdZsC7ZuD2lxn4+2W
mnv4+bgPl9p8F5aH1DqfZ3i8KcA91A8HtPJag2PNFn6CmaXbotsU3jxS+B9Jqae5
lyV7BfvF095qYcUjhHpF9iyoslZO9ke1v13UswOo8eh/s/gqiobFOpdYXK+OHQvu
swWbEl7yBTfpEkW0lqDqiWxe6c7Vl5W51sLR/CDkxyfUu9J+cZLVW2qMu+0RXsm1
Ljvir+vQFL0rzQ8XR2X7BzYTY1DPkz6hky++XP8M3umttMqSdo2C8Gg/JGK83Gv/
lYrd3/nz/9TZNMas6YqTauOrm/+ln9jvdmxIUc1Q7Vjf1IMSyW2IShfJ2jSZHa1D
jnPPsbhdM6Pbo4HhtzJ5HJDDGHchIe3BQr+7VoiN10tOEEuHe3HTfT/4gZc6MfF6
fbYmxCq5WLO5kgGgAH65+1YvgfqYgytGYb9HbABTM0SWTrIHPEYfaPEzD3IhuqBf
/Q/lXaGYXXtLNVAxkcwEnEYxXHi84Manpk1FuLy7ThJ/IwlTnGXTzgM8tD4qezRi
iS4yssfdNQOV/E18838F/F9DEsgvmz1aSmbVLJDnVAjKglfUFpOdSREomzhf8Xk8
nKXMEpi3/1TjCbcu+3+u372FQ6J3fLNKc0mmTS9r1vCE6rOtw6bCjMzASpTm0HgL
2hehXn359vP4T6SaaPdEFOhHMGsdG7E+PKElJ3aJ861tkDNuRY0p8n+hal/qcCTy
eu39k4JC02+lD68bdM+gQ/bB0hV3BirFYm8WC9i54Bex1U0exfGDckPK/yRcSmtr
7jL7kmcwxUPoUwtqRqC3hFHyzgfVgeMsJCAMBbUmYuAHdEVpkAsp1HKGKSQ/7AbJ
Xnn7KvXMJEOD6mooEO+8MrOp10luqBgqUBxbLhVElmfDAh/3ypDiuiQEL4GuzCt+
cqu69dLM0agCV1b4tuPgl2FnZZjmHmlee+whgcaFyCYLiERpvEOw9jZAFum5RSVz
cKvwUmHtMG0oJjZ0gEwR5ZS12UtrEXyiskyyPljuvTS0UHJ+a2QmAPh+NkIXKJxy
ntbrWeqOo2JD4WbQ3f4k6n/JFRG5c/bXFwp6AsFXVx50gcaDYxdzSMLMiYAUy1LR
0rEEWjCZPQyHy+zsE+e8MC2ZdSOqKb8ykHXpASOFQO+kcabH2J/mv4bbqr0g6B/a
VSG9rRX1dTLOvYQsvaD2ZkM76AEDWA6k3oA5L1NjjGwPHK4gPkQtAbhwkrHaGLxF
b23Vp0Vw81SIcz/M1CHHXLtXhJIk5LG9HBeIgDq7KyIo43IFnu7cDPiqxcNO6LaO
r4AucWil6kdl8QqMZvO5c+89zaDxo6L8Ro1KqI5CjJWEzZnXmoYqpcFrQZsTP2OP
tdkWk+cfeVQZ4uuvhhhYYxslsGYJepbRQBQanslExW8p3kzodRmOYMzWuWqv8KkD
f+Avz8TYe1ydxktwyct7iaNg/EOEHOO6Rkfyd0N9K/Sl0aoPthi5GLVXQB67JDPs
HyueRh4dDdCUi03NYufxPSnc7PFInkg/GCbC84wrJONNf/Lqt1Ps+KxMgLQ0qK/p
nwQ2s4mM7GfqajSDgn602ZRgfbBrEj7R3Oc9MzYI7yaPmWCWM0ll3rqfSz+KO3LX
TcPa+1Gg1vwMq8iMb4G/hEOAyfWXFQVBMJrSanpx5qZbrl36MVxuOR6ud+K0REbr
1GjUuiDpbnMPb9offxELIoJew8ZbP2qLrGGDbq9Rdldss39+2DsSFeu8CkpYGEJG
VAm5DlsYkMAK6vNcXHkDZl8ONHA9JDcSaXWqUarEtHDKJuNBXUyoffybAfY9tG4M
wvi9Lx4yDrgQAamT3p/Af5OctXfcIjv+/35lmgic/WwNZC93iLBV4xDsWHgGftIj
E6+MZSAvW6y00VCLk0hXWR6dqVnMJ7nmV0OkA5lY8Prfxb3M86XACH8cqltSjHRt
txC2v/NfbqhmxuQ6QOFUYmUPgunVWsSHXlaCTd4aEmBG3dyP5SvybL2WDMsCHJFx
YmL2wDx3n4RmQlWX72f03i3PrybbPOsnHrdZt19sNHxD0+69L/XuaA0FAxZN6WEw
dgFLL7MR6ee5X6FFAQ351bOj7SCYKv3bC23EZdmR2N9mj3AUZIxPEW1stU1cdPsW
xS1dcNILZqirf63wQATk0dSPxvXVbD33pU0KUbTew2BnmcXIJmVyJlzzhRjYePqP
ycCRmH9JYqkRo53RDtFj5Yu3GAQCL1BkvE0p9wx2GANXItlCmRh9YVkBtJaExCwY
sHr80dd529UsCl3bVkPEqZyYHhVAE1WxhJQe6RUcDM7mLQxvPsi329QJhkuDRI9+
peRs1iSX9z4Po/2dLQyKo+N/BT12L9yxAaUfySiEB6zsoM/cXGldSgsNpel8qop9
Q7KcGOaNp0O0FrD5jXfGJLvnPLdrcBQU82gb9pW6Bh4zKZw1keNQioOuGqILW0d6
NIzglxpXr48ysL2Q0RcyU1AVMwKC/T2051DjZap0MpeUoL5ipFyLJ35YB9STODFS
DX+qQK17hD+0/lyHOLwSu/jJa25TtlZhSHviVV0AZeg00gUblQrc3GcKo2MMnd9h
CbSvfaa4a9FR+oc3no3qqtBqoX0AsVIaGrxsMy2Q8Yw+Ta8+lb+5RvlrYqV8R0EK
DEAm8kdGWqpMxbpN1T2GcDzNsbUhMTcEJ4VgaLs2aHkcqgZCVtKLhbm1qHvgpwDU
jfRkDGH5+YWFQhB7xDZQa5uUVx93BOdEC+XjxWocDDOc/+ZKkdYxdWNOKu9nsj+f
NHWQTVdtd4QS+N1tXAayY3ufEV8l+2FP9Ze4HMWiiIKmDuXdo29kRDN9kOeLn00v
gXMkdLnrwD/sY9NF5nWRnFLeEuts9TC9DzgahjQVBYuGXN1XAqIiHEb0X48BAAw0
0tI3/QV57uuhpnyHQcyeeTPe5YjnLhSWD2HK/AqGQhGM+YNRX59mf3KgaUlxCEj5
8ND9t/CgvAxo2ddW2m8UD/pDT/bFmD6GDMWPwA2+nG5Tgk3TL6fC+jrFqLPG7IFa
J7/jkU+sVe3p4d8z3LNgMPkS1rItvdrrcmbQEO7NunbhuDmIHbC/QAhXWo3gibyy
Mo4sevtjj0PZsa6ks2xmBVtUuivxVeURwQ8/zMI+oraQtrirjnaoLjzyCxcRZb8Y
pa6bxDsrsmrP5qYxhdgpj0Nt9PJE8XOIAPf3fXL6DpRTRpT+MxDPJUewbTU25odk
f7IS1c+owfWwSwgNfXIacqUL9jKgOFZXToIwAYXR91FUdX+OZ+7ouIRZDFOJaC8F
l8CKxpyK9yrRvrRvZ1qB1cZL4IDtfZpWndZ00y53Rf5wHa4/mzePyjj2ASl2DVtw
iMBNCC10R6lzXQ3vVG6O0H72XVMeG05tknLrr3WcGrutJDv3DAa1Pl78UM/eN2Tj
wcOFzWlqdON4bswfZtJ3H10ammDqQAHKdpjVZthog/A0QJnGaGXWnnh9Oa2zTBXu
hdi7VKsBpLRwnpLInhq9w6zRfeaMjK+03oyR2QgdyvhUMn9N9Up8+MrIf0HT6TKJ
2O3tsvsOSQitDJTeVfM8hmBKsWJpgKzRjArTzO5CLp43kHfpND43Fon2ZX6JpL0u
3/azXbpG/zPBSyEvspeoYMFxcz/WFRp/O2nP5yAFhmbskl5ipXcfMqdEG8jKSv2G
S4G6i4tD6IiCvH0+rOfcvPVe7PptucwJbsPDYhzm+oomzzR7SXMfM4Ohrg1VoC0H
88yYHYvJ2KXftoBL0ZcP4aG8esjC4WCoVRN/XCDwxtn4AaaELzRryFN6T+9etzHC
iWO5Ox7q593351dyFoIkvfn9cId+RcJRVz0M8ETwvULOg1MQvy4G71qzxr/SSlGT
1s5uVTHgs3VXuvyMrBgK1lJqN1s4rWnIRgElQewa5ZmRW83LIAW1D4PKx2uX/0Cv
UEpmrov8318pJp/2GlklgVBRWJFL03POimV4PBUHgtmiqY12gocvE6c847BaHHtO
6wjQHVHFt24DoHIfHHmnc5gjp08wJyJPJkQrad6c6pW7tYuN9SYbr3MTMvab9bqU
58LfEU6pIlRm5OYJLCyyV/VEclCoUN/RQNCfVtc5ZrfZKhyrZt89LLb2I+dL4wUz
pSeRGWBfyrQsHJ/HqTENVlAd6U1AfXVot+f1zwcgtB75QBtWoVESaBf2v4+USkCn
TAv869s/uOKlZgXUeni0O/5UylmUOKUZM9HeiYUD4/SJmmt1QBgPW0eknqZqVJSW
70K7FV6faiwTFQNB/pnRDKHlVgbz6/OAd5yaWj2+QcqraHN1oDOFkafcfpXVAYq0
2BoH3JGIDYCWv8j+ND+iIWkWonfIotOZvlktQi7W4XBev9cBWMNoWm9J5uECsaRv
hoycv/ILxEg5qjTsoc+Qn2s712XGKoQfoEnj47lYAoFCaGbCTTeEdKys+wIgchcE
IuzJEXO1JsN8U4hmowYfafC3BcMVQ+KPT8GGWtjexoHh8FcPODlFk7mV0QWjPYDE
//y4cK3Eug2GipdQkLk3O/e6GT7icevlRfWiDeQwxRHQZpOaq3tyI83/7WoL3ZBg
SVCFRhlfhk9Kj+yQqXjUSlkaROkV3PziFYhM1NawDtPtAvxrrHSYPGnOvYqb/LPe
Viy8xio/zzoIfJbWs4VqJ86KQqgfPeO9C4jpGpnVzHxbDr/EFdIpufDU5MxwQtvW
Z3fkdhzG0JjPz01GkRDL5Vx3OHqRWDPs4XE7BgbAClxAPQdNYMJqKQQ/fQHI40bp
qp5EhlUkWqhwdLqRPJLUxEVOk9/R/dw/tqypcex+/i5JOmVmOR/spoSBg5pTPbP/
CrfsPPY1ic8p+/BZlBWhKBv+oLkJoBp6Sq99ghZrGjCYLjApWkwgPMosIynInVo7
7qRxtCD5J+kbHhBbDCukJEjzgR5jjYFfcaTSBwEbnSRfee4DNz3eIQ32l1cRK6ce
1Xo/7dZiMo4HL+yuMrd21S2yIS/pCEfRSHZJwXjds3DZhZ0RBXkv3QIfPjXqljmo
rn+jjkemRknWhxhENsjDOoEl3wfeCCkucDvdJRyjA4193QY7PgcQ2TwnOfSWLQcC
QsKEiFbDLddcRJJ/7LSCLNPRgotOQqOsqrVc4t1FQOxSW8lrvLXIx/DfRnNPJjcl
fkrcwbyeNEK5+9wZxG6U/zhzNkpSdihJmGPj9ZDAu5UCmtBw4M9PA7pTwsiG7Y4P
+vz/UpX8CBh4UQ72DWPmnV6rkhPFSfd4N9/+Jnq+vEdhefX7kFlOja+S79wPOq8M
PaB5RrPiCMr9n5LeVQoKg/2ofYa0lfbAbYTzpWfIutWW0+lviuM7frFqlMprZV2X
vE7SXULIJoLflFcWbUqHGJwmbKW/QgaOo4YlkGxoU5bkwTdUh+Sa/lajj+i1bnC0
fMEi3HENWqtH8jJunNNGIjMqVPr2WDPkJHAA2Q+Vzu0HO5aJJg18BOuofItW36xL
ggdSrmWXPG5/iSJTrWMXI4y4/ejvpAu1scmfqnDpc0Qry4nZhL003GNAF1rdI5Xa
LN4QD0tn9vetTdHznXg3n6eWJgDnL0BKHrEQYuWxtPqBBF27RIaEW4QfUemlbAER
GER9arPfEpnS+7hhskNbVpVp81uoJ60d5tCl4L8SCYkmSurKp6e8euNbVnXDjdd4
DqykukTA0UDxoxBjxtEoo9RlWw7Bzk2ypKmQKbo0q+mHxi6KJm7VRYq/FfvdPvul
AG7OgMIj61C6jlcxeejEN6GlvkbOrGjuxFlbXtkqdBVPsI4W80/q1UReb6SFsDVt
iOSiRVShDtAX0ianReNTx1mfjfW5wI2LI1TNP0a2lcB5iTUKSt2Ri6zVoqrjc90i
TepkaBvp+HjOS8k9y8k+Q77I6gBYFTzdt+xYJqEjni96fC3TuOv/N2pBCGm0sw4x
UkSGZk9VIWW+D4e0U/pi7oQucZuY8vj0AmWnJIqbCO3P0qNwrlnZyFKoj5l6bwmC
OlgxEHCwITmK7LO8tTwIKKC7dHlTzvPwBXpFBgprzqTwdmYE8cg9AvRXZt3inbHn
2jds7FxYGN11SmieaqWs9tR8MWbHah2qVqG4mr+hYAFE/vaW5tgoR+vPsMASgxUg
6oVxUATTsRw2xAZnnFxxZBbKms8znu8EoJXEUHroEnG2cClrYGhPMC/qIIU+sdJG
tq4TUsYfJzhOjFtOfrZgqrdOjwco9G8wmOj1zhDd3hHJ8fEriNjDnlWFGkmAXlih
FL9a+jyehbE+7tw/AaUt9SpJZdY029re/B8DxTr9GwrEkPHpYBIz6VEw/T04AUGx
8i24JblEUKSryz0punCrBFbbhzWGh17vls2hn7555vDYtSfxl375Vd2Jw88fIypu
AxiNxwWNQyLfZDCm6RpgHW8D/siYBHzyG12Zg2dF7uVlB/Otv+5mE+Xz7Cr9ryVZ
Y99Ga5p3bF5VHeRtVw7WuaEBbQQ6aJUFMzgbUrtcwkhQzHzqKyG1Mxd2BAMapcnN
+HPAf+p3Vkz9+WFJ3MiPhQGb/S4HEgc8hJ4kC1xTmstNApUwxErLvalDqj292OKA
dnqFm1lCCxx6alxPE8Y3uboQwt25CMDDEhwIY65QuS+k+Q+DQ9ARRf3MPBeMr+LK
BChrpkuYNZwWc1kTXUqJLGyDUDcSS3Qm2YBxbwXdZOfe1NfChyvA+NuJsIitT8ia
3b6ntwMWJBCGrNW0F8pBoRNXydStcOIiCBoKykjzH/QUpFb/3TCnM1SqAbvPAYhh
/cpmXHH4JfSRjAjig2KLw5Hru1+Wcg7CTR7R63Rx0zg1eEzQI0/ncxw3vI6aJh6z
dOSNMAzwgzQi80kF3OTodb/3SZOh9mauxsRJ5tiN4NR4WIjIEy4+gpP5WgAVgxEN
7cm5dvqgdNrOsfA6rqa5Hb6BEYfFWmpN7/ruqhz4LDH+k5vgFQzT/FKhWFXS5VM0
friwqCXGUKefE34U4Bll5WYG9VpIesgBSrdSWpiK1VqV3ZB8RDKTFxtkdOGH6zYl
f0RvyALfe8f2fCkvh5N1JiMTlV8MPXCwyDO9+3RCyJED8EQoWb3TfvwsRaOijQEf
UCKRsSl6i922kiPnnbf0CFC/FDWZMWH3o3BHuInzMctZKOw74lXAdFozWiXhLcC+
U/2tdChz9oqmhZcCul/0t6xjcm+Uwet4MpAoiNRB7dBZ8ZjbZgx2sWDevba51tYB
lFf7sbBAlU/2pAjnYKjInXYhk2bQ5VPVpcBOxm5i+S/EzBg88MNPgsm2XqkJmWjL
g/alvuNB6uo4yFbK2qiP0I4LNeIGXTt0LC+E52/JPapncY5n/l7CFTSimOrQu0gB
TfTlSRuo3PlQTSBRyYUKrYVL1iwEOSOJRiBUX4/ZVt9x+8kGb6Q1DvY5nI+QQHcl
fZrlHgQdsRPy954h3b3mkJhVxnMvzM7TNC51tuycobabThR9IwywfgLF0q48ldhg
pUCOf6LWLn0AJ3semW3/J3+YTwSwrtc7I8pnlfvGyRB2Z3x0QbzeoD/+/XI060Kp
mw2jp5D/lvEMh03P4zSVNOnT/xWEYct9PyCCmOyCzp2WpsBnfU6sCi8pZIB1t2dt
IWtxpohfMQUXy/WwArmw4I2wMO+Y5KWOu4YI4h337EF+QG25j+E8tTY3e9+daZp2
T3tqVpF67AwDP8EuQBkmgHdTDchGjFnjR/jjFg+v6EbnsvVK/yTHsJEU4uCKzqbk
7NW8g70GaNlmncpb2/OuBps3wslCZy83sT4DBh4nefu12hrlS8hzJ/iQOoec5S44
bgkKrJ8wtFiGGH45JP3tMwKLtCLzvt8YCohiiErf8KUcex8DPYzdCO/CEwkkevkx
fBYOF6Hkq2ToEmUbJ/t7fgzQv53Kro8+dhz9K5y6RtsCUBe7TlOryEYV3ofd3biR
csMiQkeFryagXwfCj3qWHGPcG2qF3wF2+c23otEdfjIwVC7iWAy74QUz+rz47dnu
aMrQkcz7KhGlqZNApWl6r2e3fh/BPrasZz6hJDH/nqOl24e68bOwqnMBX11fDhQb
x2dQdKBCWo+WBdoNv3QU2BFKiCLvO+gk2RQzUpo9JZ5of7bTuwZFSFBwuFS6mR1T
80XL173gv4TC4IXlN+1U5DFO4khK7mIi1M/Vlz0ol2ZbcAbU/TyHXDpFITZgzHjv
vvYJuo4yUVi62iFgJHiI2J/IcznvaxZ7xXj99c+Y5t1r1RZ00XsRF/Sbi4eqSms4
7zs+nEloTPSGWco9nHBI6jz6Uq+XjcA6fNYjUnHH5JZPLFJZYM8ohK0diEvxddVU
1Lh5H8F6uUGxo1NBr5ennWzaT9E9O4WmaQ4rgspnnW2Ou78y4MTwBk9a0TEu57MD
Nt9FpBQVH/IEebgFAVPQGhs7oB/6L1CguOQ5lHdZf4snRdHoWsv2A4GKooj0Znkb
xbT/X3GBZ5nN5cjOhPCSpFUrdEKG341d1HTJjZfz8HPmP5W4+4voW31CP3eB84TD
dtYSsMjQL6itOVPBciBFEvN5MMqZUVssYiR6JRUBKHhcT2o4zaCh32HOUNZAGAaN
2C9GtXReUR843oiPt8zxN+lWvbGBmg+780nqZGht5ZLXC6CZYVM/uWspyPOWqSzq
EO2mk4gRLm17+Dh9pdKvGpDpdqJ/RiCz4VreUWPyezgCqHQ9m78Nd8CIOTxdj8vS
56Pfo6DRoSag76Fls9r+TXVJnvB9bZx3qF0N6Mjiq2WfF1gKVi5mqKd4OzYdE/U6
DuMJ3FF4KM3uOsfq/e/O8MJir2GAbdRMinMsoGphL/LgKCjcGa55zyywEc3x5/EA
iIiOHJlbXPaHsAwfUIJUcP9C7ccQqvQaIkMv7EXL6SQOhuR08nIa2vJpEoeR+6DP
4nOl7y0+VQsdpGaUoFQP3SO6maPw8bUhn9zYPsKye6jty/04EDNSzU1L8n/D5sc1
D60jcvspv+4XtN9XV1Kt8oK3EagQl7aK2an18Eh+VrOGZHH4oGFUcme+cf1k0x92
9NRFNQrt8igUad8w1C0Mo63OvRFRCLnRF46CvU/+uLbp8i3R4Tq4OWXt6NSXbEdm
fHw48KMFiNiimHt8fpiHTJrDs9m1WqYdmxJG1taM6bl4lqyXIsepMIU+OoofVIIa
tpm+nwZHrIL/HK+kXgbtyQdQpUIOAURtpYTD7sFI4Qdr5CzMyW7+c2VBM3j8rLPO
b0kkxNSaoE5IXw+zw9gZQSMDXWMUL5FpDilJzAFT0M9T7XQbzkOs88h+mTglX0UJ
zvZ7OFRr1s0SydxXgo3OlGQOep5IXvRia8y4u307g8Ng38mPrNeknNaY/skUFlWN
k+Fq7dWiyfw8s/o88bMlREBB5S1wN2RQ9BwYgscORy2LGsNeLZ5AjixKiA5JYDpl
LljpGKkO74H4iTILrlo64eJDWPgNnQfDax6AARvLnkqMoUNekzSfxu2/18VjiK6/
4qBsHI1IZncYjEnOzNKFjOv04yNmwc0F8zXNZswjrFzDLM9RbJ/KOeOSiCLKMSOA
QppPg7I2KpUuG5XbdESLsdpfVDbWBidH1/GplUl9NxrZmDIgZeNXOTZ8rRaAfcnj
yePfrIWcRalualGMPprx5QB9FTWoPYrJxX8GxTbqcYd3648tmeZU2qpnOLgBoqkN
e9fLG96MYD/j+oIYPuY9JgIxiu6cbUhEnrgq+GBvhPjJbAGnk8I9vfII8A/vysjA
VVaq20U4gfgjJW8WMIx4xXgI533sk7olz0kV7UUhOw0lJ3SEel+GF7LyAtIs/hVe
HTXromLAmLJIx9wN+jK2DHJ3bQrfmhUg0CExQ0vZ7bh4ELQ/S+OIz6aXNL4jtHdj
bt4WAe5uZkXXEWz473TO+m0Og6nsWL0fIgIgODcTEfK5Q0kO1Dje5LotEKh+hREJ
UE1UUu/u0rlXCvYHFjZBuCFbzsbk/ep2MARQ3XwXPN+DdSE3nRwVM0E7osml6qUE
/UicMfhFntFoU0bleh/qXFZTdRLctOoOY6T1R/Tu/ZSybxzkkWLjjLvixnP9Cs06
CtywI/jNl54Um8FCjR1n6Iqvri/kWAV2miP+XlWlmPmoB0x5XOVHk3EEWMEVMq/v
n1Ik9ti3vCOw/VWLtN0PWALI1o/qGddzHNfNZ6RP/O/VDyusNAYmXzgyR+i5pYmC
J4ehfHYnS8J4SEIwJppnseWRmel4A1bPB/JBEogCL9tsJOUmipF2VGg0N/Qo5Ixa
rfcnvTtSWfq9yuyupOGgnFFgSgaFgiXz244riLFZUggLUDi9EWyv0eQyi8ws3C1Q
5McWXHA0iTRL4w04iIarM3ylQFwQgvzBB1f+bMvivTQfhmC3OQHcMxPXGQgQIlaq
I05hMxhcmb3LuSBwX2BEaYiwyIwA7vGRTvDxNaAgE0oiS5u8sLVtU/R/4n9gAPQh
mEj7oq44iNGVlSTuj256uihRQ+1I4FIQpNBXh0R1h9GdNERk4jbbgWKH9JeYtQia
2g+kbJdITdhtliQ2PvXSEHNzzjOpXE9DmeaRFoELt3wL1O0vEozSwMGwjKTeAOVh
r/ELw9acA36AcPoQMNTCr4Ryr0no/dTnQ1xSGrIiERAPRvhuyg8NwMXk12IfPVfr
FRvIBefUk7nQPkEpYQJLBGwFI1vlUNstzKdj7axiH4ixWJbc3AkwuE9otG9CmZXB
vBi+PRRio5PEg3vAiZHEFGLBoIVurC/4uqNTPBN5DV4x6D2BAkNJlcwe5h88pE7n
BFNzABpK9/OrkvevRlDEUvotz26Jeexo6RYQyRSwrlkwclPGucvSxW62zArc7TUR
1afEwRjoOR/y7sFRB2f7sCLMhWfKpnX8GyA2I9SszgdCGdXfnTHv+fiZL+t+WNok
GFj8KpGxpWNvHr56CL2RX9yVKYhbUyov60JAkkxl0aZAMWZLJkSS6yGBXoYW4ngI
NIcw1Bhb2NqTgW++/t0yCjW7t9XBY9uLG8VTa1JtgNup7vlFhkz3xq9XewGJSejf
gZcbtP1xAl2qgtWXU+RKCXj7F1HlPu2C/1QQOaSsFyWkF4wG9Yqjgx0mLiGAhwa4
royb20gENrcu/Ywe0a1Q2xlNby5LH/PLdy+zlT/uhmvbIjEnO2n+VWhPqx9n/itg
XoLt7izTcaX88nlJwgFIvlllm2/sIu+svVO2J+QT0N5cE4lPsqD0cfRKJEY0/mbz
NntiEMmKXAiMy93wG8D0P5fzopnTOoTbidI2RsjpPOSgPlPiDwWyJa56nVwVP98K
ReuzPVmkX5IfI9LECZaMuKiiE7GeWBflxXWBQ8fefkSfCw9iCxW+H74jwoIh6kPN
Bj5OlOkHgQlGqCyCrdVYAg+W5LHslLjEpchx/TqZikHgaPVGIn0Vzz5cbrZ4s6Jy
6DTfCN+xhm5jRHqgb7UkBs++JLabbWOFNP5VPdC9XzyGoUBZXskAax8gTnHHBOGu
aKoWiXuhcA2p57vnZFIbAuAKrWVfWsNcXWfQ5W25Km85uWUeOz6wG8g8UTQ+9uyp
o9Pczi/5anhxlE51ZdVwWAAnq73RESDI5sKCStdYgLGTWUJT4J6P9Jd6zVpDto5Z
98IIXQtCBN7xiPMdKarO4mgIVTiNJo0wktyHuZTq8ERk9njHgHKU6PD0nKgkCnfD
auZbDk2VNMEI6egNuRiRh9VH3UjZoia4nMBL9/y9Y7yxAk6KZ5hTcnxPy7uBd4ws
UQm5DxRP1lJY0NfuaoPl16UXCogtW1UbQEWJqVd+CbzLplHe0z4cNt2o6saAtLOf
xSLgAQUgpe8bgVo64xyLBywt6ettGmzMcxyg/kxnKd2yVOnAuqxdiHsMp1eAsXFJ
LYmv9MCktSF86nybquFSVP1aslCu2aC02oH2f8OcCbbArPAMehUtQsj0X54i55m5
+ZvV0YKWYrf0pGYoxtKRTLFSp3gjvDjnJBh0c5tXvcizWoJOfSWdTbKoPYI/HeRH
8mZEnbB7HSEQWXlTy5cP70I3r4YDKpiQkah5M3+gdQ0rNvfYhU2BE+ImmWLfIFkf
2y1PiIA3INyr4cxnk9DRoH1lSgZVJJEVsQ+9IW470T23pZk9+yRQY44wPETvUACi
efp4gnUDdtiGm7qoZVBJUbOfclFxU+BaMmtmNnOy58qxWC1Qsi1f1gcIHlVxDhg1
N1SXf4eWO1pMZLdDqYmHQCLUlXmMOClZUBftUhWy52j6dTaKsfdK086qnurvxHP1
JaNrmj/5wvXJpLfKG8lSKrtNtyhrT/ApLat/90xoD1Qn5zm/uZ9dFwDPSzw5K1v9
83Ze20fMwg2kdD3oIXVU5gJ70xzyJQxMavMYwKvSuBcj8Py2UdZtwPCzElIJmZw2
fduK4S3lNEm4S10OosRhEy+XcYYo/+2jWU96dW33M4HmsfDHVPa3Z0nPWYe3DBK/
yQP/INbMt8tDQjgZi/Lsvh8n2G8ILmmQrJ8Wec64VSDHxkz+j5RdELcvCDvXM3sN
vuaFqYbvb3MDz0+w/Hp2XptBDFEYXy5t8iF98BxCISj9eKSb+6DWkYMpcZ+orPcP
D63LUk67CObwSydWIBSNwsvRc1ALaChTJk8NSEGqFnlBv5CG4pY1KHplJzA6Qmp4
fi9sYsQoq/wGEbRBuBu3kRJ6l/FMBZ4uPEeKCb/G8zcLZD5YGrXqNxhdcKxN9gRD
r0dBp5Tbsm/9IY3CuXvF5Aez2054pEagX5kM7SV/H2Dh+mqHsMJ8e+bauk1quY38
2EWZkBXTnFcyu9uZtPi3DLkQMMgAwF6qli7W+9VQlYlMH25n7jxMYCBJ1ZCWLNnQ
6hptgwJaw0h1taUDT/KCyjZZX1Rdbnb8tsR4LwtYqJUndLR5F8r8usTxQOoYpuEk
AaiZDQwbkQBZRh97+jz9bdKgnn3VCKBpkI5eHEqrsJh09Fse+pW45lTWV0GoO0u1
26PIAjYKWsfby3ZTnlSRVDlk98NCoNyvaxDk97hx7Xe9sSe0VE637PJqf5BLTZSC
9ZlqZk9BgnyMZOz9zc7PR5kPEGq7ybYcldfx9MoPfIP1oIm+UhjjBMiZNY/Ms4P4
2138DApMStNlSVVHzpey156hI9aj73hefjyUkTuXP7Doh47zVF2zEccpr8sYJPLI
VD13NpNkLUREHv23uBzk7DLuvw9HftGvA1NWFhAQJdPdxOFaEdGb8OvGwOrA1ikt
h4phYfb9KcRRo8TSdR5XdpN+5kwHO9BPtxUkFjg5aa42bIBpFNqEpwNp4UTPUWd9
oqf/DTN/Nm9YkEWCe7CBP3KDZX+FhZ7mnGnqppwraaCjeaeAASWVtnUiMGTzRNgV
vx5tgAKREF4QtMqQTq9HzjSEWzvG6S44uy5qxccnIr3LXV9kYmVaQA2HIYNSePuz
9rMnFVTdEeS2yT4bWJFI1tDSwItYXpJatYz/cIDbQQt5GXRmLThCSa9Jii/ydIGX
PpZ7blcC7n1vTzwLrwbYnwtLkQOYS+pfyPmAmculAtqnP771QKdLKjvc3boJ+Uuu
+FEQ6qMkAUKI31h3bYVyCpLSS6xFQL/UupOr1Lams9q0sDcOhnpP1LhclY6Fojrc
ilsqvnfitg8iJkZi7cHb4LRndsNwZvMVqVcF15jyfboxNK/sOYfBIg0nw7VYR4pT
mrGPLYPXVHYwxpc/1Huz7zR67OXE5DzdNlVXhevEHPR28njz9WRb/ZAg4gBicyw8
JuGhzWlnjybSzAtzsPR+MLj4M3/R6PSlQhzV+m1UsRZvma+9xOYAZbBc6R4UDJZY
6LZO/yToyE7gQoH0pxiixm2ErSsQ9uwrQu+fYqjrWL2/76fNQZu2xBB6CluHDfCB
EJLi6hjqosuy8NckEbNNERHSfU2OHU7BXWLEGvZRiJHYQOXByCOF3ZdxrU73HVJp
W9tZzWEFUziz0dE6G205+FAmaHi2JsdBTKReEa5hXp8V1OBL6hvEyM1wpJHnZFhD
1G6Io/g3nqFhuMM/Yni5IrrZscgtBzLvqQHayvBesAUCHuzQiETgzwpGPnpjFOjW
VwZ62wtq3EFK9Pm4v+2+5OxwP4fmHPXTfSlI2ZMb0Wt/PbWS6IYyZqimIC/8YR+i
MDllqsJf9HU5kRW3IIwRalwNfY05CkRRuxxPNDS0hBZdcCsv61dq6XygQKrKPTks
rydiTNNI+ser9B749ynv6g+OuN+TtCaIdHFDut530kyE6OBGsRRbM6J1WnfoZC0f
3jeDrKlFV3u4oFLrYMKpA5CyWDyukjGrV//iF/DhZMVdTQxrx3Bw709vd4hpa0wm
nFRko41IphO33woKJob/GpTIMqoHCK/aY169dxn6EKhDo731UvUi8pzDU/6Yl2Aa
vqPWIsLwd1tpYc5wBfLrEcNKo21kGy/NTNfTGyZrMLMa3YvZnDqzS9gAYG+NfcL8
kknbmJ/rmggk8TB0e1aVpZRXXB4JU9Qod6cmh37/H4Sf3ot2/DvEeF/ytVtDlRI5
anUsdvnQifrjoCAfJPAE7vX9wkhYClBXqfzNuxLqVH1+22VosDKFgnuetmcMuwFS
7HenuF8TrCQOlz6Cu7bfzbR7l+1IExqTsV6Z3vZqPeO7Y9hAoO49IDZJx7fXpNid
tTJl9rkqOY14V5YrAD95xN0pvxyh4lQHyGFmEuKGPkgsRSjSVoGxfnqJYCoDCC+b
ruR625yGvcPBzpMhdF0uxsPEqw7OhdpaavXtlixGdFWAdaA8QKw+z0afh+oDS9bC
i/1FLhyRTe0Q16ITNiuHeXRJokQszQCzsSAvth3IyAiHfBryQ1h0YowsOxnnvSYC
mw1H+C88zd94yy7FRawvw2DyMvISNvvYtmKrdvtculO0F5tXx7OtbFpua9xZONEN
4gL5nRTgdMfGFqTRv5O5r7CWHyFuxjEc+gnFTTIsC/g1gvLvNS4AZfzodewOZ+gD
rlrTdQnbvl9co8FtvLiLqSOusnZAQg/2pB5z1/uNpnbzAtRpYKyHQXQ0XoPkiV9C
rLAHUXgTbxGUk3JGM142HbAlLgS8CFEkp3HoZ/HQ25XhGOkQUHg3YDzBuwPtfUrL
WTIzCOTelx6SzrNybUZIfRaqqA6aEkcsxsFP2mj9fyRjbeXBOydMX3fksC1wTWf/
PodoF6XaSDaW6v//Bw8l42N6bSHvvMSk50R3G49L9b98v6t41vePJTT5VuLTmHrN
6tgX/+YVw+oli6v+9OHhjQuISq5fXwUf1sF0vjNTs3ViutcimvtspTxa6JnspQ9G
ypb4aK2vsRa7QR5KXFXhYu2AKVCnT5vJDkkAVajZTMQSaJoMy07nVVoXj7FMmoPT
hmI5YhQmmDzCpq7Y7BK/evaw/3TdmJccO2JWM5Yd5J56LffIw2HcVh0fO3P7i9LE
4MCyk56+vh/w+KW3QKjtEIv6mXF1NYOsy0fm9kMSOeUXbID5762OOSpxCXwGISrE
/LrtMFr40VmKafltYKk28n93wJFobPyWZcnFQmGfItKMg4OYZCzrh8JWlDdJO9Q9
vZz4+iSvCREKOcEL3K8emnYxJJd62RcdIadJPyGb2YF2OB30Oqd5gH1CmP1Bocg+
7kbn1viaRJP9gQnuzq91DiEHS9DqI1t2NGCOEi4Eb1MK55ycCsyCBIoNM6i9ynsl
PQQwZA+eCtshx1URA1BGGV7q+eeEr5AwZKHx6d3WYe3l/U7dGiCb3c5YUS0ao7iE
KmgfvgTiWd4YpBHHcn47IGG6WWErgvbq6yZRGYvCy+wqKR1gP4EOlaqKiDpNBnXS
69L+ZeG8GWy8CR304zmDxXaPsigefr/WJPH2wKo0L0E15eowmACORv9LPvHWqxCw
bZVxVuWvFbkQFNofeu5iZZ1qABGZ12omAd/Mpalj9BoRPGWKWDdWa9iksQZqjySj
H+fBvPAdwMv+3f1hn+lPwWz2FZbgQOm/P513+kRHeLBMfhDveIsADojwYusEvs0K
A7+od6wU5MjzliI+ydV6zgLzR97RkURsTrI+iupayg9lR5d6NSDQF8O6X3sqSr+v
fAbU52g5gl8Pk9RwpXvCwZhtEqdRxWH4osxNtU2iXfJX9/QmU3S1JPEg1N8Y6rUu
42afK5vvB8n2VNC8SIcPW61Ehb66srKEu51+xav3AwtcjdPdWFP3hjaGjjBKe2aZ
NKqyG5RnwlrJWSXOTpWAJHF83F6QU+HoCW8S418H6nbJRteiDFhKPlyZKiD34G1K
spOE9F5xcDbfUy7Iue1+F/AcQiCpDE+X1hi0kDpW3rxWj+NGISvNZRMEUu63YPVz
1Udxkp202gT6vzOG9JDf2ZGKzrwziN0wwlZatVikkTO4CsfV1hL0cW8kpzXcG+Ez
Xiw7h+gwbm3sgi5h5hO6QUZux0lSIJX3EnuORMMYfc0YAEKxArXVHEDwJiLP6l9U
aY94wq4395xLgzU6SwMydqrMBWCs2OtfsjBLbwgGClIuWAn8ILtImzdrEy3t0fbY
BjeluvvGqagZ98I+2Bu5/ydQrLAO7QElsJ0Kzr2LTUTKYzSBaB9VFfFJs6jZXHPs
yn23zjH9M3QXdc5yUsmNWaN+ce5AeOzmykGlhvMsY+kK45NFQlWRUaT4KwJMekCn
0ATkq54mYvzbwb1CJxx5mgPk5t38DxvK33YUvOM8+F++YDi88bLDTJmpSI3WQpL2
9b1DKBUpnaEO23wdRsiwaKEt4ZDjRe/bNvPSTd6ADxYmT56luTLXwpt6Nzscgjwh
HZ7D/7fdoYX4H0tbOwIavIg/PJ86MIsIwoZV38AZzWgEnmb7LeMWXkxrhPJCF6td
acWiupYTJ0L7+bLWAVkQVQZtlAuR8h4dh1qK43HDxyku0vJI7svbzPeA8HvyQ/Fw
cXD8xeRLoxm5syHZxbiQsCPryvu96eIyTf8C4h1AWvFDd3h32jJ5td+sQVI60H0H
itCblEHgkY5pIRpg2hZPCPQXfMSF48rHpLbtRxb/6MZIm7c6F5UBNvvei8ht/ooI
wh9vLX0OWrDUA5lz58MD/zbbKI34gGWiDnT8Z4sdvd98IVa95OifKH1OV3csbY9y
Wi3X1lzT/g1pMn+eMTELB++y0QjbekvRcwa2mqETfF0ZOTCbdfGNz1EcI+vgb5Tj
bJnFcrfSRkQC/rC4qCu0pL86wHbjKKuTeIGkLZUTpkFX7TKaAb19vP+9HWzkgF41
aRtZLa+vVwiP5WnX6h9AeziOqvVpdDsf3llZeprIU4UU76xLUvDPYwLLNQFoI4Kl
1DVmGxF+t8QjeRMvr6uruZU9jj8dPj3bI6/NLurCmrJY1g3pPzEDMKDmMPlJ5rzu
qMWWgmsj4D5B1j/lGN5fImGcu4RViIqqTbMOM5tuhxt8+c7aHblcZXnQ7iZX+w4N
atngcByvCPv8mtz0YdJx5TkzvI+aXdAOafr09iBIjQI2BP51L/JhisLDD3R4++Xw
Yg12AXA8FpeZGpbaWKuBJ+ysXJgYPuSfeAq3F0aarz/htOEVcBGsPzRXeIRtiMPM
zWji/sLFk4EY0xsEBSK6mno9uepdzr3/HCmdGHuw9+ZpDEmuZi2xOUoJ9YDOuQON
ZHpofxlogevE0g/HXsbkCABG6CrdGlByOPvcX7dDT26qvp2iFifFS6vNIdlVSjEz
8ot7tPyuwkxeslXD+ALt7UadpMspQr+/7l5rMvpMZP92kojlkMVUzYVhSNzsn3tt
sruKhSkKqIkgvCYPRlO/tBewl+u+h5fSTzSiBoNGH0tAifG9kZm6ZeMEzxk/vz74
zrSu9CAzlKqfPoCJu42T+euN0U/qI0fKO5ooc7LoOoOwixMCwYFsKBl8gJ9dqXgb
WZTAKol4T1DdimyxSguyXj2RC7WA9i8KfcQanRUrbWVeVfMNuxeCv7L38IzCqSlD
OkdGgToK8PfHy73xeHMPIwf9lMcxFfcdBOd2/uZHPlVeN3ScnoCELM8cJ/W4s6Gk
7ve4skA4rIEp3LBaVm+wutRLUZkedLcZHM1jgAd9Mf6xDeHoYAuw+yve7Zkf3Ax/
dmbYschAMWY9DCW92KwJxbE2t/GMN6WzkHcU1H06bwRYIVRJymJlb78erEmHNdiO
0Xq3uZDWSOgMj8CXWCifpVlC1fPNCUfRcEjo+98GESZoszDEwGHZISaa+zixqI/F
XF8feOY4AXUVzYzpGMvAETWh+gQcAwa1Y5upkGz0NA2Sb7CVVk6ABTHtgkjp5h8z
MBO4pIKNRVLVesDGNOkkt51tLHu5/qGdl8PhuBMQaTMkm0/s4zbhTyABoBVr/Rr6
mPkhjST54tn93Rkxp1JXDZVShvxNmaojK+VVPMNaFC6S86r9/TJFed8E8x/VC5/s
5d1GgT8kFPB/KYvnHsdlnnGpeR3noYRIXBZe4c3exEN2d9l8zmHabX4mha65ylls
EkkpeN35eKYZ5nxCO3w54uHHGtf8aYgNJbmFBHEW+td88nJOBR3dX1s8MF5mLXM8
AGNWKUnAS1Hv0WmJSDDHfxL9PWQEn3E8ono8JKyR4kTHklqTNIxH4HpAooxQ+9Mp
60nVtaxt0XsC9YTjBdeAxCpXlqVwvb/RCAs5v2jsN9GbW9VIgW9tnAeV6arJpqqa
dxOF54RF+O8TqRGxbTk/Y9WRxB/Y+Iyt4Roxupxox5ED160hQPwlsjreoD2bvuOu
AHWYSVjmEgOnI06grDRqC9MHReM4SLQnDi+gzjSjPYsQbEhcr8rMbjwttNrQaJQa
J6RajDJ36gg8PoAaiQIZR86QxaM4KCjCn/+MZlOkGz8h1nJGZIotCF4orYlURaPF
Xui4tpbd2GoufftRInCFSyiVRaFAZNRmKjtxdu4VnnlxHmKL+3w3/rUKGiQoG10m
ZM//u7+OI6Y1QzkODHmlWTrH6+WqThfB7ozPkli01KYqiFLZa9rzIWYaoQhd55X2
lDG3VGm8jZGjcM4W1iOYHMIZXn3XMtuITbsn7pZlpNv83bMhsta4X506YBzZ0rmk
QQWsBoyxpq7c3j3rp/918bOQtkLpLMb3OOMdBGIdy/xI8/0VEouDkcsTd/A0Y22S
aWd4yLTVJvYSgT4oIe18v/wo/03l/XafRGyVNB+uk19jdZWUTnceUOuKznpXp/Rv
NgfqnysidRV91gZxxZtLUD+c3Dc4Kf28QRrF99mDF28mt6rycCkVKAExoz9hKPbl
j4V1npo/Rcrz8deansZwBq15mW5zvWAbeVm1ENsKnWD+MCpZoI+Det0DjB+omAkp
UKBuABsPo48BP4bLrYRjJ3rkM0PxOqKTfM2aLNGGT3PO9wqbyPF+L409WJNdqTLg
BZwnmi5et4S2RcElG+b2qvIr1oi/vxWIANI+KnGRTYKevjSrhheRydGTtb33bAV9
CzfitHEqeAfvPk8nTZ4IcLD3wn7dGDc6RxGpodSk6mHWZ3xuYUL6r0qojlVOCuZX
hL60nx1oWOxl/jVNiiNVfkyJMpoY6ISXLW1gTG4rZLigPAKHaDhU4GIniXxesvPC
Zcv3dCq7XlFA3jbPZlFO+qTl3Ez4EcyqBE5nLqVSB2dM5Nj+kw1CPb5GMx/NHCpL
mfTtmpkBWokavN9NgohgbvS5ItFsy3wu23Jtrq/Xabp74n0IOBHBcB+PUSZCFBJU
FiLDtnYKVf+5x6YUnk5FJqyEDcGj3q67Pxj7Zc5W3l4uhnuIvm+v+J3uEaGnIdD0
JKqCQjhGwk4aP0sjePQMt3B4uspTW8mO53/F60w4Db6mg/DuLyVJJ2mF+6tCTw2U
kaUVuv/nOMVG9NL03DxEvYDXehuaMNEpVAzf2BQfiW0LFmokIZ/Nzt08qochfXic
ArvhJZB+Qhm9PzmYDD786c30RKHpNQBZcufZivlnf87encv7vAnMUrqDMIxj8KcL
1ZD10sDo8Mu0MS25cR3G7l7sv+794QYwGHfYfa2DaevtgHkM7C8EtViU6UXwlNat
CArvNlkP2djguQFFrO/xqiX2VcoSwSoX7czrRI+/U5oEzMaaGARcITyJbj7Y3FxY
78KV+gYv0i+RIz29hy9YuOP67mvrK4PmcrBQrqv0j1H3CPe9Ld45cSZiyLqyx0Dq
tekoQByIB5kq5TaK9Ykbsf4pAp/1ORUk3neFTTAA2i7nR0PfplG6OuwLHU1i266h
7giyhRcBf7n9LOu6YgNusia/GgFpaF4xKaaTM2snbJYCPXilqZhh/5WXt56F7ivP
Y/Ao5B+8jsVa43+IR/YTCqxsBQ0yZaBENsjwHZkdqvEa6hmjUQRyplAs0AuzY9FJ
S/9gbSaZ/vnyfQg9XxcfU95qeriXgsWTmtFUCLt/IHPZyIAAxPuXvUjFK9Bb4d0S
n9cOGVbsGeXJhFcOlXAnxqsV8/MloG8peBYS9vNdizC2MmYo4Fn2Mr12v3qVRRG7
DTNM/2XgHzoJo8cQ1jUduFys4goU07uUi0j7QuN8VBZBnMnAoks5aK2cIrAdzLok
4dAnbwGP23MFSe7RksFuMfYdAPu1D/KmDq34O8tSD9jBupro/WvAc8I7RonebVJc
T4Cu6gAQhWU/2iMtdW8u1b0xtLKde3PweanK7QRyTykPYHnDV1yLQhfonpiVnt/l
W+rNKwwMNLp/K3tmz6n4FJnbjqTOn19xnYbxcWbqC+pSgakDJuqHddMrZitCl5aK
owpMd/lIen/Z86unpDNZE30L/l/4RRaP/Y54uc+QB8ImROH0y3PGgo+ewZDijdh+
XLWlPtnhBCzlPw6Ar6QdmNE0dcHZRfP8ZBO4fFyC618NM0O2ThwXlebtxMR/4bNd
zwfh3tR6o92DMy02U9fFQxd12v6xi5ASIf0hnv2w3/MBt7pUNIk8s6ij2SyJIgM0
5nrFj7XUKKTs0WLUHhQjDPwwT7lVsOUshfG/hMwnWQm322Z1Gx4guBklolmBULMR
e/vV1XGSg6QFzXAD+C1R0KcVpMRZUAXsFxe0ZA2pZvVVEJeWQd/xB/T50YXSlcys
BcWvh3L16yEUbv4honelLvLRSFBSHo8KggXkmBenpamVfVtyKnfhh2f7SEzLa7fE
r4jkHL/eg8Ru84N8SxZo02qW43GsSePY7s0aOkptCk59wtXqWo+TRuhxOPCA9be0
YQcs58/lmcFTYSyYZ9vTHHqDtRprEujhZ6kTuD0XMOsH6l3x5OgB1sTsLF3WQXFM
3LibTLq2CoR5c0+2S523q4yGoFLr1V7zSxOYn7AZiPHX6tUA/5IOrzaBqRErm7tu
sz0LDR7lVNhBtgy6b91tYI8kx7Twu4G3CLefQw0qJbDgBg5mmRaFYnKjl5xuodjU
L7mOLb52d5t0+NtOnhzs29G1r36bG9A1ASfLN7D+15rRAlXtqq8qYCJPRuFs+bnT
j6lto/FL1KgmOgTWUHTa9LGJl3K5GjfaV2sv5krFjX3BY11EAgMpL6OY2WgnZpdF
m1NCm49/4tjI29oY+19u0phmkLoaupbuPe7kErL6UZA/J9k/bBzVCV+OAkTyxRDx
H8BL0RwBk/Un0UqYl0yhmy208Yoe2wwhQLX6EEStBLYgcNq9DYYShPeu189VOR5G
h+rdlJH7YzRPJDXfvFAqVRQK4J9BPsEYKpGknKYxWy/5d6/kd9MmZEdedMyEfHsP
iJyw+pU7XsDq17PcFGq+H+Ti6nrQ3uAgxn1drTSjuWMxZs+J8kRJLw/j+s+gFN57
YUOeCzPEH2RNPXAI0rIIt0OnYiPQ+FuMdZZ9I/VW2+ZZ5cE1EfpP9WXaSj3jv5iW
F4S91A+0C0EoC/us/2cO6nkGXDbtIBc65SbWHTd/0JmUS6dNtnjuQZYV584TB1cY
Ahr6vgRQTyRKVOtnHJX9sd9xKvuzaw76o7gpnpP6G1kLnDOAS/jkkm8t6+QSCAVv
Y9acalzZSk5aMfvm04LS4RdaRaYhuay21Tl+6oHxajXGotoACzxhmPyPNt4dtSQ8
A3cZP5GsuvBbJKTZ5p+GgQ7Je7FSww+TkbFcjove/XuT8PnxFmH0x4YJTa9Opw+J
m+4XpDivDN6Ag+nL6JdUMXMY9bDk+rvDYML6h5IHcvlwwrz/Vp2UbOizbbwZ6+FH
RiWaVuo61QoIBjEtJvgOpl+A1GFAptLgrxEgdvfSWikt+e2TEeclGRVKhpcODBSZ
KoMcIhZkoq6A4V6q/oQnHqQwo2qbi9t3OQjphOKbjlCZ5QuOwNgkdNsIaQYT52tl
435hq6KaRovrwFh1BKaS6KbUy4udymeJG3fKEPk8zzLjc2hQGm5qCNclDfYOcztq
e5rrfd+MKowXcAesYeLiHkrtY9Nilq0AiUTxHRDFq8kxgO9xUvKI2vThukThHJui
xc8Oa0mMMgBiaOr3FHHU4pFqlEfP6TRFQV7WDQjU7waij4HUrrULjced/jc5bXGQ
v5NMw2dPXG3b8Z0IzUNRYyuRNgeWLD4psev8+g7g7eDRQ81aolW3255sgR5gbeH7
FQqNsbg2Iq2j7irktiv2kGqttHjztZW0CdhUg4a0UuYlS3XGbKQBSG+8EXM1qQUc
1toVgZnD7aJs7drBDapW1rb/ExPSoBBqsAbzLQN42Vi0R0/zinncVsy/g3AG8i2T
UN/1WuOpKd5d/kryGFCeZU+kNsMLpegnEOdXU5gI8arP+jbjnK7Kva4qJ6UGa0ck
13bmXPsKGebAtzIufnIctYKaaS4GKRJfgAiD64WNvcnvs0apqRvFQchpjpqY5YAm
ZhWwZe0mbThQErN1S3KMN8ODpUtdGX0qVbyNWeH5ShjfXeSWV6zpwMFbQwmhmqif
svPY+IxJitpA4a4Q5r8qQGEc/aycniLmqruOAMwXOWexirMggZUR7eIlUPmcHuev
ss2E74viLjslGtVJQ03VduZZAcTTjxUR/FaU+e/KQtcBSlDxQMaObwRWQgo8mhNU
+VEmp+nigmljKNhNgSn1iYmn5a5KWqYiD+7T5UyZor/2Drrc84h8WT55HEXZL7kO
tFnS6lSGp3odyg9HPi2D9nr4eJwhkc++PDrqUGGrscFqIr88WIihTFoSPSZ/J0Xt
5rJlVK45mGQmbhGOS7CF1yQseN/SuBK1NyhV2XLaGjPIncnmAFH1CnGSkwLfPE/E
WjlQGl9hrvGypZP3lpxKtpuVA/01oKZ9kevxHmTc6vORsYYoAOIYVP+Sfo6sc2JX
uLDDEWv1A9fePj3McAeewxoZzmsv9v8LbE/+wjTRdmKoxFhpTRTfT/Q436B3Jsa7
vcN/pvKbjbLXYa8UfHD4cVmcVOvmbvsOYpzQ7rhCQlXOHEgfe5v7ERTryyXjjYkG
cwagtDUUobrmVKKMY89Lj5wua4CYeNMxIdBfqvpjNt/BwcHOnQRxDPvQ1nl9tWYR
5wMrchBX3yD9jWQID8MCdaxALi+ip6Ks6x1HEwudiyXyEd83iNj3sLxMBWWf0kfQ
hPXcw9jrsbnxKvomOt0WS3GtPzkuX4FjpePtib8XVXavC6lu/uFFOLu0C1Vy0Qn5
2hnXPijBSCh7DRml1RKpmVVj+XmWuV9KhP3ClL1lXgS6d6apDVKqAzsXmEphjaQP
Gd+H/ZbB8v8TrgsVQ6Wv/BrK/kv6mrXXcLQHL8iFgXCX8GTT3g5O1nkX5GsD+FDk
jl4McOb5kAPZbRUM7rQD/66aP2x9LPcxbotpG10+6DMuhBc1FmaEVWyXYeWaJDpY
70lji2RajqNdKJYBLTyHknL3pRaJTtFX7T634cKWCXV+pns+R9CrwFkRhTltIqVq
69/oNkBqQ0SEvHnAkjcdDPQRcsHZJci8qhpyiBU6kpmdlyqBYQLo+B9fwmU4HYxY
/wIV3uLPgr5XRolc2CoM5mqnQSxFJ1N0jeWNf7Ym3pYARNHewBCPgVIMr1yXLBDg
Y4yPcRGT0Xmco69jek6uJS1xHvbYhT1ea3NWrvqV0pqRRKVw8AOhHJsNCJ110oVB
cJEOv9x4TuMF8isXvHLQ8ZoczO16u+6iTb4lP/knabyNeEaKXPRD3RnOyXGEqSHp
NVyIy9q3YTPq9rssVzA+KreUnbD2/VKsQ7GhO2AVnrQf2yMLW/75RaALvHd0xijE
Qt6MtJ28R40ZwPKEpVel1+RlrUgVlqg/h/4divXODTYlQ20Ct7vMA/kPcHJBSwro
8QJun9iCTXgSVWeQ3XR5h+Www+xHZltZ3Wql1vvqS22SqWTxWRSals2/HpZGNDOa
AYue3Rb81K7q/YFbHQKCHsfzinMBl5ac3AyQqZpIKFK7V66x9JzQ9OF30wwzv0ll
g1pB6O1QC0N/F14kPiCQL7+KQkVlNYmadfAoRf7aA5hEiwhUzLDISELL+EBk+USj
BIHuOf72l7zztskbslyQIvVj2yv06oTvlZ+xKrv7h2g6CU8DyqK+MF5FhyU/Ho1v
eXhCXc51y61uZv2TU/zwsHLRNcTXP9ROxjDjCvqsXHsWEHnhaEzKRPgdza/sAhhD
pO4zYlwErEG+JrKUu8GnrNnefWyZpSyQphyv7XvFCDSRMRb0uVT0JfgCLF6hYiEs
3AvR/MvVro2ZD0Q8yvDMj3KeCh9bejKXhUGYvT8izhAk/H8GGn7pTDtUgo/VNjrn
CAeoCS783lHQJ5C/yuv6F8SlSr8cBRcduL/Tle3S3Q7SypT1AJ4MwSNGZGVEn/rQ
047tzXJorMpG2obZMRm7KL0Rc/fR9gihJajj/NgpJuAGR2QccWFlNFNFjxMlBhZh
orj0cGvUE6xWnxfDqS++RYOlwDNaZePh/HaO657M+orMeLxn8nW/TW1/Jcddzhk0
xjvd+uPfzTTHu9hXWzNC9Fgj6qbPvQREVUvZFszsMyyp8L7GdqSf47vBFNJnuC51
gdJOytwJDjpPkaog3aVuh8LsUZAEGqoIYHUx99fQzvQxqiIVDXEEoHV9YWgsRt0Q
8o/0g12YMQe9506bRMausLjpRz2zcwe2RFihfKc+h/7xx2pXhzxGIBCPC6i+wGbP
ZNMZKLtAR9iFSzIrTiW3K70R0wycMrkzWMuRjdaYMli6lImGCTPN1uPMZ3AFoAP+
4aOEN1q5vrC7XAPrHZ5IPO3Rah8mg8R1wlgVi1+dXEByi802cSx+tH4+CcmIy7xH
fUoRE3B3RGsCAgfU9iIjVIqELyMtBZx1IOdFTZgGh1JL0QI1EhF2uWiFdpMezKnJ
EFuCPnyRxs6bWf1+4cGylpwOGyXfOvDGi7csR1NShs6l8mE7+Aap6QeueTvT0Q3n
Cnzi8h/NYJG6a2MBbkausa2Dy2BY5K78QY9kEOMtRdKA5u7aCfmKtR1E3NfaE+RJ
GHM/c2s5SyVaxD7MjFGCPUl603DMEL2/RsxgJW+CowA6b4WRzxw7FZGwC5GyJ3GO
HcU3sA0iPI1O8MgGyV/6DgZiLPLkPMB6SNJzYgqwwTYt/sqpr/gG7S0MXqF73WhW
CfiDLKTl1kl2LY2KAU9zMRpi0eIxLJ/VNsTJMmmZ/w2MDOm6B7GuvGrmPgc/0A1w
fQZ2s01G5l0V55RzHLgjjzrkGuCFJZgy5liVcHtNWLstvaJjLju5ZsJzrupmCxCE
tYgIheOGGW6rGOGuYV4Ed0bVrIYgd6LqiOWO2B4W+7di/BQUuJqBQX75Bdgdy4Se
bYIgpD4YxpjA6D0QO7Crbgyqagj2o44DEBFsjZveaISQ/jYzL7qFNQDImttNp+/3
vnvo7rNm187wFDGKagj6yB/8Hwxm+suNRCpKdv2kD2peF6/9LiT8F0lJxktdhsQ8
E10+KtjKv8f6vneDOrfFB01KVYgZdaoioEBnO9XyBdTzMd2QeGQn9ZFkXj07KuwG
/XUSGhuUMWesK6zcoXIMA3Myr3dOtc8mgBC/dOL7nXn+kdhUVST+uyX2GAaUrNww
Iv/5iBiUHHCGyLH3aX4/71+JI0pYxy0+I2+QQsCJwGgcONtOa7LcWWHb66O+xfgX
gwGKCYDA4rphSvzHwmEccwQGUI7Am/1snw3cHMMtlEoczEGn4u8KRH3mycCr0DMA
H7eaLrKaDnxXYvlqjlATsfd4WqTBxPUgUHCuKoBbh2NMBqgMujOW2cu+86gVVttB
fXx9lGKX1JLuAe46kih2k6kl0ZaN1CFENh+03nJ2Su98UyEEYYu2/jXSZcALyGup
fkIt5ebNykvRy+s5VGqVz4SYXpRzv8bLBKMS8vzo3LsOyYQePOiecyz9hMqWPm/5
jooFOmzs7PUZM1FxeWT+kGY+qNq/90j0Tjyz5N9SUVxHjNNv8pdyPXrrY3eBkQK2
1CeiUxchL/Ge9QKsF35kr3bnjkiP+etau5olOb4FPglwL1nw1YfGP6JsocPsnupb
BhVv112bb9wXfSNgEWlehCBJX3BvI8uzTtggr8QwGGWUS1XVTdHlzSboowoIr7ZU
6NzBOpq1KqPBBffTYWYv4Kn6ywC8ttYbXafH7YIs67AwRc2hEGY885wdlNseZe4N
jAyw6LC/rMWIveKF47zKl7JoZKw65ujNNLYwR2phkNYQnjV/zBhL7S8Kp4DZ1xGA
/sTf2xk3vkLGNJd49xm7wpCOUzBTRMHZmqYNzcrxmLzJiFYVFNh/zvlUrsIEUnjW
TMOEpBNS7/b3YVNVnSuT9fgzfkwrT608LvzYvE2XqkB/jGWxAvDhOvuICCEKaffp
yMPrDiROqo3l0s2N5dH5C4hd76+0lp4nyR1p3aBdaEhogW/yMMmDqO/YO5kqTC6u
7QoztR+fCaSQD+USjszcAM0zsyLx4tPmYkPzPH+rwSNEJO0d2lAhFvOMz7FCAaiY
hHcIDqF5LpoivX9aTQEN8EtbXlXIPh5kf/UGUAhKTqaSB2vWqMYm5eX+5O7sBZuP
mYrrFOUyni/JvvuQosbccreFYxAoYNnWzGD7rMwhqYaUnDLK/3xE2tpXQxfkV/Pf
by6irfyZZXhG9T41jaGOZwl07z7CpEdi9hopfdFH7awI+H24Q0FgddrYxHnPz1tC
XUrwUfLeP4hcEc30Idc0zqSCWYiAcCAsjYY+TSqmvNivYRO8/09rHLaIhCFsPU0h
eE3Pt6JXmJhCOjQX/Wxc7V4e57IcxKUxZvFmcmkYa3Ark3TA2MiHsbke8adi/UN6
r5sgfqrm95xcx1nwb4Vk6qbJh1beXuD/r5ldSp7m7+/fo58Xvwn/887SVfSY9iSc
0nGBTi58z+oDPHgjwQzhtheSXgr9Q/Y5lJ7TPXhtl41A66dGTQZjizYh7QtTS3CB
54zi3U17aNpbTaJXNVVO0XyxC1y3+HqG5HoLzqMhqnAco9GGnAw+hbUtjxfXHZQi
PYRzLhq3RmCQp+Hrlv3uGNrrITlNp87cMwRqzHIHt4aPI77hsL4aH6QVqqA/HJkw
8QQjR3ZTNF0gv98HuYUKBSajmTYxF0yoiyaBW33hx+9aa8LtJoQS6+3yjvZ/QUWz
7JSwf7V6goYzHeazP+VunpmLNE7EWumdEtGNJQKkWY/R90NIECPGhMo2cGV7feM3
hbKLlF+jzXgSGHxYXlNowVqydKYavo3gVY2nLt0BgJkM4fwUzQtJKatdi7zPWXTn
B//EWcKziYrsdUqBhCIxAuqk/j8JviH6uXUrHr/6vQb2MrY6OOqTi3VYJnvW57Yo
e7dHjEJX13fGoSOt0Hbw2zohGC/v1oJ0H+MG+QA4sfqmqRoKkLyiGL4g7zWO0Uzc
76GX+u2eHFIhq0xZlp5OgBOd6PheCcnjyrNN4Tl/+ot6MMcJk+5TwUzFb9dltOfM
ZXVjbHB2E6TeustQHUpvyS4Cfsr8ssjpinfhkkhAVj2V2j8xxJ9IRRZbNFRxfmgA
Qkp/5WX/HISRxtyIwFt8jv9vsVBrKZ/Bc/B00TzNknHH4vr4bGT/JH+7olRikxtL
yxbvhL+dJg7GdKSytO00quqzivAv4DUjtG+cF20GMt8ct7G5HP94AGVue+K8viw7
NBGTQDQx8WDbXSbNAqvID8HkOAIBjfQJbBIDJXjypTw0joK3r9S7eBdJLFlf5TIt
uXJ1S89AkhgMMulhbAwtk//+L96ayADBwgl6wDtIto/bEdIKLi+Fjac/xuL4gXir
h0tqQikj4NRVXToXGE/tqFkSTznmH5NJOALAKq3DqgEeqR7bWD319ihXbubmwDcj
wT9vCaz+fH3agokVbgRIBaOFe/muGVA4g0Mm28EvT+aIUWDVUaENy/BNRc88FxC4
kC2NH4crpkEDoy3n58Xa9G85jCwZN/L4vPHg/ZY4Cy60gdusysBWTaTnDVPJVjr+
QlUOViSySenmrFgIil90LYm6irFFW/CUVCpOXSiYIIJtIlxlUpTuvr1TkGYdPDuJ
sNvn/w6DsSyg7mkIwVCQwokREybsxLj2O1bNMYrWInJJP+iA7MjtmUoStZGNFovV
CfVDsp30PIoxdSyMFitnRSj08VM8z3NlVQl5EALIo1rvwxVOmW22RMbl+iEzkJnH
q2TEugAMkkNtyg2Dw60w3vrdb/RyyI2ovvKYA2zLK1GE1jQlQi3CanHOrlIlEUZk
EOxLp6PwWhzk1pQw0to1gqaALKhRF/f6knSRcJftk5aUMCs4WK0yAnH4We8juume
0virzDB1nh6nFnZdaVEcKymbASa/jNDUXUm9t41yC1DLNUEF7GK3j3IUAoS+vYol
kPIRdh0quAHNSL++5KVX13KDCpn4FjOJPgE9tHuI6e3ETbqwoaJnmSERSXdZGs3f
hT1vDR6kvTyUysVLRqRAL5TuaQ4Jn3wsp9ApjtlgZyhjIqcey3xFOu7hBAYGx291
lx4f4jFDUe+1KL6WhNkBxjtmm7w4SyeeL8+3T1xNmvIyqQ9W2deQrwMqljL5c1kg
gsppBlnD4pydqPGrkQ+1oYZxEQ69YvA3Qu6jQYrV79d7L7f13IjuGa1KpdOFE1hX
1syLMpiPzssrbTXLqAjZNbma5ikVZ9iJLXpYTc2jC6YB2fy8bs5CZf473EyIcv/u
mN962AWC6EeiVfhzT/d1/77z3t9TB8bC5HXAYOcWl3m07Ju9uqOxjCjzAFPSP844
6B/ggxnYQXZKzMxGPoKMPNgVeNYBKp9j+TZEvXAJH/9JkLzSm4OoZ1y0Szvl9LPs
jGNEqdzkBuuKoGbJasPwyZ7vrGUSJrCtKbAGuwhnQFqe4THC4MbHTsX6bGYQbuci
Z/pybPLpZu+HxzAgPZ1bDSSjgITfa5jHw64vei6dj8WqwOjU3hkk+u/eKcWdMuwp
TsiOP1X4plDOtj6XazoiQYec2mAMoHOmjC4kS9h3nY/AkJyiJs2VusMClFVKe7Og
bYEV+DRS/mMDYyc2ELhtVzey+xWu00GOTV5+ZcIS8kSsc8Kd01sbD3DX9RoI17bS
Yq+VGAF8aVo8zKjrvDcQJdz8gbgcDjxLOLnwiJw7TR63B8GrnqLLm3I7c9tw9FW/
rtEYYAAEqPrGWM7K7PUWFUSv1XlGZ37vkkomXb+JVGxYk1IYHCToGs9o/6XuQ7SU
gpEt1nMrwNW9BYa7qi8VxcPRJ344sX33BejQEhtQyw8HDNCi4aisXHL/GF/XwaLr
2gmzqshZ7rWjLmcrO45pabKJf6qWbMUzYt92ynIP3wugwYmWM93XgmznWpB4S5mG
loW9Zf/9T3/AWWywNkLDikcOOqIv/82JO6EY28Ag8HaRM8jl4wUYuQuLJgmBBTKs
AGal4uVpuwDa7r0qnkXtO0AJcZk/8Rogo+/qYk7GejHbVO8zJcRPWpmWnSGB1xvm
dpcaLhQxJXBAQHKBbZDn+qBifXCz7Db6Ioudwz7w7FCSCpfUpJYXpsvd+kVpqR+Y
XIUwcrnCtf2iTO3/8e3W5G7R69Dj4HxeHXHrs6WaWerbieJu/Mv54ugjJcVlAiwi
u/heHwa0A/5HLKK2VuXAgsbVzAWCKRn2kWrUg2mpGX0QFsKJdxgJrZq5y7D2M3Ws
sMF3Qsj8h/VgACxkOs4tz0xoYN8+YmL8XWt+V6lKbAPV7/5gq0liwwQOen4vDKi2
Tfj/1+GSZfntbyMUz8yVPhTBeqPRqqW6ai+vGGECvRj7fSyYeiG1KA4JpgV2o5lf
ZoYPubhNRdSQDXq5NfBBvNs+fYjnoTzhOpisuFwl9TEN54hwDCLO61JBzebQGH0P
7W3RkqW/hjU/qMmxikQnJ3WBROCGLmk0FkwlR5H4EVgruh/v51kmvZ1gBr66cOg5
MgAEl+r+K2nBHjO0F6iwhooVaZzF+uK/NScKTddWbZjVC6E/pPG0u2vojrOWPDRv
+MRJxgkjAxCXBnhSpiA4fJ7gSXDyHDxcg+TV6nuhdnSdy65pyumJXfwKOzj67quj
r89gVgKmjr0E53nMJG+ZhUdBk5e0V/UUdXsHC/lTLjSQZD9gzPkQrXqcYyp8R80t
T29dfnL+LBO+9eKJWwtioOXqUbLBrkIvqr+C92kyHFgaZd+fQx5oBbvoVYy1CJlh
NhKhTgrsYBZ43R0xYjPxhgNrf52t2a3Q4jldhI7IFYIDDf/KacYwYK/qrhGkC9TY
+X89e1uh+Y7Mssi+XkLJltiwWGwybZRF1tjujpkKtCeWRBiyS7Y4lFNxnOoiV0Kv
KKqTXG1vSuWpwYsINMDDjnMCsRuJ+y+Xu2ChYgFscukdJ450J++ed+5+QE6P+qia
HeMlGVm2bpEDlxcV16UNtTqBtaJgE2on3albWKtPdxu8+30IAAez0ecnhFRHiNYJ
uOF/ghmg2VCYryf7nMbbyr5NaonuQHap5zQQXXDC43dqFkK2LKiwn9yYS75cGQDJ
eTP18c8bljK8uWYj62wCWzQVQN5HSNadP1EqqkPEnCh53Zi4wYbjDQGh+/ZPlhxH
kmc5WQoOXj2UXJHrmiqb146H2fxIUjx6+yrJINOJJhBlcgRTQdcKc4EKHi8WxvBq
TIjgilIcrmL7Il7NizcmdEoeOyB/c/Ej6eNLbqL95P++wVBPQ3Qbr6ouaLAoN60O
pimxw09NFEJgBb5fu+CAKqDJJ42zxeU+8Fx8nssGBNr0fBuw6wdxx2otqzR76dkU
tmatABY2xRhfqiLReTv8wqnPCootLHILFUeTREv1yUoDn/ZDc3dDIN/CmPyYOxRG
C3s4lvp7pImWaqbKfQpkMt0DXiUmyuwOSQYdAEYBbPPKqUiV2uk4Bz/vwnTEEOkk
IF4alj5puITICF4S0/7FHKmCszFAAFVfQBJGQLq9quPMeRnmxSVhv9fZTVht63tg
LWqx+wfB3e5x5/DQwKYHDEAWKz5Zq6U6674LjiUlAsg4YZNgimvQawlo2mzD1Q1X
ZwxjvuNxLmCNsTqTDX0/ZpGHy92HwMVrpvwlzvHM0EVwVl85XaejBlx132AN8XHy
w5KGszLqagzRlzuzI/6mGTAJmz9y1F4sJJk8RwEo8Ieh3w/OgCqjVhjwEGTNobMg
INJztFgo3cDQeox0V56hfC8rZafyjgMbhVAI+CX7aWFJFVvFMqKkf5Qq6IblJuta
/qJdv+K5FddPkjLlY6A8lincZ+OpunmG286BYntOB0MnZgWdPZfv7CFGJKAA9xsa
avHQedHns7XfD+NgVzMbXc6RUvhmgz/tsgDuDDcRrNgO1M2wg11x0CDEfXOcOsRk
pnCtcXZEKavjY+shpWzcufTakxNHwL6/k8V8BWQmMD1GlHOaY7qbWLCbbTy0fHYf
B03I0ddCtdwpzap9bAVuc5FV891rw7sGsjere5Jc3s6BMQEz2XPqlyvF35TS5QT2
Beq2vv2H9L4g2zXSeocazYrya5BZpnH4TIOmvN+Va5OdQa/2R2DdhdYrknQ6fNve
zQyz6jHSwqC2bdFYtUePisJ1dVlce2B42k4TeoH1of1gaENoh/5hWaNYS/zpCJ95
UDIPIKcsMNGWh7pdN+N6k7kuGwkqhefl35m0v9aFh/pR3fEURmqvK1MQoL8foqDm
F/R/q7xrvaKxwd5RrrPUWamIOlN0rFGSNntsYSu5+qKf3DO8fhD/MVprV4+fb6k2
3DkAuLQVMr/d9cyHxwXgxX4Z8eNomdKHel2k4LikkkGRaczKM3llHlfUSueRk9hR
+mS6g8h8bHdkzdN1rL8feGPg1ghDFGkSv4PVx8+ofa9IPUZWp8QXmNMg8Y8T/yci
+nG27qC8nb0Am8izK0FtZNaV+XsdIHOjR/2DALNRSSPFq27cCiX+Q5QCSucO2W1r
yL7POKdJhuu8R0Mr7pk5wigwqRlME6F0YplvpBtq7YEDggGvJkovNxFN8wS7O1/6
Pd4xDSTeFA3/LlOqyEoIC5P/dq7FNTBEv4G5RJzvO8jDDWSiIk0UH5FyJH4hfiRD
8p3tpPeLCtdbPyN+olaitAR7R3aZgnWnBlBO+arv2U7wA7B0kkH5tQFrhzswn6fH
Gnqg7Iv+9HuMUboQpFcpPdUP7+BChUQ0Je6FJLER60QWx3tx6uB5dUOuOMUlM7ny
2n0mcQXTe60tz/3r+iPgZUyMEHCkPQyXdd+A8p9VIPf+bS/ByFE+aD64PsolckhJ
KwPXksiD5CeqsiZBq9uiS9CMGIm8mo00Cbncw34gy5QU9I4kBQ6BGhjvsGwK8EiD
9K1yAg+kg2Fhrh581ME3enHB19NGQMPlm6zAtFlHKUEBwLw56Tw/aes6Ip2J2iLl
I2omD344ca1S2I4qs/KAb65zNA38RP8R7JsQkD2jFEXowjzMK1hf7RAe1a4hBU4b
soepHtNm0XB/Y5IqKNT42mCurHp15+rTKDYeyAHETxujDTjimbed7VTwvaMLlJ6v
gCQbNQ8zN0zmcb/obeQTPGnsOYwdX6tSnXYhKVvDuNMLurVTN0NknpTZl/ZpC2+C
l9xtU+5ZaNoorx4OFxshOShlmkbj8kMCMC1GMX++QifnhXVYaysnmXzQIy+1kTa8
aPdfiJ8ZBtmMm1buKJz/jRC+owgQqplF8nJsG1O29OVPeomJ8Wl2ffYKJRC8S8Sp
Aeim9aM+t4dSJzk/lhHwYXeht9+e9OnsS4npfEzdH+cxZlevyN4T5TTzwRhdO628
JCXGXBLiS7mW7RJYZz1TX5qy2JeO+0hUf1C1IJFe4IgwFAk8glx7JFAVYUNeRn0W
tZ1rX3ZXh5wvKD8vZPJqvtYulkRyTHobNJ2qHRFwFMbDSwUeGIpvJAe01d+wKMo1
busrkJpxwwKuVSOXIzz1mgqy4+2E4ZO2P5zSGRr2w6VoFQN0YYBYJK1ENfzCpmqu
L6ZKlTE9iwnaERJgexsN+tAkQ3wxs3U9/hrB5bsv5L4xYUN1OdxahRa+b372azTr
Aud6ZLuitTuFOnA2X1Q9VzROxtswRdIKrRHzDmnhwjYK61Y8tK3a+OtEKIroEvp3
2T90sGZF6qTNxTx175GHi21SMY1SiHdU83fUye/BlRx18XSJEqjeoPKGsXkGMwcf
3yBH000qxYGFqtxrjKiqabkTpNGveX4RfE19o6DMgJE6KyYerKCqCFDwCAa5LHvC
CpOKGOdAJOEY7xDo+ZqEVQLZgLfmlhqZzpi2kJAlLQsEWU4A6W1NKVU9Cm8cS19j
0aPtuEQloLrKlVPREoAeEMf9zwTynGNBJlM/PM2H66YG+AE0g2058k1JjoglR/+k
UAPMFbiVsQEQl9ii0MKgO73ZnGY0VJ5ZSN177gMeQSBiN9Yl5zMehOPh5+DKz5oE
beOej0jcRCoD7IiPTc18w9Dye4w8uTSrfDS199JdPCF0eGDIMTb4BXWZoxqHnG6x
B0RrICMCZfyYh3R66hyn++lYpIC/VHekdJcPcS265CbZRX1RoLg/oGGGoDvrnmpm
zZTiGXciLvEPNuDU8hXQnHBsjy6XqxFpCSmfV8fHjSdM/TO9Ibx6ko18cnaI+8g2
a905at9CGaZBlNJKbQMrG81ZQd1YiSiWzu6xNxbhOnWml9Yea7oOaxrZJkL0+sxT
zoiAqm/U6apNoAREb5bmBgNqUL+JRuaxHmsX3+SImJl0B8XyQQrxbhQLjqDl7B5i
P75pl5lJv5evvdMJofhC9WaXD22W1CXWRNx8V+D5t9VunYwDNPN7VIjg+AzLcTMI
cQmA50z3PqLNG+E8xJCSKxtEaHsXN5UFJKBMQM2Tct+YlZMREOHitNLiXlA9kbEE
/ocqH3HrnrR7rmsmqsqCcp4+wVhbZJ3jf4B8piirtnN1fFIXwcS0YyH+Xnf8lrt4
HeRymHVK7efoucfnlRPFGfJaVe3W9d+qrulqdVevyoDma3AOpzq5nXwXbHxSeMyF
6+OBdLMt/U+Y1ckzFe3XulSho928CeCJtdewKRtr95A4gY2P/K2BTLCmO8J3stN+
6iIPXS5oFHN91p4Ms8HR71H8f3p80x5dDuEB3/w6MPM9Ro7/SdodxxNlFWMGtT4T
fcbuaXBY+iSFsc28FOmj/c8jcErjkn1EoJm0r3X9yAO6jkER9gUPHpALD/kADXoB
P3x4L2vUIiolbtS0Yhh8ivKplY4SJhT4nF39who3YGHNRLazcCTz8OzrhS/IfoCW
q2+Sf2VTHoiPH3hsyDePOdXp7AtCYWNck0AC4oC/d+eVYZBhEBWvhUBNBcn4MFBc
gA53QeFRI5VinvyvyLL8/nREVhhjpofo/myAJxDf2BaQBTofp/kZ716UuOC7JkVO
8U6P2HHUwerUwW33zykTlSZKBn6x++12k5BiwDXIG5+3nx2C/L1kNCOZn7adKCuC
JqtT0eldThjN26vW28/oscDY+QXsYg0NgiipFABYXb5m572CxGsw2oIVIlDUdFFW
ooJAKpOQgwTAcumpvGYpAlclDiJIFT6roxvp9W5yOeuL7XClY+UGer9M4mxbI3Bg
/PsjBA4x5/4RGByQ5LZYgMCVTM2hx/9aZLFVB3JIzqJI9sEaCXWGaIbWU49hRHEi
PqSgsBD/4SUSLzeDV865nsy64vJ3LXcqveGFzksMsJai23lLo/n0OBBpTo5LyOPe
q0ZL1k7/Je088BVZTAt0w9d2jMGK2Kxay9xvAJrKy+VbAIH5OpMZXNp7QTXSs6Es
MEgIRMM1Vpr6bZ9PqcrQGE+bY742r4j7RfS60wcDEDlhHYTuY4nWNRY8Za7zZuEG
MEQfY4QZy97nEozlyEp+3eOf1jGgZwlTTKwQwRdMgPv1/zYHuheHR6gQHYt/DY4K
Tq5gH1YQyFlesfjHrIW8PcWz9nTbmwJ1LMh8AQVLwAS20YCFCy4W1LqDIqrzhVxt
Peuwt3GxY06XcIs+Thl0STWSZf+p52h/xkDLOuum0TfoZj5YwxUowoFmKSdYnM5J
hxwFb1g6pV1Cgm1y6j30hd5PXesK5r6fIvbIVSsKR6aiZNQhEOSN71M+pHHyCFnT
+etwvXPH9JS5McSXJsQQbU1fnviFFyiiCvwxE87IE4XtybQ6m3BrpGFOelMZ24OQ
EdXDLMvDbVMUVHxA+IrONh5G5A8WiUnSIFZ/+qX0Lnnqf7ZB0gZQ0wayT6UPG6yB
x0GYSf7itwFglmleDih5K+bn71ltxnBTk7VAc47lmCyIThLj4eIGhaz5szex7J/q
BEmBZNF90rd/YDWfTWRSB5j7mqqOCY49DyD8tm7/5SpYXaHEfoFhiiGCPqSHo6rd
QqrL/RpMboMBV86JRXIy/r8qqsrv1P2bABZREGFKDKPIPtyaamWL6j1JZ9GPJlqL
oUIiMh76eb+qLU1RnBNUHMauS9r9YTJRklDmH+uKjuzDxgOZsbyfy29D6gMTX3Ke
/cbET4zbF4h1kb2vcC4GbxQMXUtKja2sBlWoKpR6+gujQZy5A0imrJSG7vVLshpk
ejmzG61RzEiJW2LEyUbe5r0ydTo9FoLX/rgcjtKpUsveXG2pIlGc27UR+cL2+TNC
qHeBgZbOGGXEGV1Bx3QB6TReQW9tHdNIFHPGSDU6wVh1lqODtC74XKAKD1vAxNiI
FVmaIgWQ6yJp7vlUbWHG1L980mKGnMiJSDyQRovdW9+iCMBK+42NYdg0qHWbBm0O
IKqk/VmQUcGuNfiLD93EPcBZObPbLTnApU85xTUV4TxQZKZdi/GK12KPSRsoqdfG
5OH7ub/wXV9DLVYpAF4/tCvfKXDf5Dy9FjpzmFocXsS0lwMP4RFA8gQoxjCj1Qo/
RPzfv19IHbZptC9qcTnMiHIkUAFmrRr6mOd92f2LkKiX2Wll0zyRT/PwHWRuEo7V
QbFyXSiVXLSUjUAOHtLDEfpB6ONcV/HIsdYDaGYQ/B/SlnSooQJ03/92SSxEitOa
fEirD4M7jAK6VeZNZ4VXI6Jzah39dCSxxhiH7EwB84Ro1mg7/k1OqJVFmkcJ5kY2
bjRlT4ZWQZdZpueBhgHgXzpekowRJ3+RxFNwSHvKw+RFAZdS060QM0BeTqx6gvXa
qyAbDKHPqumWOTpcHakCfhhgDWXC9bm64/oG8RYtj0ATwY+oVTjw87ZcEN/WMkaX
xZclhUBKHv4+JKNFwpO+UQnCXWX0WI+thYHpRMY/9b7zGMfVzcMnxGZ/TdNype8i
PbNJz9kYHI3b5a32mjES8ScQ7Bw7lTIzSycVU8bWcoXSlJKFJF2okCQjQcPSknEd
JSX8e7iT/R2RBFUOhkKo8QS2AgEWjkk5bThpOvjdKl/zYB1HWrS3cLVDru1mWbUj
qrdNCFWBaNLumEXsKT4cejoxXDaozfCy3Rs9V3Gmgjvnp9LGUUKlZhacD25nDW5U
R1cfZcuIrLfapLarWdDY+XkQQA4OF3AZA0NCRukoJKVed2hcRNSRyzeq6Q1twgO8
ikv2znPu69peCuRUW+zTZgwyAHKPDb4oCZOXSADxKzrfaRvtsLV8odUriVJ7XsoA
MxE6ufzAk7Fmg8DqJ0YGnlZXjuEmheOOf4mjQNF9fbateISx1jhNYtNMGJQ8n7cx
hvhc/yDNf9q+De1ll6dv1jmjk6KFZMfqHYjlniBaaAVs9qHbUMdLjOkHe9/SrMnG
2ctPZnCeTzAN5+VCtHkH0XW3tZdhmuqqjUUgWWDiroBfVNME0cfi9VTC2ngh1Izn
2Fss6csfZnsqgx+mshywe1cj541/1H+iiMekEXJz4QzBU/0acu08H4V8MO5XjY2+
ZjRQO5u2eqCsKGJgUggqkXK6+e9x6PPR5U0Ahy5+8be1W5xSE4lBEZeuG+ywEhV7
h9Br2Jzree0nuKgHTwaYIOdQH8fvH06nQypT7zYeSlfsCCJnzTiRG3oW7izvzvKf
1BL1TBPQl4SeKG2hbDld97vljRVHqZpO7apCAvcIHAco3h6NDVQCgtHvV2VV80d1
hPDZg6K/m0er0qzoGKR7aoDWu0baKpsVV5A891ceGBh02gDFjcqUNDMkfsq5djyV
dcLsKN9sTY9FygVc4zMnVOSwXHHl2YIvGjsJsyiZfdD2fydKVqDAU1h3in56z0lb
z+x14fLVaf556e4PN76yhl7DsYBpy6Xtc0LC22WBBFKz/tc1W8dvbf5gqW+4FaD/
mWrtWRrwIlMEHWIsQv7s8VBk+4yFCnr495YkWQalcVfwf/QgMchft+0ldF0U7i+s
T6SWCxIu31v17kYw+xQSBSMfmZWnJAYH1eas7lkhhNJFxb4qaDUiy5rMguhzB7mx
403KjZXknD9twKyjTjw2NXMoS8iKsqdgZJkRPw6U0ii7rc1RGFBRk3/r6Llab0dq
KUXMTA88S+fNWEco61DoVuGdNuz2oaciLD6xyXWTUXxszVLU80LSsNMU3GO6uazl
aV5Pvlt9SRSjXcfBb7f9W1p5FYj4QMvZJfp1NIVeoOZ3aAaxU+qRgCuAgQCajLvf
Q1s0f1LXFIhZ62U8e1nK5YACABsiw56s/lPyTO+0ZCA7oRRD36B9W7CZ/RdTJOv9
wnr5d9AXlAHF4ORhMabaBcvJNzIIqQdF2uI9HjxQNTwi6jhclxcBdPTsPlwxq80Y
zn0gY2i0uKYElpL19786NoHNz6/RKoJ6BSImI5ytfaWnRh0s/xofw5j6rH93kot2
8RXlbEM9OBH09zZYoElyf+qh9Q0H0K0wagmxg3eBPilbcfs38+C9pUcKKQLv7z7j
tW7QTL5Wjh+M2BFPd0jcNkKYk9nYyErdLQxeIddt6l5KrverWSEZphL1jQswlVLF
p9lEofrh34vOU08lTzjGRuh5KuSuj5I37c3Ko+XiBqtaHTocxqLgte+g2+4VU2wQ
akghJQtNTbhXiNxXc0RqzRcYdjMoAb7LEmOvINEcHRk1dCQ4TFKTRwtu+0JEtvQe
bQw3VyPIARn+Vg3oMlBE6ZoGTfhwN1nwGaEu+r1s4O8LQZAsZN0UIOamLTTsWR4T
K7tDu9FBgA7Tl3/Mzn6wbfhILq09HRJSWC32p+WDll+BB1ylKKLyO7yQSKujJpVP
QPTLZpg5P/Qtwo1wb4UuISbIdCeQt9Ixh32LP690YhWcDq/vnkimIJTBi1rwh6ne
hpSNeAtnDzRQC8wBB/AtdzWBOW15riIT5c2kc7OcT1pSv3i6d+hFauxSczXdspPB
/KLoHi7cCZkl8gelPqPv3SyFIUTsBxBuFfT5diU2bHDPU1O9dCpCbJzWwlk+2BPT
sDCPJY31WLVihL1qtKdbsxqrmJfas0G7KFyC83KA/BHrTtUuUIpVophVojpzzSWY
L4koU81Nu+j2i9wU8KY6GB6RdqPHX1UaJY7FJcchD5DiCQehtbDLRGbY5MfSO9uQ
WxCAYssIeF3MQTePSOhEqBffHpwcWMdeMUSZijT3m1NwKo6mc91roGuoGSrrtUNb
sVijTunH4FNBoZIimAG0ouxQ0bNT2aZaury/1MCqmfsGFk09pxGMNvSONF87Mpog
9J4ZwliWa8nm5MbfcmsFbWKGHvvBKlHJJri+8lB3++zQnMLk8nYoY1SIzFSdBnyr
ljHqzP5TcOHoWIn5brvtbdKoSjzL5G4665OOmbgqlciL7/6xk/etBMfzJ3ak+2da
cnRzTXKG3EsyGj9yKT+hqkfKOQh/TBfWCb+8QNQM+rAlPPgQOEZi0Soh4JRzIDlU
VI1THjGj+SYlktV5IICsG3Nv9L1sOtlmXCbyxHfsN5DIN/+LRX9S7lvqMh39v/fo
K+bOn8ZbpoQm3UKRI+zaUzox/m+e9lqG1TWScIfdTmGYWn91c6yst34O1dfZ/T36
H94Z9DQa7jLzWGDkQXnt9u2s9PZ18Bc8bZAsqIO2bLkPhlnUnAjP4YevpXK6mjM4
uugNDO6NNdPtbJm+gHnWv4dvhZyN/sZD30oPUcHZ6EMo3B/3jawwI2Tu0CRFYt+i
4dcQ2nByGld3C+H6I5ruk6zGEL+GmeXz6R6izWLbv90WFENUlaBiBzpmmNO6DYNF
sNyVcM6MYvigCFM/sFCapAiMa7M0VwRpOxvC7vkFOHnrT/BmQuRrqVReMEkmVe2u
LccCgtiQ74tN7NkSgjnmUFgK8UmG5SCXgl1PqC4evTFkJ0PD4xLVw+HkpImAPiL/
3Uzi2W6rGSYjaL1Elyjeb3KtbeFLokszeQwd7PtiqvYz9ghg5ZHZm92GZsQn2evQ
rQquBv76v0Rs8w7++oi+vlbzEircerL4I5nh5wfr9MyXfUtMZo3ExbnGJO12Y1ab
vrlYnS3H9Uu9Y8hCvPR/4Zk76VftpEzZafjLXs6x1D+Xc+QxhW1IMGzlVx4L8F3M
VajEiXYLr2VpAyolqWgPEqBueteQd72PBGxMNeK9hvAK0KZMGgNiVlw7DpwC/yvj
JqAnQi8EWB+RMduZvF1mAGFm7U4wtjbvduJwh1eYOtPpSnv2BkqJ29OXhZXBpDQ/
XOWMYACXbP5lKnaj4q8Xr7oCSbDioBNxH3q/Xlzni89QR+MjLawEp0n15ET+8DUb
TwLyOSnTceuiJz0Kdwa2yabbpvG6qxRADTG4dkRE7UXSu2RKebU6f94Yszv8he8A
I7r7Kag0n1Hqm53RFwAyh/8HMjaXGDWm719uLk63rfBlVmqbw4UxXt2yw2P/FnnL
io09pgKdZ6HqdsLqaMsx221uYphkXmeP9P9n0Tkhb/Ewks2vtaZkND/rh7G/ghpE
eCPPAnaae7dyWFgN/TdVPqzxWaJj/Z3dN/uvYHY4NUV1M+eQKFKcF2wc54TciMRy
85cFtl0sKojFk6036AftykfOrY2+0ZgpwPxhxtTMOxkgS8C2jOCUh7TgCRvaC/xW
ZFEPz8zzAUCQzbSfxETx/Gxy6qYcvZ+NfQ675qvCdf3BzHAMiiR+aOg+QRGSli1i
6B/rNk42VTQxtbNcGiK7FBzPTDhm5bkN5/TYHDyErmeS/p/4NdIvJGXFSp6V/Xvd
giBBP7bRDF9jm1fDXRjv4J7h5BBUx16Qp/ySMSMiRWkNJZuCADaP+UBP57tN4QCb
/X+/XsI3ky7gq0yzWgqSh0teYuGuFfokCtduCW9iGFSioaF1ZkQ82gpTsuWUeqbX
h2wqi7BXA0jcYuKncAoElod0ZQPuP2qor9kai/59x/4VNmwaraTQERzFz8H4/Qe4
G+E80RC5oS9JJ/a+Z2Cjm+fScln4H3AI6DFYgb8GU3dqyM82+vdPoIg5a1uQFv4b
Ynn6ySc5oNAIsn59E7THUONKv+duS5vH4fKZm4sJmPbLTehX9NqeI0ue2SOaJfzk
EeV0zKOC603dyCAkt7A0tmRAEG4nsSusQJx//V2hfIfb2iYuTQYOU4DDZRC7kStd
gzJwLiZOQPdjUkYRm4etHCI3cOS1H988z3wNna0kcRrxPKzrBVADMdkzCxyYcW9Q
o1394nHFns1xVVyKhuKtfMuJ3EN5rtzyXU6x5P0pxl2VfABvAUcXjaJ+HSEQU1Ew
n7NHVVLQ3haJneQXT6vSxHTl4c+bvQvnoUBr4WTuCzaLF6uQwHdGYV2/TVoY6rhm
5GvhG7DlpOi3i07xsRXcOL3WEFBxCjOGhNYYSBIW7D7YF7c3a75cE+WFUX3SOpFw
XTroHim6H+uB38EZO8pCmV/sRnrnJjWoPrhwRNpnFozvjKnjb8d6PuollGPFHs0L
L47RNViKA5vV7R6cqvvWAkoMpP7J6fd7ROYG2yq5v1/sWo880nZn86ItKCW2WGyn
7MqC6wx/uV0rN3MkIQA4SYDn0aC8vVWMJ9fxQkIMuRt2GVlnFIcg7qQQctTEGU1N
tEIMNhnbgvZoJPvzSNZ7fyV5jVApxPj+td+9tvHAk2/7YSpx0Jj+YUh0drxxTTML
flagyjDd1rd6K5rwE9kFTNQcUgYZwPmAMCOKs36YkaTXbg+8goEX3+vzdQfAD5qt
M0ZHsbhR/tKoANfIX2NO8vkrQkqyYJY5QpPsXgM0vWMI3qe1sDUB1DsCy+fpyIsF
B8NuXiFVz44zrK7oFZJ0NW6P+Kt/TPWtmTGPo1lPgFVa147XW3OLuHYm4gWp7sIu
QntOWrXHKyKI6AzfYIWRyF3TRtynN9r6jYuypBX9+rL+DMGVzngaCdud2Wo1w8RZ
kaTYEw4kO31HafBhGi66K4g86ifvy2/j0FMkmPu7RJtb79pnFA36X/qbuv1kuABJ
ACF5wwiFp7RQtMwmVOMTcHS8+DeCat7ZNeOXWkSlaM/P+T4P+EaFveJ3dwzT4A8v
cxJCsyIuGySJMEtdURnI10cyChRFzybxQLrTZKh5D5tmFA7kJkgNUnnHLOdJln1u
F3khGXQqU1AyNQwJpnt0mewfbTTQVfh81Px7VfxVmx1zryX2YCtbJhLsj+V+IjEO
NPThzTIXbYB5vTYt/r4FG9YS5eRqsnP0r9kBunb1WKN9f+vrHwZ1CdivDol0SiSo
vO63qwGeZC+CiH1Xo/L8ONOuMpbqvalfHKxZglEW9nA7rTF9qhdTjz1RzqwtbreU
q+7IuPYTN/beftPf8+uXPZFJVAFc1wRooKGiAeVkwaOi8H0KTBjZD4Vvp9twhmhE
bRaZVDpP5qvVnNzzjVd1zBxytM8BdgOabfhKeewdzLZ8gutnVJkRqmzG6GLI5uaR
A3z6z0KN+K51/EePuj0A0lY82ycdO4BTgDpvwZC9RiRHnI2PbDMsp+764Qhl48bJ
iEhiw4UXervnUnAXVQ2OR/2bZLBPfcGeNmJfqwUSaX3kyXNH+drDAHMYhbs029LL
n7BE5Otwkk3c1rQ/zfzuFTSH6qwUakPdK2C3Avwvd8hEySUMsbBV/anx6lXWUC+d
LH4xm/5GqjJCLU1uVlroyjKlEQT/2AeLwBBpQH1jqIXtZVjCKohv8N6LXPzRqVqg
OdBXDKUoe8Ih2YKNsNxhQciKkLOHwyCs/tsOJP5HycYsoCBMZ1s7xhl7Y2CBpmOi
7z7sH1fIi/3YkJI3q/dVdcyeaEYiz65I8oX5hxfspfaAD6gMhqysWB67SjnDnF6m
yILGgtvMbdvxnfvgmRGwX3Mmd4Vzfy3g3QpSFiovhILg6qYH8mp/Fdy7GyrUyRwj
2Ss+OZfgtN6M2emOzBY0djtSYoKATG0vJae6ZhSSHk8yjN695YGRUev3L07peQMs
7RrpEyMZCO/r2DJGP+pDia1qVyFiPC9uxJRwS0is8QFdVQ/OFZA3mIkMxPk5dcJM
fOzNbUiWLIqqH0VAMzJD6jvtQiFri4kPhIei+XTmEQZ9luHayeRlBTVTY/2uQBf9
Qa43EnSZ+QrWZWlqOI9gC2/AveP8rjND2T38EOFHeE7G6HG6ISOCgnsi62KLetFb
1Qln3xEoidENjhAtCAwLnpPhQARb1qGDpewzeF05X6YHouZWJDU7D5CNMB5+R+dB
XtfWk6Xrv8QQpeuFktSUw1oSI4dqpKEowpuYNjlzsMyw68fGbBf2/B4NXkj4iE72
wYY7IJBfZLXFuq3jkakh/z+fo9Gon/6NTQTvrCoaK53cbhy/lJDvGgb+biiXlFYO
M0z9d8gaTiUCy1vGBBjb9BUH99ajNjOPlbdR2qaA/AqaAkPrfSJC2AQkJBCGS7Dq
b9xUUC7c18Sc1eOUGD7x3PZc5IdgBM2du3zQRzG7Hmc2qgPwT+f91jD+AaEz9mgD
ox8QH8jIq07vG+uQYH0Cb/iEw6C5+VvuLPTwP+UmsqvHncuM8Hk5owq3aUpkj1zF
Ma9F6HyN6ACf1PM3HRjTjMMzoWPsS72szZcNudBGTfmqx5POzQwMJfV+TKHI9jqz
6TN/nI58dF+7xYdA3gvJ3p4awApBkZIFTswRELTEmiAsIe/Zt8W6soAg8y/5Zmtb
pEoUweS8bm7wQUt2HLZeJgQKMJOzEslYQ8N8FSAdtl8MqMrOlCHzJ16akvIT38hp
NTFx002viRnZilevPTTByXGIy2M5JFhPUGBBOMXVSzD3VC+YcEtUaR1w018F/VVQ
tEvH3Iy9eKhuEneu7i2rS5QALuPQGfKC9JgNe/ubgk1HVW3Ar5YyUlCy+CHasG6N
rremlBAmvqkdVNPYrkOCdp6WzFwMAa5oKVkDe0W9vK8spmMNGB0EapoNrSQw/i3C
6Tg2LPuAsQO83g4PQqLrej2SrBocJ36B+ME3tCHP9lG9XkmLttM3RveZiZDjO2Ln
nn0BcSBVS2KiNkz2snqhLb8+7pzco+1RastEXwN0Jqh/s3Tm7O4bc1rDUmkwcyDm
8G+4KfcdSnTW7VK1cOCwQM+yG/4mRoGXHQ0oR1DmIc4+HPtjb7DOzRmf4LsxSAzl
eYi6ocZvV8uyBGRxxqmJ0nQi5om/EChtvw5vpBoAohz04hQCp5rOveddlt8+xQYw
48zYBLyMF+pH5lyVh3dR/DoSDzE90NB+ziaTZXaX4PpxQW3r+xUYTSYh99pPjkXS
sQu3uJW3jjl8hpCYLTCLVon0kPc7UOpj0IWsAXSFeHmSVSj5R52siVmbxHQ5JPgj
cxl+z/pHrd33pzAxCME3RS/LuHptu8BZJU4NBuJGgA4iKYr+MClSIo9ZsOPh00qG
TWY00HiFt6RAOj+/PB01hcbzdD+4E+N3H7ioRdGQJvOZq/s0cThXavDYV4AzXpZJ
+AJUCvTeiy0NtizKmfVijmteB0ZkgCxaEy0CpMDymKNXaLkdLSMUMPrWHl00T4MJ
7Gg/R2FkkF/kdyA2y1xj6+Lc4acocs68KnNktk/Np0nbmgPiWYmGmWdYzq8fnFom
vSSWU/xF4Xj6toUFKLIZPZWQyhEZkYETjdfSpUEe6vQ/f7JrIImIqrEi7z4Ohw/7
3hoTo8m5ld+pvSyJBm6fx54HDWarIx2m8XMToZaqJlSO7Mve9HQjcZtmRe7HQGhB
PcS9afuym+yEhvEjvgdr4DmrHP2RaeLgcPZWM1lY6vGQz6IAPvNC+l2/rUTkTLhb
j3qBlHG6lj85zfKmOAnW17ySZRS/wdlT26dnW7H/Od/0I/L/cFbRDXIBhuFx/aDZ
JxBN0CwClBUTfWz2UkFR6SVxNyfM8KdJM1Ondj0RPfAQoC6EO3occtrVP20px3TH
lVYhUvweQbVt8klT9+g5yCBOygHnlrIDtLH6N3fn2IanQu0VEmwC/iVCK8I4JvlQ
8yaWaHnBbZrjhAdfJExE+ARHI/9b1EApOhxjf4+iLBsuM+t63MoFgDuOcix5/Qlm
PnFDnXoK3JqkbQ5LhmmzdGYig5i6jzU59E3AM2xsZZZggg1FpgAzcHRp+Xgav0bc
3z4t3+UmVsCEMtRlHM57KZRoTY/b6YVwguy/Fw9JD1Gi4W5iJ4pKROGmLhkTRllX
cpanfTuymuk3kph7xP2OVioixbq7d6CmgM5tDs9cyRqJNVHd7k5UjeUNAYsMCBQO
hlHpzyrOhQRZNEyzO+QXeA5XrPmOj9fKpHJIi7xVxALmKlQWD3AO1Y9/2t1SCefj
zW7x0aenw36gfP4W4eH6eM1N/Q256f5phH2KiJKF2ogPxHU6lHAmeeKLvHoDM9FG
OXDhskrwLdWQOrdhoXyC0KKSePx3b5ChtsgGIxihvmtPSKdnAKeHrMdCL6eqy/3n
CC8o9WMhTPvfYP2f8p7GKij28mEovGeW+ZQlUG8kfMJRrshkRe33m6xsaAfNB4Dg
22Iwk60sfmcjpozBU9UTqP0qhwiWcP6FGww9/s3I2oPEjnHgNHzcJCy3uUe/ROs4
wF8GuTmQVd5h6hvUSLO4iWhwGmGgzUVaHLeKOHJ+HOlbR4eQoTu4SiWrDctomk9X
pL/0IJ0inT3gG1ZH9T0NFprAcp2rJMnkLnG1lAp1tGhixgAH5QRjeK2ue4yRCDIn
39PGxJQ7AlhjptU6QDzYt82BBJVSclp89HQXExZ2NirtP99+nxfU+5+H1baREcdG
qB70NfUU0hsTjr9EL3Ue6HlyxQhU96MpBHPqOxVJSDWn8LHQFf9hUIlYofzEXibh
um5ij1x6V4lik+LBbEzpZLdFov/SJU/Zyfq5IHM/9TkxJJeWxpSKA/OMG4zP3aj/
t8ku6lPIdPHA6OgjFyrkDySmIKOJpgUWirG1fZdeAP8z0a/fUnv3MicO+Eu7c9Br
5Z1oV+hdfJFerDdihQ9Pb7od6rfYyBOFpBMmclC2SsQ0LpCe7NaNLh+Sgcc2zcVW
o3mS6Dqd+rA9mR0amz58Ou1d9X2+P9wmSr0RvrPLKVceh76euKvTDE1hj4Duep5M
avtUQ20FPLrkR4cTZvwx79ZxxB5TQZg4PAasdfoic2gV1GSXbfmr8lPSJ1JE+tGt
fUISzoCsjXFdyqxgD3VstGfkAb5MpmdHqX4YjaBJ1/OL+RDLgYPmaQTthBRWLvNo
7/L7YhMgOaPV+BuG4R7stRaWtQqh97KH+P1J6C7/Xzsl4M8koLHVuQztlGzuAb5X
PvFXuJ+uee21yU2PX8aeQizbhwyjjZX4hwCWhR7QXNJbOsx8gaMi0StuA1MxXui5
jfV/qAjhv+Ruvq+wXmT0feqU6FgEHYwGApXbe9XuJyCPYdVJKXvl15v3K7Gwk8yo
sar6BX03TTRC1RiZ/5ZSwaS87Fh1vSq8dgZeGGvwYPWoWd7JaJXVL0zybOgoIlFj
4EokIjCUJNOr0udmMe6P1XjC/4cPVBEtBIO0CfbweHhmYpeGYtQyCgY9qPXOITte
1m/uMGEzMUlywXg1OfXzV5oFBCyMjBHNnM4KagrSbfc9aHwxH88AkyIseI1Uh8t+
M3gZ+qGqYXdztYqcS5lrnhpLI3xScAQhvOQ74e6X5UXj2xi6OBJ/1qm+0eJBciSQ
5MSKPJ2eYWmSlCcLISXlarY8ECO62hbrlAfDlCdj9ciFykeZ7Ba4T8/+mtiOqFu7
Afd39dopjjr9tuOrKvPh+Bnq3o9a/GSKBSXjEs9UF77lbD++wNYpBAjy1AQydteg
nzNB8KZIk2QWFOU0lzJMhoufwXa5UA5q0qilBAN6MO7dLi3skanz6nsF1FhB6Hur
dtoW7q2swqoeSbFJnbOYVqE5Q4RAJ20sK2EHL18CJkQlMGeeuxIHp6tslsGA18Ex
6Bq0aKu1kpZDAa7zXh/vrQEmOxxqxwnL+TiXVAGFnCfn8BznXpkCCl2IzO6rFEhG
M5EJHY00/5/SLM7vV/Kj3Lbc/3OE3zgt2t2phQsBmxPgic5y7I7qZOD/ZW1drpDn
glYBAiPOU5UdIVel4IOXpLNVtNZeZ7AU6mwkeiVmHPRbEpYoKDxO9LqX7GvUNN3Y
6orl8V8IuAL/XvIbRTt8kIMoZCT7b7nP2VzzP+qSYFog3VncdvBYcXnY9SGKhySk
O/XZoxuKlX/+KzeKYR+B61hfXBRvcQN6VRVUKHWN9S59uLowlLoZ/nw8yXZFUGvk
GJ+cvQWCch5Ivnd5ESzam/dMQnaCyk00N11FqkwhxqTxIoddQG41yfJbBj9Z8GIr
Zqosp5FcO7dydtMDdsbWUsyMfVWJywz/poiheTz8o1ztEDZqwYke8ElJWJMwZ8ns
SIsPC82ipqaFuegAy7T0OIXBuGcrIyE8r2MelJBftccyQ5gZsU0NMLKqHuKctG6B
sUvtph1TlutiL62e8Z7zyuUIoQL3D88eNqsHasHtBJD67LyB7UOduhcATvQQVABu
qukAVfqoxHelmAdbLBk5mj+API5dap0onttzawP6nKUdPNLQoq4/lu40pV5hj3x1
J/ap1r0x4xMHXz6+sgmM31BdVHOFZpf5xI4BmOpxUHEFFf3ufSnr7dZN6bGbXfTE
S5EWQZvQcckCdP5H6bF/EaLCnxtaOkT/e2n6Rf2dxyAafFrgifrTthrcz5r/Pqo4
pYe4X1BpJ91vZpKrEFKJW01KkWn0JqvlSHxrbWN6o1H3ZQkS0aqKfVVGiL/upe0S
o1A+4MRd1hRSpOlujQmlni/x+c42LZUPPF95og6lDeAjOdet8aBYBPBzUDtgyBSW
a6NMbjp1+wU599uFWiD4JT2TuP+ls79xcOpTeZ1boGqPTnXf9C44C5ZIqJ5in/v7
rf+QRbcKQ0BpdWwSo8p5AkBtkLB7ousyZxMcGPb5ik8gXOpgNF4MuDGcKcOTWGay
NlpCSQ0OiQo5rQEPnvE1qatFiOzss21kI3KMPBq+ELFF+Wn2rzW4NkblTboJ7FVr
o4AyTXX43hJbTGNUl0HqIMXDTURG0aK7VlEZsqAD4bEeLwEXIoq4U308TfuyHx0F
Ca2nokeF7lrbF7RZyvJjGopEtfvriXxgv5o1kzgOdtE2Cp/fAJ5Qo0EJyK2PpAer
Bxb/QjPg5m/xF+rbzDhcAG237afJbCRkkHCJ4n/5xr8szKZtpcSkbKSLBriBUDxa
Uw+UxAvTMeAPK++ErqbMlzrVqIVZIW2gxLcvUV2WVZ/iPeuoEDxmO2QmVYDXVu7A
X1VHWd565MDWzE6dVyZimv3/47aB6PeTpxtQXEiY1pbajiu7GP5mL9lUshRlFM2q
kmcdQe7lyZ03bLbCGD4gcnJUw02ZOtoIgp/A4DI4AcwRxtIa6z5bNi1o58QNZwTi
AZ3NrpHc3fmh1TSMCOQiArTk3qP7nOcyKeG6OZrGI6LRnkMBnr/cLPlO1FU7YAUn
6TRZeNC1x5RhrbQ7pbZsIKN0gr7UIxfjLoX0JGV21D9nY9U3FYA8NDWS5A/GSkuO
HRnhi9Jw5M96BZViLVFapD+9U1GCuXWycu5JyEVDEVZnmaP81b9dfDR3SVSVfFAu
D8hPFyDIuKcoWEebLWkFNjZufaOl6sYc2rLZdFc2ifDrY1qKNNlzV7vNQmTCqV+B
BZzFGL0c/V1p/MoippqdzRnm17vt5xgOSr6SsMpQub98qqaeLBzIgDLG5mm94IS3
X6ScEfEUsUFS2DLen3RFrcIMMNuh/0T2hR4dfkPZII4QMo+zYaXkmWjQS75weC+H
u+aahTAdRJ8vprnnoDZlX9mq7ny+bZUNeKhKnvlSoua+ad1fqLGkpmtBiVycHBy9
Pems91md6PjIO22iU23autMY/UDBjLZpw1KPIeJGyZJSlY4IQC9kGwSob7Ck3gtn
2c2PenI080DvFjbGdUNEbBQQWsOtW9PbLYDtmykaHG/3SIQmmUDplMlhQWyYBhUX
1PHNBud8BA1k2VbF9GFZmOK2m189UHfp0D2VkxhQo5SAS8xwmhDUWOwTJFwyGFEh
7T8JTedBUP+w8FEN2E9UuNb+BQuIf5XmsQy5sh7CSxKf1irRr3XQf2AyMoa/cxkY
jw8B17KBcfUxZ1oOHfYHKXEfWydn5cd2TLqJZuQYd17/MbgeTBa18R8W0Lz1IhYI
cQD8u6kZ248p2ZGfUkM3fq07puQg9k8/ulMaZlK9RPEUyUgVj1BVtnGrI3MiVeMH
rLh67UYeka0oEn9AlbrbYhrwJhs0lTfRFpj1G9lg1h6ExrXhQOiJBJCcUmhNJehJ
bOL3ay37fxigrjzS46Z1qlIfBF3ioTyG24YUk0X6CFxT03t+dabvoOTQwkfr4Vpg
sShS4Omzb624GfBW48qp+yqAc1kLF7C1YjUJPF7TFf3Bl7P7Gbsk40zdB/kxaGx8
XVeERG6Qui3N6JI+WERhSv84og0uVkZr+vaVt8gCikF0rkdkqXBcrjvbBPv8OQ05
+jWGqMR3brkaPS62FnHo8kOzHkmKX9Na29pbVAOwkncXM5v1jwPCUfZPd5Ra1o/r
It6FCU/OuI3LGEEMYu94SkKBPuWkQJXHmOQEIx88hdRlPYAwW6UtSxBdv1vmooEz
n/xWrJ5OPZVzooGPu8vgYgrYs8fJ90iRpBRUMa538TgCk4X/bH9aJbrZCGTPGWbl
bfphZELNDuJoGfGft976dfDavBaHaW6wT1gUOQF34QsRDT4N/1vNoSG7RSXdLcPV
lJU9bHZnYXn8dc9LJlVL4fBe0hSjJbxp4oeGgkBsIhD8lMe/oAlc3kAOWXX/BO26
a/eLwL2EcNecUzQ/D4YxeyfoiRAeIsffVSZzjgmDEvBTGmCZILwGD3tTIL50s50U
e83yIGybLmecwHEKRs/4gSsf1U3UTINyOCTsP6Tr2v3KQigWje8DvSKQlcDv8L0f
9AjxEYrbC0hCFZG3o/9lGGrfu5B3S0WK9oXIdDYAUHAf8N28TNT7e2kDmoEHkHk2
YaKmApO0rRbvjMtrPvP9zXKr5vJRVHvJTdDieYDQ9qa0mNjTBK/dGiUizOCL37BJ
+Fl+xd+N6n8P+s77ISxrYQYaWYnnOoZElj/mDK7kVWp+2qSC/CwmPMVbdyG5ooAT
s+5GYKbJV5VTuN88k8BGigLmVlEUwAs+DGoKR4MDjys1ccT6Enk9FrhYwvQio+dT
NtqZB9RWIBDdXSwzXCdowpzf+FMYK+WjOObNrOiHCP0Kzci0BqUcvAB42jG31eYA
EywyPt7c3Q5vega5mf826N3RANiq60Ff42oka8I4Yinb4e0mTZ0JHv/CSIYEopYc
WnJkk2xy9X/iSfjkhEEptZ10YtfyCLkOSa6dWD8cedNTyRDSjS+48ZZ7pjL/pR9P
XEM/qbokWujvqZLRuzZREbzBZWSgrCNhVfREKAoj5pdx/JJ5mZ60PjfOPyH9LAic
EBd9iIiG9paANE7gta4RkfTUUrr/oK71QSz+fvFJQjfOc3ZHKCYrtcP3vzPdlb86
X1sPDiHlhEO4/HIqhVns17ZxHCOEpVTZtWG5ZeEiUJTlYVE57KhV7dkr7FP4851P
HFmJq2cEeNnPZBc56sH8/PlagP3tsluO0sRLqjTQBhCDDrMCkw/38zpOdeCkLben
oGm9jRZobVKDlXhJTJTWsRxA1Yt6+7SoZBqt8DtayqxjAI43C7pDhKVVMXM4Y+1r
CAVsLidl2PRm1KG+6C+7RVaVySCLU19N95v1sq7mlLWoguhbPYUuYO6yLnQ5UgjS
7rTl9BDaCKTVndP33yURd4MD+WA0WTkS8tvuMVC1O5uO+xGr0xlWRESriEZ7CfSD
9Y7Dwp3JRZU3IvCtUlh2rv2Z+EgT0FDYRuT4svscGXwmUEDVKBqGjx9l9jCjaEFK
edbdx1BWXfARxRcIXiByQ3nqcfEPTsmdrbp1RkuhnUvDpw/PJL00Dx6UdbVxPkZ2
qvHWIIUKXHI5J0jycuz4vxFQowsjtVX1iV5njlG7usMqFcFd8I0Myx5ChUi8jgOz
6Nme/9RI/XczI+ojjthnt6MO20GpaqXbx+6OZIonvfRF1PyPOgGU8gSR4q8PoFv4
3lqAyQjMPWM89tOoENFXuiMAo7jHxE19XfDRgs78fH43MP6PZcWU3u1lf6eHCU5X
EQDpfaG3/vnEfye/dbyMfwZ/0dEBylYBmNq67mLcU6Imi66UGaCMu9q4IaqFmX45
rpPLcUQuZMcqIr4sl0beLRBj4//OzKlNcG0B/gR8wJwI2WFAmCHsLXBwriH3tSLy
6mehpbCq4MS/TYhNHqPRZ+BYf94Hq0D5gX2gqdk+X3UsmFM5PBYcBbZsyLBePkC5
Fkdd+vvNNn6pzp9bMfW11Yw3tYJUYdLTlt0uxKFqvJ/OLxD1Sm4pVzQYXw9nPvD0
s1Eka2iR0QgZCZJ8HOnYF9DmCjoXwFilc39xM8YaHQVA+QMnTTt0mjLb8SHCNWID
OMR4FFiNqINlB7+3iQHvtx6HH7o+Mb13ewLiGD/r1zzjdiw/2+X09qUr+ZWlIRLC
EIksXH+rm9qGPjmRhLROpcEJ6Qm/s0Hd4QT65KRSXWwQzctDokyXZIwWVfeaO/kT
Bf9gvi1eYioEHQTPQMJ3znwvl3vVVGJMzpcD+6NFL3r1jKEoO4lnjQI4qCYd5lh0
agczM1hVtcWWc8cqszyKLLKH0wM8H4DpkMWtNFWZaff1EKSgGqxqPL4ezXJFjwl3
7jR59eRusLC8w//mVgl70URG2vxbPvKK+E5DphKrMtAJTMqFLOMxdrO+BeQjpCir
WqG4PQeNKZYXLDJzQpnPSzAPFfzctc6dLa0PLW3F8NyuGQDQriiPGIH2akvHBq86
twkNEIayoH1qxMPu4gOyXmmo1ZsY2IBif+tPNqbVKx+22XYqQpI3w7p1lHK4fVzf
zXXC1XJLMYNwx4Dn3EC1/LdstDoDFcOMGdapwIkxiYZQ4+u3bnKIQP3sF6TsMZRn
qWAzEkPE4YiNoQ+4OfPWhI3ChSpql05maTbeuMwVK8UWem0JPMBzvXjcTEtizGjs
OB4P+3c6VtMZNbxMO+Q5G+bWVzGgDklJWYhRqUkxFi/QSg97MyiiR4f8Vzh57/Xr
kxWQRa6leAjhpun7m0RuQtUILrFaEeMXloCf0tIgPMPAtafC5vJD1DDMx/AX1JDc
RhoM78OAWgvin1RiZ9WzHFq8QWU9VZY9O/hhUw89BwmzWz8J6BppGuw6U39EtXca
fa6E7lIxlGEbSYOgrFzrUW9qnTmMYcIKboTSv7tVwW3FGLI6ei2TeWuPaAq2AlRM
1rKzB0U7XJWiQH9etckjvVw52JfPPAerVBMz96fJIG2poYatyD7o0MgTZTouhf8V
pWG5oKxzm+hbl3LxruamAXX06qVTwSjWKs01wiclNdTROW1fH8JwFmIsLxY8yFp7
uEyWrMTB3cl46B2YT0NpHhCeF+/z3jErYbqJA2dV1+7TLlbayqAEURWiTwg6B4Wm
ykRnRx3oWVdd5nAGbNnTYJWNZ/1z6NG+/wn/6W44ubAZY4mu0jeA+xdyB2QwVCcy
lAbSgKVDu4H3fetsYKyl9PRFS2bhyPOZ4wK1bpXOpavHfgxl9H6rLI8ACnXp/8NW
36nyk5JZbCCVV0WGQPben7P9YAwZ60ZmSe39UR0LaS9j2URRHMEYEPxn54xcO6yO
Z2I1UIGnM/46/NZBu/ySm/eDAxuo8kzxuLKQ2vZzjxdliujE2APUQHQYYTd8LkuF
qhuKCtBPRQdUna37Jr0lsySCoXjr271/7x29rnbNXG2cC7/ZLbfXeWQgQZHxNA53
VKYE5ILAgS1RffxykrSAY4+NRIMw6cPT/lRWVS7n7/LbRGTq6/4Rdiy3n/VKyWeK
6+WS1aueXJiL1NV8/AWCRfz6kEH7Yo3s0pfRh1B4MT94SedqTdn+l+WlxbWnVFOv
J1DReDwaI7KyFwf7a6svD9if6QSZXlkWFcEpRt6r4zy4gLV2OWVehf2mBGFhXBza
okAeFpfon0e7PelX28VBNhhUVFJ4K83VgmHc9qYlJ1TBVAuw0gJQv29ZKwfEtXfb
/miRnEwcOFccsT0m82uujIylAqz9qj/fdNA3rxz6MLYc0t5yusv3p/QqbBEXgIyr
o9VXCVh0MJE0NNeyB3OD3+zGbd0XPPQw+XgblzXU+sp/VATh6RVMN6FXkkKhoToE
tDGvWKuSrKNLhPkWZFJbYHbGEH24OcT+9EfQ+Pq3l6MgdaIdrR9WHQOxaq5m3b32
+4ORhyOjvp+4X4J67Apbzn8+4x+gS6OJYBQ+kYOQdy0eP8uHlDSrgw4i0qtNhdxT
v2vVbg4URp2WxJ/MWqb1V02Ia3YEn0+MsVqtuj9HAYVP3LEc47wAiv1u/rTcFC0Z
DAoPHeJtKOrw2lj6d1pP570HBZF46tDVJELvPPYsvPPoJaPwPmPCUDCCoyicNjyi
DdNBBWaQxKgVFgsW2hU2D+mvFlMo/QRFV80tca27Xmc9PB6r6mNBR2LQNpZd1rBU
0JyuKv/RHGwvYvOB8yEmRT5sv1lxa+EVJEVcWG+kWK9JOdv4hTA3aOA1JCtR6eYn
YVjOQHWgQU3uD0t9jr54NisSVqWhK4NCgwEf4blWBsot2GzAwOVT0xaX3FY5hcW7
qNqLCmt6YOf1CcttQPnaBEVITS43FX3mwl3lhiD2c+10hWjFdE3YcW4dSxZejQ0j
INk433RDrh+kW7hvl4XBNuZ+uxlH/FlrFU/MuK86j1snh7dYKZUIHjekwIfz73xX
EdjzcpG/aCd/LfoHHeuvhhUV6/7Q3+c+H0q06LnPAJra3Eb9O0CW5rf+Aqe+qp6i
HSH37iLM5324p43jLFIOorGJ1r9UEN/oDjrv9C0KqW2bejEIjiHiOWSuSA9IA4m7
Pvz4H+MLPwmjfrLyyjGIbawXJmw8kBD6F03Wv5vzpBnFLX5FV6pjiqTZ30pbQUS8
902FJ7aWrev7S8mUZB13gPt7fXt3TBUdOp8lowIXXg3iUj3lk03H4AHL7cs3kv/J
fDb5uZ5TxNlCkLZcr8fZud/hrlVou8xvqcAjzqJMB6Ze9qYj+Hs/W3lX8WSVDf4e
EdClCYRsFDLiR28YBdgrBbH5W3vMvWfvsZpAY0BberAsE3LgOZSi5P9JfcnSNGYG
wB0XrQGUcT/I4J+mrwNqdVUgIU0ceD0TBtJzcIFpym1+Q/exMFP9beEIBbZRpxS1
hgU85bGL1CTa8DGTIVnc98f1zJpNK5wVVDa8l2vhi1+3Y4bwTc/5I/zrjFAqCIXF
L8i1iC+uVsFIayG5AC1tW9TYski+X1Qt/eYQo9N2JE6Bt518byU8jMIAVlypo9h0
gt9uH/mCFEFEWHlOuq9oIzcrQOcRw3EXC/ic9Op8xR47N8r4oCJ4lRfqZ5dMu/WF
5T0weTQD05O4XlGcD71egHZiNkkJx8bIibEfoP1FghojKTSQgInI9VE6eiHEJQKq
0ywGBSXfOyruu2pXSuzTPFqkqxnhHPIvOeumi9xAwNnXK2ywCQ5YqvDblZCgEzWj
nTVtlcJtLyksfg7xqvXEm25pT4dsxWw318O21lkH0nExix/dIpRUAuutjNOtBs0B
3lALggNrDQpwHaJTv/BJ1TLNzxzD1ik4e/MhXXRRtNVEfPVKab5XXEU4NFvuLvhh
x7bezieJM9ikRlE5k4MClaiuAmCxR7s8MQwqi1rff9My3Cv4PZRb66j+czReohYl
VayHZP+EX5Z0RuWyvsngQGel2jnGT/aHfjRxy/aM70qda41ixJI1NZSXZm3ASfpQ
rq8FPDQxviYRNA5t7vw9UvzheqN5LUL0rWoPGoZArR1G1vvMQGKJzudAGQqbTb+j
Khec23TIR07h3byMn2MEobi+P7CGl9Fy9W0tPLBfDFJY/af5ewLEqsQBGwwqa6Go
ZaweXygS+sGZ46Ioncgr5XoinPFXsIZcEbycxvCAZRkwuOXF2aLyP9cdZinBQFz+
0CPt8XLunqIT2B7NF0V4dI8Fku7FgI2M+MmEUg4X+6tuix6yhYpr+LfCI1mJFsae
UcXU17rprN3gtNXNDkTU1LXRUUqHLOvLrZ97V9v3AFV5ieg6JCLWphEMGYzrR0xO
PQVn+k5xbWDZHupLRinYUMdYg6YawU9zixi+c/LPZR7F71iU8oB2oVdir65k1WQN
ihsUgLGUtdfZTC2zOskLI1/m6VE2F6ZHK5FKzZEL6UgM4tFp6HDbT4SLvJTvwCZe
eVfd33nELmS7YRMu9z5KRB49/0s2Pmd2iWgcXRzjp72qMhfQq1euka6ZzIDW6OAr
ZjFU8dELamQ776uS4Q2DSYOByLhvUSbpnHa4PdYQ1YbwOyszEQodAG/zuDOlv6lB
fT2uSnakJkwAvoOecQfPrENNXNQD2q5upps4i0Xeh+F4ug9RxmTsXs40SBMed2QY
8BuTypEQkH0G3dVZHfPDwaJAluabPwEhDengCLyiChG5GhdOrL17YyIwg+ZMEz1O
0xDtZy2iP9/5q66VZrlm6ODsrZFEd1/6PP930ndHo4nJcfuT/bMvZSCUR1wsKsZJ
yMUo+/Jqu3/d0Xse1/YYrPSjP3XtHhOFeqmSxhCad1swlSvmPo5Ajci/xxx+cRjI
48sd6Q4GcDgG4nn4L8RawfWj8Tn2uIue4zHtV9DzrYObJG05NpZF4fEm6jD2fNuG
wnVyAbURGe9pLGztGOS8ajw5AhH7aAa2NOoFJt/mVXlyFiykOqLQAQJ1PkkbI6iE
u+bJix2Qyyml/dt4sYTtn61EhfEYmMXh/zM03TakOWaOfwjnoPd23jSwh0eXHWuX
NDXTetY1o9l4swnFAsnIn6XkqJq8YRDQvgN4gp9ZTDxcQ2SA3pyOGul6SiESCZmi
1BoWZwFHjGNTfBYvj3XrOsBYrqPkkThVUyZxzFRmIuSE5x782QnMjB/tv3kqVEEa
ZRXos8pPC5+V1FFnJDtm1cm4FrQgUAwlKq5npo5Rtdh9txJb6MmkdY52YNOPsEJL
rvMFmPZGTpAQxmrA9fVSqmiaXWV4B1CMs7bqPRDrJcN7FQOEqEYwMR5aCFOBl+c1
ldqONT56ZSbg4bB1k5FEo7m2769/toKCIMCIPKDL805Fzca/CNXGuQRENyUFZ0hP
G8cz72Ryu+jFHj8ljIGXecSkVD7pM3NFn2JzIJMGRLApeyoFIpu9Z4U+18z8GVv0
Wa8q5AKJ8abwhFr6IU+DUYWJdBiEnPregAfgNEQ5oDdgEXISvXZ281WENoBjSOd1
8nrLBDKwI76dEw/lvMrkTbLEC43sYIrr+jYj+aYjYPjAlFSu6BPSDrsvQ8/9j+lF
TmZBUd+6a2gW+ytfRIbf711V3O7COi+rXcffaTvbGflwGgWI7qiQkWdJ+nh5me6/
Tz1N1EOZXJKrcFAQuJSp+n7nLBDarhgib1XIyMNrW9sJrqqYcxnDwcNM4BAxluYl
Gy8uu7A35J68fsvL87635fhIex8gJsUhdLwIlQwucLpgkHu3/s+Ug5KJSe6FDm1Y
9o/4a+FoLqvywLRnAjpZ5myLdAHPkjSNb79tT5ovfIkDxAdKQcZjwlOrQQfwQYoh
DrRY9g01N0Z2yCZpsz1LWTiI2K8fWeztbjuRGRW+HTPxCZYTBYxAUBFSwGaWQzc/
NujtCv6fKk+U+3EQ8cRmluUvpMXoEsX1TBJBoXSIsBkS93IAIuLtrto/PdT6ayEZ
4VILIC97CAmiBSO9Ghft9T+YforbOuaHAgUXXMkaME6WdX8rcXzD8ZxnKAcYmDdR
8J0UhIGuhN9pKMf258L6IDk8VzFVffzTYjfEVa585T1oRCKt+liIFZtuoiPQbu4S
jHLDU3KMWR7ozQgnb7RREygxzbAbv8cFccntaq6W91CpPDADMm3UgG+ug5Rl0+V6
U6dFaeyasnbK4+bkplzRLMRzvdow4Ny+XGsOa0ZN0mhsfo2SaEKvwhHzSyYVff0G
R0RRy1hI4mE7ot5OlYVc6zLoP2EANsoZrk8Rfnc+o1wbO26cIOKleno3xuKc2PyL
8QKP9RED++F/3V7tx6fqgDPjpVtKq2oK0Il55+rcYtw+jUxvBSbZhGYcGGf4UVSE
Ca4Bw8losFBq75pYTmEcH7qHw3FVAvuP+YLeXzQxVTTD5pvIs2eYvALuvkZJ2XmS
dYzXOFd5h1jh78KnpivOrd23Hl/WcbS268jQ6SArye747Ixg2i9ap5GLKctnNTUJ
6BEBWUVdDikB0d20127T9hknb1UsE86+Fjt3gL9IvQZWwlOYCoOTWkB3mgPHzyXS
XuN2fP+BBhfATRS4TmNZj+DZwIBOZ7tA0fS2IGtx18p9Gs8QcoLoTj3M65AcEkpO
MgztHVT6jS3x1YUnuSsKzcrcefdRwn4O6ettwh4cn6d9JL8vqTdVceQuPsIIIxEO
5mcIDKNBu8kzMffsei8f+SRIbKBlt0entpSacmOT3P5Y1jqn0W1J7nFahdGnpq2z
s/U+CeGODB2W5DBOfdTyvsmShucloR9dMZqITWZtcMljPU3kEfYu4BPkXolWSX/B
EFeJe3gtDWnWeh51jT49CAcl/kWSRwie4y+kK67JpKGIbApxIVwgkTtXM34FBP8i
bcnxgGkD861oRiCHSEeSHdD6JBZQZGGDsEOIIlLNeyQOSBOrF82ROXK9MsW883Sm
vUUg7IBTHTKf2MGnlYKQ0Rut2b1lrJfhaCcnTi1+Vm+uEVjPmdRba5g2g6FyCQZU
1thyYn0Gtqc2+4GxmXM+LKKs4b3MbYgraJ+4wnoTxPS3x0ap8Ky+Mr0g5f3MK/Uf
yXGKF2EVof9GhmgwoihHXsLVKKzyneKWaPIrVjKfr6fbkUoDiqXf+q+HKbiS0MjI
qPFQDBiIUKiV4dslUlLyz7pwLhpRJCqAEGmxUAAtkaenZx7DuHO+5/B4izFx9iG2
fayetyXdYiqsn+xvJ7Wweq18vQRKdci2oX7jdTFf/VDCjrV1vIuZHwFtxcn46dNp
e51SZTxcUo63FsT0JM83GAG3Jh3emip/VlV9LYNaXr8+o16eA87qNlK1/9dYHvZl
CyHd3yKanCsFwZ0IuWwnP4WRJCwiCkNp77nDCAuHdAmqtnGbAWQowYoxTPoaB2l4
J/V/6ccJUuLfO9X7jUiHszZvp9yOnrmmkJJmrTwgaX6inPip67F417RnpUWBy35q
zivYa1J76o9+c+aqKXMIcP1d4g8nf20dS9g/Zy1HWRcgnnsFx+0RPUHBklPr9BAk
TLfa6N+EKibn30uq58i7GoRCfiwHn3QftQngAA4pHDm3dV9b/7gCu7LOZAFxgKaY
FMaX/Sqn2i/JDGLpqkUzJVv/cl1+j2tQfuh8a67hInhu/Eoc/dGJV0ueg1OFtp37
OF5B5ASh38F+m7z8RpztREMQZGQ7ZFwovtI4YK8iknm35aNTI6SJkls/3RqKj1Gq
01gZEQFY2JMIIkX/MVMO7hCUKdHfZ1+B5FMSn9s5GGTvkAZ7cevqmASgl6pO3Fft
up39OzPXGRt/+4tIZOffZaDBdddrISiGqWU6GQGs5gEUEBDgTJG5MMNZQTIgFc1g
NSm/b7+GAIY2d164M22jqW49ZkYRLLjC7moFASztrzdJt+Okt7afXDxrLOCLAXYi
t3xyu/RUcRhHCMUZ1h4AGwloZ8D+D22uYGT1X9lQe2X+S01PvW7GJ7wlaHp5p1SY
GZCAsthatLEHskaib9PRUwBdX1IB7dqhFd6JRVHeUfAbliQhV0VDbhUSpVYJnQdb
jv/+shHZ+XGueJ8tvntatZUso9dvPp7lq0rXMdU0MD1AkhcPwQhf4/ChbLRb7F7A
kd2oKN4uphQTTmHmbahReBS3oPAs+8/NEv4bSHjC0skixPb04nQVPjoP1XahT6Yd
T0ADgOAgxQh4UEJzo+uTnSyW4/6jzxvtEXWcIJhO6xbK1iWFdr2n47aWk4FPnqsa
J+aiQl71c9t3zUhMKj0EzTW+sj3b/pzC9dH9fsbsWqZM1wyaT11LMrdFE/SJPtJd
eeVPia+C4WsdmteiZVa+5ulJm2ZUTZQSUIYvKw1pJQ2mtpbjyOm2yqJA022NgRxQ
0zO6lYP2n0DWl93v1U9mgJIJeCqe05V3aZ/2O5U8hMp1gubWoA2O6DUWhOMQ7dmL
Am5hIIUP9X/kMHK7ohHiC/JwZF5pnQGj5Uo3scTZpVat/7j4wHgQu6IaQ53gXkN3
4hFMwYhPvF4OtOUNuGbVnaQXa/7ARsxnBPtoHk+w6z/yXT8wB+5LOli0bf2/OqoD
MCBBwbXboZPzylnCR0t4VtybOASTlCGpDQUE7UnAgVAGW323//mx1nuf7T2VUoPj
gVxt5upa/spGVhrrv2ZO1x+2N61RiN6JA1yGwulIVcqVJgo1ZR1CojfTZSk4jLqd
wsdYUcOICWsVP8dAeC0v6j3jmxWSogkebvxShoSvl+miWwtGyNF1fFm9ywxleb+Y
cSIYIqIM32wBg2NZUG92uYOLnJEPNHo5VoJir6iAWopoUKVSpWmKsOnAc53DRUfV
AwRnfv/0fZDkIsQ87Ys5IySJ79Hc6gFBJdSJ6U02qUkS9cf2UJphvXNFv1Ojymor
vNjZKos2OCOBz5/aOOj9Ds0pFfD7/LgeOrI0RV+HF80Fsx1IbfnfQ5V+6KWkjuV9
izBTyea5RLsrERpT/hs2WJmhVedRG6469hLy9ZWe39/QJW6VIlU6GD1H+TjyPBxj
8UTpjlyhybBPez1de9FTwlNT3xvaXANWXyHK12YcG4JhLFY8DI3NAzEfYAP5tAot
uBkVwO3Vrnbtgj9xBwwfOGTnIIy0ESPmp+R981zAumsAonjEwmWosOpu+GwhfWdL
Oc6eLcuFE+eNLSziFZEHPfRWM3H8e/wZheBcOUhD6WFn52IJ/NFlkKvb/cepZWnf
yOKqzRoNMfpv8ACVW2jpCsgcOPvVKBJZSRpUL0ut13f5lP08tWHh/mFqAfZEFtDL
4dbjCU4n682bR4YDpBZto0+Aey7NyPjXDnTf+bXyVSeN9+J0et1eu47qXnt53Vo6
hlI6DYRj8S4Li6AATLmaFZjBE+TTkzNEYFWyskCWO1C6w1tvwbgchGRZ7Gsrsxw8
E505VzpH6kKW87lU4z6gqn1BcBDKo+5cNJGAHLe0RDZuiuS51W8bIJQS/4+VoGnn
7xU0wbp+Pm+HL5EHe6ljjIWptQ06k1sHdH1Klo6XxuoFkBvZP6ARJYXxPCMnfwzW
j/qllTOw41jlCPEol+1o5CrbGl2xUtNT0MlNRuikz+AJevdft3/cdTGbWnGW+oZh
TxGd38XweE/EBV8T7X8ILk0+wpITK3ri38i4BnZuX+SE0KHgF1gnSPETYnfDAJSY
HNhBg+kbCAhWkJf5nBKIUKpIavQIxo/eqlaL5QshqIDvPi4vUMQczIu99UEnM/Xy
TxLcWakRZs+EiUhv0IufbMxjODii6Iu2LM4zfiTwnfqS0PgRNiizcPb0jh1mNrEm
ruSl4nyN7s6+Q3L4UcGxdpld6B93+Ibh8/ZALGFrOidH1pqGV3CJI4tO+hQrRMdz
HGEuXDSDnkyTraSFA77FswAgCDPtdy7f6np0Jr+CvebZl84yOsb5Fhw7s0OHkL8n
Vq/rDExmQSCgyYFcj0cixVarJMpFat/Els7oyC+Gx9rbndiWRySA3NRvedpNxyQN
v6pxUNvR12Q/lrAInaRoji5VdjAetTgW9LJ2Q98q4O02R2zdl8xvS/CyW+rPd2gD
+z9k8lLVlnB4S8wnMP8F6minZ+1Myd8vi6jKVN1x5AJQTZtM0oV2ehtIKSL6ZJ9J
EgXJWcBf61RTzYE73iFgnmnfD4IRPPozQpzqTkGS1Qkjz7PjKuMFMRu7DFMZfnEA
mfBc6R4BUCbBaNIqlWGjd/u24mRLLl/WS/4iFKbqi7WzHogM+7i0PgLzHS92+/mo
JagT/TQQnv4OjhZR7bOySFPl4167rw30Sb3EMRlpqaSVC/ujq5iRM4ecro03GL32
pRnKKGjkfgyd39aJUracOLSXC5QFI0WcJQpn0zxSUiM+HWf3QBejM9GkNFKMbZm3
MNsorUD3p93Xfna/i+mah3e6ilx7TFMf6yd8P2+rEoYUQPulhDknbKseW3cMCQM2
mg4SAie2X8NDSgtQr5FvN/r4Fss8VzbIY8cBTZhBKro3A4FXAI7IhLMvrsjyVjnH
5MDPQV0R2tnmxwXFRC02OblZbSqPdvm8iOioG+3uZZGOGnMVOSPJBIxSSF705ge7
55rMAuYMaZa0Q6/EJAMXTQjUA6PZY2leAG9P1N+OAbiHB/8rh1T8j/c9u5qdXdn/
d0sD06wQyfqVAe7mVId35cgNhbE8+u1P8KHEKzQccLu/q0ADiUzWlDknvuUlVdkh
S4in4vMiyEVfhpZqafXeZ9bsu6bvk3LEPkkkDGRZl99Lw5vYCeHRb/GwPVcuuOT7
oVnP6cD+OKJRZ0dIkC+7CYRNbvXsocNfNCYDdzmsdYvFLIqiY3aSdMS9gLOS5WR+
NAJBG5vdWxYZ1e3uKmKfScZhOrI1qk6g8x+UGRsx/i2TdRYQiGJPHyrZwC1Rc3dm
ncvvj4YnPcWXKK+dbmVZLWf5K/AmpGQZqLA68jyzA5B/Z8CJoFnNQ/xBLmigYtBL
Zl7Cj/YFUV+sDjWPGPGNJlkeZyxPYXjpBP7cft1qe4L6wnrol89DHw+HCHJK93EZ
GE06BJg+/TVKBgpdovC2ZBZB9m8JB2gmPIaz4Y/imJsmcaMr+rR142/RNBr9PQyE
6dir3Bjy7+4NAAWMKdBtFlelHEy01irSDyrR4m0bCQMXoojenfscXLC0krluT2Zn
jau7NR4nZHf34x23dTJMHyIgVs9OSfutNytAtwguoVFxzJ40FhgIM6liR5qMEDMH
9SrDyjI+fzLmylswcI97GwGALjcuHS9bUDjgDt0EN5KyiwTvIUvuLDEN3CyatJK5
MohSweaXneSqN/69XRdJ+rKcOQd4lmddTC1p+mmD7uhfU2Spl+eaMkBBOrCDTcQP
rSMYbmJh6RyTh/Z+kVQftzeRcU5csd9/hft3ZtUiwrnilVHvJL4HaWE5KKyR6R3K
uO47N5MBisEKbuLH1JNTHLHnjjmTvgjFNpu1FvwmxvwBlextMzlXa+l+yiwAY7sn
WAfcbO6CRDnJv2ocTzPSZX4itbxzCI02mFXKTj3aXauFrrQ+1vyMyxl/Qbd5KijB
tXQXhyckPA98C6Z8DLGz75DXckRa6SdYxpb+DKOwaqGKWGS7qrp/HMHxNltnWuEM
IhCvVq2VmpPL1kgnADY10IUo7+aWYnZu8BJazpnUaZRFbO9MAIN6Hpve4LV/0wwE
2zEjfL8OXBuMMHYPv8BUlGbGB/lWI3AQnOrlJwJyYWFUMOhcYhYbX1zFmtCtq1eE
5uElxtbd994c/gshwbggmi6FA+iURX9gHqzIaSuOxMjjEzBkihsnZTtSJWfrBWGQ
X88CudnKMJAu/AOURFGwtnbL03ZEqt2oaD3RCTjODOYGdIgKDB2+vWg1kYHChs3n
g2LCce4FGgAAzhezeOCHjbMKz37fdn0jRhL90q4Ub2TYRCjPqZWzeMiGpUXToQhW
MaHt1hvoTD7lCeZj0zn1rBKVz+o54UJONgV/l8neaHSVz8OJOQkmLBEhdEucnLNx
OAHoXe/wDAZTwqgdoKNBSnb8OvGSSbVEy98oZIICL6qGPXHkRtKLP1ZgO+8JmsDI
pZv58JRCOtN74JgDvm6+PvBo/ia/JF1pPzi6xt77PcaPNZ6iPzb+CD/M6rzeXjCY
bfnHD3Rms96S+AuxDraapTv8UQ1v1ruAmmMTUavcxcdstlbC8oKJiRiE0R22Vcyu
5tmJOgaUVxUhvMtxtdFgIrVWt9g2Xbuf0/quExJmcQ2ZGsBWhnDqyR12eqTesP4S
XjTZaM8VnVNNU92znvMzMLp/So+m0CrQaINtQnlw/5ZdkUGu8jV+ipsGj8pX/MYu
0CJAik86O60HbFOFlV4XPmSPPE6h3ECf/Ew5t5dcjtbkWry0SbUqFayTVmpsCRFl
LJN291fbI8LL1HQFsn8P1rgFte8E2lAT5ajc1ErDR90a/hYFFHQH0xdvdYXnsUm4
EiPkD75+TyIDMwViUZ7bSH4+ai9sTtKPdFYlV7dCiMv16jo3lFxNcqvSNra8Isf+
LaQZ4Bh5/cY3Nmv+hcBNBX8kuN6BFYHMAR3DGUXbZFSbqlsvz1XNdJlN3Hg5mZOc
71540Qy2vtaDhtfgOMMC1fIpPB0snBtjIq5c0rEO/JPcpXXp8x4YipTdw4Fd8TDM
0C5LSAfp+ZYAVCExYXlY3g93WwB/bzmb8ws7KdS7WNF0ySJyogPaCJ2GiB6J6ma0
O0GueuTlnN2fEiFeQy1PnJiEafu3BUi8uQ4SKTBfYRFXruvHfnYnDpleFlySvY7j
RrwTO1JTnjAiWLCmEluoEv4LXZvVO0iSrPRLtn7KxqD4YKcsnjHC2vuKz0h1jnac
/pkNPyQ4NNi2gKUZcXPqmP+1xvuap2f4Fz8PIyIGDVIV/ow4dYSLD1BjdwXiIle+
sXt5J0KKoliAtY5xeY/Xdkq3zBDb7UvG1VDD50sWyOyu31ei0XlZmsYL31/17sO2
7QoedwQmrYy3F9XAZEuA+4phCkcLBfkkg8Rx18soIlGoGO3T20dOJnYEMS5yx94f
pUXrH1UotjoOvxvRD6ZodpT5P7Wt4tFzfugKkIKljtC90uVcAHCSQid0hlL9WBor
cntFUPMOiVdzMUl0x9pDa2I0j9kWpEkLGOJSDQSVBRCpc8ZQGf1urlUt7ih0jU1g
7xghb1IemNCtOPHxBahogWRRveAvby+4Whz7aSLvNnQAGvYhfOIrlwm9xmDIExKr
xZ60QYmERoOwmGTBuBj3LZuuDGdZ2fBYBJZOhEWOOZQG/YOzkkcmZTG25RnzhgpS
OkQDEKSADqul8IttW7hKJFh2aLA8DM0jUvuEBv4PZzUuw/ISpG/xtWxMw27p43bu
xcHdorWnTh9rReXTKbuHj4CTDzhl8mbAyY3L9E2YIr3pghTy2ByMSctkw+4cY0Pc
WpH6sz8qrT63Smon++wqqZa8g/NxcgUDvL0UUm0NlsQVYV7Wh4gL0PBsqDTRSyP4
AKxP37K7Tl4wRfaAnWb4hl8qNuhBS0Y1brSPU3gOO/kWU1WOPcpa2mT9bsy+qMQg
RuKHzBUwbvxulq0+vqSF4KL3UXfLxdVOWbM4nE38BNU1td5BEFMpGqsDc8AimM9O
xD4rcNZHHwm9zftw5svBH4pkCh3CrwDmlpqrQAV1znObSfj5k5WfuOdLRWj4HXOb
iPwKyvkyq9B5fRkcA3ABdVGZitH9Glv0MjX+Ni0OxbLPoJib629KZyqsSU2iW2u9
IzxKnjQvNG6VrS0NxIk0khzfSeHr7kwISIk8die7TG2Bnuh/WNJ4bsMWhBXXpopd
JudwAfJ+Rv507ZB2FuQnMJIvbNnmD5QeCX+DGc+zzMu5OWQQhUBhj/qEk/GAC6Ov
saC/Pa5MxIS5HqEyC/M5OlHux2HhDUH2aCSblN4DMGAXH5lu6k6V15RyaNZeTcIq
+8UElAPsEkR5vNr/B0GiV6wiJZ6dybJY5aS24+lvb8mIqMipzEMixzOAOiFvXobm
YWVqpSg9fZZsH5w28QDH01WoUJFjBLWdNE6hlIMZyLao3Zv2SRCT2uLokYPJYCqn
ui+Z92DhlkaDN7YYo4yTnyVCheGLITaURbOWIHTyImP6kbbILj+8t2tBubZIg9PL
wYC8sXSqyK69LTqyige6ysaaOlX6Rq3lTV/s3bs5wBjCltAwtV3lzjYE4HkjSctO
qsGwfHrail+VglscnaPc9I8iuPMQoAY5nkdKWrHHFa1XBhmz4Ybh4EappSal9XRW
CiSnYCYZTfSg8LeT5F73J3auuWzJqG6y75Dd1Pxt464M9F0BiYxDTMj0YzTSXLrX
Iv/dqhR8DM+SsXBgtSL7I/89bIVJ87umGDVSRIol7BxtdfKlUN9Vaappo1q9W3sg
IRwKr9LldSNPZxJPOBX8Rx2eBV2cizh/axItRNKFZ5wgd1zEZ9ZfDrdPvsdiGHLp
5tPmF+wvyBAbHXKICeaJBuFxZK0MmXqJI29zzs2MMyoe6jm9PvAKva3nZtCtdpLn
op9PTnZaHtz5v/+QH8rG1MTY+r7U+FtV6a+mUVv49OkZdVsXWTHmbyhHrfo1fTf1
C2WqVTXCdGnkdY6fIHeQV8sMPpyHa7QDCFJ0Vb1ITB0mv2bs7wBr7TZIlKW4Md2Z
Ghm3t7AQJOPG1+6l7nWEeYG0yUpqqUW1V4HFYZptaRHCP0ESXwiV2agzDYdmASFK
lSGiAqydKHW6ezde6MXD9W4xQbKFRhKM2DE+eQ/nEkDDftywZ2T5IG9qKuTnPfTh
MO3jAGV4ZSdsJ3lhxiSknLCmHfcOvOoXjIVvLQfF6Rg+DXJbFRfqTTr7ZLGhPpsi
ejUXeWswbr67GHPgQg43lSNY9z+JOXGjzY6JYaxIP0dj6iBRY8+D31NWpJX9290U
wO5IWENBSe3cQ+JIk0oO6nSI425KVdgJbo/YcR63tpnFgIbW02Np+GCdd7mFBqpA
1hHePg2BYqBTif+AItZq6xjYm95TG/pB4o6cdQDc9hVq5LUGM9mS+Cn3MGKPwFKd
M2+ZMvFdTy8T4xvdxjCQ5qyVjua8Rw/GTt4M7FpOm7h5LKy0k+GeGx3ezdnPQkL6
9xKiXvHnS6h6pR9dppFC5YxnLV//gAEfVS0eyLLSfZKKU3T3S8h3cIQcUSwTeW15
hRDHfQX9Lj/Zgpy1JRPPKGt/1cIEpSyEHklNy7jI2w+AI9c250kwRYKJc48K80NZ
gzoJDarpLl+l4Vjpx/vV2uET4iTisuLSSmUIrbW+HYcPH6r9Kod4i7TCj3M44VJr
9NXKZPcq3HNk+NctR0TPjmF+JvCCwZV80L20+4rsaSmHhFVCY129fU6H99vua1EZ
iNeQVzdiCLc+AwyItwBYC3ASYTdMBxio7vlqSrPRk/LWxUFHXwMDmu6cosVEu/SV
77AOLil7PMrQswtk4dWlyf+2dt7rREa5dLyrchgkBYvfpl33LKMrEnKfhg7huqSL
jGZ+/eoPEou8QlYlKPQMysv3U5m1gWbw0PdvxdWw5VGQUFxiK0zMnT44mfgf4AI6
Ui+zIoIDOh165PfRwGzqe6K4ADH307bsM89bymdwI9RdEH4nSBz1hqqPGcaj+rrU
2Mv4vuMrqM0aXRFWk4o3kMmOG8+Kzpf5K9+abzRYk1d/VMGrwf8h8g0vH4AQVHqI
6JXS8gs+yshzlnw8N9Tf86/lZmDdvO4sj8MBIluoMJii6+7j/nTpFlMje4gEzb4G
jVTYEXQBZbkjWAxPc5h6f2xJh6uWcZD4MJ8Y1gZRklvfU9UG7ifMtO6Zwmw+k/PH
Nhc12GTd0lKFZ5dsR0QDayhvmEnTSN78b+Fmjycgd/EuF3VKHeXwu4rlzeTHy2On
888+uHgho+DASzc79AGLFIgOBERX4SkQaWk6nU6ntyBeDEqPgHDiRm8kxsYwTK9s
ICtYszRjHDZJhfP7SflPbD9i04WQ2qaU4divz4fQmlMibHQa73ZefXSqpFUClP0I
KpsR4NMQf9PccizkLoC2v23NHEz36TfODQasYebd0R8h4vZxMxIxWaN8BukzmtuZ
1URVrcoIEBK6fIhfHay9mvSiQUNAjyw4vq7YhnZDGbU4NaAb7vg1jACASNXiwSYW
lQMswnI01ToHd4AspoGYnf0pYSwBq7ozCs9GyUx3+7wKO+09DXPngcg9GNIevUdj
agKzRF4trO24rBIdCvE1z0AQUAQEOXuMtjItYKdB4d3vvTse0K3wsq5WxvJNb+9J
/Vr0l1MSmQnkLcN16Tr7H0CAAYMdlYoruOxuogDfJ+TGUSWER0h6C82r1JoKk6t+
yXoMHcZySmAxTUELc4vePlWHbGFBdU5PJm+t/DzlLN7mgHaxiUEsrQ9POxNBndOS
xEs5M4WLdt3RLQWBqgtM0lab0hS9HFWwdnI5he6SE5FchVYsz2lt4P8uBxXM/TEo
+NUp7GTKsCFguQZ7WDp/cYo7Zd8UTbhqCtPjP2UjlmTV09ZqZmDs0VOQG3tbx0bb
CPEjqo0076fkl5E2Vh0c5xceA/0RHrdc03+5vwKbJpaDyyQxvpEIx7wK+RuUSL5c
MTJHyihRbqRLjlq9A3SXGrOgUI9jJYBHbaaRQ3EesJfJVYgAr9wzqWIK68sarscX
c49kpirLO9GrEnQPcCZ9Py9K3OotSWQiGwSkz5eF94r09O4vWPTk4n+FQJ15CC38
RQdvjG7bRse3p+N2If9VyejrdzAD/0BoogsyQzB/gpx1ggat1fJ9CDY6abbK7NrW
f56AZcz3OUiPh++Wd4sTSMpDCKVb3Ft1QVHmzao7PQ4E6DYXoe8JGU95qabK7BO9
9wWjso//GAHn7FG8/gcWImUPH0kAj5nilVvSGVajGjHBJ3I/jl508fLxtW84jltR
T5zM6rHFINEw5u3vVz4WlWWp3tr+BcFvSO2FkmkayY7wbFj+/D/98tuaTMJxt61J
eeA685vkGHMh/zB7UN7qKgvWl7pWJClrCt7UPIMvP+d3osFy8j9nOB6T8vlIGFP3
VLTsvAS18SELye8B39AYKPHs7gHh/SXJ8mzL23Ujov6Y+Hyn/Me4YqgEvWFMHe33
UnEiGpgMsW5rgl+47xz57Ld5XlajLNtUQwgIJDWLPvgKaIA6pxT1WKlhOKRKbNht
Im1VwlPKUNauR6SAAh+c9roWdMJQyJL5i68disHzjOzIDd/FPH67cmlpqcp3j+rk
mjNLHgWyfh7h/99QpH05Bk84oc+zlOPYrg4BPzGvdUeCEl0FUmJ9wsP5tD/IKJCF
2BA8S38wI6YaEY5mCke8fJiSj/CLFQgOY+H1x+FhRqn9mNlKZVu6Gp/YPaEjHhvW
xHLkEchdpHd5U+I/o/AX1rDf/QHy/h+WK99G0SL3JXdO6iQ279/AH8pAuBffoLrZ
vdYHHmlRqO70bbNm2E75qLABI+RDcrbeg2FGBwKbeR7O7cquGEzHogvS0pFw7K98
zmwPplwqUDkR8/+FY/T5kv+Wnkrn7bwOgafnDnDNhkoWNGfGBGJb8y++X3H+uuI2
cdVP2G2CcG6aRA6sJZCoL6/CAL/Hmh0tQ8ODudYBVhyypc2LDU0ZAqyAkuMSUy8H
EtQBA/m/WvyTcPvLJjJV7EhHnPRAJPLvMTg5XwUiaGdk/KkWvDKLX5tjsvYvhs4r
Vy0NjsF2a3TxhM9KZSlC062W54DZkMeSbBhrSnBJcSqqynNHLlbvlg3W8btAfn6t
ZpRL6HsQZyDufHpJgWcctG7APkPNiKgudGmMlfflmFLNfRBGiZosEPyuhik5DDUY
K4jQCv/aIwMOM2sSvbHykvz7SKW+ASjbwL6fKxx0K4x1AwfGFUYzoYLR5ZYqWWZL
BBlfovgvPtx5uyxZ+mSiiAwogoHy4NvZVs8CC4upCYVg3fNA1BkoBDd3SrrS+NVN
ID5q7TIkeuqCqXwn5zjJnHRT0iopQjow4XWRhfqqAi11T7uYs6KywA1omTxxoZUc
UEiI/hNFAGM6k24CLHBxkHsscRfpoOaiRQuKlBz200G+nDkpcNlzcFEYH2AF1HDT
ikkNfVf3rrivuDYCG1nP7wIAZBsQVdlazxMsf1uOw1xW5fHKOJzUi3DHEREQkp/U
as5C84x9g8wvrJtf2soEKT5VD7F/r1f4pGxKI+39CPCAm8+3uEfhWwNsOXnxDt/m
hmv0lDR7QV/ML6cERA0GnTdbYbofBx38Gm9V+XAFHIYrFc3ujZsyZJ9S2jEw7YV+
mQxJFoH+DszCQvqYCE0plePlCtDFckAvKVl6wNe09vif1w7lINQ0E9o8W4dWGLyw
b0wGvRTHy6BdU5bbyoEul3ssPDGVY8A/OrAulvjmRNG9Yv9xAhRC4iF6ikGASffv
qcVqpFysYEnNnGCbuw1xMfG4Lw6zvg0aNEaZN8fAcw+DznTtGv9Ld3lp1Vjm2nRS
DdYw1FDJEdXshmslC0lVZ7Gd+fa2jfhivsSOba1hvlWCXPPcVgm2c5sZP150Mc/j
BkUKQU/OP8iMVksWeZc0k7EvoEfmgBknQ5LsyBISSuiAkoG/1LlzziEeVhI/J60S
1Jpm15B3Pqog5obZwqNIHI74fBDRZH6dYfKPBFm+NS620FdnmRY1EhjxSwTvQBaV
l4xu0cWNese3TEm96jPgxvQ7+CUv9vrqelJwKVgbjB17z/2XWS3jaAq0ZglN6z1t
/UzkoPoC7qnZ/Oz37BfrOc/044tjvBZf/HJGkRc7C2+Yj5V8MoPkbLBXWcPKRsAk
AisG5UftjHzez4S6/AktCPAVBip5VJ1KYQb+T3dg4wSszm53m38UgmoVvT8wKw7E
aT941P6WJgOdZN98fD/igkfrh9VnSdpd6pBfnWbph5BLa7BNTkSYk5CWbHtlQLj5
DZvAasjXfvvRgVdWozEN/o0j0uLdgevukvWAZFKWQOPYO5aF1JUN4cYiVfl/jMUW
OO/U3PZbFV+t7aQ4zZTjftLX0AO4A+fEFgvh1LgklB5KoNfqwN6Ssav4yxmx2yT+
ABtEVMEZKibYqq6EI73NS14dDgxGY5Z6eNJtMJiX1VPEL+Mtpv851VS0oqN4SyvI
fcJcI+gKN8rLj9Dag699q9LLi6pM36jOskE/29kw/bYeqvvVW8AS+iRsaeSpW4NB
FryCJRxqV+SeW0JRB5mqEkgVPC5fQwaQBWiYhMLtxq82zSjRP/ipEGX7ahOW/BjL
4AnIqO3cUJJvThf6nMbBcNCHEKi734Dbd8r1EZqwDnIuLw4qy1adc4k/+yy+a7d/
c/vTxdyPswB0vatCZunnqGgom9UGQPMY4lvT62LnQK8P+rpVidZNftUTMliICQLk
gUQLmZByX06+yP3R2l6B7qcdThAhPtmkDNi/O4PGfrbOTmxPHTZPc7V4GON6qx5w
08Q2M2cPwSO/q04uIkXhCZ/1ilSTYqQ6hmsGtOa2FN0DcPUSREFmpTijk2dMI7Gx
gv31OgAM2OT9t6iXMBK94SHHcGU4AC0bumkupxBiKzYHxQHdrxA57ZDTspifn/Yp
bMzggsYh8qVyRFAbR90u4T9vAgzRPqw8Mj2VQDxnWylG/4klHUCR1AB0TwnXDTY2
2rys4aKWOarGn7OKncq3WxwTyav50EjKPWBjX1+L0LfX6ps4LwdbxAQyyPS97X8C
VKuYEoSiTsS8+gAtXYvkiqYLGeUMgraLXRbycR1IaoVvWxLBldsTgRO2wn6THGEn
YYR1EfNsOZD3k92CqpsM+Fq3YGm/rINQQQf5IpUHziTRJqY4RDvsX42hjU5oph9d
V7O6PgE1b8JgnOd1O9Z+VGtsbVMiIdSyhFM+wKwF5mvvzfT4EZvn+hbdbLs3F82p
e4cFDfJaJCLvd3a35hMbSkkLMNM0YV69ialH+wmBvzqDsdiKK2lgsvUaQyjvVyjS
mAd+SmnV/CPH3OYwOIiYbX4283siR2hv8pqSCvUEMZUhRsl8G5BCuN83zmFa6cYX
pxDvj4mPR6RvOnbn4MT72P4Hrhb27KWBOGh1e32lLNe1cE1dM5G9QyelCjYiHrJk
HtAzaNiuE+l8F1am4GYXMD8mbEvqZfPXpnr3YDyAGQQ488Q1vhetp2nWSpJYqTJt
v7waPfhWayHpnmjLL2dAQN6DUnbYMifY02lQ6xzDBjGhUYt4XVQhCXOVU6jc4TWM
dXFk/hdcjcTzt7HP1b592AvbAtf5+pixcA3dA6Rv5IY8q1fazkzBOrkqYESExy0C
SNRrivOnaJ08H5W1xocuxppM+H2/CAtWXQm3WigIHVNljDX932JuhpHkHPF5oVMY
IunTCZrL6iV+YvmiOnOneIShBG3LtXS3bBCXAGskiYrXukIHxB8bUy+1ZCtdEWBR
FQE1tF1Ac8bCV5I5OjEPKYqGepzVa6ZRY7xBoKL0mYJ5Ks4qU2+BwR0F8A9I/w4D
tlZ9FkW0+h2OgjMtXJvEEh4m+PINXCEYI4NwxXMCumhAcctE87FQ/Q3OhqVPA17v
sOD1zLZ805JKprQXHmH/JKDLWYxE47gEKPpPumAGGM7KCNLRGHu9c8H26kKLKWp4
SNwA6W9jMC5E1pgK8oRg27NvM12q/PEKzx4DhwqQvnahrlIvKd4P91kGREAgQHVw
OtM4jBtLuqTDOjrfnPL/DOTR1HUuFit+7EbcGUeZFiBWqMwAQTTjyZzrL/Q/Vsrz
xXdX0ZxuT/8fZ9ybQqJTL9fwirxRf7Ena1JPJMwKlEREYe6JgsxokiwJ79/ezKuq
KV1wZ60wV/mVcgeNAiQnWK/bFgJmlCvP1U34IrGDfll7vK6y3HvyoyEk1gNWWB0o
/EKxAVfKs2LuljgrD8R6qHYduUF+sVG/JkKCTJMdSwwxPCN50g7MUx+RsIB6rMtH
+AHfE6Hw3pOqZlYCG3Vpv1blCO/6fjDkmHU+r5lmBb56PGskClqLyVaDqtQA4lNG
lopvA0+xtgWDV6F+Rb8Q0M8TNwQm+GIEl7ygI7cT3LueyaL53IrvYM/WdIYe5W7p
XZ2MuBjKNMmCBi45jPkS4hE3RC0p0edD0v/8scA7SPPDiS3oGHA7iYwqUGj+mXzq
PoBaVWargSBg1DCq85PS1GPGdymlIpht882dLrnyuStSMUL7QvaJ4Jy1DMJVXQEW
s/+zyiYNU27Bjowrl8htpGQrx7ljnbY7G5MBhToXgyvBdnqJhYRAboChLYjMQHQm
arYM9zNYzMUPB+Z1US4OrzfoTxuaQ8E5GFiHy2t3vYt2Isu43gV35pFt0UJEDWlx
SJwcUIO5jX27ugbj6zj0M//aemIulmsetBvRM4rH9atqPhq+mehaL38QvJ8fB191
/IwSuMTJFCEyTKpN878PkSBr2PoByCrdTbNwomGbmgmXR1OrFZ9PvXDe4SQzidB1
aXaGMcnTGGqkt1Tzu+oXQGcbHXfhgvAZorRX382S62od3jNfxE3T3PY1x6QGtiYn
PIMeiIKOau4meK2dtZLb+vjzcl+Gy9zdbFR18UOv6H47Twdnxcqew7FLezAq5Meh
/SsFaOd5Ws4741EFg1XmjZnu7aNbii2ML2iqOArI6BOUeYDmMYPKM3N63/rnug8g
HVUdRwPG3TH967B+iQyXdlPW/2pGcsHqLjO0ylMHAeJgYz71zeuPGrixMkGHn+sv
u9Ixzq43Rxkijy4BBxeFVmEvm3pclftipvgl5p3mkDzLDrrEPfHykIjXnv3t83p9
rODyqrhwwh10tOAhv5UowrZcfA8XLDYu6kws8ndlz7YSxANFUlz+DNV5fROV6x5o
b7LUoZ0mfsiIVxPGnpToxgQobpe0ph8swco/sDsIdbYDqjhp+FoZ5UvMn+0a7Lap
sgzIKeM7KqEY/7bqyXNIjQ2NT+H5TOcsPxiq+n47i7EadTxzmkavqERpYiDI4psA
4WwSH+ttC+X2wej5CSjFygPf5E27yeDCjNuC4AixSLxzYHXyuQOPjvUeuyNdeHDP
kHaswlxGP1BctFqkmgk5XJoVfsA/OQZozW10S67F7ekvnA7dS8lCqRCPAqc/c3We
wnrLbvmdnQ71RaZXZrq6hXhwvaerdoP8kkQJsfpyAGA6iwDLJztUFr32WSPcQrxs
tdm9RhZgwFGoB4LICpAxggirYkwE0bkmY5jIBPZZkOIrrVHiPLjH9KPhOl0ZYkwe
l+5sxuMHRw0tAB3Zi60j1kfREXnLx3o63AjcG+RZJGua/AiOIebo/uNTdpFwkUQB
oiaqOvq6w6hV1ZMr38qfqfh00MaA9QL/gRxSWEsDx+v1tixTSamAMahemzHNPEw8
UKm898PsXez8CNZ6kF/LS23tD9j702ZiH3bonlrr5jTXsbH0qPcfBbNhdR8IYu2u
uj1+pGoxQwdYFFceaqUQxX0Al+Ctn4zcNtdgAjg28RM5LwHVmOdZ922hgtDUojxt
UEw9PwcnmGJT0tTHUBmlTOJ8lvBkSQouDzVYrojiRnx0Qjzwsc5ZPVnsVRtbvfdi
3LuyLiGL3msvYDIKvhBkZIYBLeu97qlnKruw1GXom6Mv8APfINzFt8F8aYa1uceL
aM+DtpUTg6sAv6x5YBDajE9W/FwmpJLtuAvW5B3AFogVWNGC+cw8fXadMPoUjznC
9JvyoPd2U7voZoLt2hB6R+noBW7OVrLc4ACthWJSiLTyGA509z+nhtEwGzTz2KxK
mOqPXpBUSjz4tjjyvZyf9+QUjFb//YDe2t8lZ1iLDkc7MBeO7K8eXECxYNZlTyKz
9q6MQjsJU69RLpX0dfJLUTk+ExY0POpOefRR5YCuRMfek7Mk8ZLLMJNCnzcIjKb3
jwVlpzF8CbN+cwYvdXOj0BzjR6Tn0ELkSakkpYpMOqKx4VGIGXiJN9qFPNjDVARq
yfA+nuCzn3yfGHqmJRVbHIuEbek3SGWiGvVk95XXtdPCCcQyBT35w2VIt1PKYtoA
eVMx35lYP9BIDfwCRjk02lBkvQM5QT18r1ybUXMk4tr3xzoCtAruVgqMl0/nFCMy
7Lh1BP5Nmg444M67OJ5jXyw/Wmis00cGySoZp7YNB5/uEJjZR78ieKCYpAxK6StR
UrfgiPVFkwnn7Ur5ukz4Ybp8JcnQgKwwmetelaRfNPtZMUiQHwx+Kbdmz0k0TWCl
soaNRpbdYlHW28w/8snXdKLkJl/NkNyiSUS/4NfwM2Pt0121YLCjc3YAfZOYdy9h
uv0d8qbxrnZCFvH0c7hZLGBGFjK1dfxXxicAFQuqa+0flGI15RIDonA2GRgstZ0u
HUebckoShw7kul99c+MWvpi7CvqhLis+J3ji9AiGd/Eo3hmnhp8WFPcF6moRKcQ5
HnWaXLiEMuJ+Jrvc6QuBZN1vxCXztUVSlpR/bMm/6RwVFfPOGlxQQBHtiro9QTXz
cfS3FF21/jU5OPrT8fzSnNW4eziBJiu999ZSKgrs87Hfu/PAi3Gw0WNhMyMJyiuG
KPlki653BXG0a7oSiYRCs+e/UQWj7ubOQajg5eyUaMzRENcvvSJElQWG+RnbQ74w
dr0gOs6F1b/Lg5SSFKGKJDimF75tTMdWov8dwyMybgpbtBh9pHdlDShQlaXC1e3m
UygOPoW/y6Y67z56/uxZ5/JYf/LITgBvocASrg5t4QMYWqUSpLwqZ4F4qEDCPug5
0dgIKlgemNSDPi1E0qF+JMiHwqbiyRZQey0OMW8Hie9gSMwT9txPsPfKUQ4DLrR8
rAa21y+hRpyoLLiDGAdCkafvdJakCASRSJm1viDVKBN5HsL6ddVC+kZ4J/+lT5Q+
dKa8DnM9VGkyvbU4vFgBDbCCZTlhcdB3K9UzkRxrc6eZrua1e9hmk9HJ/OJEbvTj
xNCBqkDq94qupt4izZfiIQ4vLCmN8HeF0bBSZcD7b0aSQLjHzVikuO5YWLeMKDZJ
gWd7DdW7P2hlob3JP7GzjlYaGSME0RPN7r1Z07eqQzu+c0cYoYiFdR9o0PlMV66p
eiwOvyPd3jnLlBsHRj2BaYOHXtVITGW++Gcn9SL8ZZw5zZ/w1qSEbMTrPm6paUqd
Yle4+VwV7ibCLjd7Ks1QCGrrsvNIYroqCVxvKPtYqQErJQRev8QHlu5sJOjNbsjw
9YewvH6YiL6hM2uZS1s8SIuCcaCpikaN8OaFvpbk5EQ+dvjiM8eUVqsvaagm3eV/
4Bf2ScYYMdHTJQF1OuI3SwvHtYKJsd7VpNPf1/mFEqtqoWy1/Ju2MWQ3RZBqSXff
QFHIIItFxYwkASk/2E24oM2ud04UkOzoPGhc+P+98a1UTmN7XwH1sKZNRd4BtmrN
ZeEpwXHrmZJLqSbwplq0U/9Do357jv8bJbdB9s0Dko7Z075BIWrMlavJB/mg1eaL
MNaLYC6ehgJqiwDEd1ytLm5B7lSr8c3ozXyavLmMJY3ThB5yLz2CHawa8W0HToMQ
psd1N7stHF/o69iUUcuS7OfBd5x1Fgqxcem++Ub2wplPidPHB0kI8nH659dpCERp
hfNEE2+AzsIyhn/tg11wBU85DHSlKuHR18qpNWXhRt37yWnpsuk2PbAPUOLERgYT
8Nn7n8BEV+GoBFSFbQcULAcZsjtY0Hij9BZOY8ldFu/mkzAaGtJ5a8StQSgwPx5C
4xten+ycQNrSL6HvkjpjGV5jrM+73hHKUy8BiWqYJ9sNodLanTbE9OmEeJu6iPbS
RID5LAmRLQPRmfvrDEfoR4aGWHBOFNCgddtBtXsAoovTxFpjilHneUBp9t+Fk1YR
+IXewl8X2whZDs7z/bAsht7JLJ4NBIc8JIUvlov1ck5B8eirNKGlV5arSw/6sZtV
qIvShWSH7pzWjyqbKQBn+2yAteKUe4Wc9cmKIRR8FWX8bNRTqltgtZVSqP5OsPwu
mGAFWsjGDSJAZBayJHh57FZK84IE95xtbngi8YzuZQB/XzZmUgC/cXZvk1GxE5BE
5Qz2BUDa97FcWh1LbxQiOWpVeFRRY4Mlx9hkr/mWxAqdC6mF5P+E5VdXwD8QotFG
HVVxKbSTShHupFOLIVG3xVd/P7atqwMfCJ7PN46aMStNrnb4VbDdHCrtAevS75yN
txMIYJHmniRVVQmDh/W40rvQq2CPRQN9fYL41E26n8V2acW82A+6Kl5y48YyoI6t
uE0LbIrq7bEz22ea5nFa/6epjdCOxZOe0dUqXDRSLYkg5pB/0EkQNSV+O7D1Wm9q
9ims9FTJS4P63LMZEQ14OFs2RWGIAMtBPugR3WYohKxiXWCrWwXstBimN9Pm7HGp
V03wzO0N8AF14txNReTeeOQzJsGh5/qOCAE3cFuteOA4hCS+nG1AXmgvyFZeLeD7
AViDHaDHjnrUumA8K3dNqDJH6ijTboHXpZ4UT7ds0kAf9AQVdWKz3l+H5qAa/tg+
iDvafzSJn4i4yV+sfHIJUIClHwqiL+s1vfxmESiufS0a1v4JjK7XADqlzZuNuoLR
FBDMw95kkTeCszUDhcNwKj67cq70jES9ep4rsLC/0gdSN3cO2+BgfgKcKjcHmlRm
bmTkly0qdZC32D5HQHGUNwppU33/dBEf0uArMK5NZE6nU/Qo3NZNn2s+RbSyhyXc
PJZZiHGl8SDAMdM7mljw2JGu/eoIYEBOVn0w7XPUOFLvQVMOijQUZFcXDL/LXgwZ
Le1U+ktdWqBDm/MKURwCXY8IVjqNHQuqH/Am0YpSYt0auRtdafVrpnQ3UtcIs4lJ
pMl10LO0CbH6UznrsVMpo2k4qoxVV6pA0OVNl2LQ7+5lCL1OWcR1SOz4wjkHVKHH
ijcsFoGaXcB0p7Sbrcb2Q0SkLPr0s/fGDqN/JmnaaPMzOwiMIvEYaRCMDONX3u9g
YlKNfokBa7Um5YpBHEQ9qQ00uw766Avl6Y2CLVlks0i/L6JIjGctw6gHfGAeTL+W
BouUsXccBYpJYb4BCME37ThFnOh926LXYKKuQEj8DlxiKQtaBnfVnCVYw6ze8PSw
9LEb8Tcxd38rFNMWIEtSGEdnIYN6FyTzrBO3L54gYqtddnHj41cLBb9XSoTGALys
sBoKMdWVgMhEUjJxVq40EUnTyPw9FZvbVeEbC4gzHJU5QXUnUZ42Lv1HDFwf0u2t
TND+g64MOxJlTfhth80RPwzNI4hwzU4rfCzs7BVf/ohORcXiS4J2jZCihz1xZTXM
WuNnju3S3E3K5p+LUqs5y8EgUyh121Lkq06c9xzX1bwYnMi5FiJAJrlCIgRrli7D
2WwbEXMj2xkOoJTT4kh8Hd/awvMDU01tedpSzarTJLLp3X+IsO4CnZGnSxRrXAvc
P6cCw98jUGxcXPCqa81zcQrnoLEC9bXbXjSANoYwSWHg/A3rEWu3gjJ4aJA/NgwB
DhNeubFETi1CNCYawbID02N9NK46h6MKxf8ix+ZmWLveXr5mMuBi3aZhEE7RiDTW
by7bpw6oRbWhi88JUFPSDvUISp6jRjb2pbxTWUqz6FwVUaGwjbwnty3SVQCRv8t8
XG5XHVTxd9QhG8vsatsutv/o0QZYlfd0weUuy1uvkQ6dwiV+VmOwN1yTR0LtWgRy
2pttqIRUGPWO17enaCSYs8DbKBIp/+V5JHZTFGuRwDHQuvIkWrMBE5QgrAVkUp/X
Mc03FF7362MNVoLlo2ydhM+JycWrnEUJ4mGf0gPIDjqxHPoO3vYqviczG+0JRlur
UbOqqCbWheJ6KUpUl6mlzUemQowS9wU8WoAN7vqsBasGISPuAycTF3uJZxw09CI0
IV7bGD2vpxiT8EpsvXWpP3CJ1XSVApT18aD+AblLTo3721zv0LgQzdPUv4Dvlz1y
ZH5i1Rb2eTfJZLDHbDmuB1sW5hXSsBYdM2Os6nzciZ4UJJmZcOba1duZ4IdFL04H
WT+TgG8PVhHHuwT/YLsVx1hRNiQ4ooDgSC4t7SisBngXp0N9f8aiAvFB/cbFOIBG
CvfPEYu4JPcqbDQBtzE4sxifVWLZoiKZep0KROoYAlFqWZwheSKkOzdypN9Du3/J
DJNtpUQ/zQAfrMjVH00DK4jYiiHKCQlRtz5fI2f5HBkb51szqi+fhlGvUg6Xfn2v
AthAcCIuEDnFCEIvQz+ZZo2meki1750vl1ZaSKX3wFqnBx7P90ZImtxapRy989ui
aK/ad1q61iRf0FKNIUDUNUYdzuapsjX6wsV3EkZMQokSyxmd9pojEp3cJrZ1/tyw
I69AEfWsuwndTkitVs1BZU0+cYgGMIar1NJg2Qye3CSxbnagDb2v5YjFYvBQV5IP
ovOERwj3wdKrv1woiRDraLMAe67pZF7sSHKTlKfIESFUp4O9BpvfopPPm8hVjXXD
n7uhxn1XSuMSaZf2822n/4CENNNHWdxDk7lgpWOhrRqQTnz6isilPi0Dr/WWvTvb
8ng0LJ1cJ7VBjfpPUjMFBFJa7U0BouvuuPe16WyLG1fJC4paLclNrl2IEjjpmal/
txmhpT+GvZhdQrifV7Kz4ATkbcvqbEqOVSnGNGj4xGCo/XdWgHssGiBQBHd84w35
jsIM4AIaaM4k5ZOxTFgrJNh/0SqfO5PFkA4pM3ckte4vwpYRnTEA2UXJ6JOz/2VT
Y8ZWDGAeheWTBnRiYVU0xJ6J74z89ALhzzCjFFJp+W/ToFu1bN/LUd8jQOtuf2Yi
iTUwOWcsJilLemCV8rDBmzMfZJdTvCdYVL1ZoSygoKtmyM8uSnkjcXtYFKSoxqfq
sv0fD0sU3aDTdDWt9ApXLwZiLsk76PIfQ7+RGDPTrz7O/xQst46X6izgb3b5ptP9
z1+I4dk5wuUE5vT9HQy+McoBRIzN2PCkZ2oPm1x8n2BBKnnfK1nzbsfj5PybiCLg
8rW5JmauLJ7oL7WeXyF32b6okO8HVkCfzwGSTzCJM0zoFx0lWt/tzjYJ+0fq2pza
zvAAFQV4DDoY5cEyhnb4T8f6O2KVHy+9H6oMV3eUEsUS6ohjtLIVVEr9P6UX+pl/
N4J5qYh0BAaCY7WFx4kUq31DhwZLfpIqgrj/bJv4eeSdWOL1mlAwB8u6Oy58U9AW
2+B9Gb7fnxiS4AYYt0wGOdkyd5lP2oskhdkNYNicT3VVUhvvMKAD21mngzX2Ok7U
wk8lO9ZYS38S3hrOSUsL/FTl0E7ExQkQpkk4o4+bd6hX3lpJwI4LjqRDZLV1V3Gn
CRcxgyCMOw6se7c/QokUvcK8+os0+IUeZTs3VNpari2r9R4t4tX0IEBvgs4hsH9i
JO/9P67Qsv0XQUAbpubkqwdZdxkwy5XtxHT0aHpOj0AEZp155/lf5WoD9SG/hsS6
e1wnVADNOICjeVzwvMReittEA4lfvrWv5sUinGvTOHtd7PJzGVj3vpak3vvh7Rmc
L7blyK9qCuGDUcXpCpvAfgl6jSXBNshuYHHhcV6NfYO7c5qjDec8iyQPrq3e9XY5
Gia+VWUe3OlmHA5bqvqMngoaMw0Rr+uamho8km/hnQ3Fg4b3JV4EownJteUZ+oDN
qQbEVcL6R//KrFiutwxRwpSh+/oJPNOJcQszljlojoRSJaC5KsA4sGBs472JZq9o
hGHWFmQ0fZOSQ5DWqseM7K32uWh2CVNCjzTiTkWA8bdYh++gDM2gP1IbGRtp/LWz
xQC6jD4khGH/HY0UcDkAgxykDnHl5Z0DLhWxmn2epc3+DGJDMyDrbVZh7RPbiK+x
MXkVTjIQO/aIYvLRC/IaKqAIpjCkWPUglC3MXY2BPTR93AilmFqU3G52mARD7iRO
lIp7Bekl3GCRcHax96fclSH1CshrV9u7dH9aWcpUIwEVGcsDVKxbtmbsUWnn/xEx
bYtFDNvPL2j2lWxwLYCZPqxLUeSGihed9ML+FHyG5Wr+wE2D3vpHbQ9HlvE200PG
JN1U+fRCQyS20ad7jMQh/R4S8aYvFOCB3/8jaW4ewkaO3KxKSS+iBRJdsav4VACw
qfKX6zhXnjBIrbOHUkN6bXjVF+0tt4tbw/9Nb2BMcspNTy678n/RZhzBrJn2xGyU
w3Ymtnzu4BtmOZaPvdLw3EfOQC//Rw7LzVG4JKI6MKo9LHER6MqcYGYeq5L11nD/
YsGxB4m4ul6fh1E8H0yIT4xD0CLAI6PkwxaCeII/vy1TZo95c6buE7+7oHEl6Fuq
3M/7bDnlGdvzqxzvCFOuKyI6r4U6jnO3xV4QwmQjPmcDlGhI9yM9zU4/hD+88ROC
J2Wr4X2swKIsQXk/SYPVHnpmMVGaKGzI2g+FpAobhwbuj7ALzZj21pz9yuQFasx9
yO3ZtVRn6L6XcK2Aa3IrV+oLHHX0bPethltGIt0pwKLvCD4K6F+pDdRiLDZO9T+E
VEss89ldBBGMugvOEdDngS8S4a0t38rok1akhEelpLe/lgMjo4JFGS7/1jB9Kqxz
gR1UQQZUIf8JOjtBgNIuT2bY/pp5NqyhbDBr9IlBI/mn9Zr6KMxAiLidUJ+hBcSJ
PFN8bXSDsPIFuURlSy7IC8W+nc6iP/6ko45RHCjwNfit2X3WkRo86umLWEgcQinI
1+mDg/d1Cy3Ba0YfVARkyXu+DXQNbEPi8x7W+fkdIbGSWZ64cYD0bqCUe2D7p7v7
2LlaW2xzLA/RyqkC3tDtuzOQ0RVhli5zBwRyGg7aUsfgfxalALtLO0ziYhbnSwWc
3qwpYGHRM2xNBOrm58hS2M+1xUaNkJ3MtjmUeNsZ4g+hNOsgiOUZ03VNuquBszwx
zLVTcraI7I0Zdy1qOzkp118GM7v2Eek979QnICCdWdAahHkEKIgfNcr4EDkHKPeI
CRJP7nPl/rnKpsqSn7p3d5lMNl+hKgCC6usLbgSvV7d5spfaH+qjXIxduVuMMWbo
24ydEMtU+PB1U60rdByxULnTciUKSohpDnS4z64ZSw3IZcoDZfdu7yPa3tEW9haf
UsbJr+HJl5hRcl7SeCTNLEQ46BKUgvRbo9CYlq07K4gqW00m6Qk9d1YUOn2gFhsu
vCbuUMGv9y711OM3cIMRsDQVcU17OOLQUmzTgd0oJzESvI9eA5VnKmX2F8CQkFr4
Yxtc0a7zhgAgjdKOjcj64dEIrLATWuq8qWF3nW6+025uFpGeOFxKpFIg0l2HUINv
971n4JuIOGjidH3qQYTD4pYMzXnj8P81jdYeVITod/NaHHMQtJHTNWcPXODQTFY8
LO4VPnhA7Kiy4LIE1SIjfuS0VwWocPJBg+1vbxZFKSOPx6nyEDpWN5mUeufOva2y
1ab33xoxQBqQV2zNo3wWBmm741NYHQMAMxCHrv3XIB4hUiw/zOPnYTPRDaGukoxt
y+YePELTAzuq19jHSlybwOagFs8u63tuFVNE3ouNRJ8w1qwsV2Krm51KIdldHZp0
sYK5EUhFsOb1UyJTiWO8jC7v5/LJrvYkl8hTirVXBIwPrtfrrem2xQXXZMu8uOE5
4L0dddBzIxbiP9nk2NIClg2KrU5DITAULEV6HDm08DhQf9TDVxasEb8COkTosQU2
3LgoAbTpkfgR/rKwc7WYcykwyowO7fezt3fOWa13FgBbaoWA6UecxbVXPiwmUmTi
kJ2hU5LEihigU57HuR/21HHECcHhA9AuLmXB3/ik5DMgQqlbIAscfEvRl4XgeEkc
gTK1ugBNh+yyo4BJI9PCRsDbLcmXkwEvfmlg6v8NIQHKVsQQK4h/TOJ863vT3s4d
jfjNNf2qaNLu0ZF1Ir6jckx9W0QaoP5x74Q1/FYVRP+bQ4xezK/poBq6RtT1l/sX
RUGN/me4zSuvDoyeqRV2R0dHPac8OaAjzxLrafykOTE9bbpmyJWOArWsMt2WCwKQ
JBH9dxQ6ASHXeUNdsXUth/GyZGti/yqGPie5mSd3je23omqJqAhhUfG/axCVKxiC
DEQhZ90pnWrCSb/sqYvWM2dWpp3uCnpgLRBUj4Xqz8VxqUB74hah/7128HmUGxgM
ElIi6R4Psl+5rsEiS4oaVRdM6GElfOhDGGIRqXEsUw8CtUs0Z+UO9s4+mjrvA+Hx
bqOikwtLEaqujLXfBABRZGtjT2UULy5Do+03BXcl9JosPV2q/Q9NYstStls++nhs
Y56ZhN68kHUdTs8zXkQnzZkwMTpCvilj2mvtAOTvqLasptx4vsFJYTJ7KsN7ZguF
kSQM8roSmoK3zh78JTyImZzuJscOFmyN1/rPq5US6Fx8HskdJP2AZ4+VuzoVsh28
ODBU5fFuP8VZeWFrH6AgnU7P4m06UsEZTA3+6Ts5fOnBZJYqqgfJ9BcwHMs9buGc
6E64FgN7Jn1nc0gkDb4/ZAdi34paLFHilNLR7+NuhdI6bgBe0zKB7RPFofkJ/maM
V5AcktATJAyoyZgLmr6KSyONEZI7jN+aia+4tOeiY4ESirUzLPOKS65M1GU852A0
tf9cjCJDHgUqUqYjVvBzEY5LPgzhtAdip9VgOWG9/MHxmqYAwN0J8KSuIwGPbvqW
LHkNvdH1hJWj/fwjCkuGgo7Gg+ABNUFawUe+61kHeFLGTLayWowc14rVDBfQ9jLu
9N+sAG9ivwrUhGzFo1NYy6dtvyr5Ob3p4t2IvJIfRxLhYxIdx8ebp1UVmTBQt0R4
ZuHPZb83UGYI5l3w06pz6AYnxL9OVqTdblt+59hfU0/E5/nNVPbC3dlqs4g7GIC6
iHDMoU3qUEX6/wQVQp+wQrHJShhSL1LHARHl1ENb0mLxI7WUMksh701L+OT4QC5N
myAgmZLtoCF0DSRcM8NrppwVazvrf1n3zkl9yyFKSZE3yTVaXfel3rFgZEoupy3B
bV2/gcvTYqH1W4feoE6z6ck9+9VgbTidM2OhivFjCKRwRGsWuHBxCxS5fl4IL8pT
CdVn7znOV7GljOoPB7WN9SIhe13XZJij77ZaeXv7Asw+eGA+yCNGLUWea/dI55F2
9Y844AqOCWTPLMciC8IZUtZSZr4mWbWAilvMYqy4ay7V16uGo5xzSK+ltJBgbxpM
VtR8QK1KAWIPMQ3pEqc71wqh9mbpxtEF11d1VWTPcOtrvTAyulGcbwCYVZXqfFEk
P7oJyzsGzxy6MiSvKbm2sXpgq44rIuBmUBuxrVSTJosVyNHYd/Zgn+fS68nOoFX6
9779Q5ZS6LheL6OnOxkb7OtMEYIJiAPVk3GQyDhHkCS0+XUvNGDcfH2XINzDOYhJ
1yMPYYy4YAYwYICe2hjX/DlQe/OgVfTZQSomq4l3kDKPwbvNBR+sGuOyRG+i1cHq
59OkXE85UtHaoLzJ5hzaq3GD1qq2kcXbTOytruq0ngMlRwf+KXZai1avedxJtpsY
bpK10lBAsHBa1ETcVIxQNpSQdenytsYQsEC+rc00/oG04ugX9BEnVSo6MqChkypf
OSaF480ma8ZVk8tpiIQ3t9Jc8XaZUuQnXG6MgOEimHsg2MKOBUuLhlSW27jHDJ0T
OY1epQlBoEI1ND2WYqJrfFBFVUI3DgJULiHuKCePaDRG62PKz4FWce5tfpebhjzt
wogyCsK33MnjHwU7ZqE4DaTFa4KPHq8JkAZScSckNWcgNGXXqLWn2J+xrMok0sjU
qkhUQp+UPfM4Xu1T5UYVyS9M0Jt6wa5Vr3mO44+3sEdXsCADUx5UK0hiXKze65so
SN8RPhUTEIV/eYHO1ABY0uEomGoRU4TdRSQvOsWBBrs4NZsrJIwy+TL07kdiDmLO
ceG8NRtu4Ylt4u7F1NBSormdoeTvV2izZUpE9TuJheov9xaaJD6RfDIB6TwQEvjT
LLk/smTwGUC0beu9MIteLN25Ov8twIO/bRjTDXyggv8sRSFD9u3wejBDFJWLRhQ0
BqFJWZalTyS+nz08OwNzevAy0jJesOolfYI2UJVJG+u0MTUgTVqw10gBdirQkDLI
MUJ3VUAy3uiZOYR3na201ZTk9nrFFFsAJU3TgjHx66tcYY8TvFsHx9ST2LlunUfb
mxk54jMui+It2yI8qvFBZs+ZMihx0mWXsbnwnzNICduv9apKlQKxM2YmF7766JtU
nCjJ6rgBcKa+fO9LuloM2W8CZF+NHv/GQhOQiTEaIfFoAW6sz/YOTK1rRHDVEEB/
WKjfj7FUWPDO1BQICcwdcN0uQW+YGrRXtyta9gXBSWHlXdvQyX68VV7uvVYFLAID
gWPnBkC89ECFqne2IFX9fgVKQILoSrBwSKKkPJCwpopqTiIgjxlLGA4ekdV9zxHl
LbEvoEplfa/X5pMvSVBrLladJ/wggwXb7EBRBIHEDnvQ9bEjJq6aL4sQ9+N8UZtr
mvf4tCrWNPmugvoXgD636HWSqh3IkjEHd8QyuNQWZrhpBttRKLILbytsu5NieS9G
QWSwo2tFJz48mhHcPpSUIJlsGc5Tjdn8aBO6G1AR3v8FtMKMM005n9L1oBL5mwmc
rmW/PKLHFfKYB28I4H85epUslDRzIGnvBdARWm3AHriJkZaIm4sXfm/p1kw0scc4
CL+SGKKJDVcMga92Mc2W9UcqMY8DNl0VHoI7J7U9sfZLaPUd1Zc4/wBeiFxoDQ8p
Fa1bIsGrLegiWFYFRi+MGUbtW4kyvsmYDxGQ5mCglX9ltCsyeg1gpkuT+lcB38aA
idRhrBFez4KUTNTv7EByJ+1+lXN/9xA95uYNVKJPNMhb75UVS6s/R3OBuO+aJWNI
H8bFIgfVQRM3OdQqwYU8yDsBPAf0/61EMQ7uVOigr8Higkui/LMhWSMCMjQU5yZd
yOCrB9EMe61jByGSvySBcdJK/DQOGeHgFczEVxnYuQXAVvEAV+FdqAxcbs3pwNSr
dBgUxTEQegDPRhCD5S02FanbJVjk5vuz5rwpi11aKfvYMJw3RGgpw5Mhmg5BpfXE
+3OIDKNV26779WpAG4IQ3tOONcwlb561jUmJUXAGQdGyEM600CciHkNiuh+wblST
qVLdo8wBYV4hrVeY8u5XFAOCX7ZBWCKzVtG2pq2bQ8JRM5Nw8ToXWA4SD+4buV5t
1dHv0LmvO4dI+c/OKeq3En1EpyRV+VGdadByfdjHhQrrvtHFn+5++Pqx5TH0ViI7
gGco8aOmNFkgd1mo/fSnpDCYSqi3SJeXIg2IJM8iWlmQhhBW9l0+Aav7HTwALXlw
Xor5as8XMgbAkPDyb64tZtQRlrv4HWj8gJEDccFGURHfAsoRFAu968UtbgrEqgs3
pmHDoqXemlpqgXBaWg1U3HnmQXQ4jrjGzw7nk8r2aGOBhk13R8PZjLjFaGZUSjNe
c9N7rELBosCT1hCiXjt5/kB4FThATNOwmnEkCyOXWlUYnpjWMXBcHmNhFBWW5BRJ
B64fRTkaKDbStVIUDECyqFStYQhVz58siGhvMlTvMvm7qXDQNc/hhRRIBQLyDul4
8W4tf178l93IaMdm/4k9VVJyEDr/hSj7179WNOiP6ZZxhW4v8me0HU3Xikkxv2ID
tnMJWEH3kRZjQVbzHRKdpmoKqX1UtM6KaLz/ltuW7r5zcQLABJlyH9Z6XqKZtZU/
whrnkaoXkK2RjZzcZw3cadielOX/v9ghBpf3IAUffN9qHfeOyCRg+5oIjyWeJ2tv
4kZuL0k3yJb24n3D/yhxn0IAAcMTWAt3tnjCqjEklFEyYvtjrucQYQmnJOv79W42
jkFLaBsa22JCpnX5Dch8ZB9Aa4XZP4FXdiVv/TdE1oCtKaaA1hb8CrvI4aOQYP7v
ZwMK0WL2vck7KASL9DuVZ40lBbfPLhqzzTTdyI8Ibr1dnOgoXVaOx0YP0SNpGn6G
joznbZybkAIvtDrpWRtG5ei02a5LV4axPKoDJKespyvsZqi2877p6YVz8At8MLAL
JHaxC/LyXGpeb9OKBhn4NY0PHJzOeCXd3CJtR0qgfs75v5uCH8ZT6cQMPtbLCiyB
O8iYJ8SO8rvctairVwNJ5NacVo967bEnlRNFsDWxH5ikryVwi3TGNJA4PHtxLRds
izYqnsh/Q3GrQ4oBMy+FApZg9PnB0q/roaUHTliRZ08q3rDN+9PVfsfZrY9aX7fk
ULmqxMitirMn/nvdiYZZqnxDVNzHiRvDCVbolremK9SUxZbu8I79+X2usHyO8TEO
uKqYXklb0FgEV/xNh+M0JEHDQ3UOlwsz/F23NEIzXK+TAsDts43lhtL5HxkFPH8H
nkFYvxIGmHqLZzgUo8j6k27hy8d93TSKJsYTkhBXJXCENUg6sXkJkH/F5KMdGj0+
SK0FR/1lH956PWDp6PFS1LdF8IFQ6qJDlIPlFRB+JbZdQJ4DqiNwEcawOufO6fi8
5iZ8GmmLyYauwGulsYXITSCBEiJ0lnimyWrLqeDLWZduAteGLw181cb7oaiIei7D
v+DomZ5T+MTPY+Pfh3z6+lbnqVfsjVLmmrXWZ/rw5La5bIXuZVMbG7WCi6NJFrBp
gqiyh0tVmnyVbYx8Eztzj8QSzWXVErDkP0cesjpdouFfNFKRCrxKwuUTrrLq7h6n
pvxtRGA/lT4+H+NYHMtPlPkqVoRfZIzVrkLpG2WHeThMHYsBh+SwWVjUZcXyV2l6
fe8Jknx0s0VL/9CCiorjYB2HJbvxG8Yi5pwLOvu4VA/gEXf1cwrcGiHEcPNJEXj7
AIa/vLMtu4/CtpGEnokcgl/wA1EJ1hEZDq845GKulqtlcFdqZTenpCBqe8Cgpbt8
b9PhuRU0bYi+SejT3qk3x8yDJPiFZHprMfkJhbPobkElPv8ZRyMZcmPqQWtI+CTe
pKm6aBKBZy7VCySyQsEgsN/Tf62Ht34yhdFqTNUApFsMB0QeTDANAMhAuwJTilVA
4dqu6Iwe5Y2ogHm3l+xYbRNRSbbwFfdia6OSD7Li7jjhE5O5KOaozrZgsNvpJXnW
zVo5xda7w1lRz+CEDKCzbqO3xr6ooxxTyNSSSVCtgl8Bk122oUVQsYtV8CtThD3k
bfY+c3DAoF2R9y6HBeh7c2EAjAF2Cjrw0mPTOhMTTwL8RKbKy227ta2wijewABZn
9QktOP9e6Uvu9rQoBmcGBf9pR/dAbG3XKO1s9d3zQ4MYFm7MEkWJyqvADpw8L4hx
qpew8LAAldmgui+ctGJE+ezzcLEhTG1ED+Bu7riNGaygLRjEh8u0NXtW+j8SvjlD
albgwm9mvCztbwvmIUelZCgqCVezwAlhY8NifQdl3q91LnPoqA5xMOSE9i4PoPIG
HNnmutDFmZWTA7/tzAbBLZv+rQyQZkTAYGJFTMO7y0dbV7Pkn8qk3CoRNH7DxGyn
jQYCUGeCD2mq7UACz27n1t1E4T4MvS3g6MwZ30Go2QQMBlb43ohovSjWPwyGVhrf
rtwvcM9j6OJvoeNne+6Mcc0c+VtgUk4WTQ4svsJ3pqzJUPnmzZ/qRbQLx8n8afT1
VmPH8paOowHlNvKYwvTZZFUkMEiJi3nNO+fE+XvSu0FErqPSkTsmoVJec52sVdmB
hmwbaNBNlIeHOkFGAxpqc/NhID9bBuNxgaofsN8OrUve3rYXFj7WjPNMBtc729YQ
E3kAaHbhKxs9KCiErXd9Iald2tMZ1c4j61qAkgAiRmGW9PLsCE34JXdmrfPCpyOv
pQzJ5VK8aeBrDiW77541JDKD0R97akDKAIWYYVi9O1Wrvi6c1/DyTinVn2myQ7od
HwsiVMd8/h7Eevlsh0jtqv6SsZodhI7/UBYOLxkJ4h8JZ16Hw+3DSQwj1MYHGGUN
T5k5aoffdAJ13C7uTzGrKs2JYcS11sbPMEOP/UoMPgWlBzafl1ResxKcjDntp2OO
1Ip5qUO5Ah0TPx8iXLaiHzNhG5zYtxpEpT3C+gmofM9o7bz6VkBh4BkTUBoFtWV+
BlsfLmoQ+lt/zh+hHVe7x7/ajeM0pw1SFi60w3ZnmjjCPVNCgKT9IC2GQjDxaLBr
A3nm+4C19Yg/K6+psCaYwMWa/HTIGN5fbmb9XNONX5RcgM6+PQS7vqb+JyTCArZ+
DgwDVEtci/5Fv91KjjF9md+JuIyd2uGijZ019SC/ebwVxWbZ/pjiEX9yUvIWaiMK
j5FseVvgQ2iINfx9AYPLypcaeNuRU+XPrPw9mc7zyj8aX/b2b94APYx0Dm8HPAhA
5j7FtjtN4fDj+kJEPNKboRN5fX8Fqg8X93IQhVKfek+lSZFkG5WNlV1MtmRNsJ1j
+Y1GyMZqseEa7njQ9GfUQK2K+tNuGfNSmDpUo1tu8Rwfyrc57QQt/LG4Ahr3vkDp
dgIrFRxlPFayXE2FpYaDXt+U3PW3ahQfAHDeNul4Mvzx3tY35TA35+g3AR5bjqJd
OmyaLtXefNcxHDR85xPDCuoRBzPuc9q7xFm3HQq+/TH0mVqVFViS5JSi1OqKAezv
c/BoJfEYkpH1pGN/K0xk0ya5GhB4Ly9C27u8C96nDO1kXRTWB+u+ufWV2uBNxtz1
Bjo/5nul+T3KNkS8+p/VDSppK1Y6py2fl7XckaXro43wNaWhn+RAKstd6e+79Tck
zQ2uItaBS6MW2lMTMSaysgfiH1Tm/RxRLHCvxE+aCC+ObfZHOnrwBR0r5s09QgY1
0SYXl5FNkAauYIiRFxuE9WzZwIRZdYejWUDp5FIxzlHKz2GQUJ7FKbEK3R+oVIjW
BvBARQ6ipBVEveMw9ZrZ6FBUg/+jSlbe9l9upclyp4PQax8dXwEtxGsh/7ruUMQm
WC2/mtKVGOoLMOqx8UqBipfwS1W45y7Zqt9Ht6KPi4ujJ6xC8jHKaYf2pGdev5nK
HSNbVNIfw5dgheHWlRHOTvyoDKbx+kNPFo8l/8VN99WNX49XTlt4gAVnPmMetelC
xNcZWSZTuORTD19ujFp4fguOxcitGd5qhpBvv/XYCdUOp/FBqBKOiSEyWFCTgviU
YBEV6rcffUMm9qBmtHjfXtgoqBN5mscMdwdC7GdDVUDYAvi3prRye1wh6wPtsQPm
oGCge/SVFgdGprOQsmTNfJmI2qmxUSsRBIRTnmwF3km9stG6HVcHS/ftwgzWEXQ7
y/07aKeOKVFjF5WXFtFiveSq5DFwlDwDKIBmX+ItFh6O2rExhHXawEgg2XWv8+bM
qDZn47CK1gWGWk25SNfQgD8G60DfaO7AAYe6MUX3/M83Hi9etsq8RU9FMjZh7Cos
cdcG/wXhMCu6gs6gRq5TT5qk2R2s0izd2mK18hYuhqSsYLhkb/UrZk+m8SQDSI5c
BZKq6D1SIB0FxyJtQYGZOzSiEF5ezb/MT5RJarSm10XGMDcfKp4LaWoMY9joDNz4
TdiOEbJ5UQHtOspAoD0I5dDQJhjgMRvVLuZHspQqek4Pz0TkSTFykXVU1vuORT4w
f5jN55XxSK7NYSqOxdALwQ06RyOPDp7c2249HDoXRQhN1alnQVLIL/HKt59uy3um
VUWadi7PGPwWQY2wjgujszZcw/E5yCJkKUPHCtWw7MmveoT4AfvJFN/8GX+BWsDX
CphHa006ZqaS7SY4kYwX4TeDBjXbBJgWSY9VXJPLdzSXxeA/XsitcP6HZc5sJfFt
0rjDdnzCKsh0qS/liwOyHP++8mZSO1V6cKNmVejMcFVlThzMtyWub0h+mGwXLnJO
50tBFp8eMb0X0ovUTPDPn+9+Ug7tMWBE7L0Zbqzc9EQAnASJOyAT0WGs76rwFGUz
zyo7P0QtGJdieeI/w/GeFewav5I0jc1Q3ZVDbq2/oYL2oozDmBKvVPzUyWNCSJ42
vm+Gtzj52SAwk6K+qZrYjfEyrj8TOcPwDWeLIuy85TKU3X5WAKssHKvfgWnOkmNf
8B12Sk2FruByotHfX9mL8velJ4qpDjnBwOR+5wfl2HH4g5eQh6FZaJLdqIU7EyNa
ZlcZlhyJKaiJ7upeV8dlF8v/m1pmQXbnv2fiTTYdxDdLjuE1k5zjz7UDm4b95piM
jswQ/RIbaz3BTh8sg0XVjyw+yaidyVrC4UpPuzCrynRB7aRZY1uH4/e/aSza5a+M
4fopJLMN1j5l4b1sT5T4npZfeIrjRFZo2F0dFna9rKcIIGfVlf5f5Dtc0ePtls/d
iLL4GyYKrh+cjDe+uUd0JmBsOgS4uGF8uOTEL16Yqta5o4l6SsmO5bHyDSxjBDOC
9NOIlNrsrG/iZqvmL/8N5lI2Yramqf+ItcOpjFcs4oVieTLrA0TBPQAbZ+2h0MH/
C3ItRoHGUzdmHKOEpJbLJsooRPFz4IV9599ZPuI5OzYMLgSlkyGW63CcrYfgOHfc
UpVgiJAY67u3/fhP2JGZyvdcuWSwcDr1nVOxZNKfg4AA3sxjNETA23TOCY1MUE7J
Kq0AbsT1dSpqNans9vTHSq5geabO90XDaZ/gdUAD1WmO5g1wE+eXo88VwmBelT4U
oBP59Eo+6o6Jo3XXOk9FSzTBNMfpv3LHg5vAWKUDfuyXzWHlpQ048gNh8z/cXVih
00CtcZqc2tk+1HV2W9DB2dMzLuQnDnYgPOtYFyVRx9g8VKFQVkl1jvQfVH7JJix/
63FJ8VEEB6LpUHSaQ6yjfpJOJymnQYjsrDXYw5Q1d2f+fsLKYRBOveCwpp2gbPLR
coqr7ziQELLtHNOhCYjy6Ef2i7FvtVDXRuL52/YlG2qWThmdkBhgpH7tLbnf5mBC
8mkTjePKAzobfDdt3RbdwDc6in39xXzEMN27Kb9kPp+HITXnmibxFBqQPxIX569/
5qt7dAY39FBYglISZlK7tmEl9FGblGIX6O4kLQoBc8YjJZUBVkSdQAQ6GblXlRKA
oeeSpAzvBFL7Z7XelqbZiuU9YEayxOkU1eXddimR8XiBZWqX5I06XD8mVg+Pt3ru
SPcDeSBUDdj+UG7S179ferBW0Y8rtB2B1LnWPBwhaTQP8uEANIFia5XeqzaH0h+P
bCMdBea+rEmLp4ZDECOB0IWCLQ/oJSZVX7cJTwnSUVXnsibVVXBVkKci9Z2gAwsL
tXd2J0sdCQscYpdV9hWU/Fhj8VLNAlnHxC+mgLVrrXai/wd8Bmmu6q/lrcSlRl/f
cT8VqCu3i4c/G2sPAdcr9qb9CyN3tGotGSPM6okXHHIeAKoZnX2w9Y0DmNr/pSJx
QIWWc7Pj4LQuZ4k3F8DNSVzypeyUHyBGECOwPtxlBNYmgKOcJcl91p36zaWRCbIG
wlVHq/+cRy3pHef/TFqqlXOGqOLCfVGFcY4aWEIzmU/4Bcv9xPVkSfAGSpZ/3nQ5
3FgqwfkADyFsHDZWS2BQ7UUlYm7CuLn9vo66+53cfWmSg26V5bNXTA2P3mD/R3oO
Ls0W5qhyZoDS8SDyPqQkzZnWJLvX9Hn5C8kxuTGvJk/mUfyAZ+1Fw+KrXRvEcxRB
V2K7nSxQjQ0q7Arc2I0plFmYO2h++ee47TS7WEsc8D+0FeMQC4CiLZEbHATmoEuT
TQj8g/mkMdY3UsLztiJ73VNtf8K5iTb94wwLsd4beGHEUwN7ncoYYGao0yl6Rhl5
WuH2EiC2G6rK3IwjVTOlMWm5+r9ppZOOnwv7oOgn2oLkoN2AwGxE2s4hEEbSZY0p
QvUaMOrgYxg5yPqCvTDZC0k6sVB1wDvaQxsXBPUnkMED7QOugZNKfFD0Vw+aUlDJ
yZlVDBVPUBdZUXgBcFcMU2baS4pvO5ZN8QBnrHBpBg0MUu0gAx1E7Y2GWSLMuUAp
rqcg15KrRYtsYvAFVhSS+wIwrdLhp5KsVHyz4b2RPLkGxYjdlX2vAhRYopI+RTM5
q073JiFjM0LR/POBntGX4uvWYXUj89Cmup1edxApRD7ADHfruRlwOq697fchMOnH
uVrozMOgqz7V55u/db9SI/82KtvE7K5mNvGnqem5XQV+h9vmS0kFOs4V89SFbwgY
5MLJYTl7i9/t2JTzW2AyreiwgqjiDkFtYCNHHm/vAwDWN6L+TBXuVh9YdGQBQ+Zb
UU20vGJtt6E4DW1kuuKiUXEe5SV4TzAnQcvt3rdbHjgreX5nhu5nLCV/qn19CbTH
hCNKiwAD1K0nuDSGMPMQWJXAxv7UMggPMRwaso0C/sj/vC4qeeaE/CmVJKgkBomK
xPbLfnI+Cx3HKOPLD4oB7XgLlXgEX98phc7AWIGPb7ZN6zPTHzv9Vohnb9DpSFG9
AaaiStUG/xY4XE9QoMy5LclVwKETysb4Qy6gDi7avKV4v3oXJAiF3isVgWPjIdOU
X1bRzJBZK1QOumkgX/nOm++MJaBeNJoU3loYzJL8KNNX4JKtviLWXsQBVpyl8vtC
LT4gm7J/2nXaeeSChb+SZqUw6bJdkpFbtxpMipbvvtPC5d3+pIhmpeFkOt/PGFsw
lWFYVpKEzZkfQR5CHoRgO8YxFWY+4by8vmQlgiuID3pszkDQ9McC9A82nJZvG0SU
fIxpQpkM2aDUQC8y0iVUgRbap1CVr09PPAexBuF5HQxj5Z7n9PBd0SuVnVcGcLBK
4PzzPfJobWmUqMyMkJPo1LQuy9i4clShKFK93NWiFJ9Ysqr2C4RKbLXcCw/Q4nJz
kpCLaDwN6odopeP2nEyOxQB4tNK9Racsv4wpXRfwMbi8UuqGsIi0inItEoxJdN6C
v4mXDuWd7wgtzA/mQ2MYM/loBK6gCpUMosfuM41SLngvzCaJlyFbAl1rvspdL0XN
Iq5NUjMYqVkv5UK4BCX/5aThnIj/HAi9XIxRDlEtqrpXFiXZB9ZIqxh3OYOkta2z
N/5VZqnQu+dv5OMI6R7f4+rdXo+EK37GB2X61Y3IjzntB5CpZ6G8JRtsVVhjaXPY
udoIiKMFVRn2i8lhmbu7nRy+V8ucYL2FfyXHOeAQH0MGQ5ftf7bSHJ2GndNp8r7i
KMxfwQe5O19ToAPMIER3D2B59hdZyhfklStaeVL/pNubXWpCo7FjeViq2LRCY8VP
7egn9faDFz8WCRdpHpW1tJc01qIkQXsvSbDJmcExc+mEQby5cPTAJBDz+xBvQn6E
Z6QXZ0ujwmZ5VDLwpaHcXpzbkaQ1SvnMhjikRnDRzCmL+d2iIhhZpLDV52rEHK/O
wxqxgrF34OLqPc90AyNEyOyCGFvgXIuJdbnl3E4R7zZ0A90ALnU6KePb7fWss9Z6
AYnG6BLU2olMtyq5lZ+IhZTRnT4ehPtRpgdPv71Hhfa1JBmHmZEgEMq5EqaJvnKf
iRlVv4lVXaRqXAAzeF0QFN8AoNlgJiwv7ye8uFz0ZkdsJlJrSJBEi13FTO4gFXC0
V7w8/GF9dvNAwPFMJGNEIU4ZVyz9UidU6nPDYxc1LsJtpsuf4/PqooUsJQ82ihL1
5OZNb8pjXTBTZ/WIQR+4tqp6KP+b8P8plQAlf1H+VAGS9J9ppD+wRW3zEyuJo9OX
Lo9ZoxwfIo/RvMg4IqpvkjM9rV3Yn0xsHBPco+gPGfHVwHZUhz7X9oUlhXEq4gUW
Jxw+e0w9Ni31DU/txbztsFA1RwOhHjpvPyDjxvIguO/qrMjH9OC/DfgwBbddMUy8
joL+DjXqGKh8cqpEc1MT84wAXsJB050KLkPu2yhwGnWV8MmhUmPzn7w6G9FdLyEE
DRby1oI+IUT5B5TB9QUAGaMVAT+1Wo8Ytr6y68kDGzlWyqUpUSX71kJnMaogiy2D
BfthGU9kTWGKVivWuY9TFh9gXqk9ubasrqZqw8KbBbL9xd3zOvs1Zi1VI8PtdAjr
Fjf8IAmM2RvOWPVAYyYj9VGY5niFpCYU0u2yUegKkiufxwZ3TgSD6to9TEvPa9sM
Rb4/HKxFJwjhLkxx0F0OqZHj+gdNYWtD0Fjg0FC+Uo0rMrn+6JnV4i8aEBA0u4tI
MOgo5m7R6kcDp8ZUxtHEqeG53jDmMM0mH+53jffNK3NbKRp9D9s44uP0/6qMacQo
vlx6KDggXfu+kaw2cF3GB6EIBrXbffvqmBngd6OihBwQa7Oo1+oSxKkznDlp8XNz
7U31uZWSCjF9JMg/IZnfJLR8YqUePf3nVLhCpyT/cfz6mxar8OKd4Sd4wf4SRuN4
eioCkbtQs610OhoKi7FSC0a7Mby9SPL3njuq5hzBlvoc5AQuA2B7gehSRTxKxz+l
qRKuyOUEqXgubblpqucv2w2UdLVkr6uUOY/D4igFe6X77s/sLBIJwW94CoQUI46o
7Vje8CxuNgp0z57EFzE/meM3ulwC0C5wMOwK8/kiOwY9tu36bRULh09dWUUdaTys
uY1syqcksEid50ujDohJVt68PwX6R9XKOhSjvBiXCfI6k8Nx726v/49o4IfRjcEh
O3fBTCbbRrtBcbmp2yD544lUwmS8hljq2zXjksrxCimfIfO3oIknti+s+fO5j5Vg
bfO+HPpu/zeBzCEfuAus++PcfVEtMut7f3waOYpKgoSiUgWqask64svBeFWb4BLl
PQ4gA4km+WMCcX4F8lsd8PJfSq1ADoRsphaIA0+7gV8hrBhqIvAI6zobDu1NoIib
x8t8jBqYDivemh0p9BLsdOgCULE1goft1xhbzqzK17D3qcFbYr6Lav+vKQUURaUe
b+jyOdOY7D0rUT1MT+HEe0NcgMesC0SjaC7YNgX54ojhT/dGoKISlLGfGYtxX9AQ
j35/ixxO7f/gyoShRlBJpTgyil9GD9NxO2e1lO/UFDP01tXZcRr56bOMNvbIgKvf
560/3PL6ZUG0q0NitnOi2Jx2dP9j8lz54xovBO94ScgM6yewLdHe/pkULYVW414g
0pShNWiaCMr2COaMYWzB/uVrkNoNImuUNeKQ7xKccQXUXz3sl2cWBRy9/T9+G993
C58IAnnEZCXYzQBdSIRQqhNwpGoiWqErXhkBwRPNZDEH/uuszP64PlFvwpv1rDQl
Yrre54+C0IIOlxoyyyeMLIgKwqEr6/LYS7bMIeBMoE5QrmuOYpu0wM+EzP5p5lrc
urcjP6DnGPzyRNIDIr8yYLTBC3LbBv8uMRjaVykUd5W6SQX3YJxfCZAjpVrfx8bV
LAFGK54jwpiNncdLErmjVcZlF1bp6OzJ5g/3vc6Qe4xPWTZfV1ZR4j/klRQ/kEBh
3+mh995Xjr30anvvNCFVZgr1Z6BBQ+Bp5WRzwAfiUkpIYI3kOI3x3C44E4uRu5HM
b+tLVKX6rnRpdNkWnqbQ3XQSBQwRospyJr0rjUwXZFfDxxCV6DBh1LN+BtqXCcxa
I0v0FdJ+9wE4JflDHDlgBSFTfY/mECJMsSpTu9o/gxgE8w9Z3fuoc9q7G9Z/sC4b
+1aa9LdBlfRt5FODBHNN9RAT4zpnSuNjs8HfcjxFdQqXc2CgceonKaA7JHkv//xh
ChIBujDY3V6ndAXqZk0ZZMmmLbajRge9tgrTc5i2aOVLfGXoCIRMg/IGQfuxMiX1
fr7o6HoIW+8Lo8+x74HYUcGxUxwKU2Tvo8VCVPW7bupNGNzFxg8FzIoPqfSbZTsO
GJXD1fdlW/H0FwLZy43u4/YGBiRzaWIFhk8mWZJwHp7IJZzBTGi9DZNYLuK7BM6s
KbhzCo5VsjVNX7MqnICHvDUlaNox43aBGezHhl3wxvutPDHrGOEa6QadV93aInbq
SeGRBMfOm7/jhj1Eu7Fa/h+tllLlMQYEegwJkQvYbbS0Oxr/1u5MJ4wWwn25qyMQ
PiP+Wn2VVGXpz0Uyi8QDX1/+03d6/WL1pglB9M0S3wdByuVsv4V+nKz9Twudr+2i
nV2/agiiE/zHkljvTZ+2TONkReMsNheI7rMASjyDzTvmSL/x/B6U7Dzyp7CObSiM
ul9Pm0otjR1lXBDusZUXoOZnPiZLjj1et8Tm3ARic7wQODNtnRizyX5ZmqGN2ZzC
GnDIt4RDSsK6Scjt9k0xEr4xkTQjGAD1vySStMs/Ej573cgIc2pqZ5TEz1QrRaFY
BHRe8rDocqdeoOZiY3U3Y0Dq0I3UuyHrO7VOXYOJDWXoMuAHiJBZlMZXhe+rmYgV
HepMLb/LKOOkAML8efG/TaK8zssIObW3ZpzefXC6rdlMchA+BNOxuswRbMXLPROh
/SljEazagxl98zfCMnuQ/FqwBTbwrT44Qe43vLdb9JyUDbZYsjpEtD/iUDOQZ+PE
daXeMoijExkeOTCSZV/KSdKMIBr/jwdknrw01X9InGGQcJ0FbMaoE4mpoCcT98a/
doaKT7pnU8C0zuYLMBy6/PST6TPzQWegnBZT31XOgs8VwCn++V3yrEHYTo4TvDBH
40nO2E8oTw7llPw1Q4dauv/Karj4EZQR3BZH4mdqBjdLuieI7+Ey6uzEpi48n4Dm
UgozqX4KOTBA6JJv2Tj+CCMOXhS3J1yO9HLx4doOJwRDlQpPYmktOt8dU/YT1LCQ
YVspl88VFsiGPabH3DS+303CuitqnXI9/koVWJ/z419rDc+EumtJYBbjVksqDpeh
PHpHZPzDhpBu82z+o+69i1xgbx70ep36CUefuvXh3OM9pKnFb/LQRTpIsj9H8Wp3
Tuwiyzyp9ZZLLSxfnHBtNkrLelgeZESH4SCNujtlsmr4M0FyjvTROBp4KiMlMqYJ
ZQSar72zlB5NXfdqxEBJL+YveEobLSAFCjezH/HClvm0I/1t7nrvj/HeY5KjITX4
zFs8/jWdCgvHs3pK/jbsocyyswV8X11t6uMiBI0e2SHFGQOYTuN5NF0xXHeGbYfV
AKCp88H509vichOqkVXCvrb/9ehTwqBuZgCctDFOIgC2bB7dpH80oLSkpZNjX9Ay
S4bXsk/288yW5z+d7MUbARgyoThWF0BlD/Q30h5Zg0e3UDw3cX7HEgjXr+WZlhRg
+mFGenIMkYxt9hJeNmUz+cJVTum+5DoNPe96M+0UP281F088ffV/zVSeKFnJb9Ph
UFPM17nGvQK2POhH6qhmhcQNc0TcL8G1cgwYbT+HwkIfSZ6OR/NVMxz/zTeEOmIN
a2O9ZLnt5TrzuRTT/z0MBSVgeu4L/ApRb3LHThRx4AX64Gxg6rykrOuScdjBC8Fw
6YNAqAyrbz10j9gZKQ6EtndQZwrlY0ubJWkXRMTiMg1vrsIIJbiFP6j8Q0PxJMxF
JB6aDf9atzJ+SUOxoirU5dtksuUwnoIDw6xmUilsy0IXQjdk+ybXiov7mm9H8bEC
BncYFFK/KeF3w4R3V/amttDnIv4pAJXOtrfTevpbCa0I2Fcz3NdCArI8r4W+Z6z+
bn1qTF52GreEGOd9esZirLroc+MCloqtHSEF7PE86LEWBNzi0BaAExxX+RG6LUoM
3zZoLyNqrkQsWo+HmpOVaOSG/yxlNPaP8JQCcFYfJADg4vNXquaczFq1h3EC2N81
sb6ZyNCIdPv4If0vEevRDdl0wLcHdfDSrqDNzldarrQW4+wnsZ9TUr6VEQIIoRa7
7iL6QNbD8c1A7+99qshWL9cyBgRAeaf+ujO5+n/WnKH6tDwmMD0pqgttV/rXbczM
i4G/1cn/jRDb5bD6CBQ7i/Vvi3fH+3RvMMYOQzjcQD+AZLGfQJgjiHcXN+NCE0KQ
K0G2TWMDEzoOgriH8MseRx5ymjDnmL3v9MQqTpU0hgRI7hGIObuWNRl5j/Z+Odod
2KbNn75+IA1Munr2KYPUGKJQtfsV6TTvjatFByZ1c9cd9WVaR4Lk6DdqIM9GwdV3
zgFdf4sqo7+jLEehoOE/wsNO/vXAnigZoMUV6Yn2aY5x6k2ObKrA5spbLRPYn7wM
tWCoVjw/NFdiLwDptnH8rXdcqPWa+rcWUDMPGQtLIgDj9bhCnV+w3LWAzLlC6FhH
yftnuPzfpjyBG9SZsgyGEQd3EKFWMWM6s3Oz2HUbAsSoELlxMtdw6d/TEqTIu8sr
IcNIw6YcbFiLey1eR1gw3DuqZnIq2VAOs5E5OsXC6VAzXB0IxPFFUPkfl/mgqiV2
/oEx8gTlsn0gVsl6luqbDg8I3N3zzg3Zm4UABM8d6l6WRZCxfigv3t/CZiuyPqhG
pPswA46QzQYyUEWm0a29BlHzOgl/8ggc8DONFHeGDxfAFs561xVbdkQVLj2IaJBs
KDb8yVYiSK8x1ZTHIRqu1+J2pV5WdGFwpWyUUHYcO2EkDPnSx4K99SXzHEwlHzIW
n0wEKQLipsMJcGveBlFBHxISZs/ocuXLRMa1tBQ2xqsvn1dNCeG/zMywMkYm9iKm
jH/kiBuwhLPE1HiKEFD++G8zfgowMtWGISV3LKsZDPvxIct3pcEUNFqrZhuVwI+8
XaTdhSHO415wdPwM82R2dd6hmjmbPmskApZ1Qj1pK9RksK7A134JIzz+LVhv7c8I
0jv3j05CAFH8hUAsJnJsAh38OxIIgM14tRnVmb6KEGIYSkP79YhtCj0kEwNXBhRE
gW9Ho1sp8JzGI4KqLFuU7D1kIGS2SBK3pIsluhB1rZsGz/EP1MgAQMZ6np/LAHH+
NToBgxUlXH3HR0VvJzJRQtZcxd6gPX2EJF3mQB6IL26KmDQ4FnIQK+XjhH2tDK8M
4bRZf67kIe6emNtkD2HpRhNmuLiJa5drKsnK6lBtbq3AweDSc2ZA8F+jttjdf1Ty
FEo38Nee8qMtVNWovc6TJq0Qo9+3D2AmJW2reZzBryAQgaNpnRE5C49T5vEOd+dq
PaxF9x3OT+UeAzv/c1d1BskudfQcBYz2OscYsB24NK1sTLffaD9VTVdPKrhEdBrf
ZaEA1nn8buUQSIFGX3IgWLwJ9naBLR/nziBeGj7sxz3CFAMRrpphQZH/8GgjY2Kd
QfnEeMBDGQtQ2X7ylvT0zPVQQtzY30l0vFfUSLOvn5fGfMNdNK5FyqGG2I3cU7lm
8oHSdISavB5BsfJEGMqiqBmdnkPCjhYzk4N5yvTBL843/oveGmw1wTbmOQlC/3N3
qvvzLU8F2JU5YvTd4LV/WJQhjR4zgfen5AhaeDTruJJjDubhY9lpORbYHwOFak6A
b2YMUTtGVWfV3NkdFkkH+HIWcLdMdwNCUmOf25Kq+f6HQZhhNhPRvgeS063c52Mn
V5InQqG9PQKoHA8YdnTS3QNz2vQjkhg3mHkLGe/4V4t4L8pQiEv3rBQYz2mNQlBK
DFmL6ART2gC/+epkM/QRs8hYbQbKXzZCx1cLHbbW/XhmfMnUfhcplSdgdNip9hkW
YktgVAnEMRdzAFq3Tjh7M0od/BbHAt0cx/pp/PFOGetI+BNO6rE2xuVMDDT1MLRl
PoT0xi7kTv+CWFMmxyO0SFCtWgn0gU8GfizTyq39vJ3JN+J4BS65te0R/YmCCIK/
WLT14OSbc07wpbae11QBw/wiFvoQUkvWZK7t6XvNVXWhcqRQAOECtmwkkw8EENzh
0aE6ZfNhwMa5JdlAOKpxX0wvRzWplbNzZiMg0YptGXU3vu7Y+U8QXgPV4X8EWRn1
pLBPvNzBo1JMDNqTRfQqfTlvghfDPENqEXWqucp331xqPWjABjiKOlpVQ0BEDqZO
XWnB5Epl48z32dh6ZaGc1bnGaOk0Vcm5hiYVkgJJtfcesaBspfxriptxPBv88o4y
svm1qIy6f6lM81V6gwea6iOAPkleykhHWZyxWUqjRmMMy/WCLuata0rtbe7hQrKA
w3vmwwgavX/lJ2b4cxVpPb76TkwItuT8hy6GSEHVPZ5Y2NKMCKbRQFCrILGRoUXx
QJDFXzPJHnTmiZyofGUJJ3dwD+YXDDlYMqeszvEUF1yh1/uGXO8p8cmu8F6ndgHg
dQZ7y6vdcc0AWXclp0D1STR6rXOqjfdOQeyVVjtMfmGuLrxQPk2d8qm9GVmQNif6
/W8zFFELLaXZbZMb/y73QwQMiYwUmNne/q74JCxiSvWjzOjOrQIpiPseOcG7Plow
QpoveyaX25RGVc8rCvBhjJmJAniITCOh5HnepDgkH72iaeicEm2bVjIB4pRFBI1n
SizlGSHe7epNgtFDcRQLCE74m9TuR9vEwmy0o7XFiSZ3iKKleCYFfy3jQco6+jsT
03Z0oGHgJ5knyvVnKEDKp3HaDIum4ISc/rF5ubUD1m27ccBEYldJsTmMy15NsSCJ
QD/hVfZ3q/9vqkh6dIAT0zi3rquYAE0+spZdIN1NmwBd46paVucTQabRvZ6MH4y2
Es2RcZHaoPnlSrQaQ+vDSXTymrrHjv96BcnoYDXnpYHybSAVeoM6r9zEIZ5up4s9
tfEdPGnfihXlBGfT6iwrG0+bw+0KrTkNk/W2XwvbpGqZtAZiUNtKl481Ukck7f5B
rj5VLRNtkZJeyqwiM1iv1e6MHGkQIZ+PA8qAdFkT+MeTtJ4E9DfHXH0flvO325/k
8vmwEQlI7eN/3nSTbbnAJIs/Vc5z5JMMbKbZ8C7aKf3JMHE1SPEwZuXDvoAhAqUf
QRFyyw2Sl3VVSgf+1tqrR7OAs3mShIpx4DylmEc1XN/VPXrrD524L+U61ivyxNGj
wYO3hAxd24WLYlsPOwmUD/QM7ldhZSpbVlDIXz7ksM+MgCIzD2DYk3ebi5Pb541s
bxp3CxEFZOayROeyVyGD4jssOz4eWeE5nkfZW6ga/+GS4dIKPQVY+nH0lzyhP/u7
RzbbVccFAXSb+WCtuqLdyWrDM7GuPI1f9/8p5F5bX7jc5Ch6jys6VT+rc0miNSBi
e72eDC4dpKwB/St1+Hd3N9Dtv1nglzNIVKN8NDiVUNk/on8gYH7inYanXHe4rfaC
IlHrHdzn2GlOU08WJrZieUSqO0VAK0suqWtwRsgQrNxm/Fpv9RVTgUZrjvQdDTqo
qibtRUC4DMHOtI7av9+TlrqWG3d7u3fJ332Kt1CZCI3ovEvZNzEChK0y7I3QlEFP
GlLDpIIIGW+NJeyJoHriLDJGxQRaUx/OGrXAB3T4wEmw8Mc2UzANvr6zEUja1kbs
DrfW+xVgS8SqGGagI0SnkWAi5dZqDrprwM3dYrwmDSnCejV/sp53bR7K5GjGMu4n
ifCvI1J7RgBvbW1QVED+/mH3I6mG4gVgVBrGE0gpXOefGMwTdN6DzfSyKx7sxkCQ
GruajGTTZ/GcNlv4crQ86o014QK2K90N2llvFcBcXgc6DfQdn5sVUth4g5goFZYy
mJxbrMbKtXGddyzesotFPt4cqyrQoGdL+yPe02YCo8/tewGJ9p8bU9zYZgy3R5sg
WcKkJbLRXMtMUB9/zKHycePvUxpn/MDpfZ9ePqW/PeDlrgR+pPy5HkRdDp9oiug4
eUDk7xOBBW1FJqKWQ4jdJAiqJdeKYhgbPpyufbl7sLxY6b93UPxBaLKOVk2XZuJp
E6FIfuaey6CE/F6DLSMaVB+TKBUCytz166mJwzD2tbJLlKspWmVxkhH7Og4ss4Ol
D+zTdpySvSxjD+JDzmsA1UiEceInXN0zSHrI9xDEYGF9ReM9yI8E7/BwNnGUtxsE
2L6Dly1qsLX/Xth4sM5N8vwcRMu96eA1VZo8E2+YKZtjW2bdxi42hnK3F2HSVNLk
A5YDCX+H5k61m4dr5wzfofbaiSL2MobYxigP8m8fj+L10b3PEeJz1m93auN8gwnZ
VFcw5OirtW03n47DRmC7FVGlpuQl0w01bXAV6OQAGLifdU0EKwk2afCBe0VXncvb
eaUQ8IbEs07DlglN6DsZaXkT0dnCRr+rdS5KJMNm+vYUiCUrkuthvd0L9yovDGy0
4SaIEAtOChXUckjSqtjPl0q4exAMkIOZnwXGUlePjg0QC5Odi9iRcC9z76zhhLtx
P6EUIo5xDSBJWTHFNgGAc+De9AYcrVQpQD2cjd6QqD/1cp6D4r6rehIjOwBRjUwX
26bne0tzjPzpC2LT3cj99rz0/RtZVIyyKh9GRU6jzn3ooPPmhjOm5N8L21UUeJ34
cvfkC+yLDFA4m+2tgKJgd4+8aq8fl6UdwSFjdI1djDEmrut2fzl90twlSPPsHdlv
UJ9GNa8qdVM3Lgdz6Z+rdBpsPNS7twcrGtIHl0anJukVBGFaJiNnDaImEHm+MKXr
eO4JLoVfTXV1IjMn4l5rRwmNgxgPTig5ZFjFCjuq84fhkMB4pkqIo7H+b820lkxb
m/fByMQGoKz3nmZfcTt3eDTQ6NkFxRPmoN0uaEMuWzqCmvluznhIYveRA0ihM9k9
h0hYC92pcvK3B1a7p7E6y+EPGHOCdGZEIM3lDojJPmoW6RJDV/I4iKMN4hneDxHO
OH2a4SR4oog4b9dxt+CmtXIF8vb3Cx6WUz5zgUES5jtP92CmACzWDf4ealug5+FG
W/cQYcyCpA41hOu5HkvcZYpp+IYmr281VPWTLD/mZgH8d4ezPCPuh68+vhojPKsQ
wo1oNzW33CLBgig81yspqo+jlnV9vhp7SjMVxSBxDghCaU0WWMY0lc6L33sF5vAj
KRtR8KhxAgY21xPTV88TpCfmSBvWhZThI4bQ5cdvkGfJx+PgTzBZ515Utc1IBRxc
MtYGa4T5S3P+tj+M7ik6NuE5zH/eVfBiJ9GsPBhk4eXxfi3MWapMU8pqRM8q6d3d
HZPzSwZ3Qx0KNyAs3AdZPpW12CYNHO6GaPSVjSnXzNxVVvIMPyl3O1Y5pdUKWUiU
CMNZbxtoS+I5SzgDh4JBPuj6Km4St5MUz/AVdpKMLBlOPyr2uTiJy50fKvwWMjZc
XspF30bAGbJYU1aKLFzj10t/Rp7GMY8D6Qt7lB0gFhactYXNXDWq92M0DmKq5Vxm
fMubrmdaINmSRgdvAqcRNVEAEK0oxZazJmk2a7CvQBs4aDx0C2qUGK9mdjcXunBa
huOQx/hSLdf8l9sS90UkUjTPPxG7Hw3v3eWKPzRIqU2/E8SDYOFQqjzDQmqHzTwQ
78ja06cNCgJLCuIMb3G+R0dUrpYR6n9oqfxBBo1XnFGmk+ddBO4i0OxX6wQ9hSco
AMqMrhsTFgyJO5hWmqz0TfH0W2ziil3qT1z0NW7wV+wSgWeukt4TQbMgAusFHW3T
bGLlAEprFr8Mi1goliFBSj4m/0/aiVsWqA0Biho22MJ8tts7Uavb4kIZuLkbixDT
9p12CYSa9vlAnBiw3wplwe0isgWl8bLqV1W+0REC8OATnd1MRo+SqdH/5qVJ1AeO
VLen2ZHXgc9lTybbB95guaY68C8BqrAFgkKh7kCUjdCFMOsr+uYssQ4pzqfcl71o
oh59K/Zb0IlYx/J2drwcxGyucDoEuPU2RDInW4xJkuftD702HPLWwk63HCNA3Wu+
VkEoExvY6oE1kHl5fgkmMFj/H2sZDqrdXU0MZ7x+azJX1s51WoZBp1tCRRwU9kll
uUZLzhLKtcswKmcgT067lMCv74CPDm5qA2amkdmQKFm0yVZaNcCnd251QSvaWc7/
gjCQs95EaNr761oUiu3PEIDTAXrWygN+49SSF9nK5mNXjvc7/alDZVbrBplUHyYQ
HZHWnp89GphS612enu/TuAOHheL9JuULJGVILVgECRv+r+utlxDL62W+AnNuSRze
O4/baDg0R+OHLpvrwf2hw4ZRA6YUp6qPZTdGNnpXZBD/7gyoTmELUKUIgeb3q+Lr
5/rXqotyL0lnQwCQgLIrRowO0ZWF1Zc0DyDH6Dmdrjp0q+zll47xm42KnNRtzlg9
qEHo+zHa9g8wl4Wkm8wA6ytinn76FndxkrOXo/+xUPegHCg6zaEfNQMZNXWWMYvy
ykdtPCoxVtUeaG1qKRFvG1Tvl3F/F8/MGYzdxyNnilsnq+5Z0U/JAl3kWGlfKjn7
0HBfTO3b45PEPmOUF9qC5xopc3ki4Z98FnJmHM2KFsW7p5VRG+Apb+sNaL0lTHMW
SuyMMzSuY6zwn4UQwivtPcfXrjKa9MrWP71kMbONFqKig1YE9RobH2uIfXCHKtQy
VdSkHlZZccfEacTYGpwBq8e2KaKNdfNX4PvFbiZjH1TpxloIbm6dN8DkuFmnfR1G
r2ZB3zmHdUkU0e9aYyBBQXwYkcoWNaeUjuPZ3/sPltLhKvsQTNKhOvC5XN3acMZV
xGZ12ZEXKqc4HLuNu9UG7hrj7wukUi4NHKSuobC5qIWPXJNR6MRBVlRUgr326Ss3
46k8FvHfjESeLe4vDhtYoLkbZcoOV2qAv2BkL50qQ2MB6s95Je/vtT5Z+bSdQtpz
CmWjB8MOphm/537rvOeLKxsohbdnscnkwmiSOq+ODjabj6e4Vmupg5tlv2aKnqZX
awJEORp6XuvZ1BqSP0fy7h4MfsO3WOJ9kDS7Q/hEUUHVrrc1ZoCFPLhqGy9sK7M4
7byROBIKd6ENls6Pit2OBF9wP6muHuOC7A1Ht+q22KQRXhLBTaef/8j7hlAo4+Y1
VmwgUYb4SNxi30DH9Vf7ONf6bmYpAgAhB4FJSRI/9Z4I5Yuv/ok5j0snb6Kr8r4T
JpFAB+Eu8qoAedyz56y2YuL6X9mstjQMps3prw6W/tHBdkctgFWM/rHkzhuKrm9B
bI9gOIpARdqwjre8ueIusNB34WTdlFS4GD8QtmzKl9BvFtg+8sVwY96UaPo+vVTi
C6dmEY6w9jMkAP6bWin4UcgyODfUJEXZ7FMJabR/vMBPXJ6/gv6gjxv0huDYQJSg
zNLFFLSbyAkfpnW8KY0IdDqGXPy5PQ4f5E1hQ8+6Bmz9/MlbtvEpoA2MHxH3gadT
OgxxnC++t6xhk1NiwDYoOf7mxL7wS4tcBNd2w5ek3jc/R7vE7lj/K78NojiT8iV+
oOtArSXYhehufPeSgLnMsFMdJVz0hBnjg+oU8B+UUAAF1dzc5lj9oFke1zi7BPTQ
/yW0GRwPtyVGBuX9FxUIo5H+Ik7PY8u/t6P1+asTTCHo8x6iFaVT/uwtL8wEf22B
w0zsO0FTcMLzUfpnXThMm+Il2b75twCk/wf1p7UyG8h8Ilkl5sOBxQNviWipMWuc
8GrG3ovUF1ZWJ8Vpzd6hJ3zzzwT/7UTa07k0IOUvX/TvY9rlm4D9IyJFeUKdoF/y
ev8SRkyubsnnnWVou6l07fSAA5guaoWqQ0pe1EOze6F/1bhGw9De64YDvM5Vri+r
V18yv4I75bWPhDL2pRJ6NPpr8Umsqk7y7BFrGxy5PeIiX0YiWIXCVnMjfLGZxVxG
CeisPQuGxOCkGmZvgWrAsNG6l1qeKwRBzMtXRAiTlZHCh/qRMUTo9U92TM3Va0ZJ
SkyEV8z1LYWQvIcQ4zMUvlgWl/crhipY1+9iP7Sf/UXmsWicuDkPmYk4X0YS9/Uv
z5Us5OSPH04OK8wnPS4rC9akqb/lVeMWSCg4rsEhfefNYSyHOJqErxZPXFRKju1g
UrTlnoVoMwowYCEjKp4l1tVgGjFHR4u2F8dKNFpPj3UZr0InAsAM/gBYAN4mqycF
XeW+RVlC2NbBJfbRpiP4feFynYdpedoVu8c/DqccaXU9rIStP7/TQz6U2pmHyPPX
KvAjEeimCNt70WsgbiIwpo5KWKMQ7oNGjJx3D7rjVkNVs3LGxFcRyNNJm/RwF6fU
xVShOFcLpFq9oiIaWktC8M9Iav+Bu1BukqZzK+t5rp0pemRagPoW5oiR1o3/1ADT
MB9ui9TeHxYOVJWD84lxQz2jaiOK8Q8/dVFO6HweR7Fz43G1Ma0/sq4oJ6AvkSlh
w1L1x9znHM7kxkrOoPovvD997w70YFsAUTX7yNp/5pD7rooZq4WZUHGLdRMZ3ScK
rs/pktQfTo3oKFbbh9/CVrfpvVT9ScjCwskecBFBC0xIzw0vVdb/2tlNyiLLbaBm
IAPoqrBCiTMQOwpmP5VKnWPmc5wbLIMEdmGENT8xFFc/o8jjUOXPx+6QUr9OGa00
pExelnAd0Pz7MqlRqJeksdW8gs0DDjIkMo0lkHs/iKGaTWHa7z/G+VZ8TGoiNHSR
nVaw08SUYNeEb6CWOTGVctXDejWBpRUPOZnCjNhyTD1tb/h2wiEkCWMvnVJJaYle
dHiR1IOBpGHd+KX5hQatHTzfbSLHUmO9sv8tjnY+Ga+ZnbZegEQwze8z6PJyTWjd
ToOJX9j0Oqwl6CtjVcqBfk11NEs3LO8GY73AUK70N0qLwdCt1WQagkOEDlNcFOrq
c+4T/2tCWii4DF79lOQJddExvE4aNnuls8RXHpZepIpaJ4tC4rjojyJDHbWcQe4F
VFbzOLbXFagW5jK6s8zYLTSUeosqM1RUJQ9+M9vjUVXg8kcHk8mzIe74ZXxJr4Vt
HEiWpJO7FK9+0Tj6gfIS2IIGM6mdelMle/ZBsu5UMaX5cr4uqoPNkrkE0lh1dYW9
4Fuwe9yHDbd2UkzpfE0G4T4QmmeTa3D6MJrRNR3p8GZ06VoIABe0IXznUJQndgMh
oVn/ej+PawqOsBHfEYivU/EVP0fsYubvjzDsJeyPWIwbdAKB48jqSAQVONbkkN85
+DrBQke3rktHeSSx7+U9FfPqlLhvQCrnKjMe0o1y5/87eCGvJoq8mJ96X1rjrdcD
xLr/rXykaJtKBSVihRkYCGsmyeQ9dn/cFoRTNymjMwp/HJHYZN7WhBQxJE0J1dc5
4w77Rt7h+sGlBKR+VwTvXkO3Mi6VGkih3nhI9JvZdHlLav4P09F//gaNY4Z2KDDZ
0YjdEtJXY/O1emIBRiVRsCRHVyjkNF0Nv+dKqoHbgUIuwXtf5yZpnYT/+BS+HJ6I
D+i8r2ZKOhraVlhQCOcYpG0PO8wprQN1feXIBr0cfWjV8lAfdoPP0bIQzzIH9q7n
rA9Cfw4LUqA0dNSM2foKpJLcYjPIAxpc/spGSQT2iBFvN+fJNFuVNb862ESS6tCa
Wkp1AcwiJ/WJLyvafbboZ8rbXb5rBsWPcKbEUd61SEI6UXQ15HH0gCu7Okvst0Ci
xc1WugQjIZAEy2/vj+YJF8Y23lVunzwXTXubMSHpY0ELW1dcDAarfhNzdSTScVIh
t7CXuPNntdmzknNj10fOWT2wuS2xeT9jc7w/b2U84VY7UXqbp9IAHK4RHYdGgK3r
NN4STG6JG5kzyt6uzql63RE/2dIme2IBsCCMuaLNpcDAz+I3tqoSvaRZjzpiT939
PKoIUwaaLyPXLQz6o5USdrfLbpRjNrnT1mJWTOzzeT0qG84Ats+vEMVonqxokJkz
84LHjajcdv5GYBFhvMdQzqBHnvVmHtr+A7qtLQW7CNI2V0wDyQ8NPFtW/5Umlceo
HdbCgmt+9a889rqOXqgC4ky4UKw2uV4qpFsjfHLEEdv+uS6FedqMjTBlhjSIBIGk
tbSlPYLuBxtWw2kGWkSxjrr5SklpuTyVngOBYKsVFa+C3qeTer0nRso1DDjdh1jH
rE7sFiTFwaFWzsJ6LKcMtjgP39TyaiDyMhIKccNLwawj3e0RYx5XqWVpqJ/X/T6t
0sT1qi3O+UDT/r8wKqC+LY6epngouaAA4yuRFeZxeG2/Gc1IQoLe62/+w0e1JAPm
lTU5Rcl73NyE3wdoZon/Rbk9Wh26pE2zCBwbVoibckRMuziZCEsVX4voyxaQuSh9
FBT9cx8Bj6o9l8dnCX5WpTHb77g0Ze7xcldmPkwKzYFILhtUnwTV3Mg0U40G6zTX
o8NGJlUWeoLvrZ90dLeRByM92FqxLQufzdQ9oudmL8TI1Dalgwl6+614HBxCCCdl
70WOTlpfSJq4vDNwOyf6AM78J6fjPgprq2ehvTzCiqpreOzrNGLpzDNuoDv2KQB/
fVr22BvlNWd6ylm2l6mbWXo/51i3FoHG7oMDDB1X/pzU6P2qBXTsaEbY5FgQt94L
MffzimML61Y5fYt+zwInDvc5T3ckcUqhzIux3dXo5oyLY80D2NJpkV2JM2OgdV5q
FFIzYw6BVk9nEEBrXOBZCRtaQvBGU38YGexMbOupEYlblu8TRubre9aG2+aVDPWU
1pfBQ+/6d7PGi12FmVDe3s3lLkvklvev7AAZlWc13g5YEws5FjWbeuGuXlvQ4izf
iui216X6zQYWbJoKD8SEdhXiVNtqKC8vNpSkGB1t4I80W4+Kr4tHUEeSyUW68VXX
u/Fb6+8ZMxaoeMQ3NzuM/PGbT52NjqCuMuIJBLVeiBVnVEPxcuF9JeFo6Do6ff3g
LFqeYVQsyKIo4O8ulnEPWM0iBtYIWOznsHLukmTwzvYCErKltgnoQRZKx8/VONbm
tMU6oI2Ub3zKtlelE479fpYdRaPrtkxLHIkeXPk2TQGwrFvli93gxknmFQ1Egqb6
lQMv/xUch8cNhahhwp+ZmCHun0ARfNkfvKIJW6Lj7ge+2cOm7akNMvf4RLEtScI7
jY5JpBrn0d7rEREmp2War2+zSgzl8yGcHVrkyqyokm/Y68bnmS1PlEBEJr1uX5BY
yUIFfQN/iKCpeqRw/hYF+iMQyrHerC/oc790n8D+hreZDnMKozIDOuPXCjBGPTzI
/yd+oSL0KhGqm+jxfkcfuNkmaeKyP2Gn8JJpYzDkGc1s2OFN61+n81aR6hjhGNy8
rrx8j9zjx6uqiH6z3EKuyXr0ZgQREdTvcr/+yt1ZgeWlEOfN38b/ZIZzl3Ckb6J3
ZWG86JLUfeoyQLPqq7ZilkYS8hGGXVFeuiy3HPhRoROuYauUaAPKJRfQQl/YGB0k
yeo90EcrhGNfa53X/orH89qupG+EAcVxyjqk+jZuCmZRmMzeGxYzTszgbnTrzDnO
ekABPRoUUTlG/P+LwjqcQjmkj3BwTG/lxBHgnvV5RK4sHpcDeqyavlzMCUdVLO4c
pY1pD2YeGOzwC9XBKKMVg9WEwi4nA4u2+UgYV1ccqiHqt6V59kN7XQ9PST1s69d+
mD9VThsGriWdhRsio0WF5bKLRv+2B8wWSv+Kjn2d5bOxPIBMwugnxdBvuDaH3bgj
gmXcHkbkmcNdjdDQ0KoVHQ/Pnb8zhknZsJMRq7NCFP9Qhha9z59E6ZAogQIc9bYh
Xm2SgbUmho7Msps9FkyzSul1FqyZHmGCr+OqqYq5j0SuOJlSj6k7EwIWjMEzL9ky
yAPxUCvCSfcdAveZ+ZBh4jOMRyKIFHNel5p0izaabLKZEJmRx5ZgcZklO9JX6wLN
A/gcK5opMBIUfOfdTT4Swx0ILJWIvauDa4T8PDt7GgP+Q4esdGDHkv8jwQuhQnrU
wsZd5fIAEqIu3CvWIe6gket7ZTuCahHwybrVbwJOJ/2KpU+M9mCgzH5hTmD7bsrz
y71mctr5mi/IELHCL3rf3GFBAmPCd5hKbni2iAA7JOnpgn46af64GfrLmB92mWR8
m1uhQJX0PcQbor4Py0QJc3Dghm8HIs3rOJQOCf2oslM+NgbX0xrsjnEE01vCouFq
NCx7EcWv9hkD7iMyJw28pDfbLV8lIij0t6IFTCx4lXj4BKPnzPgeMHUwm09rVUdy
Rncwho4LgzY22cS2uzN171lbDX46cGZ0S9yEwa7q5klDxghGJ2g7ehy11b0ylDtQ
mpZWugGJEtBdkThSiRbshaEZhA+6nC29oS1DGqFQa6c7G4EEmDrT4VcbBcLL64/g
vJMrkiHrR5HQhInZ9lhhnOJf3tx1nZ+EfwwA4Je7bo/ysoC9GLvt7WjY9a8z5K1k
H3NqPsTRQran/XKq4WULX0eaxaSWg10f8QZTOBzvGFCwRi1uFANuvQ6ncg7emh7w
Nm7x7HjDUdKarx75+2ew6wCvPqPVn0j32z1eMdxr/10bDRuQ65PiHQpIG93E8Zg0
mz9no1fc3UJc8gtV0I+qXINVu9ecaArdUZbROqYyCx4cfB5FaH5wlbQzm0Rk+sit
LpPS3XcNU3Nv5OHau9fAzxeOkiP2VF8rl8GB6y2cfFdoviuPDEC0giWEEM8nzlY+
RtZ6tLnmLIhDmmP5mfu66TAEp5g2vcL9IPKOAQNSr50Sv5U5o2m3kcDhOxHoBZPP
g1x2eAG2bdwBmOW3aAAwprXo78QLyLt98Vi82zKp3xFWqGxuhfMlhf6P2x4jqcl9
oG3e3R3GQ/vp5wvMkN+HFVHma0ZYvW64U5lOPPDXbpYGDAV3dPCFADdQpA5Npx3m
TemRVWhhcPj3JZbvYEimYNgNS9h5gBOR60m8hJl1HvHyouzki7QVjXlejcbAlxL0
4QmoEy+d75I/j2e0HZh2oeKKtqbZVM6mpyaEFEJfLVBq/ONpR53dhjI4/4g9xGzC
9gTcnEWTpSgslZaRWvf819Akxov+mDYDa7I1D7u6XWCjsr9VS0QhKVLhSwL39W+S
hejRyvfBZUCgQ3iUEe9ElYN3XVOSNL/Nvkcb+yBZEHJhsEVpFp1QSkiZC6Jixc+L
18ZsxO+tqBQZInswHROW5HJCAvqY5nUSzfwhnfQKaKMc3Vt1EMY/EmYwMoQww2d6
zZjLMmOgrxW8yjNK99nI0xwjo24RhNnUlPFJxLWRqZLQgD/3/61m2bTfMhnJhgnw
gm2aBbYxBA/NsyI3dT3Uq/oppCnmaS1azybT0w4BSTsRxEPw5N9Tv8K9+8PEFvwp
8Nc4BI9JgYBXlRjWYQ63o5hDX5ZngWqnBUrkyBTvIxhxTKfwgRxia//clIKHvfZ8
tMUAFuoE7qtGyInzOLPRh/Xc15NuCbSewTN0nx0tlke7CnXtFSdPJpv4/Hhd+k5k
aBH0FMc4KtsaLuMwXh73weWqR3Gl9kvsTXtGC29cAxrdbuGzBBs7F7f3f0KWJl0A
h3wXbU1EPXQDkrwt+C2gZzhi1Ec8MXmeCtisv8XtQOzDkh5K2GcnU1z1rpqMvdxh
yRyFj7IaoLFZYJ3Hr7cKQQifoQ1cDuyNk+hLu7708E4bbQ4MTP/pUeNNeKHN6uui
i+IsM53U26jbVeu3svimEWDup2VwwJwlvhazE8v/IC0g0TN4tT9H3GaAjZac8kxn
10dTDXvmEzYIuu66ttGMnBZYL1JvE/54snszma936VPC9aDCp/IpqW4daFCK8CCM
TRswZp3PmHYV72Y6m3ssY/4fgS8/ObLfQf4fm2ZulDWyPPQOwOEUFgnI5S7SO7vM
3w/gqup+aNZ07HUmIkgrR4upGgL/tUkW/kYjw1EAPqdqEXroXzE8Jadg89l1q/Ol
UDXtCxGavvWUuWsI+h2KUwmDQhT5X0fiUDGpg7iizztEwOdiuJs0TtYM4FBgVtZD
Aj/rM1yrq5Yo/9VZiUiHBQrToY9SlW4BY5D1XcHwJn+m1adDhvItU6baPCZfylb/
ek/VNGP+l0OMx9Jzta23gBIwIZyNLapev3GoJ2EK3pZU/x1rfQo8+cUJlHsy0DKF
/EMTszEw9uZYXWROYD3xXwvJsRabioC5W+tqXm/Sp+toot4YwlBW1noVt5ipR/+j
2VtVD8a2uu2macVHWY7kSB3/I6hB9gzDt6t4JgFOKGvCnKpCdXUx8/LyBcSA9pgQ
FLAc3w2Do0+0P4HwQ+nJ9S9thOJBjniqgFmG99KIoL9to8OV/EWIFs61pev+bsR4
/1y4DSuVcEPM5cXruv9rUJk13rL2IKgQGSQEikHoLZ/s0CEOJjBfaB9FYPCMspNT
1bbVfAy7csVOuN/5RL5Nvo7ygwqqy3ckBOeOxYKeQDJwtxknK8ajkiN0KI9Rr6ai
9Ui+cvKOceFKjMLvC7oTcGrt0QAAaQ8liQ9N0eqj/72SVioFuxOtfnWgtLbmWvzo
ft8gsVqz4dN9zK7FC6O4nmkgVeKH5sJeQ/cAMq/Om0V0e90Jx4KaoS9DnPy2sxuG
BjffqBlmO+wRpFU0VMy9J7zKK95V//XkafNWUcrtgx+77j00i3/4JXMEwQOyECkD
xwXclPTnfLOW7xZGhXBckWS00d3vM6ZHbw09qxATNCbXU64WN4KNTaGEUUoPLmQn
IMf5MIsy1Y554jTSxO9Cc1v57HEXsJcY/ej07WBNqD5MzUJ0/fmIuBG9RMmsghAS
YTcOTo+iOcSfvp0icqdcY48jWGERZUuaRN5MIKmkgnn0suQwgVLFTxmsH2swm3hs
a+0wErtMTX1AbeCxbuCKb63KmlhSMVWEd00tXKwxJzsVJvjE2m/OYOGhl24t/hlE
UvHTsFIdOXS++UqtEfi6kJmQwn6kjqbX14E9ONuKJ1a97XK43f8nr2t24zD5zHVc
jbisWrvkLV1/h56DhGboQldfF0HxhdR10WodT72fq2KX/TtzfzdPLS0AtjQ23OdY
8/6NGL0OuJKwLI1X/+b96IZZS+hNFtgAojwY5LmdZlKiDbJitwZ85E0oupOjv2XU
nZEK94lwVghmUKgMeUihflK2LupdYnprveEdgz80GY+NsXYNshUh8VPpvoTuEfOw
D8+LMHb963yBgU2fdYSv9aRuWh5Z0xMYiJnXZa6/702tBspc+wuK/E+3CpLVeM0L
eLscJCwCK/TZ4f4pA/QZyymO7fSFX479SGyXFYHrB9mtxNhXkncvo0bg2VfAIp0+
fttH/iiL1bVGB/fTUQWmAC2RkgWN8h4b5yt85819Oc6YvAU+HtC/ohyspyWYUwZK
M/xPpjbQfRDOl/LLgUO+bDp+7UkRN/6JF+Hge7yzrUmdcVCAYspgdm4t8OI/j54T
ucjKcdWrzwsXXurVjKFNW3ECmUA//eYExjqjCihBq4gmSKKRD2jtOiHydU7a3WHT
tChahTE1eT0FTHylZqs+61m51+rMGDK+JtJItoMuZM48lj6OuzTZmjKHpZyOfOX7
vRzrDoch+C9vJmPV7nTRBF6vAKBp5jjMc8/Ub1/ArCyDLjV38zLFNhSBT2cnzLYe
bjnRyHlYCNNGmRkoJiT9Vb2fhMedPYBU+SysFa0kG2L+LY72JG74vJhWkuCdJWMA
i16FKfGUAYBDk1mdJI0L+gey+EmgPRLErmmjadL8U7uCIrw9TqF6Y8d75DhHX+vc
b+JKiFJji8fc1Is8O+1I2iYYfKo/ql8bK5MTnvLKnr7ZuTBnzlhhx9eARjFg/oVV
m79VjYjHxjn7kzwfCiTDNj9akY+dLUkTLDUb6d9xaqigLoQy3N+ti7tNzWindjGR
9qQNGbiN5khiXrzbuJAMDfXul00UqpQEP8hHc2N7eIitD31Hj18xtazK7XY0msJy
jSbYQuuFTbz9cYy3iKok4QLzEBGz10usKpbAvOajpwNwkdo33da9j1BysACNvcPh
hdVhQXmsdu/yPcP6dGpMzEPuKSZ6SaoxW0aN6w3VYXvGtzKYGq80wbnYWV8txNLl
AKBcwuEMXZ2KJ+3JJ6APe6J32dTQYAfBU7P5OHk8l+w4ck9xY7JWCKQOo5H281DG
WIXscBj/CtD4v+17qTUh1rWoCEJkm+xRpD2bgCmdg2Rw3s+LCD050e7H2i/jyXga
te6bR27PRgafvLULvgX4sssJV28wtQ117G3pjdAeDrEi0IligJAkK+e1BT5A/fQM
/0WfkVYGVAgai+dnZKVm8iB9OptIF1SwF7KTzECVITbMxHKdxNKbLxvbW3XHfwtY
BSNhPdtEEZhzOqnfppAql+ujSStOQdbFsZNUuN+p6NhNMeVA7tx8YFajReZc2+bv
6K45phe+1RJNEBNTMpVjMA+QMWsZ4GyVv9hYvjS9dR6rBe5SYVnP2dUBfDI5IrGw
DyNL5oFT+mi8xXqWcfQ1OYvV3likYsDTH2YlSdOwrugnEyEOXZYKMsRjWUydxSj/
MTP5ZAWD+qvBMgXPA3+czpytxQsrcs08jBq4Q2avko3yadG8FuhA/rL4bolU7Ejn
iu8bExbLPcmwSfOIne75SLd9dkBRuMN8pX46AXcVzolSrvGNx9SLm4HoG6YaYHx0
fz8CncQuFs1hcZs1ADgCEXTNSn9SIjRBNnB+OEgKE6YDe6Vn0Q3VTLQ0UKWkdG/B
eiS7NHRk7nD/VGN/R3bfuxeWAck4CKqtwS27u0L66KYe3rqSHG0GwVpdX9Uvqn4Y
+pDS6GSKmSzBl35IxB3VJWeBaWFalSUEm1q/ps5AifB4z0nMzmP7ZaR4L8B4Q6uM
AVIyMy38WJHuFALiYLa5lpZm9NUhohbG5rCuGgAuHvR6YTM3dgc0owLrj+oavAS7
HOCUvYl99wx+dwm3TiYurkVboXVhKYONWOMjdHjYUWptRDvVtuDIGvMDwagBa5AO
qbzitXSFuTma0NEBh6HwFuDGqtyQjrkhcbHKpip/xkhC4SwlgG3FK8vF1xVaJACE
eGGM9Ux+C1iHAowb4riy13OlO5VymY6P/dPqM2vJruJGxea0864+pRQjKWTxcVOd
xXqrVedudUKS4waTic8Z9Bozcqp/pqnw0Jdz7hAeIwDmNPsfoNOJogwTFliWno+3
RUE/6kFCZ9S/YUM5ium/ifvImnfrjsvMkg4xU4CINiLCRHbqDLcnsZOxXvv58sAN
8hZDNpnY9d8YXFwD0+r4XHbZK5h988U1nmwFod1tMGCRrolz9o/Rg9hqGwFhlIKt
LsEmoIMCxoqH0lpRvhf/Jh7h3TUnq0J5CdBrd8+0g16fgp2p0lcY5LnQGcs+nvLY
Y+cA6MRMFz4e2aYjqcUz3Tjh1Icl/glVODCgsiiZdWhBiVVBDluYDn6OP4j3tqoW
qbba0JaSWAMkzDkTRJR98X74PuMlExA2HsKSWmyDCofIQL7ou9kRoc9aTdKxBwCm
pCBtIh6zuNVQXGenq7DvVGr13czi36brrrnAxwkmmKZXVN2vtiMXrgwBKDKNGNvL
5Wu8wzEUwRe++CqHFmPs7HNzDJD0LjgDaTwUjNyzuo5fDmKAP5hUQzxmSXzpon27
7zwhgjgx+wtq+rAsyTJg/JjMh2ovFdZN3m9ZIumYwpspx3VkoZ10wvNqrry0Icb+
kdvY9gpVLW5SvmYVLtzcLxDR++E/PiXh8CeycF0eiUHe1VnE/fO7FZwDDMgQUuIC
RA5GKF4wPzQHi+qRv25TNDmRihb+H/9rAPBV5gObmIOQ4TmX+dUG4qaEIBAtWXwz
Ad11xOAqibLQ2DoQbIhk+l2fv47fhqp3krKTRxEFerqMfH9Lxcjv5dee/WUfl5rv
Gnex9r7nQ1jejSpYCWu6lZmn1c90KumKwxZZqO1oqqB3VqjFHSs+5rpnB2j+g7fb
qcY/Lro05lyM4r5ofqJa2gApUHjvT/1lE8FHIGELwvcHXcn9vgAeTRc/iMONy/og
/CQS73K7Y/NKV3R4hNhiI6cwWfgrsV0BAe6P1UyiC4a3zvMnmXoGl6q4dalyse3W
InDXM1/X5grOO13gO3ZQhnSXeudoDu5J44riUT+PwYK4Uh0eizPh8LyLmiiW0nGa
8mPwTYJAiRSrZ3n2TeVTlIpyhtKfMrcHYC5YncR8rGNHndR4pLcQmIB9mLxj1n+h
91EOJuJIQPUPxady8kbXE4rQaWFfAiMpf7cZiRyYNrlc51BUuD/t074RiqDsyWwe
oqjt602xZJpeCLWOpRQIslvrk2/rhAgGHGGERnoSpknuqSqsASpQ85G0jQ9ddViG
TgO7qPL2F3i7o6n7Zu4Jqz6ZGm8GS3hBJNUUqk1oOuEc05qnbCxq+s+Me7TcfigF
04FkFE3ww4FblAAVZY2y+WhSBoPKVfGmciUHn7Vj1blJp/I1jyiNoKVb+lUBLJfJ
PGZa4y+dgwxq2T8iAlS/uhUN3jBS/Ffb9OBBe1R4+AoFCT+VOnmN16CRWMu0fz/E
1D/Ytu5+zngiuY7KHfOvdj0oTPOqNs7gnpR1lGeH97gJriz+fYAZGtGA7za9/Jx9
/LX1nKaSdznnrJGhLvnpIT2DtlO6eDh9Xr+fcPVRhArEvncCaip19KB+XVbnTfSK
5Q60UEPKO79uiIwFHCzNiT0+TszIrfZWt8hzfx69FchOqOYr6Nl/E9PPuR70EyMW
yUX9m83ysO3qAybKjSpIcn+AeJnYQcPMwz9CQldHRtEN35OCIWxXYtRAyX83TzaI
hU0y3EDbQODJo2w1F7EJjOUg9WOrR9zPn/Y6maAzWff94opH0SctN+Gmme/mcACo
biscB9KqU0jnIPtu0dsgMBZ6KRhY3UkCzVPG53OdtiP8wVL5RrVvGOLAEi6S3E75
dm/6kQ5Cgd51AWCeGefWiGqi8/1tEjd5Su0I96zYzrWaCigPqFY82NnReDsnAy8d
sIpIXlVl/qohHdeujThqEyEIbgCT736ZLLJycu+DvN8//PIBUq/43mLWkHx3bbB3
0i0o60z07s++/GiMFd7pYNNch/gctjO5Sc1miJLE9OH4lGk8k2jtZQ16H9NWOGMa
ewUxwHPlVsiRnL3gdy4TluhQepnlr88i1Oftt+4zEq+9nnEkrh65J7NrtwMpZjHq
5HVSl7HB9LkqGHbcIGLoCVYuiEzJUhmI9wFHDn11ECIGWR9rTyeHchDn2KIfcit9
8Nvye7RZpHS5chTHrRXyH3yTH5wstpGkuLQtluN6cnycZ2A/8M5sVPGR6k8Cs+95
6HDZF4qeSjFQqM5ZSB6sJAm1JH2LT5ES3dsTboGrCkqFtrSm4aTCoYM/1sFA2R4L
UR5rLkYPd5HCHwl9XXnIQ72+VMthRoATjO2aVVsMYtJWPSm0+eTkQ6geViIVVYEz
C9hP6z7oYP4P4XnNmwFrRUv7IRq1yFXBY3FGnYKwAxL9gKwCdiTM/Kdk/bevQND8
snSVEnolmdeEef8Huzh4N7CpP3njYCJWYtEPEDbB6ATdRFyOv/ANKKt875n/cCTs
RnM8ov1ZT/oxK3eFZNz19ZLFrEeYszZ1JA+aFoAGSn2w5nF7BYip+VxORbkEmWKE
uEjVXA5Tc0Clphyh6/v4QFsPNs8KfZ9zi3eSdMzFS+w0A168wx9EXmAmjCYV/GIA
IVFDbnSLohButK9ZxGc52GT/he0gcQBWc94lixR26tOOO7g+fxibKpnKYGMu9bcR
H3doUfYtNFT6Y1fMMQ6bOUwJuqy9+nmM4aPxb7MjhuO16Bab7y6HMVXiubbIlCWS
EhlSv091ISW8K2X1w7N5VdPIf+7NyedJY50LuGvcutxwRW4kx6V0KkK3H0y77KrP
nYh9J+DUIULGvEKDGuCGkk38WRNrtPJ2W6PPQifvv6nEGHBYkXlbfz6Ngj5eFUdi
vc1myPVyO6f03d0YC2KyY/So/bq9Tg613RK816peq/cCnaICD4XcL2TsPEi8zwEo
3iud5eeUU8gj2DvavhgA+sbabdkEejkPVir7kNIueEX6VaPC+8zaMkp1fQNNjkH7
46f/LqfA/gJge7DQ0b0YaLpSJ2dHyStQMWCnNMnFlIvrc6C9Mt36a2+GFqYadnOF
iMh+oa9Nab7DIPMgAM39LG/b7LEPETGA+hN0z18ahiLjq68kxB2pZqJRNT88CFjz
bJmuyCku0FZbZutHcfqIAJeirUDs4TBSsOeAFq+160pJ3zEqEiq2ag6WCP3ar7s4
efiyXaeflAvRvexsyfN5RYSNU6Ej+gycznfAJPSXW0URPTVGg/xq6asUxgoYifwE
c6CcARz1jVLo07KDhOdo5cG/FurnVRmSZhnFXPc8xX8uMINWJWeYuVIbnn1zpLVZ
SYmyMK7KGrbmJ+hy+aNJIfYqlxbpY04FFcrFgEepdcitktbnVhuLNTvCfHy+4VzK
mVScIFbiWLgRuA8wG42/eqM5vrWJteKLZDOrJyDLEgabFUL1FaBwLrStc4gmIYSm
WBR2RjQJHG/2Zc1YJ9iOV6UxyUkW7FLP1QKannkwg6iBmma6g5YfWV7fG46LIym3
1PwnUWHbYkkSpO43p1qPBzzpKqCbOb0GjILfqlnQupmUJw0iWSzxVR4UPASJ2KPQ
TkvP5Y5zPxUyJHYrIVCMkFQ29fMyuSA/1ynUowYp6Hj9vUh60C+tyk1Sh4k9GKay
2gtXyLV6Zh6s9+eMMndnxbZZv44jpwU3HSbFkn60VoWTeevbb7HGHnlycbFiyQFI
VokNQFR6EBA6eETWkQ85QJZW2ZUrkErdKmV+vLxdww3iuyGSfgYwgwKsHSeZiJw4
FyYLAljqkHp30dp3b0Z7MNLKysoUwv6Fu6pWL1bJiE08P+PnYryJE75U5hAkPRdr
iZsMRL8nl+ywLuL4L3JZm95Y0o5eyWhzxX7rLlEwu9sw3PoK9fOL8j7I8hDodbFK
Esq5K0xxBxNGTwlaOK85Yigd6jUdBHUK5cQJJPJ5fw/qQoyP6fRkRJwkyqH69xoT
ImAXP5Ax9Jw8MIAzZUYQtCcNqyJCWkyy1DBs/ZiWwDdRlArpCc2hT7fhZxpHNcD8
Ier7X1Bh1KPiHs8GISejYa4hkW4+sezcnh3HD4kG4GM6By3HDMxjMg45EKRJgz7V
XCYF9PIq5wH8z/J6N2YhpbW1IrTqs5enOghpCJ7LUpsT/xkhPC9mFR8ZKdHZulbK
TRR1VI1dQ/PREYIcqFDgeNFd5d0IYlvywHy2PRa6hjg6MRL3xM73+ik3fxU9xuBm
gaMFMjjj8Od8N5Bo9sv6zoG8ccJNtGXVCi6S29sZq62Ztil6OFJVh0TlUXGQzTYe
QWnSCx0TROPWv7v/+iso/Orexn8TZfru+00Mlbw/9+zbEtj0Wf+VlCBR7Q8pdW1Y
eAjAyKj1HcfFEL4v4d86QdNIErzUYjbUag9GDPofWzQdmh1SB9d+FMqcPe1zTDHp
P4hz1o4IZGgDKeNaIdnrsnBIB8PoymmoSlVTCXD0523Zfi56OyqEbZQ/HGbY9TWO
O1nkz2Dn8PlyFqTbX2Z90iZf7ivlpXr/Jx2LNpqC6cCvfKG8PL36ZFrLizn34X9p
7I2mnVCS8g04GfBCz7hVVEMINd+YR4+IsknU2pcceKHJrYfDcbeIjrQk5sD3ZKj4
GJU7glySZ6Xp6zzrZViz8uBX5vpRgFbxeaUoyObvOvdy4Aw9037w4MEmL5hicOTN
J/IAJL4PmjIEeXtuuSkIRlRGZ8rTlJdA0+jHs16aInK20NPPTMXkHJInV20TaRrh
Pwdn8SwQHs+p2myVrnrEteLy+gndXxVr2i6yWILfts4EkEZM6uZaG7FiZ6dHe9go
PQKER7rvUGViLbsVAn9NFuRri+Ixquj/qswzfNS/dTbNNOcZCQjfsN/7mBrt81Cf
JMzqWkDmLkoR/dDOND0SStrZMxzc71JEuK2f3oy+oppSi8y+OQz700fbuuQBStzD
lGUh2jNWrISqTrkxdL3+tJ+l6kex15jWEkiSFrcUv+C0z7q7JLUF3q23XRDjBqMb
qpm1Lku+l4sYdAH73rNGKs1s1al7XHz/5C5Cpzu+BxycMZBt+kH/fNSGCdNHiagO
mU8kNzI8cHKp9w077CczpfBrSwdxB9D+GwHR1eq4mQlqTrMpOOAZ2IVCI5FaPlG8
6bMOZYvEwcxeNduqHU0l8rzF9AIci/gM41aZ0aNJEoEVhi4KyYEZe6oUQfWEPcLx
iI4pHdI21YWgtXrAQ42TPFa/ryW+1bhX/wp4R9NYfK8Gn0v7XZPb1xiZURPbfLIF
SjtxvzrqsnyydTYqWkIPgrz2TDO00MkpsajaGzXyeErg0DJo58iTh+pwtGE7gvS2
xM13jgF7NEa6Srzw0eqDpDmXkG9BlmJb/QS4QJWSUE27uf0fq6vyxLzW8akXaaF/
x3sluXLiV0su0t/syGNb5ifTip2URSPo+NiS3kMIKVHmhvgI14VQJ1aB8Sxsm/L1
OeX+z0WiAeN9sa2eI8HU4DZs83F39MlcfDL+qNx+fmc7NvaYNCIIoADDHmZDRNWs
c7b8iPU57wmJ/ogeADcptjQaKqmh2edXQz88Jgdme4uCwUyI0F562gnwXB5bE5pJ
226RGXwLMZmilAE4FmHcbTnFiyJloCmlCWQs2Fk7W9C5eDOta4Bd4uwFlaVDtay4
VELEgpNlxGL7hXxvmblbK0nS8865kMYlZ2tsnwJW3Z4GodU2Irc8evL73eB5Dczl
BnKfWd7j4SfcHHIf7AZ3Ln/jGP+EKMFrXsGIY7W7/W1x8nBv+ynmgq2fdjfIMgps
Q07SsIjKe9bUtK5e2rCIT8HaUOw6womxzH8J6MY3K74vRCi8E9wNVVI157br/I44
rXno9/EryEU32/QBZoVw6H+VjR/cWn6qAsUW2SeF/On1ic+efqKCoNwIIRx01qCy
cFYZ9QwVeYQX6bqy7MlgA4yPRxnhmkCDGJaHtgzFxCKnFfdGatuBXmp4csU91VJ4
eNG7xZwI+v9XMTNh5wd4vx9grysN1XXPUMZ7iYXEhuFsMoVhqvAdB0ivw8AG52NF
LaBoY4hUaCzj8/AjGDqzBZ1Kif7QKgaAZzTKAm/IZA6NFFEu7UfYWZCLuCCcGEu2
DPS5UgOnuyMBBfNi1+LgS7IS8fqaCufnkbO4p9CEULQg1uEJQml7oHyzujombyPN
EhdrOzvWN8S1IJ28roGmoqFQCy3/5ZsgK+R2KDHDRazYG16rKHcdZcM+WJiN4FFF
Ex6VXplPnRrGCRNH8JiJe1+U+hRFAcfctY7Kdl/3dFVHJ/YUBkl0Ftjc67oWDDtU
DraKe9r3X82Ba4V1ujgtFt2B675uPamBZgK2BIcUFy2MR/Oa8qKt3r8zmoyovvYr
89rvywDZMJTmPVpWeCFBOjGUG2DBLyErRnvROH9IReSyGE97Cezknw3sI4l1dDJd
V8C0p6GCkz6TZ4Yjn9gNAeg4yWzICreluOX58T3C06qkYSEjo8BkDhkf/zZJ69FN
QCWRnRqJzTUIVvb60iLLCLdMOYU80oj0ri9BwUe/l46H2KCClsh0T7a+KzSqa7vo
veVPfkIV1z3sKnYDr8WLHZKbpvZ7gDL9oK+oKXLgGpSsiZzqY1S8g5pQc+5+QSyw
CTNesVJm9HbPtKL0ZarfCsvD83uw7VFvmYVCMvBAuNkHZ2DyfEMZHZfIwpMKLqgJ
/Aj3SucCz1ELo558CzVORKlTHlvGaP49OgNV0366vNK7Ih2UKBj8gLLt3dzlf1AP
lZ3wDBoeMKaWL/xiHd8p9ChkuUMYuG3fVz5PBNn/wACNlw5d2YOkjh3DOjSIqqxf
EXRZSFh1w8FEt7IAeBDdr0xRVKNUy6fSoh1/5MGeV/EQeHvpYRqWSrhoJdIJRRA3
VM7IxGyT2PBUH+iTvogpxe2kitlI2c3KlDqPmcv8ENHTsFChtblLKy3aUpBX7/va
WE844uIJpmf1Zm2pqO7fqs+oAE9M0/VNI+86HGDqdLzUIUCAi1Pt8LwLNIpAxzlc
XqYa2j1KGP2OZ6AsQ8iUaiY/ImPElZGz1yryJOZAUioweoValhmvFzxvO3sBpbtD
EUe5p60qs1ISsHN0+2qaxzYSd8Zs8Xwvkith+BYquXgm5VjyT8iPgwfy9SO+Lggs
U6TAG/Bym6IQzNUQDfsyGOg3pEmCd9sq+Hhw9MFAmHTADeoL//i19/S+J2cPafMu
0qpl2S9njzWQVLTfV2m2maXGN4QyHc3560tRJv5UoWu+6oUQwgkL/2ZOYvgDsWzb
k/MWcrm9WMXeuS867bIegJEfLt/mYrgiBlLNEwy8Ldhxcw4w2VwA6ZnM81kVHaG9
Em80r1cjYqJje6Q9Jh6DW6xoA3GVwmuP/EAJq9oX4Rdc70PhaQJUmn/sP//QkTIu
EfteUbJHP2sKF5VrcoHQgmXViK9f+cBY89qNJP4u88hVWcsE9dW0jmJ2dKgX0Qc7
9rzM1t+S80Cw9JOEqO/VEm6B+Ykc92sIMe02qzZ7o7EIw4UlxxSeisQ4PthBrBI5
cxcjw3LrnwJ1LwBDnVBHf7PaP0gqHrVm5JoPb2x4jUppIMlTJRE75e3WOH70ERQh
n3jjyZH1IX6nh3dtQ5Wyq8fdLu/ckOxOChJEIyIIUceV7fTX/z9GbSx2QeXRdyf4
eUv1zpEGfCIpNPNrUsERT5bWF5JFzkRpsML4kjbXLXw9USkhLRgb4CA2oSlit7m5
BdtxkVhqrjbm+gGkoT10b0ists6242aSi+4tJu0iZAPR2fd27ObrdcAHshhTklMM
8kCJmZnkvNV5smwBJlQMsCgYe/8rjHY39TjPdkchZh16CI3JLq6GM/DtHjrjjiwW
bjARtRIEaDdxK34AHbKmyb5RL1D9si5G1VocGYZj090Jn8kkYS0hzd12GXCZha8I
tQINGk4HeW0ZJOSEbmPg+K8v+ByDAvhZpS+KQiASOzTGMA5x01fiPLbGZO63VIpc
yj4t9QQeX0MvgaV6ye1Mv4zqiHALAPwsteF11/Ftq4sKF7FwWTfcX3gmDgeAfeYX
tyKOq4C212RJ+0yyWPuExOjrkcE7ql8F/xW/zzFLG32wdJ58pUpwlPuRWN/7r7aQ
cNVvsPhiTn1e7iDrRBO29PykG43erCu00clC2tmdbbqebHZJPzgqfuT0L9Onah5L
09czeOQyZrfjJ3JVnYa6RJwgOzCI9ZEMfKXowLPyBWcx4LkwLWph/vc7vsQ/B7OW
xTpnqk7qVQanspU3zzu+COr97CUEE/r0gIl3ZmSg51q8mM8fV1KQCUM6wZfFD7z7
050FMWpYhVTWotNQMpNuqbYpB/3Jo42268/IoZLGd+4mkdd7N0nAp8Shb64fmHwq
9M7q/u0bqA0Xt57aOMd74muqbXJ0YfyXO0pa6IwPm4k3R9c71j84PX39X7NHsUCM
0ua/b/DzGNXaNs7rxfsHFt1NkEFRgHTQWlOD/a9zyGmFBI6R2WmaTvJbTJ5BB7Ty
H/qF+dibV088Mmrh4yjQvq9/GDT53UAmcZfbGiyU53xMy7WXqVZjQOs4qxKB6eNV
dWq2t82mzFFext39LikxGAWx1EyzDmLNVQhZ6HyFYsJAkZ+0MUXNfl2JThKsGQLl
MDR4SL2tUedd96Hm9MNFjFud0hWrUoeDkvRTA5EK1iNmIxZ1XgVBxBdDfQscJ/hp
AXJ08gJ+n5DR/Pbyvb/mD4Z4waG8q7fygB9vRx3CoHrsDHgNMXfO05QZM0b4TQcL
I8E7HpRgscJF+eLK1bx+Npwe4jvblfxWQGxE0PoTpuOFzBkNUS3zWeKyTfgQVhkq
vI7pmFKQxBfvqDVwlu8gi6e6rqdG0Rnv2yVjMplyRkVidx+UfQsqxeLmgOXmeLh4
qU9BZNDR0oHpw3at+Onfo5qJo9t4zFN7GvW+BX6XcJQPIr8juHZ8nAF7Sv7MGyJF
r8EOjAwtq+veAAWUylJkUSi045gAxRcKIg8xHp188l7AOVWehzqBtbgQo5zls7YJ
sJK4BvGv6ey0+14w0rrCIZYNtJzkqKm5idtpQqA71Kxnjqmgz3fJ3VJLV1zvtA4L
kUDkHvplSVI+75KU6bhiCp/zcl82q13KMvk43zy6HPpw7LLxkfdhmeoc2ohVt5q2
uS8hbTuU0Q/5BihE1IPgZN7+inwvOs2f6gwmEEqwfZfHiDn6u+VgIi8kKmJwVtG6
V74PHRJi+s2vCCRPCDFVvYBPlYhDh3XXEaqUdkT7K2HKXOG7a46yGNfeXurDIeWp
9SBTZYxeohrI1QRqWaJoKRZKug9wZSKCMpM4/7qF6NRcXaWFCONmxHSwMvdE1ncw
Q3Iq1QbjXiouaVDZX5L3X1ZOkVZMcf5//SkzldicIA09/SdIwJEV1/3/hxnnrDmi
R8MREA/ZbpJqYjGof1O2+Dh/jCutrP84yshHIEftFuOCa/CggymRQT8uaMU+SyWc
X4qjMJoVcCH9Fduy+lka/wmr21bIiwho1sMKivrb/Z8UoXsjFQuLpQMMkho7fjNk
/2eEiWmQIPxkKRpTC1hYMs63k2czwWs1jCq7/S7ZooQGu0/vGJu82aagOXPnJ9E2
UDVnFG8b7M2D761rxkhTl03e0hXVbsVXMEUQxcvQFQzDrvUpzPp88Q3iuYXTTy/U
5tLozujMvTYxqTncRfKQx3Xnr5jOtOyztJyDz389Z68zJkETIBTVgyDu398nhMQX
Z6h18IzuxBnFat6t9wbpD799WJxzoFwOs0gnUy9tRGnqAANiNLXe2ZkwKucQAyC9
03WM4SqAivmW1f8IZZpu4kzVAafi/vYEO6UkPvzlmmnswHW0QZbFK/djq7IpDJM3
TzOwHgLWfytOVheSZHt7cvKbUU1MoDbWgdBhSUGTpqmgJyW/1HGcHwZ6EXcqdJKZ
lkO9sU/q/FVog6S2Dh6nYIzJYHdvsuou6uvCL7nkjHt7nDXvinBFV7gACplqwmn7
LcRhedN0Wfo+JnhtxpLZg4Uy9iDbBMS5NF7YFFJflWaxVmjkpm1Il4TOdgDvJlcf
lylCYCjca8/yXqHM6eYdeuVu5qZ0BRhZWvO3wSk2GygSsCTpgzx/ph9EIiLSrRnO
KFWlRmuCrxybR3v4q85zh2QxUhMBW0Ov0yoeosGlBV+aIQMk/Vn43qu0AeLUW/hG
f4wPSY6i6rhbn0w4LNZ0YbKJpUf46Jq/vEe/v6jHOuhoxLacgbmtAP9qmvAq2QJ7
6tMF9y80+T+2S6PQhDsrSSL6ApIzH/1GbHSi1w1Dk5jebgacJodnhwnwMqNmQYVS
4195ysaFPuhtWEXVvZML7c55QmuYrOZRrq/advqDemQSm1kQFNk3GnCrXdXrRx4X
/2FyBQCm5z7cl3KYug8SbjTNQkyblSUGmPmLUGnx0rVUV5630UREHA6Fg0Hcpe8u
DKHBpv5G9k52rmfHdFoulamtN4Pa15tSOHbquSpvfI95SigXo080tmZwSwgCqdC+
VAsQEp6KZedC11gkFBCRK83QTSudIw/S31ZTubUI2aaGL08eHxcqr8UrtZu35gEP
MpdyleMW2EvELLme3fJaY6syh5hCipj64oL+BmnonwaYjubbXhFj5LkBzSqAhK3K
p022Nu47HQbvc97tRTwUWQDjHreHK7+sE9i/FWz9zRPXDDT9yznoYUN2PXCFzK1h
6V+E3NTcGfoWkvUZSdAYrI0TErX4b/OZ6zhJz9qc5ggVSitP+j3TVcY8jK605Sgb
5ur/DwKa8ZLHsnVS/A9vK7Tx7ml4PGj/JY7nmwKOCLKyT/bsjwHqaOHb7Zqi2FXK
C+1wqdle1roOk+9AYKBSZqxnVo4lGASgkCytBqxc2kLDfEAyrtFcgiBRUgStdZeZ
LUj7t8UJp9UJ9DAzqO4CkM69KbkOva+3ww614TzoWdZlsk+2IBqDisomSL7Brp6L
lRMyLSEzIwcAtEm6YP/JhleOeB42OxqHdsVOfPPvw8otertTfaFT9d8Lfqr6B7h1
bLv01VYD7ZEo0vrHML4caLa1O2ocHS07x/RdMxVtulFyiEiAgwj2fxHyKT5yC5AM
XJ/++lo8wsju3khG6GALExmXGkoVn9SXfTEq6+scEb0dTciCXHvHqJ5E8VBEL4aX
ZxHv3ZBLeo2I6C2Axkx5MgcnYaIDch9I06Avf2toLX2UtN97WKZSQyvebd9pvq8y
Xgics2HtgL5mcRA9pCVQjmzBLwA/6OnJrVowwx4GGUi1EzNdZ6/J1VaQnJCeCaEY
/usAtRBt0wm6zdtVVfPZ9XxDEX0s/Tg2ed4gQVu3FZqb6+nR+E4DOY3HDQpta+kL
qxI+eA+4A445oF6cYQbl7TDAFz//aDzAmzNk4HVrjs/FwveJl4t0dS78OKGy6NFa
c1ItEKk0T4FZdqVhg72jIeOyE8P5DqrE1sADv3Bj+2hgrP7ULbJAyUHqYLA0p2dk
HIzzGXoi4vmArhjLFkI1re0Bzjxzxo5NUDhSai1xIOm0ahUr9itiCacb5vpOanAY
hmS5x4cAE5AMJzaSbxySxJqD31i4T/m4+BkmSpphpd/OWeGBDjtWYJEyyJTE+6Cp
I5+kTwt8xzVbRQyh+QDL+saAF4a6Dvz54p+POyI5lUXrryAp+onEqTGd8xUSR7YF
qSZ5oeWD5swHXOrJrlzBfvkwSJ+0oEhNqZHntsohjDYsfc6XwzDJqUDtcm/IW8CQ
0YalbnG5MGmKMKbWYBOj9n3x5IQuiarfRBT1RQbaJXUaupI2c8R1qIwtAtjVDoJa
bqrrwlKGFSzifYnhpCGTsttR9gaDX8rO4GEMykRwd6FvZtHAg0WgOU/XTQtk2Tbi
+5gaTvmu2Tc8xhKJdNfWdLzp+qhvGIWUfWj+khyAPf6bd4E9bHzzE1zSFFJhuObG
Lp/e6G/XTj4tKXQBIoN81f7linzpSozONPbVmKR+SSmkpeJ/pHMAaR/8j+Dt1kf6
EUb/mrgWFYWuIl4jQO/hs45lPa8nfGt/JG4vXOUm28P8QI/VC00kM1aqxCk0hEq8
NCsHn3V28Kt2Na++iYaG6lNkYidhwcXz0q8XXk2MONBisy44pDTZt6P458sF8dqG
LJvH4XfqMjMSykXr7SbyNbzwzComXYnQHdl4e7X6YYGOrfATQPfOzUL7ClOh+BEn
awNeKKZRRHNgqj8+ooSq8dXrWAcjpD2p9WNfwLCGed7vGDs1IchB/3nS0LF9FjXw
7t5pIa6JbW0gnLwNMFah8I2y3Yy4TNxgK7ijG7jGRi6NT4hjZ1hS1/tTxviFaok3
IT8ID1TbMJqHIPJ/iaro/M5jkKDecF5MgmIS3WPkl9LuPx8yNyHjyM/SYiq/QxSl
iR85DVV7dCDqNmdYjtpk4oU/ctGrMPWKWURIi+KGE1qlEART/OHOatSqHK6kDlZP
E34rygKm4nbKznBbszu1LMpEWO4v8RtxgsyuXJ2gGZKY7Hv4u/pcMfwfllEOfy5K
OhNnmzsM9ruMPwce2kdE3KliTrXXwjr7zCi1jibm3p7bZvOYj2TcFVJ54Epj7GUN
VWtlKgyQu4bYo840Lh9Tw6XUTuwPnCo9C/H4GZffU/h3TRNbTfxzAZB66jcOXDtg
NKQo99BhKA1bVcMTwpbxtxWWSQRFg0Gn+/JUkSeNEkJmWGddSY9l8pTRA64WQX5a
3OtrtT68DZdKzev+MR8ZmOdWVgSCRvMFKh2bqNWOwWSXou8RRT3xf6aKhCYZ4MLa
pue7MJGB8cnp4ecE0+0N+2AzqE7pno0OHVkGqB3FDijtLDkvyBbaarsa2cEuQSp5
rac0O9vuL40eTdWqvKyac3yKW7w/qf+w+BksDqI8aPCpcMpiZa73dCci22P3Zp/s
r3kh7CdVoG0M9ADzJsjAaTQgDiP07YQqA1tIGAPrEfcqKglKxbdEMbThe95eW11h
ICC95VtNKi8ohtW6qGNRI+y1eQifTTz4RjlB4Jywgfz6IPoHO9Ctfdtz5KWOhmHj
OUwprygmgtyBZ+7mRxm/vZGBNl7zOufMLnG3q2lNHRn5hYZwnmZVNrMGnrvh+9Iw
DkdmLynOSOYU4qYbhHPEBQy+831INhtD2a49Kr8UaVyjTPSa2mAnf6lsXlq6cMBS
Nsu2NakQO4trH+HoECAbTRG/oU678MQlqRf3OomlpIGAg8g9kWw5F5yrj1DxdG6e
t8qvj+ODXjua47fr4rO4eIOChdFsFpPUAuYeb7k4zw8w7gk+xLJHh+aD6iIjMhHx
vz9aLIoWMa+invQkw+0Zi48iVHmGH8UF9V/qIJcXWZlDxem6zx1l7FZczUjIWp+k
BxH6J8HtlF3PTbTsnpr3cqQeY/ASVorYYoWA25szc2mZpQ5qwom/4Qm0T0AZy8nw
0QaTdaR2bUliiWKwNBcnjXXYSpa2iU4dEZ/dh/3l83EbqWGtScBkC6uS3qOh+ade
7BO6z6cY+QazF0LaeWICIsrmHNAaanr64rPIX4Jkvt/hrPYJkaa55ABXcSEmj/dz
FlnXiHnPiEn7RXb1iQNGdyGiiyR/aP4tV0glrq8480ncmPqZNLyvI9ThYuJNyMc/
EQs4JlzYWd7nU8oo+ZY+P32kWnVVTV+XnD1VY+LK1EqmxQSDEIDswFhtyEdFqZe4
76yVhsV3D1LHmHczUoMas9YsiZ/wAhr+w3sQpzpk+haFtnPwPswru2kPTrpjnll5
7wle6SYuR2OiIur8rlMMrRwfOfcEWMyLUbppofPUoNXtwLx8A+XLI/9OD6YvpyXU
UG2Dkg3imkPtNPElHF5gCqOTLj+zo2qs8LbPCbdnE3gHIwecPDek1SQFIrIxzXAF
cwyugPLqRvGRcg9IkuZATnzuMg2KD64l5OWHi3kDc8l0u8zeKYQ6wZAQO1Y0jBD3
Lco8AWZFMvkW0Tk8NZPGxgqaNnrLC/3H/Y2pMMP5fKLmdCwjtsR30WAZLjWtSwc/
noAlIUVYI1JQL7pD0Mmf/8DrZCS0wcL4wHK7XLzSjF4pAAQYNFdMl9cCmntl3OEp
NoFn8uW7Qz0APkhUoseKXizMgyISAkcd10o/ya2dq7O+tOgoZGI0b+oEEPrEkbGE
op7tiMoG/wj96OADV3hZlX5JiN4qq3BExiPZ3aOqVvepkUBqd4/uOMbTAf2c7Yyc
JY1Vawv0icI9TQOCIHEFpyVzolCRBvxYpBWKa+siWKMpj0Ngf3w+iRismow4gQbd
E0Q9f3iU1L17hvOSBiExeXcA8A7NyA6UKa1VShc5ossxGgZTln5rj1Id51YvGhF7
mQ2MGwYIC0yP+NmQ5b20HD86B7i5A1km5ze/1dKh6a3e/xlnznKHs9sM0GQfzNZ0
XmHtfv0hk+wEO6UcptpTT9C8GJgP6niWILF0/gCG9EWzmmXxcSAd8ANqWbmFwgYd
Sml3yG1tMKpdaUNzb6Y8W7IUbD5NDO6iXnqhaQE0lIu+m4qHoBg8tLqyepjoLHND
h1N0CoGkAVPzVB5t+96o5qTW6VZQUgHXHFcYVf7cOdy/G4gUJQANdLqeH8Qym1D3
Yv1egz/oxODKmp/sbq3y1E+XzIsLCiS5kr3yPdZFIUtwitRxQgPI7wz4CUwSEviO
ia0qTNHpQqrUs1iwDFOhYk8X8ul9APaUMSGgt1rMwfeWlKoeyf81Q0o98P8/j5LH
yUf1wBe0mthxKWqrz37a3E5Fb8BijbOt8uYvHmDDA5i9fs8pPsS+oThu/qRLKnjE
lH+sCko9MFsE9cPr9TGzqiQroct/6XFvQCJD7jdb86P8q10F29gqKIwVicu3DrmZ
Pz4Y887vnqZnmjvm4Lplni1xOGHS/jwIYVH+hHXZzMLyvYtr9Dw+ALomUKYn6OOB
QeTUQR6Fj8wQVTwokYfmb9SdS2bXCqeXE8tlpWEaQXHRclb/JqLeq7J5jgXv14nj
9GXXCphiSpiwldeWMqkwOBd7hd0u/kYFFrli3E/msx3EbckQ8LMa2ORee3dGI/TQ
3emMGblx/FcZ+a9qk+xidEOrnCyJ4BsFlghqVO319zRWKAxssKRVzToO+CQyUTEC
/jI2XcDoensYvd+tYvwsV2Juw5EqFudgWTmE/nXAkFntch4NZZIxgiVZltsbG+Gj
pWrRiklI0JgWwsj/PO7injBtRbesUHHKiHGgSTXxoN0Kyn7ATqlyBueb5Avstr8v
HJTmgE3DzkOa+K+1bEpg9R/bT9UiFT2oUYKNn9p5GsYOd7IxXhp7EB3CwUsUGjpI
6C8ONeyXmj/fM/FQBpXPQMNqY/CEl2RmtIcf+HUd0Wb4L5ll8xUjOiru+N/w4s2j
T01+azAG3e78iBuhlmOmbD4Tg+PjpkbB7aAZekptMztJxpklNZ+g47T2PhYwVNGf
0X9tc/z72ioChZMomzQp1g5/nqWHYECqzCsQXLdbsd5sqxIrrl2FRKe2hhGgmIim
ypKv1SIB47UevvnZe/U3PRsBQ0f/EumeLgEJH7Fb8RlefUtJl0FTatbXZh+NrobR
VDoff33vr/TtnEmrmkNQSuGCewKzTl7HlxPut1CYn42KiwfLKUG4X/TZhiJQt4tX
5yGmHq9HyzJi1e43Zsiq4c9PXaN+EksqsHy9Z2YvZERzDI98mSjzw+8m5g2MrZ6z
OiIIL+zH0p/8YQJ7hUh4s5RI68mSJIdDQrurUYs0byvXg4youPqL2So8IrgYzjLm
//N7GDWRzmuR/NZ43S5EFMDEM7MZTFj9ToZd5Ki7k6wOhC6IdsoXxCgkLqtziNxu
zFgZmhKn9xGYPvhAD2l+Zz4afAlZRlEmft8YIXev0mRqMMe/b0fSFNA8RfZZY7/C
gkgDUeGq3nPpxT3lcx5o/u+NJEqDMVo2HXkYRM5XJ9VL7Zhbaj5sB1szAH4l/DZ4
Pz8sDG69nu2biotWRTMpK8MKApgDC9vamOId2hTzsubLvPUfeCQRql6cuf5X0Zdw
U5frFDgTk67Vllaj8Sdb6RCdwXc3TDhhJ7wjyLhdzafX+7LakBe75Hs7xBWC71CA
YIhX85J1ZaN3Vv9fiEm0VDt8iAuk5vYvDaBoopH0yrvOltW7qphnGutJ5Br2pqbJ
q/0DNHgy+QrZmXZn3fwbwEqsVjhgAeOjErjwLneSBL4u19tWDjxxIlBkWfkQ3fLY
v7/2HrGXmyiB89XeYC/Ew75+ph93+iH4dU2o5l6FZqE5jfY2ghANe6lRI0KWjX4D
f+06xmYON/hD3OaGZHStarcUmWp63Be/jT+XAQAOjYvoWxkpg27ZuYHgiYUwSiwY
Me9AtU2NyGkmPgTd1BksBi7GOHSt/mcn1KfhKTQddwT5HEYf6nnU/rcsRMd6hm72
HFidD5dOXLqWxURg4otNWpczZr/wm92sb/OaAzLUIx0HLW3gGiYy9KFSj+OEIugE
3Z3Ug/F8uM4PyKigPgyFo+pV91woh8qdDei5YfZgQ5lpN0e9JncudG+cLUyvbbNo
koFZUE+6GX0kv7UFgFC2qU0LE97q59orhzQlrqXpqVCpG7l8nHYPWhysYUvYG75p
ypA6Yw39NnnMn79YIz5lKTm5SOni7YwPkc601YUZtV0y0J9gwn/aNl0TM7tvexUZ
FCjM+AE6e87RjLZWqx7icfl0R7J2FLTK0lSRMez1TDsAECG3nG0TwHHfn7e4zgXQ
mCCcQd0+KQUgfBVGx7E4yQAvV02FyU45GaQ1Pa5wvy0QC/ivc6ZLxUFFYoExpAfH
ZZS+XEUxhRM3r9RQF+xFJdRue9ivRONw/vtRbt0xbhLKNCAMThSAKOxOY4Z/xccb
ZNLZtqU7EdBzk4VWV/d0fgHFaDxW5N1C+9SkhrO3sd2LggKCKlc3P8bhN9M2eUWi
ZGcmK3kdFpeMldVBTC8oPrw51QHB9ZFbcyE88kGvLB+LQHOaJIE6Xk4PzSxdFFFY
UfvJTZVCI5C0ngVQpzyzgyO3iCXISeEjoNmm9nBL7mXm3d8XsYuDdolq45/HbEtb
b85UvZMcMORSRmqOHtf4+7sE27H8UmzHmMC3hQpeKmXIaANjSonLL2Utkmh8hQv4
NMxEU09X3EEJYY/FtWnW0Z+0hOAnn9tNDd3/lUK92OtqcnYf55YQWGEUxALQKWGi
PabsEsHN6dxONo8Mkl2Qyajt/Ou8TDc7gu2EjSTaHsl1kjuh2U2TyqhfDBcRrwZd
w9AkZ3jdUkEW/M4RanJ+d3wcrpotz8OIbe80AwZQU6pEI+fUcwo6HAyRlr+xVqfy
cT2DUaEt2mRfmtJuA4ormQeQt08gZGTF4TCcmPqrUH15kbiV8bl8gSbKOYU7nTLs
pKE+I59NO0SAZCyJFP7HXbKp0oCIlVy55sYSymBGXaph7ASdcAbjUsnYwNag0caB
u1v/zXzKsaR1iboKNUiL8cLMwl4zTtqhEOWw/Wrebd/BbE7UXi6w1Y0chesxpzze
Esxqew8QdB/S23v01WPdLvLhwDYeQoLS0devewK/RMBHi2bVxQ5NHAutKifa5muN
Sn8TELJCO44h49trlvFwHON9f0V7uVpnDrSQQo0JGJdg+xo0eUzIAMaFAhy6/cEQ
m63JUC2m3G7YHEmP2s8w1MC1+5zUOyy+T9idnOm2+FSSFCwGKThiNLev8ul3qNlJ
jhHfMsTaXGlv9xoH8J6YgHI6teaQfAK04fDbjyhih4WpRW/NNBF2vz8LRIgHi5lc
N7XovR3HPbzEp8qpHAf8TxnGqeLAK4AXQ5mlI7kAVEGr/cIo/zMBr8OAXUiWfCy+
vWlfBRfFsqjDIAtsTmIQQPwW1c2SpWUiGAJkwyHxNqNvKzdTICRIxpUl+m5KHJwA
Kl4CzOWXovfcICVtnXwWuyHUTwHYMz1iST3P/EoqTwCU+Lu/DUVoEEq/XJ0uCICL
6L+wnFZ7bgeZp+K4rVa1yAugQhPMgBcjqyfejbVN3CqrKmWr3if10lFa5PP6l3FF
JbYsEVr5nVn37bHfzDUcqmvY4f+68zIa3TeKAVg3PaROc75JxMtHXE38sRvvGq7h
ytcArSbvKc5Bvz3Fe8EZrppvzpR0g+LhjJr5X86NZNhi9mhHstNSDdGvPYcx676w
HHEkKQe9N2B0ciD+Qt+zkZXViWQSHu5kYNjk1C3toUpOpvpkohOR4dkCEZK0E9Gu
Hx2B8D7S5wQHs+sUtNTdrrsC873jqekwo3OS3ucWTlf8zxw5WXD0WJuulsiGhdMs
BrPFGNRsrvjabSYUvU9Kdbr6cu0jp3Hy1jQySqbtUIR5EflXQQswvY9XJpbuCqG4
/culDC8HbYd7wPo/vmqw052P3+4oaI7wlHkpsI2lajXPlMSqV9VctuTcVldWoLjH
zwhwgiDzRU6uhE3Y4PdWAac1+OsQ4wZmRz/TiQAOEZqfzKWEbSDfWbUGmgF6bT2E
LbreuJaW4pNdwfrQMXyN2FTol7YZlk+IkQ0Owm5r0oFU9ysmYCyHhLEnTNgKb01K
PkTEZFaBbr+9JolWewFloCkl7LZOgYUGY1ioJjMyfA9zPU+eQ/cABV3MQky57MEX
vO7HKdqssmzLtp4al3EXFKxgjPqZgqadzVGsFbL4m3OQeh7OaYfyfpFOL20Ak5s5
trknEazrDYKgRoK/dfUWOAgOjnYv/8OnN9GCfi6oG7o2i7Wi3TXXGR4G8fnE7u/L
6+Q+0r1qGXDGQfy/dBbLA+4IDirubGunleUlC2xBzVvnc5tEdtME1JgyRUPbVN/e
pdF4Xk8d7yEOQc3rmKG52XaTaukxRizapXFivcSGeHxniJPFNNVrt3n/6Gj5++iM
GrQooCmeDSZrbVUjNpXKzzzNApm8lIMxzCfClDBRcCUW/XoWVcQj+GKFG9rMUVcc
oNLdUe1DWkuH6V6se2vl6iPmUic1cdwIezBHuVbavHXjzzN8OxCh233axJUPJr6U
rRqhNG9XB9/UOPuwr4G+/HJvzYgu4tqa0lsBcvyKOsMTSgRq+774TJBT0Er6n9nN
Mj8n7uw2fPv632UAdTEKAIZXyZEG8TPl0yTT5dwH3kgGybrvS6pC7H0dAxpHogjM
sj41NfkoBuXYU79jBMbqQJ+xvfRJyOHY08Zru159LkWs9btH+77+iE0OaKweBr6N
EHY8ZLbq+GQ1E84no7NvnAKNhZmXWXQ/Z/QYwhi1rH2a+RISj5kZn8f3Fo3rH5G8
4t/k1bHxeyX0Zxh8zQ7KLbncKAMjE1idufSWc3PYHD9dvPqtxGaswkVXGSsTWOR9
tVoJT07lXcYLsGDoUp9pRqyNX7jm6vldhzj9+54lyPo56F5SK4k9wkXXPu9SFcZu
1xUvVzzYqM/aYpKOeQXALWSizWxLohGAeEku00pIZlFAg5S6+rHuCMuFAMnI+9mb
bYql9yygnpGKlRSCHrraqBOi97FRNaulGqchZfcIDEL7DnUQERzCAsa5rEvSNUdD
K7XUK2YfC30Ubm17B2hHTMQMIhuDhkTq2RM3ccxEJaTqGiOm/devi0PIsIUjSxME
3Olk1YTwpJf/AMA3/kHUahbFfIConO+EH/HjNyw+5AWTMDg/EAnOFg8vEotJ5C4g
E9BAeNK5YjizX1UZHG7g732/C4TmbT3pv6B5DWtnLBWHob4GTU1uY77dc4ik3pR9
5I1U2eQoXbMxwFBZMhp1mJGFFCnDlcdNNDNoNuqtp3fk6l9FaZVyvmeEm/ePK2/s
HsX/zHJdOi6jTierNFTjNtAcohF4/JLE0V12NqeqTPyx8I+1vw4HHe7Wn3bHP6b3
zX1Naqfl7hKZjf8wLUogRVGYgj++3m3w3qhI4ND8JvnkKqCxnmbiTGFl00Nz73Y/
gQhwmLHCIwpZF0+ZqIMsklQNYmYrYrM2+x3Eqbq3Z5bacc5jdPOM3JYbf7KspzdH
zVQx8vpi9BOqrkZiwWY+g4+9wxC7nscPCWPaoRsPs0Re80bugEJqUGm9/3Snzp4v
CTyyzzJIBlvO72d3H5r8jgTu5wL2H4amG8cdwW9L4+5rauST+4vUgMhtpsSG06wJ
6nD7oxwFh5rPC4SRtXWi0vca1WiKvB4V2qW9H3I+OTjWmRX1jWHp5w+KpSbKy93q
hZ+CB5h59u0HjDl4jT42EhmuCV1chEgh/7AgUMN0KFN3PqMPDTfrWOjV3488TW6O
sDgy94P2x/lmwoLsAfXjMTfPI7LoQ6hMXwv9StC0CR343Z8vkFnbHovHV5PcJHgM
Gggg5gUsJvWikCfGSIoUPUkQWIOiokBkDAg6f66GHW3oWxmZ9lJa3pPykdy/tA2X
aAtyseBnYqo49MQ3tfPYnkmxN1pyETKIKeVXkiuZdmAUxMz3KO/TIuKmsgBhX0Xn
wtkF5g3DMR2MnspRpB/JNg7zrgDP9cfHPCjl/pHadpM71Gg0j3di4rgQDiq9Mils
zvjeI+D3TwhRK/KBE3iZ5t9o2SGv2ZqSeAB+gdaWSubFTY+aJYBrpLcaJeLzS9O+
c6+ow4v8vkhhC8BWl8XknMwEVIE+SdEH5GXKM4xZ93iP5xF/W+7vgIZMQ0sOG17Q
nRVh1yn5PtK7Q/OHxKoiK1utH9uEqYLRyqfZhqQYs2auyz1gxJXFbELtkyJM+5ud
ECjsiSQKK+VzmYz1uMBGCm6DK+661higlHrFcFEu0qk8bWxUX/iGiPoKBZWJwJ9W
Ym0JNuk5zz11lG20qJd/dK3CYby2jF9J1QTc7jfCbBxAzhWMKwJJ7GLN9To4qkYb
7ANQmTXcR4YwgWXagtYErc99uH3hx2A6pKIq0B052MlOadjp9IRI03Q29mNNqEZ6
QXhFuCrDxHnimfFAP73YFmx3twp2vhX5K4CSkcPbqmS+OYvvzCEVVxYRsOWy9uIo
bQ2TYBNAUcSBBCZD1HcA8ycYf/u3SVbyhz6yOK/dUX0oVUcb+PqX7Xh98KKqzJ8c
Ulg4vOjAkIuQsV9EtmuiD1/4XoZX+K51ElZemTGAbnpKEUsktE/zCK4L2DOKX5Xl
W/YV6JxEyGkLy+FCbN7XbhQlkdIk3ZgSBvAhRw2BqLCUIFh7wpRGcS3wFNZr1mjn
H+KmXJiCxq7RauUWTYo+X4RdgZWh5gLK3w0egRVzjziq3rHQ1HwUxQ8/bCo5Nwdx
IeqsoZCdk1G6iZey5ZNKs/mYGJVllcS5XYERyV3nD2Od5YSftZK3bp8fgdWBylQC
6HoyFqHElms0gNk25W0KLfPoo4V68xmU8vbbml5NBpVAsWXR0UBJooNn+egdk+vQ
iY5LRpjCaKJiz16LCoO28gR6m3tgyEEdhYZNB2VErF0S5T4F3qXUYqbvoUsLd+CX
apa0GRQESbX97VmKt7vyURIEyT3x5mysJGH+O0+A4maQolslruyC1rL/5hfzrGmW
5hxu+toc11wJypLogZvlusxLubKVH8piOo4oAO2XZafwT2dXaclPRyGoHbMfemW/
mwgpRjUVoL3fxCzS5IYCbpwHmfHW29Dpj+C7TTYtbZbbK2chF0a+a3oNg8lRWOg7
7hwVkCXRw2/JHcQMpEBptE/LUkvjdvs+Ar8W/KwqIa7eDfTlMm/7lRIj0AXWm/nw
v2UF1c5EPBA5vyQAi7i/9zdIcC3q9C7q6QHVlFBUO+uNGPxsjin54kxCQSr6g0Nv
GC7Vzdbl0ke4wg/K/SxSaq3j2aDrb0TLPFOVgmCexCrshKpU/dVi1HdRnfnEBJcl
wtWL2h78o91/j8vrHdAT5/ATrg6vt9lreKAia3Ona6INbDmnYxhls9oWnDabCJNi
ax9kmUeJlkvwggVyTOhAk6+C7AvFH4rwyes4PlS7EGjWRjhuOB9eMzS/zgU6zSl+
Bhei3qfnz2UEs7Ay54OIYV7y6WSzatioyoxjwAVSrgG90FxTbsWC+sEmkgMnTBR6
D5K/hXn5DJ0YIwZ6HNP0kF2owgCiVebYZ+LbGr6K944ZITlBpmz6LOoAe9wdi5Az
4zZsbaN5JeH0OBrKKFa1M8IHaUehdrw0dzOdh1h/LwqxUfIa/SC+ps56VUGkPJa0
bNaolOMZHPdv7mwbgtEQ1bww4rmh+b26TE0PLqosBINDcu74wGNAOW5WdvAfrk/+
FtCoZP7RzXLk/V8fzy1jkJR079d+EcxHiht3wL4nyfqS7Db3Z96BULATMwMng9pS
Bq8XnvHUq9u5g84hipxvnDPZEN/lGOULTBlhfkIEwC6/aRO1F35oshdEJU0p/a8e
QM7yA+tGLzMz2saFHNtd86X/t/sNWsSTgx4Jpa7G9IEVkwTUM2+LsKeQv4pLUY1Z
QcKDAdeoVvgZtqoAh9fkUmN44VKzzW3TEJ31bM5OgJqWhcH/W6yx+y6hoeU7hXR0
Div1JmKVxuRXFHori/cTs5A5ItnJdES2yY5xwwLJd3cREUJMdKTbi14asqB+K7bh
FuTSW2UPJGV368+rPKqGICeMCXz+L6XjnRmKeBsrz0WS7s6I9m3mDMkx05hLPxpN
f+y94djPnDiVeW5W5c83zR19ctp+CLQvL+M/fYXZB0G/56aedHQjIQu6ZW7CcxWH
ZHtRChwZK81ijNT2MgimOPX3p6ELUclZ19R0DMN5rXb3Hp+neyJsH3Bnce5SI+NV
TgWP3nWk1cci708IOFwNX8FdK4pqMvBZA56myjXxrh1UTTHSaeN6TFvbNLNQ7+dv
XyCk/jHDJNfFJP0edHKmrGRRrjyVULjvXNmsCWJmU21l6sce92xi3Uk7SSc7UIrI
+YlAa62oqDSpL4xutzwQf9BIFv4tm85c9olY3ApYmIlmG/dbto+101GmQAc+rXwr
Zrs5RcMIdHPUdFFEhXmfSPG8vTcdlhElCxZX/6015Khw57AdwCrtYKH+5FS6xpEO
wZ3TxpKWK2pJGWl96eu9JdBwIChNrP4/7DJvPcb9c8kn1RdkcJcj6b16ZZBKSQ7P
ANztpuL2jDgUks1GNQjwfD+UfvpV80bWdN4IFJhdkk0trn3sEqOKyL5jQ3qmSMMe
NqkpTfb9/K7054+mo+PhWS0NJyc0F8etvE5CKzCL6u/vxLR6BMXXMKbfdH8uMbrb
tsIAxPis6qlbBEzhaaXSByjsA603aUs0hMiDAq4/TADloGyQ8KWcIK7mzIjmLb4b
N2NLKGxO8L5xMWS5ZE4m2uux2BY7JU4btl/vmBHie8GGI4cA1S+IF5yHt67RZ3NB
U15hSbnAwEfaMTVo8JB5+VEOQXlzUu4VWKLhfE3p0aghMRX1v2Ofy02CMPSobUIz
L2/Z8BdYVVoKzravCSPUDQTwkLbizQu8J9myf4CAC+zHVgKa4rNsDIGkmGolcL8v
J5JIJzgGvhdNWnhNLaIk5EFEx0UmRyoECqi+VPoInfDKqT2SLIo1Uwk4+44sZRSG
YPScDErgL+q46b0s2sGbtguZrq3yEJIgJjWWoWKSk/gtTo4Z/ai3S4cHAkHZng85
obsDJITG/fQR+LbFJxtH/vGl3o+VqM5FFYDQtnOo8YC87yck8FCPCHaJyGNMVstc
dyKmUxTtS4K3F4pH+ysfkpVAWEVVsy4Jukz8EBRb6eI4pSz5O2AzGzYS+t2H2uwy
lwQVOhOiUok4XA6yYu7OAhvRWAsA5tviKcQPYD6zTlsBv67rnY/CTBaDLpvVaY66
4CjxLtvMYpxF5Dltpcaac45n1nDGJF0Qtl5/qwGBtJVzOaNwoEeFNxkgvHwfaLLL
2x9oMzXbIzuQvDFs5V2/sl9KuxtiCl2QwujFyhRAGP++T6CdWd+mbbhktoPM/J5K
+uHP15NEY7vxqdnqPntEWwPlWhSoY1NSL02OTmW3lMea8oqWbnbllt1Tuw984HD/
cv9oCg5y46doHpU0oiV0cf3YYVzlzwtJKIHZBjoRkM8UPU00LOY6QrXCTdiu9MXl
kJrNQrPdZfLlq4itSoPBx8kP8tG9/9lcsDHiGdF2yeuSq1bt848voVI4Ox9qkqc7
fkS1RtNm8Cy8AayEBNG5x0k122CZRnPWw+FqWEY20EMIZHHQJG6oE8Yo27m+R07Y
5Ngr+Hs/Xsu5iei2zVC4YuPzXcFNHqSJBZYwhCe9boLIjE39mDyX+Rvoxj0faHME
LyUBvM4WO+O+mrBZO3ddEbl/1ABBGf/0DQ3V/P/x2NrBrPZgnc3zyTRh5+fOc3CY
81wz8iQaqGBZOftV9jm/P+zHCBUqDFjsXIIGqAkPLplmRWVGp4YfcQCUeXtoXlMc
SBif6MQtIshSE4KFRni68QJ8AEPcMg11neDMb4boxBhbkmcj3yvCVzmaQaWbtMCx
merWp71PTJcKVxoKc5vkD07lrNbT1CRKSmcK5e/kqNIn55hr5oAAcAI1HXBRGK1+
kNT5edOz+4Z6dcHBFAElVC+ur3Z6A+WaN69Z42PjQK22lFN2UODwKQRJ0z/JlSsF
yEvSIfwl778ydWr9sESWekYty0Tzn+aWXV6por6Gsra2W3jmhb82oIgFgU1DIdS1
O6w4oW3yqman+VgHJ9XXLdnjpwTdmGIV5cFXs2Eo3uRCfLDdJECkFzMjbNODvY0g
60eUFwYTg/PlWV5oimQMT+L7hFQnoxiMPBpvC+kdp4qDq5h7/142DPdIARAdyR/W
xbLZC4adricUGU9QUbhQvyumgyoMVlVHv+Av3iAsYRESN0M7jZOGj2Q7rMXjBx0k
DLtL7rQSKebjRpfaTLzshTOLrw05vfwUN8EGcTEPI1Rj/nzI9Ny0LAxhKgTnYO9w
Azb4vXE66aqExpvfDSjNF063nnQiDv3mF5Ss/M352fNsiFf6yqlisBiLIDbQ9Ay8
F4uyslsvu5iTgPFeXGyhGC/AaW6+vLQjRlt2lRMbCE5MZWxH1zke5UsH9jnw+Ih2
9C+heQ0G+LWmrwqEKRYPMA1dR2xRb0YThhkdiEpeWbCb//aueQadH+UJKGyQLPkR
4MNHwuJ2Dah/JhRkrjOvWJ81viRBw2q9Aof2OxbqZTNPGyZ57DYC/Q220qEU061G
8sxy7JUhAOxbbIbZJOlDD8x7zeJ5UAZuNMDK44yBB2LJeCUsumBgXBzNyxlYVP8o
L5TsZJjEZuO8oIIunO3eb1aJz387kZTPteMAxdOHzIQHeG+Kg4DZC7y4esSkGkKr
YeWmjIo3hlkVgym+nEcmwcyZnwjhLrqEV1JD/tjF5k6mRiNKslcLh4gnsuKoYDIR
03XYCYvLVNEoM5gA5lx0GoG724d7lZEIESf0ll83CTqSr7xxegHgoQbul005Nb69
zY/jhUnNRef83RmXtoKG/l3UIcMRPTO0sMJA8hszYHf3MhuxXX2rQ5tvBRbB/d/0
o2zTYUUqpyXMIKAtP2SjrftmDknqiOSmpjp+zPVWgdkYODTZQFtzSYsjJH5l6tyL
cKJSxA4ELPELwWVjj9VF1ihAbyhw8oO46bRoSRVVNYpqRJgtGm8UA1q7SXTdPSrL
pbTBf3sSv9vEdlARt2LyLcBJptzkfmWkxI2sEHtO+42tXxPhTuebsLzCcXwKervq
N6itZ35FPPekIOKH/zKnB9F1KSc3GaxTTTPacbo4f0qsYo0YjGu3HpR5ByPMqQKO
/NEslr9NALJREpcjAwLmQjjG3hf38wmTykjDAPCoKGu+9PR3lMU6A1i6kLPa7R3O
j5lk5X0sXuEMEcGJGgPBipOUP3gBMR8ZG3e9KBmtGY/Lgl5lnpCIhEhc7xRlPfxM
uWR8JCTFpDyuDRqdBYYxm3DVeaMgqTz2mGtHuCWgG7EMoTQ9ZmUXhNmG6Iy14xt4
qzHDKcjMyNwB9yQtO5f0vmLl2iEV3vhPwhRDPqBijYUcsjr1UP2ByVeq4KKUu8WA
/5qOeip0mylQi9UNTpoPJhOKn4kOFD1Xygeb8/xDjJ0U0YedJTBbMGW0Ia2HU75G
hR5JCiq+ciOPWy295HqTMf/OdoiwQ1x8GISCNyoblII+uNHLJ1MmSAZMFri+A+oX
8jwC9aOprNXaZE1jUYPEm1nlPPP+YkBqoMG/F7Sm06aMYS0LV7QnCrQlwy1dRa7s
6SBLBNHMESpN92dks0WghJDETLKlZqS5QPpsdSAF0vBqjVGGUOpAIYMx0s8mqHKn
SHqWa/Db2VNE+8yBX2drLjLw8EY9dM6vtd2XpVjKMUp06D7/fPisC0DlSM2OGL/I
MbsNw2Mwj5AvgAytopD05ud9w8ZaJbovqFz3QFe8+27BefpJXvgnLaiX+wYknbXi
LG2foCCNrfBb80mQrXDcbVEl7i4iLR0CK8xg3iyX0d4QU7GXm4g31GIgcyNkAhNN
HwHOad2pzCs7HgYVUVbEmkhfpKyPIw06KDDUwrVk9/R+zYUdtaE64sRFV29J+3Oi
vISlic9fggidCOLUhQ4gO9S1XI8HGyWh7AjXs/oKKBEiQ5dgFRvckp7Fwdsu/Yd8
Qopb4tBTLHRtW0jKMCUN2GrUR63r3W+2cRgki44fVXuMytccumO3jVDHQCmmwMus
7SqZ/WU36EU5kIVwGrAOOfBvBBJaAUKTq0u+Cxw0h//tycTOLe56z3NT1lMdzZze
vOCyPBCxGorv3TC/BN/cAOrQGxh+Kbxpr5JPR43W+X2xbrSmhxK3f5AttnDR59//
oRzAIuTNfXWqjXhGZiHZN3G+XTN2EFVQsCjxJEUadxbjt9HxQIB5VkLQLKExNwBw
z5I/wq/DgF9PCu7o81FTCyoSZxcaKxRVdn+as910368iEjdm6emVnFGFvZjvLwId
fBPTXgIIqzM4uSqeSJ2WKQdRZZBU2+h1XK6cMOQe+ncZQF2CXK40hnv6D0ucD7eg
5EGaGKIfMhS1dPdNrxYR1SBm32ELjzuM66gVo0mEJygxpeEh4mvMbk3XOAe9aeVT
JiDUmmCva0+fvPbcyKiLXKzMnAEWE3HFHv38dpYiSn49dBlhIp2Uwx6VdeTswDx5
M/3RGzfQYFvu5eJeIaFqbxfOHHr33tPS2GFKBWKb3Gc7LJinhJVplLKzLU93eCbB
rP2er+r1kPdbm9yjgn9U6O3NU0OPt9WNsFAcehCmJPdgkbo4+Nbj6BrURRLu6jIr
Oy7SVZczUbLZsQLJvtG6QL6kI8rj/uQx0l8IfHAcRBUc/CHRJFaZfG9YTj1X2MT6
SMXpLSIs6/NytzrHqOJUuc4XTENTeY8IggRHyO4M5L200rWuLnPd9R/ueobT5dOC
43J4otZelny7TRf1ZtdrsfMS7tkoDSBW1LP2vQzJnRtDq1FyXMj0EQ3sqLU82LDW
oatmAKN5EJwMss6uEQOvjJsA+Mk/GCWnMag473ULzDM21UpoPpwzjMA0e8eNmOyX
Huq7aB8oYUUomRO3TVopurd8aB4kPNxRsnkjQnPJs9RmTGNVPq0HsSdBGIl0BSb9
o6kqqorahTtsYTsIU/GZLmbaGgxkq3nlDXv1kIcILCtNv3VYRR/H3myXsn9vBJB+
uzXMnyP0rql8DhW7PIx7Uxu+AFMg33D+u2ro6gqbMeNA8zUNnJm9dqM1tIhKJpH4
VZbiX362yB3GlUmYBIhGxbr9kKgz1GTPWKcdij0N0NDgfwvIuSV/kwi0CQc81TsI
SUf6zKerl8lPG1AxV33a3qyArQE3W+ym3ERCURw5FRksbY1Z4rMrV5eTLFEd/XlJ
q5JTWe55Zv+1lZYD4ac4xHYhpwdozk0LvfBGIAqPQO72kuwG6/L9CtBIJ+NQvjo2
9eDl/znsFAwnxc8lsb/Fvyph3O1Ld3DYhydYGV/nbVc/I8qbY93mCPWaLhvCsqS6
hLW3uWIErCU0zs6YkCrB4hpqrc9vTcty5qiJN/cXpcctAVaH4ji5YSPKCvq5aMuE
XC6pyP/eUGSiYMQmoO6b58lVtICQwFv7X5AJJUBjIJz24OGI4xQl7O+1+WLqdfak
lFRQCK0vRMKHUx25CmkuAuV7PHEZ5Uq2WzMbyqQaTi3Egn+ch+jFY0h/qhbGiaZ+
J5hNFiTKDrAV6vQ2RLMguRh7HE2wZh6C3KNofS/SPJUmmOC7tBdgrzwP+gJ9tgFu
95LkqumEOaAiSg2qBVkWHzsM/mEWgkvBm1BO4cdaSlqW4DU1RTtB9ACtGL0XOZu1
1uPZ+Wc9KQks8/aUyi77+0rsviMClOPeSHX1aBZVRX/3X/GnjA+tBN5BkvCDns/H
TRI2+XVzPtqXE1hzs0JxkVFgdtIprX1HJXakkFw1zK98UEullNsuYqyZHyD84+r+
54DgfCOtvnzki+2AKhAK9saQbzFr2C/ZP4GHssAfm+9VLLPoT8TQtcw1Pjx3X889
ZsC1gYfr1TxlZyolY1AFd0Y3pc6PRPTaz5fg0K6H2zT7+sy/mtnHjuK1AcNP1TfB
i1WayYoRM3rxkhzR1k7IxqLzkmDgx0Zbom/H+Uq0Gqdd17CzOkULmnIk9yGjAWOl
5i8hk/5oEPJllec9l3yfbJw4c7aia5Q8TgMWOjAWyMoGlgDErJzlZiQ79kJVYXhO
YWwvyNMSVbZivktFR9oM7Nu15FTGFYeA14BIKvpm0OY6pk0xbQwmzaoda0oJ7B54
V0q4UNJEmg8VxAUc7dC9rTXsFY8Ur1lkjEz5yuOG087E5bBucfOK8PVY2+pTdl1/
bgoXytHbj2HAXlyUh4bXrvPROZ1XPQCfLhrJv8ZZlxq2YqZOL9IYJKXjYeIlBYfC
JAmXQ5r3qJ9kzLVG9ByLmZHlM/Bc62dEZ0739OshaTAxp88xaobK+qI2fDgD4Kd4
hORt3FMhvWwTmSjqLIp4sWR5GwUDEjlRdXOOM68daOmHp4E/8npxZzO8i693x32F
r51QVeOwOU1YI28K/+FLg4YFQkVMlxAEP/YGUfkjHrsotemOcCleYOjMkMAF3wrT
pkVxECWl6NhtIwemhPS/nCIUljtSiUPlV8k+DFqZdNrKoO1RGBB2AGeQn4u+HjuS
WDkQI42TGiYu4FS8ej0flWMyKk3YZ7XpkiDIeOq58IFVitEvZcBP/DV5lQjVqjjt
MCDioJTdvogZ9Dtqkqe+8ffXEc2dP4f9621idCAJH31soQeqRuHNnaeSl7iTuQDU
/4VAufBQoJhAmAqsqRndcSdge1sr5VNnRUkI8AQzxhqt4HntIE34o/nkxRxGALWm
ObbGD4B9/MlJg4PpcTp3/LMj/M76ChN6InDQBNrhMrzjxeG1hH3x7GlSdIXph/pZ
Hf0P4M0ur5jJCe3iT5IITjCRy56GSp7Mfw4LGtELAzzBeM3BaeM8h7fLe8HUS8Qm
XfH7BdcQEd8HESHrJcH1dF+4CpLCdx8lzmuJg5C8mF4U+MN8+jCKyrM60Te2tEsR
qDTXxJv2yevaywq4Ztkh26lmIDXV4gg9MNh4t3Ji4+ojvSZUpxAO4951FfZ8MglB
iY49B1QZdNEcECC/ip/iILcALSsyJLyILX13x90XGjmRSR0s9ibxNUzfsefw5XYT
92vL3mytZjmptm2V1BbvNw8vTUx7XbcV2iTNU6Je+/v8SVUvBBCzhhr5bdlcPbtY
oFavKf55CDMt9wdq4reMFDjD4FpjGxpgfoWuKKTfvyn0TtTcWTTZcpmBTqSa2Hlh
EmBTHVKK/ji1otaXTFJ/w2YE+CFK4HqDxQ9xLueKTLKW/S893xzN7VEyhsCMunyp
0YeD2cLDYpWv8qKyNwxOayiadyIdf08F0LJBZO1CkA5lZLppP6e87rJc4C9Bd1JS
h9/tXF5rH4LRcf6xniCiRnBRt1o/44dBdLy0UqUBas9NOmNNI6j5yYebqWCAFbtT
BCNdt0WSQ6old7JN/PI13L4AKpuGgxcQicVF7DK9+Tuh2Uukymhz5Dy5JUbnqo3k
lpaTNH8KL8wN69MR5dD1YB1M1urF2ch8kcCtpDy1ZGaamg7WgjcX0gBuh3kzkbSR
4tXm+lRxFsGnBhXBSObwPVfmMUK56oWS8tXEPz6Gp7khK+Wd/UEKtmgMIYbGrsN+
qvq7h7rP7dqKAWsdlyi/MkoPjrOgdmIU/gr70Nj+bcQUA1XBxVTAOLbBFbSRdNcd
FULPy0gKRvYtE7GG207bB6PLZws6Xy/2Szs7+Md/aK3vp9Pu9yHFuTPL8yM1h37s
A1nJR0LHi9lb47XRl9sf/t6fI+w9Ota5iRlj7eW7wVdAJZkJrVY769mhIM0RwucR
JmzmgskJAcxDdPFO5J9GFo0dXc0oskUslkWP4cQ01FZ7veuf+eUY5WidLsWuqpox
beRVsVdgLjRSFNDtp8lhMw0vB+XdLpbycdrda/79X2TgetE6Q4SruQWaT6kMGr5Z
fefgsqpre7tp5wid08VdkwpLEzHJ0RBV99a1SmKyiVfRN+wVQU7G/9paJiO5+ox7
VpNmQUg/+kWjIuEK4HTncKs0CgH+bUXNdxOXJNyhLIGZNjfNeaQsSZMc5OFFIU48
zf2APzclJMXjAZ0yb238v8dLX4fx2fOT9Syw5J7NHohHvuELZ+MFQ87/Pbu/Miae
cYByMZOk4RfUSBDYYLh42RZU590vTcnPLL1xhwvvsRRu2WvohO3RmTuU9+IaZXAu
Mmv287vwSQjUXupfe1Ok431QSOGsT4OpxHvCBwFP5CK0/WSoe/k1Hz/vlJ6AL6++
1QITYyPCfM1xBj6cJ1aYrgw9BEnzUaTVK3hqpGni2g8q5fdcxdOld60HReY8vlzG
aUEq2carseuxHcsJ2EIqoaaDTLhk/bm5mCtW/e4SX4uyg7nSkJL6eXEjK889pk1d
wwwkh1vucbDmlQL/B20Twi6nMS1+o4Snq+hqfOawyMbibAzaIi9Rpf5F9yzfJ63C
7ugtAdrd7UPRlRwc+pExH80wmJrP4rZzEI8zkoe9F1sFm10+Q2ib6F1KrwM30Tfu
5sXYXT/GoF1Niv2daayvzVOUCooFW6VmBKU7pJeSTaRRJtl0RCGjPZe+lQtqxB6x
u46cM4NvnWfEzcFyuG0MinTYqAuP2Dz4EnXujhnXDizw1HwjKvzP6IMW0LjxJnSc
e4wlgsR/tB9m+kW/6F0f050yKH/+ddCg8vgKoK3zP3/I4q3JwIJtWtgrMPtvqjBy
V7nBKBF3loDbuGKnKX+QZRhnRyzmlCUpF0JEbC3BPNL3foncnH7VWfBc8pYKfV25
9wgTiA20fXa4iFctyoc1Dwe3tSiTHjkOFGupGs9GCF4rBJ44cACX5jFbZQ9UDeWL
nH2ZZLezA3Um9OVriR0ZjyzOhAdJkgucIDiNt2l427N+9GhI1t7HtRXRK2t4KOqJ
07G/Q4ij6mPPNEyl+GHv2RafFUzyUWtytXazeWpK1kz0ETlu5nlFMuWbS+wX3Nr0
PfwOgfpiPKCLIfATNKxzzvXyGbPy6ozKeQkEyi2RkSlRKiNgWgVX7EBDv9ZVj5PE
wV1JiEtMS5pJiBAmEwoXfHUxftG6NSRYJSO2u5KYaOAjhGTOCLsm5jvqO28H3v/5
g3IaoxnnoNwkxDXZcwGjNjnBMp+xLLnbAmlDj5ztFaQKJDKlK/ksCAwjTpqGnS21
PjSDcdLzuDH0smS0ziU3BbiZVqOQmrKW1jAIiq0OfbBhJQ88PGYKEuMiE7nqNoKF
vUIfNYs1Z0ejLEJqu5YyisaP+veGEZNTHILH4nV0qkUwZ7hv4P8LuBhkUOWw+PJw
rdxqZBraSpXQqtaNQ6GeQYKz+o576rxt4DzXQRfRN6LK6SR57B1FqiElv8QXyAC6
ItXMwlC2RlAXW0VXRVbJEl7PmvL6M1XKzfrxAvZb+R6wVD/CZTdIo2gDXHAQILGM
TcV3f5XIqmmvlanTKDdXOVdny46pgz7utyuVgTgkr12BwkviCNN6BlzSS9huSMhP
8uZZhwPJsiF/iq4OCtnxME/YDkphbhhcdmMY8Xos3n+rKrGvW07Mz8trcsAc3mqE
2j3mxrj1/LvFJMrDno30VsCEUvmD80GTYTu1hqIjwUFwsqR/ZNKr9N9FkZJ+F61y
cRKOZFzbFnOwVJ/NDJPZtM3MXa6SQtzm+24vlm63IteP0un1LgQzBNWF9KsDlxQl
OSs8ccmF8m8FFn8B7a6ZcHcyxBeW9neOyWCFrc/01AVh7iXXJzHkd4IJgAV362iw
X8vk37YltZ2x1ElTmvk/O9goe/N06moloqiGqff4TWrfN2KF9wvPahEOjO2H3nsp
w0bum5CkCYE13BGqMUdwRv64g6F9nDGzgsnj+bGD8nGFxpeoT0gVCRemlW2VqJQo
p15OV0eyP0O7W9rAO7lRm1bOYQbTsXY6FiIqyoeVJa6RyRzoVFAJpowLGqJTpUi6
BU29+2jjWDynx59dDR1L8Y82AMMgZr2k54eI9pXUfUcp2bd9w8CTpAglSfCgJfSy
dR5aXEMO/wnE5tKznW4q7YVOhVpASDmhbEuUGrCqlL4A18gXCqx00gqqdvWaKgEN
seusvxvU3YhOFY/0evlCgvmY2Q+wOX0rxzry3j7L/5znUkaEs6BQXsQJPH9k26WR
CwRoS4UdN+gbt3pw9GmX7oNayYtIMR/NvjWLQnUBveymf2rGLe94rW1kuxmIP508
BKMiNrsNzBa4jpGCC8alTkLJHDPY959JUM7QbRShypIXr+T07nGizBAOIGo+DmLt
SYo8/HqI2ZhBFERAxtQauOLsK9b2qeSu0kfdoG+0fAUphmq/fga7lFgccstAytcT
/p5n/EEaWsIemdem5PAfQJdlMFX5LblUzxWYMy+Ito//5SPRlP2nRXl/lNF9Jk72
2eiM6b6i8ytHK2XxUqBzgCajMPu2VBfz6+w21DyNEDvG7pWbL9zb0CyIpYa5oId5
64exJD/IpKs9fDK4WNooYwpvqwRg8589czeL5tEINiUDyX2sYi7oJw5q8X1osyRw
N31AzHRHweWKlwJqG7aKcIHlwPXgPLhb0EU5v3ty4ad77QE9Pshm4VZa3p56BA+g
I2DY5bRsPM6ViAu/+gQ/chqnS5hrjqmjQ+zmWycLNblF210FitpeGuEXU1hL5qCO
Qxs3X9PwXkynZPsy1bSlhJRQsS8qsm4wlx8yxQBoKvu025BtKpYNJ7zujc5n5NMF
YwJI7Cgefc9hZ+PoexXFgJf/R83K4OsxYZN+SdA6hLbkCPyTssVRerW6DmH+WLCl
Sys4KCgpCCHAL6YCcmTD3vmDSi4sSg3TgX10SI6I9Pqi092z5556StJwsvvPymyz
M61jqszwkXSUg6sWFcmacw9d4ON6dxFbKC3DRO6Ncp5wmpwsbRBun6rtC8f4+zLD
cgHktITc96U5my5ffrsb3GjLJpT+FNAecg7FF6ZTKfNh6FMw7G6lmoPibe/OArfU
B4n53xn5dNjzBkOQaNcndGiHYcqJ73mz2Ny+kmbMGPNfhdhh5F62pknYcMGf0YAh
NpVCS83Q0rkeO+Kx7zkh1GQMqFsYom2qSN02/MHM87n1qj5EqxbLNji4ZMSVtj6z
IoszkVmdjq6SBY8q9Kib7PEDdhn+mvwbjBN05e/TIQLmNTX+6lSmegYldC0cC5+y
Gwt9mR0NTtGs2Rqy63EwrPMqmeom0C6NntZqX6D3lz9rzfQncYpjG4dqMnPH1z6n
2O2wpktopB1CM21TC8QvJYLfTe7dUJsBLEF8isP6bvQhpeP1VBeS5KJ/1Wz0HewY
f7zJaMYG7W8wQH68Gao4VPj93DM2LFLb/cBUEkizYuT6aiVxfIL1GTPOcYoc+O+0
rGcIgSrtVz2U8i6JQPwUr6lnivhrjxUl1QoLkH8VfOo9P3rG6zHmSOJGJp8S8lcd
/NH90trXWCkubTOHOsLsPMoUwZuM+a185XUYwqeQsV64Cg7iWBBlmuyN2NORD4Zj
xsRaTWDRJ5Nne6uPtAUCx/fi/1CnKgzZt5WhClR09a2oQG7wDHEB3oIceCjH6OPV
rrZKd83EYIHZAHkYTaWaFQwaP5tbQAuIOSb9i16626cYDNnv2pg+Jt3KAQZEq/QZ
2OryqlJ6R2KuTbtK3XPG0AOX2rgeMSDxFBWAAH5aB/bpkFhjCp8PgzMA+puC1BOX
MyNvsxY4Op9J+53+qyOXv0acuW93iPFaWiOCP/QX5Bu3ueW6f5+2h1nP3fCtQJuZ
V8tZwpOolaGDyNjz54bwnxr2rthPz8oaZ/rZ3i6lyKG2yqI5zjU6th30BvFNhKWo
ievnbVgV6i18XXmRJppmLAEwKpWh2n0I1kWydQbP94+ADNakcdJU2I5O3V2AmmPH
+YzNj9e7/rDv6ZumJTgmPiov+RlS8WmwcTHVEBNt7KdubnfApwBbKPNJJM9AVNe0
GoKtjNzwGah7t+Ii3Cui4hAffgHYdf1qOToTjdSNXRUUz6fIRtMZkn/k6OWpAEgq
PvtngeycOKXkuR8lkSSAJ6tMyQaAVsnP6KD5ljkXBz1C8SjVqi6hB23H+DhAcWc9
bgw1zsTD+CaSwgIGMAWN48QeEazpl3qU62VlJN/IESSAKU3/1qLje7Ua4Crrndki
aWaG2YzIFIFA8qNSSo9u5zjc7/KtR4itA5FB4BSPx5aK3pxyslNhcVlsQGZJ3Ikh
I47k/zPwE21FxDWWfS8t7lD/yd9/F1FHwwwp2qIug+qcPi7YZkj7FeCVQKKNlb1Y
nLhygTAMu4puWgB4c+b+jXiEdvI8yHGdPWhj+HmfyuJMV8Dq8ShavPyJYbsbTvo6
IZYwWdzde788USDfW+Vv9Md9TPWExvAMxLC9AMAITyvazn7fL0hyuIgf4BAENidm
27ZQUMdjM6GP4Qb3DfCrBwu4XUYLn5TrIbw/8pQaQyW/jEL/ftWAjYj1hXIxg5+Q
IsHWJFXrhlOJQDuopqxywnQAzx4kCu42czAIdlglWXvbybpaxuKggHJvVSwuRrAT
WWzroBh8REZVLaDsklPRONHvbFoK7QG2qXTEfD+ITXi/w/QkXjG/MpsRrJ7EsR8Y
5ymp0AJWCA1YE8m97Ctc08j95x7i9PViRRt6VyiJ6UyEXi9EEZLn5YCncCFIfcld
qs0KBQGS8l6GXSIZf5/CIJSYc+U0I2T7cYyGDD6UpGpg0zHITHuuSJt9DxD1y7pF
yeoJhOP0uTOEvpnPUOPobVWPeghRQ3+BFLRSCudKxUmRgiMf2BQgZSHQf9XH+05C
LnAH0BcbEmwufzIO4nSNWP6bHtwdB6L4GEHmbJJBkx66LkZZ6an+cb/X8gQBG8BR
c5cMrJw+nWoj1LLKKLqOdEuim5GwApopUW0R9N6GIiEwmhcmxtpHxS3b2cN5VWrl
a2SpN2rKmgSumlA1Wpj+03zqcREDgkvAtzH6w6FVoXjpgcGMn49jWO+KoPPUgzUo
pH0TmcmRFU5bTqA7xpR7niAPhnEu0nt7vvh1cuVU9kwEQBkWeCiy5p+94Lp6YLxD
PN+v6ngbniOSiQQLDwFG3gbyjPKuLCJ12t/c+x5Am0usk3LmuUrSYn8g1g8rc8q3
MRsIViShQqCTdTj50W12JAdI8Zyn/f/yZYOLCxCfd4amsKZQlj8Y4iR3iZviSszV
xH4pkYmH0aLMwqq3RGWoR5bYY9lNEeLyNyVhpbzvJSfMSRYO8UILQSIQ9TDd3+q9
gZbVjSLveTAz+7bBgRv00EdB+y3U+zhX4V98+ZMkCX/MV82kCCdoopKZJIaBbnRe
d8em60TJo9Qf/RfNricRNSDZXvZrfK+mM9YCvxT/15Rn3ap8Y9HnIVdOWhdg4yfB
snDtQto/Y0iXR4Mt9l+KjU/92s1DLCnle8wXr4SqXhk4pJXoLJeVV3qvtxgM/KMr
G4IlcNd3jvg8WZNlbcIU88ypUVp5Q7nDlT1PMXIhJ1CvxZDXV+ZlPnT1FyMPzsay
ozdsyAhsz19LRa9XmoSNHKOLAMfiV0zDHXY7BDPcu3bHKzUIBbt0xi9edwz8mxad
LAEG7bJjpG2K7uHcpT5uLDX2FuFeN8ainZnDUzMiVNM67hBW4hF1ZYz6rEPfmNIv
+aArVRu475XfavN77YE/ChezFXaVo6JJLELZALPLgtKB6y+H4iw9R9AtOuyg1wd5
XkeG0nGG7WGKjXXWJllC4AYGbQi3eLCHDnxbjCLSVxMRIF3xSZeGrRlg4ys2tv5S
aB5LPKu5SYG/1byDqnZtC0awTpam0BnZjiYKJ6JhAifyA6rTUfxvRgbvURhALYA/
+vrnWkyv81kWfDx4TB6vZEGE57T2tNd6KeXOZIGytfgDxioMkpNZpZa77PJFdu3E
ZaE2wk+QQ0PXo1yOMHyzgZfr1n82C/b4fJ8k6OiwTZjD/psHQ/7XPWAb6xrLgG42
00kTZRrHqmv7c089kkfma2vTDxs4DxBMmeuE34CtSe3I5fsywLFiHXDdrMOg9hFQ
SNEATI1b4ehJ4+lFmzeKwvQPNylFsI23e/RcRqSANVHsrrE7Qnn9Ac2mgttHqQj1
/EdSCtvu4+YXmRXbb0PGbsyZJBWSRDaLOWaRg+xZ1CnnfeBrBzq7anfl4A8mEm7X
f55ZiuxgsEq/7cJ6flydh/dwWqtHlVbG1A9yipWDtnYgCFfPH6RCaHIPOH5obxX8
3xd6hRiClkj5Ubq+7MO30GxMEQe9V0lwoZgaYCXGbpM0v8C2kFpN4D8PisgJPfDu
qk4lSxv7JXKa+Y1Lj8ymm3gyf4zPiOg2R7xmm9IcTgmIigbv8jRlJMLId5DH2AuR
1KVLpBREqOjJzMAHYGftPf8Nxb7O5DQ7fblrtxapZdBSfHIwSF9973dalWqULbXp
RmTUBxP2sxkz+o+GeLb2tcNj4eo/UVVO5jp7qRggXC//JM0TCaxFXFeXdnMXwtxw
2xDNNPba/KVHpEWR4M1NTql2vfThUFZSyyYVmX5q12UslMBTxt1lYQvElzyP67Zn
86wRVe7K49/JskAgDRdLh1Zc/D8bvdxvMxS0iqz8bVTbjSd/klh9xCyqn1fNOL3L
agkig6c0SbOzT9clUTvCmO3W5MsgGFH2x8ZXpgdT5/RlRlQd6u04xM8Tf3/Ud1K/
2hMAJerh4IWQqABRWjiIyWZgUlz25zJDGvvSyPEh0wlUY8f6R2G9XdRxll6baYza
pMV9VnJpz2gGjtx81fA88tbqlNHafJmhe+jiIDIk4HX6SycyI2WGcrh6GDvY53k9
AkHdab7MUAabqpFYUHzKnfGtG922WW0MHZ2W+uaCY5FSTbbGytlfKOtOHfrhtCkn
WVE4yYXUPdjSs2XKlLMMGC1aNj7CIascyvs/tWHK36vzGr6ME793mUMm5HQho83r
f3jwO97a9HAN5owEBiFI1iQCW6jedWbpdtGl4/9JShU6yC378iM8L+bF/NhY4N8u
OzbwPxlZmyTTZL3DTxmygySJbf97KQujtwL+y68FebEqLsKXakBSWgrUnjrCmkLf
8Sz5d9rfALYyh4jPcfa425LxgG20QqSlzJU6eQYNVdDocpcL1NezOd1d0o/rp5Py
Q70xRxk94HZZF3pWKhIdbOLWEcqxMZ/L28qu20938OuVim4mwLJ7B4PCaCH/QWIt
6nlgOuYPqmK0tUrRlX6i5+yKXsQcf4doHcs3iahWjh+eC21nnCwP2Xj/0jAQY3Re
1dYPDSOUyGwfvpgdRm9T/pz5vFxJO9SxLrdxZZPUU573T0bJKdvo7x6a2kBivBVe
mHHLeWE8NC5Zgd7GwbpXObb5O3D3LDw20hU1XSKYcwvH36AE/sfGAsG0otGHBq0S
yKqaoL9/OMgQq11drA2SQeYaW87JST8TvSkyDDHms1W5Uyq56LaLU3jhwGSPil2U
TEuTap/O94RDpdIrfscSsuUJP0UVCsz2207siWDJf82bGABIYli+s2nvT0zag+it
621QmP/1a8VQ2Kuxcb3Pmb+HFR6OmByshv2Trzn6qRsnUZ3u8iknCr6HyKntS6lm
HVvIci9yvYvZW2cLrkT1/csx1XVk2bPh/KGhM79Ets841leZx4aeN7YbS48fZuz+
Gn6RA8vHyETKnwl/beteyYNTJC4moeMN6jtidubBh7nuVljOfHUoGgYPz62hgc3k
rH/k4bSwCDVuH8qQ5eX62YwZ1OWJB0J2htUYIpcguFjDFfjrwQnilrQM2rnPtta5
J61PYn24TmSoHKt537yVGVwNYEY/5ov5phtVLytlVj/Zu3PGQ2aeYgSfyOVIQftV
p4hJirR9KToaqKWEQO6H0L0VA+MT60d+sYTgSF62zcwg+FNmxPZkPt73tisINFhv
CaDV8xgVZKsXtpcpvrC/pO78mwEYiy2lOQ74NXb4hMrEOz+pIIJbzDarrOGMVzl5
SX3usJqdSeGwT/oWutLnzkrYav8VUCeR6lObjfTWYcv0UaEKINNZ78VS7/TOLAdy
eKirXeR0SAD66jpzzZ9vK3FxjGunr7uFO8VCw8uxApbv/OyoPmLgcg6f3NOp9G18
N8ntU6p+fqQvm1rJbPI0N/WESF2hsoBCwJJi7lehVVm7fW853nLDNB5IiMV4OaHK
WzoExCVcFmlssAfubevBvnH9r82c5prO0sX76xDfQdYv9zQHeMhD1BnN8gKFYDFu
6FGu/T9KQFKK7S9XIOlNwv5J3VjCmnsQ7t2jTLC+siaj7xU192tjtfrIrJqnxaIH
RkV9lY5HOnN0j7B9+GSL+RdFzI0LNmLp4Hfxy+zULJ/dnamoJpuNv/Ge7fL95RXL
hs7bu71FTV4SD9m8yRp278gCnzpn5SH/ExqYxjoigqnc38lsW2ug1fr0PgPmDZ5R
M6a6RUDBef73tbZ829LAiUjHSyQUB2jUCW2DqPPMnZcEgQa05KahileCunMft45l
FatecKKoO5hUfsh9AIsQm8NmPQMtYpPQl7HqH1y/DvOVnFX0fYyxMbbi62VSgNO6
qYpvzAsHD9bAdLjiAuPb3afiTRdrYCGbAe1ENxfxcQ2+yV1/3diH+lWD3aorUq6v
c8ta/NDcl5toyJ/JjcQAiNChZUiFgJsGTKpAjtLUXhtvAIxsZ5pMar2XBbF9xChi
DP2EvNc+IWXnGEN+w8B9N0ksgZWErz5tHe6i8prELjlj68P4vq8qJtiZvo4AjKYi
LiemPLNoph89kYIGtEv9S9qMMVTrYbCL/HpyCeTrF0jnRJm2QzxwNqu1TI3I6GZY
Bs1qo40NVOFc8JKr7XPHSOuew6GGRlFx4Hpy/lvJhtc1OsIjp6f5XcS8U3nNWliU
DdvSKTIp4dHNJyNdXsfhCk4IAd3NwFmYdbUxE1fTaipjgfHOb2HniG0K3A4hI4LQ
smF9/znVZHvoDPaofxUgB2WpqJXmzzzNFp3QCrLIWEAG/P949CX3eOcEly/ymw6L
c1l/kEcLTbeKmxrBM4ADWaQIkfvhwTFeRbFF4c/gTM3kW5WqymCiU8CXBU9Vdvjz
thGfG3VHhLLXK/PVkj61OlpfcE4ihUIJ5yom66Pr6F+jMMf1DbxZkIQeuLhuNCPV
VI6wsYa/IlkgQLgp7eAV2qQrGe5MI3N4hJVg/BmWjMdlRg/yUlr1YSlmH14RHBdd
bJTCda5ThgU/9G+KJexMVatj0pOix28L23sSd4xREpUvRRPE9cDD8BIwHNs2JckY
U3rqbEV1jUPJlKVDgpQq0+gPiXrg0Jxabsp8I70yY734wBtDYlUUY2OJDD1gpEmn
GaMDrYuJMCy4obVywOAkFdy5jRavgh5Bjq+3Ojj9Nj7zq2/RiUnpIRtnpnKfMqDX
k8SJ4SFlzOrXI/BVAgx7D0rpT0gq/UkX/HeXbt4my9hip4zhJwu1j3JdUwKOrKMY
DIcacgFGNKVeCy55lWbrc5UyM7h7wt6C4p3vLu7P2HmCfiVUVgtUh2F9OGyrwr+N
Ww2GAjGs2zYlFqpSobZOZscy3ztHojcY+b1t+59wLr5PPTvglDB/lRGfdsAKwHZT
FBm0pW5/TBJkOegTdlj8K+stVpyJGza8nAlN92sYlfMmdZtRKwLmlv58ahGebUZU
NTaxPjbH4hJ310485+k+aTudN8ZqoDyjUorV096wo7ENDWGklQUGLFKMVyg50f32
ka1AZybxPOYDV05jdY22RAJANZzeL0NLs7PCbATY1JhjMSjudYP4ev+Gu1VvQsKV
i0s8Rp0g5M2JQHywCQt8+KHRhytyYMndjsEHoEKM3c0CpPFi3jsbpdl+hWP/R8Jo
A3forLzolz8tzZoNw+M6zZo6WyPYGvNimztYmuFZQLv/VsBxJ3tX+neLq5WYW/6R
IoDWfBe/MTbMi9JAymhYlZbtBKeaspmoP0m7H1BnNKUNgSzGPU6ywuTm/hXdku0y
OQUjxCCh8I19cOHWST9wNZBtHul01PYp4tjVWVq8cSBDveLGRPyzfO56JvqjpkVM
UuYlWP5+QfWySiT0DDQVaScrCAH7e/LS53deH59gmPJCPd2p00RtaZwYh0vZ8U7N
Krqrksbx2X3/twZpQdc3IxDwBzJwL4kebvg6nf6vJFfMgEAuomkYi04YueWlyl6F
9fyV6spDTYd1yEPWYBB/oxYXJok+uLdPdQwyrXsR35nVB97b8rEMzwbdtof++YJg
4tiVS4w9CKFAiRBpSH4q9V0ryiF4sR/RUfsj43kmyqDBlMhMAWId0JzLrlzEJhv9
nvheTUfbFrd7hPm78QmuQFGUNPBgBQ/tuelOvDLKetkHuOamPYZvGYCU4uHsGNVt
tU71/geng+Hwpgdc7UZf4bYidt83w3MnL0g7PWex63HnN+Nsr7EeZiCUC10/yg6R
a3ZaRJmayYOLWQjvwZSi3T6uPFZmwAFZU/WP3l4eJMXhnlkYuj86RKMgb/U4lJvk
BKHe/zItNHgK9W8uEAS2SO4G5QDTz8fOr+Wo9bGPIPRfvtdpAwvc6MzORPtm7os8
R6/qHDd3m8N6ZBkPxGrQTlBPmeHbQrVxtKRpzme3pEb7siBQ60lnXMtPMVht0xNz
Ll8mF4ho4ns7scZifnv+eb9Y1fouPohE/2PvHIfkC8vUG4EeKbNFitglbwPG2SHg
Kd3xbAcrE3xc4bt2n80s3Jfqb/kwNTke5Vb4qeaKM4n9y5d32+6lPv6awUXylyrQ
sfYRJNw+lu/PcT5BU1qLeROYgyhKBAFLRjeb3wYNftxWx4OfBUkmrNlGE5BdA8n3
tfTthcR1D4PtllMoCgzKMnH92XHzdXSY+xCeR10gevmWtC7G5q6ml2Q6h1nSaYet
BM8jT21ysqMkHPuZ7cm4/ZUZZVG5xpMWaoOrv/+bLLoyiEf/IkiaudZBjFwFVebl
LxL+aZDRaZNCTTvSqkv+pXeTp8yQ7yFr9TYk++BMXLX78wFcJ01e8Y0HAmVNii4u
Fk8VcEoF5wRW/oTD3RwCuxzIrwRQNYdhUcEHOEA9w4TlvghUGL2mT34cjh0gxLr4
h0Y+684CjD7vmKwerkTyvToC8dMrXTKC/Gays3guTTHAOT7075GWrWUYHXcEOu7E
gmYBS06aaFV9m5s2U8I7U0qvZ4XTR89T2QRJx5YrWx5BJJqEqI3twEFWQDQDCzeO
3n4EhdpUCk5d+h8FShtO0wemJTsSVHVkA+fU3N6a7q53Pg3/Q4+O/zrIZTWy4wyg
8ZpUtSfcdzSFn8FtIQNnusB2gHoxj6TmrZuSq+LMkrAQlCumGcj+jTJjHBZPPtIN
VP/eb5DZ+zJT4m6na/Q050aIcSHK77CQop7ihXvTneMW0aJyFM5D5lZZbJag68MT
XZN6Ir9GOhRylew+QjlYZLJt1DOxdebSTy9mGwDGXNPmbhC2Vr+fAms/lwFtu//+
4DfvHiDRQIldl5ICuinCv9nzsyVeFIzu1IBzSG6hGa0FKQOObJROM9DTd5x4NkUW
dNY5t6PqPFdy9l/RP+4Irm0Bg9TX89HY9qvAVrbGRO9OoTw5Nm98+uQMWuW0usgK
sWo9PRLJ09mjRXDbcQTewxooYFnuBdNeDFV6KyooBQeQbmpbfevYEICul4gqmatj
rPpp7eAtsDc0PV8od06JeBHxJjUsc+Gq6y/cPZ3SsuKNKk1vYzaM1voVq5ikJLhQ
mqChRHNQMxW/kzZiXPDAROkkmyv9V8H9uJ/Evvbzt7j6hNJ83B3zCoZGgTF0TeDh
gcFumrucMm4eqFbzkwUhcm9qn7ouR8dXS1/LvApa7pMirxsqvBgvoI40B0iWx58K
0ZUt8gV70YcEueT1P5Pm2gXVjtG5qo9QwgNr5yvVTVwJRV/L1k5N+qF8wBlptNwU
SfBR76yuNgZxZtHihHGTO7oAU85z0Tv/pvRC3uuVvkZpWO2LTSikh02M56vQFKuf
k6GhwC1h2Ro6qjrhAdlChsU4u7YsqDdLeC0CQF0iz/JwmmPFtq14214ipSXTFeca
TjGYQGDyrQCaeCg9rLLvfvhMjmW1aCxugBnlM8dwoxmn1tBekH4rzLEh26TRQOHe
n1tVq7lxS6pwgJNs5pPBIIl/LFvdSPdvRftu5QXTLcR0uNTX2R3zRfz3xvPfrc6m
NS2fptAAsVpjf23n1ypmIfjsvhH3ZBPeWa4O4cgwwFQxN0ns+eJbb64c0f2Jf/mo
wWrce1/xsAawv6XUB1ANb7El/bj/6kw+GrlaI5Z0TcdoyzrdwdK0ugbe9m0JbmmJ
j2Z7H6VQsqVFzyIgfsE2Zrl44BNJqQwNccK6wCXqd2c+7kWdhvGtFVGQimZPRcMc
tGL3NQg0Eb19wkXvH3u5Hs04COAP9Ek56API+hlKFIqwEe6ZrOs34/MEnyzV5ugd
pxaoXhJj9pKQFYF/szRkvlU1OeBxk6uILTDJEQvSm6GkFLG1uS+NmDw+TnJJRxc7
IgE18USxbRBRcQaaqPg5R8v6HIHuucsCxkGTBAGERPjsbYbQ2C1CRaSb6zZrXrqS
+dv47F1gatOwOCX3J51/IhmuNBg6kFXUx+SN8FJz7g7s5Va/ljM9mZLlbOPxcCaU
nKHQ1tBbIcBAL6Znr+I59OBdojWgKD6ii9KiqHgvCLRsh0sXLglYXxFJl6BHwDhL
hIn7pUmq0bbvEII0Jyi7goDAfjZKCM8FeRkFKoqfjyZvDDvy2uPv1T1dBxIhui7s
rDCsVnB1hSWarLLZYo5YiS7uZMyFvRoiVZstAhHNR2/sChD+9YJJ9aJNAWTkmIry
gQ1bg2IhhnXF8YIvDvU1YwTwZ1CpuGjRvrjghQDQjgB4kwdrRLBB7vzw79WVu1Q5
pc8jM0QL1tvkp9BAud8yNzRyw/yz7c6pyOxLFe+zFgpwdwZdVDF43F/YBrGQC/gi
UduU56t6T7xKpL4hdHfL7XBLo8gJ0+N6osSvx68DELLFYDkd8+Qa1UhMuJXs20T4
KeFF8CdtxFaDCzGxq3avZ1uR8uEN04rT1Jmz25jYXg2/X/FXfPavwnEBFJU+62rB
qUzJCOirjIOzXr4mR2CFskLXPNIRrr1KLjxfGf6Hei/upwwL6QcU5M4iqJ4L+Co5
X56E2VVsXpk2+JJXvHIdImiKdbVb+mXYRF+FezGuzemHn4v9ajx7/dJ23XlZvgqJ
O+AD72WVClxmZuc/8rNK9op26YkOnPVNdhG3pAVpiZZ1I3rLkJoYKMzsTjW24lVz
HzkN0HTdUmwdcheOmsZsXoZWv2vjpnR7UOWd4H3f6evAv/EsmWLE6MkevHOdd+EE
lAwUED7QZddedUJ0jAcst4UdNbA/Ym81N2jgFcNQtEhIrNW/HiGaH43P9DPZcbE0
O57+Vq0sZ9W3wDVBNy0gz9+soihHz91NMYI81MBIVrbmefr0KrHxwUmYUpdxqNYT
ieU0C6kzN+3OqykBn6Q1i8lzLXydMBZO493F58sHsX3GZ8atbyeYudQUftUwtqaK
DcGLHfAGUm9EjIbi+o9rhqL+im8anqEZrf8EyQlRYD3d0k40aqB8600CQpoyzl0W
X5SWpE4HrkftNGVFd39S0k4vWpRH7p1Q8yvlQ2P6pRXihZuXQV5U25o21YcAJfQ3
PdCp3tAvY+8gGNdQ8f3ULw90ehW3Qd/N9w0AY52nv+MoKDtxvH1BcLyeHhwlOBWE
q213KzsLc/rjnNMueo2X7EWd3Os8HFezwJoWvGdn2fmzLpgGNx+ug8C0mXV94s3z
g1/fTXhG0p5ytyxAAKBTbE1hnXHEhiJ8oeYkjsAD1fw/fkK4wxpMQ6nJW0VD4nLF
6g7oMNHW/Mwby4nR+055JTOYcIhNrLYeXmd+wm7rbHkC3dMvbRjPmKjE6ySt79q6
g9dGOAU2gGjkndrdj3s/qCQqPT5+liTUO0/c4G8ZKRHbU5NSYUcTSm1uW5zLBRZP
YmOMFIN8vCxC7nzErE0X+UxC2hW/wsZkoQDFxwOtNU9JYFyeLRZ1fSbRBeRdRywW
NHTpY00yr7zUsw40nej5Yw0mGVxyBwI7ovIvZaXrUodLxQAXOB3sK/UCZehD5gY1
cBssUBdMEmbaf1YU1TCyfrQ5n5iw1uLN4TV6z8jGw1lIlr8/WmAtEx/PMgNqn3ND
B43x6rgSu/M6LfMRsMdrYLpy/sU2Oz5JoZyjN/DM2TcVDRiRbfUUfkZLUakXzXg5
QiIUbMuWwWGgbfUMS1WzhaFChEQYjHI+ask/pr9vrgecujO7SoNyIts/eOsh/hYp
sLP66y3KH8F2IWnD95PN2Bx067vJiKPSM0aFfjeCQknZEF4Wh8qEGfoAApOEs4CL
LupodjgLAr3TTZEOxcpcrueIXg4+N16HyyTFJlQg+DqXozhpp2/NdZBUG43jvDVz
wHzP9xQr6dNfUn8BbVU0p/usUSLouPsZaUGyX+F51ulk1scpJOt3jdfN/919xXig
lI0ZAdji3ukB/cn/GLL+D9BI050v088pJCXw2pEhZURFYsedSWsNJZgc3Xmz+kaT
1fauf2r+Wpi2vEKKsKm1wQmoCHp9F+GqTYiuUNm3Da+xN6hORWpOqdeGb5qRdFFC
MEux08lKNO/FNdfu5JOCl28GudCiVJYGYweHH9I5PjpM4/uyIkjd9DC07CevACKE
ZybfPZh8tp4MWnix5oByHJokl9EVxTWplxldtbds0CBqSGxQ4w2iMPcchpGaOg35
DKK0oPJnhAtxWFyWUDAezUL5JXXURaxKyCUuD8QHNwg99he048EY3sH3pmnFFxXE
T25YUQ8BU6JudVZd3yHeDbDq46t/ZqG8IBGEy6xLYHTTLzjE/c5yj8XSiEVXvOWF
5azMFYbJGR6JbLZuRO6mUyGkCX2yy8I7PxrX6uQzWCQJ3rwFRj4CLUvomDOD5E05
q9T36k2FEDzy5bYKuHHkn9F6gRsbIV6/kT42ocqO5h/0GAXHb+ds12ahGCofOUkI
xKOrWKrMNvPjfyqmrsurnX4YsU/H/LX58Hig2nJw4elMdmoJZA6K2ULy7mRALSsI
jGzvKm9pIjf3Jfdua2lPgtKwcJxVVjirXEc5yimuQsCNp7SsggnMk0twXqO+3O3H
UOUn2j/oHgNOaaSyJTBLvKLvs986o1UjV//Ww6R5O6Jtt29v2EPj3nvUJbHn/Le+
UvL+2QYsqoABPz0jDxaSXflwtKdmIP907iKeyvsG0zWnV2ad8z0k2vy7D6I/wJ05
lWTUEtEjrOv1fGjjo4Z/9vF1yUthVHpg++fnz5frPpniLoe6bZJG4K2kctJFB6Bo
B3Ri8HAOTHR4x3eO3BFDntO9YtBxqjgbZ5vBj8croCFihG/uKzJqO30WLUXALPos
UmsoqIGMSXgofQ3jDpwNr8bZccQDXZl9rUsjSHl5ix7OWUp8SesGtASlR8fAEDZY
3DBp5gDJ8hgwDYapcBV1t56StzlCIMDVrpixJdaZ+FRA0OsUojxrt6sovFpyNiEy
p2n4LIdtbfz9QhMg4sdVa/+iOPsBan33SFNsmou6t+UuuuDSMC5inQ175Li7CBTw
e4AAa37UoWwH2lkQA2C3ppYi+jHl5Sy1b8j02tEFw/C7O7lGStLzn3GyRnKpASgs
tFKWpfoErgkVVo5ty78sIRfzDyXcKfCLJMvEwabNtn3NshzoAFbgg89J9z4qc1FC
uw9fFSkMVc8q0g8xwzuzcsjcFcPRz90SNMJ9U6eDuh0Fwgndb/5t6K+k/bJgC1s4
F3Awfs40siVmi9x6DFq7OibYKzaFi3phrIv5cdjXG2pOHVs7ZtF3d3YfALj5ehxJ
3rH+ct2Ut2/SjApvXr7Qi+tqV9rEgtaclHoxCUoK8hxCHGU2eywee9aSxfpcTwJn
A9C9j/ldIF+G5vNQr9zEZBoYUsutm7HD/JSLbVeyH+VpWEgfZ3J0+EJCmHvcAIts
G47OIPU/uk/KoijYCq4YbWysUV03/e+s8hK4zLqNKTvE6Eovk/MhPB8y7Wvx9MiL
z3NMf3wg4fJjVp5HhBztnxJ9H0EXUjcVP7vg9D8JAQ02q/Z0dMv0lCNdmerbbp64
jHIykBgCSBwK++8kJgRoTwNRolBKcUa7NwIw/v17qT7QBn3/4SMez36lA+jYGVnB
VC6i1mOsl59g9Nw3jD7dsa/Yry4AjBXjP/l5CwosCBj143Hd0m+YL6tm5XbJkHJT
nR1XZIMLL+b/vQmgLsK0Els5ywYtICoQbvsmMFZ2/HYCCZ6f6cZYEqs6iMNnYcLY
K1CbGHOgWgRagNA3/4RAZDMIwP9on1vzn4TB51p4pCGO8SeI1+hUbBiDno9rHXBY
96zmhMwiBSP21ta/W49rZ0IWeiWpcwFfkbewEDUE1Waxi8Hf/iNr5WjmqTdCct4r
deLmP3+vFQMHL7FwznFkJ30K+dmAl6xUJnIFrlhdA2wPOIzPxiUW3LrfrxGFrMKq
I3E62lhdYXcXKdQJoLBpSK3cCwH/2ECJtbRyzTNMTkQlRM7H67Y0X4xEqXBzgTLp
3/fFTc/vpqmgmh3vwONQ2r1ioiX4KXoM9UcAsHwW4OTBJvQmvnCVhWJKKu0AYDit
tVpAb4KDKkzX4xeEzJEItP58Ao6L8tTj+pFCWrJb++fnDhHgC96gHCQ1vNAAw2w5
2QS9GzdH/0LMF+ly+EFCjz/3urzfOLCZrDqmMjCKL1ue2KDpdT8HR6m2or7P58Ln
PhiXXjEzNJITa5wFQdrRfBSKiHmkWoFozYNw/JajnxrAp5bvfo1SKYf4lfAntg2A
e42OfB/Y32C4Yb8BYw/jtk+cAwdVg/TO02l6QWpkoSSVBtUmb8pbOSseJ2pS1rP4
hJQMKjhekShwV6QofcJMA/Zk5RXOdPwqZhUdIY4TzaoNeMzAnA2Ij3xLsyCVfaex
B5qXMapGQECLyTSZwsqTzixmRbA/YxTn9V7vgJBXM95RzeTNs2YRfm4e+Ca1w+1z
DR6G/wjPn9eCxPEiWwSKaEpbIuEOgyvZR7otuBLBU7BrzDgD2dLWeFC66E5aP75K
dHm6VyO687ltZYYQgkhEClRnuu4EBzjQnGybabXVKFb46rFaqs45ETAABzRvRGCj
GhOso8N7JPTzR7inAhAQSQ0uhWA0fRP6ZBZcwqcF4yv2SEz0mBxxQEd1Koi9Qjt3
sXwjHuyE53qc+kCk4KUR+0Nz0KPyhKuxtWAt+XJQl4JQU/xhuYoGJSqRyopKq+am
5KY70St7oK5dKJWEUJ4vBCBQQc58D6I59cirLu7WTmqcb1/73uRRSHrSmqnyDd57
DGK/p6mgye6qteUab584lBmjctvDIM/W0RhkCzLP+0pJ5GbGU2crsnxZUgB0WQIi
PWMeiDNqW+KcY0DmtwZm74F8Z5aSCYVyogbI89ioBvVdTTtiQJmAj1Bk8K656G5M
4gv14C+IPMrjcFCKaUrmyNJnC0PEcaI6GBDwc5R6ccEhxhw+OjPxcC2pSMS8U9ig
JTy3qs0zD6Cto1efrmpq+BaByV34mk2zVl65J9GaUVpB6ZijD+2pWmqgCcApoi3L
vJsHM/3knq3odc60FlVGD/fQ4UmrTvY8IdV+PW5T77mKRtVuwWolP6fvEgqNrG7m
1eVD9TGaweAYJPItN+SKpUV89jdx1AkK8QSS8ttRrNcpAhqZVUS3T4YLRS95rNjZ
V+brkPBbdIu7Mq/u10U2C39Z57eZ40SGEGc/CgKizDsir8uv7VOd2tZ6c68D17SR
z5lrOMpZEgS0sQmQ1RA4dPY9MMw8HHrfjD00DXsscJwqlxuIeYokAFaSserzrus6
nMAo2CSKH5E2FUBRnlh+yL+KO1fqGFNX2Nz++N4OogKPPQtibVAk29OzVpxb/ugt
5REzy7mKrADbU9TAzcYwY5BxRNRj8wmTGGxcHyaS9ACFCgEgdbnbfVCOSj5puhFa
SBUDsWT/ky76U6uJr8JyQsSVFlymPFIkBdZYEOa0Wj1GsUc3a/V2Fcqx4r43X5Ol
RuZUJh5MHcBZ4+rA7vl1RmV61OtIkC+m1AL4DsaN7GM+BMHodCHUPryPPu3Q2NIp
PKqX8ebADAkjEZb16tcafbZTykffeYgjK4I0yqEaQVvZzK6XB9l7tGSLWwscXEPg
ZNh6bslJVT9UIsxNs4gJHGKCa4bVMY0e/0WTBGugRuHVP8enSQXPOzIocM7Luqh0
9a7dF6Obp7SpFugKoMiKeWcPY0v+LWerV0vBTqN6IMn+iYokM0auinS5vn/rGNl5
ULaTDPs8rZsVPIs6+AJJkS1WxQlAq7y6e+wxQ41cWRrtz2j+bYIo4dnLk5PYk5dG
lQpzJ8si1NYS8RZ1fKx3BDWdjgOVE8eneEz9KmbymxwzHj+uFR8+lYOJIsNjYJKw
ytq4W+xaR+S4bFI1FE12A2uIDE4ASWryZPi0KoPlYeTJxrQAtXCfNeFRRoG2MfhK
TgLVa+aI5vo1xfZ0MNqsnZu/AUvkWpgSa/CrX3nUB8mHJl/a/Z/NQxlPrkmlLtqG
43fHBv+qvkd7j/6MRI9F4OYeqaNldfsu385bJW/irYssuZT3rZdd5pkgl02nnmG/
zC9wUODfNnKxctLEsl/TKlsb4l+5PWNcdHQdrKbisDNgtbo+1mUcMJEfM0ZIikcy
BaP4Dol2/PQn7srraUPYUeR4psoySdBOHDfeGxop71gV9Euwvzd7IDHhJLMI3Ieb
3uDQ5VGGGSlsEqVqyVt7Y6tX01JzWzo+VkFHB/o6mNdHuqNqXPk0e742aAD9TUcR
7iUU0oCCJFqsyKSVP0Np0w3Gs5yyb4bhK3oWBnGI/0pFV9VIiZ4lhot24wDPk/C2
8dO2nlxfBYYSa9k1xAlkvgwJ8my3VK1LBfDKMSXS6rFkozboW7LN0T3z+cVW+uyp
u25QpmF5NsZHrU+LTOJMh2jlw4vfbK2Bp1YeF+ylZ+yT/5zg7rWL1oEI1VluWwN3
mT5CwSlEJDrNj3ZNUu8Hs+J6Sgmgtff+lJK//uJAQZrbMJkWlP+73P/sOlSRcXat
OZ0zSq5PGpIxUDoTLJBQFKJKbvxsxlg/FtdxgdqDhzxPP7A4EFpoPeRnd0wdQZ+z
+09aZqqs8W+zsAVy9CidqcRgj4OVO6WbCBaU7F8lRh+XhqPiuc7RtYu5EWC7TSgT
D53OWHO0P9MLgDnD2cz9qABl869NYy3CmaSLQY8HO+wHXOIZ47Aepk2v2BkQUB+O
g2lKXumeJ+vZfBUPK4UJ1lml/XJiCcH+bE4TvrcEN3uyHPHUGPpe+IdYOVqBWaCD
u7PGk+GckG45ogIYrHU4dZRCRFV0hL4WlDD0yR/ABFEbBUMNJeqOg5X0WHsQElok
dO6/14kpKW/SHKCWeKv/exoOZ4xI3YhddAoaOadeh83csEw5hRucbewXFaYnr59j
3otiYgHvU1RT5IVktBMNO1lpufjgpxxOgFbD3rmFOWzz5idYTnCEYWe9JzVxGdIf
V72I+0AoVubsh7hyGe8xkYF5v67NoK7qZ85sQFX4P0K3RnjiwRsND63mjdnDCZa+
bbfF8HKmQCsbixFqu2Y/6rKsOcVTBvAAZ9ETOzBv6ddIgP6GBLmYW6YdpI57SNFs
fKQ97UT1IpvPG+iwM4SHWar97fG5AH653yfrE7HPC0S0rY0qUq45i0QXvUfYPOic
MJbCYGxdZNIrSG/5M86BuIPk/izUsWil045UatXe8yDOSDzDcox30svZ7Sk1TRsk
GYfjJnLnnZVrYVeAZp2JWUKeVZrrjfreR0bWmPFtKeKoDBOqzN9/3VIb80VAuIAB
3gs3rbE75wE1Oy6zsCDNt3cjyQPcifQNn0ukc9qW1MLv/Nm8SuId8F59xQtNQHkj
Nlk796wWxBVkJyLKsbgqDkGSkyD2TIlPXAdCRSQ/G+knU5k+vlHMU0qQer95A78d
VEILsuPycr+l5wHfu2QrnuVVxShiOmkdFD65p8KUzhNk2tqwqHjor6oQ15QV3dao
+jUo3IjdyNqTUrYnISae5FrjRutCa9ZqXvzh0pILIJu50xsxXWVBZehLP8LA60dl
UMF3kkdrIo+SFDMfouCHxCHQoEN4H2JYIjyx021xC6LgDICA8p15d+dL8Uc6CBcV
oIG3lZ6IE7bLGGqgAZnnur9AvWaQfVsuUVgTXmlVxoOsckP864+p04Js/iRTvs2w
xJ3BetaOImaBhBQReAi3kqfjt6bBsA9WqUG8xJaUh9cP0xfkaagg10JFUzZ7p/4k
1ROtbCW5/29xKtcG5bowo7UJvyc+gIsevvYSTnFCrqpHrbNArMEvUBoqFLLKEK5J
zlP2rDKSYctHhPajz7Vzf+uBI9B0EBYWxUTU0sKLyCVCKRJPwpwrlavE1/o+1BZq
dd0+86OZY6s/XxogUNWUGl/rmY1JIPThsTae7d3/hDrSInoSfvLqsC65e3DlhoRQ
9i9vucntMzKhARDDPYfLkpfIlMjmQUEFFZotIYgH0EstpF7VO12thCaZvsQl03WH
Ahq07eVJWhvX/Nq/y0ErK7W9xNASZ63EHrSBZP6DQIQiEop4quLx+hB6ftphJey0
8aywf1v8Za38oFIM8LFtKt+uvKIgYPOEMERBEufB8htyK3SarVPXFRAHmie910+2
aIkmQjtmScRgzYYcXf0nKCyt0B3QxSSS56AK5p+uH04f1KElOpLevXFWVGja5cz8
VK4c6goH2DKkjGLtmHQkb1h49nULwYmpDGC2yLvy+WR59kFUjJJ5hWHyLB8YYTOH
vW0GiNOsO5fR2lvzE8qvrBhf9HlRYgyjcNjKXnddXQXQK4Wj+l+P/gXxC96zGVix
OS6GEd2zJMkcUfizwv+8MV/Q3yx79UxJFKI9vfZl8dUvP6ABAp25IQ/amZ9/2vtd
7RNkhPMaSL6BWnsge4pyLn5kZRGK863ghNvYC75VodaMH1x7onilJ4kwzn+fbrC/
vDFEkpuiAoNkcZeAh07gDvEsijqfIkoICOaFDZPEmfCQGW/Vr/KfV4UtOvvYXhx1
uR5dBjVCkXO1Jt+FbD/4EizgXJrPSW+So1YL5VBtbKXjey0XaOLzy4wYKIpYhyGT
eeKamBZpRkM3W3JjIgAWD7HUjqxlwU5V5hUC0gjmbTooinRnVtpVc2m1GMMKbwcW
19p/yaSB7/oIpHjh1zNjzc5cRbNCQ1rRnghuUNlycFdjCu4v/H6Cxk1e4h5WtEpp
+QDlrWxPZIBD0rji+mQjjYKs6UGTUjWWQf0F9oZcyZkBcMLo1i2WYVhh8c1QrexC
63D5NoregcdHIOO85dn9mKakgQXCA15DRjoIj8L+mXRHlExMdTZBo4Rs9UptirsG
u8Xq4DgTirOF41tLJuYcItgpi8F8AWDIXawsfNHjJ0mJf/QVlOcLELaPqowByszQ
Qwx4cu/x+JjC/VcMC6ScU94yoy3VT4zA/jYXvjqhE2BHAIxaNxfLD6b5dPazYaYg
UBoDi/6PKSVJsQvVxkYZPOgbxyaOI1O4/dPYzzu1szB/0gnIGltHOaYFsKUdlDwx
ABFVO73Uchkn0Rh4SYguS+k4qFYtJf33L/PdxczBrExbzMMTUdPMT0U8KkICBAJx
hSw3v03FhAu85888kc+g+lOxmUijvXC4SQSJh32LWQHX8XGaZNzVbmTjrd4UHa8X
u16kz8bBKJ4I7vavAShllVppx98KpjJSlqh8+IwwICNOC57eYRhNkti3vcV85tyP
LWZ5mCiCOw3p0B+lRbL7BFjP4+RUUOybmA48fBPUx9zMrVhdH5q95COGUNcV71RN
eGbl41f7w11NWBggtC0nYkFW+U6eiTUoujEvnqFNF8HU3wlqBwdLHZENz7A2kOXh
XV02dvMtKq0yjVBJbv9bVV6yIENJ+FAQk5I0LhMBP07CD3/yhJ4TPsAK3f3UTDbm
mUio/I0OV6agehwuBaJ7gkv0PIsr8qAGM2aXyui88EeCKkQx+LketOuh8hXjsoWe
a5Q1TSLzIV9IXj6q+S/P3FvhBfq7RnDkr0ou/GtsV0U676O0WyYZjPZQmt1Ue/hH
PSMnqgs16G7PS2vFlGCWMjKite8CqIdnqgi43lhF8YetkElK2td9Lh4TCmZaRnK9
qS3zY6RTNv71ArfiSmsmjowBEPYWbtLWQfca+E9JIHs27La95VlYqO/9Qx82EUVY
5eLgy2a1pwDgrF9tGuah/W1lcmtIOxJXP9vWtuFhJu0rfQNV9Z1ymK1yoxLLPR9G
CcsaZwpsRRa+k9kbiokc8PyhTmifYPLtRcvOQI2j+PPWvpfAIbGzgrvgpbKOso6x
IHbxoqmTANIHrcTDp3vij0/Y7ygOkRTHHi5hqf+3NIMYXm6OQjHXZtXu3F7q8cRq
3lE+5ZnBb+lC+tD62rVBC5cGDyZ3UfcRNnXwyNwfh40ZYUpwNFWHhHXbDjTC4hzB
BNIP2Aoqe1MAC3jp2vaCeiIvvzQHWsXUxueLMwykNkXAyDPz5q43vF5iwjxbdB0w
eJlwTd5ouyXZfj7pI5IB1lKyjtMQyi0YZzDT2QkzrOQhZQFsqRYipZbAgw4tpvv8
v/i4VJwJKo7n2YQcOLaaKzzPy2qOE5+wjJzVbXrFyt+NY1d3uIIr7xDM66zBQLkt
YGIO1pEnmLi2OMPJrRWEL68tiSrSwVj8oI31vQwfL8OD2Ecpuz6+oFz7yfEKlFJL
buhwBD48lO2jvTnYQ8r2IEk5HpZl2bDsZRY+qN7+rF4zBFfDXTmeUgtBeh02a627
qQntWofBwrJWAsLHfpy5HQNHbikSYn5uAIxWVPoDbBtSbs5JVdSc3xcgtAEZI1VC
mcnSx/hICr+JW/Hwl4Fv8UCW0i/dIlMvH5PXQ8eZ3cT3ZUA6t3s5ekPxCuzSGu8S
RSOjTQEJMnRgQGePtnZvPC+Ml7i5kH67z5N3O6N80Vn/QK1CY9B2cX5E2ZPH3tRN
SeyhNjBIDFcBNzAWrlNrM/LtTGjvchcC//+cXSkCdN9mfZgrPExJgfjXq7ogsWzB
vGHC5sNLc7ofWrQhC4bDgUpaFJj4KQgmA5siRKpaP8m73ilFUyZIWXy0b/YUDMZE
WhekAv0Rz9hwhzwApgbFWewHP7D9xMwtmRCrZ0zdS/gznYzxMm6S4jPkM1pLHoVv
RX9Y3hmJXtdqr3Jr4BQnDkF0EwDZzzFCXP+GIVMNbGpjUTaF0ZH6dPxO4evbtKE0
F7FYpGNBdf87NGP93QBjeTP5dy4hzgL9Sufpa7/JKlKjtKkPdD7+uOJV4Y1uBY/Q
y1LLRAKgQ4PpKkkDZLf5sNGnwiqSHiB0L3tmq2qVR529gz4AYjueSTXkX/5tyXKb
mcF7sqjel4/PEmYqnXbk7Wwg/oKx0O+f7F8i4FfrvPiJDFvl5rBLYvxo4mRfsgee
SylICd0VqAGNBpDPTfgijRRkcbW8lEWoLN08UIBSkPKuaGgi1Vq3yqy0+keoqzHD
6tsy6B6NU/SVNxsHOy5+U7HIDwaGlZspk+FUH8RyBwiSsA222nFrdSNcJR8XhMqn
nUOyC0w87fyR1cswrscBjACs5FKP26NXNynicv3JBeHYV9lT4l0gohm6mr8js/rK
0/GJ+efPF3aByiB3kAeUWFZtQxapA1mdqaSJEccxpTUqptIt0NwS0b4g3PDy5/AA
y5K7Fp/8ykMGnt5zDSHboKLEzEq0JYRoIuS4UmOzxTm4lVhwYFcrEne4yjijFfth
DRshofBXGwKwaDjMJYVV2OY/lipscVKQvj0FjuK4r/SnP5DQKu19+KngOc4D2bAS
U6PCHXBuZGShw/khMNSH7O2NZcQtqI4eAvh0Dv0wNLJtzwkXPMG0P+uutFufqGQc
iqj+0K77uNdcbn14ZNTCCLFqXna1/ukQpZ17Z1pAXhrqdfNoQbHbB3GgAKx1pPLt
DfXXCI4F9ZtfJWlQZXoHr5sBOSWLbCK7AlbO9raZkvkMr15EWPr+4ZM3znPGXKIO
IV63RhZnUnjrOB48uCSzautA5LeayxF5589LUm8BrbYNJOZrGoWCNrtqdq5nyk02
iIzSPljmgEE4RMplpqXpv8OAVnn8Zrppi+jqCP3M3cW/gjqjsgi4edBsWU4K94AN
jdDx+yoP/xCvN5YpXHcpNoI+GOpVNpfjeFbxHVZO6o6QBOAYdROTo6RhbAetfCoP
GQIRpO2OZo68oxN/GC6nXmKaoC9B/tXXJAkZHyLxiUkc3wmWJ1EP0HY5iOgTtv9c
uud0Nt9l9RFCUOZVMoJKMZpPMzP1JTdoA165iBqIUzShfn7p/aZ0P1E2X7WuzqeX
oR+nR6m3E/RxrxP9p8u1xPxJVjiq7Wpjn8EzyLDBIeRaMk34fafNl66wHkhD00sF
3ZA3wYpOkUCnoweSoVMShBhVraHZkEYbJxd9tUBjfs153umDbbJlAUD+4u1dPC7W
0OsG1H6tREIr3amMqZdKEhPdgMal2NufSdn4mhW3T04f1RKZ3AT5ZDNz5zj1ehD9
mXnb60PA4bxlH9FJvv3jpRdv7iQbMtAZDJACjPKGqumjTWBXDwpcW1HNpOJJ302i
dSn2wNnHBN0s+1yGVIiDkZPGspYugvNqjCgcxji5AyiVG5d9TfXqwrbE1RtO9Ieg
fHiwt+p6OzcS6vQ+kplz/mXvwIFUiC5uUf0CpMP3wQ0TW2iXrK5JJInNlOLz4iHC
ayx/Pkzc+w/67z8wFS/bRiSCY47igUmj+mEftzn6WlwAJ0FDnzl8rksm1a4s2qUQ
usqGPyNo0YWS2edg7o86vF7vm75o/YAcZxcFpmiyVBo+tMnCY4NdJz+ImA5i1mcm
i7vcG4NlZkH+8Ucq8vEPY0dGFz+7gTJeH9s8qIYVAT6UnTmy80LEOoYcQPycw/FD
6GLZ2z+tHngyNrfKo8ZLaJPItVgn3nVw1TZrWbLARfmPYY+H7W48/A5bGkMM1sZq
Ilzw8El0qkW9b73fg6weXCmGzDqNHc/Cv+biLMmaXbqfR5p6DGNMx3CgyFjZahq1
SdubrQ2MpOHCSnixRNmkRazY9+zH/yTA3TDh9B8digP/5kchM1IEDPR8zDCSqdR7
bBP9q2aTZMVKEk8eH+zCQerEpGqSQE+f6pNwIJfQZv+VCAAK9XLerIx8J/SbKxaw
bf1Z/d1OI2IjUtmrdA2pYcKMFsgrr64tyv5tbDRtuwhDrk1hL6vvzw3o388W/3Fy
Ex2N09PaWBU468t6NDZA7YtXVxcaRGoordLYzF/jhY0m0WRhtnRd3wLSp9vm2s+K
iGFisCPZu8435/o2aIHA91+R9ZBkG+Wf+quOyRVfzCFKe4q8s+PD0aqv7oCRt5P5
LnliMEeKXhnN9mvap1mpdhFp92FFDtMf+/ckCuACLY5ZBJi1cl4FT4riBCqOOi0N
uFdr+XdVqA4N2juc59ngnD4VvLtxCXWj4OXpUzFW4DgihG3gY8PrCizDK5ZpqEsH
xrXmgJAJ4f9jSlqs6YeJA1e73agdVTdJfNwd5tOpPPHncrnNlMfjrd6z0ZTx/bXg
nsQGm79KkXoHWDmmGQ3A6H/q1qvuQqcTuck1TkB3GQ6vWZ+A7MLZhv14K74dKt4H
APNrL71ZxOy763aus6wKPOmqlxOa5qEwT/dGT6m1c3u0W/z3EpDdiilk4vCjPTMG
PF1O7VWtoqdLeMT58fCGdV/kGLsTKQfyTqBvNBFoUhnTiceq77lqyfv+fOa1F56R
YHOOgb5NYb1AGI2EvTnj0hlePmT7DE4l9ycu6jwsUQd5bop8FfdRnJJa3l7W1biG
Ospz2hjM+ptsfhFMSjw7h5YQDVaxpzaulEroNM2ZDU+DKgXDaD3LGoXqAMKDGYWY
lQVM7b9YPlXFghtzN2J4+6uvuVFcZ9pq8Y1/qlrr5VcELkP3jdbJ2IWh/Szk+DCI
zaUnOHJVxcvesZF8DXbLBFtvMN2O/5ABYnMKikBDYVoO7yysv+LURDfBA9XmvD6s
2i5oHh16zDAY9OVB0OmyqroxN7NV3mF6jlN+9vFmePZBbaLqIiF+b1CU6mFPGVn7
E0sbeB5q7zp2mjXYa2ClJhRkkkkXGM/eHxE6BAV3eSiPWupR9+OnQ5Sp6wyBjwoe
t97a54OEflvDVF/yAHgL4553qa7PLn+1Erq3qFpO88l0aPJazTBtcC1Uep5E+icd
amyv2xaZAm711ydXW+2uubYpgIX6r/Naq6fsMG/cpCf4dCvhlw3o4fI9ROzfiE/B
bsKEhXBVGuOqUX+GeZ0/7eMgC03m9SUHZI2q5xBS1tnFBZb58A7lsWh+HBU/Ecxw
CGmpJw8CJHuET5QEzGQt3VlzahBgvAbnJHloqYWq8fiK/mHWSNRPd/3FeeSkZ9yk
fGWoIptemjDHJeZloWDG1sSgxplDvfe5ZbjikUs4kvhNuh9y0HxOmgLpBKtgHz0s
bz2iZ7yP1qqAcy+c9gdRNUyEeOtJyEt9qCga/u7IuaUTZQml68jFAllLdxrUY022
1B/hqwxkDuFNzki8bOncGHz/ResZ+RmKloTq40XwCmo+htKIfk6M0Jub8YHfaXYU
zLsp+pziYlroE4vissTnEy9YLOAxWD2HKCldpMJKoturznmLAVRfaLd4NbMOgLIf
5AEU0phsU8YX3FV3K9BzuK0HyExmnU4pkCSA8Guf2L4gW0DpVKtOkvtK8MJ5Qjju
2JCVpSMiGZYa3s2ro4sJp4GNe9+T98zlseg1gjbe3nO5jykzjR4AD2Pu80TM68rc
RwmNhjDoqaD7EiE75B5Urcntf963vSi0FvJVHYtJ6bdM4j0mUAq6wZHVfksmaN+Y
9q+MLCsTFKUt+Oj1QPBbXXzKuNkI4hfdmBcruOtXxHG7Aon2QclzWqgnnqhDgPLT
ps+zMLO3in4RiiHffHynbg+a40QgRH/ZmHgMtP5NUcBAosInXHfwVS0N1pTMY/qy
crnT0ZkX9AvoyD3qgTfeNGy/HHTFoDWuoj3GBOM7PL5LexRAJ8Kem21T7zS2QJnf
39cAEgbfcvuZrRLvcfwpQ56NK54L9xPBoFb2OZmpzwDhXwFK9Jhq34HNQW5crZ3S
qt/McrBHhoxLx6wkCaPXsu+SCoVatfXpTQ1f/t1KFpY5VxIT9ZwSc3eXWHvOIi/o
K1Amu6Whv7qIwvnWeLN2Wras258593LOxIYlMwVJOo+PMx30vrDrpUxvEydt40eX
cMTfb6VyMab+EqPaRRQPQR/GitM1uQIJ8wPdKonewKpIjEHUB73VDlKZcLp7YO6q
r5IKjuzBGl81CAy6oUzIg9Zy1pmllKE/qYcCQMgduvl9/FKG13nOHmgDaEPomrlH
3AtY1Ami++3SafNhyqzLEZxXSQYQq8RdPC1qLPj+RQjcUGlCtXMwdvmVcboW/04S
0Nxq2WWZ8wJYOPhCwdfR+m3cj2WISn8Ele2M+zX1YnQsCrih4gntCRHd6IbVNc6e
IlsK0oH4ogVLelT5U5CJFqjgMRwDAvpP+grFFj6/GojSqvQ56gl9qiQRBscVTHMc
xWw2eONdPJI5ocTveNwD6E3QjTa9sXPS7IgorJrsXUTh2Q3kx20xrGszuKb1wEe0
M+Mf1mLDdEs0u5+Wvt3zOOA55NOonLyKmBxhK5qFAA+twbBlAx5zaidS0jlXG7fc
cge87aD5gW5FYffQqB/SLiGMCYk78Hr+qrczfR7WL+mr7IvjAYgnDZ5st4wSVEuu
0tUpCPRYWOD5NDbNizPvhCPNuQuto5WCyxc1iC0Lq9Z2y1apgIzNu3W1h+/VHsuK
LEAsyPnxo/0Q6CXmOSkrkGCrER3HArQkpUCcHImSGNmSBNTbRMYN+G/9Z7WDnzqb
BmYoHFu/hPY4S05s+97A2VslvSPWx82ttAChZZY17A+kb54GwyzubDWypzVVPh1M
/7AOgBjVViYa4fgTiO3K2qdZcOhinYZ+fQhzTqH2NZvG0wbVW0iCc7hjocXEWH+Y
uzQg6L9Ec7NxRSEtciYeyjcrFV51iGhw7Jz4+69FJo9ymwfnBjqa8JDVd5BnoIXf
InjlTi3/DubLoXIrX0m83fQlAU/jzzfjSnyVVIIQUxXcgQ3N4/lhF31kn+tF8MvG
antmBRuYCviqLWoWmo6KCMBjg4U7pTodo8AB4t1jf6H+JyfWvfamNwO12Htu8zjx
NUE01a7jxcCuYtVi5+FT9KN6PnZbqEOH+Ye4JPeGBbdyU2KzyAXasL1mkHMIz/ZB
ejvO/b2trsV/O71Q+1q1DHOdHx3za6QKCckSAQqd9fGcC57EgeTbY/ahUOY7qUhI
UoC7NtNpM0Kd2ugkeRqWaG7fE6qUTiFWwG9oYuE1b6Y6B67igSkS9uzISE9vg2/y
nqeAoAiKS/aCE58YkJicDSN7TJX45ZFdwYskyjUtHN5G0RBAG7Ai6IQd3YHS+R1M
9FSW1Iv/xSxTCAQnBdyug8yig4EvN50mm/av+GQU9uNZhNWBvtFvACSOZxhuhgNE
mJ2QMAPf0rWVrPo3qFtKC/IHrVtqeuuYOlipvkefxgcDdkpO/WqRmpLPgMZMvWrF
CtFUS8+n9RUXjHmZa8P7wl8os6lZkACxXVw3cc4E1PGGMr219VDLPrZoaa0lyZIJ
IiC17R3LJmsFb6372joo83N4nq7IH1bcIxXTkto8/AMxLPI0D66ozVWlwCOHSNAv
YSRHaDiMsE4gWd7m3XQxuhy/WurcIm/44ATN3sSQDX04+65QOBPBP+u0JJ/T8Zxn
+yxzSPndKsAzdrNmkupEoRJiLA4QLCjJqBsNcjEIcdgCiXcdzBIX3W/KKPzQ2PM1
hEfrjSvkQgD7d7bXLgycX3uKqK0OmRDv6MWQrD29T36CXBow0FYlWv+eW3y+BmZM
SrOWgnPvtzy4cm8TR2VyYMJk8zre/xCuCmIyZKItvdD8XePrTavB/0AIXZfojMje
2hsMfFoDA4OBMu/UF2NARzfx+JztlKNSx0ITxES2+/Hpbp7REHdjTsJRlZNdDfHS
GzULicE+ZZHfg5+03SnLoidZiXwa9F5+5Cx0ijDOHCiDuVyLHiCoj2Z5yWQMmRVU
8mTiNPGoH48JThtSMgv2qJxIUrbK+iF19JEA9KMYwynNE1RhieagIGdm/ruWanmf
GkenhBRKl8BcvE5y24DX2Idr0NevPXhfrdng/Yiqw1hBzQC4wQvKfcbfdlsQxmih
PcB3emPs00C9VuB+QNkjrn+tMepQmt4w2g1Zlx1pFnEfqV7IWLVh1a2XfKd2ChAL
nk9mDDIBBsMH8LrXatoZ/z9uz75c7ZwSiLH2tlfRGzKll0Y63xRkT85P4+6vDbtU
cl8DQpNVQfQhjRdawDA6kmoJm8SdwvipEwWfgA30Ua9o0IYOTKL2BXsNipIm5BI7
elBev3gJaO3cJrHjzaeY/+ZLQoZJvfNDcyrMnr1UQMfehOhK+CPAQQUtsyB3LQYS
LFFBYnSoYGx3/hJ2T+oRf1vl+kLDkeoN9qaXHY9CayRRd3lOK7KzHsVqxPSH3HS/
JSWDCYqYLQvO28i6ZYzY0vRql6Tj9IAXl8xA0fQ4pLwxrX06QZA6jBLM8ZSTLK/5
2QTZ9qrohVlAhqPcyeBxTErb+B0GlLxhfo8HBmqw5mbKVStgrJ2LARabC2x0N732
+yjsmTb0FHjMm/C/FRUIU0Tg9CuISnxW/2FwELbEcVSJmHEnBBmct5I8e1GomWVk
/co6ouGpeajVaIoqTrawSAZc//CV7rlg57kN6iOr3F7JEC9VdfxmLVi9QAMEnDwJ
b3/sipgxttgrP/SDtrXaMvM+K0zaVF2ILDtB9eqtI6oCxJp5aDMmacolfynz5+Iv
UUeUkzxvPjpIGwzWaxHoBZuBYJrT9ygt09ocJIbizJd70PLLqExehk1GweavW12p
Vov82HLKHrN2TLb8ZJuIjIw0AL/YBfq5g8QcP0Dkp86Wjh2msZlhRtvffoMSmu6i
aC/Hvm6qa+61DszqSQLpluSMvTIcg8rT3verPRbRy+Ft5hU25YOthM8OEXkt/yeY
1SS1NXHgyKA9yk65daQvp+JLh4CXDfY96Z4AJ1hkusGc3Oo7SEjuthdlkttDNNLD
tSysddqQCsy1RczJu1fx6GDOTvjKtc8R3AXev5iR/5vR1P9pV62GW/BILKpjiPqE
xnK7lym92vVSobPgj68RcEBxkDXX8mQCg/FXRFk7NUQ0mgXw+uMbn0VAy9eSRpcr
IYgGHN5M8SkiCI7aCNXKyLI5fc6mAci0Fon5hul7H6/aE9rv5AUU0766HuLtfoGS
y248p6/bE8OAiZxgzblIrAdcpaUs1nzUiaA/Ovg3uAOFHipipvebGIKXcTwUjsme
Sqk7kDSKOTIsXtNdNEh0SjAfqismOYA/DJmnuoU8ckU8aeN19YXY1rymXZvSdYg8
tYqM7i4QQIHjAlh293J3dKwNLGaiVIY7DJYUwA3tk2cYbdmulJd7md6h/0WePwdv
SIBPeIbuokpCxpS+rWg4qnqhFr2Fl1K4tSj67OIAmaunCjqCJyQ2RQw/y+RzZz3X
R7JFiaSrEwIwnR4tF9wpDl008en13QtxWEolwcsaaO7fYu8e9hKjaFPoW3cGxWwS
GyBnPYZY+TW+bmM5ewLOYwxB/qH2wW9ZFYRVIyGZQMWXmWZSwmWPVAgVjFTw6k/J
yTn2gI3PvmmZnFZVD/MypecAsRXjzJFHDKt2Q9IfngVwmfzMJeBPnyChq58iuoRD
cAFMNVjXTl1zX0Z1dm0TuXdvwT9yRgh0BFEHuQgkWGEtgFrKfcAwTaRc03ycx8wW
Uuo7vZ7tBM60/Ei4Fi9yNwTzZPr6XbZpqo6shY35bduiuct0wTLMBhwyjDv59T0b
Qo8Zyj1j2BOMzI+5JaIJgyvHA01kdj4SvxyY6ppnM5S1oCsp4LQ3yLCh8rUJDODm
gQ0BaTQLyP8sTd+UsaBeg5v5WleKQXXWSxXElROFJOC5ETD2lILTRdQiZEbTk0h3
+idgiwU943GsXEgeZMW+YsfoK8NJNJWjZvlLJpfNGZsfqYT9iVaA8JF+OxMhVO9+
VYBYbL8aZ/Cs2SgChv7UwlpGA4qWhp5BOsQNho4yGKCdId123mltdDUK2onSLlo7
/zxamGQD7KkCnxELbh+m72iWH+Uha/RQky+vOFOixnEJLpx1lZ16dl6BkDPDm5vm
WRtAA3u4dTnBOuinf93+ElNFarNX1LuqTcp5Pyp34xRsLQ+TDavZxYUqdyaQwTwz
bhaxILKbbHe43ESEcyR8rpIydkH4mX506Ep7nkaRtMEyGowfh1Ok/BVjsS6PUwOy
D8AAl/fn7QtprckT9OxCWbQgYdIktAoWtq6SNCLg+3wSJVR10PZNR/npqUfTxK53
dCqMAA0veNVuEZP5wi/Gr8f3Qy9Hn5ouxd5KjpJx67HlmCmvf/OLJ+rSJS0RBL9R
FmwQXiNVQSRGL4jmRdgzFchOyg7T+Cl86L/N4/fo+z8ugXu/elL5Z5qHjcOdSiTy
yUzecYqAYS7PNutowa5ZVUoyJIf5WGVrE3JI/HVDZ2eeVN7Ev1odnGCS6wddfRyx
39t7R8gPDAEn/kxC5+kD7744lDNuRxxmpTGrFuTtVuZB5hwMuiV6IMc16w19PDcU
0b77VS2fT15zsr2Lq14pHZsGYoNoY1qZgLsQ3MUnTBEjSN8O1GjuxM8znY3f8XEu
qP5CeD8O3qfdWKbFcVXuucJMiOX6fcnKtvEh8/0MLab1qFa95Jri/nSL5WgBIRvf
ZIMPyp35yc2bOrxfc7F9HULwW2r+VR2wkgMC6aUHYVVPZEMVaUPWy46Tv8uJOfAN
Y2eIbfgC8sqD83ZmIGJfUiTR/zBneN1KYiVoHH2l1lLai0GZ/RLP25ENZbK1wflk
5bT2SeonH/Pk1U/T3TWHWZa5+GDS3v0kdX4MufeNN4zkik7I/b8oxua8uqXKybPP
loOWGXQJFN2wIvVaiTsh9Ez90ng22txA1CvE+ellv8/9hJX0mBsmlXaaAcwxm/FT
zgHgtutBuEzDVbkAScijWqwtnqlQ+jcpNBe6G7dhW588xiIvK0YLx66rTjSGO7z1
DdjLD5uBIVdDn/LXmV3JwaeXt31WlfbAQdG6cWgm0aqFVPsT5tOfgWJRuFfTpopc
se13n88s5/B6Aw2opclhsHOPiZleM2oWfd7HHOoDzLEtii4LlnLCKgEJFKQpW6Mt
scqzTn6b9CYfp57WVRL5zGqOwiVUH2gO+Ov+xYWsLeyHUUJ3RZ81nV+cET1CzDuT
vcyAb3T96jTYJPGJU/miw0++j7OiogpLmGnjEMsUA8wjqbDj6dg+QYe5eFfvM+CF
Ig11m+Bj+LsOMxqEmKGEnUvxE2bsgOWX+eJ/QuRjC+SmzvDxbqzA5BZju/i2L0/p
QQtfoENxUx9Yvrm96iTaeWBp3HqQ0R061wUrUM0yF4kRdJtWB/H8yc7CtsqoXBoz
xUW4DyrnK3cMb8EARmM8krJN4lShIAQSZZvWn0rY4zkqwdacMY/kV9UTTC7wgPTO
Rm/px51uUXQj77/42tid2ePEH2u+kR47uHgXJQy1TyPw61vuryD02OOiDezuDCJE
uja07tfkJ7R1KuTwwPaOUE+jmnFeqHlIWADICTVj+/z3Ur2L7JFcOtYN1uzQFU69
sc57N8FnbaYD06coqX17MGkBy6BGtxSIkLMjMpUquIaU0CkO1PxIqh/va/3Nfcd3
2rnPP1nJ3BWi0mRhGdui1M9rR8GeZIhYsEuenGomiZQLcsO5x8Ad0O36/suoCJ6+
garvQXC4zR+9lyQDT5rBQEwF1uLkcFOLSSBQZrr3QPt+XSydjT2Nbg6SL35zHBoW
KfI301v0qYjvvFDJNwGfKsGMlLKHZJTuc/Ui5uDxf46gk8WStNYfxcHUdCn+2F4I
7aiBlVxpOK3MoTZkKKjZ72ixoQeGC+qrpuPqVyDl4VtZ9qSex60my4mp3JbYg3Ah
TWiHK9Ta22pi5nuH++b7upONyzS1RL6w2RjWU2kB/mRtrmP0aBnJqhmGVRdEpcy1
w/j4aLdPn09KAhdRBtVeVN3Lgr4nfzM9KhaKZmhbhVy2gcjvs9UXCyxEbE0oiiZj
5/AZ+xtsDoYml4LJjhfEy0+Kng8fpn+Jb8zkHomIfyr2PfWv6m/M5PIV3gfKxIAh
MAIOjgXKnnBUIxabVfvZHi7d5jNK30JJYScIE9uAoG9szcT00TVU8pzLVFn+waL5
ANzNV58dMTwBLsR3PGQWbL9skXWsjIb2nVFVe7d2rKEgla6kJkTHAzFkdcG5BxZ6
B3oSn/D/orX2GVKbUaEuSRuf9TUEzoJO7VZWePZ2zMlRyer6gd3x4lhta8E0ugx8
ThuybMtgiB3g26jnzOBAIBDwLv80wtpGomGs4YTV+glBzBC9jMEGX2bCf/hk+D1c
ekSUiGz2pe8q+Wd5+LusrTBa9SwPnVT6e2Xnrcnu8LWw1vjB2VdfeUPJYlmBQh0z
N5mTuIgLIwS82ljOmsdka3txOJ+EiFr9agPKyGnjaA5XFkptKkd0fOFUFqXEvpSD
KYto/GK5BtidWQ9s9ngXJCTo9RzF783bMqCGYmdRZN6snOis0fmem2Vgf21IaKO4
DKj9q/zwPeeJFIsn0IdZfs9Yc14jHNdg+olbjcl/kE/rszKBhGDqujEjcXvSRGFH
JiKN3ru4ZowlJ4z44qqoxwI3igqcQWLMmnJ5jircfHwfp7HArmV/pHeDzu9Muy6M
MzCvbJt+r77WhoFvZlip7cDh+qX0VAQFEeCPF9B2re/8yykh+HfwIeB0vn2MJ2lb
GdiQ7a+TgOG1+ogFQkkRr40SWSWrwMRwIVsioXfSUQMhCVTBgARum7pkp8T6hI4I
KJaHyx6KGj79J1PtI3eSgCkyJq/iTVcPSBalfViJqJQSssuK19Sq24f9HBs25U0x
6UyzcfxGPuFgxaN+/UCEM33WraNYqInV5TqCrxW1SWcRKg8aSo5oNF0c3Xa9cD9i
lDeuyeCuAYKqKEvkGw1mXZKp1lJE+ZAJEk8YgfqTyr5kUesrwpqjvEiglz6X5BeQ
cGglg3GVLlqRLomvB5r2Rh6cKrJugkO5YKskvxlw+AHbTbUXG24iwiJkO4pk2rhb
9KQm+kAvz6uNcwQlNkIpzG7AjaJUyD6kDu7DBu19SaS5YWkkf+z8CS9+OAevScGE
r/0RwULaEsgNwia3LMm6s5wKlbCgQX5mLAqfHN32n2o/w4tLZwrVqobYF1cecSRz
6/688hjag1a37K2KmhyVSTq2/2Fh7L+7ZjkmvEIdaY5guW+ogQSC+gkabJgPSN8E
T8nwT3B8PiFdqRkUFlhSysXmSr77doz+Cc12ZYMErt0tMolCuck9cqkA+Iq6tcui
SrvsEH1nH/BOBnOoKYTibjAFAWlkd+UCZHRf1BQxj1ilpW7AXUx74vwh1TLZ6jn7
d22baMlhcMCufE6BYsAD2u8x0dfIkvtAKUveu4EkUsKL7zPozchKbaYWPiud3SJW
+6PGFpwd4yBH9xHXJfcKVUxF3FBoDXqAZdO697lu2am4jJ3xynvREVhmfLZqs8w/
GILqjbvaIUaupwU3LvpdWsiW8yw96h/7pFu/7UPduYpr1Kw8DnF50sRfoPMlMaUa
e8PpI5SElJPC3HSmtjHpc6eFjnUWvV672aaZapdw3pD6/qG6aX7ptcU5pc27c7xw
gvCVQTj/qyM39keAYL+uzwVKMw8PM34EM0qR85xnulByXeUhyNsg4CDx6SXAOv0P
JaXt3bRUE6IFdQ+8WsKPVw/tSPjN1y27dlmDcKR+CRE5XvmffC/rKhuAlW/AaSor
QR20Pn21x1o6Wr/16cYGPHvBn9NJMW8LFNXcIkVcsoe6ADDpYi2aNNdN71VHIr99
q7C6zxgI6jvyZ6mhkGXz382CLEu1MnW6jEyWxB5foAu4YkIaK1jL/oO8gTPTR5j2
uMDIx5UN49tlNbz82/hrQYFV9YlRGqZQOXCQQ26p9qIheLoqq4iX/lzq3aAKrDJW
sMIe2I8cKS5IxdTEIfIAo7F0Ckv+ruYSlxWiCFwN4JJOihNBb7tjDknI9nGLj+wQ
3wa5hbf/Da3goEtk4dzNh3pFT1Bv6mmz0loElOz8DrF3DRWvQaCTAgoj8BeSoE8V
w+yK+dB7uWI9Bp46DAikt3blJNObDB/YVBxdh8iW3Ejb7et9qy1tEafNC6jgJ5pY
WIbJ+fFHmmFMIoovtr1zhrD0MbJxDr18e14BR1iKzmhA7flyheFGKlx1jUibxyay
wEeO8DsbT4sDbi0U2OmNv0Y5x92GW6I9jxGgCI2hMlG6bF48scrFNZQS6sksbPnm
NPgdo2jbqwM1avYoiA1e+EonZfGe7UvKS8125u5JaQwiQta74L7+1PzVOppUmPuv
rxNtVTc1KtTHVKHGT3ZkQeY2XF2ZsxrzSbHo0pHruBv3aZS3OehJ6W8Gvu9UQonl
nIVuv3v5+4t3emgfY/rOT3hnhT+CBxZB4fzNFMen1DxNp+XiDJoRKEhhFyBFzXCB
bTlLNXE87bek18I4DLP4amJQEjeTDPI1bQtOi+RzxQbx3Onh5wxtPUceGNl/3+F/
9IMQ+4y9jt97EA+zz8MMnFFvAmG7GXbZH3TLfDqWRXKjt262Xx+ZX/DAtNStANsj
qE9Dm7sMDu2txAbr0BOKjh65iM53yJH/R6F6HRQA1o8CkVGNSBkLYc79GAJBaasa
cvyJXsS8zvvBudJWwsht9GI4E/xlYLxPMPcVbCg9Fuu9V0rtOVxReOj0A8D1HU6p
R4ZtDVJNpNLTJBrYgFG+Zf83TM2dbd7OsyaR+vtQeD+fLo0MDVsIr3hhOAJVCwIC
xOsRWmjkYLdJKgbrhKd+/jAfvvrsvdNct/rs6CRlNcYJ9rdxJBLVTNsGE+NPa0PZ
Tfw/rLOG9+1iwVaW18mImlrpkLb+zNkMxmS2F5uMyfv2j7PjR4gLUbEDI3HmCOYl
xfHoLTDqVsmXvcLXPOZXrctaiI0A1Qxjqc4gZ5XjSPw8PA8wIEUOkD/A2xGydPXF
/y1ufw47SsyOEZx3KLsDvZD2ROsCKmKBLMgaS8DqqSSV2j7ZJzRDNqjIOEVEBQvf
Tn7rpu7VzUvmOb+pvTF2RydzIJDC5EqayulSNZ/2QDVc3fiyt4zSoy6QxF3iH+SP
wxCthkkTHU4wQO+yjPcATeodNs8/6200HMJN4DJ0EWrXMuaK4ufuzHOnTRrA3fb4
m++xcndo4bSEm0h+bYeMNa182Y2eAKpFmkOmtC/ZBs1zfX1zg9qaIj+KsUPcZSfo
/VI2ORQBbDnuHLacIvcZx3ZCL1ZvIBvHUfMKF0pGsO9ESpIkimFmd9wEIPV7g752
iOmv3Tq1sxQ4BLD9XR9imLkZy+vgkJ4AmIY92DnCBEv+BGYF4rwbeEY0WptPNVBk
dSp+UWLRv9p4+I2cdN/hLr15Nptn+W+L0mAd60s6m3FKqa53odHBymtWWbHX/5DQ
Vj0iOB9o1DK66Co1eONKcD9GJUA57hZyQR70cyHc8U6AZAbrcElVDyfxbSaOP1re
3teGVO8L74a0SXdcIeXCZjojaLAApYmTji37lp9zdZDjVfMNrCvdDxmcyRvjOxgV
Jtz6+K7eGdFa2EwFpX7+dDPqL10AGhcrRHSXaapTSznLo1ESf3UVXFkdB05DdxOc
ToH5Z4hCoSWagppjceOi9oRZD6j8EZwkQbks1gpsKYHfLF8lIxvT7jmvbDz6EnXO
s7F2yQ5QwJtf+ugdOeGILt/w7AEfFX2K8X0JP6B33P3o6lVkhdyV10UAlMJk5tV6
d2Hnt4EtcImHsA1ypDhhpiyKvoT4LfnNVxnfKq2gW2cDY9R8ZaAYD4mCFLHHGh+s
zSljbrMMeLzNacvK1bgb/vylp5/WUEf5G9UKBpnqwrDqyk+Z+3OuQOgAcDfABMbA
1tbIGdk9LCdw341fCo+LPyp4cYN++GJnX5vOROTCSxGYmpe2GQoqyCCRhs1iEU0S
pG8G3+2s/MC4WAE2pAkWeJVwOtsnR54UPfyrSweBnrm6gKym4kCFyjRN2J7GBD6x
QWbUZk5DrqTjJu5yd6W7WAgBpk6fbEWUA7KTKY/H/sqG3cdRNZgtxgE8LWt8aWPF
7cB/g0LyfzyGRmx5ZKZNQrhjtI8LAvI10zbIMVVc5L0ywbUUZIu2jvpcatWO2SJl
O7DyWL3z2aonjUpnGZqaYG81DvX7ctvkR6f0nijmFJO1RodREu8Gcih9VTBkhyee
wI0Km9obgNxiWx8dOaja24n1DsKNiGWZ+rheR1nvm/4mbnipIYuL0Xkb/Rp/Zo+N
fxjz3Od/xBDpbvd5FFhR93OJkhg1kB1HzInBU7VVxw0tKvL7zNHKVcFdr/mY+fsf
nxo/tB0YR0kktmRBRwKDApcuLloU/jUeMYHCErYMKUvY5NhkRW1oqPurlpTetvEP
yc73ZX9Knc/L7OBmG+CyGIQpj9iiSFI9zAvyfLnC/A/XQ74CKBHrQ4n6pamDLLw+
NL6pAiy4e1uhh5LPT4qBZ1ib7paGytWHEpOwkhEmnPKUE+JfbT59YrHDXOIxmkxD
0jOQF+PGrdDej2bpMl1r2geeT8ftJeFidsf+DZIWx8MJS57klLi7hCVDYzN25pmn
FjTIEubPu3mzeO3vSS7T16DX+CtORUwA5UzEMFgpQekHsBrT/N1jKlB0Y5GXlqoF
+5i5xMoqXRJu0ZtlXlveEWxSKpO9ypscMwUD86bZKa57K6DQhVU39LMVdLpnQ6TV
RTndc0M+EhG8QtQavrLG1mi7Mbbn80O4oSYYPFnHQcRfogW0R3kFYQyQu4Y7nhbw
L3MmfG4o6fJ+/ajFSn/tMOQcFiqWwG9L3ouMhwYSXyGPUHXrs4MGHSTxh1ssr6Bo
awbLKN7xTdb+Sm/vm48P7gsanH3nuxFNuta3TDl+8epgi1txcMAryaxbL+n1be1K
zvSIoUx0Q4m+yUPzsUesFmRVWzFCBPsU6k55waRxj7Lp1ABrL6CjPgkDW87Cm/O/
zjVqgvdfG4IAN+hndSNCve96vzxjdma5qST9p9EH/bIUIrv3T/AKF8HJ88WAWE95
9/txtHtIYgEmFP2R8o37+qLtWzHvAOuFXlNgPib2Bfj/lljrdOPsd5GLTSx2UmiO
owHiXacc5QUj7tto+JozGRkQfQYi20mG/h0DDeQBnu3WdHY6M1FiKcXen1nm2ZNH
FlX3y6cxy2nrctlh/3NrBvh+B9Q2ia3ONk2h33YbU2R52MlPHwkzVML3eCQEdLd3
B/kutktem2YLPsZCm3XOHncOTEQFuMk2z/bP5Q7Bp6iG93hT7IBXMt7l5stGP28R
JL7nR2jLnMOujJYdb49JszdnXNUOLEElS5gcN75phs/gtOQ8jWw+HsvY2rIbY29a
c36skSh0ulwLjh8/k++y4vezPj6OIml3TfjTEMOelH+3tTQrTE6A+u71rI93+HKA
H+aM1ySRlBr532+j3UN0JudXZe7vpuLegygWBpKYwkZi9k0LFCG9y7PikL6LUWx5
vyYpZxpiTh6JUQCEmJWMv6UPv+wSvSF35pBZY2LyT1+jZZC+cKT51apmsrdeQzak
t3Vv1jfqYXjBL4PsQlSh6QJGRto05tP9V+AzqwsirxIaDpggA6X+61vzeGAB2U0D
4UKi7EuMxHuSVEC6Uy8UI30DA65/dArpNtpueQ1G/wahecIWV/C6m7eOor4qN/6l
gjsVYKrNn/M8QkLVbY7tc3kzFkUN3lt+ASxzdcV42xqQw/DycBrRKehPn5gAXko1
nt4ju+EVu4/r3l4yPF3pk2+FIWfFqcIcYYl6yakwKE6JG7KVXmvLVeCngYT9rEpP
rQz6Zrnv8MKjfaZXy7CBZElH0ws7eeqa0ovxsb4g5ze6Ese4MkX6fHAI1O+2t7t9
nlsxTzB/hqnsq2faDK5x7eUcCgOaTVPCk6JeZEzt/2oLcOzs1lPz8eMbVIKwqdOl
aZKwcr8jlu9SiXXmiQa7lw/OsgdgOYK2yKOWQIb/aRomjuKpqG0N0dmICRZoeHz2
vWxfSxJMYvDf5R+i+ASamtrhpPnLgC/Y2taAa9sASOIU/gUCNepZmlsgPvzL6+LD
aZpE81zMV+gZ5SR4eWlYhCKeKWh8PRmUZl06/1kUAl1E5a1meN5nynmaMsiC7Cgf
9hEJMbJAHSuPWUSTyuuBPx7A2bzZKuBMTg8L9Ew1UMGYRjFHveA2kLn2Z8FlgVgK
IrU/Pn0jdomX2vwsjEyXwT9Ql3F/CSbh54rTU+cTayhMJBu5HNyZ/RBu87sWqb4l
SmOtCni6P+RbTZ182SnyaYbBL33YE+Eex5llYP0EiBxUZ+FGZNUSknuwEsy6N93n
5x0g4X0lD2gtzvVtHkwbFOs41KLcnKkExQDNAppCTZOvHp4sr+RPgVGBT799OOZU
GwrMUxftYkWbJrRQn0C5qCem11koJ36oa1aqKu7+3iHL4sF7YBu0awmd7CZjplng
vEs0tgnx2iCON6vFrRoN5U7eTJDfmqtpqyXwF0HA8Pd7SE5z0fImDCnyA8vd+8MJ
u5NPxxncMy7TdrDqBqD0cQIBl9AjREmxCWnCPpvzPCBVZwGXjTUiZJRrLm5qSpux
cEaHkWRIRXMUzs+le0sbOZgaVvFs9OAk1coMUHRldEXQDTlJFxHc0I4/EPsfaNvy
JfIaHGalOe355N64Dw4/AM7fPKIkUabM67Kg4ru6xiEqwlgMl8hA/mf9/vtamxsm
33xphYdtDHWW2JS8CkD0K2N8iTE3tROLbCv61TDNcH2qcq6mwTpF7GzjccoHnmPU
D5oS8CakmSh5ke40GRQqqxQCPfI/ehORSno4RAYE0EpwnWBHgMgYKkPD5ozdCcX8
N6EoqToL06BecqCaYfqvaEuvFWcfFKN9i9HHqtvtoYSjo46eKAPHe4zmd6F/FaRL
pAhcri1eFiay+0ToWN37Iu3qkkj6Fk1MRL4mwSM1LOLeO2XLvyz8SHxp1LLTAYzm
AcU3v/ofDnTrsz8cj9wuckhC/J7tHoouRoCwyJieq/078AQ9c1BPOBcmcCSKWHKL
u9C+2c+XVSRkgbLRoXvThCfHgKkxWYc4t6yozMtMhgxoDzQpOotzjswBWvHGVaoa
398fnAcgSVjYLWctasdenUA0EVo04YQZ1vAvhfsuFMa26CBu3EGCGg5nO1SxtQDs
NyRRVtAyWFJgZ1+pHHIRQYbAbc/0JS0QnbijAR+U3EzTI9+F/I9bt2PkYsGXAGYZ
iKHyP+ZMbh/fY0ugruBJ50R3WyDmuVY0toDE67uxrUdRSRND7PQ+5Ua4IJRgkeGu
D/QqvpLHztModcv2Y7QDqc+crcvF6/VY0NTxSaWCriOPCjvemM8GFo5Z/G3UrjRT
by+oesCdymnu6nm9o0EMu9ui/WMS05oLvd/wPptOsKi7O6VQGxNkUP08h9U11lMv
hyl1v3XFIciYzPKv7Uz/0Tjq/0HAI8vF+qtdJQy4hZO5PVV1/xphtcQtln2txJH/
ixUeMZnwh+OjFoSLh76Btmv+M2gx+NKlV66Q1Z7aXqn/ODYEizPtLl30dibRmJp9
e2NoDtN2R7NZEWNCn4htJqBUh9NI+E1QzpCcotoLprq1GP1OJ5k1YU3HN86AL3O8
U+PnwH0jTDu325ZODc6gyTldCPaveL1de5QZHtWNQHZavtD06s6496JZLNuTqGFY
1yCIW7a/ZOFhvFii8JJt/VCYsMAoXW2WWdp0dRNiK+WtwZla8sJLkrKaNN3dzH2/
ry4ZEZNRZ3hH982Odek6gvB6zQVWJum3Xa3+R7EX+OFeWnGxT8SLpxYXKmWqdPq9
M4suQ8tlPgYi3EOaydhKJtvqO50QdhSXwHK2iPLKAye25nu9dn/mA/p04iwpihb3
MaTFIv9oJ3qIgb647Fr37R9fhohHw4xbOEHCBS4qn8gINZFiDIigIBrkOtQtKVcn
VQZfxiCkpxaOOrRq38cyImYRrGUF1oaS3DDM+SmkQXEI1h0QqaQyCJ4m7T3cL4ZK
YQqgPbt6yziUrkDSKb0LMgDzHsCQ1yKcX97FYKLyl/oVOhIqe6WOdaybz9bSEsbj
wUM5hieQeUwf7Ntv31O4oF3Z8F5R1f6VxoZUpEWdC/wLfO8nxBq/E4hQkI4ZHygZ
o98cGqqRcN+Gbxo1HukRnXNzAeYb3gbWvkZ/po36nVoCZZajZ9krdXfZFPJ4eVVG
yGssfr9lsaLKh4zUeXvo33cOBRN8Z3BQO5/qyaCmT4Fh8qSJxww8iB1CLi1K2ei1
j+V7J4TF7rwp0bhIIF6jw9SS3YY/Uak0TkDUKElNFmXOYKc+N2224yQ/3kXX4JG0
HRqYzuoPyLarUSt7SGYYoOgtQ942M563Smr6goBaOw7c0Oxuux5PxyyyHo7EeTBX
eFhuvqu+2Tc6T8/r5n10unwmmFt4gvjDOriWPfLR2J+ueaIS/8hUONeoQehuDEpK
yRVh/pIY0je2APZdlSurl2vmocNtNEtOntsmHv3EJJqdIeejVdztlY8dtkecQGXA
rH3vUnxkGTRT+YQ3MfKRckG98xZXGgqA/uPQMuO/N48xNH9xX4PWJlXz9g66uIGO
IdD9RPbT7ei6wVGlQiLbNeottA5rDQrjXtFBAL3hm7JsHRyBhPwCA7MT/KT7zejC
p211z5fR8o8KUgzM3WNnQOZZ4WnhIU+Tiwkk/yI0x6vqBMyyqnFkL7rqldMqKTC/
NgfcqAmMw7Ok6M64QzrmkNl9ITltg7k7fyoyNHsl+N+duIHSylt2JPRkK96fkiMz
nRucn2yjEPNN5i4Nh2S7Lj+J/4emrkAS7K2jJi8PzZ9qGG6UOmIzWfIazb9+z0Og
cGKfjp4nwVolUkpvUjZxBYbIwXTNH6ZFQdWOnwS4DPdDMhIW/BbTMBbLrPchU22s
BpiW/THA3czCwYUVcuV2UMpFB/rht/v75eiviMXGUN7swKzJLCWACdwXXu4zB18Z
B8R6RZt7pXGexxy2qUFqS4ZzgGzTprTGxu1mBXmStCJc7hxQKS8+f2E05KGB/ibC
S2FnbxtIpQuAYDsBR/YI2UHSy2JLs7sBwmTSUtdZihrKL0q9OTfmfNbPNGBxifWV
zMmnRdUGn1mnouRGKuIgdFy2yzUgXYNG2+3hSsDD5brAszVBJsjQWkd4E4rUrO0D
jzSODWWJlsK6AbARN0crb1BO+xmOjFNAH3qTQma9jwh837cM5Nly+9eUKPxRc03j
hXPKIKuXILUQnS8QTdG9jgi5I1Wny2C9L0ntgSmEsMoy9sozY+DsVs+HHK9ie2ZT
Ka37WaaUY3oMyMtHioYhVfANXy5LtMGPnFjVqK7Fs9mL1KWcvfadbOGRT31xjWar
Tw2ty846iSvQxbAImQFVNc4tkvf6pS8dCKjGaEOeust2wQ3s+HDaBv2FM0XrU5Qp
ESaiOLUiQ7GkkBGH7LZrdVBvucwnnCrWx1hdCoktjOFNhzCpNutEW/zcb4zUtova
Fs6/vDLPXEHGCTeamZ/Vqed7CAVo5A7FrYfq9yjmeM5EZU7mSy0b2FHkkyHT04z9
NIBBU4UtlVIqlDJmiv1rK5kQtb/NvFFcIsTSn6/EHy/NfD4N+DVyu3ywEyLjv+na
SOw+tGwTNP/jS//xqBizzI+odKCbzbeNpN4Eub47aCoIphwWqUc9gtMdAkQfSNUZ
fQ7vWNN0Nd5TagRjqKQb5R7g+kUi64lwxuZvA9oEadZ+OD7n2LkoxTt0r2AV9S48
0J+1xwMGpUBtI42XjGCTxgKdHXHqw5ku7mbDxmEWxV3gvfSlcgXv3BtursDW2mBd
bMO6NAmwR9vjulgcMBiNTfLTie4XTwkQNy5CyIyM4kPRvE0Roc2k7k25mVhtgeAc
Vs79tdhcnE889ulAB3aaAVALXhU8v8xgTwszaKFwCJZSEj+gDzIZsHYKIVK7KGUK
kJFQLpyjWwcDP1a54o88cegWXIjuDVNcCQuKlueasERRQpVB/8etRxpBmVdmjuH7
CVLaNMlT9MXJMTKrgU35DBA9t8QhN7hXszhZNhNb2t+yoWN3C9S57Fle0pGqLhv6
V4p/erVNZ0Zkhs6/DpW1zm/PadhNspj8uJoOwKRRJ8IObsW+lQaferuPvIoX13SV
QLPgPr3RPXwB4fAiJxdmholgtgXOAvCX7+wJIgS8mj4PM9rFlqCOX6BRqkMgOJf0
HKh2KQtGPyM/2ZELduju0zHSfc2pMxvK97c2YL0j4JYZGRye+xwOCfA8R3b74UZq
nseVJ86olgFoTwZYotXIimywVnAkwNq1C/khVYle6+E1npG5KW505uzMnAhUzR/b
GY8aTGeCsjg4X4c/7H3va+n/77te8W9ERSuqxXUFSkjmJhxONHyRmJa2EeYH8U6c
P6pZ8V7nFGGgszc0X+TzjlnmvPVmWkATcvR/xNbzr8IoKuTFWUnGPfmezLDd19fp
kMwhGMwy4O4dwkyD6q5+59HxXdRyezxUOJCkWdD+iq00PNB8rCxDAZqLcF/LZFze
7LvxhgKAYJfsxO2Kdq79hqiP3YvljLmsJGwT1BS62c1eHoW3M8MzDVTK/FnxnnQy
9FA6ZDVix1a5zZZ46d4c1RLtHNvfgponjzAY1UXRpTHN0F7+FC3iCdXRlytI+kG5
fQGhYr3t5uql9L1GLeTdHM0RWunp7TS3Wn7KjZBmciyPVDlwwYnJ/HzK/ZQ81iH3
nW9yuN0sg33cTux+weVrQSFPP3RRxL0lHeSFMLB6bnLIDck3FUc5d4KDZ1rzuwbK
aT4iT5BIKWnTbYPZHVwq2JEBxzbQK6RAX+8xTjxRYzhRNjnPYxINhApgatILuigi
wh7eQzBjCP1OUFn7GrmAXTXEpQLeAHY40y1Rm/+tAHjx8nxZwjzTVvgILMJ2tmAB
p256d526pJtpoJx60ESuu2Iurea9e41KIENeeMlIfCx8HCXqN0XDp7rEaXy5o6eP
M4mb2Uq2p54lyK/SMKDTyXeJOi5U+IFgAnefd57yqTZ0NXUYFs2KxLWM1+uqiTrV
le+LJ7f7zCeV6Em13XvsmUYkFKqDKGXLsO6lkI+H11UzzN7VQ4oQ/Zwwy0dOeQzL
+MAORgWy1MZ6dOSWSnVpzpZVqTGVUI4NEQyD/+eyYDHYrspJGM7o+WUSI7i/2/no
PICLsovnysWamW/7Hyx1KE4el6JDgk5g3GuUbm7RuLNmlEjE3aoL/87c7W3J3I6D
rBWupP28VRdXNIQKAtaFnEZnTAI06DYkfo1yWonm+H3QeBDXemQmfNmXW5ys2H6Q
Xnrm/UHnLTIOxpEjVrat+epSgilUDt0f7l0btZxu1lDhu8tCstZkfX1rzvh4N5Hh
vjFkWjGY5Hx7KCBLzlf6Xsm6aX+F4ilpt4gFJfKtM0awz0a925snUBeFMN9zL4ch
nNqKXiWGYgZZs6g0MB+sKbocXBqPTGUvmYeUoMOux3MOK5XEmcYgr0/kkfYGiCKQ
kvud9/wph/s+kXFiSrfMEjkHHGceJrK98ZiuAJn9LT6ZaC7rhgjrQoTJuZEeaa91
mh9b5hk8vE2D19+4VYTu3PVROiktB9B9ovYn4SzQgIwe2Un/e3ZKmb0NrByuSXLs
a48KmGCJc3WYKRbEmNlSu9u/52qjeBUyBe+/SsasWVOO0K2XeIW7taUbajpcRjIN
depzjHwo9DGGebf1W//bSGCVQCak2b6BJMfFhaZPP9zNlBU3/KpN0qf3JAqMWOnv
gGRhLN4WdOwrEnuUbVTcpXq1lu/6TduWk3M8kKmkNjKR3brC467lQv2awypilxVY
z5h/BABgHcScTjpgctxnTF0NCB+VFPq8Hd9bALU6qEwFuycujDmy1kX0G9aCEGfZ
9gxWYGGbfdfmDqL68cncLq9tnugcXrx71D2qC13+CyxJ3G/20M1k4O2OxT8VEfa0
nCe00w9C6m4l3qaMoUsgLYj7m34irTD0pCiv4qsJxKt0faYQHTeIvzHvtp2o6zkv
SiywX814JCuIVgV+uQXTufkN8bCsLOiK5kbjILqamgL/yuSm0Pi3HodvDQxO1oE1
eWx+6sXwItz+wkwIzLYgG3JUiYA9BTJWMpPZDJG5PWGYcA8vy8u5fomIx0xabh/U
UaHPFv2mUhPoHLr/ENcbOEtkYhRJQM7TnnJ1qSHET8QVHPhZmhh2GXzpoPYuRUOu
3/6GK7xBuqA/MJV2lrC4CwYaP5pQZ39mSjNCiuvIWMiMk5H7NMuLP9CSsxcePQ70
CEC4sgsDRjy83qXznhCaJ7Kr4H6frb2jTlbtc4TlvHFVTjJodDbsjkXrm1knrYm/
mUP0Qafh7Shau/uMR4PUAAm95wWAiPP+0NDraY5sPEGAharFTY5fqw6BJPTv0uEw
d9zZ/vvf0yWk/1QTWHMhu1fyoiAGLjNTG/HAFeorWduzlglumnxbGLjPDsEhdCSB
kEzPTLrn0UGjDnrUNDU2Wh/X2r6m7990pI8iMAV9DRRBQHN3EuM8xEPzjSndrTUK
mIAD+yPC0szBa7fFNt+rX+OI80RgX4pmLBum8oKzmBMTm1KT+xXO3uBgkxdH+MGp
3IdP3HEFjiQhFSMuIuSFIFo06pVWlS6Dg3l8D+0Yt8BZIr1C9OlDPLqPs8DRiVPx
9OA08v9wfe2I09mM+RwYrcs0QmjyVgVMbFuYOLNcb9oitgP/TpwR+NEkwbDN2GH5
/WfyeB/EmbRZMcpdmn5stEyxze5ICR+/8TmbjKVf/HSHjsZqeNQpy6t5OYfEQdo8
oMGorrDSuXsudOE/2N+udg/7ZrXj4/JZmILi2LaOeFB3fMaHj8jS2OnuUnTqFPn6
9D7oMo0syj8MRFfZU0LsySshUhfHW4rIixldx5p1oejP8RA/tYDEUD6XeRDSYCjX
WaR3VD6/tKtlkfJLjiZyKi9oDzfXq+DEEkgKXx6DJVt8Y560rlZ0VN9WC552jhqz
l0Y2Uccc/k+uwlIqWTP3h0rvtGWLJuBcu6rxMbwG1GER5jNpupiHAZJTXLvtd9Sq
hz+mW/VxpLzMipOXwXx8El6/yuwxK2GeFtOAVv/fmBX1SnWmXdB6Tb+9sz2WAQw2
ysuVFP4p7O4Eualv4HMqZ6YEr5O9lXBzhs4zP8+Jk1/ETWTogXlzxjXG6g85gD9F
8NUCcGcw0f2FRLB2gOJJYA2ig3J9HPBGrSBZS8Ct96bQJF+bKuETbP4XALlC3o7K
0sbY5YnfyNCvf/31e8zRoPFMTBmLX9Ebx9Ld8HK8sj+0rHUYWqFFUPD/GCHptc2R
+DmxH9sL4x5GBCPweQha8x4L9tLuehbmTPc8rgXAs9n5epiGhL8HVER/yw2IHKBm
vSCoT6KyG7hkoF6VCMsj2r+0Wor9TvVNYgnzwWa95V70lBrdFmywSydNSbiEHRbz
qT9C0k61rA972753CnXMoTiBe/c9m8mRE1eGG5mStHtBp6+ZMdWQ5Oi6QmFKsjpW
s/4MlpGexly+Uy6kjpuzEIgeXnslVIE4N9/FcAyZC6KWlZPgg4HhpgDACREnU1g3
M0PFqoZYZVHSKLh/3f5OM+MmEPnZGTdSc6fANUPnQ7OpCTaJTT8ylzUrCo4d/SZr
9yhONA16HkIlvpZtpe1P6rPWVObkrGvpraQuR2Y52v8m+EQEnJhTx/MDh+aVy4KN
DGOD57xLVrub9THEw+wqHNjnglGQSywrrH7Y31E+0KHiEC8ElH+1VrNvD74w4elJ
745zfryjAiM+QnMAVriJCbauwdzldY6IVGQJBJpMamp7alqqf2t3Q2B3M6iCeN1l
c2Of/SCyyoYVA1s1WiIawSFg7gObw7nJ4YWcW2gEz6/O09PsbSTxUkzHagZn9dMi
cKuiL7m1mKEM7DXMPB89C5CtPaJ0k3TjO3pDsrIvH9AjNuhFlMP+Bk7h6FTxg1zf
/8FxcgiwHRSvScodid4pJu8rRXRPpupS0g0J6goe18LaXkh90QSOvSO0DkcaxJaT
ZWONUr3FduNd0vI9FvC0Zpgj8Pk5c5zNm3sP7nhRc06P/8pQ38Bkn9IHkfqthfom
JIOEEk5tfpnm7oZFQxjLp8Qpr+zpTIzQbwIrypBGRlASgEdaiguB3rrgjHIx4fJJ
lrHYSnNqpC77/csUgN0xzYDXpkJfqwLMrtG7LnMCwlDCAxtCPR4sDyjdEo1zoUlQ
535ztXzFKa4pvYtBmfX4xuD4Q1NH3NjhE6e+92wKM8PpZIgNkxhUvbjntdh4VSuK
cMUrbjhODGOKEn+WRNzirqkaymnNhWfx+MK3jbbDjElC8oxz2K6tBm5V+LDf5Rkp
6wpXboHauyNsGpiP/DHfepFtKmXwALO5W2nH/4WuuJ9iwyG9wtyRPaqF+Q3+6xPs
k7jlr7cSLPtYUSKqJMY/qgAsTKLQaUCxvC99u6j0xqHNDEfp85GSPMUeesxXdXID
G57yY/hLxWiGrIun/yLVv+EsVYHQXElNyyd13e5fopFdXrFv3uyqV5gamW1ImTYW
Jb1XQRYEycLHqun6ch026utpSr8Ab00E4VLtBdUxVAxljYd02gu+jG5yXJ1rON1l
R+tpY7XwTSJ9jlIadmgRNkyhRLGfdFLBvafQaaMI3czbwyZVWdcnM/vosPEcDykt
Mq0l4yb1DoU7QC1uffwdHPlJ6cLVc81UrbsXI9e8UZW7CYMS/gdPRfqRKzXNctHP
4JuMDQuo3/14VehC2r7Exd0cRIvD/5K+wxlSxeT7CvLQTsRJcRRS0VNBmkdv44xH
6QPtU9QmiWfUqon8gQEgueGJXqd+Lusm4AKrw2OFohN8Lz8ftSzsTF1J96E/TbZY
XN2LatkJMULDNB48DZscieK+7fky089du1/+L8CpBKSyZU8kaP+sRQ26qbmvM9EU
3p8WtGRpHwtRsRq398aRVcFm32p2750XctteP3AI79j5h2D9qga9HMK7vHX/lNwc
wQa1g5kZRm8VL/mealiPW6SgbfePn88hhY3CgfmR4y1UY/lxcCX+x0PYk2G0//Nn
36yFV+x+sSOBfc5dRBBIuqnRYkuYGahhRQZqEcFrbLWGMs83XYlIUhetYv/EexrA
iBXGCwx8GmNAOLNm10J2pUup2P88g4xhoKjv1PVSZD64f228j1lVb3ZHFOccT/cd
+R/YDo1ZR8vZSre7GK8mH0aEUZ+aGNm0vFHKA2wPadLZ+MnOFGwm/kDPBN/3nsZO
/tcgZpbA7bp3lgTsivETu1DsrooIQkJLZNNocY1/7SVvcOBXXXKKKZFokiUSv44k
9YDfIeE8hwv0TziHE0HIgJmTMOi2tjeEqcMZqCspXbHz4/R9ajCSalR3VwTrRGwI
zyklo0CectbThW33ZKq8LUYjh6gDUJ9lwsrRYW46IfD0O86nxcx/z566E0JQnaoj
yK+pCBFO9tK+DJl5I8VPSG3Nb7FuFJ6QPX69FZx6MXTopSXsG5ABfKPAmSscHLO+
mqnjHu7QR+hcs/p2qprt7iLsQkNorVI8vm9tbPbD3b4eJR7tSpJsICGI0a1ysGf4
68no7K6PfMTgSYm+5jpItle4sj81CLR5CvC2ljZvalO0sfBpUxDtGhr6/z155qoG
o+QxqajAzuk8jLAj2nOUND45rf+LD3UraaEo1Fp7qXhLw7ND8861cpK4L7B5P+Az
YRTywPOyWx1VQa1na+tF1m85FaAhvV4Blff78cLPg+4vQK+KZBqdW5b347tDdQkf
ZuszCKjniOQItndb3/zK6Q1EbyESeYEBMAuBWOEWQ/Wnl3UALRXdtZKBSRmD7FbM
V4CsZClWRi3tiMAiwulh5NDwQP77vlVT/2imRxGNRP103gMMASaeaeOC8UZUx2M4
fOgvGAUCAvjqKYQUZxk66rSaoOCLbV92i5a6Sgf/FH4deYmmKSvXorBAWIkLRtc0
vPECpqR/8z9EZ90N/ke0o2G7xqiDatWFITde3IVzXk/iGoIh+RxuCfV2bP+o6Iwe
sveWzjL5g4Mivk9x+Qf6xfwd6JWYj6lNDj0RNHlYkbsp5yEy5QF28+ehaLbjcehA
htkcXpkbgmjLHcy5bSouDTy0W4ELq8a8hJ1el9hCWweeYcXqHgJcQlmBh0X7LLGz
LDBWwiWflIzR90uLk/uKXU4g78NlT9sPXhbGQK0GtEJi3BGlk4OBB4BIQrYBHbn9
O92gRKLXMkTwsRslQmsrjCn9i9nxrVDCMHUllQrcxvpRV1g9j6TchkS5tMPrC8By
Sda1yy6w8vMmNIydId0zlV7hPei6o61C1PwIJKC5S5IPN4ESkrldyxomQJTS8LRc
FsbWUhiRh5WBzY57CS+6w3ul8Kp9SmM0hXQUV9gFzuC5wvVDwzKg1kU2tAqpiVMK
8B1oT97QA05FK6pA6eFJQ9oAuFM+kVNKm7logfTaV8P5YYRcwmUrEh6ACd2dh/o5
Jox9vvwA2w9XXkFLeZtpyAtL5RnHL4TPECjJLtiLBL24PP147IhBE5eSdO6XzMQY
6+iC1l4CkwmGZp24pstUIwCqQojPHrw4vurwzp1WZYS7mXz57GR8oSS+1HJzdJDi
dww+cNRqveRVi7Ac6vBooB/OtOJcdpzPzC8GWGolM7ux9xqZ8tq6Kjy35hbolG6B
Vp7i2ky7BYn4l1eefbQ9TkXUH2PJzgLzKM9Iqkg51PcgbbSSxOVdqflAFgITCGrU
3fni8sIeKmtMqB7Rzph+tlsu2hiRKBIdsSBPe4bPXubesBvWOLAeOe1DWwuZ2FAD
ZSz1wrR7ox4YbJnA7yJXWVJPo/RXbHr113FEliAUm9wmbrnzznA+qaT6/ZNdtMmq
ON8jTSfp2sWf4J5fRSgTB3UhVhJH7qbZBOny7zQrIAuOTy4rOwoPnGtxmv3mNSok
cr+YhC9kFqLtmvjTRp8dN9TB/2ldXS431vdUAgSii11l1qqozuyH2tMN5ZEPfrs2
k4L4xHChr2QmUXHr+ij39oeE6u1PglkEAHJTmLJ0i1ON039MIILtFPuYQf68SsKb
++5hnzdg4a17z7acKVpNv5NYXGLs9rTLHxvLjomXYccxPZbgSRD9/GWD8+DFaioB
0XQ40tRZwwPqvHsMBJlKHu1cuRvHC73sTyD99QzjeZDiwUq+U5EubtZ4qEPZzfmi
sPKmECcGlnQKbcKCByIVAgi8EMgXzGJw5Hap3mNyV6OlWA9/2gZko7zJqElqi1Qt
010fRQgkuOghcMM2/Qz9/zGX4CInNA7rrMMjx50S5+oohaRYYpCaTTIifrq04b7v
rh06yzV7cXUJ3XKJgCwYPhDB3+B4UftHuBPctn7QeNy5b4kL6hp9LNatpaM+kQep
ffpvJvDQAPSbyMt01Fxq1QlYVdJpRGZKA5qMVs4PpxXOE2gJ6MAEqnAys29sciuA
0UO2XyAnE6OlaKA1VrbLTTdTz9c41IVC9t6tTirl0L9tHxkXTJEdXSkmk2fwxH0R
7XmfaQKmiBu5nKuW4tOHaAiwf9qbcVoQDLKUtUGbqXHvmq5QXY83zE+xUcH7Mnv8
Rr8bANAXd4Phfyks8Q0fNPWcOf8RDOT62VNgmxvlDDnPYyGxXtLtj7x7pEgBsXlF
+dxLM+IiHMkuj4rowbYhiIRixwTuFIUWgV1BpttjBrXFooVs2F5VImGx47iWuQ1I
BkEd3yVWMeiXS0Pe0jGmwKs3nmH04O9YAAkIzs2S05Ew3yxsBZJo5BxFNFa97KGP
C+ibyf0DB4v6ITyIZB3wY5rha/eoNfzRi0tymyBv5ktasP5tWwQmU7q0jqLUBKX8
8ieZnV8aeHVtHdOF7q4noVVnkUNOBFyfuJbIKI6b+PWAaJ+quLPSBcljLp+VQ0lY
3xTATTxZ49pgUt6fkNbdkVyYt9NIr0xk3htMYgBHY+c/ynMviQwJGHsaLL9hgqgx
5N6BZMfiad+MHeuYtMf3y9inBm2yFoSYa0Es/WiHoV/fJnaHZZVN5Lig13MVH7JP
RXNHkWqJFaSxKuVY7279RTISgBS7JRsD205/aRRYyCuXoRmv9Ug8g8CXkOm6gCdt
XhGwBMXxDTz1jKbahTN28foI65xrvgz2tS5XhxUfKCiDy6AS/1LuwSXV1itU4Fue
A8QSEDsQbK6JqRfoCRECGWdED1478jOrK9S810c74Hs7rwujzRlX39w/8TO4+ZLN
4dE0QiUXZyhQ59uGmeq8EvOIwnVXHJnLfCbwfqzazF8CcXaEwNkj1/+Zwq30V+k1
pZvL7NnCgWhOrstwGBPQpJAmnGES7uLeFWIRYdVgDGj8yf3ep6IH/6E/X7mxOCVe
zVoTlFDjWrb819wy6n1mwsJt6KjsuJdKdvjpmzJJ8Xumi4TvJ/F7ULRGWwVqjwj7
frseWl23/Mp9Vx4L/Dv2JCnA1xBms5iBJCZj6HAkDlGp7YBjAgAvR0WOqW/Hhu6s
MmTDoXmkxu5z1O24019w3iA4tdW+g+Y7Eax0HDP4NFbo9dH4NV8RoCGN3Xfp9n4d
Trmzh7zcYV2nLp7bIH6iPY7mg6IG4uQdOAPUhlysWuzLhG17NAxrdK8y6S65/n0u
7HW7+4osUmIVS7MoEjqBOGzyjKsui6CljZ9NL0aNtfNIgC9hPF4CyfuVUkkL76bn
G7eoMVe7zxxDy2B7aDH81aL0IuIvzZG6Q5+P8odNGmEB9Ycy1xYGIOQO+16U1lBq
b9Dg2RWUEkZOIoPP1D61KhZZg+fuAYsuau+TZ78Xi2njg4rNdDzeFI9oStSWvwJj
1NYIn7n/DfnWdmEuOVMX7VrUJ35zlFkF9tDZMS9wb2qOI/v2oXbq9isYtdLvXT/U
jjewx+xsTryv7Gxzu4T4ESFb03mgk4EyU5+HUxFnwBaMch4/JeP7zh+lpZCUVsmg
6u19VFH66gwgoOE6R+xSEaJVDgS/5ArAfNTOyfWKjP+KX1KOed9LYGKUjmSdM3XJ
b0SqKTCy8SVlYCIZZubbmuhj801T7/REu7TXvvGuXxjBoSv8bHUfXctcgk5oDJuc
VV+N+2jPpJmypu9CbL2zjCU56jNzNU3MykK3Htyn0J/qEJzj3e6fAtILfexA29jA
F5x/JQ8/cT6w0DZ3Xr0OU1VhfwAATANfNhJZq0WG6ddLCZ9rjokMZ+k4clJgEJXO
YQywJt+1shnVhcV1CocnIPXje4rqrsG6LhKChxb61SfzA85PwH4wRXvYChaugpsz
wL6t+nvnm7wXQqvnoaj/kPBqZ7Z1Kb+5DqivaJZW7sWQhXS90E+f4v7UgyvrgE7M
/fTZIQCLdIkC88kzWdg6mqtsecXmbNfZqmG9rILE4cmHsaHnH6sMuMMap2v/3Z1q
ZASh88SW7hjCYCveu8Zq46XV6F6wdjBzuTx7QET5rdb6kDGfYu9pWVucqxDmEGgl
VeEKoyrOs2/yUv2GendGjA1iZfNorHtVnrAz1eSOpiq5VH7NAkrLno6M5ZUT5xpe
XxfsX9aVum0j0OSix4fMgfsTWsia8bGcIQY87jPQPwoTzlqB6NUVn2wpzQyAonJY
1kKO8DKScadz8S47c4JWvGu78Vj8l/raFuZpPmzHqXpNS+zu2hwnFVzVNxlJZPr4
F/aEr02LAcugimsBi7CbZ7DRZdHr35tU9b7PlawdEr6rQFr7xckbys89Dyu9pCsO
lPTv9esTEjQlZhpR6LUBdlG1Md5PqeNy26VNHt60AtU8KkP8etQhJ510Ec7Gl8z5
/xefEBlY3qwrdfAdut/C8ZdmU+Ee1eHrgvVUt8hb2I1DFPSmW2gPRSwWowS5Rq+C
+ZMNmcNgEFVv/Dp9MQqPVNA8GoaKa4R/a9XLHGAnsicPgD5PSERMR6sya/xA3deh
2XYmPjmt0A7m5JFoAiK6PUj+qc9Ewu4XZsnj8wJN+hXePG7BXp5WNvE6IoPTaZD3
NIMVQMt/KMNSm01YapXWgGQ+Aub93OpQvE+gkS6G6S0aargPnRiHqmFY6CdZSVUl
ZI6DaJUuiaIlnH6OrdbHH5jRbzOHWc3LnSMKhmm2Nz42q8/Tf/DG2vaBTc7mW6G6
K2aTnt/p8DODBRwekyHR2Zm35VhwkoXzyGCPtiHDnMQKN6OqOjZE+3YbrXHnn4OI
AXLtQsjXSHFk9DgOI7T1QBLo32yTw+ZJMsdx6NGAq1xq6ENmEGqYcZ8UC9XBMR1G
Zau9kKKDwCK92BPibiNxb8nuPKR1pCsz37pO9gkbwXHN5PcwETp3hMH1krO6iLiX
IRFa0wdV77GwyR31Xe49HSUppn80fp03wjUZ1SZayqPRVvNkxj8mVZIoaqrKNySb
590qgtiSOrrAb8aRM0vRknLG/SNO+v3OkbC04dFbqeNUn7tkwLJGWAS/xl33Nlbg
tNkoBDnzemQHHfoZgfVWgwjoVntsfc9szFN3hc7htVNghTrR+IkW9Kjn958PmOns
FOob16wqnURaf9rbTN99Vwc3lIs9aq4/ldk//T/WJaK2jHKcMstRb5cwRsjjnvs0
/N2GBoSMG2xlEQccM140jF92qvHOkMLxZH0tdTRhtqgEAaPq43ggpJyHyQDSR1at
+rRoQqyReAyPmwgh3fIW1gAcU4wY6cV9R/ovYkuCjtBS40ogmiYWBWfZ+s8BkVUg
4fv0QViI0m10HxPiMZKRYZp38wYixxwzuOXZjuT/gBXg21FBq8F21lnSsNyt54ae
V6FoqXMhOD/IHSd824TbkzZEhjQ29kocYXwTOu03c5bVQfhbL+ofL4mJBpJ9624p
2LutW42hTCL6/nC4Ih+dzb20rLcdGy1Rpuc/vtE19pAhVznHbLeJywhBlrFch6xu
jymKGOUoEGgtPIRnipT0tXB7ON+kLc82qH32rUFifNq9tQn4L0D9uv2cHo9gafq5
hWJJjOjuIkE3U/neqZSdjm6bdm2q5P3o+UrdEN8zghM+jwXO+uzDMjm7xcdS5wUj
Q8aE4L9/evyNA4DIPWBcal1kvS+LuCZh5ob4qNEfMByPnEw5oOV1hwcrfX8zFljJ
OZjbeqoWqDfagM61mC0BgUZEZpMUTUTSTG5x2dIbFzf4XZu8pxcba2UYCU3KV1GP
3uUFsom3UTYnCZddMGNnfgSsuATjrGdlI41VuChtkmkLSik8NzvJKR5OtvKZ1jtR
D3TULl6GvroXKE8LVf+Eu4gAAnvMUfeh7tjPIiGmIu4OSasp+Va4NwFbmUUfPFfk
DXi5DCEL64o0mmJLK/0nBelBiFTO00kqCqEZ5DxjXbhRwq6pKsEHSrLHEZ3Bt4mF
JFeObHLK8fw061VeernapgVHp4owFc0yvthV5FH+WYjWaSGrH761Z09jOaviUayh
TpLH0iSoP1tSkjSQxdo/fTFBbWXMPhhOjY56t/1P0tyJsbHdYEQJGtCD3uqgo3r5
hPn9iU4yjwc99xVypia9EHLVnNEElxYlhcYkhEM5qxdbUHQpOXkdlIcoEnihQLGC
AYHPV0kIOFemlbcbkT4ZAR95LmFNNzcheqaQfaFiY8xBBa9Z5Q0/bRYn3fz2aNDb
ph/MO8aaeUe8XEq5ysFaXFBRSGkWzFoEwuVAYrk/iUudmkR6bCRniCNPVcDX6tp1
mzrkajjgpJsm6dd06smcU4k2BaihMkjATUj2LF55cnwnBzRYa4yVAibsJb1nBxSA
aVhCuuc3cWbWfKWRz9naWmpuvk5iuE5/TrAz4S5jtoJ3vIPmJzM7O1SKC1oT4G1G
eav98QYJAzVMfdUZXElgfiR/ebUZeIkhF5lVfrH9zgeP/IwX/N5bROpjOw5PBF+c
YOl1E4OMQRrIhNyTuqKB/hfFTTGYMQ1W1apt9vwea+U1mvMrDXFu9FJ8r8xSFjhb
77f93mQRIPagvY7S4Dj5CxlFyDMZohogIS+NqjB/qfcUZEDuSykK2Q054XG+Qx7j
73UHjzLCPzDq98YDKkNyPeh4l7aCFDk739HnPVnJvUSdoXNrCrOdUVx47qfV5DyF
H4ePUGUA8fdwi9VXlrL55y5WnS14OOBFMflULgkg38wwFb74U2CZnKweGMm0ryew
d4NgAjrd9ItEdJECNgp49pL99OFwayroSYZ0egB3IRQVXlNdcocIv2CUpkbdpq9a
4I+T6bh0Ohmqy5lUU8U+xKaPlmrFF84a3gIF42vMUX6kK4Kk9sfC7fiEk4iGXUIR
fMt5Bnbmelyj6oZKw1TZE7ZoaaSU/oVud1qLsFYP3RiwGmaho4/wG1+dHwznaZRE
atPwUelmdXodWNT7dVTOVvRAL4+zsT5LYS7/MhjS3gYw9oqvoO3HnAt2XoY70/Ov
arm68jZvl6aQxTfYsnNlLXqPClBg+NC/8BR5QYRNDxiTImWkVWCkXIhX02zFQPQB
5PCXwVyTw46Wl7Hrr8p+/hy3S5Ok0lj8F7EKnMB6F9rwh9rygZ6VO2yO5cK3Q58H
Chqu1ucOLacez45WO1RJpKKxmn67csvTztMy5lx7cyxDn13tplwm9SlRDJ7ZKIwj
qF+bcyypHhGsEM5uCaCRik19rf7n1KrLOvqWe7jGWur39X0yddCPVWHn84s4g84C
2hHT/H5kt6yr35QlHkV6KeZxMN/+Y2FY5i7juV2sLmYIZqCXrShXX3nBgDKQY/39
s8JGiQWUeUbni6+xGxJM91mP7smz7hmW4Gy55PY97BpLwLpAK7zGESYfh3HMnQZK
CJNG8v80DyItShGj+fxZv7ttjdTy7WSpCvPRBD9CrW44TsxPX/dPcPN7A1W/wB/J
8S2+rG8ZhivPk5J+ZQmYnH796DG7ltprTsQYZvopAOSIYzFk47zbEJWQpbICVMw+
036DRXpEgX6aSii9EaESir385LldKEvbbIB+Rptvl72KJ8dDiQAkmwwE6nBOnNP4
cKYXwNopbcMMgTMvgqNoWAyyr3gzDlXf62qyzdk37ZVdSVN2WwNPmmH2wGtg1nX/
tdaQauwzHJVaxpFHEWMLKbzcptKvuEw8hwiJE/QSFdxLiJYbEFhu29L4V2OH8w3j
X2bQ5QBWhStis7J18g6kzLnVlVU4LZNBKxKvnCT/pWis5Xa0z8AwV4n+URgDc3DW
Sr+pvrGyx1BTlxWho6zBEqYcfbhR6q/gAlc9yQ3B0eBweavFEuIB3p1H5Od8cXqW
C7rBadFbbwd+xnMMBfKm8v+g4d/dyFAO8AMCTtHldmFERsi+Av+7l+8NF7prSfPc
1IP2FF/pzz+YPGx5T2USiBd83N5Us78BfkBfSbG+tvBYGOL/gMZFNYu5L0d1Ilwg
wp5sHC5FqXnHzFuKPWFB40wWbV5YrPycpDQ5pCzpKtOPLi7WiDxS7e4GBGKSQ73F
Bl3dLrSJv0j5s95JnuKK1yU8Zfw9XPfiWsZZlLlXpYHlRc+O3+j+jPB8om8oO/vC
gS+3jYtbTvsPTZVFd5+/uR2LscstuOanZnHQ7o+Km1rnAnsASVjF7S9YSqpyvnqN
JNlJqb8YLhXLzW6IAstPNjCgHgmMDjSUvvvA+WPIxeSXu9c5l+RkrAjm1QC4heOM
yq6QGAs00Ih/wqlfuLGC/OpCDdYAuMHVqkGWJEEbNNt5+zIKiBsJZPk08KXcSqqB
fVTbbNHswUswDz6W0KH3oIS4VOnanEthpx9buKyXx/1YRbsoQ6plBTgnZ0AmrmDy
2vdppgir0CEANsXxQwdz+GXGE1McNkSK5jDcrX677VZLGjHh5KUumJl20DsksZtB
4iUMQuM8HwtV53ePflBrfznymVbXKKM5ii5I8KH2ulTPR2Zhn/9pYCr4j2+vVKQq
PoE1u5gMRMyMXab+xFo/qSLWguamv20lm0zbe5ocBqqb+tfbLABsE3YsHspYCEyz
XuIKfXKxqO21amfFpCEamN8MEF8WQzv4RXJjxhVYR6PlwWyr+IwppWub14ys/sVu
c27xcxxSLRL3r7FgyPafW9OZxgpXRE2csUEYVja96mC8u3eztsAI44q+oAiDwvDd
EqqE7W3q3DWyLuGl07HJF/ITlocim3PoN4rKTdPoGlVQO+iQTXyje5hmf5KvxIMF
p80hK0cYnMMhUm8Lx7cQICrL0AoUyBI3QQs2h0kauS13msT5PHeutzdnsdUr8Z31
C9Xf5jrTdEJALYL9jdvfDwkRCY0gORnLLUSpUygn1BPdv47KtqP3NrMXl7I4Zojn
ETq3dpbn32S8NkyB3vkvuO1NQmWTlUv7uWHFmBhdYon0PBLK174UQzPlXevcLa3X
kJYkFjfGZ+feprXDXvbB+1p3OiUaqn0Czf/JNQk0zIw9v5URDYGd69nlEOizu+D0
+2wQt3Uy7Qie6Co4S+JXHsbZN58VeRdvDdTqDXccr3R7Hkk6WPt1Va/+aZGLaLcW
W5F3VkaLOXi0LfAZM9AMvOS5ArGIdhey0DWv1TFo4VSTKqXTDmONpijYa7t695Vs
kAW91SoeQAa0ZU3tja5W8ZYIDlYwJ/l+sUIYkQPIi8Y7SmD805aH4O76qd9IZ5j2
KsEDaYn9PJCRNeaMphX1JWpP0fjaHGhDB1w3ALlWxs2p+U9ntB4Va0eKawwvdFl5
4Ie7rTyFqAb9ItlkZCP5I2gl6ptk0G1ieewv5O8BtubgL3P8tM5skDkx2weB8nHF
e/p0IffIrHSCLj7Hvgm1MKdMvmsE3gok5gZxE6O2OfxyLwhYAjTSPM5tj2nOo+Ml
mxOA3GHGajpXEH6sws4xb80y67M3+92x5MRLTz94hxv9nHsm9CqZ8BLvshJ9zKUq
mdc1XnA/FqVcE4ePmkfWgfK0vPOaK9KPABmRhTI1z+CqsffNbX0Q8/fUdKXawwpv
6fabSViWnQGDp0CVl2n3fvJ3QdWIKwrUpwIp7eCGuFJKuRYDpSRyzp0UB413JF0r
IiNnJbRMOOFgQglnOno7xAZtEfFKk7i/HB2r2k9Z88i1iwb5Qgjpp1Jnnpnjw61K
Eg+la7Z36/biKWcQgcd3+UZasiHT7cp1XFHL1CR39fOhq4RL1A4X2h1q43kHFDyr
xXhLD+UKzSE4AzzlCHGbALfqObI9vrltfgK/ntP68Ci1gI6uxMchC3bRTodIB/dk
l96mk2NwuRoR+1984hIXI4ncDF7el1iocALgNsvC10WKEAe3fnxXrTD93Z9dCnpJ
dXGRXseIyi9d03znxP3elrQtLmwvMv0Ekm+F29caGkRbEr/uHh+ZBj51hbhGWWC+
QNQANvpxmo/SyQ9r0v90q4Am8yH5x52R5zV4Ns/T2gMU4AXr13XWTpZeqt7f1zyT
mKyZPzMvBOaATd7ik8ewjm2jX8OR6TtHPqesCDaYjHJv3NE3FiT2NuQtm3kRX8dy
LS/m2jF145iW0UbOmv+UhRsCvh8hVy7aw5BmVQjsgOwcgVhmQHDuBBc/w1ArpmLU
d3sqjvdK3ljgkXpnTGYW13QtuJfhJW8F38RJ7z4r/mdJsIbJdkVeR9clo2RGAYRT
rw49K9POZbTu1fpJEVGXGAf01vj+mfGgLbKAhFljYc4J6e5jIGcBkFmVkYrGzXir
XgJyseZdfjrFYzd2yC3oOYHaER9G7YlTy5i+T1jxpSKfeL3Xtcmkf6m5jBdD7di1
t+9LAfYpsPbgzQaTfQOSLeex4aUNmS4BSTL6B1zh+7Nx+2S3yod+wvSly3Fzy1TN
Sz1neVYEv0nbhdMqm+qAOvBIDd7b0/UTEfk7g4jfDCMtk+wERhp6A4t0fQsEMu4S
K/FupqYj2MQ9LRCNzKtXD+UTWDpTqMaCL8WPKaXx2G95bekX3aKAhrcrO68ZbJku
SgXzIklxVWkIV7IsLelaT9WkZF/6RYScNFds34Pdm8BuOu05mklMdCSSBYp8eAiD
73kuBlfA6leyeGiRkcPPYCeXRZtZTBgCCLeecD8pB09HHOHy2K/yHAl5CrOK3iwz
+PTyRtSxjnqGvQHpZIjxV5QsaklVa29ogzbjDgUyYSkafTWY69hM4GgX4YboXEKb
FUKkP5t7IkowZSB57VLHePeEi5uBb+dKeB8z9N1Oi0N5nFO/KbVCHXMx1914jfpy
2njCPMqtR1m4AvQa7HxAh434qQhQ9aLFOX3x7dwivWsUpwTbztpK6fUpV0CnB9rs
rwwgu4XvB8vbOW9zr74CUfJaMsOZD+mir/+LUwhRgZbp8ag7G8t21qoCNX15y/Hj
0NZGiGe0sLgZrVwn4L9PFxQkDb5kULSAH2llap/8BjSUh5WvVCBIlnQ+DLqpxch7
aVzSCZ4QYoqfx8Sr0fqbyVlIooAP6EBosplyQ9og1xEYoWcHP9tKSZRAMbJ6hca3
9JbvHgjhvkuDnb9om3wusnmq/1Alfp8qpcvc6CZ2WTeD1oG56Uy5d0gXrDWMVeUh
Fp1rBdtwWr1AlxOhICp5666jvTvEwBssd6oZ1kv3Sua9FGwJnwqGAbqJ32ZyWEBB
M2oQDj+MK+NPhAXV3RZapkWcBUmxSDVg0cyI0HCwTro5SZ7MVl1bWFp1qCsfc5dJ
7UFHjP0zTKmK+qHxxO3mdqYA7KrxEMbk89L0Kn+ZXlWTB9j7mPA02e02EczTRPRa
u6+Ao9gI4T/Bqa3rCDmyJipPIbIgpyU7kCD9M4/nBZnYRWPYBrnnXLYpC+RNj/zd
04Ke3kAAy7GyuS4pKhjIBDJFTiXpb7AkHusax2ltfLOOvc5VlTcULVASZBYEloZ3
5MflbxD8fqoU1aCXbVatHb+s82N1ipcU6Mv2yDadGp7c/FOYn6klaxYexXQgDqG5
9LZ2RK1MjeENjaVL10dqHm7Fxre4ub/ZhW6zkO+k7mLTDMQAgtsViFyK0eib2TKI
eLJY5/5lxeNuaQ1/Eg77lzqA/g3JcfoeShZFlJslpFjtEfn3baZ8v253QUADEVHi
Q5h3Zi4T52XPL0ce6BAehPZu45nEm26je9JITUFkMjDDwjgKON3+6IcDBBKOARIC
GMMNBu1pQh7GFsqE6c3l+yTQ69Ked4f2pISlePM/o6Vkgkfl12i4tQ3Tis5IZEb1
DzfiI+2W8FdzhE78cL1g/CNsBPqMFs/4c1tbGllwQsYBztl1Si14nSF4JpXMKXLG
hOHIFY+4/iyw6T8rpZ9CYBGW9REzyNor1O0s2bnfwk7fB2i9jNdjlbnwAqvIRmIU
DWlqhVNsj4DAdcJJQ9lnZRdaqTjReBw2Py1juT2CbytBL1/dSXTRCUJzZXF9dzDo
LtwHdOjtXNbrKMNxEU2hQudjfJpK0lW6ZRdxvfzM6faOodDhfdkzpAmvejcbrqxP
rrrrgvUIWUx+VCf+nnnCsB4X23S7wqTF858kkWSuT7p5aD3dF0SYENK3lvP3GY7p
U6LFIm6jukre6NOFvf/O6ZT5tyZalbkpgoXvJD501QIy0E4YR197pMcTOutdY2IX
L9/M3GwzU0Atcc+ZOTEeezWNiDK2jC4+mAirnGQ0TleaAkgq45gtht5TFhJewzId
myb5X7G/m1KEvtISxf5f6fjZKyZNc4550SfNZBpqSAR3jd7RwQH7R1cYfYFyCcnx
HcyarybjWi32695WI39GsNrwh/aaqzuILdZkpI5KVqWX0N/OE4jDsmjaLAFju6G2
+uPx5LQdQ9j1mTSv6fDVeC6joCClaQrIyDWR0WUX9F7xpJpJKkhLHdTpSpkmlxBk
vdwaJQRsUmgfix2TsIECTL4ajXBtdCcElOzhkrODVMtQXVCYe0MwSfmz0fZRPt3F
hCPV0f19WyHwWnOXVYtAcs6iqY9zIf3V65tG3WN+FQx/Pu1XrRoNigImeTzGRfiu
J9YO3RjPAEoRYv8E545lDNVSUiDxMFgaDW1G7nGqrdcfNG4pEZmcn0SxEqztlJGE
q3Aw8n2afP05pAGe9ydW0kO2rB6cO4hl15EocHMq5GNy23MHd7ltoJ1/SObgrtmO
7JgwxK8nbKWae80+3/BfOghfDgiRCSIr+vheGex+rF2+rYovJjJt/X9iHidZRO16
10yRNNu0l+JFR6lTDNqd/rGN/H0bU5+UVrYVN4HZQO8KQiMQ/T/Xv7LPbVWqqrPh
xXEsLDrP40fe/GrY8j9CBMvkwfHA1r4yBh19ksLIXs+nMwuGPxU9BC6GQgrOPnwR
k6lUrmInPehZ/rSAMVxT3Fe2OrlmkazqfZUfQP72CJif3szNGVD5z9V4UMSQXIea
M3gRy524QHZgYoUgnGtICYSQWsTMqPNI6yQkZqEWocBsCuCyDlgHCvLON+XgSNS/
MgvGIHvwdQU3KcqOaDrQFp2WbikH7libWnI9dStcOkapyW9Bn+lLsp0Vbt+ZlHMs
oeqr5jm5/1xQE29gBeFNnmiEzID7E4JE9gfW2UhoytQVtssWGgvFAcImTtr3Tkjl
WiKNFBj1QeN6AnAV/DMaRAs5BWpW7xsjCYcaR5/XAYwfxSPrVfHzwwLpMELqQAyF
Qeyj+29WqTE/TNO8MBJNfcbdNKwxfNMr3/cupGxDvRgjUeBOY3jQtm10/vDBmO0s
xMUEh7SA68hToKBY0rpNjpugcYdmaBcMDd51iWDeFinFIak0UpEOUvQOvhGvw4xO
sne/ddoT5J2CpXoZgCxZEelVsVTRCt+GWTfri6EZiwXkNDaXYMRIn2NyG9akvwhR
3cUncNhHwCeuL2cgI7cb2cPO/zory/zWOxcX6MWGNNv38AK4CdE4NT5SDteFZdbh
JOkZTcyhGnty0kLoMkuiiU/yHbD7jUVg+4hP2I6qu22ay7UOtSBjdFKrdM6i0gem
bS9Jz68FWvdLIAffTZIoTAIeXJJWTkEA2Z4xM6MpU+E7kN1z0+beQhK7CCVcxLao
DG86D/BwqzAUOr7vNvwjKbiYurFLoLw+/Yl2CKWQvO13tSV0X4pO1Ji5i9Q6HVCk
zAtLJeOYvVzOect+T5FYniO1EleYLVH094HXEPFXu2tf4jiw8DTxRwmwpaSX2AGZ
Lxco8p4OGvpruoXAUsdNJ+NaTXLFVOJ/e00PozDfJi5n9i5cBWVx9o4lm8c/aGy0
0khUxlUBgbMEiETZh6WNVAn6sA//mdk2yf0Pr4aGqhryIE9D/PGMRCeGSC5NG4/1
3pzZt1H5W/8Irm9IHqX6/KKYfrvNoY15NeHRRlJNmQOGsUGzBPGdcZ2AI7LzvNMJ
m9kVNdbS+D4mP0o/4T5aPFxCDx6xlUG3i7P5nEkWkCLDcuksalNqUW0r/gJs8XRc
Xnwmq+BhwFPHIV7Ye3dtEQ1sXpZYRQCimeRXoDlEgAu3Pw3sHrFGAwj3DaV94YDO
hO728stCAYvnsrQ+IB5tixep641TaUkT7AIDz5wNbDqj9lGI3iEvBv0G1B+llfPe
nps2Lru5YmbUKi1qUWcP9UxgHsBVyRWUi8ZXsgly25xp16eWERTU50wfkr8mwgz1
/+Cw9MuUialxNc1ei8uvNxTAVOyMJrQafkUE0BaelffhnRzEQWVVHWxEYJJuvGyi
ndI8ng+8d/7s8vB2IVz+R82h33rTin9+DT/0nKOYgi6vbVFPdu0edAgyGGrf1WDm
GGxLYzQd3vK0xrr3K7R6qalTpciaweT7zx57X9vJvpyyRfGrJFSFyc3DMUYhlJk8
sr8uDninHTlDEQ+d6vsHGo4Ik9pK6ON5EmA6iuacnI8r5VtwZefrpUdPQLG5Z6sg
ssBpOnmiKQ9+tw4qXq4uy4Zh/Qs75tpzuz9APXVQL3jDqtibAJO7ssFiHYIpTXgh
I8gczUFuRu8KP/fH4BnKKYQuQ4i1S8n8X9PkMBiB9Jki+N3S0LbMYT3yvYwyTfSn
5aV2CXln/8qriS0cHuoUn3lrZw8pStUNtDVH77f0GGsYveUFZTfT5mogmz1R2aP2
2XmNauQfq8LNAxjWTPDlVEkZq4IXpzZxCIwzVetIK3sIyXxYCP0qBquQ80X1sCWc
uOAL8ALbshjFKMldCe+dzaJ3DwEJpIlmY30bPXQJeV/SIRYSyYK4n977WCudA+pz
fxzwcs34zsYwF+e1RZIupHgqpDJTty3AlIQGdlx7D3sgXJIuv9zjAGZx4+xD8u8j
ley5caQ3ApeBrBYBTFpiG/Tefd8J9Yz+VPD3OxFj61Dhn7QHhTfZnRHRhQ4Tvzar
J946oJrm29/rwnsqHTdAFHcoPyjAqCK1JEK+nc+F+gSOdk24i1eyvu8BLs1IEI74
I6LGg+B1fVEmx8iKisY2PjOpIHLfIaQt9hti3vIEwyd5uZ5Hvo0lAsfPypSB5Mun
Vi8sH4buEg6Iakhykl2it3106A0FVgiKyyH1Nv2cq9xn5mzNrgdAKx9PUjyFd+fY
MnVJMBeVWaZmOdXZq3JaCfDotzket6dhB5rwlsr5RqjMqnxZvn6eOKLajdK7jB19
NySpKEyNwWnvfXTovZPAZGXuRwCQzFogs4BEdTgkS3qSb+mlIl6Ba8fJ8j0qsnM5
YndUAhXlwQKiSld5akFTYIvIt1cnPNjETndJSDPyOgvE+C1/f3EW+9elyRrNdpSr
HHunelLWqFP17UXdqhTcWSkuJHZcPutWlMaURrIWpfH55yXpaG7nD5XxaII40NEI
a2IHnC0/SmqaUgJJCzKP+J6UNAM1oLL8LvE/MzJK4kcRcUkWm1bXGSdw+NXAMRCd
ykWdsxAq7ErbZ1ujfNKR4eVnRyhR2joy0CeAXSJk+rnjJD3cODBIEKYFFA/N/C+C
oRnZMKGHSNLmpNdrDuiGo7anW0aL4SlipLQ3uRz1Yyo8fxqCSezT2TD+QY3IzcNc
MkZ3tkKyiKhzPApBm8dXHQr9acwt11PHMIqzhdW+aMuAT5nzIj4X/Df1lf6lPco5
qa4JOxJVzYZ2pg5t0KNUfkX3o08MqK9tYjdGm6Y8MSdKpZ90RXIQE8sv1B1FLZfP
fpftMm+1EdEVhFclo2yWm3bBJIixJZ7Tt/rENp0opOp0njRnY+U7nJ+X7ylnebWG
HSo+qMAqNOC1s0TGaCsrHEOvHGU8G35yCY19xagoxGRISsLSer32TK/y6m3+21Me
cLNSI2kr0nUJzzWKsvOks+T/Fu47IR9XNXRn1MAOGAddoLCnLpCCmkxTFea0WRAz
a+Kq+W0xD/o6sDMVUlzX4eCP8K8ORM6JEcMRyoFBYOPh1bp2KfZXgtYHFjRwi2vM
y35bwRQqPfRnvGVb9ghCYqK9Cng9aruD4W1W9lvYcxqBqNrSGTZhYBK8I3qq0tIU
BAwczQ6uJlM1hKjRk7HR+unyq6jZ9jGkdYiD+mCFHfIgAkV3Ummji3jHHynqPIbr
0XgOl9KBw5Xq3EgIxQMXND89avMOa3mmLQBjyo9We6k9qUYWNbh9uMNlAYFms5hd
InypiWVPES/5Ca5NVevJeVpJcAhK5JgTXvKan4Ts4oUMT5G8VDfdH6RmaIEblwk3
zzUShDRlnb+4Sb1KcgQSaCBvVwqeyMzl0FMkxopyOcA0/RaTTEzE5vKelthveaS4
ajupvMHizETmp/BZWMQhOHdoX/8fxIQ+OB1R1zwa3ELkM/B192v3mQzyxJYZh41o
kCqN/oQ4Ay6z9hBwyUEFVCVrIMf+2uTI9z9+/4t69gLoKGO2h0GDPVHzS4iOiRc8
haSscAPsXA7aLbRELApkixCWaGlQOL+lP3/ClfELZPfrXhJAuvCT6bwvjrripfz2
qwWjfft9Kh403Jrd2i7xvNv8bTBC4ZPJe1fYZHTg2R3XK6xjpufc7LPOSc53Qu9X
YbDVwzirZ9fsMIfQ/MDNtzHmsbjVqrwhwjx7xMm2U7Ih6U7GSYIAc0ZN9V8rn/Dw
evHF/DpOHhLfVowqTB6/7rM70j2fGWc0DqK+S6b7cMQirnp/2gE+cPeEkksuvmyW
93Q+o1loVZo8VWbU4xdkYQ/kPzwTzDzOFEvPu7SLV1csbCjxWDjRrdburfx+qR7j
1nRuPCFopYCxK33rVfaIxtFJE1Fq0avx2p01VzCq43spb7iDjej7w5vja0qQlRBh
dYHgizJ1wiQVAQFbZ/6HBp3KBklmXw0Y1bW5DrnJbcIBEieFaI2S1w9J8FqgMP9F
Uvclg5O7Q6LOiJjfhuyWEXfrGyTOUo3jSyZykimny8Ab/cCRlkQfqsapRQWQk/G9
wnzEysxyMDnZJ1goQY1xZoK5NYtYy864dOCK9pnvWvOlX0HMNbgwemNHevfURPZq
+7ZJ+Dq3wsuVmXOE+ZntrnL1rO5ZK8RIv2RjBU79dPiYjquFQVi7XYH/pLwZ2l7x
m8KUd7tRUqHPjCLd7KsfLMJ8J3meoSrpM2KDaZqkI/+1UFqn3IVFkKrz1nS6qddY
5WO9DDn91DO859SeH1Hm/B2h8mlQkGZ4tvBkEH99koWSdsBQAJBXiZDDy3R6TQhp
YqpRVoAfDVWLFGz4MKpQnVVWLOQBKC1RnHGc5kHsHXtmIRFs8xYLPWqhaGRDt5HB
Adci87TRyIAW8aJ/TAhnEdpzQ5QtBSsNLc1RyKXJyMRP/PqfzxdFgoLuzeQAlOS6
FeswmA1oQsxC3+7G7Sol4eFNASZ/MLEscrowhAOrC0mTRLozIeNVqnEx0g8l2wUf
CAMcY4lhZFoGFoHBRrqo8FQ6hnvBP6myuc/8WpND0bq4ptmhvFyEAypTfo/WbWvA
TMy6sGZBm/9gRgs4Xv1zVVtDrpphuWnnNidfHxvQGwzeD6eXGCeDgymeGI1bkkUu
bq+BIquef4AqdOvazpnFh+vA+0xlwpkqqfRAxuM71F2ePVkmhc8/EUVSmQnEDo2d
vgMN5yvr0zAag15o6YYRgug6aNjSCe8QYG5tF6sCFabllSdv6yiYXe056f2KElQL
WKdIa/4S0ynRkHiyVEjtfGDKpgpdoQQoucBXtVroIlzqnt8i4CjoUnnhO/freJT4
1/1gwIQK4mugVJFxEq2I2mdqiqICe6FGeUDwnDQ05wNnoSlwG+jAddrfJpsDB585
yhFKfiHHfCMRBqCSV1bdlINcqMxDVlYVB/J10RPT/qj1gW8TR9GCcGMaciXS6ce/
xzufYNedtDuSLhh+3MScT0WOh1OOb/0b+uIKbGaiY2w09E/4cjF/Q1wMlYYkfCUN
i9qwd27h8lXaicYX3OVShlCGC9/KPxesazdNWkFm3nF6Fv4OS4njXtNRCngSE1A9
kFgHyjtrTTJOLI2MV9Ee0wYP3ubCUBAd49veRFfRMmwRmLZ5n09F7aM3VRzzqJIo
pfi1wfbjsxgUObL4IN7izQ3fVQ05ZnFfSSUUgnpDKFYQFacCEPvjQGCLorrCrVbJ
nsSdgZ2GO6bo8DYcx9XyKSS0GM/g/QI8hKGDX7NtScrLCH8EBOad2G7oxTPDOs29
3TNMwr53RcdVBChj0f1+UjIN5Lrou1d4Y2Z1a6O2DtrlpxhBMhQEyuugDQI7Is/s
Lh1LuLzkjA79Fy/omCYFAjzldzE1eZdbz+n2ydbhv9B6HUYfW/sS4p9SdwOvXSPL
fPYf/aUv89W/qLF0dc+bJz1tmWy2Sp2TxcLPqhL6cclXTVcoS1ScVDhp8RChU8uG
lss8Au0zawFR34L6wwhZM1c/VeqtBGcCqqlvXnB3fSaRrPj3+wHlQDV+9O8/UIM3
gPjNAaUOmPnFKoVCJ200Xh7e7JJZb/8Zlto984xaF7AT+P6syq5EewUEsxIlxZHZ
KmgQNBqtGGWIXxq/etdwiMjat1mKeWNF3IkmbZzuzbJYqg9bdrHnIF3rz4SAVshN
TzwSFNhvYAWTJDHyM8xXnz7oVc7Od/zoL5hlqQCxIbyBhibGV6sGqN9aSLsCVQIW
syu8Fqvb3g0xMb0M9lzz1jJewF59FdDPrKifSHtGQrpBxjagwvGtaX8IKFDDeCr5
8PKxnWptDtT2QkP1tkMyFdgi3tnyAZ9FBDIUHulyRbaXKMi82U1i3mMvmC+abh42
b0RL73l2CwOmAV5S9CxzbaS+9hMUyiStyDOZVzhCsaGR+biYL1nBqhHc+KNp+sld
Q+BpGUsH+xgw/grmFD1Y5gzyXUO0D+TwIrwE/8EhS8sMzaHGsrIQSTdbFzECnyL1
DkDoduaubI+kOssOyXREMXk/Ix2xZ6OG2HmTn5tGdxeqQqZEgCC/mCELs/Njd7Gd
O9c0Za/3yWhAEzEyrbFM3ZKCgx6SdOj6frJw0MoxZC9zgbkbrU4Pa6ejDJLL7F8y
yhzOc3NPpREUDvPXNLX9nQj6qs4CbkYa6htEck5IB5ptzE8DN8rSFbzEva3MbYio
B3Gz1AdToFkYatHpPGgqk3aqgxrva2384+kN19WOVp/fS+f0JWS2jhPR6Ykh97WH
Jf9ismIsEMxwj73rbqRFSadeCdK2lCkyVwvOeponxYXmsJkVb3b9qH3jUuiE6jq8
fbmI4j+0bW8TLanz4ZvqesdzPOeluu9fWY7sgJlfrIs1ggkme2XmVcKrTaC7fn2l
bCYbwrK7mqI65zM9xMRl3Y27i8r+fPf4bF51v4xEaYtztJjVWQ+6wkAAUuVM76Mc
gdxR5YMXb+WJVpriQOz/naADFO/fCqGwvHYSPhfVCtgjx69vvb7NdsdNeuWPIAaU
UFXOYVYeaapDzrb6eyay5AMC6nwk4B2JpMS5p6jacymgCZHWNW/FcgX8I+Vk7bBb
c9q/faKabk6lFa0NEWbptBmKpPv6uzManumRdnk11WeBgYAirg7f7GEL6JcqahBt
E2zGEQhy06hR1YgskF7X6Qwishno+ZmkFm2yvA4BizqRKsW/vZ063cnpPo8+C+ie
4YM9xdoT4wVRYv6cntDEDhW72aE1Us9z0JpQNJSy80ZvnYt9VpCZKnpH9szsKrF1
0CnzSFnUl/LLBHG04HQ7zui1CeAJddFBSHR5a+7cqDaXiR6/AqX74r4JQcyMNiPe
nExzQld04z4nJrFjwALvJ+Nlt220hAW8lFCJdtEHOezKv0VPdaVjLb6uFeXnvsT2
sZ97vlIFOV46ZO5Oy2YVnfKDYyNr84CtJKjcFyZMdauddAtUh1OhEcA5BirdSQl3
RPP9lnFuio1l/OU62na1uUqZXw3MxOY0nPP6VrJj/qYrYVvQPqYnX6VP+U+03+Q4
cO9CrDUCcc1kzSN8labm/vVe+Ufm9JD/nlPETmai06XsqAgwPdEkj8kr/WftYAsS
t5+Jk43uPmQzdnee4oTuwl2/1j3Uy0rERo625pm6DMm/inRjTfk3ouxfJ+TMCvk3
M+2W48Sxowwx5XJk47KFVCshFFUmtEvrEMEQRwj1ME1PB2VglCYv5B1cf1BGSGM8
Pq6llarF9UWbIQ2ECUP0WEqRbrCvNiQu4rNafz97xWAtFHmLNF2cneXB+1kPGX5D
h/9kXJeFljix0oRMDySYGZIr+JyCHeE7xcoxPK4h/U+AdqjpxvNbxSgcJf1wRYve
dOiFueUD8JBW0GN41nhoZnOAvZDB/IZXpKxF+c2uigFAnME5ENzgLgH/+En4DImO
aYcs53LqMuKWMD6NZ/ubU+IBB0ezp0OYD/tAc0jAMmEKPOosFXD//lZWs+JpmEON
ppF92KM0QtoDpMUvPLghnhULDFQHrp7rxa18r9HSOzAQaviiw4nuZrDS1+WqSsSP
wIt7uBIyYQ6inOvv5/7aHVzVP4ZkoB3ZFH4iIs+674g4vO8vvetkZtlIkshBGqBF
j1nCsBINER8yJYI7FpD7JP3Q6I06JzOhSZ0JNyCisBnlt/DwDIkstYzhhoBQJkrW
HgGohZUdP9q+DwF/4BN3sEAsPsRcQbj4JwBvivcXa/2TAqtYxcirF1RPETo07Ka3
oDJ/fhpHvxmWhoEW8p3H/6i0oG4nMocUNQrGVQ3uZJ+x4SBYRB+P1A1CjWzXVOvn
Xe864rhhGmSbl3+RrR48mPKWhhrA/JqeUO424IDiBCXHLiJF/W7LFX/V3d3jfeHT
/+ae50rhPDBVhUQulIMR+LavzXes2weIoNpEPW/h0FGteRMQsK05DXGuWiI8ySxi
ikGnGBqggvcVh8tFP1gQZ6JV/qWPKANMtdf39aYhFDPdVB2hLKr6d9gh/Xxpp2c/
wDR/nIv9QfiL/rBlUTIKmqsO7aUydS4lN5akJUwO8GtF73EKfs+vKrwK0Pwh+UMg
8KEXDfmxxszT/bjDdeLhSBJkYeC3wcQ8B4ZHYsTKetIym9scUiNUP83KxJKx5rpl
JP22NQ7IfM6rjmqsaixRybA74cUeMTi9um6cz+PTrWmxEpG4TnxPddHYfoRXC6jE
ndWg7mLZePrM1WteBDZxJwsFg6qXLCFE4PrV6w8Ks2QSZu0aJwdHCMOXUBmHy5j7
1ViXTNc4ePt3ZYEDnqgeO25ORAVxbZ9T6N7QfSk84+3r9aLUL/CN6IMgytHFUe7o
9K+JUaw8gGQ+AI4dREUS4V3zgnvOnM/ftV/ySXok95VR+SMBRw6UiafORbID0Zks
ZWHONJOHU/mZv0kSnzjmnsvjdc0wwM1sMuclOCcQdJneAHCuLf7bFsD9Ur6+KWXT
n01Z+YItn7Hi9j3En5bgZSIEJ/+vraNZRX8fj95NP7sTDh/9weaFsuzqGm1+AHCo
j7HnjxbXLt7+887iRIN+ZFaSZM2GGShwfcK62X6BULK1g5TXi3jrFkVs2EybJ2fO
WXx+Uq/Zm7kwjM9k4lkQsHyKON6yDcQKg5tXfhgc7CRS4paQeG/+MPDtRl2ZF8hx
0E24Fd/eCWS2B20cLRgIRjwBHgIVCEL840uqf+ef6SJzGVBuW+AUwbSqCSinqTBs
AMvW9CoA9X5AKYgvOCcnfhgUNs9EAfncDcAPUZSjFpxw20ThPXuTB7nHxhuX+zQ5
hxFP3YVXDMOpxbCH7RBy9Uuq+XBHqpjq3RJR27MUWtlpVzVM2zQOLh7cqZwSFbPF
4wAXpNfHH92DkjDEsXDp+PpFmHFtj7xL4A0SQbZ7X4vbZH99T/CkCHwkmv/Kv2dl
JGhs1sKnA1mHQwg/3g2HiYg8g0/flmwNc8Stm7xspZ+lynIN9Up32XjZs184UnU7
amrimil0WH9v/X92Ov39sEWpIpQ+o2Gc+z6M0AnPmYnpmLwtDy3x8BICXj7OxBgu
/96vKqGRibL4pkhcce+zdR+39i9Rp1IKptOrRuwiRyrS87jvDCorGCe45KcfTAoT
i3IOdGu7DeSXKoF5sQL6Tud8zmvPPGikWhpwTo6p2+ZCz4oXWUZ8lfEk8+b5FOAI
aL/8U/LGJ2ibZSLw09mebgHCZMNy5jPfIYykVpzP/3F+00BeADg6XvBD3HIYmCc1
zcm+S5KKJnx2/vMJnttPHN1ppbkfd0d5xYV316YCkPqc0MOYYmVss1zRbn3V2D5u
bb+vc5p7jvJbGTB9CNpC/HBCJaqQTcd1Jp+IiTNhehXThX/GMf3ygRE+8jRCd+Vz
BfYYgKvUVcABisH5UM4d3DISFaLf/Kr0m/3Qt7UhW0iaCV8XiRJmQfD78WG8mh1q
zbnxRPHQmDJgKUKBWr2SpHc446ncr604CvgLRNSL4M6uHhRPZiwx8EOilCu4BozF
YOA/03US9aeO33E2V28rWRrEgKUYQMqiqHZondwYhL8qxT5/gA8gCRkqUGpMeFAX
pufkj47sVZm8pHakEnEh8OCqB0PYvWqjj8qz4rCBATHNpGFzQFQwRVzJ3mNDN8Rb
sITxmbNTe2IVTdivFcrngAy3yYPeVWzxFjbI6lQYYisTdwjDo9gSZhWnvPDZs9cm
f/OIoubp1cXtTHmYZbq+0E7DU3rmiTP8UykcEVe1fKpZLx52mmsUF3bbKGB88rlT
chjODQiokMuln+PqzqW4fsAqN2YLvxCtomLs+eLRWWvwiKcyKaDm4TKRVL4UEhd3
cZMdWO1slYXDNI9lxUR+Df84yGyeBEYE23r4poEZ5hKiu9Z1RdELWNkZcerqfZZv
ZJnIY3+Mx5KCEbcaefTY1t0lvEAk0NBVbkdewF9LvAo6RKLziFqGcoGJEWWkh+ni
5L+iwE/pjNVLu0kAG5OGxq+AYycAr1/OzL5aENXia8lMJAXf0Tavv6gp0H4Z5HoW
d8A4ZwlnvkxYoQkGx8JysZvaW8GR7kkaYqD/Czr95ChOLiqKxpLn9X/NLNzpnVG8
aymYHITErLjsfYS1DCTnKQP3SrkftD5Q6W5CRBM5RxQc+VvQVQjpnnu0RDPrXeHQ
K03fOVyJsElXYcIThtV6FcflcXYujVE7JQ97/uHtdekn4rpga2ZjSlbz1sVLI7Od
LDMT0vipGQdeKWl3SqVOt0z+gG9m18zDy/t6jt9ADFVub7XYJ48sx71Pmpc/FkKB
nf4EOjtb2dfvTO/hTRzhwdLfkxS5vtE7d4drXzP8QmyOEsapOZmqQvyEq4isVXwu
pzEVqUW7SoChJi9AZSy3jmIW53K/hR2P44YDsl2aHryQfpIgWKQNSbA3U4u0IMKD
02oJTyg5Y36y1Tf46d3mQP7CxvMoQqA2fowN/yU/YQxuBjI9AoSIVxW0LLQj8pu7
Y59lVw9R7b457Swha5Zt+CeH6ZdPjnAgiXUNZwmzrsbMMbW6mBoo0eDGhhDKl32N
n+cyK7T/anZS8auUEYuNcRglNiEYMm2sgQ4earD9v3Nd8nI5iuDBxcAcPF+XiEvl
qJRYqEWEIhFgmmv4SE0AiDub3Tvr4BLsmDTU8KQJeFqQlVAT0SpslQ9jFEoaMIWB
zZEYUMZBfnSCmDezpN4qUxhdwee9Ae0A46rPRpBP73NHoq5VUQINhRdI+w8G6jKY
vCOCNYfMK3+U5ddmkfTaGbGXZwcMMWeYigqofH7QePcfoTjMaEZ0b2P0mJrJRXnL
XcEnCGNr4+X+EYETa9Y5GWpzXU/dZswGqI0tMm04XvayhsBSzDtu6WLJlcAuwItZ
QdRL1iu3R3fDAgvPUysH9VXPFTFI0WejaktzChN2f7UPlEm3FE7YF6l5VMId/JvX
FX3eB1ytN4VZ5dkt1JOy36M1DmEpPW2rT/01BDpuiKeNxOdI2qX5ilCXyLGqxghm
HXkJZueY7MCEP9Bu0DzKTFBPv9FBTCsMz/X5jd/4k1ZOtFNkH/MO2sI6b4Lemt9s
8gMjOJNRS8DiFX7TOKC9cYx/i3gK+m8nVLCvEKtAh0ccn/mqzavxzeGhT3biC9tS
j8hIUqxjN5jcW11GxhZLV2PskdXTYbHyERR/K7xl44uKRKNPsu4qSfTDCd+1cuxr
ZkxS5lFjBkD6RQfcBKX74GHiKuT81QN2LyJfjRozniqZh3tf9SFQVqod67DtTY/G
g4/QYfdC2WZpFiJVKPo0havzuJ/NGi1SQCX+LjeY60DXrPFP0YeTjBx0SDGWIecD
WMv3MTMXPP5d4AgohuHDl5gs1U5gOZYlkm8br2Y0RwEMb71t7zBD+yrowlS6OyXY
ZLOv+a8D2At9FAtx8mlXRsAliG7TDQ2CZ5aU/YWHe/vx2RYo/o2azwW3gjxaalZZ
/3p0CD0aBHLW9MuTntsyltHetyVLIRT49gSnf0K79ABFmXghoLpfrde5MHVTBGlj
wMlpbAE02HF5nwBz6QaCXdhH27+TOpT05E8RiSdIzOH0VHappkzTBkowFRI3xFMf
63h6NsmmoiNKSwZtgCbAABQMwBwGU5P+skFSgHRbP08gBgcvJK/AU3pFpBClFVg0
txYDv5+VfP49F6t9kyTm1dpAiOqxhtDA7zShyRsBm843ipaWG9ywbH+zoPQYsd+y
JLBa3ojLGanPDtvJ1lV5Tv8nB+3h8jcvqJAy0RDYyLWsyttpQ/Z5p56UGSKGSvnU
xUbTl5kBi7ejVH9+WFQZESzjDHRD6CdtvSyyRPjQw8hu+kEigZpYFme02dJ/j3G+
5ifvRgppa/MJaN5grL+JbmblZ4kihFgRrDX58KcW4RgqVbUnfaQuNqDl0uoNyK20
qnJc67M47oDIi36gDHyjpFQK+ws5DypXKaoP7+PmURTCMrcoMQtPzb7qH8xoqT6Z
yNkEjEsTS6mGDCBRuBvujaiNM7iBebx+wCurIZPbdSVjafHhisWiO0iCAEI8v/q3
jsXTvPmPadJ/UwPXXp7XSdqGxzqrTc3cESX/bxwWIjzqUr6SA58RuZmo39Tlxk5r
E35olxi+dUbUFhxZfh+jbtQvEUZX+XGDujjkhOntJgCuxQfQ/4+bcaGqxopFvInA
/fThwSMpuM+G9mihGBbkUqKhOOMPXR4kJ9e9cxbRKZSMA2sjtTIKgSVtnsyUV2oE
e7n3NoKb8eO1SQut34MWWvaAhh00SLTXHrYi8R8Xz2iCFqPvs5ro3xve91KrB2EO
FlKhEMrS0XCWY9BzUgmyLNx23SqWn4szN1xu0gW6GlKR852dnD3JVtyzcx1k886H
P7FSM2sF5/vLY0mXX6AMlPX49Mr76R2u5xuCs3KGibc7bkuvi+YgVP8RSa6Sheul
VJDi+lnWqYHC0v2s+mWJQvI/R8H1+Q/zk2e7EsuzG1qvNsPWs4erGdZbVv4Mq41K
P26lLpYf7EgqdHFF4PWv4XGq2/w1N7iGzaxwhFJ282/+6VeE0njKMsCWPJoLzs+K
WLEjumTbDld/KkJC0AaJH5YBItB1VpB5dOjuXM5fkTqsQDN+hOycJUS0oli5mJ25
GZT6PG2Hy+Z87pEZkkgqi//wuN/iVpRMuiZeoGaDpNvAzyelky1LLV1ntskKURbi
J6Usp0J3I3Q7PvOKJH84BHC+180owrq8GxWduGmHzCIxpMbOWsPm6M/XZxMgtVET
6FAifzQvndBiWM1kWw4a8uH5WSfdZOwD7+3LjfGoDqknpZxVMxXFqtyAi7PpqLjL
x6Ui3QRCWuaQ5OyEdGpSJI7zd/xC6dGypNCbaGtdTwu4eCe1xnl2Prkkiap018If
Q85H9oKNujBp5xTHykm7NBwrs4hC5fcS46gmNYRHq7ddHVhmDWcaVnZBOA1vs58q
URTnlm2MD6HJOk5ofddzZmGXVwWGCwL50y1HipbjkKjiBMwxlgtEP9tkC72/Y/tH
/rEMKTyBtkOt0Uvp94aDCDETdu0/oSQd5flo3piuHKHYF8N2qG76bSBS6ToxpuKV
ZN3pRnq13X5ucAXRt+AmHPSz3maAiOMIBL0/r6q+HeACb9oghtq5qNL/XjRq7EQx
HJUCTdZfhpMwphisZgyFEGzyZemGs+fE7OynC3sjVbtPJL/B5caOcCbGbR2VvRmq
X6o8o+bgk8H2mS7PGst32CodLmCXwNdu7P9fhyRup4zBVXOEoZv/a/76dCfqrMoR
hU5MjkIQ69fypHuhp80LoC/Y5Kc93W8k8uwEclRxuKO/MzspzHFnikQ913HkbIdV
eUox7JN1YkBXKjCZDF/joYH8R0QUFJQlBwZPRrMqAJKXzwgxTRfa10x+fDGrRB8r
U0YNHe9kKH5dJ2N6Q2aKNql8Tb/3W8fhMgMqaEpclvO4r9miibWuiI1a5tWbdCHm
spfbd/CNwNav6FxF9OcpYtpTFZjKYO+saXe4i7agzTOVnlvtyZutRkwsZpY1q/NP
qEPVO5TczrG3r3+4qXJWTcsGX6MI6sd+dOxf3fRbzdT+ajm0/goLM1KTD1iEL/xD
kdJDaKeGitBTyQzhPqjK1qvtMsN2VuN5VGE/vBh3oDayQUyyFGYQGJsUpepcq3tZ
tzxvERrscIX5/mVZi23JtCD8eL1bsNNoCKYobBCfm5nt+/ezf1HL4QpOKIlkfO9j
zYJ3ZYuOuzt7Ff+c0sIW4c1zrjbTNS8SRfUm6UIHijvwMSMGqS5LjqNw6McO/ANt
RfrBsQnfOsXSc5Ojbdehm73T67x936nkjnrz9eT5+A6QAIG46rheHobNnXQGADg+
UlPzh4ZtCXUVc3pUXKr6fiFlNB+A/9FXQ47XlC0jl9hYYeVhUPq2+nfLEBr5Sykt
qNk1tYrOvlRO03WsBc2BEDGYZbtfDyJiv60ZNQQWwSujSnzBwP1bRYC5MrqG8AHX
lcu7zOhEnGt3Bk7KiexWenkG9FZBgPs5KGTtZm56RHJCbDQDZmc8lPKHthIHndjl
A9SYmv0NvU8x7UEfUuwGjRsXCtrW/0RIMTstzm9xo49Evv/3B5FXUHnngqkjb47b
dfjS5ZbGbhaGevFRtSfwkS96XYwQtCpoXb1Ivd1BvDIbsJOBXHRIFSkuSGCXYIEK
Ze2sFvq8iHki/NHM9x+BqdYZV95GbtqgYVlXmndJt6MwfYozDZ1pztZODFf+40Mp
jB9P8gVCBfXNppcfJRV5l3po0w6KFSaYHP8rb2rXSo469ea0cT/bC4DAq6a/DcyR
PnXpAS5zbY2hkA+eiRVUh/hE0qkMORWb0wsRunjT5SdUmAkimV1cOJNmmmbb4apa
SRoXv6sV1DT8+75XgODDT1xEU3rhH2nrB9sKRy+ENx4YfJIWAAYqy9wYBUwS4Fm1
FTvPf9L/DN5wqARa5viLuwQIvJpDyfC9ILz215Bw7GcSAVUKM9ukWujhBODkLWsU
wUCzzC4LmrRa78XTZ6XpJdrrF4aYSAiTUI+3/j3ALbN6XhLZ64NRsXAjOa6HAC72
tAebIi/N5N8f0IU1ES7vCX0mYRb4XAUsf+zR1rsT7ezIpt7Qt/zfYoVJk3MYK1Cx
3uhm+s/4wCKaIC2ddL4Pl4eeLKqpZVmvMFSEWv/3MAHjTKL0sJ0PZPqaPrnIRN8I
RKN7FFAbxoTsyrueKb4F/QgsVSDICJk5pv4cF7hPF1jmBNHhOinOaWRGOqJ836Hl
CooIjvGyyAhwFc4a3f0adobrXnCU6tGFrGqKGujx3qiFgiPIt2nEO0TwPLGsEMYF
oEVeR0MCKRhPKWUagcOKRBn+JO+VbZDP+soCLFuW67NoGzV96UcTMbN+DjOPR0dV
ugMCERIdzBKz3VagwRkGXXOj+fh34+FS8NYik1jSXmlqTdkesUUQPYixrfexg+9s
NimENtOMHgoW2uS2eAoWS3VZyuawMAgfBDvxy6uPRdoPY60MDY5+TNu4HcIh6t1m
lWjsTbwtjx0ULyNJ/XI/WUcf9qB34rxTN1u+fWWZC08NLyQ54cZW/+Joc5FnDVDo
OVmFL2m4l8FT0yLLQPXKUjJ+iFSkrfoZbkqvCjfPCcxgMIOHkdib/jI+bErf6V24
84cfzCr0eaKUtvOp+b9Rnk4K92dDnyvrjtfe07w7m3opvk6k2qvNRGuifouAk3nI
NUwa/FXV/Ivm1ejIW+feSFStZtumhGv9cCAA91nyaFCE+ARUIy40LaCh5D5DvmPj
gPKlXyigoCto0ekGwkE9t8msY+RtvRRzLmHx9ghmmd7xQDV0cy+52k2ywSaApf8x
U0TyVopbGEN7qPoNv7vc4VTrz9P0J1HJhDa7e1qtCCdd6pm6auJYRQZp13nnrNzF
yp7CzYVxntZYEFmntHPfWZstQoBmCi9riYTPY8C6usJYdWcnJ0qAv8vTIWjBqIlw
jTcIQ1bLKnVggERwOxpIOlOjqaYa90Bhzc+OsXhCPFvHVyVGigl10GpvKeMGo17H
a8r8nNIkzIUqRm5FoQxzg3zc0h/AT73zUyiOwy2lFR/gJHduSQCCB36L9JpSJWk9
KiJCgtt88cCu45ekBdijOJjAPZCRJYcDzTsjcnxcXYwHztwdh+wVhuUAtEXaY0s6
l5YXQn8BSRxT3mZKqlHo7qiCJjiynGaIVFDgnSg4UnhbiCK4+An1FcjqYww/volR
hBsPhAxDneMegjXWdhi/Ja/ecg1T3K1TRV9SEK1wyeCJCvTS0Szev0vrCx0HjyPV
kIxYVE5o7YlsDa584pIn5Xpnoaev5o4SQJ9fq2WskyMofhAsTr3Hfa+wyIFkWfRu
yXnFAPGQq3GIIh6cRE4WT3C6tr+MRWvknNRDTonfcilgYoljBVJEJUo+IQrogn6k
wgsoMavJ8c3L6BGyCrqGyr/g1s+QE59xb2fyr3IjU6DvtIO2efasAARKZFzH+8iI
JBQ1/ZxRvVApinbTBdB5Ia+kl8+3AYHPNNmPLaJOm1o2qr93Qe4VUZEb3dCyQfzs
HpyISxVtelvvy3GV8EfSpyFUVbkrOuSL/60u9i/nHo1z0lHvG/FmiQQ8QkLOjePS
hba0Fgh2ugweByFFgXZMUw3uFnFiX8YRYi3UqaaCrq+lr9BFMMEr8+bZCU+WhZ/O
nNelcg7BsHU6acuUPs0v5IAqxVNXC34eAr++lYJkALD6gp5FLY8R25W5c13mKUS1
nhSCkocgsYQ2PMXHuPlFMT665tmE8USuDo87w7zAeXf7uD7xiM+4QLsEaE+Kg7p7
xF1yTAwnUn9nd4y3KhAdXOijFHef2gWZrRraBnIzZ5dfF+G/sWdmgjMSImJ+UJdI
k2NzTu0ofTQEQM/JW0N3AbAF4TuEYDnrVamCJNjmT2mJLW6z30nX6z8H/YPZaqqR
4fDmBWw0zGUWvPBDFBa/rHiv+A62tHQ4RdnjluFuTagzdtaXDLhhoi0ERfgt+oQg
kohHJMSTCe56aHbvjyjup7m2b3KTi0rmJ0QG4oow+vX92788fegg7NSqIQlES0fj
cEiBlr4fj/0OnyZbiY5vsPMR/98YVd7pKaLygYaE03zeNrj/xGnNhkzoN+ap6LWo
3RwolGxcQFXrO7AmGYageYcR4EZDHDs0KIowH0RlkTXXrYIhNlHPQNUvAGTj7hiD
fHeDb/mZ1KJeQqIuWZCLk8fn2tWeUfSJXtM5/V56268a12eQpeTTlnXRKIND+QWZ
YejQqXUezhGTxPQuQPw0GSwaYrdiCbZPQdDLQ/Km5sPtJIsSJrLMslTZ2Ggwbvu0
Ld/gpI+Fh5NduAZO5EAIUpC0Kt4YFshe8dXsjD4CCJWefzD7/lrxsmmFaO7jL82M
Ff3G7R6LO8ct5C0A6OXKzoEH8WHc6pSyRBgRe3FffoMOBRjpySUBX9LzeT7fIYvU
nKSpjx/iEdOKaW/kJtAy1FQFWMGur2zl4mSBCsR+R7JRqi70liLhfqZG+o3WT36Q
oq8trYAwdNtlt3r6+0DVKiu2SRyJsSI1eldHdvmYaYTu4hU5t2T+Y6A7KGSo9mDj
/ToUkOYWpVqXkYi2mt3T1eiSNbkCH4FXlDvd0Cnyruval6lVOYYa/kh67rhALXCR
dWL/eytepTr+fCxckMxfiBkL3wYXZyLi/42PaQ1H8mHls6spJ3yaxHDcSA6kGryn
vD+0oDu31fv8UdNTObu8jHiTqWOWlG4vQ4IgS1ddnu99dpVSmlXR6P12Hk6vTQan
1a9CZGfSY5JDlCVkIyRDBPxO30vqnq+812buIyS6klvA/wBJCmuNheNn/2XgrRWK
XQ9DBnQp5lpTC3ZujRFhKztbgxe3rT0LggQp3JXSYRptlPPQDyyvSmUyJ1upvR0k
ot9zjhjmCLw0N1R/0NtPQ7Jt2mn59Pp+YN5xFNQOawptWkDtKBeDXKCT6koAuJzB
Xg+is4oJzvyJbWjTu/cqjkO4piqePBjcyApZ8gd0Oyume6ahENVCesaAmD6BA8AV
AZV67f97hJbHsdK9FevnOcKOyYVO4D5B7eXt5w7Zo/S/QoeipuNic9gSmqLDg7T0
r6/dd6/lPQF3wvnA0AbasebIb2Nz1fP0kBF4BlBj6QqweBPnA1CzNK0wMj4caRql
Qb/zHOA2+O+5NsgVT4zvOFNO9YUz54JQahsCB+4h6sY/PNAzszfbgN6y1+/Q/zGH
s2lzgJKJhpB/nEQBPvTor9X/rh8VJpNHCRo2mDexLF+z8ic1NQ3BocQb0llR+fU1
hTWhpnJxYWCSI6UtLH6O/RhRkQbh8m4aW05RuVNMq2Fz29iEGaPPJ3/sVuk5LFg/
ESDFbHxpA9lnPc90rmNmHBzKMEVsA09BeCLaDDFhc8DrOItyCxtI0CS89OXg0Mln
/gvcpAkTTUgc7LzTh/8C/z7/QGyvK/cnehZeS9utwiMQPfm0mMq0SrdxnLmyDn4F
FFWPSxalM73zsq2EJa/e9Xz8VAT04GdEJk/B3EjaACFBpEX1cO87XOhyanYCQSoh
AJtsQo39WCFFCWb6zQfZmHBfAnzTthUP2oAsctf0CAO0YTWQ4YzI/RCJXQBoBFj9
7jgpF57bqXRKuzYISp+WJHiwm5+rvCdGSFx83wJww4pSl4T88EXCeaFD+b2sN63E
T3dXW94Rg7fEMgTN0CWg/4x+RMVPSfI1ZKJGxfClkbHuh4lYdatYYDYW5MuGhoZ1
eITZ/CYJCbALMPNjpb1ulTsUvNTDovg+iTu2XhO/YItxj75Hb0i1rCBAR6VvASuq
k7ovkw29uBr+o/gpI3BrkGOL6i/olvzlEPRu8zK1vfVQ0RN+EISmyivhl2lKux1B
KG5/kumTNZN+y5UJB8CrOCb5pECw2RyhkIqNz2PJle6GHAjHvBq+58QdJQvEwNkd
3fWt1N8IRTNTlsRFMBkXKXvqwdXzLnk+FI+BgtLYJwpeVVDDlxekz8T8m3FvtTuf
pq7rlrVb85ZKMZViSXoW3X1O1aBz3f3xOj208mLyhatYDOlfpIMBOQEHxvZsLT5k
9xZInMP34bzCYceL3nQsXH/WzlOfqeBo9Nwr2eKUE4F9ZxjJoqvX8e4XTHTzLwu0
Ki5fusz/Pa6/gDP5IF6C/dRHXNHdAZpu32kWGYZ/4UeGeYJLb88KZ5DsPGhJhGAO
ad+VpNHRNBuqtXVkwgj4iXJa9EWyM7csHXhYAxCXztXIneISEjGHwLA7Wg2s4uIH
iCquG9hfLP/jz/BzxG4OZtysw1kpS33rF/Hp6Sw2kZrbadU0ZsIr25Ak94REPSNn
U+QHPAl388ihBCqNRplg4pk3OuOEQdf3yqPvqFU3x50CW37oRPY3DlR5rEU5u0Qn
ifxjcTkhX1dgYIOMHL74K2H/WK+WxFnNCw1nk3v89v0v1dBDH8IyFZuTOPSrXPHX
zGr/FUP6Bpnc2wMzqxzWah7fuqLX6t3MVbxX5Yz62E9Ek1lvu8Sxkbo8EjrTsgJ2
zvQzzvEaLivnXL6NFSTM5P7EUl41z/MoNC+sOTf02qH5OajRcNaA1dwNa48/bKMj
b0uRv1WuQ0JTmN1cNICrqJ3BYiO7RpSVd9cuFkFvFdvZ3994zF8ucmZhYRuzCVFK
RN9wZeI2bO2qVZWV4hRQMXx6oY7ZMzmg9t0qK8RIb1zn6Z5xujRCvo33YcvuATop
nmYUah5L3b/JM+RcZt1RilnLNF8HRpoyYBcADtgmvyrRWMbtNWKeMuK62EMTtACZ
pdUHXy6uRFCrGXRWB0R/SKi1peo9GD3pKsM/Tz859JO3EzDs67phYM86qYnIu0vY
nVRdhOCEsQU+hwQLVQ8RFlIDAGv4PE5QZ3Zj7P6F0ERd7Mv0X7qJgRp1fncOTgjn
+GeY0g2IjrByVmD09GY2ZRTuo3HxOAjc3hXCKW/h6XorAkBRQ4fyTPpIky6FAqmE
qRubEEnA9JhTOmqOQGnYZsikb6mMgSkwUIGVCLdLvhv8pUiN5YMEv95LV1FDbNwf
IQ5XTz3xCQS5HZkCmpcI9xWqHPW2DukXgBqmOLXx7Fje42Nl8S4ON6e4iUkbX6x9
ghIJ+YST3eTLcjQOvgWECIaaixALSFXBTGaOGGnK2v/LDUS9Usd3KlIiqMUGB+Po
7ImDORZ/n74GPF8oJVJ4GP7Wuvn9pxhegOI7eyI49oZrb9eSyqegbmSKFApXdms5
xY1ocs3OfvwCNTTkfsDKMe6JM18X/vxOV6YL+LTDu6sGJxDAnpSDWSjopEhvTmTp
U+5zFb14hkBbCP3VDgw/WF1gN/BTd+kIDWlyVKfN7T43VGDbCmxtT2iUG1d/dH5t
B55bkX5Nd9ySoKiece6YXQXhQ5UMvep3im0e8RDy5ept0cS3qvY2uGwYE3PjBIgX
nebOfYQNpdKlFvLQS8illLDFDW5Gn82h+nBMVnUX+ZiQfbW0L4WOX9mo25AflqDD
2wmths1EcQABQqxr1lk7YgI5u7JtRjrONSpi4QLgxe8L7hUbqNxJbSlgT5VxFtNw
tmcG2VtyTqtrb443ivmK2SpWGQnLA5Wrwl9P8SilDbw+MGiJ4yct2/T8e1yxsArS
npmCmpuVmYxy+J3rb/MVhYhKrWofJD3x69htLJjQhA5jA/Ddo87upBeX3CbkqyjT
3cX6OEbigPu/Wd6btLkZVPr0S8RTCy3yASEsgToRdctw4HyW6T9w68mBb71YF3sb
kpRKRWRYKOSg/q/VXd4dD89zGk0N7QOT5F+hp9mdwUM5OGFyixE5tTUO1qZYdlGN
4Bl4sck6CkjXo2b4GZZBlsZxvMHtHEOOUGtM8FrkFh24RZ4iV+08QUfICKotGGk9
X+NTkO1gsJgA+E6sgYyQRoHUiLPWlj5HG6OwcqPINXrA37W4Y+T96oH8r00kFb1m
5HWn8/YzrG6+VEFUk+73Dccwj0KTCQAIv9MI6b7fiPDCY+sUqZujDAUOxwIjExur
iebYuFaCd0zo/z46XVraygv1wI88cptg3gEd2jMR6/p/jxn+KqokOTXDvy9Oxg37
rJSUTD0raSIeGMqXESQv1vdxm6nTEPCBBp4fvOI3KCiAe2O6rBb3xkVyApIPnlDh
pCG9A8o6ggqkpYmJGnnBb2FPa4oBAOFq35kumqaifSTGGuPdeyF2frFDI04qH6va
LATJZWEw+m76XKbuEqczRLwubcRapdpncoYs3qWM0NZITIEFh9N/atUccT+Kle86
N7ZM8WsOIc0xMPkCEnPG8sWpdvJFvIJT+udrNE4mWrx5F1Qvplo0o/Esrc7oL42h
9oLEGiQaS7MzeJZ12TmOk66eesqkZ6bLVw9cNHeK8VwbszFKwk+yjMqcJfpsx+RN
57QrVUsLIvxgPjCYiDw2FBL2SdIIsObFEEGufuCAn3h3UnQHUP92GqIP3g6hsrWh
KX7dV/QXhClMrtwJHEaa/phP+Lygpx6M7dHgwuq5WfqjMFuXkdAkgJPtfcKczTTf
D7JIVHtg99HYUZ1zD1MU9QX8hn7m4pgr+HyP7ffAwR57L9GJiOf1p9MYMxOSJqMh
1pXe01+EuBGG13Jow2WQTG6NVAx4dAGxGanZrsZ4jRDNrMf7RAyoMk2BRiUTmjSY
XhMQ6DBSTjAEbjzwuyZrpkvhKjlAMuXCnW4JRxBK8EvIaW7d0nl0Lc5CHpLwpkt8
NzrFsoSVlRhxCzhrdHM6bL+Ap06gB59NqOLn85YYL/nvWovnEXUvHAqzg5jIBA++
6np/Rrb1SL4n24FpN7lczIXkEHkWV+5MWH+DwRd+I/krMyNkm5zWkDOS8ZtaRwlA
H8nUryL/q+XIWMkAYmY0tcZY8TYR/DeOpTHJ51kGnSyUpq+aJR0G63pFiVGSML9p
/YlXU2TYAKfrg3U2SvIhE5N/wnDIZwVM70/g+gsuZomTDF8yIKL3rYmFrR/xD6/q
oSN53QNEFTtvAbREywB8rGxPhiqtjgVZWALoSBqKzmWALYm6DxTv7/Pv+cS87CYh
oFXzMRx62uLPMqrC+4bn5ec6ibD1+4VzY3iqAidXdJfRr6h9FZ2C3Cs7csfO1IlI
Jqp2SDtnY1PsXdmEImG44WTeqZ7ZcZ+UD+K/sd/Fiz0LX/OKkDFdBnqVAB7K06Yz
adDtj0Q7BhuEhb2u76QtyksVPV/4/eTZiIe/bLeQCAkmWRsl5Ve+Hp+93EO0cJjs
Fn3Q2QR1yeq7NQNzM8UVEnec7VibSGD/pydNVdtSGrNN3QW68tmGdwrOTDJDSlw6
jbdBl9a/PoYARArvl/HO0s+TCbimrVs34yD77qwAwjLobM3y4LOomzzNPFI6aC1Q
dV8LaR8dCtWwDjQYVcm9Mck51u9cIBEOqtQEQ0+OnhA0COPFIF4Rj59aV1V+prrA
f4u9ec00fNok7E2NVRGWTr3WxMBY2X2RDf7fAbq+iJlJa+M8kB0uZvAFqBO5GCfu
e4mQ+A7mIzjB8VN9RA+PhG82p6PDgXvISbAb3L7DY2UsOyAaSen24taJlJqtfOgR
eUelseCRr02PGXZOymaBYJTe+W4H+sQeklK/oFg6I10ajiEuM8Ml2OIDUAl0Fu+F
1FGla2upywsttpratfHYNG5aGc3iNwTgvSXSsUyJZrXhWYSeIeRZ5/MvElepkZwo
vXnunHeIXwl5NR3SWKQ9Gl8ibIoVWw/7CffhM5AW3Y5vYymOIytS5VJ4f97PFuYZ
BjxNNpSCTVQYImxzlZ8v4wANA6caavJKa78eIEZLiWz1h4tRGd5O+yI3Q3iBUjb9
RcxMiGHc3nLvdbMy9muDJHrhjjO7WEhwkEt9A8UEu6jzzVktaP/RQy3r/OZVRHSV
NpixGLha4WSO4+hGTb6ZdnsR6ZniNVNu+1Y01eqToYXDcOShLVeBJQC6CnOGRZZ4
16VUbdNZJcIkfPtwQyWhFYaTZaJTiycWD4CultaKzn6ronvTIU2XDY4DLq6NpTNg
knGRTadScKaM+b9FxUJnezg3lWzYF0/COvyLGqBg8x34qGQuzGEQ9NRdJ0o2Ckgh
eF7GNLgYSNqW3b1b9TYJq9Sc0aMDnP7sw+YJsiZaE8+jaLdd9VAShNO30Pp1dZyc
cgyQSgAkky+ijeJPWz6DcIEBcVpLM7wOVmEQ3k5i90hClbhHjCkjwnpcLDzvuWAC
0iuLhb6Rjrm5twAJWDc3Mo9/28ZvhLM8XSfrhNoCuDjwQuLXX+OkzjK1BhR24xR9
8cDbHHPMMpsoPVSqpaQIqaHsRdRZeXLLEkovnDI7C4iIpCusQOOJF7HW0dbezEsv
DVH8pC7dt5homI9T2zYfe5+/JeWUdXZAPwam+Nbd7KZbdvURVc4TEw564nYSJAmZ
Ed6YhXI5VHkLERwhORw+BfeFjsFctG5O7c3d6WJWaYi6QAo0q5CPZoBT0LKPOi3t
ZeJLeBgSIfFvNENn/CmrY55jjM9PUoyMDT7TEz2O1ZFzUNfSkCVgTvClIzFlXn08
LhIDFwhibDzMQZolZaamnCWsIQ+v+O7NGLwDcvsbC2PjBCxAeoVLCocXi7zcUziB
tCYCAhERMAkWAmVGkXivhFvOO3Q94fdy+V7bWKTl+IF5jFbw53wUltFJDFjkMenL
j6L6/ktODLUucWqIMt29Ugy31S8PFmgTj0smfAGHAN4VGE4znZfxFPjfP1Q9zXw3
1zLcw2Ue+d/UpNfet4z9cUvdzqnq1Z9t5eMD1vsPJaBPKNMiiQ7lY+Z4bZSwPiYV
TXqshvE7mH1kyJKaf2+IyzTl6059YVcH3GZt9IBzBqMm2VmFbbv0X0UWsP6CbocH
AOl4ZevJIYOnexB4boAtSDxdbl7vA8yJ92H/JzG3I0soRxoRyYPMZ+G499HqmXs/
92frpdtGtYCGtY373jctT0ubWIe7SlORPjMkl4E0Kesxt4IQjJNqgDUshZwOrR4h
AOP+LUGSYHvaeyy+9Qb8bzhjnPgfuOxv3vQpYQdvs2FSkIPey8qEkRJSXj5nOBfz
ErTT7BLqkAdYo9sWfjvNiqN/z/2BSwr/1x4MbF9AbtceceP3zzwP6mPLMcopbot1
RqnM3Nnf1bKhXtPnQDA0UEfIxSdQoQYlL6l4p4SAoXCR1qRQZcQCUjxongebe9iW
Y/8e+/2Bhy8Kka0aw77IrEfSDzT4EbRMB5syJkD7KuytdgGQETlyJCEh6h2iTEUH
wbJ+h4Px6H+VhmSlmYQHLZTF+juePHZwDF6A6wb2Lym9TiONj2pJaey61CO7MnPS
eplqf11Jl6LapFGR77IpMj5QrbUbP64ZTTGYw1eRcrABlkGoMnJB4jn4mqKCmWGn
6V6boffGc7BxUwQirXe+x9lGOBRVJ3QQjwQwW5L/woP2S/HXqBApUO6aIECxTI3Z
28fLOiOIf7vBGv/lZs/vfcydZM2mG4Pygr7mkhygWXm/UGr0F5PYAKQp9Xtf1wg6
bX2uDE8M/V7z0MJNurkXXqnp2OUR5K0pCcBLdw7w5ZPH0ibigHDpm5a3GGXdK/54
ZR20dST2w5crSDTGOCMnKmMDGUg8sV9jk9FAubRlKg5Ty2HcHr7Ky3g1kS3I9GAS
XaK+A5sjKNvDdEB/Cjxb1INC7/P6vMjRenWPH6qoADlq4TgN3A7EMgYTLUEYhFqY
2DpHAbUXVWRQ+XeNKm+2NHFpEdPrKVpWGIneqUota0t1k5U3t7orXKOSIqH5vKbp
XU/QrOY7KNDomPwqaQI/jwzydqfe7x7PKoNxkUzAGDvY0ky1qNNnoBNwD0vJ/Tmg
L1mFlOspGvm+bgiGI/tky7PD9cRg72Tb62os5+yt/S0NUmFKFYOzRHsufvURbpPt
s8iCT8QaZ7zFdN84hwzFczXFV/72viWjFAVFzvS5X1KIfL10MoDmRnGnQ4fACfpx
8vMXnfJkMZOuIQWij63cphXCbDtFclF2D50hwVieH5wbcB+dq9XHfCkGL/ku6B/A
VNtxZKHTEcs2owtCruKO21C63DipoPL39NgXayJ1fNiL4MPrL1oZmfBd2xkGyeE8
L3GXAkOiDUo7VWzIno9tghtoK0o8xm/APM8KcmhRQi/PVgubYheFkr+ZtOZXxIdZ
1PUtmZQ5IdV/Dzssi7sAYb3D7Rt2BXyNiFw/aiYM+7UFN87gm+8peg+7PZOGAWG/
O+Nz0gkpSyJZZn3teRyyFAHdQ+MZhI1j7Y/JXG44UAuAqMTbHkXBifzPyq1A9eEG
E9GNFIFCGPa+LQVrdOzhn/xKFy/cOyrU9c6KsRXWHvgK1D51aK3Erbe6iYgA0es3
Qao7+mAozmRr9FC5IO4z5jrlkjpZ5Ztf6P1gIVgUdzKMieGUynegM/JG0zCx6ofR
s3qAYtOhEB08tXZ+F1RmwYdUqecTAEbEeZ2napH9c0BBUY5tpOXpwbY+jh9GthmD
G7Dd7SK5PREAhtGjf/KJIqRVhhjA2juRqCbTEk0j2R8yHesqM7AuN35+qRtldyFD
YYhriackXuZ+hMU6oSaKJizsR/AGpA2LDPnxXwIBMKdma6GIKMIyI6vh64VTZLTo
/5wN68a/jBi8syUjqGQFP5v2YokEB8EnyjrLa1MgQzkGA3c8p0zuT+bbXJVsT+/g
DkyJ0OCQ77mensTzkhCX2nVIKyM6rP+/mqCLRGx5gw78sgltPPBi3888r1XmbPfo
/7ACD148cAZoe3TsIuHulHOXXYKS1rTQz3M+MO7euZXhiOR9UjnGzBbCcfUsSsrp
lhC34Getip4fYk6qRLPiT+ldfmc9mCGewtoMZXJTcMEieBPFQyDrsZXp6habfNDC
nusq0wQDWWkzTZOrtfivUL9VN+7Ltgb4UEnLcfxhQ1CvdSY88+c1Xxxu9gEhuj20
rpiyWEeUNuDYaLk58uMHO8kI2xs2bOSELKoj8sWfQYx7mog2KIy4rVWSODhdxkwy
JgyNUiekbwi8W8SMBecs5474/znHqw+z56FL5f6Lbdo135UgPio0c+UlGSirYgP6
7MJjq7CCyFc4LRgpKklT2n5+u8brOVHLi2ic91Lnt2gJ3w+oiSE2LFCoAkJb+hu4
zXcEZFIScYCQ1Il0a92W27RSyRwdtsjZmQ5qXL2cVOMPphiXtzaWApejiswRBiRw
yhBXukPmD+ilgx5UqZXmkCjBvybrFR/Cl3oAUqC5mWwMX9uXmMfHYj56sYyLSSyc
CI4osRkHlSbUNax/eeuP6OOtEuahds6apThxTvwTxAzroOkO9e5w1lbqm43oqvh9
Y8HoLbB2Iv1Ne3HuHQMwb7LG2bK6YMQEbZ6nYLi9q7BIz/W8PMOAE9OEPLGqn5LC
EcqMYfr9asbap51sGfZHrNY8cJbzYhi2SMhelEwrfoMaE6v1fZ4OYU9whD9AwlQt
J4MjFx5nnyvdxp+lbxYCVsyjSkv/DbdusWOlthO7OzZ/KN//fNpwF3ES8quTO1Wm
0DS/bj3nxmHWMCQ5iAH5ZPX7G4CPlKSXsiMa44VQ2Arr7Wv+s1HIgZ6ltHtLBPPI
XZQdTJPTH5UNEmjC5ORgCE39+OGtpOWh2v9AoI+8tLPPwLFreuAAIt4DfYLceVX1
eRJaHYEfhEiXdIBJcrOPC1Gny1DRmZm7YgX+Z1EhOyxklgHN8DMcTrxQjGeeu9r6
8I6KSMFSz7AsTvr5AuqUTG0AF/tmbrMKZqseP7KtUlFr/2nsi6+sX6Dc8yLvWBvB
vth+6xwppzD0ifU+a9+nl0tLt8oZRC7U3dJT88nB9zfLKa9O3LgBcsKHbL0Yk/J2
UCaLV41o2RXMZLMEcvVzUZ8qkCgRBmbYgLpeNL1wYOBht2uEP9uteQ46ly12L9tN
uiSekoskxguUST6mX1GWG8iyn/kkZSXEeAhngAi32NgagRLuDu0pXO33ovSG6VxF
gazavDkEbdWjri6OZy2K7l/XYA0pbEhnlJYRaKHbPmLXgnh9eOsc6fa30HRo3jY3
ZcXSZIDGplpM1FKzW2kovNL/Alq1vnD1M8KX/w8IiOMRaG2Z6Q3oNaXIzpLyQnYP
VXRYzmqnIL04PWqnjvy0434ng1QvqmR3hwFcTYaTTRFaItGE8Yf/wJhy6Y70PHu7
u8THtlP0JfFvvpLp9wpZVVEsGWBnIdwSXK13v/45gjnfBfgZLfAp51e7x2HuqqI+
hSAo2o118XbCJL6KCUdYFPwsYNvVg9gdoykp6Vgz+ifksh7wxiImOdU80Lyp3gpd
IkAO+3GH/K26X3BtmLPWtG8WvoxLgTsgst3UwW7TvqapCcZW2qKP7X7C4mHNQIyN
OS8B9/4VrpBjurSTM1RSBItkXmbSdNYJat/k5TmRNTmGWXx23Xsarg+feLQprE61
jGVU4+AxegiHSGqptu/SNhQif81/UUO43dbJHRI856afAgVwtLD5Y61E2+jff65l
y4Dhs12LsqTVyStVQR6Qix+Pogu06H36TNTl6GGVD8R/4F8NNqhWFiTOm5AJ05a2
Ds3GM1N9x9ET4hCD2Q7Jrix8JYwHru+6hR8NCYVujR5ijCN8+qXQz+o8GwZhu8Ba
b5BN3FYLTOkJPMMbkECYkhkXt0aiyC36ofl7n9Pvmy7WFKJyv71HmObS2IUIKnwJ
Xvysx9OiwOYLU0lr/sisS1A5lI5fzcKnD8gLCtpsRPjId2jr20tU7cUixi/nJV/M
II41fSkRxhLCHELHkdUKdwdijxlMD/PBwJ7bP9gcOSlfG7f2adTZKWz1cKL9kThh
0sXWVCmRI9nbEegFKNv1zudGJJSqtZyAUwLeVVbhrazpFNPvaQLlRMaw3DhD6j21
EpJB60kpzxsJxPaZ80YB4WYKtoSlJbH1xH/fp2hRVzURK/FkghihdzTWSk/2Q4jL
FQjZ3ikjBSVXwpQ3/2bwj6E43Gx4Tj5hZcfz/rRWfSzfdZNS1s7qkKWjjjgVQ7wM
TyrwRt88qd8il2vnDoKKh6AHwgN2TqiKr6zzi7Ksl7BT8dHaiiyKSo27bCxUDqTv
vOSTMptH3ddX1HQDoanetJWZEx8wj8yHEo3bX8UVfs9Cb0vVz4FKVLh9reUzQABJ
vvVLzB6L7GKkKom7gOrh8NssBJwu+INYNwXNBX8san++VbhoQndmnbL8XFjxXFbs
58XEuiqbSxzV1vTPrYsT5AGs6BVhEnMsfsVU0pVpUWOAVD4ihsUY4ZQMVtRh2rXP
G5rpDS0pLPmrxr+1pSZzpcMLBzzGk3F/9rxpu4NtuLgGPXuvQrJUHyKpg4H/z6a6
OiQsQnjDhX5yCMI9aUszxHHn4i3/Y9y5wjuJlldNBsSYdooOdfFdTPbyhq+AYQXB
ImGqh/OhrFnxkNNLinUwvsK/3AankL3pA30Gv7NSRKVM6o0p44FlCtJobptaeoxm
psa4MB6C8VIbo584KZHb4x3zEUUHyIcyXcOeB7yiOeYZfuNURbIazX9CkPEY5Cou
nOm4R75klNtCgb7hKF4eE2MtZGic5Jz+31X5UcLyO5pHtjR1AWa9NQelJCJyM3Gw
PmAnX+uAOM00ALWVYVRVASh8YxBrg7HX5+Fa/nZOwMpHsQOvNov2sqH5HhmNDBwz
RU3qHjUxHpoIgtHMJKR4UCbAzl2rM5hMTxaCjsgLERNJjYw6Gz0qVyp8lF3YEuvB
T3vJjkavvkJ8unWnzg4Cb4O56DgbArjj/D0VngXDJwiW70tAilMrwzykpujPTfGs
Ts+pILusdyuzz5K7hZvCOBEBaDDLmiY93umjC6RTFcvzigp2LlowRFnaA38sPmx6
a7R7RifdzWmZdfBVWatgDNdKeovthLszZoXgqVC8IO84LitWq5gUMWbEhTNU2gfw
LNLNvQcUOOdqgb7hXks3LDC2WOSnH8r7DrhEQv3YIk7oGIxkUm37me6PvhKXCR93
reHFUw09JrGZG4mq4ouyMkn4xZ6N4LT9dAc5q3y5bF0dbsNIRy8ZReF4/ZIJfRmi
ubNbt6cW+Xaev6D/jbXkz7RVkXdQAZ2IAkTkiU71SBFFI/mEGDmZLLLoAtTfBNRV
KjPEapxHgFiYzQ57SwHdA8IB8nmDszrcYKfJFM0SCxKJYnmgup4/1t+XwGZd2PHA
PMR0/w4T5znHBhmQkvLCA63mAadGK6wbcAODjfraPBNKnuaL3SQMYH8C7fcjKVsX
sZrDz/+B9PP/p71tPMDGqeSxrBR646Ck/BkcaDTsE9TubXq49K9B/U1gnOfMzwY7
5nac58CCv8kqokPmkIUvKsVS+ow6+pI/wqA6MUckaBIfWvau43Xtq/TLe7+dY9BX
LW57qWd4rbTmkbnIusJHgixeyRuIha4hclDgmt4m2QJXzb/6Zr+Pho6zOTXf75dn
uAJ50i82QlWylMR4B5XSQFb1z1orja7qBCNpcUcms8JzaEr1K4xgUSyz/AIY+x6T
cRWH5Mz36BW2ffBQ5SthNXNucQDYM8R9ozkPPxp6Oh7emqfjl3TXtTYsj28Bv/On
HzmWQnCO8MYbAg3FTiJFkIsNtY1o43v8X4avw/1a2TgkyVDqZZNdCX1ToPsiMkAf
cTLsTyIFiGENHJvmZacwP2FSYHTutSmwXCo0xXGzxItdXBVuO6eSR7I3y7466aGn
9Me1KMYxMIGgnw0fmcMGZZRk6M+UmDenv6MFGriXwwvH9TCJ7jUAr5BiV7Uk1inb
8R+kvmQGkI1QocVjcq1sv41JRqB2hH9sTAjmldSbrhPnhIZHuzpNXjU4Hoe+bFr8
j74ixGtst1c3QmJFDKqM8tP1WZ9AxLXL9YVNLGjtdvQGNGJFwHrJrpW0BTSKRnye
k/VRnG7Q4UfCECLfb63XyM63LPYmGOb+/ulS6uTsIfrBGURR3zYkIMhHBA8VmW0K
eeIqfIdykXO9/XmmjsjlHAL2NMaX72TPpzWUE7npDlz38OCIBP7Qb26SfyDTAoFl
v9VwbrsiadSRtokv2HJGff8/mdbvHA/qADakDhFPvGXCdAk8V5YW1nJ8B66A+FPy
yYAHKh9XmHhrooljunNgtvjGAgI3IiCVzsyd1/aTRFQ6BsKpA21fpuiisgAcbRWa
VNxAcMvNMDvtS/Y5/1BLYY3qqFmQi1xV/RovA7GFiFkxD6fKM0t1XFH4JQnroJWo
w9XwceudqEdjNJvnRYsIdrZU4usZgBnugSuVM1MXWMpqJgAEMYpcxXTI72wTFT51
mUiGTVDEehWHtwKEAjdWffmSLHW+Xh4jk8X25czPXCyyroX17ODEo9hYIERUu8A4
h1HcWPN9cxrB5PE9Y6bMVzdKnIy5KCK9Yk76slJL+WhUUIk8uaeQf/T3yKYKRB3U
uZwfDa85LZIz/+JHupThD7STVNj/6jeV5A9tFiPo7NxvVJtCmrKbs09zczOvK1bl
uej7gbe22ijTt7JNYQiX0wyJFORg6VMXuKcDdH2Cdk2B2UToc/XLn8cYzkDTzXq1
uLVVjKrvXv9q+POqX3d4z7/z7LYdYICmmFTr/6R1p5JXnQoab9j3UOmruUCIBTAx
3/6peds50TU7WYbSfYGXb0sFKCWd9GLx9RApKvaS49J95SXep2FUccCyXrfeRata
lxsQmOII38RkgU9mDmpU2tPbgRXDK9kTzMs2xvbfcen1Igfy6aTe9ySXMHt1TuAo
vU8OnM+xybuARqANxuAr0IW4fGaKs5shPbd3nWWMIFTsxvpcL1MBnRMrMdL45fhd
5ESV/d+JRTys0D6jV4gvmnfMd7xxpwig1Ndegz2L/vjA/QEOpavnRNwxYZyowO4D
eAeufK0jYs8JN2LYsZfMLi7bJ3IjL3j0A9ILiLC+N/Q04U7Y28uSmASithXiQH5a
XavF/Awxd80X54TQYz9orF6O8DJ9a0+zem7gERTiOAtxccJvZXINNs9td9P4YKaz
wvyoVd6H2lsFaxoswDPHiyLvu7M+RhfPmNwyRfxqvJ6rqysjVGIJxV784QcNVzNU
ozubLliBCPTqTgybfEFnLm9+Sw8h5Oly0PBv0m/nsFfCCce60uLEFEmsmr4D/TUY
KUPJsPRcot6+dN4tceno5/Hfw4VuIw9zd7JHpr+CVsdXd8NBCwXMCLPvDsUQ3RpC
0Ub9ondkwPt15jPzPCuXm+coGQOMSh/5dJ+ap0LG1wFPzqFCqB6LsE0kymzcZdhQ
a0OMoly45xj49rpUWFhJu0QDr3/iwexeZW8Lv6mkCbbvcRvJHxXPqy+MpcMekhav
4TFJUNCZmeEht5oq+lM84DzlDyWkeZNUVWyjLnsGPCyKDVBmSSepY94xMd6v3HYO
FfUXTvnwcRrInG0U191Mxe6tbLqxwAHUeKeUiOzGjOLj++vJJzOev7A2mB1a4/8q
O4staxt9rIeNr/JsyuXIsptIzMk1nLd135JuyQwOKkfOSFn8/hRWeP5UjocDjLcZ
XvuxrpoTITpKhI6d/EX7lhty32PBHRo8DWB9euZezPaX4D7QKjqsN6wuWqT7AMqv
oaoTNz+CxBr1x4UTnnH7huSO+2T+rtswLiEE2BGan4dn/8VTfxqC28sKrX1FfufR
jS/5zv51UyDBhgT8v4fVZoZy6+Ox5t1Pe1tOzpZv3vnQeF/jbMnKjdrLnwxYRyw2
Pz6qEMQICkd+QRF2ijkjGQbHrngXcT9PNuqGQ6M2zJRcyny+5Vd9wttVfx5Tqnmv
EyhNBERxIJaQU5N8vAi+XDvf4Z2hhoTd8cNrhJQdF+iYPPqdO4JJiGN6343L7Vz1
6URxpjc1f8en4QbhG7rWRhq5Vq10ToJKgDcJIooZj+Ewcyud5eNLZ/drxGp6GY/D
DJUZ0+OA3SbjA2k88IrtkV8wQquerZeAgO7kWr3RvfvuteVKpGxpXU2xmzu6pXNQ
f2Uou4AVZxFWZXBTxs/fpdMymQ6K/Gryt9jLKeBxollxDWOdBycWX/nMlpQyMNeM
5XxqFh9/49WpV7gzRuqrd/A5+I/i6zZI5PBf7FtVvZchn/ipKh2gv2FTjohD7+Hi
CfKQmrGc4ZviadLFGE4N2AnJEWDVW5/lpXHIYzAeqiPLbYZawno3EF5MQ7rD1dFS
RKPr+Cwgv6B+QT7qhQhmdt8NzvpqbkxwHPTlqu0tdR60fCQkX7ecNJ9/aSLKB3Xr
sK0yOvl1FKIALy8MNmbwzgySsOIuEbRdaEfas0IaajaZBvw/W8w0oz7aD9YhAwTH
v+nr1BBvVcrglRg9o9gIKy/wTpIZDG2AdDBVgncVHDz6PDq8OmSEIZg/4erLXE9V
bBc6IRMqna1b8/Mm6MxxXYM/wnrqUH3CySl6pIbcibJqssDligloRcpKan23G5JY
7dULLZ0cRUbJ8x/8Ho/y4OK5BV/lvRh29g4hVvlcKxBNvITZHgfXJ8qEofVat9Qd
9MjJ4jVjBOjHlHzmBVTY1hcX4ERYRbzpPpmi48ORmamuEesfPq5eFiloSw+c9RAR
Z/OzrI63MmQqRalGMvpzdnJPPxR0VOkhxfo+cMshQoPJiAz+0x3BLjYKfwEOYeF1
aH4npzewUzu2tUVbp/bZgNNq3wMoEAObgoX2Aa6Y53cds69RLsqKC6EkIgtjP1dJ
WI6fJzuN2qh4QvceNkttvxF6WH67ddzNlTY3xRCp4HAclretkbe8h0/x1tSNNBNX
26AKKR1wXNWhhy2R05hP3M6vtadkfj4vw7ePRw2GuoN/NwXeOd1NXAY0eWiwUCGJ
s+d37kmd1X69MU7oMY1Mloj2CYrytxp91lkigRnTjl1pPR3YXWaC0KLZUU3JkfP8
Lax7YJqyNTmSYHaJANmWgMRYjG7hZD7VIka5t9EPHDyIsmUZhO93tQusVQFyUhRi
mu5SADgeEu0bov2LfS9VLvUGaFJGh2ZwuGhpWiNj5kT0bFmqqwXl6BrNiHYEJ0JI
J1UKK5oXXZ2rj6XzHG+yh4M/CKh0l/zHM+M1ghliItRESh3LcqIAHe4SBQHV6nNp
ua6pAvh9pqoHukbgID6iyn64buDptfPG+p1ktInsrwcRWyRLxaN9bNDXV2TIvh6g
DQS67CYFbDgkDmMrxMdGMGK5VEk7ostmGVgBOzyrlxLEHcP2qxMzCnFzx4/22XtM
vRCM9gzj09QNFdedfye7gfxwRSb9KcodTSRWJPpmY1JVqtm5EsrTWNuZHFqcY49H
fMpghj9Ul/a7Yohr/7FnNOUTz0HItbKKAuBaNeOVSQPAQl14WOOKnlTBG2uymDZy
4VprB1ophTt0ETFUzXu+YU+8Iejri5GmymxQ+/jWllXnFSbWD/RAS9NI7DMlTNWr
3RJ5BHJyf2EH/haOTRWqoo1SgZ8mxQsqJr49JjzZiYz6NsEkwbDdnv4ZHoBtdr6e
f/VKgf6kdUrW0fsItp/ABEd8Oj7SPIGA4XZ/ziqZe7Wsl8Ba1CK8bWA/9MnvxQqY
Qp6j8XcXgb2U5i5jzgAZNlU8hu2+2ldYJNcLE3776aXLPL9UipXcV+tpRJjWrm5e
8QrbA28xUszdDioON7bVo/48vgvHqOzqk6NNOiNX9oBUAkQo6ICUTkotc7KFqKPt
pRv21BjtQr1H3EUgWX5ykZBQaDph8DfYibVUpw+4hm1VZe9Txb4ePlECZ6lY8DhC
KsHjlYqLhO5S4M7kMjF9dlMzr/uppZEy4l43xxaX/ODVwn7E+kQJUESR6sFsrO0E
qxu7Lqd/MMeo38WvIJHr4PdRUZo6UmIXkwYKpOK7Nhjc/h5T9iNVh3BluSafOPgU
i9vy16xA4xipEy6QcS2GIe9meAflL8KHTBG21JoME4ebj0AzT2PZRTOdcVeNQ4Bj
45F4vhHG1fz68gzq007Z+4V0a/cNlYuAjRiBUMqyxHolFJV7haa4SdrAHF4rFT9i
EYZq/+1GpEwoUcw9q4NL60waEkSKrI5TGoXTS1JzKze0QcaOz62iCkJaccwFkAog
alWwGrBdatb44ObfI6tcsmzre9RTvOfMYGMvXVvdmUC58adicUvfW5yYoj1gj+UZ
IVtnIRX5y6qRdCHiUswzNnpHLAmsnfGKi6NaPIwMgGCaPBzP47uUerJKD7oMW0eR
sFRocxGKoAc8KPc1hCkqaxmZxtumlSq0VvSv6vBSCwsub7Z50x6+YyyrPTM7jaEs
LuHcz7wtsCu8jlPwt/57y+N+9xbhfQ6IZC8TiPFK0qasPg1UFYowqJf2iGxcsIn0
zbs0SAnjkglOECtnUnrqLQOuYYTd2l42O1t2q09N1MNuvbTLu4iyDzTXCYtAyUb+
DKwt8AfdEi1OWiKb8rKXiqH5u8QFoCDi0EwoIAikTd+mRBLg2iCPbfDQgH9FsdBl
yfjLKITM+VN7JUEaUGKpRLk/geNR2hquFIJ3H5chK8pfEz7h5qbAVPyvF3MdFZHU
eHiJOpxIXeZ6A7rGkQTVwDN6aj8dTObCrAMzG//aRDhD3BogS6uiHtCJQ7sTJM5V
TYNWLbKHR4Oz4hi94tVRaYpc5h0n9/1TMlhNF6eY6WTg9Th0YeDTjXhc7C68AFxa
DvBeLqnWd4Npac3EYLNBYfo981mjYsPbIxwJUtQCG61VTviuYEyR76JSt0aAmbAK
5dPZ/D2Oz+FrJHkhHVxjR9YNm5MEpEX4fJisVvonu+6xMNDPdRU0jeydGDn/L6Qw
HnFrioDeRos27NSWcPQ4XYftMoQuc1j8Mm4SIj1o8SjOcGkPSVHBIKf7WIxazIcx
rJbwQWvHzn7/FURUYCyxJ+icClm6ApUuZ9afgw4rntQeMjeullrZQtl9sZf01/f3
rRi2RiR5niHWm/7NVBKyINqRYqyKS1fTTuxYWeLPJUIzU83OMBCovzWgimV+aSFG
dF24mAYSMXDLUqO1Bub4jIewvikZtq7xKT7UGHdGsgr929wbZGSuuOQy+DBgP8/H
ZjLUc3EarjMgxfWyz38YKGaKcDWbvPiQUlF6CZj0DhUuINP9UiSFGc4VEq9jMRS1
UWLGn/LTU+UaPkKDzyYj9pzW4zBC5U9rljC43MmGk+w7JD+gTPzHxiQe7V+91eCG
ojEfnqFW9rsLgqyRnmVutERRda8JmikRTms/a70UnyAJ6GLxPmLBbYSYAT9BiQxO
s1fhmWY7N93CZucgkjUdW4LXw6q6zv0NxkCOPSsLZsRQWcb8Pm9Kz1IcyoCz0aZe
1YDSn+hcYhenDXz1sedwqcryDiIfRGJRlDxRwUIPvbCXocC4VAbLhwzUMiHo/Ww7
RSAGoppY5QIk3vux3Y6m1njHko5hgGoE043Iy1AihtGTSCOd1r0k7uQDILnNIUKQ
rtD/7ncYd4b206aROynsTu8O4ECOYwVT4GR4hPC3aoUzM6XMqzMeJ5NyKtScG6NL
xPOahtLyeGLQr3uaaosuZcfbFVW/hEc+Mhk7MG5n/jy1XNMIFOj0uoF8girViGXC
KEH5CxaRvlVo+Ruf43WX8jnDG2G8Y0EjSaSqF37oQmVMU3/85I+j1PXxBKl8f4u+
dnDgvpHC9wc3d6j+SBsg/7sMXtNlwhDmAp2xveeJZ1UtS1B7wddrZbanK+8/jQXL
yiXsw/ITUkskCY/jkg488uXxbNJsLfuf4vuS1m8wajlLqYKhduJOzh2+skOGU4Lr
ahwWVjO+gjYDMnC1SXdq4Wswgzmihvpz1qUHaBhgk91z2VC8X9Ht/Vhsvhkc5pgm
hy5WDdaLyK5fW4n+u+q0o5f6FtZBsXiuYO+5oj7qmtBZzOhLS2pKgiAwgRz5Isiu
MvGdrwEaWDLSbsf1ApJPsvt+7JvWABw8JUMuMlm0LCOwEVxQu2bq25nU7CD0uLqU
3mB4DRMdGuq51+JRAJOZ8EyYF/AtBPP16zhM0A07nXafAH8k+s8qZjtlkoRtoD6Z
rCRzvo8L6DMHXV3XFwiCdKzyf8Rtq8nGMKcGxI+BKYyj0l7vFR6wAwWfY3e99BFa
HqqgnThiC/UuPOA0DNpbzMHs+AULWNmOWOqqSZMuGVAuON+NmS2yx2Z3ciiECAJ2
SIERmDzsmZBAtTNs/PL3EvI1WSf7p0G072PWH70DQg7sECz/4u7MgQYRZvw7a7OM
gPdtNiRYr5n1VvegSmRJHGaY0CgwlYuv9Ueadh5NMevBSlJ22CETxzDWfceSadjX
qbTO0DK50qliKO+zvbWMFyGi1y0/m+n7cdELmj7ULVZ4C6HBaPZwHkQpwAIUh8cT
XsekTqygNMUGnlTcaCncStTth+uzhpEwoAhl2tx6g3eCXkpI9vsoMpC9UuCFgLec
FQ8TAObx9H00aMnwgiIhE9Eoy8kNb8G4Zzpk0UAVCQTvCBYyCCX2HiqwuAwj775K
e8SMzUpAykqIjikZ5XbucENPbJaBbmvCiIMiguYu0ZBy8Hxr8ohQ4grmftpUmliK
74rYGbSWVUcNMLibud4nM1Sxx+itY7tDM1m1tHdLM3yWwct7sTCUeLR058ATJQuk
Lw0aNu8Z4ExaALozbJmCaINQ4WDZvd5mga8QE/PHvmK+yfAcKwT4wfNw6ujD3jy3
Te69paEbk32zLzRyCgKl2vSa43XpSIMmNZjTqV1BRLq2g1s5nnOPQHX3oIk3/UHj
P2zASs1yE03051w3/VHNIaIpzUv1YLfJOX4wfDpa+lBMEZN/iuDLIUAacXR0BkWK
UyZIfdp7zgummTH0AbHn+lW7tm0pQxY3aOSZvPF6Enx2oiK5AL3Q8ZqfQXuJvm0T
neDLHJEKcq5DqPQAU9nuQP+r2LTGJGyD34bM+Z0JXw7tWSsqioodw2ygCx47JHWo
JP+/hP/eJtEEQ6GIEx6QYSad0q1toey1BcGgjQaureJSed06+ha9xENbU8qULc3T
biCZir5CweGM80zFFybLhUuGH+7XJxXMA9XmmXhCDjVK3Adf6QbxINz2SyDvuLjn
fGmrKJOzT6m9TsUj9Ht5FvDK9G7OqcRMSLLQKADGaYrAXsbAplTRYo7RaYsByCZv
ca6OU34mB+unljyOalhS6YNw0XC5JY92emftRTg+G3yXRXVH70uExtK4bqneoZ69
so1uctdsgNOm+cAMRUkBPayzgVDAHCRzU6MnU4jkgY6+qYpNKx3pLhStax+6h8yC
6vHBcMys2qPJu1sJDV08CLcBXAaKnUgM79qT1+QGv45dpUT1EAeBHRbUfHqwPkAq
ATe+O5iaedjmjLf6vCMzHlwp40/dH3O2MtUfk1pjRXO8pubdnj+vcI78xGqJOIVE
+0JGir/JyqExWJnn6ndFBj7jWbXMKJ92Trabn+V7Of8bdtrYNhOEPxlHqlSd5YkN
Cj518froCp5mJRY0XBghBCXs6OiuHrjLemCbr/3uVThF6BTyR/DHrkpyFWgByvz5
Slv8ooR4OXo12tRwuIwjDjX6Adp5Vy8MfRWcAQXtSLiUx2dtJNC+uE9flOhTVKsM
wsf8tb9q+FNjKjJnoggnmFvAN5jlhLeTgsh7TBje8F8yKSf3ShAC3j4joMEOVrhT
QDIS340qxQWExCLwCBvZJcMD43sCiWpCCdwDxJINoMHsOpw4CcffsiT1WGPcQ16a
es5yYMAamaqBwo8B9aNPj8JpGi7kE63i5t7FPZK9svP+AanUlrFiVyxhEhgTSK2h
VxSGtTSD+Q3kNaKnvfoO54UY4e/nswdqihDNbwJfpWkCy63Pz9Lbg1TJjd/MF6bY
phw/Ha6ncF1FQoQYa3rLzpp97gOM/XU2Cr3nzDlachhCkEMhyonR1CKRPdMSovQN
PlYOHdV+2gUt683sUrQtT5dLa5QXDby0dxVHzLGYFext0doBf4izUHhkU4tDqWga
wVOW77VcpNEldGBVXcTnkjeAq8NSLLqulxGWvpQXfsuWSSfrzf5dCpL1+Ye4EVZk
ZhrRuvK29HRJQDDDDWpVmaVpbtY5vWBRfwYRdISilCFPfRHekZmNM4qv4o2v3QaL
28kah5AJfw6H3T5iOW4P1zb+yzpMKE7dxVw8fagnLZ6xOVCnHArkIrJWTVRcXRRZ
5XsmDpjPvL4KF7hORnIZGUzBiIFMxpxsEsVwgd4bZEN0qd3kGJOivUsY0CUbT+mt
6YVKJrXQR9hwdO92btqAe526k2KGqm27vC2ElDURdj2HG+DfXAzkZsUbUIzL4LGD
y4faxWVf5AdLiKx1zgMGjw6Xb7vCmFAaq6OZY3ppB05i8UAQ62cSs5EVTWDGe1Vz
iCeyeySGAXMv+3Nn0TvJN5WGsnO4UvIeRC7gRGAAwxCfD/eqcIVbFnJU8Ovbsk5V
aTEUN78+3iN89TdLbm6ynfyFGz+82h9YT/1d2Ly3yErah/+JlPlzG+WFI/3exLxl
0sZoYFg4F3p9XtJayP8nVVhHO70casy3HgtU2Go2m258V4qtaJPthaO3rF5tvBmW
U3ONwT1YEETPp6jXrXeRvoqnDqQroIs6/0LC++JHWsT5/5RaBrV/tbUXvLk5c1XH
sq0q/Ps6Qkcc8Z6kynGI5mchJ4yOuMQwtwzW3BjiNV6+oyKdWiDHlxcg8yPLUhU3
3UFqNJlxNZiow6YUP6Vn0tPSR3eFGxnv4L2bkKgcUMrQNIM1xgs3vHxJOJYTAd2x
QuE1+kt/j6fvbemUbhbJ4KFSF/bt+I+iazlz6OsbSviskoDq1U9Hjgty37LwH34F
H7vidqR4U4mQnCSzDiWF+ES0FXGF20/CTH/y+4+3gc74B1eEXJ0k71BG5dembQYV
wXj2zNDBA8H1Aq3YYyBwi2QMwbqwUgH98g3VmYaesBppOEqIHc0zGhDrWOyB3R0W
AHByL8qQtHP3jQzffefoU4bu4JCEmigYaGDG3CkjplcqgZ0QugbHZBNH0rYVDm88
b7FNPGs6VnrY77V4+aeY8BMWsqVM2tZ717Qp9VubUy40RXZ1o+/YzsJaIhiX3eZ2
29wEYb6gvwBzf8GG+haiENHO+1D6uMEkuGuC1YfmzJvcmrXdHdx3CapQTpUZNhws
TX4taNmKGRgvrT2Q0U/QVfN1ix34gxs2lIboxfCzxeuUFyDmPjYUdwGhQC84ukr3
AwS9ne6eY49bnsKbFoZgLh9d8gsKzMkLAct2Ywad/RAqeBqDwr53mPxSqNkeiqPr
eu0aNkh/Y350m8yQLlZXaO66aYOUv/J9AlPAYzbvlVqhlp++/qCLBhvRZoaC7yDe
ErMydbsRJ3OpMNLlRCGKfZoAErVKJ3/vJEhtBpOkWyohJrklsjJu+M2JLAI5JKt+
Zxd71qLyyKSVUz33F2kAbfAHVNAp8ScnaKVIwPDpK7JxCQNCD/eEEGvbTxSG3ke7
w1raVXKByuNhME9y/EWzJuuMsWqxMbgHCILSJ8sTTUHLEs7FSNUB94CEm57mPrk6
azbPvxjgNQN79XZFG0YDloQKuxsBMzwrqVo6rt5F4O5dYPMWPXBUFS9qAOHpwHvO
rTGVSWXNilslaw9wyYZ3yNXRvbYD6v79NC9iU/+kKpX8QtZ8ItbIfkOTjJBngiZJ
trDxU9hh928sT8FEXgOERJHaKnaist7Tw7jynyYHc5hhv1wavbxtSLv2QzvZQTI4
Pq0I+zroCL7uGYF23F7RIRc6kif08q/siP08PdqIXSiclX+X0MiH7WZiK/2LFtc5
0+zm91RcEM+E42+D+IXhjpwV9mLT9p6gelt8S2hQfeT9v3vnKOoexbKEQpu2lHPP
Dt/REr76GApNdyZRiWZIGQcySicNhwU3ZbqZCrodVUqp/gYvLGOHBju84nNhnch8
5QGPjkzzWlcUSRvGEODRFBkznF/stA+JTrwWeK4kWysY4skp4PKxWVSM0NY+YMe9
5UWVbsijsZmLX6W+3M4/Iz6NVcQTfo+1FzjTkyW/hkg6qe9FrXwsPbqGDxx/nGXP
sNcyh/vFf6KMvRpOpI5GDKNyBKeXO4XbBQoMknA9f/8NCcpVS66Zk/vwLQgVTbs2
8v4aDnmA12YB78PLW71845eDlFxQwiJCNzF4dT2WCkhwvMAlk0oWelXS7VpYKn8K
J0bCfDEZHXUjNh/8WwUIJ5VNT3em0pTcMi6m1eeyEZHKQ5CeRwnrRGjti5jvi2Cy
qBehQuM40qaVcxetA3z8xrXEy/5gpoYqLcgFz7dGfQsa6+uncblm+lJzIixz6s/q
GzDLxfdg0S5j9kHapGgY7WI9g5M4JzWOtSaY+Iw7MXaa0+taTS8dWAJ+SbWtzmxD
Q/3lKfTqspaTK4zIjxGhVDseDj3feVEq2LxYrNVCF33SQSi1bka7SzXR07CDRWMY
R41SpGUbOwykxTplJ7u6Pof7kkxdNINDadTO8aK6RZBaChuhq7gYzGaDBoBB/oM+
nbk7tBD9hoEVZV/T6sE3khCwMkU6+45JvFtMdxlo70A/3AlEty1MqKQLUe7dCf4d
TvLdrC3ick2nqv/PuC1+IO/HWO03krKrwJX9/hLOuhGwkJ3WqZ4nUx5bSQOVcGgI
bu+kqsNuVg5xQ4mV+BWL6QNsv2d1Af1KN0u2rNnQE+PZybNm2HJcHMo9Pt72bBYM
3UE1zgLNXeK5DTpGXAlZuDKxNRJjMZEfiS6gAgDeyyCR86D3SBKimGubjWH+x/FI
4hLfpKN7Y+3htnCvzLtX+N0LcKN0sCShFWKjZ9gv0082Tzc5JaMkWJNNVDWij/yK
wpBJytf+ew82qplNEY+GQmkEchWuDueaIvzXEoYTySPi2/YFCBJEBGR58HsuXW/a
OoF/gQNUrM/evQBTvYDoZJggtg42Dv4yYsk+vGht3B87EUgho8+doBazthhDFMAB
C2F2hWRpUqmL4jkEFTq0Qb34xhuyYwuk6SxBq504iIwQCE7OQiIHTNaEcPq/0CHg
J8VQSilOm7ms/dDrcc5w0QtFB7Iqlfuce6nzwKxCkZWWuF0456gTmtp8yi0Oxk/0
hctdyUSin9FFviC6GhONIZyNpfqxAdBk+9v36QgYODGcdXzNJaOmrcIAOW0o5Cpp
RPH5NfHnZGnTsviI1xLy491mZLYAloej0Z9wNwe7vDs0p22RiW668LUHRZrhp6Fp
wMj1o+Qq8vbBFPbZ6mbCRV2XrHS5kL1HqJqCBFbU20pC2VD7qFc1QZs0U/DC4AqW
y5hP5YxUuh9FhbfKqxfTzTc+rHm8T8wqTisXpCrum2RhJKEowb12NySsN0KhzmO6
NQWDo6/lQLysjm5a29XXLRV7B/6k46UpULvtNl2PUy93ZF7DKyQTEHL7kicK9t2X
IdgYOh7Y5fp0ltYJfU4piUFCG0siqSfEkxHmk/Fa/yZBO6oPgaa3hpQwLs9A8Aft
/uoEbNTOR+nuGOWRUMrHog1CiUZyJnYEfj390meoW0PH/O090zt1MYXsUMIrcNDq
H8Tq2RN8o37H15hAwctuKnhefMldQANe4PC2z6nz7VYBnmNQppEArNKf2ociX1/o
QrL+I8zW0kD0taRij7acp0F7zESUsg+0f+dBPjUf66ekQYivJbwRdBBF8KdZN4+7
uBCqvVxlBPRhFUkchVozwQPZeBDhwFFj054itWTkvWAM4n6U6E0RuDfYkBIk8Oa2
wxLpjWLPvFOVE/h475lIWVAb8AJLfJz0j7oEOOY8SUL/kGWdoB8y27Dgd2aM1VUi
A7t0HTL7/pVKhTyvEHQCgrH/RQBognH1BHoJRqvZZsxPQha5TaZsb+2rrxUJ+srX
VQCnGI+HAl0kHrQIFmSq/+1LJNA1wPmKk8eEdRKzNtNS8NKj39M65mOlvuD4o5Tf
WZMIwKzNA7xdLbNdOO4w6AbZOqGfoSXktP+fYame0JxgW7xrdURA8h57oBzNtG6z
9RolYiH1Jz3P1C3rnjbf6epU4KOUfW4xSUQxrLi2eeSUOr/8R/mEQbWSjxDDCqgj
oyTCvtFMAUwblN+7qgrlenjnOsL1HISL5qxELYemkVa8DwStgTmOHho58/y4g13I
G5irB/TXN2rDWiTEgkwWYGdeQarkVFsPtNqrmIu0SC3+dxzI0NWeHnzKcNe8bOXF
jkdb/9Frqr+QRqZgKMrv/ulEISgym7bDMCYj4jzDP1J10EFK977sgeHeuP2h7b3t
M8zZZ6KnDg4ZQc88zUmXWEtHyEAVaYFjzr3WHlhxcZMnlJzWdh+mb+/m/ZbOYyDN
l57uxtdGURRMCm0UaXZJT1oATrl3lf/ReQD8VDzSk2fcebLzMs7piap2OoVi9+IB
vNCgiTzL9jFTJ8ARWUfwVgv086jDQS7zNytDvW1udqqtTbKwKe02aVPupB3iPZY7
UtFqCb/J2pStMPfl1EVgkZBoZQTddJVQY+7TUhr//INkHCS1OknxCqNfeaDuVX42
vj1lTnvknDpmOcHZPCoNT8XPMfV1iBehd40YAPU+JUX2/4FbngG6htAx1MHwnv96
50JxO2bHNY7dczgTMHhk6o0By7DVLkrkDB+XHzE/eAhVm54FUG3uGy4ulZCLb2zI
eqAXm5wcLpXKoslZUx4TFc8p0pCIg73ANM4wuN9rB/9t9bOhfCnRZixvoaXKIQUv
a27arMDuFlmqXP8cKdN5AwwNMxUFnU8n4yk7/Q8TO8Ee8bYA+XGKiSq0Ol6ygsTc
w3qYurrl4656qwhRVFbQv1iGCOI1oaWo6+n/E73nM4Qu3faFAfVl0B9Cz5+bSJ9O
jpgIFhJCrOp3UiwsAehWDVcLcE9GN6Yfxk3TM5d+jkWF6BOBy/nfv0LwpskI93UM
ni2iKTzG4ixFTuhyJ//PNwN6R54rul2x3VMeFBH0oP7r3YDt2ZxyEq/igT/+LdP4
39yS54/jBpqsOtxJY6Ko74opMqtB8LsCui7kAqLIUNfHgYRAFSmmbXmruHKp9CWH
0Hd4zcl6aAt3zukKIUB2wbEfT1FI+x5xF8sblMyEJYNFeSDWLB+1BhWJgl8KuIyh
zY4rF+fQcEq6rw9S5nmlhALN7mGV+0/0gvJ+H5hRsTJ1KsZxJcQUg+AVxmznxNUb
KpOvlxah+5YDgK8/ir9yXrS0ng18yK6pASqkEkbFSRQAh2pUSpaKZrxLv1OL9+no
WhQR8Z6J7NW07kv484mbABzJsgBY9cuGiwLm7vLpLNGqPNPn3Gn30mmE50URUJKH
JiK6F/Fw2zMW8MhTOoc84rzjkkX0cPgr7D54MMwRQvGeAdRU99pxkBVQs7gTpLTA
dd1bVwV4uwNKFWFgEfpOW0VWoHSR3Zojru4BcT2r24InHfgEjJHqNsgOTMg5nGp4
JoToLdeX6Tj5OTEFLhoGxbmntep/GAUwvnpyIU2aQ9+mmYfZ9GVacAa8ZQShbOX6
WfdjYZWdbMi+93mrE57hcgeNxCbF8OUTrnBJsXA4SACbNYYtA7gyahQ26pXyOZh8
dVWTZ+s1De3PaeEPKN8kQlvZAtpS1Pr8pRd4LjRYVG3IPgVnjNDyXyQpBUCdckrX
u1vFgxL+U7u9GlMci45rPVaETtZacA9RCnWE3rOenpxPVMHhQeaisLtA5F3CL8ln
oE4zJvTMycYsPKoDKoFKr0Dc79x+zV6UEt3ZA7I72U6aVffRuV/E7BiGDoCOn50T
LZ8axqsphQxgw5wvq8aerQ4xUEqebbH7h0E5m4trgtExOyI4Axu1jeQs/1WCDESR
quzCZqRDIXODp3rn382dMaotALEJ8npMNwaM4t96V2H+9wZ+yUs4xaW/J3EeaB9q
YiTEI7mzVJXfLzQ44y1Ig7EHiGHxACd2uJfTa/G+hb6I7hthuMHbSzIXin6vvnj6
XjKh41Y8pUMWCnQ0kYmZCA5bhbXiwZC4f+mMSIVAbSAdCDQC9FTB4srgUUMjBS3z
gn5nfNp8BT5ieGkusXt4nXzse+ClvymrR75aKt2ouPycvL/wui6+c6XgZoiyy5Zb
h4fVjtHUVrLGPWs3hDU7/Dzu46EMhMHBNX/2q9PsQYfm2qNcuhtFItWsg9tIh8q3
0Ogn9rI1Zmqx9VhGc/PEjiyLTLWrvUsEXhCg//SyPiwcglbGc9sHzaUTW3TentMr
7LZn//jEs0kA+vGaHAbXVPQVnbV7Kjik2OgcH57Ryu6rpgQ1jemy7PIzk64VfaPn
UrTjLbgNdPB4QrKNt7DvPf2bQbkoeCLQ4P8C1yoPVBbpE9W5BEVoynFWLz7xyMEg
q3DAsuipFe8C8K5wCdh7nHdt4kW4YjbLb783dULsLDQKsEEC/AedfuwEEmQHqIAY
J8Tt/ycXRJzurM411kUmQs4nsAr2NXiGg2PHjduyJreDjU5yZYcXcr5P8PME2ygD
/zIJb54dPJFEC+f4tk5NcYhubJ9tYaOAX5Ke9qB5ocfzw/ludJ1meVUQcU2Xv0nn
1xXQpIUbhgQxFhzqlfdWFFrbg+1jf1ktcafO+9pVt0FUsJpJOmvu4ObTIdPU1aSE
2Br8XKX3V5F3MODwv8b7+IgaHE8yx10zKXUcbOciYXI/g4w3WgSydzeDuqV/toC/
5CpL334VPGfPQPmjdIuU7TL2L5bhL5WxczaFa8G65pEpV7Q0ZmwBZbXENVjJX0rV
1ptK+CayNhIDR2PlwmTi5bCsYlq50nIWMHASUCRLRJLqQqCSVO5TnDNggcab65AP
Tqs4QJwReLvp0oRr+STVTpg5kpMYIvf7DDM/g3jc5ZSIkT1huJEk8o3ZouQCI/Xh
C+nFeEU8vSP1rZVxcdHyF/KhIE0bbE8c32tyveYRgPCWEg7zF1PeIgwrjozoc2W7
CTHxL6VQfSf9Yp1iIlql/jzw/0WGgbLiH9rzfE6OgHwc/lrygBVP5ZMXXjWcf/+s
O2o3acYhXrf1yeaMZFe4Z4/5JfeNXgQEhdD3UMPvxLWW6NaBZMBbJk0D8XNqjRje
xpLemRtqRuQoFF5sm+NIH20JddLbSfDo4ALLpMSB7XTdgcaByI+HxkJ1zIR3NOEg
T6K0JqYezrH7In9vC3le07g77iDGz6uvojguMQNZDLnPlMCJm6WFO8RttwW0bFqN
WUnSA4vayvQu9VvzS3gMKT7Q7gTOsadxDRJlLgNT1qsV+IUS2PPG02CAarh2+CEK
hzjj//To5WAda0tss/8x8mh++snQQueJu6/CwZsIx0rkOHctdVuQVP9910ke+w4K
5fY0pyYHLEIjVJuN1gfjpHfptPvUlYHNAOYPCqXdoazP2NZjtCkwzM+g1oTBm8SK
uxseD8HjkmDGreZSfZHdJPv+0aDreo3+ujCZK30jOA19E/rWnAq6y403UX6KJXuG
VQndSLvq0Ey4VdZClkmKxxGyo/h8Ye9m7uvoPSW4jIAEAncIWdiG+lrTzd9RgoKj
p+RDSMZWt+HXj6WjpwsjmRuSKhL+PNYOmif7IiiiDo6l/yQOm/yT2niOAcS0VuR8
BK58EpgH+OjJYOK9sVjE3oJN44o9EH9ZtTrxOiNgILg2uho4m7M2GIYC2ZtWgDh6
JOyihJAoUEeYrGaG3IjXss4wZuVKdhEVhq8j+34sMKyKjyYoYXqxpwhv2XJWI1tR
8BM+Bf5V/x0gdRk2Tf91N/fpNJCwyqfgubLVxZSBUG0rM5wu0RGjG3N2a6yVe6Km
M7NzZ82QmEDoJEW9Nem3Fsbu7Nax11pHvE8TM64NIhskUKQl7QNbJTgsjiqVryXt
93H1n3UAmn/2kzrVHj6ovG1GB+MXb1seR3BInaR2YBJMfAO1h3vrPTI6UsM4FzFu
4dC/EgaEykKjEu5JDcPFwVWLHnzoISuiCRPzqpqugU/xE2cATEJTpc2GHXw+zRcz
ZVZIs9M0SD2mx0ag4t26ZIcFWWkX4+9DlskrU42zLnr2AsGBw1izxPUYBnAJUyGo
yVtDe8gUAE8gai/+dsobxCTK0N8XwZGJ3CGX+B7FmUCCpn61L6pGkZiCQXL3nbGm
rPx2IvEj9ChsSnBCDnWAiF7MX5tzE/bmM37sNoqgdQI7N//ArOCCT1qAIAz9jshn
F20NrgM7mTL29/TpX1r5sxFV6z+tIJ5Xzqw3oZ2vrJSaxRblascjm3fkJY5KcahW
XN5pqDzw9RlosDBYtDIFMad/6LhP/s1AsZJxV9G7ifqXGyq5GNyEZTvoEW4E6aRf
ZQixAOwJSQD3IctMVB9AJX7aXMCzBeNbNRkCfJmUB/OAY4do0JJ4x1JjPAhb+YWY
NmRpH86t8srnYu7GSfWJmUZp9csXGM1/vGhnX5NpvYI1wB9GRq67Wo/45ic5i41c
Vt71yHlz1gqtVc4iVJbiR+OXSo3abyDG3+qYjAHpJWuancnmm8AKKeaHhz2Qu8dk
o6aPi1k7mYe05JdgK5EwrYPPnlHkPxdgYMeyyUIafttNSy8EghTJ1mcA2J4zng9K
y9hWmKW0/g3i1II62NDvVTw4CXQwufpoRwhRbXdFlJUGHWjt5rsWLqvY4a/xXE2S
xKaCvwLHn9HfXqrJxWqnBlWYvDHgDeOdvdODM6Z5BrLI+WuBDwt9EpHwDPRcOiYA
kWhQCh9Js8F5//pFDpyOypFMv00MJbXhPuTJoZU5AhSCi1r/UQQEiupMcOvIzwhB
lszalUfwv5RF8QzamhoaNRCQmhwAC3FcW30rw2cmz6uupl2wRKEY+rLVUe9oIZA7
JINvq1KxIe7Lv9s7VZMuKuiPHxpF5xuSR3m6XxIXTHCpzv7VIGwU6CiDyNQJL0Nn
0haaEiw1a/FsEZ7VBXmW39mwQEbCLK3P/3k70xoJ+jEA/+v/J09JhpF2Y+HzU9ci
tdde5kz7JlsfRZPVO5Ozwl243q4Sm9oRw1DxBzRuERIwsweLvbnvuKhGYFqZPAPd
KEFHh8arZ13CZ8KkuJeBlybLun2lsY/od/5o9jRKLum4M/QnkHrWk3UGlovtwY8o
kwMh8WSIMaiKYysci3QghSyfUj+239jqv8XQcnmYfu1yTltM5tbF/aOuIKhZEsOQ
OrS6N+X+ayNSLHsqlSU9RXXrBuZJn0UozIHeZ/ZwyWqBGymoHCmiw7PFM8UzSfMh
/B2WYiGzzoAoQyQHRqq/woLnOUUWpaTobPTtv3Vdr05tN16kAkFkoDocilmJzSnx
zW5ajQQ6hJWX5Hl8Xzg1dSlRn32ZIS57h8TiMqrH6gAdNhry6d+dv1uuOkAFlE0o
CbBtDC+hj8uagKCRTCkBervQKHIJzlGC64iPOXMSa+ru/wLxsW0U5vYWftkURfwN
dt/bN/pbYALl5Md6qfP+qAn+pOaKMcXyDXtJWyZjbpsvzLJ0M3b7vaEbqjIR3baM
1c2xhgVH/WOwv0mr0ALyEgpM3JxVC9Gj5QLf9XbsPgsbCbruc+k/HNagwlz4ksR4
O+nFvGBZiCAkor+b/vrXdr1Ie1a5SGsLzWYfay9doU9pbh5cvCsBB05vUT3mGfPN
J3hoxsTVZ0T9uOUzLRCATNsu07PzD/V5QT3Krlf719zUKMWqk4qiR9ZJ8KdVyjRk
2x9fvD+LYroUQXTXN8HreGXV6Jv1LyJW04JkpIq3GEN0nAHfSSf7W27k5MAwttqu
QRyZUfneYn0L8etX+hJ7uyFq8EqZGuxvq8/z/SlOtGHgiuDozF9GGgLe+oF9U+5R
ccjoxRC3JnxwBRpfe9VeMUjvt8FXHfNQs4yeBV4DqZlbdXpXVSOUfplgXXqUX9rJ
y6Ey9N/tiSExpL9+KoFBhbNzWdQyC89cP/RLbmPR9urIq/E/ITmsoEHPaj5XhE9m
1xeVpqhW0RsBXsV++BMTG0rxl2swCAXzQdCnjOPBGii2frj8wkS9YC9cpv0nqVQ5
rZZv+dOw+HHpBKqjzUPHETJPRfFQoKc64cbyY7N5F1o0Y1vhjNbfT9ZNuuVby8Sc
sk+2A0Ng+49mw7VMUGPLka+ByUshhpSTDs5xQtzzrivuxRA7aKQ4Bi2mUt5afYH1
3HZUIsmb9wU3KUlDZLZdSRGskolarZVAN1TU9WgkbCs8X2DmRP01KRr6BEelF1zB
J4ZVM1+fz80F0untetQ9Z3t0FEpSa1OUi6JQ6WAIH1uzHpqn/EbWsvJxIwaLYuuT
yt7jb5bWfBYAp1710CA4kRfk21l9y4SPZxG/prOjqcIYgNDrqlvO81vFepmCPuTT
iQDGXXfOHt0SwGENBFCJKgR99uPl/HzRso6u3uo4qm+ndH5I5DTOrEaynTjjVwlo
iYvJEAzXv/FgkRnQ6vmkHKLry7ZIqht7kTuggUAe6aDNbK72keXalfWbyPbIxQAV
uef7lst+nFz3MsJvE4p04DwEjfHx37goINVsETtjt5h4Ogkpb/hFMoYYpejdTZXn
E1UuRoFkiYy/gRCkNObIDqDPKx2MnQOQ2O5aKs5p/Mr1iE8WZ0jUeei5rHZvLmME
0ZkB9wTm0uTImERNwbI/zqaiHDxQb73ltPLCzBm3MBIafb/pdRqeLJoCtsW61eej
R/A+e+VCOGDN4qkoAHWGxqKU48UIMFDhg1WLehZfUoDxyLtUAGm3GZax5J3lt2d1
jBfz/UNzHanxd6IXNPHek6c59KXxBVyPIlL/MkwgwSdQnzf3T8hq7C4hlriOUSsU
cM+9sHhdXYFi9+NEYDVTxJynmW7yQc+kpYcXIdFxY67iOi7JTlS657j9trB3yFoO
9cfpuIRvPcldalfOh7SbMJaowxDWXtgH2iP6ORT98TJyTkTcMbSRlcBUZRYk97Db
oId4dzrTMRtw26TgCagJv8BrKwGz3dtskm8x2Vw9SNszaGcoclRqun8DGvwPgnon
t+fjb2puWBowTgHOlfSmAEctqlSFx9D2yPSJf+JJBjGp+IUxY2249jBB/zB/W954
NJ+oeweUy8xiX1pq/oMVBHYE4IMLxnioaPDYeFzarVOvYyZsPtlKbMZ8Y61zvYf1
YoholNdhrxGm6vs9hrA7SFDBn3L6c50GqBf69w/u3Zy2x7VUo1muwDhsqFpD32So
hLX15+Y3Hh1GkZtiwHobfwQZ85QOS8dckFt0uDH34efezIKYJN9n82GmUlt+GiPn
foQUcpaaRksgLzvEfjsWCUvd4EDWGudI3Ib6+L+8Xk0U4dEB/EgiM312bX3Dquev
mCGXHKuF6Kz9WbMNbKBeT+zo/3TSzhSZOI6bOrOKSPLY5CGjv1H1szvQlnQGJu1m
Mzbn5SbZwfTc/TwBb/0uIs2RGNekiVkOGKuYEIWiz2z5R9i1NepSOvk6qSg6j8tk
V0FWHpC2F4WEY5FM+/6LQEaO9aOgQE/Zh3zfA8B4ms2FI5iuoz7uCOEFAN2q8y6h
LvV5FjL/ss8cdUFGGgvkAlDhf3P5kCSRSKmy83lnxCerjy5PyEyV8qEt83G2Zof/
Bc7WoyzqrV+kG4/R+MA1qcsExmF8N6gHQsDVOlVyYWeahz3vF/vLKbCEJfKlOJvn
20lKzr3tYvBGvaOWg/8HJOiM2n9ly4c443KRaeh1wJJczzWFKGiY+KGCjzBy2cV+
Ke3dRfzYDxuSNEuHiE3Z+iu+eEI+BWjkVdhFdTC+vXy6SUaPEuJMR/5aPsnwp0Un
Ejsaz6WNYvIIHBkhPDy/XX+jRPaoGHImdW6TwVXivXbQJOlXQb5IZr7WJ6ezJzmC
FQyzzbYdaEBi/z13/2bqDwQXLxYksaDTIUBVBw/T9kkPDdCzsvfjVo7snL8fk31T
7QpTjAUhkMQUK96nLIavzHY0m2Rp0N3mZDwBC2hF+IyNdvnZoEldfw8UWnHkKM+B
3b2jmca/zVBUn8RW46AooYXWAirzwhFZRw9oY9l+PacRfl0bFvC0uAxyb8mVQlij
FPa1/osa3AOXkj/lBJb0q+kJrpMNmn3Yk7oFnBrg2RoVAaQcd19E/vfQPkQvS+CK
aPmc+zWCn3BDfMDUV3l4zXf5rPLW/tjXUcQkD3fePaM4Qdu787gFf58Jrbzvysu4
95BVF2O1N1jbW2ZbUTJ8Qy445EDhTO+ho2aNksaKntjEbKXTPHVN3VaVa5GVuKHE
DrSaRQftG/2raR4+IBoUMZ4uLpCCxCs8VLPTTsFz6pK+YZJBFiPkdBhw3RwFgf3E
RYaQ4q8zaRTZu6ab0t4mm5eIiylRqR48PSh+ZVPYpENNJQcVek432kfPlT8eiNU/
l0vDp/KaW6y6gFdJBW0bOARhwUpBjIq3BKhvaZb5F2cwh2Qu9iai/QyHZlO9neI4
NXYpt312/r+Mthueegt4ozI+2AjtiXWueIMdGtX0u50+yhSXjzou5aEUtcI4eM3Z
/qhG8+cbZPzY7bApA95Ti7OqIUd8yKmMkLRLcdd6phxQzjnh+qD6zr0dwWzEOrPq
OA6GZJjnqcy/mAY1PYuKK59I3GxT9PRoonwGjWe7mSs/il1yXKQf7xPN/++JyoEa
lTzNHc69pAYVU8eJ7L6klJwc3qOEoXYBCtiZSmBSzAYmcBUxNSCTHgptJfoucHnq
nFLI/O6uZpKNrQTObGVEVjgNvkYqeFy03i0JUi+pPRfatW8k4CYDdDa38V5bm3pl
WSHZI1Z1uUupByAq5wS7wef2ecdp4dnhL+xA7OmSwMrH+B5HBMv9R+LLbPl707j0
rGf9W4qIXxzgR7KZWk9WGQ2wj40JyTfCukj6QMz4pCXe8IEkdUqtyl/HlODnIACq
ECbK91KTQuFWZP6R1lAlKTmuPbUPSyo8QJcRBuEBnsmZFV45YquXi+rwDFjC3aBs
ckUpEl8V/qvfA8T+dXQbbrLCgqXA8G4fqXjl84YNBrh4qyt8f2wCdEF6A6ucvNLO
iDK5OfErIh6VFHL4MaLhfYnI4Y4HqYITiDapzA7PukPNU0MwQsQEi920PxEZK0/1
mWhppd58ZxAp7Tjzu6cbq38iaRE6EDXa37u2Tx6XbD4QxXPP82C71DCDMzXP7QwA
3ABMEyTEriC3cycMhcq2ICdYEaxUItaCHGmkU3ccPLcxYq0tt3L2BsuW0KHplUqb
w/GUF6DLTvWw83ZuNhl+VtcelghHZXRyA8vD65YGEcCOY/dykGL+6d9kK26aEDxT
UY5rnYdtEZO255cAMwUtliBrjslKPFjNRjpc6OjtMRa2swKBZ5VqwTbCSn13IF1S
6pL+XU0SKRvCLHSsyqJDry/UGOi12L8FUSzlOS2aOA6AyVP4iDrXt9ZL4VOa1Bxj
jzbVuId7oBs8PF9fgxvIfRWTAL++XEQqhgDepYlQmRjEcerQ9EusTzGTB8bXi3Um
E9SvZ8J5/7Al/sbEailGY5+k0JBylV3Wuv4GcVpkWOOLE3bn5qf5dILwzTC+2e9Z
b7eC3rK+we2OYjphf0t32iBLqmmPKOcz7zgjiR7ZT9ol48Wr5CqH8NbXl9sWhRAf
v1/GCwP6PrzYq2js3yA4KyleB88fs+Sxud+V9W5JXU9JXGPUbie2Msmn0FHeI69f
+KJBSGVo2Fo7ODwfRvtuXuWOilqQhZwU+y9wtG432iZWs80cnUbZVsTyMFeFNwWX
6ZrI1SUEAlWnjvjomOAZfMm93xXEX3RRD7Y2k24QclKf1ZX1OcK11cmgBc7l9TkU
nNFdLszn9EzGHCGq4t/Zp9jLqsyFOpdUv8irPPDVYYeIV3OhN3VjzXMd6QvvokVq
W1oyD/YuOhi+zNim6IGM+T4gOlSvK4eqRHIhkpvASeTtWnGaIEorUw58PbrGcDhG
MtWe73PL8A/6G5Fij+20l3lErl3kHOOO5I8Aqbqo0uyWqXm00DCn9YMyztK1Uff7
Nq4by+xJsktE5j/NiuTv42WdMg5Bgi100Y2WoMe8D9oKLt/rORQsuz3oecfstJot
LqZ7ugOTazkSiD/BJ8+YAYUA3VMBe7DhbJ7VdVZARqIy4WA2ebCNJhIzkWrAL/sM
mRSQmo9Vos0hBkBF+WQimKseuSVJ5kefHFI8EdNTwSrWaNRTzoRr0eOr3owpgI4/
+772MDFzV1V4tCM7/2OjMP9Mabm3/LQEDnotKO6Kq4m5T7WaoJ5YRj/EnyrtKHOy
KsbInz/l16NDspiLlf5TKxRvyhVikfQlFD2ZiHw0VKK6vsdS3vG+d2t0iSElp+ig
JQ5v/fcIsYaRxiL2wPZGaLioU7W5TqcEeGjivaxajbgHXHbbAp3EVBi77F7zVLTb
NSPLl3j4MWz2autDhMtH+m2ihRvsiOolltAOzd/8k33d41Bs/++n93xbOd+5IjMl
E8IoJ9Omohk/4A/PLA2QqBJqzPCHj+zRQ2Uu55ZzjLbEKDongCLfiJgHuVOgA7ff
exl1+HrCbgNXg3tU9PNgEOl1vUXrMNNrvjw+3hpFFc9/EX6Ji9QqB+QzNS94TJEr
eBfY2RRKg0weib9lHrC3TMzl8LQcO7vfkuNEDnJ58XcRgABfMZpuw/r3AqEjrr0j
NTcPnyFvx8LzLPsWHVKTxKWEBorgPBxKI2wCzHhCkcMkTNL52xhbm0f7ES+8+588
9yyJZ6V7cWy4BhttsR0wyyI8WYh8IpcV5h9Mio98Gk9N7R1sDbRt6vH49Gb+bDtk
FBMieykhADGDIum8fbgnY78OA9pEt8PCt4/as5IoIwSF/R9wWCBiRZu2aZMgQ4yl
dLoR7UqAfwyjmeXd8XpjOw628UG0zds0C/bx9S4cPyy6IvUH9Tgzr6jwcQ1srvOv
O+AXAXN328exen4YmyEMjNFHEoFOMfOj5EEgOw8ExpkdFH5bUaUJZ1JC0zYD5QdX
94m92m2RFVlEnUt9O02PmxrCrlMopvD6xgd/iWVvNF62fT7oPlMNe09xbqlrgCfI
NTCRVMHXW2B2nyVXx0ooegNEhHKMyTJhp+R/bwOqUu1yWwWX9k9sWTsGqveidQev
lKCSv1IfqnOBFbLYaGC+xkTJUzMtCSEA3j01PvgRW8r7Rdq3qx/sjo4fkSy+ggCO
XxqclchQDikH18RE/V6V0W2YQdLLMgjYtOAEbTrTNe3ntiypMa4h8NbmJTQiCZcx
TbBQ6T2eyIUrSIrLW4O7/Z0dOiyaqyKv6ba8tzA/0t8gBgmE6BlfDnPDqgzg+UQr
5BlILQw9exImBO0MB0kcbIBn3ppYNol4zJqOUxtIJwvW6AKUgT7l0P/OcdQZhiH/
Ht/QC0Sens6kjmnY7HwX/1jSBWiMbqZofCq/53q7kNr5XGWnkBRmN63IL67VthR5
nZUV7dYXH+Rweqq/tOlEBghT3dxt78ITJrXLZ9gSI4rooTdDxAmxmxMDI+/TI3Jb
4o9r9KhSSCOpnlDXk4QuDi3iwaPB8hXzRJJPpE+AFWSdLCImMt4xHOBABo+1zwk2
fJEoIofjkEcRZpN+1VbDe8331pAC7rgMrcmcQ0sBPZF8W8chSVbO8ec1JOHm4Sc5
cYZuR9oZ2oMAN3o7/CZx63mFZ9QXQi0nc+WRdkVjDVrt/h+Ao6UmQ5YU7X/QQeKu
MMbYkol1+rf6c/vrpBlRm6OlNPXhyrEvkwNS0xUA5uztjKkifrRqla19GQo1MwVH
9l8ZtEXY9GDk+4rTZMy77Se7sBLecPQI0pjnztErYyY2M54nK2kMjT2FeXWeCFZW
X3f5tWUdWlRt2nrioyeoJlAmnVYtWGE8CkT3agbX4xVLAUteOlEgmxZPZAG7Zx3i
FVux0kiSY9cmr+fz3B209gWoR9ZexscHclciCIivmf+rq1dcKDmDyNK8lU67WCJo
MiMoepyMl90h9cve5sm9QaJRKOGzAydIELL8fGL4gdtHRuTI7/toEXz6M3RBAvGP
9t8Ovy+TDXB2SEd1E88HhjQ2mENHTZ4RNk8RhBJlfp/VjFXDTmJW1hSEosq8Vdz+
oViirYR4cL9bd/ZThJphJ27+2wtz9bysvKg/O9WiYuQAvCI9tFqZXFHm+cw2i9H3
pAWtCaFW5eAlUzoVYXbW/U+ghZrY5UYy249A5t4/I/fCJyI4c7KFEJm5meL4grTc
8tEh7oPLNTDLfwtiT8dTnmFUEzBevP+V5lTSFG3+I8iq1J4ZetK+3mkC8HJ1R94X
B8c/33zi74Bs+u5XOIvgWR4hZZnqLoX4t4Mfm7pVbMFqhmnjntsRqNwS2C3tQOhN
bafrrPpIfuNE5UT7l4plWY/j9+v9dw1nvp67jjaKXDbC4GdKq+lZftXeHdqcx/Ye
a+r+oDHuqtqVgPAd++iwpN85E+Siqx3h0ke+6PU4siuV7/WA/v3vf4PRDmZd7cBr
3EM5QTghCQK+RG7t0/nEA0VyWsXCUdVA6cXi+UEVkHN26lgZPNGV7w6GMJGjImPf
O6AzvurcZhpDub/zO6Ri1bpnpLZ19/yGN13qdbRzH+9k6ybq1arsIRwuyQGo7HxH
A1gDPr+JwYae0rJ2qXGXEJD8WarNZOhdTnQed7emrpmn+EEUGJVNXb0MK3GmH/MC
WKuOWp0Gfwk5YrytLiyuNk7NivBYeP67y6DhHYWqU4Cdj42EantaWjOFFWg7GX7G
Ng9ZDXPD36MU7ek5Ofzva0u6qjJ7w5E/92EI9r+7DiSY3tjSA0pL1ugzPhDsSesw
nd0+dLVvpr+Ah4vihkYk+L2799bfYJO9Af4E9v+Zp+QyrZhXFIGu3hOsS+qwHq3Y
FK6+7EWRkjJIGpQnlRhJgKo8NX08LanA51OtRYdYTWNtybjbi0w1ldXUznZ82llg
0OmB5VYx+ejQv0PgsHAdp8XlM+THQTzXSNbncXEVCRaGxGxaU2Ygcpi1aKfxsIdo
tXGWdsPsAgjKZlQpywasD6oVaKAXb7XlnSmSv08+O1sbaEHdlHW6VViWKP1wez80
wkbdXTEzQzRE25wS17InhU+4+miBuCQTDqQHen8q+ZYjUg96Yl9v0n9arsRTPm+w
yL4bqJJkEY3alFx6eJ28uFyNmaRhqDNGXyFJ7GoBkygsF/1RojiKM1KhTW47UJfc
RWYVnq9ei4AgiiaEY0FXdrpUAxCMm6u5+B+q/th6JHh9tMlgKqwwz7439FgK0QHU
/VYsu6xSkPtKStWCeCN1X8a7cVmWy66yF8fMYzsDW8c7G4+3EFO2BBpGYkc9SVYz
Jie/FMkwdXI3eywP4jtNLjPd3tfByYWijVI2VUk7odVqp8Zsov/PdUhazB1HH+/F
hIctroXyeFEzBkGzvc5UsvazGGbsPOS3b4Ofbo5LUd2nlJNLXGGcPO7Wuvd7yjkQ
GOPmP0zD1Q7ki9oj/TjKUWwcJEFQOAqN8niEWi071ecsJckE5qrqkCBsIAkwK7ej
FtsiwZ8N63wg5O6CsxQkxUEgkuBZwQmeMkf22X9Rs6P2MmU5N9a/Dh7A4084G3kQ
LDanopJzj+vJfPNzzzRsXWwZqIuV5SFzp72tN6eCj58CsAdkZozYrE+2gNy9oiK1
lj1aeu+FifzQ3mhygrwIRZDT5FO+7ub9Bh45lnwTX8RypTryFFPeM26WzZijbOoe
CbAUkUxAo1wHycumuYKhSlLLX9UhiYl3VmUM6tr/fraTNIoJbhqsfjqYDGLaaDie
jU/lGutxJWymL12jh5KL5QrrBruUSzFyLT/q/cd2EZImAuXlHLMnyd0tXHl+ZCTj
inzJAE/Y4JZEcsZgtwhj6DyWJPd6VNxrpq2W5NeT2MltKaQTlJ4Sq6C2wheUREYz
TRrAltAW4ChLi5jaF9ZWKATBdG8it2j/WrM0HcB81vFznkxqDvd5WiBE9VBCjD4u
ppv0wWL8xCvq5N/gAaLAHVqbif+l2tLXx2EptRbnYQVDEXV+LyKynIb405WZpkXT
b3hhDLIZKgU/ZDEzm7MuFr0dd2rJjIDW4xXoP+Fu7dPzv00yqMVWHatgpnAMJCSs
zpe/o53YMD9VUlXZmGgBn/zAvVivXHQr3LngMcOgmOcLHneWL6GtSkt+zaBpnIqr
HZxrDG4ZsxVgvPz/oVjUvkvmRhmDjHvExwt6lDeG+fyLKYk7lrk0hJsXAEJyG9vm
yFoyWTVeK6O6tm1+CknbtTjbSQWk1n7tED88nY7MH2cvwIs8fdFGma6hJ0XSeNVl
4GIRRV4iNBHhvFhKKNZjDW7m1wh3cGrOSUpzDr5P9KIh00oyJexvo90ETnoNumwT
mF7VtRlZyE3V7NzD0FQo1uio9ctsGpiO98L2on44SN0V4gcwQtn8RwnSg2QEYXf+
QcPBr77uM8dSF/k8de/2anMQG74fXAPiUxN2S3HyJ3a6HRkKSdWt4qxWtfVBqwKm
uwIp92S9dzzpsnBpmG5zLowqDkknHxxtFwB1I0XL9u4a3JmDP/efhjqEACzTJOTX
eYixnxe0XuYmQB1GOChhz0fPPi/VoGiklCz+grKF9pH0y40Ueeeu2tM9wg3juG+Z
0w/P5EFM7BgNDuD4KOSuTT1YwPHM7hjhO+yYFtrBtSO3L8i/Yo0VEdh6JpT5dZHE
G9dPiFilx88sYVq1CJZMS3lzcWc6G73FnA0VJ1Az4f6nT8JF7i63yJRPsUfffhBa
ro0SLKFLGXq1r66TKETOhc7+lkWVJu1fHbYJzGRgO/YhbIxlUBdWZqsY5PaVXQ3S
oQzhQQzaLBu/7RCbTff6BUATmdQ21/VizBg+4/nW2GnOOK8QkT/X7zz6SmvPMaCG
HqBfXXw8HKjI072j8JifQBl9xSqDMhv1hjehs/1L5GMsFk5DeYhzZNgnm6upRIrW
s1cxnEH0eVJQTJ2VzvtjjnFLTLLosv3S9NR/3p3C5Tw5OIAC9dRtN5GGulH8FgxH
wrZlbpcmElZ9sdtQ1E0+KG3DOAWv5MiUQhBlMR5ijsbCXf1A5+Aw0NNQV8ntxi2T
NR8hr8vz7RHdODGOlRp4uD4VwKaUx6wxqyvLCItRLd06/nRpUK+w62zbkpHXYy1L
Gqxq9tql0DbMQEJLtUQIQDNcLnTtW+mZ2kqlsXttVDmudvpCghflqEYuqoiu+fkP
JU7QsEe1AXnWOH6RcFA9N07arR6b04pnpHPNHH+9uF+IxsqlozaLMUHrCOS9vgnY
g1f9wNX4yBZDnNbDOHX5HAHomYEmZgIoFq7SWI57hzKjJ3D6ZON8vraMARY5vePI
bU6rATw6F4cZ/HnqArGvXUKLb0X45fneDcP+TODV73CLCoQ/HEgBXiU/tJnzii/S
X4E3VgS2YgX5OE27936WNTdj478Zkowd9QNFNHiJINRmdgzqwxO+8TQnWyGYnqc1
jHjIbceHpp+K365dy0164OD7gr9QovKgiz5KCAl6xxoLatBCxyc7lbUrJ3zBtpE0
hT2eUSZDs8+uIAnuLQQqnNeAa9Zyjq62YttTLfkA06BGv8MGllvQkOg4+F/qIORB
cpB5LFXFCjnDZmg9rVri5YPqq46Aw7ZOwMboC9/WaemNRTBa4ZqSNqFEOesd+gg4
Wcei0Et9mX5Elj+YA0aPT9qY35kHvk+JBDiPW9/ocm9t76Imn3UIlAbpM+5wced5
uw+pM3SFjxFE9z7oZ0pgQUxndEFZ5R++I3hxpefb4htCKHbklqQIhQ6pZK+3jZMd
iLZRcLMol+mt1GjX/0anCHZ9X/tBNtwpKMyAZxOTVMF/quUY54R+vDJ73vsZsTSR
gAOees0NjMaPzASUcov7BX9WcDAOUhtRX5rRJihDf3/HsN/CNu/MMApdflBfRAMd
ktJKfo44d3n2DjvDAVq1C7GridrKux+rygtMUl2ZJEj+rlSXigiSK8aYZ9LKwaFK
PSqu3q+mZrt3L4cvJWeAGtL1CU2jdBQQxQkvoId3yx0syhZ347uMcV8Eqjzq6Aqu
QbHkveyBAqzF9+vjtVBQ13EhkdOmJdPjyBbNu44ZL7eI1yNmDyzTJPz5rvUVpmXf
waaZ3Y0iiN1VIGdMwiwjjatzotOfIYPQhuE2bFqt9Y90Sf174JhE4lyxvfZiwGAo
qpFiVIm8olkHrf9xG+HgZXwGiSP9BpqO61RMXPmjqrRyNDMnW5qYoJ1rEwal+uGS
wAV015dIf3Ttu4ZeTh/4tMEcTmAekoPFLQy7A6b7s7sl3eks2WLR0jecH87D9Vl6
Q9pi0A1LYP8RUO/2CGjGmKpi1uPwTEOvpMSAOyaJXr/5PKQjhaAD7m0P3PbmSJBI
iXKgV2dPRz8Tqofs2v95nx3Bje2Qc6O/3VVPr8QymAjbHku8Bbb4alPjUxKWXoi/
TvmVloHKqxhb5l6Bb7ce30fwyA+ic28PV2fp2XwIw7F8MMUf2Fcy/yAR4dRYsFn7
bD4MzQls/Hc0AJuEi5SYgQRmTnFbqhQQ9NZHcsRCJLICht/JamHulU08nLzYChO0
/+612jATYNxMY9W2pCduqfs8WY9/Prfcmx7VaBs7T5+KOK/fVfi7/uKaqSR8G90l
8a0FrIE4wYEzhh8+4ciOE9sVdH3JR8MXt/arIhgY35z/HVcm/tDsu48f/3zNxU2B
MGMhiOcMUKA2kEbcAV6Yc/U+xM+A5rHsaDvmGZ03AAFq+6eWhs4UutJqU+YvRebo
eSicM3n++25Vz/Ac+OCmn6PgXgvndI8N8kfPlVw6zqW08g0AdA5+POcPHDvtqck2
43h39nyBOF9oBtlewUBIBX9HMO70ZVdMYHfpJe9j5QVkfBzAmSSpcrS/5Ynz7Zn7
NvtDWbJ4fTkv9qV+/oajIT95TRo5BhC0M83Re52MfJY+gx4KQ4XRYfK/IYhxda0v
ADuqSxUvMkK7lCchtEHQcelMqQGYPul6BBNsP5oXDXjAYAfioFOGkheJC8uRMsGK
+Ql5YcARDDdLw7B1XWU+Q8WbYYwd+lXSrpwVkBUgjTLDuKwfEKfBCOyEpsSZULPY
R1n70li9dh27Xy/WfOVxCZbRUsabjKx7U/W3VqKzG1GZD+abF5yTdDy0y7EA2GPW
hJoCMx5e1Kow9WYAQJy/UBmfUaQeHp4r1JI2WbYX2H1aPGv0JOnHZONrfxlu86Yo
fjwgUq8Zetf2SB1P3bA6L+usAWOQhEW+CHvIozJag96ImNtixtfkgMzfk3G2SnRz
25Bhr+SKwOV3CRCS3WcTG9cgZCZJGKikfLC9YKeDG4015Nc3iwCygTs+Jv8K9oaD
jIoPBDfXNY/opjNidzAiLdBupS63GIFniikk/47oqPMPtoNyqWt1K1F3Kw0SdIzC
x5QlTE/Vu+/62j2zMZss9prajcaNW4V4RzFeOl1+1/eXOOu9Ap+gWBG4s71MSZyM
HvtTUY8ZNLZDFWJA7sBVn0dBmTnh21Nbh66G3X79KXTp9XrK92S1BrgyJ56Os0UY
YjVEBa+EIwi/9I4p3H/Jd1YpeyUAvlalv51KJRM4Vo4GY5oLwuKnyptT/K9BfujU
zgO2Ygq8eWoD21aHhjfCj/cIlqxJW+A8JzXBIv2WUwhWWw0wjvnjAdDI+wNn1clW
B+NYQOR5/2NPnV34OQPZ+iJvzQUT3SYKtg2rWjE5XofE1zSA3md0oi8mySixJujc
qZ/dkhqwFcgDt8ONgN2UUEwYGtR0YzV6q581MENBj9171cq5iiL4mTcYHNj6redj
5sCuc2W/8eJ5akZCK6J1S5Ui5mTqPAgMv79FVYgCH+BgWce3iLI74zSozTV+WE0k
/DOea6RtApOAIPIb6nyHnjxN5Sq8qXJioEPopjfZ9+uop4EDH1xpx7IO+eDk09CA
mRGj+ur0eT7Uu+A8qHlsd10Xy5cRW26FdpiQWNuPBHPDbE8CwaemhuRxJ8+wODIB
vAkYp01k4vbxcCGXtKsfFIkE5tacFxQgbb/Ti5HvLr3oYpDdToUj33xWusZkwc+y
YCWkNi3tS1FGG2YSpGq6egEbQZFsg2ae3JqW4dAUh2uCFx6XN63vQ4lRwe33vTqT
tuT+zwyYvaTiAVovEJYmSngZMfr+2jXCqhCiRYMUQxZhHHyMfugXBRqjq0YBYIGa
V4ISVvOE/wBRhBxaq5ah7CIH1nwiw/h8wjGFabtJMUrLqGZ03Isk0ED5dvjPocj1
fW4lDjYLWOG9p+BEY0RE5GzyZq9ZgWP2RNwAKtEl4QD+zloaX6KowtyA4WYi7aFm
ExAC6972xv6aw7ELt0PhdUF7WFG1HOggA6ELAp27w0ZcAGiVPnCbFmBqQ3g9As1o
ruqzoZq1mUORuKRo/GghUqzOD+gPp8NiMDMMWkNgf1dhqGwkf4W65eL2XX5/5RZX
dWzO6as1O2qkdXTwKF/WCzjJJ6qym3af/DS1ukelMOMhlW4rGlUefXVPqFjvcl38
Zpq+4JoY3APb/Sf/4zuAknO4Ju6dW7YSzeBe/F0Sd2Y5IbjchSd8A/mtyEPAC0rM
LB5LiqqduKrN4YUzvWQN/wSrYVj+b6cgGRO/bWJpmHrQK/PjwdYsTdpDtwhe4d6O
kCVY9iXU1C6NK7f6BcLBCh4XbQd71DLBEya7NNUy/BOoBB3NvZW6L8TaP290D1z7
G3Y6LQpYRwLOsp6SCngaOYV67g5l3fo2qyKupQSW/71AQryS3FW//75pirMcjFX+
OG+XsHP6eueeA/X+Sf6ivWPTbb41oMZiEnxyW6fffkQSwUfeqZ3F2YY+nCcbsIPZ
IN6K3a6eNPS24GVAu5V7KdwyWzwzOTj+HrFBwKrTyrdLYJAHnL8uwlCi9esQmRKJ
e5DXHEESvDD7n3vAIDWuoPPHH+0p+slHZpTIWliGI/6x9JwxdD3q0QoKRAiT9Vw7
RNkwmI/i/74idHwRyKZ7TcbyBLd58yZX/V1iUGaGCW+DNL8MNlcXNXFqKjlcalp4
5Q12FuVnQ3wg9xpC3Knatz15/uFOD4vEeOw0x7XcykoDFR3BWxIlfUIJxDKjyocf
WU832gDBbOOPQFVXgc9MWrsm1Y0Wsg35xvkehaBj/u6/etwE+KP/XfXkIISjL5vR
aILU4oo36QeuyQtdpoDrbsKt6D0MqxMwulptf9psQrtJZaFAgNI6CacZ5NKDgiOI
YQqO2tGKCb47VJVJh5/bUbtsvP7ZmR1h89HYa7NdvL1/f5Qyv8AVUpuNcZKb6dcJ
ugOBfY11PAFhKldcCD6OVl2i2LScElCFwAVn2HS0QH+VL4h9gOpQ5lssF2zfCNZ0
KUUYR9yzAV44r/QQG4HNE7mgrK5nDkoFvqK5cgHbpvyvK8oQoCpCwgNevTAuy2Qq
wppO1fuM66Qrb4zmQp0ytCv0rHmyR9pH6B/kPeIN01M9LUbpnAr5Y/z9HUWqoPfG
+FpB6Fa35lGe7/xLeGUZCtMsEOV52n1wwCsQ4tTlAceR/k1aPZbl7/ZvpuJALs5Y
X04+CdPHgDPqvUF5K5RQiE2Oq4vWmV64b6rYNB8bj2XmgJn7NQUI7sNFHsHed/9L
cKbiwjcoqvnWsKZVHD4myqaCVw9sCXWevMqc9Q4/pized5DTq5owiH0SrqADnRHR
NBO19RmumUZU4C+qW2uKdqOArWfLk8AGW60nsAEJYguXHWHCSZ99o/49XAx6UiTY
m6xcGAbgCFSxrLBGMAaHpKaaxWa71G/mcPj0o1irDygUiGQUxVCeeQL1QUmM9mE6
5cBWyHOFXOnA+sBxLyHgwDR4Z+omMg/tCxndbmIDSMNc6rMhbolUkCimmS5LEZyK
PjsCoB2JylDcXiQPpdjqCc9wfkVdBlfpnNxLdhEpNLfCcEp5avGzvD5SOJuxAINl
x2E1YRcwvrcAg+Rnh0dHojVTGBbkXj/L++xHPCJYFqQ5egSizSbt1r+Hp7Q64KfM
69A326+4fNLk2HGfLdiBfCgHHs0Wud4cW7UwuyrnCEeCYwHlndF+STLK1blN/d7F
fiDvyCpsUXB4YLSYbYEPp/hFgJiqEPkhPexQgqWlRMexWoLnboYHOYn6NCYamOxc
mNOXd3iMkY1OqSnkDxn9xcdAHoYwoOZKIMbkwqW6cyY0+HA/iW2+LINmRafbKOXe
QYyC/hkGQMObuaGOY9cr2X92QYuwuMeQ8EA/h8fd6QFe9u4onJ++eAq3UCHSVC6K
xJDAbU2ryRpq9AdU0JOkotSn5kdOtONCixuSDW+1cyjyu7Th0vTM1JBw/BSeLHPx
LCv5Wm7ZUTp0py79FAtMWDx/nBZgDrpGC5Ug3j3ZtilEpMJ/GsfV/oQrUTA/Ea79
hIls3MEMkkcprWNNZAiYVe6kNgQMlQuRvMj+QcfQLaEDfOaZKnJQsEx5X4DwKLeG
ZlH2qxj3zDqHKhhDa/qByO8uXmNeYl2rPKqhabc4X5QTqEOQdEzbPOuHmWelGf6Q
vBoxkCoGX8422SqCYsNOOeWn2LdvYYhQ+OlTZUgidSVegIuas37cbzskX6QtbykH
DudpUIp4SKI+nR9o3hEPfYbugGtcMuW4zeqNMd7LLdKAV5LF0G7afIFNpiw04vQy
kVkACI5W62ZxrKJTOQFc/z8yyZSxjrWpgCmnYe1ivqy+CKJEK66lqDY+z+Z5c1+Y
QuRqZGPZsuMjmKVKETivFHRGjf9ntvhgnt8wxunoPwlOXr7IzGTkTXm+Ep6MObzp
7pqrgk1xtM9Kc912tFRNFWm8XXSil8pn5s3gIGfgYchW72YFPCbWrsv/08DLwytK
A/a7ELqFDUOdoBdlNsM7QBTTxSlVnNFkdGpNxnNUpjt0am6duyTTianr/l4hTBIf
wyUxx6Kozv3RF/TttxKxWEdVuhIS7I7bYnOLHzifokIPPfZiPJuNoSOaTH1xwFw9
3fxQ1yK38HF6z5qHTVq8aw4FyudFD0JtWPZda2EWv1ATM2xJ5A0RUw0DRXSTJfdK
l00LhgHC6Wb07zoGJNX7xPbeaOLRRyvfJej71wN6i9pIshj3PYRUuWzOmCGQFFoq
/7k8j1LsFRlMdTMw+oEDqfINlnKScBSJXHp+XUK8US0CrcYYtE3IDXieQRBy7jsZ
yuQ1d8KfFPoGtEAnlZykpKNPDdI5eOoBKP+b4pdjiSxV8CT9Jycm4wwgz/vZasFp
gNKs3jsv+8Iafx2LsPRy2kdqtnapt2LsWBWLkxQGR1BJF1YnSFQiFj14Kzxel+rD
ZE1ja2Op/CrgjjGXP3xQEC0XvdjI/q9IstaULhqfr57ETE2m0KzLaAppjliOKCw4
tcvj893GV541u4mtGEXuX40wzahXfKC5fq1vrWYFGOHcrt8Nd0y7wywHpKs+8hgG
z+IFnYZDNamjMNYluyvQgVXXgZSnu34eBSbLlkqmzCuFVck7mXVgVQO0I54rlWh7
C6rgklDJtI1YADIUMEsCNg32rBU7AAaRH5ThaaVOS3Wo0QjRi/iXEjvP7nYtT9Lf
yT6bltpQ55QKwAi8azi25OKpLqHt3WJeRYagtwQI3JeKRXm/rEU3YmPyoaVQrgqk
i+D8UUs3ipsEydf14SMbo4d+OhCSkd1i9PmAelnrI/NHg+BckbGY+S6TP45Qzs17
Oe6xzRh2UwLrlgFt2YaNV/cSIPjzsiIPMYYxFmWxK4rGMwgRYv2P2o+PUYA0Ad4H
LXbxibW+ZZ0JuWOJdU3PKywfv/c99M2VP+sK84s0FOz/9ux0ZYXvDGwNfHvh9LiP
BHdR+5xYDVkI7p1XJFhHG48dVJBFlNh9q4KwW9Rm2pC/NfAqgVooD0Vc9SabF4p3
dh658IsxgQm03JXj3x+TuB3J5KpAWgzsMPGubQ8s2uvsz5mkLYnP7Sl00hcf5Vyr
2/1jOcZMmj73wG8IfQa6dNIlYL5k1/w8R3r+/4l1gJrTDkc+h4Lq6lO4lWm7WuJl
f5f0FdC4t4J5NbenKGw4w1fTF2xDX1EZNZ8sLEYV7Mqww6KxKNFBXsTsm/+NKAfK
LgjTlQNd4M0RnhZW6cvJbHemT1s/JjN7zESO/+twroTIvPcrcxHnfMCfN7eT+Fnj
X4yiCFQjP0zdCatGO1asvWpB46E0w7dPybjOL3lkjg69p88D8ZDZ6KmUWny/5qz7
o4pMCDH+aoYW/IfcYuDEPodmuc0r5g8FO0Rplom14SYUB/9J8Y9OcU15i9q9sdsW
RT74wi5L5ZuqsJiXZCjbnn8mmw84asTsCk0cJc0K4dxJZxEkmt78vk3yzUbgcGQy
t+UkMqSIiBYPzabFKxngLw5pZfPC1v/5Lqi8p2NnJKFxImlTeRQkgj6EhzTmoQFn
HC09TsYIOtYXZX11zX6aSlffHMDUrujJ31nXjpUylC3f5LzwKeq+snCEmcYMAhMd
aKUzE18W3m/LcTlf4U9N7OFyGAlyzTcgXdcCDkkYGCEXyjqr+K82Cwn5t/hJqMii
z6rJd+NaKv6z8iz7EYfWNIgMHcYkT7vj8/D4ucJh+th/FkF5OxL4iMjlCHkorlM1
ocAgMq1mInlhnzzvE2Y/wYnO3rpzdhiEOnKPK9ZwK7/uxdbwe21fGjie60F/AJ9F
7/r7haHQMgGGgQ5AgB1J2tWv44pOAyRqoRCaWcywAlm64r52J44nTpxoI0l6yV3n
YwB7aCYpPhP4WKZmyl0Egv7Ovh96tpoWcGu93ZehC/41zQ8QJ4GrkjonP5e2e6Sm
qFT/Thu2vh/qu8U8EXVIonFrwmgxOlW7kLexsifFad7o6uDMnQ0dz1c6LKfxRx6b
0or4SbiV0WTHy1Xb5dLAqZM/oqBGlfQLlCcrSGowvTEI8aBffMJzvpqlwnTDpz9N
mheE4dfPl34J6qbrLn3908/E99ZNgWqmDj/SnIp82dDe6P/U/WaP8WHk8BhB07QV
p8tCBy7Xw/aDwHsUbjeG/ukZLJusDkUPQY63sRdD60E8d4g1cagNO7tJqdmZKi+P
MTZyMqz/KiyAynu9Kefjyf9Xmk9ckxCRk82FH4OAyTY6f8qGM3mNCDt+vqBl6BUV
j/TUb78/2ULSlzWULwvlol0UFBYFVDG8Hlhp/rX62dDWZOZb3cXSJ8Q3IqtyHtlK
jc1XF4zWvbs5cRHG9Zyu78+SqtiiySNOaQGLFIBF3sE5U1k+jfuW+Mrg1HsAeiHj
EdOuCksb1BpJ1nnJmEJVuUn32xn0OjSUYIgTkpmzO29VkPFa7LhYWj2kEUifwBV3
9W6GtQDruFL0vmhM5IwaKkzfmt0FdFs4eVjjb5T7RCubx92fk+3nxT2IXzmkep4P
nJcUcBG5OL3A/SumdG1aDve3XUJWUEGh1UMWJl60eYOPULj6gIsx2i2zdbySeb4I
tzC/E5gv8Ln945HeD/ygeM5OB3Pz7pjqy3iiUFYWtYcBprXgLXrWWe9UqMbWCAVN
oUoAeTlaWkkof0pYLS92YKrAYZ/SgVlNOgafOj0GsttscJ9JSmtW4g3s4J+Plr42
qc+r3P4ucNh9a+STOL2qeYfrd75RfN/IVLqYioRGq8I7huyjFAEWNQn2ZDUVCytQ
PiZ0dZBpAo9ORcvUc3pw/JoWcnCTKs+pR81HGBDugsSLWAjo+fbPCPL7ePWKzc2Z
Kk1hCum0ro3bQhN8SMfFiOJGv1Er1LJGYXg6qi4CtwmvHxxh3oXo0O5yladRo4fO
x0VF8bZxgnvRdFeec+Ro2DZF6JvLJ05KEgHM6nLKd1bgmLvodB4IKBUrKnR1MF/a
VaLxI+MYCKbMjdpbZTBcdJWm1uLCgJmeYT+hcjQphTI6kfqhxWfPhXUkozKAcAoq
Nkg0Y/mNwipqiJJUFqETeZEG7sc+8JC+XrlXuwIqgrxqNS1L0As418iKFlsxgYYe
slCuSzTAF/UZRFOVl5TVctg2/b1w8onJKbJ9e0g3bzH+YHsAD0ywdVm7qJoo/FdX
BWLqBTUbVzaVsRtlHy++3J/o0xzxDQlDeB9685DXi1uP9eRxMtoTYm3LLRKH3hRf
nS+385oqVDozaTIc7BUP6OG2hs7dKqLmJ2EZJcqou6hgyqHzG6krDMaVNW43mbqu
LtrVXwnQn4CWc48DPW4U6PnwKwNPw8ITUxWwhs9WR5VtMjzS+aZWPxrBM33lOHSU
wj6pC4Vy/pCf4JjwvxIctlxmPMflH78BamVY9WGURb3atf6F5P2jGoODj2SgFxXJ
s6qW7yyRbfNqfZipfU1ARGmXjmiIbF2Dxm7cOjQRm53SeYil/iyQVYvdKcpRbZWJ
pgMkY9UqXXJqWrRl6RYCFtd+uvBjiKsTFPsKIQIM5acf6UJgllK/chL4QaQFoFtm
YjMgAUT0B8JS4VPYEaiNnVRULOO7DQEkqR8Nnj5Dx0omBk9s4DqWm+h+RNjcx1bl
hIGrwcHDCBWbT768NWRL9HpNDPEdxqp0+W+6pBMOQLfrLhEcp3ANezBT114IckZ0
xhQqKVPOVVXXXcR0e91NOU7CKnY7J1hJrg0xFeXmiVwg7tM5B5XI2ohGPHGiqGM7
7VXqGr36Q4z1ZmRJeeIWja1VfLtMyANrmgL8MHhLbh8/wc3K9AlaXSCNI8P/o9dj
5RxFTFm/u87/xP9uDKtw4nNhMSX23mSh6yDh7b7NIUe+00HvnIFqOOYf5TILCSJI
l4joFnFON96wPngrI74lXNSuInemZFe9YyPip6uwMTq4Y+SiLLr0jkbyM3BGnOCu
o32KBlZVJtUryL55BOHPBsclEY23ovM2wmP5TUixGoykMCgfEbHiaVP5Yj67FSnf
HCUf9796BUYxT1QR5lYYTPQ5jADMvALoOYBdOXNK2bG1uhfSYhDKdH352Xr2pgEA
yfvTy3Vkx/d/d854kZJ6u/QK7PuC2K5gOM/ghP8py8U2GYzq0CLDayQa8k3Q1ygH
58PJi4hPwkcvcFtuVq1uwwu7z6HCkmnNhfSrgAInyMIsgKo/eKPqofKE+jyk4FTx
6v8g9aeiGvNq1rHe2kDNZc2wEck7g/F+Btwo8Yav65DD12uWpqp7RXKTcmEUgG/G
YxNUs2Wtya4RF6emIOh4JLiQfKN+DgqZxhLckMvtCfkTfbFwxDZqtwCM6uMmk6+0
rYXi7jChK4hnYOihjRfSs5JIxaLtTtTru1FOpDOT4ewRqvIhgxEORvCI6Q1aKT41
VMpjacFpPRXwtLaouqV0JJZTdmdUC+/vHdccvuQj4m4Ob6158y7/4h0qEiFQmBOW
QkFXAKdH9SjL0RPgqQQDkgH8U5Yw5jZrKT4jlvovatAH41SIvw98vsNT21A/RvfS
FXU6T30DjURmhzQyqNo/RY4WguOjnVG41FQ1L1ZWO4/wmbLq9QqawAka4c2pGX4s
wgD22/Cr/PaDvWQ7RV7Mx3O+DhGRMHuP0D48alsNQ6T/qHcBLy4AmvQIDAl1fC+r
D9vlTSE89WZ0TFzRWDNCagt1y9NjhWjFUtVWJZLlDvUzkk3SczQdJGiWtOk+Z+V0
ifjnqekq1zBkhomIFhrbSJkJwWtW3Df3DK4nGO9ojq3VIiaLbCGe9QhplURo48nu
RZl+sQhtq5bOE3YrLjyHZ/Pp9aqhNTogCQyFsKPgGJaWMeSqOj4s3KRokYO7KSVo
JTAisx9G7A4mCDTDDWqb8XbCOfRsXc/beYwa3JRp0NSagW0H0PMZymYdgD5xorDZ
D67aoXgqqhXk8FDPhcvmLQ6cXZzU3UJcn102pgqpUgNTf9VcJ03OfYQfFvxkVdwa
sb9k+rhAjIGZup4CdoQRaz61oYzVk7Lo8L5oJ2Id9pswdVxDEvi9NLKNNQTGd/se
HbvIUuC+eLM+tE3mzvuHarU7vR7vPgoPsPDY6X8u67IQMh4HPvR0jpbrIgdXg6h+
doTkCNlKQJpNk5A7bigaZKQ7p54w11Xep0kLyivBXjVUyUodEG5bWfgb6N0ZJLZ5
Pt0DZvXFK6Q8k3atYOfcXzpz/fO47Xe+eToNVqwk8MhEWgcnOu9zPiWspJwQYdXn
lybsH9fmE/yQH1Ds2+GHObTofP9khx3CWWklFLV6brPtmU6C3YoXr1HdvC/BtQix
Lc8vN1Ok5/4ZSptruCeNZToGyS8oUcQrh4ISA00ou3/BmzdT9lHQYi4mFnaLK+qG
X7xw/GlLz2hWdzrx54LqrGiM/XV/K7ZaCXFXnggyzi3thkPRUe3FsacV5XUSbhUk
lCcYqctyrG5IBEmuNpP5zHTt4shsdy2IXiodHtvWkwNNdu+MJopHOhXpnIH+/nzh
HWnbNIQhTeyqMXdBDNJn16nV1gjixd/GY6sjigy7D0AVoE7//m1OJAWQJ1UNOsLG
cc3a9KzFrvWhSLrWGfXaiN7w6VS5MO+8v2+eyq7T1MkXypMM86fn2+7tO6CiUujy
g8NevQ5b82W3kg2pMP9+UA7OlJHQQKE32oA8eowihhrWiWVLKx3xOxJOOpeFEs7v
USQx0AiEtnOiMB2tbfUgRJt0FSbAhi0Fsccvfwi27UMVVC6nz3Vpas0gDHtMDY/K
J8memarVj97JraXmOJOCmCbiyLkC9PdcMJB8lj00WcGwld2T8iDcNBai85HZMclk
M8hp+WvUkN/nyyYA2b/EL0DHz1BsDpgbGj9d0UcUK4czAlj31QJYm1AnLBoc3m4a
zavkXMxhAsv8+9Y/QuvuIwqYZWsxIQcJLCi/fkK6O44ORc07dBC463m0dtEORKRj
mxOfXXB9XecXzW6ayxWgtDkuTd1ukZNq8jkNKk+8kWaRVxOonLSqseg9R6bsqAvV
1gR5Hao8CiY65OOwlDauSZUBVht+BWwE7hNKoDHvU2drieDOP6YMDJz4tV8+7m48
11QQTwJDxzH5eRh078JmW97C/B3pzTBNkPaZ1Vgo2Y9nfYKbAmSwgsg9QB+2Z3Qh
R2st0SsrJ+T8fBx2mm/OKeBlt9MsAtOMoad3psgLjwyzMXRIDInSgqUOdUQIa6lR
b3kUvWiW/Ni8fqkdxwHBN/agR3YyvKe24+xcOHAq4VIjsqZ3sU1W794YArZV7Ws+
Hytp0q0TYVPGd6X4h/lbpRUg6Ak8IjVpBWdHtkbUdYnDELWHjhWHDZcDU64gzswD
2tBOOtG6uYcuRqOMuXQWSc3j6MsWXW5B6wbgmWai3Ur/vzId5pe5WWeoBNdXX1q6
MNgS33NkyIFoMsjcF8lw2njGC1Rc+Yjym2z3VRBo2RIRBmaiYNxCU5T4wSl6kimC
clRGucLfSQv93porAjNV5SytibboHmrfuuILbzPazrzfT13RYfINW3uKrnHkBGHT
iCFXVXa9OLoFTibHyYGPHGIBU5U8kG3ElPsQPYG9wjyKCk1Yfyvof/zca/yCQ4zY
Sg2phfrz5YtgWx7+NONgyl5E4NKfST9iLCBTHKNIZKCXDRZMZxPUnRtpw3f1dtBX
cPRisbMetm9Fx8KR9HNmPARw8aR5hPXC0Qj+I16wFT95AAq95xEdnqNnluht7hi+
WRIEoJNvlMB35yUQeOmmaeSMcL8t2331zOd7rhI1or5lAXJFGfbxtZeR36Wyn0xA
jeS0x9pHee/iq/J34BA5FfBts8RKnrzu5s05Nidz7GOrMXTor2kCCdB+TZUlRMar
ehubzD3t1Mja2iatLE6w2CFHgnNYbgOKCEQ0oQ/bBTklHs8BtmQvfNQ+J1u5zYaM
yN9zYy38knoV6KIy0GCZCDV1Hm2JnaVB0FyicF7IzbnJYKR5hkMME4XYj+kKKrV6
MBlnUdOBuUJ1KLCPLEmJOdfIue3ggrK1wjnY/ftq6DqQNCHtsHfVBU4kbCCoTr1H
g3ss/mqyaUvCuclfVb1FUdw01PK3Z7XgRkcr7KFf4OCpm7bUR6TuC4YsAJphwYYK
M8sxVrxWoz0nrAeuFf46LYabtuCxNL3n1YDvpLqphRyy3WhXsNIqgR294NzvpZxy
NNzNEWXMgyVU2VsLr1xWFvUF+fweq7QMdzjfmL+9wxqwF3x3PX0gJ+dJ5Nwa1EmP
JaVtHjE45EVkRTKRfg0htevSq7+Ijs8YFPJCqkBJlOA10PT+rDSM11NeCfAAkBnP
ys+L5pSyDljLR77hJwF/r0ixR+ZF+w+q0TmY7e6ilaPkIR3fRlVNAiG6pYIvKmi1
SHo2hlm0K3FYqA1r2/9WlgM1cBFhFEbX5/YwsquxypOol2aTPp6DI9+E7UYOPsM0
ZixMnJBJzbPEyQ0zW+obTZJvvYo7u11jmH28s0QLfA8dSv8pU/siFe+0v4fGiCpY
ifK9AyQgtKVioBlav5aDEpmJ8xiYvKGYfQeV3W/SmgYE53ftEfuS6DYMhu8pijqd
FkQEpJDnuIeFd35zwKETddHMzXyWCTA5ZPvyByEvPA8zlcv4X7IMFPl0NkrqMtUd
HPU0W3qk4lL2NuLnpL+4efD4kNu4VE18motXotvoiCjW9PoYqHz+59XzHW6iVgGb
wnmIsYzP5lqz8QLn3mqTjVUHxc3NFIuMUj1RBXG2WmFVk3Z81hnqv3wa6ooO9m7Q
9kVywXu3f7u81wUj9PvTFDpUoB2GwjWh2w9YVe5tIJozSp0RprkEadv1Qv5RDpRh
jwsbquqz1E3mp/kEflvLYyzilwwN4ln7A7uB37GfyidU3T38Uvyjx7e6gMuEpCy0
uI08dfmghpWrsQ8RgB6GoQMwBIL/BlgeJ46Ju89b+UfiY6KYRSYsP6LtozgUbwBN
h9yF9l1bkwv2qge0IqKT7eOfma7DCQQoNcToslrxK8Y2XTruWARmT+7vt1UPjgM8
MtB6TkfMMxlGWVLP/aVefrC0OTK4BmQ3/j+3IL4GDVQi/Wp/HWq1W692ZnWa2wUc
Fd9fb8dlHt3TgPpx9TkwHhobESrMowVbNVFFr8jX58FeLlVFh/ImLwTcNUAEc0xf
wJi+Ef6fWbS4uU6cD9UGs0AxtjeiAiI+X0QqE4qVpUUJiRHRP4wNRs1ZwCDucgOv
wdNMqKzy1GVC6tbz33FGNU0W11DiReDRKzx+Fc9AtQicKDwEf8TEWNUbdPj52RfG
rwBc/Nc77fV2iTx68AuK/80SrBPCMCDgBy+02M5iWlW+B0LjhFYcPuQiLvOIAJZC
DYmDpCLgU3NcUMk8Korsuca95fbo2Gx38JLLbORipMWTgLP+e+CVTHgsdnMX7hDJ
P4C2ZLppKlXP7jOL+fnrP9hfwL2dVRIABFhCNstIgA79uvlJ9Y92uZGFG0WrOjWf
WP8kOIJZdGbJ02/oGvL9dnk7FwVxJvDYbW7yhjXANUlqmCt7dtKRl61iQ5t+4QzX
bc11Fgz+xZ6VDZVzG4NhdAUp9vSETEJ3GVOWW8XThkkgDsZtzLn/bQcA1qVourG8
RVuMAox0eb60B1/fKdJsM6Y/YmtoUjRjYsrF4qGIrZfUJI1XMqcf4jOYddP9vpDk
mouECp9x2qQf4PEOw5zOXr0o8HkEBvXBs8MDMy/x5WRETZnZBjSmmEx5s6UE/wBN
ATYoY3BR8MwmQT7fE6P+GmVqtfFoE695jB/3sGT4abr3kRk+lo/ynXh6STEdcVoU
6g98ByRE6WkBdCj/8FRPS6yBR+5KNWRwzyJEo3PcDFaFM+2SvMzdoau+BItmfJuZ
fszrlYDfWAvYBw+N1avYb7FFJdf6N7mk1/iNoUhT5EyxqasLCCKNtueqeVl5zoNV
vemSx2DGU7oyJl0lo719SuQub99pEyZi9N3HLbSpKVL7BHUOM76ykokieVqdS4VR
5/hFqSUctYBBOVZeAfJmPJlfbE4QDJ6uOjHwg2+qJV1C/IER4eDj4m038oLiK9TK
ACXNVIAZbIsIzyYNmqCWiNxAjlive9CDH4WQtIQ1d47w3geRG1ZbhrJ8+aH/rW8L
DKJ38JWwI/GgqmxFRrNBGd3PKvv4HiFgrABXyX0NWv7hIQqZsSRedz3FkAqEvXX8
TfpVOvKy3ffha08ljPOBM3acFcNlFTOstWt6NnWXmJ2A4qLaSSeD4VfiDEYHFVss
e6Fc/fS/Atjd3mXnfDPrY+r8V/FZtiNldrXpSq81GG3uwJs6Ea3bwn2oy5cpTyOk
aiWlaRis7SGpDs6cAUJihfLvWbuqKh6mCDydBwfO31JpuevnJfIK46WpdWEm4iBW
CyMpTEzVH+b/es3M1oImOEnM7CmF2E6NbxkibAGo8g5fV+5FCQDsfmHi6mpTtE/A
jyPL+jsLnpNCF8O+XU9rScpodznfd9Sil0T4vmsnVh/aOthHa0R4cFAB+BHs/sTT
lEn+wdevmY2OZiw7x3PNdZdQ6Q0tlMRg0TjLdYPVWiMwGAhiqwbKvLNWhqKvKg97
/SmicydnUMnmjQh6FRtXvgoSqiODd1dwZKaE1T8FwMlzZdnoxRMgSGzTNockXVdZ
raBWh2w4S4xP+I/CzLyItVf9SszWvj8xwMoJpL6P4kvMgOYCb8cYiS3TBrdTRJVg
KJfnwvlPIIC0zuQ/URQTsGmNBB1/W//bwk4W6xVbq6SgoE8wmcqc8QJljHsKSJxi
H53tiFaKA3khLOkk1Sa7EHatX/hapkcSflyeh56x+AFhYC7Yft8wFuxFmrfHF0Xb
zcLkOhFqHgXvikaE7bqd2iw7MlsRUNP8LD9AmE5Iyglq2+NBCcHVS8ev/HkhBzRQ
GpWwvOk4Ets28DP86C46quBe2pIDRkmWkFH1xKADUomHHGfx3Fdz1Z9dhAr+yM5f
gMvDADE3jT+yia10W3sxKT/hRXgRkaFxyan8O4Lcs2GqBZMUnaHK1cMpytUXIv69
VQSYWFGk7dFFIHnPQRh2ZLh4qb+QicEkcVK5bOaHLCuncPP8Z6mlMbHAuVU0PPDk
WA2YHYelwKe7ykvTcjxbq+DgQ0VCdXHMOgT0JPmLHdha/Eyfhya2yJ8ZgqywjM7m
N1cGp6Bu8NHvLreKDcYdB8XXnyL1iZWB2Lb84+Qpvc9VM35H+O6VktcMbpJ6wXbl
8CySOwQxJLgH9uP4AuV7FMJiWLL5L67BukBOH+siqtiig8Vrz8j+JwsqWNWvZk9K
ZsOGN0plUABpBvMFZUW1cQ1ffU29Cjn0vx7kxcKFJ8+EDNWWJVLrNOn+l/lHWXWB
35F3LFX1qKAugNoB2dAFHixrpXnqkJvrg4IkfIZNrMkJ+muGD6BfYK9coJIx8Qr8
qRJ5h//f5f0+e6u1pPk2GRWempSxpY88Y9Y69g5jGMddDqmpe67s7ZuPE09RqByA
zmNWyStFLsqTvvc8W7YqNgRWc4EcXxyf8HgdvdgxmEjSLKP5C3x0GntWiwfK/ysc
pMDcFJ3Pp0JqZ1deiMSTxgqzt1ylX2w2P7ZTseRShcYaHSxIkFmCf/3i0dSwtuXH
nE9C+bdCUZnKJfJaY4df5x7JJNORzMFOXi/74onjaqHL/pUY4niH2se1L9q+Rrg4
W6/tQFCpPzt2wAY846coINNepGEmXNvn00+jhjhnVM0UC1lv5KGqeuJob6roz8WI
fHpZf2pzaziO/k/+fTG5CE2IlR5BVzhjWDfg9GKaFrgbd7HWxlWqHKgAGTLJmoM1
OgJ3ZPUFoaFHE47rZC5ZxLy3uTGZv3YbfVMy/Vss+JyRTccmEODRWWBPzn3pG5io
FumV2jhBpsMSbh7LbGirUPUgPcy9jJG6JitCdrz4AVG7EXkQFoAySFi9etvSVEzn
kh/O/lifli4n2Fp2JDJ6cQlgrdmvQTkgmrT6mmMkEhNg/5SBqFkFRqMPnKH+eh3U
5203I5+59akBLhKoGa1J31nygNiYahvE9Qs22pz6a1ckz1RlPOn4HUsCv1bCZb+7
Fg9fqEmWpQFDnjossA9diEJM28o0eGaN88QzI8QFlw3/5RaiSxdP93UGVCLkY3/L
/bpXyEhWoUFYojZWVXu+yTseN84bST6i1Y/dH+GOaG/72eNaBkVVK3GLxfG7wgOc
KUFy9N/s9COaXYZDwiqEpz68TAdnxWq2mSJf+qc3YApIBH2RvohZ/AzoMGZw7Uyb
x/4XI0W6NGWm6DB7IqT/DcmkIJKnrea24M6uoVocQeXaXMmPgpyFSBGPXTZo6/43
zelQr4f7oKVu4uFWGCMz9w9sNKYlA2CU8Ht9Os0mQfufhelKHEkP0abTjy3dgCKV
jFaYL7j/RgtALxGdbcNSXyRP5etszo1FwXi29sWuRg26n8AmMM2g6WpePzOv93r0
LUXRIi/DGCuO0cgvSG/2EueM4jKXk5QIVXNchaSJI5IaMgYv7df9upnt4aFV10K7
dc21VwSwPUPRJxXNJ3A0kJxLuM6Gwm58d3tSkbisLnYZ8KZirOX80AJ7xx4NSuEF
NMpS5vTxotZt2sLKgrQD3YicsRdsf+ilnNlkTAls+oUkYNd0vH8dmhFMAsNWEzWY
zM/8YgRGWDFyVqw93i1nyvlST0GCKVmRurjeneRQsrK5fBK0v/8/AoydOf0mWsY4
wOyDjTP7Eoe73K/XoA9b7xdH+6O25AdaN+GSTMFvneTccoIVBafe3U2FZu3A8m8l
G8YXb+/O9Ccide45WBmWHbKwE8MXyD0zLapNPX4/lhk0IMJZIGkmvx/h5uNUWIJQ
8/x6vBSk0XQ699pZtO6uVoW1mNNuwj0FizQH8BDvckHqSJTeoXuLq8KJrptnFYwO
UmDQY3/Au9xazEJ7rasnDj6fhhwg2C5Rm+OF7/JwdAdS+vZ4b0hi0sKLQW635Ic5
vU9ggm+yxrcuoXolrsj5Vp9ZCEDEdv/BqL8MDBTtVDFavlubS0L9oL1HVf1h7hlV
CSQeuJZ2cFJv0BLe8MryfzKiSenoqSXNuP9zS1zfiaQD8CKm+PJoAQTYrZ9SYF0+
mZ/GB0VDC9cbDYSysKlK8DzgVxLl1DC1eP/+0IfA8GEg51vgmeQoRR0hPrv7bFyS
xNte1nbnW/ItgOwR+47Qc3ezIeu2UazO45VGTioSLBZcN/eJnIT2YrwcRIva22H1
1ZtStZTtoJ19R2NMvVC3/ySP+pDUi17lnhBm4QeYcx3RbuDrMJuqBlXCiBb5Z8Tk
K2UdHNlJIrICUtXJZZBjwHK7Nsk7/qhDa4lywNzCoGgWiAbajLFxli0f05bw7s0g
HsDzembDrCI1oMp9Lll1I3p0OYT4cgE26ee5x07nnK6XjQIort8+JCIvZKEkT2J6
bosQwgl/7F/fqmXqXqtQUextEevUeFTm4HBQjwtWN0xBUidYsj+hYxaLfRMODivb
Ztg3pe5dBdxyD7AyHCadvEi7Bh1VQ6/JS0n7WkeAfnhu4o6geLF4981k/ULOoyEU
hkpe3G/cXk/fmi43X+i4ambHADWqwcFLPMhkZoLeJAenJbE8qG3BP7SBVDQqeKLp
jqGIgH4xAkUPYGFIM1XEakU5Xx0CbGPPKO/UDr93SEqvINXbixSQ3pSFF6F6fXeE
vwebZaYqIos0vhgw5mltOJY7TNPSMQZhek9SGChFFLpqkq1jL5UrzBflPlLYSepC
GFmz+27iA/2x2s8tpzcEdzpgjDIls9YAsfy/tlom2tEDGnsxbghTvdrz7eVXkGAR
prZcG/Yb06nXLpERvxe4LEdJjU697k1tkABGRuIVtiadXzgNKcd5yEran+3Hk3qw
rmSTuqPW/GDIYAkw3h2LIrQf7dL9glWZ8S2wga2inJjzaNWxH+xfpgYGchbaZxk4
Mf8Va0uffHURYa8VrQncrz/mGT5BjVdYwZa7CxXYJhUPkQI7q8QkeWru8jcRgLMt
cPAdmrTz7klJO3hvttUMRaw3YcLcFDxItYe7kFxwSwDPcgU0W+C0F9zrWSGArfcM
QWfufD25yOCi3tmoBx3JJu0j71fG/t9jJv0j912JCyGFJ9rqyNUNBf86av5zeDUW
e2ORhlAE+aX5g7fJCe2k+FVc2dcKlP+ULvTHb/8miveDSngMfs9e03AMtnbcXWDA
Nu1o4NC/HIfEfqLcMN7HHF4EPJe37pGGVr4yAfu7QIG9Ha0ydnkz+mp9/kIRLrl6
IYj2JqbQKb/YeA4TGxHF8TLJCucfOc8xOB7uONFIfUyft25suVl3XyS9jGgU2C5u
OZl6rEuLDeIexdG5Z4sZCJa1V8ZdIvnoS9pURYEuQyO3lhbw3NMjaDkYthweo6I8
XncW0n3gYjnkJTV6O3mt52+9R2z8tqmxgsUyLt2SaKrr+7TUutyL3tFzZKcPYfT4
bzVyYxbzr0hn6VscD5T6zhqMfQFPoarLnI906IZpOUx3UFtXexWSoFU0UOFmCtTf
6p8F/OgYMrwZZuLY9/nYsGmBGJyWxlmwsnkd7rqxT5ErZo72xBj9+NILebLrMNOz
W+IGdbOLDwoph1L3aD2rVQDUuPiA7z7Bj4AIjuAr7Pe/iGAXR/PwX9eWrNQwnil0
cNzM2SLUbwo+jgAPTBTiJfkcsLpnIrzRb5zf2YEsJegNplBhEEyytkAJztAPrZB9
zrbIR9FWiwUpzCRMgLOuCMDaXZP8XcyVkknNFvsIuWARJal4KTkIRw/AXExOrtbu
cXh/fA7xvkXAj7/Bs0eUc9rPB21xUOU+P0k4ecJS97Zg/f7/u+Ku9CsrTFfGU9p/
c+0sCjc7qxacKjBQWSzFqCGkOzjoALh7isAB/eJSvy9fBg3ZHEYlenWB9aLvpY0m
stFTeLWIu7ZBuZOH9cut+jGPI5PcI+Jj63oTkMgOZwfZa5v6vJuugInHVMCfVghr
EMBhjCvc/9AGojb/umAusW/Eg0fhl8x9I8DqEllZCjvtMXsDhSvAZovEa459IaG+
XaSC9kr47f0wjBOaZg99ooaCMhWGhxlZrB/53RQKBR77AmP5wC/nTMuNLZ9nyq0k
VAqCPMH2xL9jjN+b774XVm4UZUyaxp8pAsebQDsizSIy8htQnwRXNlaoG1LmCp5h
y9ROEreoF5nytAiOAx4blNDHdyOgJEIYBs5JJE8bJKlQD+9VfsHirnJ1zWcl2c3D
VISEw4GN1jkIg6mfy4SjREKKKowcrVpRW1bQprpYNboNj5c/jDvE9cXJqSvnUjj7
EcLPbg86Li0mrzWLfjy+FhPOeDe/P0tG1CWCpAdUOhCtl4WAmI0iNmDVDcA+ejzc
n4b7AyaSweHwJvcI09LzioBAa8VTAod7sT+tCprvVX1wjMZ8CFzYIGUw+8qBbI9g
S+ncduUUhZ6EEnykQC9ATZ5ja+OhSlMMU/XoZ2eCD6lrBAI6m7ahsVo7O7SDXKue
Nfc0vagRoHyF5uHpMceXedBrkAfSVPcNbySHdKfKdin7EVh4zwgl3UKBW9rUHHvL
qgbH6wK4u2orqQiwpcwIip1s+TQmcu1mqBw/mQNxiSWy+IVSyp5zDX3Jo1/dDckC
e7/lgYi73PFLR33EjQWqhm8DgapOzg11TVS0IwUo3H4IIX9+aC4ATLByubzM5ffq
Sl3WRh+53LA6afKHycgcDIvTmmWyYKyhnzrGzMS2RaafWRbuXerB5BCXlK2zwVuv
HH0wLpcO7q/du7gR6IEl4OgCRy44t/ux4a/Z+VqZALYg/w4ZruGOGDS1uBXFwMaW
g3KNrHnnXM6UEmG6pMRUsQdZpiVBOMPo5ZYfGg07vYIbBGlr3ZBvDNvHNnMStRiG
6qzpxQ8J+H4WcMT32gSzbo4rQd0ph80sIVz1hcEcXLnIRXiE0LViwJcq9a7ohYgq
9UAbV8kJ4Z5egUzkaZSFAU+3K+YT4bM9qrmrDSNHT65H6+ZyikMbCs69zrQIoouJ
GlYCmGQCwghGz+2EsDnkcmhk00VS5SiDgcNK82X0RoJnc8umd+fXmQU4V1bJ4RYM
wtmtT4gTTb74ulRmUCZYobMMk9/rc1/mBs5oH5foRx/8NMhgbYVKpRmqlMevUiuB
M1gAgBDFIGngmprpYmTcWVI86K2LmJXdbJEvSc/uBD9GT9Tt/As5vEbCR9xSHzg4
m81RZTu9mcc4Ab+RKoX3owj6tkl7vsxLfZ039XfkFAKnFA/6jEw+n/yJeFHYhU2K
U4Q1STc0FaadsPVnNulDUrnOXliLUi1o1NeVXSqyw9evFtUX3dgNAbGjnhP439pP
2rdG4F/MGp2lKkkyz++EKwdTfoN14n3t9uxw5z+6rL2XbGRaphRBhpNr4LfDY0y3
iAht6gq+mj2+fjZxUj/En0kaqAxeJIsJReCYPwB1Q0ANWM8CAJ4Q8oc35mASn7cu
DgLeuGC/ESkxuQ2v+Nz8NGrZ3ZIhH02oI3UXbutlDA5jd0xOrneqREgyoZZrby7l
Vlo/sTNXo5UIYHymwiv0+RzXI0Nj8IWrwT/V839xczlQ+7QFt64SqZ9jIZ3y8KBq
G9DrHDFDl+pIBKG11jG0plCWLsV1Uim9s3tBX3ywS8UFggsHOTkfvjJ6PFhlip5I
gbfNc8cb+O9MMfNNsNuwc0zHuyB7gn6UaYnggcg5hC0/iaB7VMDNN7auWpT8nH2W
aUhDDWtNJyztb8rBjbfSQzKutH+42ZyBuigBuyJPuNVd+/K5y2UPTSR2ntjJEfv1
YO40fBiigUwKfGFg/v7O1+vD4KxxYfi9LqT6gzsyfUvlTAXtAWfyL98ZOeLWawUW
IhA/ELCU5p2FTWaoSklu5Y49WqAhqlelGYiYBeL259wOwkvPYNKLbZAIjyUhPUj9
dp5gaqKgAdjCy6dcEDCAzkeVraHsjBhT0QG+ywU3MZ/Dl+G+EnLqyLYaKjqRwyv3
5+sHrsJ5XYMjSekC0zibsERt4jLxXsUo2QiUdNYPBuuqPEKXvYLfb4t+GOj/48Zb
wWzMLZDE5vBvr7RoDTFe7j6/FBtY9PpqmruSVhojorF2Eyq25o5Bw6oFQz0CB+vA
plMA0IhfdT6G//quetlfdXF/aVImTDyx7IPDxfjvgJr+Z/+R3TPQF8s8s3AbNoFG
VRRakJDJiNTNkxCKfKV2en49BjAG9YqPlRXQODgft7t39/jbGEgYoh110w6oq2Et
seTg/caEJztVAjzG6lA/yvKpVeXj5pIWNz86IWWqTLHUATPb71wv/gBC0m1/zrSF
5icKmM9cIVetBc0nUbT5jiMzZbStw49vLEoNeE/bFdaj7frrtm0u82OAOrjHZMol
J0X0sIxd4FuHdi7dyvTWOrd7FzUN7wTEXOwUNj9aKarLCiacLcyNrRdEuAsaUsV/
xAd6SW78aUCF+ltGm5eEnv1NNmpgi+yjDtOsWBtsf1YefifmVKmCpJ3k3M08TxWl
Mi73Dfi9icVp1739FeTuPeQm9t9eJyP57mdLwalFzPrWrXMqoxq68FvEEw6b65tg
uGxYgpu3dDdYIwBwdXkXRWAFVEm8dv5bgW2/Ny4pr2Gzn5TsG2ekofMhIb8uU3A7
HYYGbqe9D7R+W9Dy/1+QqX8f/Uvk2d24bfe99ko5/Ndzol1DpKcQ4kAjrjf35if4
3B08wvjIokXSNQkTH3CLzPl0/n65/vc2Gj3kFsxpQB1xtBD//U2BPH+Qh77yVLUM
mRfWECWZu5A8hSviLVkgMYbhPNhJedYqy2zPl67ZCrKEyLiycIfemNNgrESqxtlv
3hZX4sYblewJiqHNDyYjwrTsQznyLZUjSJUX2LfiqOSs7WNLCPtqDgKg2MOHl3Fj
cqgp6aMiWF1zriHQkeROa35toaIgVg7jHYrO6y/O4KqNd+yesCvetBhMNoddo7lG
jIWxy8mudg1LBPI3jUwkpAQ+MOKwItcnr/xoJ9CZAF43jPq8ox7dink1FZ+X/JyG
DsQNpdzg6Uw4aUEQL5E3tJvuPRIczy68XLtpx7RMiFDUs2MkNNLRbnP64HEMHt3k
nChQHm/VVAOsgJZ1cew31IQWhhI40fXhpiakC6wfd8gm3BQxR2S47cmj1rc80OQa
IoBUfAFW/aDUvE7tkv0sRqyy8XgP3Q51xgcDRrxsfBTarrwlLWS2kRM3kGzeFuEz
hARP05opmK0sBo9IA8WXRaAuMzvTjCUckw5Af8HFvEA4uMUInc7gXmV8Bwewh4Gd
Z1mdBj9M/LHvc9ERQho4i2HByliq3lJCyX6ccBtZHMtRs3YY3q1PG93XEIEYNefN
ACFujWBY1AH6CJi0fvSS9ZFO1h61Z2zBV3Jz9D+Jm0B9BV2vOXW4J7lT4/NRrFzr
ntDKnF47I99o3sSQ/k/bSIWdaMN5pz9XoWgEBoxvr8PFztPosEoYC2EbfMbIvA6l
TNn8owdwsO5H8f6+uwzuuZxtopqtrfN1zM1Pulj8zptpeZKWJnzE+GRTB/O94wku
8Lg4i/SfCBmWDmsT9AsmGiYuKyOKYkIXet4hAHMKZYYWyEo+QTAD//z46NCm0ZWn
lN3FrYFmtp7j/tbjVCIGPP4q55GmpPp5qaBrxMmy77BLOSsHNLXp8cfu/YUo4Qko
auCBdLiF/NO5fqDE+fmncUO4VbTrvBRmpeQDzrARAwI8RVshDwjB0SWw7bbR7xkX
gxfF08qYAS7Zr1R+/90S6pCQqq53bq6RYsg0IFM4KjbeJyBS83p53/p55zU332yo
7M1CGN0T3X6KN45dc8AWfKJokQQVuFnLC2nWYq8GMY+CyQE3HVE5NFDq8hXMWYCF
v7gCOVpgWfWyea1qlMplFCpMgQDaems3fNjaleAwKFyWB78rEuHmY5d7FnJrBYOq
0dhSSDrHMJXscJyIu2h3SE1e+05mpG0v605ZB0dlfQcIMEMCJBDwK5ptFgjMFmS0
lnqisjanOfSXfzOrx3vYluMrs4UwlQCGH0kMNLsIUS/BhKIEMNW06jdNAAlgv9OL
6xpOCtODoBoseijpXVRTYWCMuYOnQAyMH4a67CbIlL/EKe4fpUDNdLEPO4c6glRN
MiJv68Op74Y54mSCMrYdzI6WDiTipOJ7bg0/HzQWIheh5+Mz1KXKfsmQZbpiZ9If
dR+mjuWFuDk/0tWVFpJl6kZA5mPEwGgFJmC/uKJbi0pqc09i1H7oOwoJE6DJcwOY
4EkgwLncsken3C2jb70MMEbQkBtudEzAs08Y8ThwZf6Ky5Yoh+IDsqqLwxknMoVY
0IgVycLWvNd6+zTLSPoFVu5A7kewxJJHqUI+HzN8mm1cz+YErHE3BGR1tFeg5+1U
73c/CevUGNFBRjY4PWheQOfEi25VtANco+rCJdzEhm0kzi1sWesvQb3DUMx8tbL/
JwlSVuxGr5Suw3ecJjXcTVIWgut4dNQNVHDoa3JjHLoVI2iL3v4xwaRLL+pdK2+E
LoWHjT9orLmuWLD50KgUKJq9MDuD3cwzMdcvUTU7yIL/mUHZLzSMOchLPMUSQmTj
DgelLkbqTYckinjAkmTEBOmnnIk2ES41yvggXzjsoG+8JJ+VeksseBI8+qD56m8D
Abghw2/AAFrq7K6Xywfc189GYFcYSmlYNcPmxLeYjnLpuww5XEf3MIn5Veh8XWvq
wc+84qS+9Fi0rkOL427EIyiaR4NSni4vmN7RvvU1oCJIkjDEUqaxl9KVmjlFAd7g
NrzG8ZzHGJ5YAQGZoD3PS+DC0b1ZN6TSzoFGWTV2LStMje9OerLJWHylD1TbQLWO
9iemTLdj6BW4UKJTkJVC5WAt4QvYVTMG6GV79aX3HidP9BP/sPKWOWekL1AnB3Ah
hQRHPu5eazWNng0g1Jg2P8VmLiwBVbC2FHDckgS/8v36Ee5oKbaxRvosaA6J1N/I
T3Bh4fZyGIu8fzhaq5Uig6OGDsMb9pGcOBybK7AvyYDuhXN4MPjeD2HvStJBG01U
AoY7fsflCA1U9Tx/P1D9q3+sbUeb0o0zGwEeSckx1o/87RwmqFqp2w5IHTLDEnxd
nQLT8chZTTpAMIzBQh06RwdoLIUfroUl0isBb0xv4uP57Yy6vfdyjDCUQL3C8wt3
RxdCklol0XybyJuzy6eXALqmVrlpBQMG2qVAwvvT4P1+hTE8Fg+AaWw19Nr5bWp4
T75F1pz7dlp7+fv4ClwWRHKGvOUIWwi7zSG/Kae8cYF/eIPebeWmCFOPUm0QOVOZ
5Sl89aJb548frDqnEF108pZ5tXOXuq0x8UaEn9J0dKjlLZUAAXLnD0NgrGODwY2g
kRlPl/VFkcL0ijFFyHTScclMCrjI/p7Y4DvYw+smswJJOL4nQ+d/LBXiy7ivbhCs
2LpoA3Y5wo4u3gkRicYYJ5EHgoch1dXodSgo+MHFWYsTdNj3+ryT+zdqn00iiTiz
H+a6kVift/aK1g0TkOVXcyYbdbKqHwt7th/CT9SVWFTqBGhiHidV3XCIIgXeMORy
BI7bWx0oKfWe0A9MPVk0fu4Jh7wBd2vujpZk9FzYa5wNZEYArFhPpKKMGFtz3trM
oQ0jZWZNeoo1t+qb9xeN8HMGE6FY1skZfQmoYii/qJCmVB76hivnKI6iF5nP2Xde
MsmouyTP7F5Z3FIk6rD1TZ/dUWAjlG+BvS0UDEKyoeULLntG/3iU/eBt9ynmLoe1
tnYD0LY6Lh+6KsUdgnTqZL2KwRhVfjR4ZrELJfM9hI+XR1YlJCWLTOW+WEJ2IepA
oIN8/BojXlLUUvt5c212yef+C28st9MbTykq5zY7fng67IZ/QqBzHWmaMCiWiQ86
VKnp3WFJQv7ionK5EbaIzzYGb4iytuLUICLdLvfH7NlVHZig5NH8MNseobAjfHRh
NrOdfICRG6sEquHP8h4Rae9LIQZ2zWWMMd0coFG04cnqg1CdpyVQ6ctVwly5zxmF
k8Bk5ZNj7pz0ajN6ocmEYL8pbf2HGZqEqple9FlnD0QVH5IxPPUJrAYPzNIf/k0A
1jVUT5w5H+BTC3jbUmmjSoAqvMAmtYRPvUDRgyM17bBcHawf6WxfNJ58V7ECeyHJ
dDRKCp3gkSOzfRZJhtDQSAPVPptw3Bpd2ROxrqHnJ2Qbg1HiQCNBeQZSg63Z8f4I
K9NMWFyEYayUaThnmifecGFHZTqjk8LZclQtR8YTPIy9hsjbz7Pc718pyPPloEUn
YzTWb6ApFZ2IgpDY2Ba4gQPSKB071rrigY+5eCG/6Snnf6LEkC8JauibhmNELW2o
6CN3KkbGY8AvDmHDSP57wqpgpCdYO2WQK/69g2oacpPLIArIxEHSxyLqLR9EtDCf
ckv5intcSV+rMmgq/ufNtbSbyH73bha9O8BrUL4uqaR7hrc7pQCDanWiZSmU8Nbf
Jqnzd5V7u5YiugIJcr0yNpt3q+qETFQ5Fs8FIhrN+YbeuyVNQK0NktoKUScsF/yd
6it8YoPG+X1b6F0hDiddiO9ULX7vjKsxN2/mxO0DqAk4z7k5fx6hU8fbWs1hBDQY
vUSZlOIit3CntuyswhwCZgYeua+KPfPRXSLAN6JKvaBvhttwG9FHhRnypcOoQEIo
GNtnHL29h7NaO+Ix3PpP7DJRt08fO5zBxCGJOfgsc9N/UO3ZNnTYeB1Vx6ejJHYn
o21Ymj2FUEmn7RfjSN6XfUjAanBm7uxesW/NmLY5sh74Dy0EdbPb/bEHrAnkTTm4
mxrnQQ8EqTjXbJPTsqRQ4Lyga22SWISUJuOPWOyAd/sxCImyBL6CUdRf3Z0vEg0E
f+eeKwUzgOYknli5xIg5ZRmmDLOvYAjaAopjvdXMy2UvjnIYciEmyFHJt7Xgxs8f
DeBKxGFF3pPVaXUFik4T3rfDf9Y3WMMkBlCzJYGbvVP+KL8bJzaz65zS4yTAPTaK
sx1shil4SzNHyrMtnFAzZfusE5n3h5a2kWD9xt5hEMbGZmoFjsCwWqNXOPmeK05N
l2o/DTTdhQpkjPe49dNfw+ink6jpOH3UPMZVEQVtlTH2EedPAn0+OBj5OkyLDovV
61ysZlRuWhBHvl4svkloEjIur/a4Ol+ae0yu9Pi3reZanAPt4MNXd/5QNdq07uSj
2ladXvWsosZga6es3xIRlTJboOTFYdUkW5ZWzwIAwllfjmeWciHS7lRrm41ohcU+
nzF7C8PU8OtNWBsr5Qi4Q/ozw7GEjjZJSqGmeR1vgweV8SnTxpf4+iPU+ZFWg6o1
VnxtOgru/kEdcnLJUH9DDGWnl0zkxl3SDV/3eqqHSmFMkITNaWoJ8R/WP9h8goho
8hB3dL3Z4fs4Mrjrxr8eBB+97WMyEiWd6vt7Mu9+f2ETJ1P7dwYtaZDJF2XU+Q/M
R6tTXjpM9KpQvT5KFvbUJM7sjSJOI1/Mu5BngoWGia7b3QmKCRJIuuEcVxAMgqzq
vkAEiqVhtblts+L76Ca5VspHo4A3dMs2XNfmge0TaKdJGbRAIvIEdQGcwWIn4Bgp
zRg+M6vOKBnxNU3R8VaVZ06Y9K91Xggi/pnrXJK258aycFh7DbMzJk4UNym25LwF
YbzKc5ewePxHqi3X2LO7QwitZugxkrXN8RRGh+pStyb3YI5SSWxOGdUYLr/1Hdyd
QxZHNFpLWO1zXB2/0dueNza6OxZqsxi6PtOU217+uadnzYiz6KfIQUED7dVyOsGM
H2yS8E7FKZjL7xHMDthxnDgPihwsPuB7mLvUHEwtFI2KAXMF47It/5AnNtR5uu57
3wOE+fN2Kku5H6Y4glbkT8SpbcRv5oIDtTEWcjnEx5j4Jh1rEnyVlNxT1VREMRrx
kxx9BkryfgQZ56z4c1qef/Iw47aqjWLBLwOOYeZ5z0od9+FzzoO4Mt+A1NO0xWNR
64+nZ01rOyNE3a0IkfuiARMKGixXlFCqwOiu1RZ79NE+VjGAI8dC3PaEWpwmTHIc
L7fgruryoZIrrG1q3j5rNpg4R8/ILDfg7qzx0GmAqZl8PvvRg5ecgBEeVzcuAXWQ
Aq43tngR5IIy69NZjATtJm8To/kJ9wvov7cKE0MWGdadau3AAOIf/xXZSstZS6zn
qMKGPRc8Ja6jtQ8yJmy9oIbzfQMKDz7xdml6asZ8AiijzSoCTGyHatFtNgXeKiBc
rAFJL2Rl92bpA3QmGqtooJboEsESY+JOL1PiZhqEiUDdhnqqi8adg1E+Rr9yPM+/
DxEDcg8lkQdz7IizGV2eZnv6sYzUTT1zVL/UmsHTiOuk2rYX9lY+bEz28F87b1T3
qRwNZnYsiHgcGGIRAGJpY9nmwvckrT1SDkyYhl6nLz4vGKs069/f5OnCYh38YFxI
2nZCl6OjF0aPNS/4Zl1qK+KC84hsLpSkwB6IwFWCZynEf0HAjgyUcNbK38MNTTkG
oAyjnL/vP90S7fd1YBfkbKYE8eDpt0mii/xMusfPI1y7Wo/JM+41rURMdy2Ejahp
eZzlJ2PiAEUHNMvbzU4N7Ybhj4R0Ct1LWpc6ja/v+AL3LWYuWjINgvUvVJG+ryZA
P6vlZJWlXsg39sIFjbpLM062Nb8NL1FviLoN59vhTfdoVRHz3Gj1oIKN4uVEvcDp
dQvDEuZWMaZxFKe4Ya6IvuBtdxlgy1Qzzfj3RoI/HdpTpvWXPCYuapUPUzj+zPPi
qeXIi1Cd+LvK3cc8xrgQOXeNXgJ+IafxWeTy/jgtnI+DIO/D71rmURZY+Sy7ty9g
RDvuc1Evt67NA1GkA4my5K5Gup1FlBOlJv6vn7F9hDPe5QWjTAVjFycUZslQeaKl
KRDLVosy4eZ9WH6p4qFKK9tv1YtqhPGTNVHKUFi2LPv37N3lckbUUcbay8/xhNn0
KVTm/KxhdlhEJoCTCE+eM2RxQquBHJEafg7AqE4DC5aEh06rkLlUlTYyUV7P9kKQ
ZiqjjFtH/nIKWI4ziidGsfcS7VFSE+jf9s7YPQ1CPn/j9RR3NcFXV5TE/WS09UeH
50gMEKMeGg/dezEROTlFroPIEGIjB/gvK2iU8v9vi8HwwlI5zhG0HrtXmTtjV2cv
ZCK3UuaPTn4ZlbWFowmcLFjNLaUgGzFSXl33yOnBo5cJtNJwPNHdOP69s/RuHJpW
DayCNbfpWUuRjGkEhHCXakVUafWh3l0dH9rPV1KZ9LuJP52qoblUJWzEU8fAsUNj
A/GDsjky1r5SbVeRqoRTzBCpItXMYE4IzTfj5uTn7kJQDB0uLDba38LjrRnEvuC+
DMW0nthrSzyRn60RJ2g0MIUypKBn7FN7Pla8zDhCUj13f+YHAPbsf+XyCrg0ndS1
nOt/cWVEXOxoBH1lhif0rU5eXK9PS/wgFRxoE6jRfYSQF76m9nk/cFRcmR24GD+q
Dxwzv8Hbo0cxS5vU1ghvz3oZBT7Rcj4gpujx5o+nxb+FEnASrWi2TPvVOokm/+6b
1MqGIilLOMRhVX2FPlzIdd4+5Pju7JJTtIDfvIBJj5xuJVRAlF/0c71j/G9IGynS
vTrMNIMsqkvJGmpXbGL6JsQ+jclUKXXTa8IXzU+/D+EnVmXKLRA7sRNiyy6LPreZ
p+GWDuHAwWQeXaXt3g3HubyonqgSm7ZcEkhWjUkaklJu4R2QbCzc01uuBMKYxnGh
Zl9i4UT0/bPYdyR4Mm7czCbzBWhTvfyVCkwcf+PnjmCeFx+fgRcFgqAvwP/DLkZo
KkRhkdOcQRlE6AbNQ2Z223QfOmYQiX0gdci3PGiZGiEz7oLMqdI5/uCRM1SSYaZz
NvXwSfFV0949HcZImhqo/CdSzmOQjzqwHzN69AW5IL75zuokwCgE8HZ9H7gL3eu8
21PqrYN5dRqb8lRbaYOxaGFO3/8PB8P4LSks8GdF7OZTrFiRUYE11netOBvkasmC
OvCgSjrLmjngul/Yhkkmnwq9RbjMYrYa33p+DarNEiosK1zS8Tcy5hM97JaUg8kj
G4CoA/KnswG8ovafOCZWfj67wMm8TuD3NkL4PMqTRX9XRzM1Nstk84D4pHAkq7mz
EsmZ++XeYKQd78YDRladagUgTa7J+kTtWyKPsFst1rjq4wpjI5t3zfOdooQA1GmN
toZPKGkDYkQ9e3X6B80FqZpjoQMw2jWmoQ5UZAN0WBtr1F+JVHVowBJrkvbChw95
1HZ+QB1jj309IpeRWFe9taoCmVsBR5CU8wydyb4sgnHadamC6r47aE+4WzoitpBu
Uib9VYRpfGh5CVmWB8R2dIktes2cFwfnhurJP8BmVtGLvWiOCrpzBz8byo9PlfiX
caQOTRPZrNmSbCYjFIfzjrBjWwu1aC5Xe/FWKz2nb6DqaA440X7bHRlWPwawy0DQ
OO6YdFukQ6YJsuer5PvAL/lxN8zHk95HJCd/MHSuj9l47O/CSs4D5JXE1VOAYSjz
38papq1Sn9DdiJ/OkloVrTCtofOeQUJkZSkVUuIhtY17G1UQHTuBEcHmSvYsFvPl
v/T58hfyAGL+4N1XCRJvSI81YAp7xsx3LTMj3oA0PwzU7/wno8AqfyPIMdOsok1s
WGFFbjrBg/6kh1Io9YvE8nfF05U5Yonix30y9+6hLfJo07BFG77l5cMv26S9yY2a
k6Lf9+ptDqXWYH/kPRz5e4nzG+Cj1KEIBvHnLiTY36sOPr9n7F1gFFE4e7t7BrWU
jnadX63fgV2+CFxRy2jJmMb+SvNeCyDeFsfmiRe2eRNLTdS6YyR1o0IrgSFc4zo9
Ux86CxEtun9Oszq0ASIhoXM9wpDU6qNVyfXjrb3Ym88ivRD35Glrdd/CqEil2/Yb
tLpb1BP2M20EQ+bL0e/c0Vi6GKqVVVwWHkMJm3YDs2ZJlZFt6CNWOUolGW1pTujB
ra7Us3UUxOK93RYigqRgE7t4doLs7XbXRCwEezORMwGFa+5CzdpvUxZ5Y6jV7e6Q
tiuOncxVZJY91/pBMPLxN2Hi1l4s7BBClT043u5OXLT0XjU+Y3dwcFasn/wpbm2j
ARrW1S3BxK+gWcWXepL/CLwW+/1/XJnFVLp/rWTqIZjSqyNH7y+kA2THyMb93Efz
/ve1/yHUKCN5BWyTpTMsN9zWNRLP/+SC28I5YTUivxRJPzHkyA17Zlz5AHyxTUXU
KQNqlqmsm+ROB23MBZJ/NQm+GqBBfw51oJXFO5D8/gnXgG192T0IUhDMyni+Z7Ff
AihIbvaoig9FaXsIBPSU5PWvRpSh6PgiS6GGhw7YjWPDnsnWY8ox0EOeCLelcXbb
5w6VNKJJ8WQQw1U0AlS0NGYW+P6vG3yLc+JqwZr7eN8yFpgbV+hkU4yODzZbjYgG
BXXiMvSHoqCd9oFj/U3CXIUEPYMr0Kk9r5gqhct+f9jB3k5KjNE3chSyt9TbF0GH
NTr7IPtC4b8/dGIwbNPq46MVYACxRLIebCBjMA2IyQvcDwrI2usy+pKEKOq4RMzb
oB32JlNDH/EW1/yx2HAkn8+Fptm1IjfyPYmUT92mMrZNowkCu/vSUfHrAIUBDCQO
ARi+DpJyVBdNpsAmL97GubAhRp1MbCEqn0aQCWy/AIw5N5HfNK6zVjqG3PErgM7k
9+Sd/kXgmJTOOHtlmKe2xaDi6/IlZUFUhM5uzbbwC/0ycRK2ang0W4pSSQ6W49tU
Zs9De2mUFjdMgRWzSBG4r/vGnU1rasjrFJhsvhr1r1qnVNYiWr8rl5bniV3fvRWX
lMSDNiJGfx1Sm3d3SHfgNzCA2CaR9Y4VvF7eGbKiII3YxWw915L9EfZSEtUu1kbP
hgYoTtifWbcMthW6HkAn6fcluBnKrVRppL3qRUOD4o5BLP+igPUiw87JGLbjH6q+
zoEwRrFhStPptVTTxvsOhAsSp0lfan0Va2UhB1h2hjcTEfzWYebHi8y4JJk0Xdg7
W0Q3OcNqScm7aM/CC5iSKflSisf6VaAxE0g3PyNDfpacVJBFTuJwLe0TmQrnaGLF
M8pimy4iMy1kVAulHm9LPsxXfhgdyvsVDiAAdUZsJQCFmahhf0wnDtT3jpjcQHUt
fXSi1zq19UPD546/CcUTNG7j4nZW/zEO6EAlUuLAZD7sSdRF2iN+/81sXdSiQlKz
8P9RVfIkbWclG3kdLdHlpl0Cvor4TnUk3VYMAQ5/5lnhugZcVIU1B5iXuE9yGFrr
YlakBLQawTxXFW2ho4PjMCVdTg+u0ZMFZMGHhLySQbe+XvyVJY7AgQNKqIaTjyYm
T9gM+q6rB14OH1BuJTP/40VxJ9w5moRZEcKo7G7BEPJ45oK6C+M8fVTzR8NFq2e5
PJppZ1AODl5UDs50ynPJb/KQ67B9IlBc1tQT3TkAMVlFdOd4cAAzYVselKq5EH9r
wsHjUDAeH+Mjg5yRN769mY2boJNHYemQxAZzaIYmCzp+jxKTnZaZPWCrgXNcWL+w
6vE2XXQZpoa8KX1IbXITWKSLMMPRZ1eDWU2v5lyayJilMDmpynqL9+jr7ecRv5Wj
XS5+HIwg4+AoEm4px0rMx+1uwysO8WO2umd/q0lDzDr4bPuQ/mcqNGBthRkJwyJg
e5GSOe6/COixnMCNSL1vvuI7QdENDBx/mssVI5gzOsEBuo96JF+Mc4syCWjc2BLe
b0GhCbLMiaHewpUwGkTrvDAayiYRl3fR94NkWvNBNfUCzwhHiE7jbgJbAFaq6/tG
nO9Bf9Zw5U9YYUEKWwqBVHe2YNTcyla66tYevQBqjOgmKjh+5i7H9fA8bUsASEM9
Ui5lG55Z3ztPr/y6lK2ZnE7tpPwuywdWWSijCFh1T0+wsfhaz58MBNvRODANSy5L
iWBVkyffYHKS5dLWQGwPdcU4stM9ePUNckBMZ/LCa9hyp8L1lz7tUTYtCWhH/xps
kTSIoDublojSfZzucSH/t3PuE0D9R7QEpQluTUsXQEOi3Bhlhmv19hOZn6RTnwTF
PoaQ5R20sIogmC2qQNMnJgIycYkM+D1t7UjoDleNSTUX9qf4pJKM4K0M/wHNYTXp
mQhYKU9fRjaRaZgWXXWAR0f04g0MF+/Jjm8oEsD32MIea8nRynMm2dYT3F34PsBA
Eog/Vp9fFci9LG53Ww8zXqrFT1Xl4Ickob7yCn24OT+TZg3XOp573ToetZAIk75o
9mwmzRrfYl7Ez1T4zScfzhZTNonKUHLiq4QOeaQJRQuSKKtDvPr/i1zX7xIL8nSV
z8tdJuymvjLiS4Jr+Mflmn5KcqZDhgH3Y6BhVYM9Np4AY1wsxnj4rgs1aibXO/dY
Nfg1FxMXOaa8IQHuIWu9hMUTewLY4gIuVlctaz1B+mzHad5QlnmhI+gi1DJswBNw
vYSUmmOYpShnudNmHisGuyg/sbQ8DzMRIF/fHjsBbrBDcYWvYWuFL0FYRIBnahGt
490XnN0H02DwHzkQfLmuDHeMvUpgcjzz0a2tbntNystmMWsXRxWczQmVzZQicCXc
8TWiEZvXZlqeeJzfmz1opw9gIclwzLuu4/iKbQqAY0VcmsdtwrbqIM83eoR+dzuE
VUV2LPVWWyrZ8xaErK0WteL2/JfplwCUR24NNubBG9ClETL/4kJuQQyDyYAPidOT
KSv7g7xm+wOX2VTBxOsgCi3q0plAkV6KmJ0NKavX2+Tvj4/GpCMAKVuxOHUKMJtH
RurR3AUkSaENNssAxmh+9Qp8o/5vFVy6hhyGXf7ghZLXMHF6tot2u09rz4B3TGe1
WwwlvCBeeadKBVjyjQcNCTjKCRp+hjBhvLTXr8BcamZWzxE2fv+rrUqJ+NKaWA+n
etUNHrJXVGaVIl5Xat718GgqPrP2TNMm8WpT/5Rzl4DX+2F/dy8dRos8gCt3NX+R
MNEI+UeEslyU2j6mG7C0Ab3D0Yfz9W+/O4zaVYpeXs05gD+LJ6x23A9hP+VfSARo
n27CMSNfx4Ogxg1L3yO4QlEE/ea702NAuRPj7ZlQNuHBU9w4ZxNHfCfoo6LMuaVa
4qVgpsyyyA2SeYYpowt3gw3V3NZ1BtHJsGc7O0G4R1AnJwi+tPhe+KRrz0MpZpN8
m+5r0wJgUl1mi7tGb1chzDwesrf+Y3Jzpe0CeQpLxnAyVCvyQlTrbwHLemcXNTnH
0iewiCI913pxat23+AZsBMc7U7rdXK7RKpAgMNyKrxnuRXMjETqU/IBRm54xjdKF
GYU8DYhoCEj9yXzJCfUa1UtxomIUc7QpUJoARi3gcTbaBfwI81yFkr6xGxP/MyFy
dj/wJpQU7l8czvjOgSPCcGzWq0NhVCwTRpTiHZfcGCT6b8qXkxSUfs3p+5EiUNNk
ZgcK8fdn2Y7FcGnQFHLcmqtcfAspM5lF1PhO0lYvTG6nrI22PcUy/TpPbMKsdBeo
d9skVQ7yXCAaBABoRiKK3TU8DBT9JDtg+v87hX9aehkb0wUqTEYzJAqte8MYMUWi
IJXB8jnN7xjoRI18goAeV6bjZyZGGfccUf/P9wrJJrtn0enZu0kEQFiwycd4F9Tx
AjhhEspGPYdjNfj/6dcqBIr43qv7gG64kpNwBt7hONcz2sjIOyoah7B1vUu6Astp
4ZAj0YxABdWFIid/97RJrCgCMMEzT2lOPHE/2Dqhlbfy8aN8asijFo/7AM4IKGiv
3wF+kxLn55Q1LnDkWvsyVrxHMljh6z2hY3O16SLU8Lj5ndUF9RMo2G9PHLc/fH9N
smRnnnARPE8n5MD64ZCgL5a1GKze+scI9kpGNG7bF01OK2IjDk+/H8kxsFrqJNSe
m0kQqYGFJmBAxZEOxUhSbtHObqE992/ESCAzQ+25L/Gp62Sy+p1H83hPwMcx5Juy
tqyr5CVL7xTCBooBsFSKztDnBBupdf6uG5dYpuV1KE+UCUq8TKpPSIq9JYPeHyDz
RvGYnUUEydzBY6/Lm0zn9DB2sw2yQIXoJk/RtvvPA0WOPqpzSaEml9Hwlne9KIdK
lgJTTuSYiN7b80F9TtLg3eYsCqE2pPsHzbwyis+dAiCzR/aCnAYKghmG+yMUhGx2
YlDmgH64dPWbAKlvyU6Dm4AYALZV1lpsYe1yb1Dl4YwIuqTMPf9Rs7mZAmxzYxdr
EYU1qmzF8e2OdwFGXQoGkP8+5L6z7PhKR1c9Sy/sqk9xJq1bGkyRvJnQNrfmydy9
fPfP28s2bOgv8fG5z0DgVkD7QdoQDEKlzTaJNxpRmPUPAyD19B3KKDjaTBBFVX3q
WV1jbFYxF3Ko8m1+v6vFclqx9W7cgxstXf26Ir8Zft4NCOSV0UbdgBVVVPeeMga/
tbnOPJw4D3RDQDo5YuOKGvlDkJyDUrk1SK5K8ojI6M3MfYXSEfixImsvGdR3g8l6
FqclKTnzh8hiZI4i3SGdsirF47rB2kDiI13f6S8mSY1hemXY/W4YQjkukRd93Me4
v00yYBamMJJCqHakz4aVnFGKX+9JH97dGJAcmXF5H9VIiYmO24VaFSDgNGIQzppe
vizOAunB3en3V9QLkVASpUVH7ADcLOGaHOee05Aw4MdsgzsZ/Xu8ok9Zpw0HxHaJ
bw4MI4bmmD1jyRQ27qJ4PEbQRjd5DtneBAgNsuX41XMFsk8tRGCbuUEHUX4Z/bX+
iGAmaOF7R926gjIm3dCDOeLCTsKcS7bCaFDvW/d+G8IEbsgCR2xYh5GB/c2oey0W
A9RCjddyiYvJt3ouA/T/VEyYyrpmrcK19yXTA6oVY4oB2lPkoRb76yOGtTGA/UFn
9zzsJvOrkRqwDtar/XSiusOOhT79gc8D2KijsRL5ZfDvsNP3RsbNtC2cEMq2XcJT
8MsRDAC842lWLlMQhHCW5jKkHivSRHmMB84p3ySNAYpUX3d112UROI4ZpkQ1/zmd
Qg6Am9vyF6bPPB0dBIRI7CXPax6iHh+14FzPiHswWPLsMoyNDL5cuxDU3MF7emy/
uM5/nPwHNIsEiDpF5PNjeZ2SDxXM/lLucTe0+V/5VISqa9bAsK5TgnnGPAC9SX4t
JmP0MF6PzXIK3JFBsLuhBU9+Ufw+uP3Fo2g87/kYAer3WuxHZ7l2IOtBi7HMo3li
5zwn3e4JrGZurrVSYqySr0xZyt+noEgZJU75P19vwrsffskyNuVFSb0vXXCROkzC
KM/OkCIGslCOyk3r+VhWP4VV6P8jlRNV9BbXJRmJGbwjRwU99kginaKSsdw31DEa
5GPGPAVxnMiaU/RX9M4wFJ/0LmiPEdbqXAmDJLXYuaeY3VXpdwZ0sSXU6agQY4yY
RKUqZlNWt/eHOvXUEjmS4vpdQPLuDhNsz7C5tIRyTa3hSFigJ5HHp1C4DU45ko/V
qdKoeOh4keIbohq2TQiQr7fv3hw63Ohx3zO0ZdTM0X2qM8EbuGmtpqkm8xgjLM60
6KhcTsaWn8Hok8MtCeFf0ca/5XbLK5z65VBfDOmxjpHWEW+DsVQnUziGbhs32U0V
wQiz0Dj1SL3l+IbwW2nufp+egORSwtvkQaqon9vhsOs0BCM4MglBH6WkHQwnD1sS
prjnLYE8csjMkXqznxWKD5Z1Ou2XJoqXrxE8zdg8vsWnYz4Dv+VnWmnEsaA0LoNc
UzAW+A2Vi0P1qXHTtesQxF6llmbEQJeMx/gECdtTBKReI34a+E+6kUoPDYw0PUp5
CloaT2PPRzLw0tIFgK4ACVjo40imPEk2E04uWCvXt7awaI2Hu92CknhmJyvLB/2I
ZuU5ZMO04ip2sUE+00eKY5x8xzEyKnzxitzzfLm7oicIVxXI7tyA7r2gw9ITvkRI
u8sjf131FOy1tpn+avATdiFcC6mIyfhqCA+nQKnVyBIoWh/pzQh2wpIFDjV4OGvu
u3jYnbsV2416CvM6dhux8n4Flz0JCNnyoQrAdJQygFV7a3FW2DuYV9R5XmT9kNEa
2jhPpjbv+uyUw43zLChetg3BT3Ux/nLQ3mrgPqPnAB74FYuHw/s+AClApv/gAuh0
2PC8nmU/BJfa/OnNpSydORMslfT17SmenXMh9mgeQCw2H0ByYXUsz3ya7SmY+G0Y
QGbLHLDljgmqJaZRRszWqybuwLYknwSWDjbboRwLkiYtVFIiw60RuMgx3QJMShV+
2H4FkUTvvyImGSTMb2JGb5YEg9RFAQw+SUkkrwlYAKCF4cVEdhTdEa8DKrfoA0kK
x1VJjbh1f7jXF9KaDXp/hp1Od2JCyRu4j4oalNDGQLz2LJevIFWkmZTF76VFoHP9
i3k3ZBfnu0ZfmTf6Ux9DoB2XVXDSci6nKOJO5Su5PF3c1LevvgW3/4RzptnO7Kjg
TSvwHUQb8RAVe0WRdoKiKbeHqMTrcqfHin/KK3mEqKJkaY2h+AlDHdBlpmkHQ/ke
3nxT9UoHLJNXwJhh2Uk3sPWeP6ss1upDe1Rw51Ud6WZqa4IFq+hHYALagY38vQX6
EZ8e9ipSaAaUzPRLo61UHQv66McrLfL8jEaBIrx181w0IYchYCu4xtNir+CUFnfK
Meb7n5Ad/Pdq/1lLCUmd8pqK6vyRoU7v+3pu76TBr4e4XQtcxXlapXK3JzrqH5zE
Z8Z9YwRkxhkRWrGM/U4nvL7bD+1l++xyt+BZ4p70pTMzgiebMAbWniNSBF6kTTmC
q/4/L+TWWLB3wlt7SHyMlFxVcXr5NEGX6Jr+WtUDvqxRtYWNx/ZVL+aDjQ4rSxad
3potM4yph5GGB9nnNDySs6KBZz+67oB0bWHTUzGpIKSw+tpZUkbu0SECLBZLUPQk
FpfTvzcnr9YJ5s1Dcux8/4l14Nwzv+mKPxa5C9I/2tT5iV9qzUePiqAPu9iqDofX
bXuEBRAGy1olaXbOtIlQmWzHlxGnaf2DnJy4ksy5EZv6cgEYp8ihBDrtq4cd4e32
JVg6NMhKBAL0P+X26XITqevDfHCz/4CIG5oTFgH1/EmeARX0nXcZf6nAea6g6h/p
x/zUwnPYefozVo1jcUQ6P5djeHwjWeCKA44uW5ZFa9uvP3cx/IzRTelTJzM98cTr
SFWPlr4fQVWcX0DTx1LGtAv1+DKAWCY6xwHH4pMSzyhtvHQxSfj22z4WUovWqOZe
Gjflfahp0FTBH5F2+iICUpuE49dMR3QxSiJMGw0KBzAt0WoRqmTT7vcoybFq/krS
klyjRC6Up6Czk7LFCB9+lQ1LSN3gHpPsZrShLAP9iiGGWMA1EJs05NV34UDtJ/gE
aTNOUy5Hgq7QZ4Fnz0QfCh+rWvIca0UnMBHgw3RN4YCdR8CXHcm1gJ+jrVyuDarK
bXahLfBKQ36L6UCTB1YYSa9Onht8UMEKm5d+Eqz1qzCz66+oCBvzz0+iOQit2J7x
oE4BlfT6Y217JdOTm8sxXyDU4kRJMwnjmdP70VeksWaLc+i2XDimDLwcV8meOAHr
ZCuwjBvF+1M/9QHRaBnk1n7jCw+to9XGUg4FYUZN4mdycrCfCqwZwqQbMKz+yBX8
Va5qnoHp0xJlw9gWsaRJt7NvoM3D2OVI++MbDhw+YKzglaVEELCWeaB4UrlGq4Wq
Jnyh5i89dPrMUZ15YiyrC11oGbQikgSFXDqtEws2RkYFe1CS+pndYbL1eWpqz55a
ySIAJdWQe2JBa2eIpTq1jlktbsye1h/tLcqjwvVpmuglPh7lVIJO0Kn9Vkpo54T8
/KEArLcmNNsxhzFbJySzi+W4cg2NgCTiuDSqacWv2VMKEo7HXZbbLnyYlak6xp0T
a37SDLWZFn/Wr+nxj51BKkx/KF2pDC9DAUtTtT9Hj0K+AJgeoU95VHGgZB+yUjP4
KNOl7AXHxsLGSAUhMm4cKSexnhrL6ph6nmL7N9AToUWKi7JHMwNyCaYXTZVGxL5B
pAv1FEH4gyR/2sYJiytO5uO/OVyUGeoESqpBfWA50A6CEhHUEYL/l8K+Te2Z6/bI
InIzleSU5nBjXQS+XhMyBa7rdqkubDnV4EfRlI4CGaWXpX3tBUe1po7t2M+PJXsB
1Vqk7+gXJNk6SPjatndklpTYzbmdd0bXjUYHd46HuYOE945x9qxFttUk9npDt3Je
7FFdih3ydZfuztEZeYBOcpr9lA3oyeXXiwHILNnKCm+u9HcTSBFw6SJEwIf3dnXQ
JMqLLHQ/k1BYT8TnI29YWNfClJKJEfxCBgSjjwHtksuLLaTUz94/bU5QvI/Q2/Ww
MWqYkHDSlWqlcoZtZvHSOkVyu6LDNR8V0yOAWuTzL0nDZqLnnYSiiMEue4vmzDZ0
iJWyuf0i+ccvRiVxVOFmvV9CTHpb7wkf2D1ydKVBcQR/C7lcxnsOybRo33TID+s8
VUw1QLqoKiULNC1UCQHxEw6yYnyiCVnj+Pv8fERsvOIa6QxDvmUIA0FrIIdXUv8H
+UApTtWC5e9c7O4wYsFvg5zCXFNamvSN7aFToZWQoK5sqV8kgGBASoy/j81cnKIG
R9bn57kn8IcnMFCHAGHSXsqMDKmO/YInhRrg/WjXUKG2gYfBgi/IEMOUc0aKmcBh
Wj/E4IM+jp61YUePPYCPYXNWZuMl8yzS1PE3pJueYbb/cHhy7jSaQgdbeKd4QxGb
qgYKVz+nmYxq4Y2KH09jbjbmOnN9cYhrGF6HHTyVdfKlvXQk1Mem2s5qeeW12v1p
rSUQ9KiawKLsyfvESWCJUb2sR97CUnxCN1TlMCkQfpZaMXiVmo9Fn5VlvdEtdXUz
jmgFKT+xaNKJ1W5dz0ufs1QiVWovN9XYw9v65DUfjB9Dd9sayAQ9nG5YdjgdAzr9
6II25mOEN6GLF5hlEumo8Ae5n6XN0xjYrOwF/Z0mPbx57XUUXsiPfxHJ431AqEDy
mN6sGflZPfov2NOmgfwJ9Zi3ZhqdQbYbJCV+IaGn6zkIogijgjB6qvFRzKuxRt+6
0hRC+yn/+kP5Ay+H69obxzMaHOTmIDYXQ2eh0QpFPGRuUCNEX+55opf8VgWnsz09
5GyJaCLAt3nlMfhbdJlLS+VIQCg+iMhuNAC/JKNMXG19ZMkkQUr3yg2Ami+uvxbL
p+d8iR3Q52pQaaiHIqtxaS6s7SX8Jt7tdm404l1m1E7lyv2zndPO8QVWyXg4TCBy
tHMZssgd0gELCFvnifAUzvVTDzONAfHJpaPkzJmdERUTXQJISEAz7O6yaC8EwOkx
MYEjNmMp9CMd6DubsHZWMnIm2e4XgSP9Q2SNZM4Z4YEdD2qY9NjMMgboTjtnj2co
b7TAMJjW5wsCV/Yaep2Yysisrbo/3TwjglBcFMYpuGtnxLceIhdB7zak3amCkD+K
OuJ8+39GDbBnhnUED1VwASnR9G9n5i0FnLGJCzQNjvWvgDbI41YWI0OHZ2gN4Up0
hJgg5JAdl7+ezzld0BzJlS6alHVQwd3hvr6NVUy/XUB+BxLAkfVMlRQPQOPwAeVj
PaeAcvasVRrJ5kZLqo6t/iOx0ItpwWoU90vu3kyk5jhQuY00tI8arv/RZhEZDkg7
4AOlinmDfp1H3ukmj8vKHjc+igOMtmFEO24KEZaijlYMWzoGuebhb7cSK6Ablame
vno3rRBTUjs94SN6tbAN9d5ir1jylOZTEeQYQXqUr4SkqOHyt/xQ4gRz3xQzAv27
tHG0PJvWdxd70x2xZe87yCpiz+/xo0KgjbdobSdqhg81tRi30Mgab6E1kdNejzMU
M4mBHA6BearyB1qtRQeNfhxNnlZB35kY/6+TP7BiHPcqNIdO3yWCcRwxYUQTYqFH
n9e4L3rp6VChHUa0whi3fDZuUWmKpYP/qabqlLES078TBEDv/zHwMslGsy+hdjy5
Gzxztv5TZLZOn+Ma2FczKuGxovVSbjcD+0o+DvadQEmf/tDHl0tc5Ng5GRtlY93j
0qqaeLqGyTCVZpsVcl5zRCgevEJRsoWnLWxtmaC6as0Ffni+hQ82wVAfafb/7w7f
fm5hc9Pxf0ckr58vwiA6vIkHbbW7LjfTnGSQ2U5Z6GZN09ib3FWJNivGui7u1Gx0
Or6SXPbXzcpEJeRPGpU/cXc8NOOHPmwoFyAc30y9sOKfkbnZn1IYoJ3rt2xt8lxv
ki/GCKMj+fHFazgKPY/WP0ZsPGX01zyDjBmIrBr2bFt/Oa4M37lcsoxQaV3beY+A
vg0I/Hz4TFOOIYxfYb6sUECtCueBP4m5ELpgTlhfuIKuHWiFDM9FJXV6LZphlhu3
8JgX+VZ+OGSPAjPMp5JafcF2WuB6a7PCgD/HccacLo4QeonBba5hvjspJese2xVg
JXwLHTQ/1Imt0HqqZf02YLxAzSZzlINpXtxg9QBkoTXUL/k6qAFBVmI7JKcGbglN
4V4ajL/1hXM7XhUa2J4yrEMdHotz9+2MetpHUZJZygSGFmQKRp+QIPFCF2sLeybd
CiY2TzNiDG5w9Jm/kMHN3Za50lXbi6KiiH4PFmADC+ENAIyQuxsDojOE+hB+McTz
xy6/FeCoEIIbt3aV0lCRPuAnYcpATZQeX5D98O+lQqPZDeiS/SCJKB0RGwoLi1bs
hLWbTLwBMtTfHJZqP3PL7iDFN5gJ0obYiHxV8FE5GFUeqtPwgDk6pJbM3YLOeLW4
WjI/nyOmI/Fd5HCcwgq8ENlDkNzPKbPYQU8dQbc3FjhuE91XlzIYscXI1tmChfy1
tnAzrJPiTgqpr/5Qxx+YaUhGm6MlMNc8GErKx69YbkYyPHV6Rwd3flavJRK8J8BT
7+TBQqMXHxC77z0yTYiFbJ6bK+4rINCm4tKo/+LfNNKQjKP3vdFn3cjyjhcUFees
rXQehW88ggB/plFLx85YNu5hjZxttVDWTc0QTcbg4AyHPDjcFoeVDH3xXWwBmleB
idIgd4szFMPLAJGwqDNFDu2SP3RNr1uP60GzEWPYFyDqFcR2oKN88JErScau79ZU
Fn+h4d7XGzugmSJa34MuPwmb6Trx5GeBLiwibLMECrLRuY7pu2afJT+Nvk5a7NcU
1deTfko5YUmjWp8h1HnXadrfFJ69ArKXxMAwDq9qU+X3Lk98Xj+hUUB9w+AWdBZZ
YUa4frNGqusjYLtDIrHuZdJM2JizximFqfgIptiC/kUlhbvDgQVBYb+cNyM4EVJX
WwOZmYxMAhNJLNyaLWlHRiZnOZLX6sEUqzgH0o5y2nzAmGhMKnrgOyW7kOdtKgIc
miMV6LtZQ3C4r74HqBG3pWhFcqkGFVcM+T5PeOp+HVzQtLTBpEmpLH6rj32fjxJL
QmK1C/VNpbm45YozDBaBNqzwFmUuMz6JFRQRWCtpy46pTwjUVtbfpRSItbpIc6bh
t08TlIvx45idTN4/1Kw0osL0VN9xhH7qk9HKAgQpsQaAl/NjzxFjQTKLTUb92tJh
QhURlJf9sKlrgipcn8BkAcGPMY40ROgZleKYyDxvjuTRiaqP6zRFUwdxApNeIm97
YDIQjJwIFD+088KKDnoofWau1Eb73mbSOaCxuYqS+px6JHOxW1FhbPS7mu7qHkvh
rJz6E9P6M+8eEIRS2Av2fNWcLZkgkAcwE1sV8T/2ZvJwjjM8EratJSxpIP1vKGss
LmxBpHDRFV/fHAJqCPwKnaPeexX+DGWCbmHfTeqwre0AaKMXkutPA0r0DGlUeVV/
2UvSOMiDdPLivvjgSkCkb7I2TwmNZYWQ4G+B86cuF1AiGOBdrmAN2U1ihlxFxRnY
az309TL4rI3U2/T5AIqo7PguZkYXFGHGSgz+v/UkRvrnEy84KFQJ1eCJxzttsxTP
cG+L84f7NSFzihU2o9yGXrN5DdK818EobNUUZIPmrRc0HLEfL7huJYIyGNud5vvz
DwLYHgflsF6COYuNXfFhg7QIS1+xmY+46go34+ujIr7hI3Mfz97cKq3v9rb3wK1J
rUYMoSQDPu2HspuovXM2OGiHoVi4iYeVSiO+k6RqjBa3VQLLPWkM05kduEExMZhw
kNBdEaoPCsSnaYUg9Q9kmQdBZMW+qWZHalsM4kElzO+LlQPUjB4K6ilHatijeTYR
CurJog9sHOAX5FHd1rvoDzdlJfZbP9jYV/yHvdnbIjc5jxQOZRIRrZS9dqcYtNi0
IWSgYTzeXrvpsHZsFjNnl4Dox8ixifxbDCNqEzgavwFsNYg3Bc+vBkwhsMkP7uQ4
1U6SH8j73OqukNNlAkDe+93K+a/TlnihDd5TE2cqKK6BOJs/lQJOYz6FAvecLjyO
5kn2M9qqA26zOHZiy1J7ORtvEgoq9yn5nWRfsp/MUf8/LLY1j9nqkQ9Qtef+dPLu
31V6N1LDKQkXt9ICiabZ7Bb1iu9on0lKrWfDiGHPaBzRZWvoqb6UbimSeawDdHm7
wf3Vw5CzF1UzB/FSGncMyVY1bNxUyx5y6Dpmmah9UiEbsxyrxYHfLVEmDduKUj/8
fvYQ/ChfiIt/7zUoJJVlUbUn19W1G4jpWXAf55kMWJIsxibkTSaivO1QEXjoa6XR
4gyHYzeY9mVzvxMesDDoTGc+aoXlvrdvmGluLO5dDStEiJLUjQSEG7MfvNNuD1OV
v6GEfpT2LeckoxCqwwuM5qBHsXadM2CMXLfP2TvCdp0rh4EjMrm5VYaBYyb3Ow9X
0HxBoMdQmhVX0WBukGC9CZgrqqAW9DjXnI3V0ATKiTQUlQ3phppZGz5Oi+mWSQnl
E/rOFPO3G33/rOiq468GAZhAP1ZO2MeUBEGN8i1U8LgPkpY4LHiRdirYirqwmwhF
SpvTW4q9l1c/rSdm0NWp9eWfJZISNzRHB9/bhi2G9ARyFzcSPufO4Zchj4/A90K2
QNen676Gf9QME1CyULjKOyQVYIryknNIp9FoVE5vbnZpg3DHlo5yfQAwYTzCTtWz
9kcLiLmcctU3/9DabVJ3NJg/IFJHBUZ2YNFJqa3r3wjGrnU5TCKYSGrPKa9P9Vze
Ws61q2GvX0QZQv5Yu3W9g1Trs78GCF6fFCw3GEWYo5soS1/RxvcvGair7PwFd74T
wdwxB2L7Lfl0LAgtG8l249QQgAIUfJjKPWk4cC37Ap1D0SbFwjrNCG5vzbck7gVy
JTMsNgZarnpKu9cP31zd08lA++D1kNQrnHsYn5EGMJ6FUH+ox/KdWY+Idk1RnjW5
/viGKO2wSwDanQEjayQEUVcLqxIhpW2HJ8VVs58R6MvJSPcAqaHfAEaLby+N6rX1
8a07W30CPZJTef9YfwQYbp91DbhAw9ZnMy53GJphGhPeBN8UlltA2SjL/ILsPQFU
LIrKXfDZwIk21xlnpdmoxJc9FMfuvcfPw7Z/dRXPFzMDVRM10mlTR2A5TJXF8qpb
Tjktj/y3jBN+JPQ8J/TFKWz16Xj6ivUHmvNOcop/JMiXc/hqoCy7TgjQOt4qVfnp
XOx0Jzd5b+ANeP+f9PaVWHhh6r5QwoFMwK+d7pB+nAtlKvfC5m73AwzLBq1YZj+V
4eM2Alk11SjlVqbohJ9M22+f8UzxeWh0C6F7Ale1fl6Bx3X9p46zOgm5bYil9fGc
ORd1Zr2p0YVbeNWFjPb2GY5mFDRq/6158ifusz574S8oyC2M3XiuVs1oDKD9pzdf
JwInSlLGmYdEPbOzeTu1ltLPNh6HweNZBfb1mUrr8YI6tPBzPNRLSY3yGYlGtHvo
uEFFI45z3yyD1CBHQGMo2r2ixvqhwBB6A6XYwMvr4WkyxOM+6C6BJeZWljGNdbPb
UuF6hnqM5XzU+Ztd9S81IbH8Ui5JtZClCw+Z2Z6HNMdTRc8lYjGdFHx0NJzzAe/e
En1kND4EMnhdHlv9zdP5sJfxAlUh3rayHY1te3+TVSx/vEOIzzmv9Dq366tVh9hw
IG4H9wvTFqZ53oEL2E3CV2zaEEKh5BV5i4xu0HiPRskuZduPP783phiCe4nmxaV3
IySjw8pyiSJU9uwFE8uM6JJrtH93ksvZ7V8HOKH/U1yfXViORRJAPjW5r9kwfoOT
G1zNCKL8NJ4HzlwdZDFNrzqjBAi0Nizcl1FigeVG6VSdu7sFxhMMQPsY9Rpq3mBo
oXJaCOSrBhQ1+LpMElJI2ZyxTCIuzy0q4d5jm7x3J8q8PcqJndOAX6KewQrh2FEc
K8rUvCvCi2N56jf+26MJ70QZVad+nK89s26q6i1pGufNf28avAn+zJjzK2dy7W8g
hdtzdcyaItOiGATQsYYcwwGzioyP8Ja1ttibYji+0zwmZ3AbSevdSsnQOuT1x4+W
fyspH6S77jKkCrdOEUMv73r6DTfGEq+EBYHscgYW0A2nAxV5FksPNq06Z+CkMJPi
7HI5ajwVP/Y2sRBg4BYb1g8+TNT8n/ZPd0Oa8rwXno8U1XsGYkw+IX+GvCN3eTrI
LCeLUsXbolrjWpgcOVVjLITOgr21TbPg7IsKQAD9uHrTDOvHEKqXTuespiy7AmvC
pUR0o9MhEM44oQ5Mf+2Lm+TR0BqO9vcsgSmvSn6ZdFlwFLeePi1mRIchtZZuV4VM
HbpzXrbVuLcNjlaKwm/unz+JI7ayuoho5ewRUgGA8L/VF0k6b8xCfKbiKzpHvVQS
MusTPbqozEwVux2ohJ9MZf2YwXWnvliMJ2b+EltRVvjNWSkC+UR+ARJcdTKJ9UYO
svUFUOD+Igpl/bCD/IuhAtmUDsh7chLfJtcoquErvdM+g4zwSbnmBifHHKipxtIu
qFCG9pxToHjDYhqnJZCfnRhgXqTfFZRiE3aBZl8vqBJ4HzsMJ0mSNL7M+vBszOre
3B3lLeamlbeuCjoUthwVw/CcKq1gPGuxHUzIaP/4mCcYlIwePJngzos/5Im9so0b
jYZUtvZFOppa/Hyk0dk7mspLsvm0XCnxLKRISUKVOGFwlZtplwWTcO6cbiOHdi0b
TWPnjLwEBoIgJ748Aq3TEq93nGe12CadHauEYsgIXvCk1qf/VpN+Mf3+bgBc4SKN
NDTwB9FO1tKnk0n8WCo4jIAoU+IC6hla7uhUjZp+vT1aWdpvIdeWAuFlzaF4gUMU
DaGohygwO939ImpVwU7aNvfOD1l6c0UZ/xiokr3ZzP4UFXGbVA8GslFC44jJigYs
1ZI2vvLK2MADq6W10TvOXwIwfV+1J50UzdV7gSP4uwCjfsBeC0VEc1QyGm1d6WMj
gM+6Jdf7gWQIcfjnLfTkGgJS1acC7S76cedI9F81FiYMtNDQmQvfoW9iuhlo0/n2
NoXG4mKqaDlRvKv+n4Kfb/BSbB8/cNKKjWWd9jUGmuCcgdOHU2Tds5srZu8HVV6K
ADxes/owNkbQjrSlZbYeN2NziiJNHpK9mEcwIUlsmkGNYn7YsCIw9lvBFVP7V217
0eQ/9oyGioobE/+N5GxgIOOxCR1gckOm8WRU9xDLvxXz6HlOE8p427WeBX9Yf0vQ
ivJuHwIt2SaPeoL+1wjNyyLTvVIRBUrOtNMXm3J9msjAopqdF1LDl3glwzWsPHTC
WtD81t+3+lrNcrANa+ymJyPfSOVq6Iy50sCmhugOsFJ2dPw2ne77a6SansEwAlLy
hH1L7mjT2BvpJ8I06+nnAIgiDqFXW6a9edHyfm+MROarWnu9go7NuHHQ/ggQt/yd
kfEQ44AZikCIGKJTmAA8/JMVDE1z9vCfzNvVonLBSnjwb7m06+jt+jdtD815PvmP
7EeYhHMXKFooFwHkssCws56r6ByuqpjQIQ5kS7H24+vs0CCBoXz11zKO/0PhGbVJ
ZUIHoYp2t5egqXCyiF36qaeJaOafFRL/PRaM57x0eUVQSLsd36zoNb7MoO4ZAcf1
WyV5AuJRf5NM3vVx2NkE9ZttOYMxThv+83G1DYFFyqGoa+yPDZeCoTXKnom/P1fH
BPNTWwce/xcgci9U/V780XYw003q91EO5x48h5/Ptas5/19nDC1X3g/tp3oIL/cy
3A/k80fnvciuZv9UiIJnG5SVjIp8lyRERNeD4zpmaJkrj3DwQGEZfGMyU8H5e0SL
CtFg3PoOPpyt0CctgaW6stXWkU0YGzXRze4YLfNxxYyfh12HmMxc79naV441Taac
y74yyf3HdMV0rgYl+Kt33UMfj5bKxVMpETL+s+NmjW+K6rh4B6XoD/pmyU1iT4qN
NBMCXXQRPW20gFKZSQZPyJQyTmf56OKR3jIFVFPEZQvc+FG09TlxQ5LpWwBsQoIj
Y1S4ihCMoPJtGg1TAFX06MtPLo6f2/gxbtd9f51e+NhL3I4K9TWTEmNi3L1XNipW
vVe8wT4/VPY4qVm8FnzoXPcEmfKp/BG/C+//7AqJaXJ3a7QhxB+uYBCVPpV7xxtE
eqQeaWbU4EEqgjat6Sd9BhC+caFymROlHxFZx/niTffNt1J4L4N/l1QOjJQ62c9R
PBTVL96EDNbz92cvbRliEzEyrTAb2yQ5Fw+AcmXT8TuW++Q9xTqk06YBwCw8NeO+
KAZ4qiTmkdCgRrjnmDzkWBa7v1L2zSsAWTPYr2wvumC9i6gK0+m0CftHh29eU5i7
ptF53C1axnXx4oh3U4OrtT8NGA8nW6yPSYIyPxxikk7pSs7Te58CTIHu2xGmn7Zd
hinZNw1JuO2dhdqfVU71edQFx7EavepvYtvqnXqn89+QyJb7hiFKHbHAVqtEykQb
eAoLsMhF58nk6O8pDpZN/qD/gN83O1sxVx/CfWg3n0XVDyK2fTMDNXFeyjzNIIuM
PdWU5+Iqk/6ucPUrowGrzbp20leYQxhs39xeEvUMhAsgNtjn/tk+Nv51AAOFWWWc
RxAEvxZzrTWx5mqAj1mUuqHuMFsZtw7UICSBfsRFkfooLH6eXnK8CzjglkCJV18t
DcLqYvKlVvgy92IQf02Hd5r+snFdy3bKI81B0DfARbjniFOkp4HGGU9ziwDzQFEU
nbyI1G/ni7I2VzYJLam0zoUB8xM4lwEtu8+6umC3dOWCYoJj1JERa4BvRW4JSBgO
SqM2lMMruv/1ASCr1rzyjXeU4JIC8PL8eZEiFRsCT7sSkm+yoz/3h5Muyfk/bWk6
k2zsTHRZpuzxWW9wgXheWor2Pylt4U0/0PN2QcVknbMzkYwZnWrCJWYSxAijERJy
9Q/ipCdv0YWqlVJa5k8pyfp+amQR8hZQAmYDYpzFvh1CUmAw36cG6bCzY7xXNT3a
0NS0NVhwO95AmgvwKIqlO6zH7+MY7MaKPIUdDsoofW+hb0/tDlkNKyWdS3s6GdkY
vgXt+yFfOeGY0q6UateHQ7KWo7l7A1aAHSR2FFjmTovSmserhxbjDa00HhL8f/xH
XjJIAcMom6x5xINCjWZKPbasTQMaTpwPGPtNsEWbRTl2XHASbYdMMvioRHFF2271
KjplUYZLyjtB19CgL4NeishodNiMYXxKuGqJgf2MX7t/PPuSjhl96J5IUfrSkiOi
1sluJwnR9tsczVUjuAef8vwfo/qH0DD66raKvHiAaOO83OydmO9DSSn0n3oG6CgW
yzVH0JFFaonbani7k0ytaH3j5ewyxu8iYNd1ADFvJR4dci+Qpbq0mEos4txcoGiQ
pRHg2GM1p7M0apeT1JArynTsQlSasq8MQVzYQpHV72Eq/S2QGNZUyj9cLa0ClDEQ
kQ4AWqWl5VmJswWChF8X9QMG9e9nP6Z+iB5lKVRtEy/bZi6hjzkaoYf4FdJzvGdM
zyw0J6obCAiS/sI/7Xmo5dNHxmFaddchz6igWhSZ7Q7vnyZ7EYukDvJPx7N+rva/
1TehNWhDwMRi9jnxY9qENbRH7EUzAtUirpEQAiKB3gQo7N9vsvWTDb4fFVM9Q0Fw
2oBo30cZ8Dhlw5KyMGh1SLGlL3Bh2235qE0SsL4YPDSpjCypzdUrGbwfAiM9v0GR
S1vjFBh2xARaPIomk7e2Tt0v3eUqbE1k+tgAm7TI4bPT8o+b4PXo7FR78vW/MOnC
pJ6BN1gYHfSJP9aiMGOeBQjTHmIhH/sx8pQprNs6rOj3hQ+ZFBrZxZSmmJL1sj9j
61oKnrSLVAxweRQzRAVL2WGAExy/visuh/Nh9WeL0vmDtJKrLTrJBZ6qrXLNRlLX
5RyX7ih4Fu50Pmuub+ZaLkXWMEcxuNkRVgmmUPT3ofkkstAlxK4YEpTdS0Yi6ONH
vLBai+jN61dzO4ztc0HbHMTLHyDFBPkF5+qbhxAJ2ZTlcmj0s+u3v8XyElNB9cLv
u982xMKU0GKDklr+47cHYLHlGf1S9k886pzT4zmmrKtlAIJECvQsYU3Fvm91YPQW
tlUkgkLFQlE0IBdni8ZwdABw8iTO2vp3WKDZeP1gog9uF5AuY07mEI6lBCSMXM5B
ojiM1B5mOQbuZtK9vSVUtcsQ7nHvMY7jxnq7NOtW292tivnwqryrKuOYYsDRi6e7
+PkC/FV5Hgm9LVClVWnyIlk9sJspV+dTk7uQuqKPafvdKFk+WaaczerVW/Xd83DR
/ne2FhBGXddURJyNuxuih9ezLBbgDRQ33H/0sVgvVqTn0gDkGqDqHgFRlt2UtWIC
HUJXN8wMq0gAuQBLCZlQkWRUMnsMX2yEAsy/RZQiVtoTWRGsFo9UFME76ZYFdRRg
AUuQY0eVGxsw1KysBAttVq5OdZa2hbN59t9ullR8+S39eLmePckE8tfgtEXSOOz+
064c8mpNOMc024x0FcUYizoZln4/zawxZvsG++Tr8kIUpzXDMdwChJEdbmblM0qm
HUQvAZ5fUuCABm23ZLf0n+VV14e7Gcu7dZ080k2CVz52j03c5LHH617MzmHq1tXc
2+HJhEevH7c1kee3AdpRWg8gBwuEA6mp5YRYCHV9j/FRKeN0G8v2huYMTt2qukx3
4fcZCR6oJa2eDKqFzDp9EuZa6fx+TTrx15FiNj0yjf/sGKEb5EholTPnT8NFPdfq
ki13u+1+Si82zSt7/KgryE7nVlLqfquo+dFtBMMA1xKOalbqleZxBzsdZsuhaXid
nBvsTQx1DR/s7dew4GEXtS2RI1JBq1ec1fwAKYMOzl59bk5WbmkXJ7xhzVmPBAxV
4tAcbnYzuCWGTmb3CJjm2lJAc6g8toXnJYylgspnEmasbRrWb1sigmJ+qtbLJPJl
R8Vh/sx44n6MfxLHogpSkgGE4Db4mVA1sTCufetzm5X8HOn5dN8gAXt8mSrbiBdQ
+vn+zX112T/wi7MmwfJmFXv9kqkgnxhbFlRY1M/wrrR4udscMcVWtW76dTj/U/DA
7byYYj9RQNxEwjIiQ+le4u4l0wZoZG9tEHUXZSdQYnCQzIi6NzmQO5dbl3VYnNF9
siaOQ0JErdFlZHKoAeVzNLG7Nw5Wxc8a75FqD49f/f//tQnvscslx/yIO0FOPysY
WEiqVQxl7UbxGZQkb8U0E8CqFFBoPdcSwE5rYDd56d0SN66xk9sl1cu3536h7U7O
QY/8jJgXiqwm31fWYvtuQ4WA1Da4mJ8pGBoH8EPn+Jfy+pfejihbcyGCiYOIbdzP
z9n0Bu0nHfDqxOJdN9/vUxK6PZHsMQ359D9ccohAufImhH3c71kzjiCFXVBkwkLP
NpIX+P0xpkIjLTfqAuqLcTXnvucZCgefbqB44Xsf8eLEDjgHHjtniMs2hlXw0sx/
O+xVinGzFsBBelzrKTwLoqBJx/Ef5tl2xLhyViV0DDSPS6bJ9RuqwLPn/gqmQ/+D
CgDre5vRu8Iev6vfqtYu7YJinD1gwfWQl+7RGt58ohf/MUVSdrTUJS+WEuNJ58Lt
OgJ0YkvS3XqW4bqNfcbtexxd/hmp5i9XCtIc4uHFJEmQyZBLkSsKda2YAMZ33tIu
gMsN8zUPhkgAm+ARONLK70aecVL3/NmcH4ruh5/Efl2wTiAkAs3ga//tcQo2EofZ
hkKf8QDqEiEXbmIm269qRlKb9/dBFlVZLiU8d4xI0yb2/g8aK5VBDlboDxDn4rs6
kd9oGVtGlpVR/4yGnYrutoNYPTwD6LDVtXQgPbHllCeuxvv3SwPxGfmT0/zRVoJP
GS8ZUya7JX5YBVnhpexI1oZMYUZz6MkseupG4aTB+LZFGf2lF1zau15Gm34SmByZ
Wpq4cPgRMvYRnGrIsr6F66XHjDLjrT6dWHtSA6FY04cCNfuAdwy8v2CM0cqAh5aa
BSI8QFlQU+0Vm6VSek3bFqGETu0nWgXsagzMvpHi+8tLAyB/Ph3r/qt3HTWrMjPa
QtYkEeOOYsEr8/tAJzDWaWIeA5K7ECFEaJJc8Bc8VQOnjFQfF3adF6WTJ/dODtcS
P8zWj0Sg5DHJwvIV7ZtGkDsYcaJ+rW8WwBKgSO4yeYk6UoXW9TPT+9WOhumqedCp
KZZcjQ2RjUxm0up2lvTNhIqJ946/D6djCePbv1GA1ZGQDMKBU+F8yzdj9fAcygse
RkcHReFvpfbqNuAlCQpSKAo9/vT4EQ2pM/q9VnaZjxtwmftD+23q0gepT1P8hFRX
HvFGy+V7wqky0qzm7Ix7h9fO2QuvrSuCguyNR1/XjLG/T6L2yMuJTumqsa9tcPP5
U4tpzGaL3mKG5wwLsGiWQkMmkiDHwWNnxVWaTE7pw5jFDkFem/dVlesUmeyVjsyO
2TNPMoDYXeAqubr72yCT9LwKfptV5juFeevrBzL0PXDEE6DbNKLCPQNq+iIf30sl
cfQIhQNrudZJlyqWLMaJAys7B3cZkDZovbh4WpPpkYprDnaQWne8WA/vtTkA+6bG
I+NgX0gxMpJkukYunbvRRYsFTXc3ECvHtBf3jlGoF2NHq/A0zWlMJSjVU12JG4bQ
i7KDj+QeqSgj7uG2nkcy42ong8KuFcol1yBmnNcFJY89wjRj8hWMlHKuUQVzv+3A
R2ilTUvxNtaxUkoNNmFv/CXU5D0REaCoDkvv5k89aiDIS9xNbv1hLgzYNBttXXZE
lNdurwyGs3Er5oBw1pj83QdJZYOZ+JRYWcR2ih7fU6r7IumzUba5I8xt9CABWBAR
cO1sLp3Brw9Ot2Y4T55YDVrGYdW2nv4WaHQGYRqDRJrwbjjIh1QCGQgz9+pKToVh
Hlm0GEn0hCN6cjGqkKod/zGDDUXFYq2q84XVulaM3TYINxQF6ObworO9oQz/erl9
ZXsDW0CzHOlUAvHM8PM+6LnGjqJP5R3r5Chv57CySb8wMqahR+O+44NjuUmv10Nq
W6VGu9hy8KfQORBS4w3NdKDH7z8aVOD8EVX9gIThfa20z/9vRe1Km6w/vGWH3AXH
U/XYx2k/WXdLMvYo+cSbIasJOL/iR2ZffYAn7mYVL8I0WjwJoVs0ojkpOHKdr10I
+dT0KGGxrjtjglYQrmz6vc+QBzBkmNoPO7WoQdCdtIl5RCa6Szv6khhJLkBtiXcv
8YpkXG/2D4zy8SiKNMOlKqGgly3udgvxaI3cLuRllncSusH0H7W8royA0GlyAYWA
mm59FhRe8PRVdQbTRotkDTcdrYeU73MOvL5PbJYGE3H8HsqEZPHO6X9o5bDnkIIa
UKDzgHHq71r2N5GZjHC+AorSUjtpb0mpmsNrYFK5iil1IryiCNQffEFoEVWL0nHs
7yDdsns4bGwbXHosq5uwIRpWqa+d1t5sJHWwhx4FAzrYH5OPQgCaYke8iO+3ITXG
3+KKTe/wWxSEX+H7O3QSODuuW16XUAmNMAIvMpapPGGRz5GN2YggpNNcamTntpmn
Ct+pLSdo8YNyDncVdMtjZsCH4W+ThdNjNLfILXWW6H11uDsv/1jNvfzj36of3djy
LYQ6wmljyqgVdhtveqU2rMepeIVM9mxTjWIbsWyV3KHZaIDs8oarNHxs5brnRmbi
DEBk5Bz4RA/kcm6SSN94Uy2pFBlYmd8Xy4Wqeibhf9f/6GHzeuInXwG0pyJXM7Rc
3jZPSsCdz6TdoLlOvEHhvT2YPXRdLFAVLZDvwsF33AVs1ZJ2DAnHw1b0mS/nyces
RUwsD1obYTjiw5eFyHQaFzcYFSHFWd5DSoopeCD8wZnR5sYk7q4Wb7j6ZllrRPG3
MDOZ2S8RJSSKCMinDzckgaX0j5lu42U5eOmtaUCmVQqO+f7DPfEmW+4uXFKgzYSk
9UZ2qLkoZCNaT/OhUkKs1fWg5j9WLn5skgu2DoG9O39EYpV91VNhsuG7P6gFvXzo
4ZZHxC8Dk2G+l0xYZOhI0KVGaAGlbR13wyX9BiQeLoqIP4QJEcFkdJ0cwsNVrUBC
52sNIkuQX8KwMJKoia9JfC5KWOLNFVPQGmQZH+uYFfmWb9SCiKW+ITdz6Ulgiew5
1KKZ2Jo+w8U0MI1OdS2EJbuwkXZI5TIQJvmnpceqHYmZn4TvfylhvzV/J6YUDU/j
aWJUSsZefjQG0d09WtTQwziwGoJcw0SyFCLt5UTrB9HL4OHMQrstdWLi+9/4Kj/R
213BgzvzCaX8MgVHgZnmXZ07YyDKQwwzZ/nd5v6VwJRpflDjvD8J41m06QEJWA5h
P64uANQg2m+g0dPow+eNFs3UvMKcT3FPw3SEwhjQ5lVdLH2UWgYNB67B44pu20qt
8lwAkwLrShCGCXBlgpS6WPrv8qYW/erLGr7d1AS/K/vmRaiWV292VhJodn6Aj3D3
ImVkeIzkf7YgJjyD5ROAq4og9AKY8gNiXa3+N41yGgljvDq/L+d64iPc4oOynOBQ
tU5uJLe74KtXKU9GbkJCahQCzlQlf5leY3EdBrLmdhQeTjuTjXxiTuh6ANPCC6zp
xoEmLiUYhFbe+w54KjGf54noMO2uXIWuK75KD2QczT8XiThN0Repafd0yhKXfUZk
bShjIo+83ies4+tZeoPdZS1g4yA3LV6+z0rolFy5fuv/yioh6WorOolqXNvS9MZ7
IvngGNLMbjpNvASyol2f81Y3zgY/eBY4leXVgEgAqBPebmudQM4Dg7k9t39gyOdF
0BUVpHjiivUkFEz+tB8Mome4zyaas2P77bMVNqLjniNv2tAWK81sbyCLCvMtDG4e
Vw9tzB/ZVoLlhS35SNxqYC2fDmZldKiCp6v7lQ0iE55GWJyqhkVCxy3HbTuUZyNO
gd5HdO6MsAkGx7iYfCzH8EklVQ4GYnCH9tq5uUhcGDTuK0TWiyRRweMRILhnAFOc
mk0JUejHpeYddfEW2OV3S8wBLJSeEqXeJbX6fraVQLn4eUcVQ/gOKLlqXsUJmXob
rl7ocoIY6mPcD2cRx/3VzTK37GF4eD8mT9svLD4cOUl251dl3jUYCGNgt+SKltsi
X2BdydE39VjYYMQJ/qsRmeqkAl++gy9/yYFJnlwPEwPOWlc1pWw8u4HJgo3XBF1+
ZktsRRp+jsoNBhBMoymZWAvGk0ZrYk0aElVH3TLr3L05FM6JS5682Adh4IWcrTsC
vNtxQPe2mxR5rl5arqsGQHIYuMbDKTgMOJW88V1JyC3DftLXJtej5GNVhzzvqJqp
lnVoQW/7GiTicJwiZ6ApmkvS38/f65C8n/i2W4do3fVovPb7eBZsm41vBGRg1IU7
2FqLQoXBu+KyJrtH3tx2zTfgCzZyjenZw/0GTr5AhaupNCupMy9WrCWrkSJnk2DO
S3j9C8RSOroofCbly7mT4ra48ZxjHzUK1RdloPLaD3Vo/UAMZdTx2aqTzQ//Z90i
rtYDr8PsUUTH+3ykV6k81aOgceOjywA+CS4zhwSHIQcKVLfBzGLNvZMQGNc0osUx
JYlybl3Jr41KUJADf7EUAbAaMT1MVosIR/Gq24NlwEp3fHqWYF0A5IuK5f7cgc+n
hWN12OIrb2g+oFsovSj4uQPJQFAaUXQes7LCD49M420zYAExlzd5Lphy3FnE9IOM
ptT37s8YDCWaZGVsuI2Da9FRHKZUt3B/fhP2YYbXwSxeQo1Wdc1iC410a1B3KF6a
g8YycM3vWPe+Wj56tEnN+C9Wmtd9lRbrVhPUw55ggK1COOHcS+bLG2Kuy2vDn8WX
9eTxFnnUfCKfYAUDdwyuKjwOPNY4qsGIX80Bjy5VDJpDgP5bbS8qQiNjkcvSv4sc
b0+kzAoUag2/LE2CYj/du/EU/JDjWC9D8+drkSavcaP47Z6ZsWsfAMLmk7BGPdYl
CaYGVSIQnv7qV6p2S47MbFgU80ahQnr8KdSTM7xtD1EK30nJ2H/o3UtLn/JCwlYK
FeEU5tiKLkWBk0iJHW0jq0IWp9mhayPsYDm+RtX/FBahLU06yrpKl8qSc0tNzBU1
P8iy/u4FA0gtctcd8RHKjdwqZG57uZCoHq8DFLV051h7SsGPGkZoLJwGE/W9X1Px
nNNyAzYuQ8jt/nRfR9F2NydRq/DIUf3/sy8kiUcmbXJHHoOUK5etxbuuPa2JzJm1
WmnEIBruflZ8mAJrBj8lyAGUNwtb8vOSbXxp8nI/qdXAniS70FCXYSTPRGZ4VRJk
SMLWw23uqxZr28MLL2/o8k6qKRjfcTLycumm88zzPdF4Zh6z/JqMopG6COv9D0RY
Hw+du4G+boB+q75KLmbEmKBG7Ci0yIlT6qxyGcOwaXsnlpSxYhIypKZrq3m1Aitu
v4RLEtI9jcR2o0GS3zyJKwprkbpyuNok59KeJTSwn/eZTxbCiKqpY1RuHo6Wwk2G
T6qmptRkOdqhDSCtJ2EYPRYVYvi2d5HAoDs9YB9AoB/iDWilvF0GyI6cT+3jeqvJ
me72cdJF3KP2r+ydt6lerkEMW+N3kPQ1isFnb5P2QnJ/VrDBJ6qLMMmziVhr9241
GFprYeC7gmPkD3jonzNAulCC0S0JMZ/HRj3Q0mv+bYKrSll41r6osIgP8gfUA6fh
hpM68W4D5TU3ga8/mnrs7g038Q3aCQw4LG20LeWU9ZLCP6jh8UPKCpKKo21617y7
gHcJfsh1JytOOl6NCGP+4T/26U7E8oY+U7g+J61CDB9yv/NryfPliY8vSQVSYASK
IKbqlWuNsu+41JrTeFQ2WpS60A5WVE1WsxnFL4NbccNDQB9cQci+2bSSLZOBhxxa
okB0hkTzM5JQWTptHV3KqfF4KPbeKW4lHveIYWKl3gA91Jm0fXgPbShjd25DGHfu
ntQz1h75h1+duFvd+nhMQB3H8MXcMRsQfsC7Y1fG3A045LTsVvzC0ijJcOLkDYWJ
++XNTm4+au/cKjfCpDs/qWuqPcI8ZGs6YysQtEgsV9VBP3sbVHw74MTGsBK2JobT
6xoyulj9k1TpDFqddjYXI5Ok0hd9oQZB6BXX7SFSd6V4IFDJm28eV8KEGda+fQbN
Ff2LPMMfO8sFOAxknz+YX3eMH5UzEijRokQU05nnb/8ocItNvj8CIPadUXWWjjb6
9QfxH8sq1/MDIxaUNK4VMo4FAod+iumEWBrdcjYYx4FPy7gJmG6YXNlyjLK0Urz0
7XpsqHjLz1gOZczSPpeyPRtuYV9qnDN65g6sZXTTTfLO4JzAuUziKNBoha8xz7AD
A05Ojh+oFZVV+xcAJzW7kKQ6a1LTBjlVTK9SJiE3J0d1J/alTXLr0DJUrdqYrf5y
adNhWOE+UqGhjv0iKGWCdnTsNNlgOBEuQcw0ZnoV/bbP8StspnzqGJreVkLCnlJD
tEEAe5HDUutQu00CgepJ6EECWCuvk8hN/sDdm4Xga57ZDzAeJmOwmtoERn24LaiP
8jfyo5eaTRci3M0SDcVw/uEUSuXq2HdCbhFXqovTiCxDi90gb0DqvN3F/IaXMT72
n2OPJZjBBvhLEuMbc5gE2c66jwg/7/l0Vl3aqRLe2oa1ywuy9c+uAmr9JPEGsx+L
Bib06cMMAez8lrsm+YS/jzb/MAAyRUoLEQR0ao0P9yFVvzcc/AmW/mMmciJKmnUS
DUbZU9ZEET5UkxsNt9hCVgRS2+qWm49D4LxUjjqz0DChKVa2AgL+GLZk7+NtbrP/
nvZA5xBjRkqx7FY1OVc+WTEzCxDT2lzUODIVSDwp7tg1rGpBvEdLK0/9ziCLpDQ9
ix+/y3eHu8s/P0M6/ktB/UBh4rKtaBXc2FN4bZTnd/H+fzJTOsPERVWuflM7t/43
XqgZENuANR9IopXLEVfv7PhfwIumYLes4Jr4mCYlTGn3M4YY/epFz1mVc7tSkFwl
31WIj4xWKnhdHYNOw3TFA7IXt4VSBcdHP7GvJBYRJX9RkqqFrO3Fc3ZppAQQAzro
cGbDNX39HCwO61YLbXHflZbiaQuknir26Ted7INROB9cxVhlSUTktwWLYHHyoqr3
lrs1Kv7hc09wwFsCm6hAZSvcCOUZ0m9JDbveDlImDrv40RhJU/NOw5k5U1Uc5DPq
+3cnPO16y9ltzTENm2D3a2IZ+UpNwYUqQ9VSFGk5qA4oiUBTcnNxzDDqSRJ89BzH
Z9CVNW+yJfgA2rtWbehUBM3jGn65xu0xQ41JkL0dBrd6KQ3DIHpvPXKABYJ/XpRX
Vax3jmg48gsDbrbbN8LqUBCGzSNYsHvSfYAJqpZpKiQ4XOmqhcO0W1E3jYgBZXGV
FxR4k1f/Rb4KScMN98xXsOm0o2Eb6apCaQpXCRonaQv3Y5Gi7Hda8k+/5toYjJYr
lGxoaTZoPm34/H/jCjwWzoh+Z18M9VuUZfYLunYSJbA8Tr5U3vLN4iryoeBT1lK9
Fb59WD1VMD8rEyw6CTj7eB0/hsJjHpgKYTJZmK31maIvymwdodmtl45Dv2lq8vaQ
6QLexQlL69M+JRJzrljsOyMNVFQxVVB2FErFcqC6yNKRx44ejVIaIs7a11GEJ7Ol
CPsqpHI+m1X0HB9tj4iC/QJDQEr+gyii/LRfIFr/6CtHl6MBlrTpLqeyE2b7VDTp
WED9/XyAB1UjGXeZm64nc6IwPkBzJGmETA/4x1HYdE4OjHkJtAs9Gp6gFgXMIi55
fWxIVHiAieWPrYqUg8crK65LLPRJ6zkvJ3qvUzpM47TEqzg5sFe+UmAtF+DBnQeC
6i7ZuLiS1z8OIjuVpKUYV2bXhFNyl0OYXq2kRbrh2UZiTw2m+DdF/1EofksdMxI2
XqPko86xbRxbs2upjoYNVZIxYlH2wDqhibXG+NllOWWFvKCTd+civBaKoAEZdUm2
Ytyv5wAK4IPBK60dJP/eq5fcOPrnobqWzLJQ71JrwH6KNegfCDbzlnkqCL+3BVAA
90XihbajaZEwlnz0Fe+UlEQnsawTmOZ44fyLAwCzRTIgTyX+W0mlkDqh/FGaPfh+
47me0W3S0DSZMVKg3CWexG7dUFvRTrP+1+QHlGzoaPUsf8acNWFrSGcE8LQios5q
V4W6VQrU+fiHN6siJFPhDNB1q71dtwKkWf6GSoeMUGXPf0U28Pd9qH/SE6XBTtyF
AbInYA6vcQmFMDNMyr/97KCu5PQx2iJe4oYU7Y+PDbyq0U04R2vy+xMVwrr7sVup
o/lNdvlRHHnWpBU2mZZKu5eYsEvDsVxAhAkuvWj1QpKVsT0fRK0MrMJjREv5zMYV
asFRAHL5IIvJciY/5UQmZHKcOfrgZW2F2+KD4tW0vjVlk+kixK50elXIUr0vx/mx
Pdcsmv54EP2wAa60Gfa9f74NA7qgqURNKt2VPxXVcwOYkxCvsOJKvPhjdL1lCVge
gYBbQEQC9YiKK7PyFYB7FFetmvtGlGe4ULJ53JUWJEUetEnULhz64CvWMmipNhaZ
6uu4gUdfOs9+Bsj0SXWOwiC2NB704AVk1Wtx/9c2GEqvIQN09RwpWKrF/RIxoFaP
71UjlzNuaBm0bZGNHb3Gu+gW32TdMz66IeSIrVXKfSxgJYVYSl+otftFeYSDT8DW
aSqNs7BDIcOVKpZuD5Me9WkXFe8XKQl7+sczRCmNhKMkRooJ/MEwEZH9Gcl3htnw
HGiNXIO/Hfnaj2W+J9CpdLE8g3wvsFrrKtQw8EyBHhTxFECbI/0pdPo1wcRlDk22
2c4PBGqr6LnHYCO61ILE+9SnY5MFHmhGYO7e0w3PUkBrpq76SDrRB6LjT1g3VuiQ
Nmc9LtCyVZ6GgHZigl1JGgK0VNmvjhB712lwaplDhJlYLRfoY+Fl4eb16zrQRQt2
kcYF9As9+5P/LUyY91IKrWAyxdevgFlmDAd7h/1Hu9giqKbNvgN+00Mrb3GTktVC
UM9abH/b9RkB0xmutghtkfxU927jyV8Z8PRxRVA8hGitLDXm1k+Ko/GFJdtaQiPJ
EMYb3JzqmFt9hzIX+ye8Eyti3KCJQK69MQmBlsQSpeUQS6iWDr2qA5S1U3NLDId8
snE9l5kGv7EveKWkNgT1Zo7YqVVmHdJCbHJ8VAi1hcJrsYu2nMSTg0COT9RNLlJn
yL4YucHfJ/K10+fJ7qJrJwT4UkO6SeXas1BXrLyUa3/qW1j53AjGU/G7sKq38Spb
aQ7xv8WOWUULDi1/0yBM0EUxmdMqMVX5els4M6VYdX7jPlav6Nh/8AY1+aN0dcZw
ko0pF7olwrz+pfoY5Uw16jonr6DM/odXeXbWPK8r/FFBgGFKwtKy9/xjeY13BFIo
falTiz3UNo67mQJkFehlGGWmiCzoLdlWoAAeQ+DQQV0/RyGx08zEF6yqNs/XZo9h
TxEAiimaM0m5nzlIjD4hc5lqpZP1Dd2KHT7TgxIRxxvWksUd3b7GIj87p1h+ahcn
jT9MJIK+0vxvETjTVaWE3xb/s8SIcTFJv4Op+p4e0lANh7JAv+G+vwk8JrECrGk8
Dsn8xH1yUV/DPMnf74RzE4L2z/O4bWmjVTexT0HyiEfKUPRwde7w2dxEU26MZM3L
9fjoQ0SyxeJVTEDBEsFgSK1vtyxxeth3aWhcpny6ffKNzAImJgZDG5Pp+kf5LsO7
0lqz1H7WMqEd5Q8e/CPKVawJHz8LA4wHsLEGPJin3rgYz63HFvggWLd2/5usBZl7
ilA1ezF/X4RD9trCwfR+JUu9KlyZtSBKvI2CiOsMXRDoFhOCGnnLcK5SvRD4BXJl
A8stBnJx6n8gP0fIkNP783C9fnYhMtJIKE+BKhxboVN9UzcIuDsDY9lzD3MjTqeR
lLARYOJCcsd5Kx6s1dvmeu7+s6XnuxS7lh1z5sL5j3mRX4HieN6+Jl47npPXMdYf
pqOyucJmNJb8ZLQ+lsUSk/dzCTQCvj3MMdpiq7kd1cBmGny6Y5iKezILe5SXaeX6
1/K4TzpZrLZpvPx62LC1lMffG149UNsPuZi5FeeVM2KXEf+A3wqG3c6gqWbP5I5E
bnS/eivqMzSq2GWVq0tJKFvKekaX+urCwQUea2bhh9cmLYKVMmWAX8MYjgw+k9Dt
xw+5BFpmvWFUETTY3JLGIoV0PEcmjkuT7GRcm1K/sTYsOyIo/Zzr/IHDjJ59HJ5T
iv/qCsZ3+P3z3bYigaVIfygHzhZyVouzJ/HU2u0ozRCpd9frWwUEcgBf2w20iw80
gnaO2UDR29iz3/Us9V/gKTGVuo0rgcoRk8Z9m9s/nGQy82PG5WqT44uqWHr/uhSs
WGk4O2cYsh3ZTE8VMzni93jx4lnTW1FF3tjzas7P/PlfjWY4SChUWXhnkA5S+6Wk
4skqvDDy0nuXNhR8QV07qZBxvIVAk4tJw7BpnMu9DadWbmfw7rMyP7fMpuU3f7Nc
ChA9qLOTUFvdlAZPkzNpW2iYqCBNN+saFD+dv4c4JiuM6YkCVpGNvjTXHQt61Ksm
b1B+ZQaiQP7KKvAre/kCsaXQclckfYMm6c/dv7vnXOB9vr2GKKaJSqPX83HadBCl
GX9rPgkfvyambVZgmFakgJEvx7mjG2JsAetj52VoAr3jtj4BIPD6l+LnqWoOpXSD
z9Ra3qVloVM4c1oVbue4/iDDetc4+Nd95a+GhLTD48vZEeRwTkysD+kDFsCFbyPc
VQP93ezNs/oTfKbQ+dfrZIeJ8fKCMRdmEpSOXiXlRgD/jWou+TChXzB0Lodv9DVP
qMGg+W8OUk5EaePTBf8RkCifjEtkiWI9C/dP+EZZhoPJ53g5QpNMWCBMzOG7zpHB
pX+3HP1ooyVQelSdtywxwm2uL6NURRldIAJx9a3VFcrWJX7HWd43Xi2Y7CznT2/g
5wjNkJZcryH9YuwmVyrW5Fwr4gesKm+kTwDGPPEaoZlC92wz3+kKGIp09xv8l0XY
ejbqMC6y4v1IamJRmBKQRSb9C0jkQReYYZiglQQndMFcIM/YetlL1jqzvXLYEgwB
kGAn4j3CC3pdmupcFZ9LS1+3iFExbppfZnk7OeMn6GxTXwawlqfc8EPcdyrlMgxG
Ev5x2KHZMXwwGp2NCqddCuAjmLabFCCHxmwV5WWvwoqcVbxHxID7MfpMCinZaT5L
uodchQFLJgrXTBj5C7ccpa5shZmrqAf/oMl9nws21oReabDJ6lEgdEIMQRzvV15+
7Avwo5IkkFdyvaYZlKNSok/rHd26UWCP5vUEdSb4H6afNwArg/RadXBybA1qr3/O
z1iUxUL1A5/wBbPwf2bhtE8IEQ2zssgfL11QESsD+wWog81cXLg/NiLLsQtBtAn6
dJvljnQqgNKdBcAjIaYgkOvXTToq/fcyN/5SkVITSae4P+iET7n9ePMylQqE/klB
d9mtiV2w1W5YbqcCwdr3MJ2uSz/i7baTMHS2r3RltaNSv8DpESiIHTV2vsQVZ8Qo
recXVMN4vDPnWY+Fgi/njrWh/PzcVjBK3fQPACs7vpBPNQ51BZyCSw8uwMcIyTfk
AhOBuOU0iXbzwiaVEHqOU0qmAd0GdGIJ9DBoIwXo0UByowEV4wDLkJyjjuHjDuet
PI53UFxa2N19Scw21kfBKCgDxfWI9zT+o9ABNokfazdJUG/8RmlHCM/boAb6guBf
lEzTFp0sNcL0GwjzGjPLsGYT/K4tlaJjtV331SaKpoMUqCaY5n3QVJsrwrVfTY/C
brNS4sr/0vMMj/LzWgIckhVaeHkFw/wvV3CVxqpMq/XqpvpKODRhOz+4ShpqZPk9
pEcUxW+v1eev/g+7ojhAvaT2NTHNDMFeJLjzeUJX70yJa8lCA2FihLtSJFo/KODG
jfuEubjDljX5roUbxFtPg587RhK9LJcOwXxNEgwwkohVxGrhqj1kiYuNJn7e6sRP
UhlY5I9kfd1yDxRNyg0MH7RUWgdT2AJEewDb+45jVTmXWBWSK30bdq6aqvQBdutj
As/Ayn2L5xmki6CjJ475kCyDTRriIN33BcB/XHtNTvvqW/Pukt2gxq4Vp/EO+McO
T8oIhPj1ksTOOmj8fLxLsfW4z0vjFUwUazFKWC6yn0YguGHd5JdR1Nz4iAomxgxV
9NvEDPRxCpC2/9iwb8QKRiiRZhlhafcdoL2emQ/yC+wTuTKfT6Y7p/1bhbkEX8Hc
3c7nZcy8+/2SlbJ6m+BHoBbL4zhtQIIK7LmuZ+0YiUhFxAGmu+N1jPgWxXhLA2D8
ubtokUGk2TbB/zEh2luMT7qkaFOcDXSH6kDts1Ny2ZgHJIoFhPYxa6yvr9CcCEXj
Wnyem1Re6M4HIiFY9MC62ygtXFxOn79JGbtBE4Q18RRUYfp+BIcA/ZbgHu4BbEAx
MWtOOBv1EG9G1CYPteQykxKXsFSCxiC/fzwZs3FJkRiIkktu5rIXh5tZWDwL0Lbu
q1xL3TgKnlHjoetpvxB3VUu8Hde9ku96b9mDiH/NcvlxBxiAMWUh1tX9mVkDCvyy
0LClz5QEifdds4lQ6jfwHhpTlzwHDzW8Q5NleFEYxs9/fHP7PvcSwUrnncWP3tgH
yUSPd0+dx+7gG+ITbB7cTJkJYvKtFVMP4ITtjL0WB5iPsg57CDyVWU8A1q3nTWxT
ry6Jsb8GDQnKbv/i9QRZBHVtg831+XIqaYXLa9Vw732bKJ4P/J3mBIc3BLSj+yq3
x3VXISdDatFIsihpTyMMY8ebzOMWLaVqelOLrLBE8q4MxOaHb3RQSPJk0CCL4iro
Hg5LqrFusOv/NR6WyKSBbXffutEiuHDhM7GXHXImB764FeiedFXQMpNT5JN+6rcM
LtAc2kVvMU5WhnhY9Ht/PefZxB8fkuO1R0PFL47lvFvJf3KXvRQ2VL3xrRmxywWx
zMdI1231sTkGG6QnHPAIn4Fu1P62J1nJhE+FwknfUI/HEqMikcKCDl2dnkK6lXVu
/tOTcDQ0nV60mYS4YyQ2XSX0tSiJJWB4vTcQAqcm2RjpXU+4zH3uAQhTN4GZ4D/A
hw4Q/wqe/u6Gm7g+zajFaS9RKTrzwtpuX+lF0/KHHFWKWlhj1QBT5ZEc3daWuHtu
8dZiv0XbBtcFz6196NWIiP6pR+dp2vLG12IA3adV2za4nclGoQOyGLrI7LwMxvr6
oXfeG3FelLjNVXtfjQPkcC5ChaSoFGx38oGtd5SsMwPR2BayPJCVMqxbvchdpd9B
37JXqANODaBQHGu7El37z78VKczEZD+stw21P03kKDijnI+QodoSkBicJcXTil2a
/FpVuTDMSECeKHL6lUYZ6QQmhfvq0rVXr+pfHg8LZ53UDoLWJcH/ZptjPm0AgicV
hPQFP7FDgbqpipZY2P21LjImGTFZULYULRZYB9dD6oNRoIg7IuKWJ2rE3Vq5Y+Np
bBWKCA36x5TTqs0VwuYIvOBywTBCYk/rie2F25Ac4A4SakAj8vWuuaoxUgH/Mm9K
7uUqDRRoFk/wDJ31kZCTsaQhvEPMbc8YDuCFIhWTmoDd1FXFPXNHezU/tU81rrDa
H+8XJu2X4VUmikobcfsgD+JmnfQW6O1G6MvkTUdkDL4TJgI3BkF3OMEfuAeFMGUz
tIvgp8ebzrhUbvh/MULN0LNyOKkAOgN77TM516LPhI/UJoI6t7ZphnzuqlKtJ6et
L0nmpR7pj318DGYuhHs+zLR3DhGOVIo9L8m4MJuSQG2Igr1mYQgYL5karNqQOakA
5WYJfgUiHneA5hFzD6fkllR/mWIhcmscsALzL+8HB39y0MmzH94dpnk7mq5jb55f
hy2Y6+p6b431UQawOaPBuxCfi1HrSAf5XNu0EjhFXvo0/oaABp4VBb+jd2nXLcNc
bDftzxErfdR2BNAympZ9lKKpqYU18Rro6y+pOqimnICxU6jByEJufhMYloc2vxEN
2u7GPz7d1QbEj0JBZjLywQdJ+AsChKAdseGh9DnA1FMQ5lTzWyF/dW66p+ZUp4oO
wZrZCmh+qe09i4xCPaWF/A1WRUkaXIIIGZUf0ePuWp7DF8fBogTKQVZzWRrsaosu
Q8ST8qexEEpgflf+G/SeQH+K0qVuhSBv3MvTvdOx+ISJTdiulH50S6mGm69CJH9s
Zwy1cUJ/C0RfZjdPyBOEXoYBCpiL3a53kxor2RfavJNV18Yqp+emLUBDSDZtt9FJ
eniS9GIuf+bNj81F3Wva0tbsWM1GwCiFg6qghUTm2COCcbntd/wYg4WMSvqLgkXc
3+F++c0fPX8ihj4rk2YX3c2ZLOuZUTFjRGYDtHlab+k+0bQsCP3lYSJKS3pdJJ/M
Tvs+F2JkCnf/I+V5aTuAXyXoHDe3UjcylrnKJBQLhfj3jC+4vkoLcokXq/Os1r5M
CCboSSBUiMemfWd1Z6gPK9DGHxpCY7qvnsC2Xgs8rfAQCO/iW/tQHt4ApstonZtc
E9J/MRkPRYBZF55LV8KyO1Zhnh3OkxOw3wHtXTJqJwbXdCIh7Zt2FixFbHIDbvox
O+XP5t9bmbDroswF1NkwUogWb+hhK0L8RdKP0x/DXohwr/wbfsrDPciwXRoaec+d
txq/t1HWYVS0/rSAV3yXR5fsCGkWNUxayzwWG5I745OhDBwoSC/63Ic3DlkCtbn2
xmEKzmdTnMcHI+HYWRA+d2JwuNAZUzVUChaAdL2MAq6Z60UAqWNrOFOm3g8QnTeR
Jsb92FwMGXcBVLpww08zi4BI2gGXn/zhzr7+mbdKC1LnPp+XBdwR1DpGhIAQvTSn
NavwQ9mCfjW2I2UPx2dPgGokHeNVq5QLcMMW13PSLUhvNKv0rHEMfNtMRrp/uDCl
nUpzIjm65kyLpPnxyE7dOk5buHnHIAO5cfJF4xgV3v+4lFu/2mf7Fnd6tDyFCHII
/iyULPGsIphEoedIZdIeRbgzQEZbQFrOcwBhClDVykKyriBEep4iFWiIllNQPgfE
4p5RgEcJRVWlNgjqWe5MuDL3hpvbILN2LLD5AZOUhe/fYR+F9M1vl9VLqhg1wz03
/CBZcFrz2y6RLLxMp288M4EmE+dl3j96OC8cwJ6ldywQdu6BT96ZGUzbfmRj3N9D
gBNPxLBiFBhcdRt0UpYKmL+UJNXBwdcGkp2A1UxOhmi5Z4qjPc7ExS+dGbarFeyU
aptoigFRo9tF0I7SDgQcwzTF/yCfa+c4j0p8BRSG1H4YzkWUNRUWHgDJq9vRNjSX
4RohlVgfphXEmTJ2XlVEnxocZ/SFyu1OIOPvyoGwZXnRMOIs05ma2aVeYtcPFuaS
2PAb4s9YaiU30dZJfYVpCc1vgPPwNsqFatRhP9/D6vXtWkRYJaE2iSSBlD9dW/hU
sivdiBC3EPgggs44aiRDs8qXIAoeiRQJVo6ZQv2l1zenpkkg6kbGLtdobPaUoKM6
FMpPHh1fB+wbKgoz97glUuD6Xhc1iWp86Yz9T8EmqXKb7zTQG71Nm4E/S3i2lTuh
VCvEd3wDlF1A/aK9GriXiswsvNeLULcHXpXvtZ2Bz3XeQIieJKcGu82+pMIrgMh5
7In01b1g09Ydj5MpoX1qB3A30gPpVLhEBbNOxWsUEmTAxQba8uB293iPJuGk2EBk
Q2TllGaE/gi81FewcwcvgkZtfvc49hCqvnyLMk9ae6R76zAB0wbNWUIoueZ5HN4y
cLKoONMASMOl5TSB6Be1GGFV39qOW/37vagXPIUIPwGBOJs3RnStwmHZcojccxNM
chQDvyE2jr+xv1MMUjTr1DdLJuy/DnNbsa8sQt9NoZlbvfMATMZquOi+2zrbgicA
xsLH7ADgPBSTNJhpoHhdzz1wBdiC8hwiK0R5KWcAonJMaRuVJyGwB4uz8FppQ25V
NaAFMJAJ21S/UTmc09vOuOdChCGeftmGC1BBrPoPlyXSyabicqM6HPl90m8gWYnH
gPV0rGtuTZnv7pjf7q5JYjXFOZxEDffyRSzsJTxW1RjOJ0K6wDPqQ9QbaV0MAw5Y
c6e+1WCvmTFb2KOJY56w5dQxgD7mgv/fXLNhg0RqfYbExnTrLCI3mrTRqQ9d8i3r
7XR2UP18xfpd85+SrCMr2bTFByE6U8njDlWY803/bFntCUc+Psihh9KQgSbd8F0C
LU5WPkr9hW97JA5MeLjYtbyxCnQYzm+ym49xys9YZw5ktWE+hbmIUPoQ/aW5xAgx
/Wc2QfGsw6DjfbdqTVDMWPtk145fTyO7+BsTT0aC0/nv0RQjZTSh4AvliJ45wiE7
aEakOOQAGfs4M0ttQfUA2O+djZBpUXN1fvc8mQs3d++1Eo9a6fJLCK1zpfiH0zgb
4azio80NbKjkc2q0fs0DUmCJHzG6Wv6XZHDAJnIH3qYWkwy/h67fTwgbzYq4AVWR
T9KbQWRsHZMaJY+6tGvz79AoDZAacjm7eA6nVcjv8qnMwu5PN30VHVnE9lN4s/S/
88Kj6X6yGwSa4YGqAdoDHrtSJkeUWOENvDhKq6cbX/4T8IywXa4pQQ9yJ4lpqUZI
eUZaQjGHbP5IPfHLMssAfoFvqyJP65w0BRY1Is/8SJun1uggRYg9atAr3VIsJu15
qOJfqiypigG+0aD6MM6FsG+FvCFrdHtpeon1dARnz7LR+ClHIfJdEe/bHj86keTq
UJzK90BtkmWaeydbYKToPlt/vLqrpS2i0ex/osPu1hdnestZNNtLUt+lcv36eAUI
hYYHJNZ5R0E6kVe2m49BZ3nVN9brvuPP1WB1McumF2jHaIHa60Mhvpo8s4iDz/95
7P3cfAVVKBo2bgh71qAsZTXaSNPsbNFYwRjGxkK4ky66YkVkhiRo4EBJvvwgFjzS
0ZqJXWabTZDHgehav+BYctAMszbKhDOYve2SR+yADn3MQsYQCvRvg5qUffVUv2uT
1FsQZxrXR74C+brO9NYS7IVOzKIMJTfHPJoUXu0Ar4kfpbMRETsQZL2aRkgPANr/
rTGycqHWWYNQsa/RP23HfuYGAFvzPYPnZ8+aHzTAnj8rbRR2aiNaOLVxVwV11uag
FHy9PX2lTPYC6m/mwKq5e5jkUajEkW/BGrOilvz/NigcM5r+YcK4lP9o9/lW2hm5
0DZWjuFSguTX8V0RSYdqfdlai5rMs3QvOw6bDBMjSRJFZxr+aElIefrpgVxFyPOW
FqLVLP5P/a2+7GkwlbxIeh081/Hl9ckv9AJ1VE18h+DAHYSIH/jyA9Mvf57uXHQi
hF97EC62DmUEPdLv8ZUseTy4zvYPTn+cY1AfqBPz+g0tOTbpQLFntlytv95/uOTk
3E17R2PIcuv5KPd4Ttsg+Y3hvH4TtKGylyRVhg66BMsmOBc5INZGqP1T7gDrxN8H
1SEihfSx9acjj7yICD2EXxe0uFFvTSBEasxsVQ53ILZrm2pe2WjnYOHOq2MqcOGB
aCO7UJO+YR8u5B6d95DigpId7oIDuV7j2wu9rBIKIC0yDSWjCHjfn4GKhRk6ZeCT
khuk78i3tmwp+BhuED1ns9UOcCdC50E+Mqb1C72uM3HQIqaM3PSOFbKqWc+RDZg9
Zi/xoKwV6/5LhTjc3IMDRJbrPPH7/y9fmbLU7Ll9QaYjGdcoU5sOv2kZdExOAWhG
XKMhE0EZxZaScFhSM+t/ljwb+uXkXvm1dk5GReFCX50jGVx/iWGttHSkTrn4O+O2
JpoxAfN/+jqHnu24avmwl8HKUt/owzf04RqV1fCyNwDIlSgj6CiFXK8Cccm4wFOa
SFxxDSpeKYk4GELzVk2uJqbQcTC/VgNNXcc4vPTRd3t4okWToY/r3p9DGAPwAlFL
NxtUWmirR67UMFkO+WHfU9agzulfZex2mliiwzPHVi79XRiLoBdZ8feX2hRpFEya
DmIp5y4BzvEmljhZlaKzESdbslPYkfUkcLyAg+PthERZHlMpeFJvh/cxIj4za2zU
vkeU5mutjXz/zjnlKS1M0D2VV0WOCyiuM7oLS/FU32CVJVELrRiyVe8lPe6z9r0S
PRts3qwXve/bTB7Lx1IC6eY9echnJGTOvV8yxGN/MC9dJaqz2pxPHRhJNw65Fb6X
K6JNbAvsHS4uZ+MYhWHiyYuIcROhkAKcFNnRp0pPDzFIDR10uzc+pFBddZpBmqmj
etEwUmw6O662u3v0b5/OsNAPB9Ug8eNpA0uWnXbwsuoAL7AdhQ72c4GKIOFCZca4
DW3Sxj9y7tY0y/MJpfdMqCvnz42NZ66kY20T03GLa2iL3I7njrQwhInXWXsxOf2L
w8ehxCF+6eDZ4T7AJcoTfCcNxbMtxROZhg0i67YXAbpZa35+IT3xvZ56f1iJX49d
MflJ5Fqu6wFrZgb3OhCH9x/d336BRA4wb5r5lHrWJSIYIdWNzeeHZnDGGbIdZsn8
moTYdgWE1jfHiz4tb/7AT3dexABH6L7cdZ3jkSHyEqEiEh1uN8Rt5Ahhx8mIcqnP
XpRFBuyE1S01pJK0aGxHXnkd5SqAuFxGWsD7C8pwkKx2to0oUg0EPv/xTIH74Zv7
wDoO4X6OLWkS/avAM2kH5O4UYyxfxL9CWX80ux6OrEPEqmH69QHhUqf8JTsVgvXQ
NJHkx1H6XjoRv7TEcBLIKRMdNBiAzrNttzd4oHa/nrFZs/CCi7+iDnBx0W6xSlqO
wKMEt226xpCZG/I9qXWMCvpxg2ci8/avPRCmLaysHgVqT2SGiclvpqBMID7oNO/O
s6cwzrne61oU2OguALxorBkDUaDvdvxoyhSQCt0YJeyScglgOpRZsA9zjesVnwS+
nsXZGVqxkG7lQUSxOZwjyiFXkWZWbek0a+B8x+D3/xu4MYzRn1mHxkF6gdIIpEnf
xFdI/BISqTP/95P9IS889j3NQbWKsYUUZMedAwefFNp4l9DROObMBrW01PZ8VprN
FrUYB5EUCvhGu2+mjC5lhfgBxfSN0hunqZjM4R2PEn18Bb1UnXhnedZsyRsXPKVn
3x/D8xJ7Zjm3r7RAhCcC3xPqosKPZ1CA7/d9Nm/hy0pFmRxpTo947Gmti+W34oda
GRV99Hlq3OgAHMBd7isEgxkEJ4r3GGLtwckEhCi4knhFm3627rhWzItu/f+co/LK
Qqskofu/04W1WA7+NKZmBpzc+KBqWyDofEAcU52kTdgw6rOpssVgNFrC1GTLVQdC
znF+snZxFLGM+ljvDefk9b7LgtRoZQ3J0gvy671Hfh7+5541uoc3JDcCLvvCuyF5
Na9t4l/rxxZjkYPZJBEJ/uP/d+LwvD1OI7iLBUJZ65qbcT+hjWIrPjYomDkTXjbI
qYakNJ/uk5LVnmE11YibpyrqpVje34ChMFIsvRNTyssWHdr01vlsPb6S5BwA2+cS
+X4FDOB703Y2YbfS95MHlHzLtSusMQmxH1iX+VQkQj2hwE+t0piMWt33IZ5eaS4I
iOVjTyc5nsCz5B9p0jGYHFMoYK/bTh/zt8pgM9qAe8D98Ei34GTAHqtEYpkOURia
73hWUOX1GrglZQVxq90DI+PV6bW1tJprIo829s5T+fmFsYJy5TxvqfzLg+EiZ2El
xQHr2DYFPNFu2sa++1ur7QKGunUxj4d+L1e9vGGuNOzRPu5zFnpv/noMdvsNHl/v
jvRuJ/imm1+pbni9eWXdP7Qpu+BoixgkAGd2k5Dr3+Z7QLB10U7aPCvY6JQrq8T7
VSFzHzIGs+q5UCgnfPsNaQhIl4j3PXH/VI8tIHWIoQC5A+rmwNCUcWTnoTshwUlV
bQ0vGpgRuS9lFyuE+s4ZkL7CDPYwfuJQ6xGW35m/5VA80aKP/vF/95i5rmBYfSrE
SXoM3oeNDwuvpRIq8CreE8X2NOwUq/KMxM1FD5fXAU1KOLvShAZFuVaBM2GAV/XY
kx1NenUMR2zLdB1hnt3Ghj75sjQIDjERDkBz09GIdlY5jI2y6eJ+p5Nz1alfGkOg
3g93H1x4yLl25p+C68CiYl9vFWlbzDUgCQs0/DuTlAHpI1skofT40iTE38H1JtGX
TUXrGcsQtTZKynA7O3sqFPnuAXffIYsYu867TKyrRPdY2a4p3hyctsqv7hrsbFk7
NPEhfYxiOIjugN2jUPUHrfmkkpeG9AFrelGY8BvIRSADxjws8WTcAGdVDmjrp5ly
e+jccmlKg2YXKqms7xWyFnKQUfq4CyHITtbQ3VAxdXME4cn7e4QhMCVPW2//9/d2
H8YUuxyPtJdgDnF5KGEnG4LO2dLfC/7kxGe+xZrwbuC6n24V56G7FYspIOaq8Ote
OJI+VfH+14zNyWZJ1jnI4qbg+FIpKn4aYfHA56JjX7K2Rz3CvbGVpAT6hp67HmEZ
ywbKrmMnGYtdB6VS5U9TmUYdX9jT3zm6u5DTBpjvuoDTh1FQ7vSLSqAkuVrmx1m3
RLn6ev0Sn6FhiDREKka+4zvrTfLc20FKvaoizckwP3fRU4AxNThPxtYh0qoomWBE
rEP7gE/BDaEE3OSI1KsyF7Ail4I+cxpEUbhefCGcWutjF+mY2AmNlQuLnw8grUMI
xHTxq2chNHfRWTKb0SDh8ffe3xvQLSsLBVMqi1HhVaG6i9kC9xGg7ImpFr/pXbFY
uvO8VlMCdr2r6TDES0TBU/DkxGUUyjLQ1gD1NriX/fDndL38b+y6iOjf5Kvo7hZ/
19s9vZUDJ1c1w57VhBT6Tdj0zAPrM3a7BUzf+qcuxRQV7Kz7FXkDhOSx++MeJzO6
sYj60tIPYAEiKIsebL9Fk4g5sZgYN/xu3r42w3xP2DOb+5gXSQwkkNJlXiu9tO6+
IH2jap+dR8pBrTFkSFB3S7WNDHfhtkf/1927oy0b720kWUV+JQxDZ5iB0tRplA0q
bQ9oaD5v02TcSKhSJ4X4K3KIWGAIkA375T7qDcXLPGGXDVh8N4eQO2n9X8p/ac8+
xedYSfo0vxkc4By/Z0msi58+vO4yVsvxM6756RyvvdnKdlV40hWl1FaMPjpjrw/4
aH0cH4wxfZq4vNFUJWw7T63EvRpm+KkX0vM171VEnPASESvrUqBgT20yZz9isPuK
FXj6VWUbqtFLB/QrB7gNcy3UD2l653mlWH81BF0ZbFAh0JD77ReoLhS+gPVShYWc
j08Q+8Wof7yq2U5TXqG79Mi0qKp0CFwFFXxFkTo+3SFxWOfqpQnOVBwTotTWaZvc
J6TOgoqnlxCUIZYWLQvvp/xqb49ysuOXsMnxGKydEpumPk8nnyaj5+QhvURtwbZU
0phEY/VFwa+0o1ZgV7lZWaCosFzIc3rThw5BGfGpBzkyxV8tNAlgAsv4iG7D9Gv8
/O8zAm1HSvYu5UDjQ/yH284SiqeL4He54kL86sfF2c000n7H6C24UhQc4ylPv3Ms
9iJ8uHoXB/YPNj6icVX4B5x2YD6X2ztv1q/wYW6ASoSpCyYSKNxzSNWNMn61p2Js
OXABSG14fRqvw7amf43oCgYJNXhnblKfprUxI1rMIEhrdjZLQ1Ry6C3b+vxm3bwa
6fiwZKDvoV/643sZLzbjowq8IO62iHYjiUo73sSE8KrpUGDrrkqUnqDb4I/Yen7h
juhMltQedNa1Y6FsEyfkhNAkqZSE1iFQp6K0vajU81sv1FCz8zxxACoPYBwSqjL4
UyLN07NABM+s/z1GufOfCMiTesBMfmqRwc0/zP8y7t2cf1rYVs7H0+DXn6hihjJJ
DoACrw2G1lv+EyOVu5TrlpYTV34TiErzuOxDBEN52VOWGpRpGbDrBJ2jN4xPsmTS
LuZp6V6kYjaJ7mpoFc2BIi04Sy9wyyva8nwlWm+b/au0NeEH5KCqTJQrGK/VEUk8
qxGRR8wg9Pt63SN767TkS64nXlxsZwUDBepwvgs4X93qPMQfJuAFy9fvtnc2ShV9
ltUSuIBg15y3ZnGq4H/8l2yI27F3Vv0w7KOxy+ngvL9dlZKCiRH275mVZDqr1fXE
hvuDik88f5fZx54yUZ9sPhcDzcMNkS/ivQxiB7ku1PBQ38HIFq1YXKXz03j//7xB
JVB0ew++Go651C9KjBMNEeN2NTsnhafsfQ0txKFIu9CCTV12rwBKaFsvTJ7yBcNT
B6NmtkESZ5F4caCGx2mstr7a+PC3ZkaSSTw3NFm//pfPjIgPRn7FKDt8XZCk1NI9
/4cy3DUJqTLznLdK3jL00S1q92zkt3a36S3HntGNhIbW3Rr+HgT0b4kwRBbx+1rh
IeXIPqU8ymlquIyjT5T3m1v5cNlLcQbQwqS0kTjldf3HTee9Qy14JUmOfpaQEu4C
G7e7Noq5YHlBAgTfU3it1bdC8XFf9gfUZ/JJKhstjTFsAcOElKH+YryL2LfGKxbp
BKwr4dnuLFvoIP0GZL66QagK/LA7e0fygGiOcZHyzm2Hqkekj1Fl7M55ofG+Tt/7
PB0n2VOoMt23iIvq8isC+7lV8HLCSAFI9EmeihCHDabADACDy3rp/8ZSKPQTUVtC
SFE7C6Dgdz28fr31CRaJ/qMw4FupJeztNN9bWlqwsT7sfv2gow+lSTA82fcTdS4r
XtHO/ZO1zAVT92gaUhzv55jGlhHEF9RJ8SEfIRC60AFskGpkbAR3moB1UFDo3722
RVvNlAVaHgk7DM9R4ItqD/Gxuo7vWm0BHDNzNecYIwXg3pVc8BW1eDd2Ggpmtad3
C7hjse7HnDo/z2xcPNCOlVpI1NZTbOWwZCAlqSh8ONcHZPGAU3r5i5obWq8Y+SLR
nq2r6uN3MSZdM6n5i9ICCONP7jfCO2NZzbTeeMh+45K9izUa3awpBQ/L5t9hsBAE
kb4+9HLMCRjvjcovyXRmtXar41wk5IQ/P5XaIshvRI8NQqdGJ1BepoFC0nBPoY1c
y0ScZbn6B0vCWTIGlWCgF6ufPsMSMviNARxCYi3u6ed8FMGR2ZGJNHt5FyXE0pcJ
UM05NW7REunikU21BauKQJbwftD5XnIvlsKE37lYZHjZ0mmap9urk159ISIh8Xmp
InRJYRZyrEhfhcQmp8ZY7GfbQEpHGjLbWL/wOZhWlyi08H3NcxUikOfXlaiagrTL
V3I/yhVu5SO/ahEkizFNwbWX/KAzhy8StoTo+fDm2aOXXrDbVbBTQk3b1xFb77YF
BXqnISGoDxYVHbu6WpKm5sUQ36VuJHxNcdjdcCNeblHrF7XB8gy+5AG46Ix8n9OM
LcE+xGDPiaBg9zKwATlaA1jBkAmeZd3R+paThYwXu4np6dE9SJktGu2sbgi7kQnf
few3b2egDzJr3QankQVljTyzzG1y08owZEgugsJqGS69DUReZa4C4JopkyRzwGNN
4iUzZFwwi3bgiIxNY2oea2gwR60IcJ2aINQO6bHB4/cgMjj69NckPc68I2hO5ePk
Bp1Dzs0pCGs2dlMe+1JxA+5u992fYb1Wzx/6DVYBmeXV/gfBVreIb1ZhY3iLzHPv
FsyB3rthWjBWxtbnQVAXOUDyvw59Sofy8CH5EwIQf1uvlsOuNhzwfjsAOKLN0BT7
CihBMal3Cx9zvOxTDmLjPOfynZGiGMBTvQMlb3deIi1ycfsUOlpqbquW8ZIr+bPu
p0pwLwMRANUFb83chJAI9631NJl9H6oziZQ+E2rqIgv1+u3tSezltUmPCnSEu6sb
GEooKi4iGGaPwL3tq8hZ0QvDF+I+Jqf08kvZp9p9G2L0EPtAvsMAfmMX5NS/Xv9y
3ydHw6/5q04neT9hVUsoLFBN2GnrgQhRL/vC1AFR/BLtoXJQ98TGkN+KqowFKw6A
XR9Rlzo+f6dF0jdwuJN+mx3xGf7X7Uj7fD5Q4JYetOCJZoVbo+Ct9YfBa6s0lpEh
vlzrv3dxfVKn1Z8Hm9QEBRCaEQ15SNJcdawY5nsQ8KBbfummekUU0UFYXX5Ymxrm
/MlKO/4IALsicLl3NpTB8BhOyc4hVApGyYSspIr01fPgXUEoowxqfEhx/zvaQztb
C+SIiAqxiYLTdVGSctEeQ6NALLD5jAPbrNnlHwkmsKSc1HATQ3bvWw0L//kA1m9+
UtId2NRiw6l0XOBK9/pzK1c9yPryJr7rmjcM6W8jHF26Dox9RyyJCCqUddXgoSJK
S+3hR3ZQAd52YG31kfx0UEdQ3fxTnglyLOArUfAp/dgKbzQKcIXjh3gmKiyloc3z
IPtJXfWR4fel1LuzLt5eY2FDxtI/rOP/4pczCmgDyS52oRqHPnUSsV/wbHfmcWQ8
nOXpZq1VDl2rTOTXqaCqaKNHtYY68sJZD6o+Js0vzCssuLkWWxqqHdF2OctKmnL5
5EIJc5NtlpOK81q9S6emE6grnOEbw/Q9kOiGrKls77/fctABCmL9uxZmyBuJsAOy
0CPS5zm49E4J7WHAlOUBHdl6ubsRuvTSffNsPaKxvo6ndk3E5ZJQ6JuRHkynD/em
mj6XNjoGcv3ZId0ODa34Islq01/a3jajTqJvz3b+jWxFuhb2Aa1fGcugjTzCe1pr
AELprJm8m4KKea6vmUPMoWIyh8qAz2AXMmmYznndbJgBLINiqa1015hzF4c263d1
dqnAvpuk9YUqlcDmyhM651XnTOiLUmJ2F9mCRy7nbjtGKxv1rEc1WopV/qF6IXLG
H3iWLO0Cf2XyzuNIGPEkd5AGECxNZaCllpyx3dz+542IBnmizG5NEGQTR2xJYIiq
45i3kg32x9syACDsECVtZaBi1s+LM1RhFKhwNGQdDrLKyaOXZ3OCgpJmwL9s6sK9
akXkpEUpMgJujJjgdvi0bJU39+bFkHPsoqoG/v/JEgZ8ZPTHiREiOzyQ53anM1WE
DcH2HZKFtAjnsD9hfS/aj33o8/6/xOgRhgLvlFtb8fmiVM/kdDfR9iYsIlTiYr9J
ObIy8zH5dDaoaV8egGG8j7cSb68aQFecXPpYEu3D/YcsOD9bPOjC7WU3FmiY3enp
rxZTfzxuxH7HlwjD8XtfC1iUkM4+isNJi0cwE0Qna63S/KWbhONdE2rWItIl+LZS
my0M0ZbNHylfB2mAok2nC77spXb2u9LztQJlmKnupuw1W5ypDQMV1yZQ5zb+Yzov
AA2/I6JQarns2RFSqsgiQWQLp6MxBTSxOk0fIKq6Kgi/I0oTq+Gk2T9VDhydeI/s
D7gZH8gdi6vo4EBVU5AREwU4xGBAFweQbqvigO2B2dcEJ0xMz74DoM+tVZwsXayd
9kUhEZffO99gyM8h/Y8Fj3A2ium9qyS7TLJ3AHVbmZpO1RYRdbEM7yRPvvbSnivw
0BhyK0MRTQWrG0tUr6V/egWQSVLIhxxZTIwDfPfavmhiGkXjf96cu66X9zSt/vKu
bz56AiHxkADHq0tzemuO/DW+qPeEyB1eCWIZKWUs+tLtKukjVzmg3EeeZBcrYrOx
ty+xQWNgcirPJUVmJqkwez4OgBXeGt2SL9K+GiIQacyOyNUUagspCgRkGfW1W66H
lFA+qDPH6dRz6KBVkf7HzWM80GC6D4V15hvW405KFcUEsgrO2mWvvLu8nWN/Vu8Y
ccQQncBe8C3tb8AG+D9J9+ZrLaNA2qe0+T5Ztm6omgrxz624s74Z3kwsoW3HU17E
/OwU4i+9wRFno9Mo0TEiaNgc811NcbmOZa5elvXwp72aztEU7vPnaiS+allZ1AKq
BPUE1s457BS5id6/IRe6wTpm6hSqmdEikbiF4aipv7rfJTWqKbJuNt+RJ6zz+uvQ
ydFf7EnmjBIeOm951z5WQ/8uMvPrERf2FtKUYMujBvoBaQ3ByClUTAxBMaxXzytV
KryRqzIwLLvcdOinw+RFIa8ImLfEebmPx0DoIzs5hQUekFgYrR9/dlegiy0cttqe
yiv7FIvgCS6Km+IUNwbzmVfhVrBRPQtA+oCaoAY2lxFeZ3sCI4QCaUAQUt8M9pxm
PHzNHHwqsbdwJ7w+VBuA1S2wuVdrA34bGMYBmUdbPkaus1d+txW0WYKOHYbwuwGV
c4uId8OMG3fR3SgJyX3Rz6Qvj+q2f2QrREylZ3b86vYNESIprqiRP2SBS0PVJmGh
p5RkD6DgqU5GILj5JGrGNqrd6joJNpGPoVs/3eb6kALOAcjag0AIuaFlcHLSCf0R
QJEAVPxuOTBelpmmuPoGQOVEI/VEM0sOyqhVaibHZPkG1uFu5NuSN0nCb3myW3te
9s1XAYUFuEsqXJc72REbs3gHnMGQHgCrTSyAEMPTJ96vKk1/mJN41EcuU4Og2m1z
JRT+8ly7NpKuUE6wILFP9FzxOV0PTUj3OV8HDwh4KL0q2Ry1KRldwWxKpzTan1Zq
uBqNGmJR0wgiILs2My6rt/4ddp+WRP2+8JLvdzx6IL1lny2TCG23fLpKtQrYEiXm
3D5II+ylbLsi1labLWH0h6WEAUzJVuwyMyXmlsjJfZgYlyGf2MRM2JzFjBS2peQV
cz4DoDR+8qu5Cdl1DNQnpizn6cukyRak2Tax4KX4jqMBgLwRfySQ3eIQEEhDkC8w
iDuivzxbLKZe1sA1mgKfMRpqKTpQ9D8hhdK80PpRbpI7ev1acfWvhFIL6u911c5n
Kr14gWZfLJU7nVRC/10XdU6PcrhmYYXEJDpRhbRUUh+Rd4jFtUwRoQf7v8M3XHR+
43FouMCOAMYfRx9zGoaXQO1kj7KS49sNN5i4EgYmCFFeQk1aK7R8LT3Q/X3qzfnf
TENT8c8dyGCJfvePPE4Hb4shFksc1bsEbd1sSmTnBoXsQhGlbFlrwxyKK4tfsoqw
cFO7xQf7+q0+yPFSzQAI+z5pQM56vHtJh+oxpzG5W4FGZbOQeQNadYeRYtO2V+p+
gWnC4oZ1NKFgik9A5njG8DakZhndma5yaLbkFHkM6CVJ7YP0GisJBxP1nPFfxEB/
z5629COFBu5ht9pGZzdU6YpJBwcmFsSnyohRpUxEet+kEY2ApraDBGo0q4zNUQH5
Wz0z5x7H6WV5GvJScPm7M8UoxcxHINOtGtpMe47iHIwMjSGfDgrGZr5dgXe2cDeg
uY+ReVvJVy677APelDZ75de6tsBg7fOOPR+p72n4Y6hvsVWOzlNmbPngYvd9QWvP
bbIVNApfWgY1vhxa0A+Q0NNRsrrO3L7/9y3ocvb3FMOheubdxgc/a67+QqtAumzi
PLrhMO+nIO+WhwxSDDqRbY5RCzJTXX4fBDuY3ja2WANnBXQbAUQE2gKy8Vk/lRkg
GSDo2Ir7ING3mreEgYqZO5Fdx1IHqZ2FWfRIKENHSdWahhCFgYet6e59bcSfLwtq
vAISetAZAVY5ei/kHX2sQkDOXqzOTkDacjO2NK6eGB5Z4RTqfXRK30UMKj9ua9+W
k9FDoVon2s3kO7c9SQbgIYN7t2syR1PyK33+O0fCA3ELhGwSpwLOhkXkjW9voyvs
lj9dsv5RQrxBr1y9qHtstU19WDgYgftNSkL0D6/2IyVXKfaPsvmFeX1QPXSTGKWM
meoRGREMFVp1HwbpxNRv7nZ5x2zcPUY0mGc0teu8R0idUmXdM0G5au+6y9ckC09q
gDApIeJuM1e1LBmwnxV1eKovgCzEXM/+Vug7rFs5+2Vk9fHkyAigF2z03hhjAN9G
h5TK0PrB/qRjf/n1qbzbNApqOPQ5F/yPwnhxaEDkkk1vsgAdTP+gX0FrIA15siBV
9/fMkH8oxZiqROiISAeaio6hxrDB5nx4yvkyQxkSCJlgRgkPIj4U1lNorqYNXNFe
9ycIHrzoplDjlMLIzMOFMr6aqBv90pDmLMQrzrSznCwNOCKmKrk2bzac9JlqyvYG
ZD1inh/TwjftorjHsGHZdWRPNAwpOpjoloEGK6Eu2Sm2wKY2cZwSUDKMAxY9jx4E
rkbRsSGA8omVfoYNipcNtICxeS6zsh4wPdoBBr+wx6SJ3bzBgIvF6sRczljeR0sE
LRM9CJOTuYRSauIQCUvW9S7Wn8oSShsfoQ4zBMDq5R4GgFIQWh7a7jllyCCx/J2l
OND+oKq2sW9wPe8I+msy8PP71TSjNtrBVlJESmckFKoaLbP6znn3bY8P9xK3CwlB
tvu+C+c/cMxj2cJU3Czh69Xi9pebOBBU/qSGGoNgQnI/1P+y8cKfYKSI0LYFvMNV
I8oiacShDqjL552kkIWqrtseRXVrFZojg/Soki9TVnX0oLIFTXxTpjUlinG70/Z3
ra9tYQuRbLdAuPrX2ErSgQlVCBond/pcuq7w5I8Wv4Un2BDzO12sPKh0MScAjTKF
ffAUOWeIOrK7Mg97C2FW+hoBKgFS5FrGoXH4HZjSHvqyiJu5v2eaoOBdBF9Ypo1N
TRKbY/TPfwyLMn0YbMiwa3mXx49sT/HkPCzPIQ5ZowSR6swUFFo4gbA9blo5vJvx
s/seSCCh56La1ERyp8ZePvOEIWSTKZenmNwtGGCtYHr6TGUPNzzdyqNYLYY17WVz
p7oIebdVh38Hb6gL/nXXf/cPORRjF8XK3gUKAAwcLAs1XiUtGDtq5XxsD6bXRex+
Km+DKhPqIGpS4sEe/9phdZd03KnQfqJyknddrBXi4D/51yyj1oMY7Bx7/3KeHJ7K
YnosEo2QbHheiHMlK++9lKF3uNigZYWcRSLr2VgvnLdMCIYUBqEw1Sd87sso1LfQ
K8VCse8M3J1/ywetLB/f1hJG+OSbVn1jRHPYAXvRPShGcptLTJudfA8oTePfO+c1
hDCBi7OQFtyWwulfkp1DuGWZOyugtuEmKKDNauU48juvGAVzG9s47/W2TDys8lUA
PhwCHwTxmAMtsgLxLTpXRIGb1XFXtZvTe6QW3zfM4NND0v165lVy7d0Zf2qtg1f/
T7ArvezceXa9u/nRZwjbUo50Cu3VW76qt9/Ak+bR+8IHmB7TXCitdzJEdAUVoNPz
78/p3RN2ondXTOWMz9SEkywh6HboF2QsYp+cBp+QBEX5j4VgUX8D1o0yRT8uiUV0
Td8jVXMb8OuSvfX2e6CnxmyUcEwGflOBdqUU7n8fQ336xUzyBYe/SoKb6lOuMiG2
z0h1HYKe8gYFCF25noD46ZZsHjx+4/VOETSBNp6RYGY1gScBRXZyUgb3EWhCBH/D
16dSTc9kWBSOQBXdjlvomO09kXIwhW9V9nuzfiN0qcIyQmvlCPGTgc2oCE3JvSZQ
qlBHL5mUnJ82Hr8xNCR0xFayu2Kg1YQAmrhEyoC8iE6ElT5HUhHoBK7TKSRfVRG1
YG5AwPqiPOc21PRuzOoC6p7DPHuUxCYveGYYVeGm+hLAKVbFH33vjZ4/8jZcwxPu
rX5pPUgZrVe5v0qjMzQQP63Z20bOb5nyClxgLKUT1t2mxR6RjuZYCjNhAIIg1LIO
IaitkS9sg7dnWYNiobTuWB/4zP5VbqeH1y1k2uEFQFVLL1ltxsbWbOAwtXcSJpFJ
GCBCwwrPSftQ459sQM4I0DhDAZpA3OXVuXjp9WBoFXLWC4aIXr6fJCgm8QD6Dda4
EiJ+iKkOCn1eZ3ZFJyV0onqZxg7zObCFCm0y9r9hFK6ETmGD1QBhR4ZDnAcFf33Q
W9LBzj5/2q8F4CfyrLE49hZPYY+C994RggOR014tyyGzLaSWKN/IfEpBRUN7qbww
cjBfhYhMqCFGmxx/6TwEK1uCi2qnSk75ZTkEWz2cQ8NPSXSZM5dBFmW/0+CQ3y1i
nQg/kmn9JlA8pkA2Nljoor5wOm2+IQq5qfAExGowvGvI79x6bJb6Ehxkt4Vq9vde
gmSqChYw0gbXUA2r1Fn+X8vxQNCJX9uncSb4tDly0BGcZv4YY7hn5LpwmpLlAjRT
w9uaZKvFX4JP+yHyAFRyS/BgRXO1pgwNcdxSZlQfLOZkKLChubtSLdREr1rnh+sN
3sr6fVtV1wJf5pOZX7U3z6CBjhSpSfTtp8suF73zhbLuWemcRn+iewa3UXfxBeUt
IvND1o2Uyqs/fmpxciTK6oHNu6HY1DjZF066BavzAhRRyk0w1WaJpGomcyirk9sX
uFPF7vsrdNdIxCBS0sQmTksttyfW4Q6DFrV+aui2cQrfoOIqJJjwY+JPfq0vbtLO
9vMSoO4DYY9HT/kpvTEtPCk6lN+1WPW6Z/bCSOsBIV/G1F1ifdd74HlpasR1mOLf
1xkkvTsIwxErRUnegWAgdRG2uoWPTIXD42QXP6cd7Xw3116C7a1TOeTvXBe1M5Wz
fcJFyg73FajsyglY6CZVMWx7V0Qd3LbNwIHg4J3FDC3SKKT7RPN2xyALirT0C1n0
7ZlMRAzLhdn7W3aTiWAhmykHPa/JbKS7RWNRkVC6gWdBUV0MqQM6VpBfGly04qrq
cOdxyy+Hm7M4lh8Rt55JKxq3/sOkaH+QUoVQkiPDhVCJ25DgZ+wH6W3RnP7grw9k
SOGKmQzXonwzHRi38QvukSLbH96184bz/tKlkwLu/Rfs/nh7joLqb4pefaOXsSWM
Q4qSXo5fynh0pN4XOx/v/I5JBHZfWSUImyLCuXvsRKduU3sVDWsto+CinaEvWWNZ
wiWCKzOHERCdPbmnzew4T3fnH8hamiKs3UmTQ/DRqLPblyL35WxcTxoIzGhNTrvj
u4MZVEsT3bQaK7Lo8aC6xvi390Vo1uQpLLuFZAH4Dx3lmSiGdeimxonr/FcpbKiP
OMy3qTsTnQQ2nMV5UIoxRUKDP3LCx/3BcwxyJu3UynvTl801Sp8oNju8iCqt9Rc3
K7CM51zs4cgCIz4Y4nzSHcrzXqiyttIlSxIDv/29rq+/7xkeGhQMFuYRpXGnzNg0
NwKmEJvErJJdwReZFbctg8uPMGzDVm5G0d31zjRcNRLWxEHpiaafVVS3LqJE2fcx
rsZHNGAU/PydU6UFg41YjJtCb2SgmAqNrh5rmKehuha/mYAAG5xie2OMK+81pufA
+iq5LRRsVG839qQMZwCQO+diVBwfu0QnNn8Fzc1EzXHtayFNUM/Y25AUJp//S0IV
+4K4sEyucInGKQwp/h/HJynQv1KgFE26HgXEaQ33rXR47/S6VlwehsIH3NEz+Ml7
vF7a5e10nF2CfbwHebUDFkjuVomub1c+/BM4rzANssnbUF6IbA4C7Z/dLCFlXxWV
MKJPLQeP6ZrZMXwLg2VSxFQ06tRIXqVgKNRObSQ0HA0h3lbeZBWLun59b6XMYxk5
dYFcCh+thMCAQEkfrnwO2skmXr3cbmr2BrWW0PCQn8+1pZbdQ4iQGnRfTf6hXLn4
DBusFV7GT/JwCE526f2SVCff3XPF5wHHbyOAamYUjTfl034Nbyr4/jELYYY+x4DG
vgroHwoKzD9SYPmq1vb5PyROfWk7jMXW9ZmLSUIKwFpxS/UmKrjUAvFE3FGVVVlc
5AjEvky0ndA1C7YTCXylZlCE4rhHBhoQ28+nCt6fv3mmQmMpvbBT0dyaNs5SU3Wz
Z0jJUuCyAybBhR0HcQ86D6ByK0NozQKfftPvFf3oyvPjg+fTg3FfYdM8uuJ0ECR1
r4DPFZetOX/gPRuktsebZyw0u2x4eE5RHAwAEcyD9rAhqNLuH7mYfaiWQwvky4zm
XLSzPpmAGxZA24bmfh81NtZ2yxuAkRvhiX5RFpMB0uRCn1A6TschrqD+w0shLeQU
5to3KLDS/c+LDQ3eDZenRtA3caOY0MtpleM7ULqRukunkRZvoORkXZObaP/Gf0uK
ED6h9FAZCkeB+pgptoohw5d7Zwm7x9xB0PMJ4IwBqr+mJ80jG7EKE18INcSGen3j
FF7c907yaKRbHj+5jtVWbV3soopSM6iMg6hwr3lYapo+c/Zwrvews8/H3ob6A0x4
oX3TIGZUlDceEN4lE5GzmetQCfXKGWegfgMwyIcwcChIygRb5VUra+NzIPzBGBRN
qwoc4pcj23aeKJnBiMM3bdsAMuB0FrpCNjw+3O38eq2QkPAITxteyfWdOrElMdfi
86L9WzcmlB4JfxqoS8xiBUf0vF3rvUYhxVjbu1BEcIDamEI2dLoWC2/7zyQn4UTN
Gc73NZjhNLfvdnVlwo7YghoLvdYLQCvoYWNtPHQ0Pj8alwYR1aUBsGGQAQnmiu40
Jl25Ofni3QFbLTPBOTiV3H+MII+IuEu1vjeyxZFPj1u/EkJwr6bn9FLQAvQaFOuB
J/QojFjSmA1ScI/Xv5lHYe3c3tQ+fPRZ9WqXkxNj3YAGcLA1e2AEyJFy4pTr2MR2
JDHqWdVhrlGeuL6IsnGxCHMBtKF5ixyFjbo2dzk4Dr+fLp1COzeLYtjVu7chY5co
9WmzGM2X9CT2zcyvY+kq662uuulOjXkUv9xzJiJMsuXF6MDLd+FFL0JKJCbXqQet
Sy84fp/w+vr7ohTp+ICuJRvcTCmT4tAms3kQddqU3wn/gl1Xbn9Eru5mebNaR5qQ
52LaaKqrFQfV382VVkksSXMQjR1ifBioS6+QBiaOAdsT2grxoQHy+PCnQLR/tYwb
U3XrCWumraJRNq7+NKtEVnt9ofyDDYsJJ+yJngZO/+jmmz3TlAvQDXJADy6ktyAT
Sc2wMriFLhG1GcdsROqzFqS3pjbTN5SigEfhvs54vFxWZ00x7ElthLLmG0CJbCq2
8R8yh/l+hzapjiCqcxRjv1tX6KLrns4LpAmiNADLI1FUwW0U8zoT+CNHxra/Bz5a
1YVaNNE2WB/Snl76H+qvf6ix1/9i4EV/eKPEzgGdRJAchgGXCzWj5SAYMxooHfa9
rnl0ENb+cL0BkRDhBBHcxfEXEeq1XPBBH1UtZgwfLkD3c7b72ZC9mONxU5g7ArCE
KybdXI8uMDR7IkjCmutQiPtEFKCTzaJK0LqWFx5O3rn8/Ibm7WTjK8zCJNv2cFDy
J3XTd8h/nhJTjqG8H/DyjAzAC+eooK0Ga4FQU36AJInKvaTzRRi9X6dGR4UktU7P
oY4NnJwcewIyZnugsabAhEWgm6qU6OuO5HIyxf60CNw4/Lb3YzXGj2T+GMvNl8Yj
VIDNqQ0S1LruLGgrkhVLF4Vfft0ek//Za6txl30oObSbaVTwdc53xPbYBoChwQSh
m3En/HsDiDyo7dTxOjN64t3OKkX1+zAhPP6oReEL7TWOCfPdp5wxyhqarhYZxKbX
gHJLp2X+bGwFqMAZGmoE0dC5jgoDBW4Ov0JgnU3keB+bDrS4Rn5rvaIUnnNMq9dk
faWL/NO0NtjsJS8fqNlwflOS5okS7ZoEAYG27B/bu/hUrZAfo+VGlhGhxBQb5n4S
NdLXb4q/MO9NQI0fUL4YGkK5gZS5mBHUvpYHwyrQun/S/7bXeugGmYxRVOuQyYhW
lJmCGZA/3+wRVJfp5VOwisHLHUsPINOr0UKN+dedQZS+FpyqDYcq7pMMOKVJJCFj
GAVtq/I9cdGQoAmIzl8GTlW8nq0Nt0J4pRm50d2aIaRB+HMtRcTG9YDo2JiqRBDj
qxHUTnNsEEblGbS0VTEdiXTDD7YbtCsVqzeEuIOl/XMmFfHpDa16TLwWqEUlUCSZ
T5/9HUhAKHJwPILW5iPev2smvnDLflwFPRmtklsfBTjbvsNfKd9wBIlRW4WZ/CSn
2Owdd4Fvf/llMjno4B0q3IoLexeTZNPtizSvv0/glhApmjnJrBqRhDVC/Xj26HOt
KC1vIX88KvL2mWpjXxuHUGmV8jYd5CWLbS13cOVyak+IulWp+iYvgaCFV4j1F8LP
FyI6spjDg1hrIzymT4Lzi8PrygI07O5wGQ4F0FyUd9DzWvLWv3XaP2ZOvP0UJ9r8
isrXK/JAsQdAWxodywkIjpiS6OYzbJavUe59gSaeiBt5ILcYixnfSSDiYn9Yk9Hx
2OL/ok/MiO0/pIP17lzvkZAbjmFXFhA9o0tBzyR2U1SpbQdoMhLgnmsyW/gBiw9h
E8/fT43pwlB4/yaJttSCCvWGmqrQJziCwvaMEfAskXXN3o8mwA3eRGMgCYWl7gdH
/pf75gBkyQzBHXIpjfBouHZ4MeL+cfjOX212Qg/i4ilapk8SnyFqcdTmo1NoozpD
BBgj9QyzTmrurWPgoElXqBuEEa/28grF7nHOSPyY62YHuspYXKqRIa04JE9wvp/g
9rMtt6Um+ZSybGrkXPfRwLgH9yGHfUJdO7mYWYLCbMFV+eZEFSn2GCcWlFgWyFg8
OCqTCc+YAFzRfToelPlI5p5LC7PDjKhM5B+KOu4PafKHEXDUoxg+U9tsHLslLZ3h
jqmaELFrUHTOk76SawlAVm11NDzKBfEZk+FWp58czhidWtv1G3tTHjlwlqeyricc
kkZLzqqcCpvTZBwxwocBMhgkvxCdkyq55jvtuzaMKywA5dDR9Lmc5pD3Uuyb1Vom
n81WuT+PAlMsq5oN1bff0OV+KW2+NPly5B0kNqdE73+HboleRyz8Pr3zjdg9Icak
wMaFZJ89nVFtZo3KDSdBWwY+P3XxWMw25EiKY0FJTyKzkOnqwRGS6oCvqbPABDHX
ciLnEIvEL2kFaFCUyI/BEdb/2hXmlgUQPncMDuTLWtJYTlmPBd4PM/O2G4UFoJn+
pPHQBA7kWYoearl581ZnyiXC7HwKEZiIv44oaFDqKpD3Q2EsZbVzBnVzA+Ibsiuo
iYad4nBEWVc0VpesUWvtKlFm26oOrmeDZ5QKLdaVm/LH8yKP6QSXJWxy/oENXXh6
wVnWvaK1CsjOxrA7hoL5edXjdlyRoHf41DXmDhdYfv4Q8Qc08WSWPqnvOiXVW9PS
L4EgrEdIMxWEzoGFu/kFIDyI4Y4iHKV552GknLqeP5mZiR74bky6Ak1opaKnBmgj
UDfZspdc13cRpNJ+z4CLFDodfEUhKx6TJeQh6D77bzm3n+AQByyJx4fhRqXFOTDs
fDHAHHoEi5OXwqcNZCrG5qa9kZsMDjJkHgLUGKdIli3Z9zBPv4+kawOg4OJ6inkr
Sb55hRDt45pIUJUxC4DRYNK89rHGGrmFOUBHt9trWZq/fb7OP52CzvwhuZSAVJMf
2rTg6nBSSW1AFaeEGhC/nE7l5VySWV+jB8EPR9jMn6mQqyh/iq52hD6cy0pYjX3i
cwHX7Bx+9gmFKoPhYxN+d9tqo6Doc9j+0+AL6tErr2dLeZq3GOXAygWbnb1xX9sO
ajYzzdxTpjR3QYU58Wm/UkfnAU9PXV7mlJWofSPN/rBoWmX6W+5JAlt4hMaxTD/s
+rIfeURDouf6fjltwF8cRAQI41igIGO/Owfiahgj0IHEel4/AMuD7XjfkHB/4sas
avadwxCC0l5rgUdmtTogfw8ypG4lrIwbDSHKMLirtg+QFexPjmU62w3c+sKGTpzy
9LS+m9qDon9LQ/T8e8Q/DkFFP3au08HRxeXsGrfYJAiYX90r7UhJGnmPbVGj0oSi
uXLsIFLEtkrMntSOE8Q2p2A1fQSa23hp0MT/TFYnA75RiiYlAmgcR4r2YEn2+Qus
3VJ/lP3H2KYSWUXi6TFm8BCTPeac3+iVYKowQE4+vDjNSqfeMV+qzL5HVGGv+MNk
gwO6ZBqIL8Xg/HgB9j4Ow581QClHmRkSk/ITBjJ3lrWr5qTIVjQxrkxiikAntudE
QjMxM64XoMB50L/ZWDZTQHfyWodG8srrc1bRU6z/Qz0Fbxg9NmLAa7tMyYock/eJ
HxkzlFmUdR0Q8m40F1ywNPK+UvRhA2kLJvOdC4zo//Sq+xRoCpme+j9tPRFzsgqg
XNNSgVpAYuRiD/sm8cECu/qgm8uJW7xyKvdokNaQuIHoyHOWp0H8eZEOhaO1TnTR
gp+CjISandKNWpm9DUF5kj2kOLkXI31RrStvlf+PmozoaCLuRp5lYy2h8QYXO4n2
NZanVo6S/0AIfEqlXzuFr6bxjMy9VrTqHDXp2pTj3Xb1VzR4Vf50h539d+SseI9K
FyncYVil7PnhJ2Ug7P6XUSmCA6GKkyFAWRAIOUiKsBXzT16NisYqKiRj6z66epSs
ih31736L6QY01Svbx/0n+JJFImdJNvC7S+c9ghh8S3jUVPGaR3TPCHTQB08yeNvC
MFoeR6acKGe56CSfvxHDKH0DGtfv7yeqp7FRPZAwWnLtj7rDmRTup6DzMouf1J7n
7kfQiYPYhhDzRbdE/1gg7DZ2w5bUy1XxuXkZB4rrnHwJy23TzJGDNtRADqB6lQrz
jetKB1gbc7vrB8aWRrxmBBxAxB/60KtFRKWhnymwIgPMSduH0E3KaBXuOy5AJcJY
UdVolRz/RIudPATYB57Yxk0qFsdKdl34A+SWjP/bVDMFVB+aGHTt7Bsy6X4jXIPx
fdb7bb6+0ZtONZgL5mfFejS3ZCURcJjdTwS4T/AtnGqWRwb2ByMNGQoNLPtyzoMg
a45dTY7JIA2XK7mp0NgbnArf8AH2iWhY7wdBBn+dr8k6MQ3RX5GLeiWXTtxsEfzs
Dgp0EZAysvLm96yocsG0bfQ29EYSwg1RtOv5LddJjQ65ChKsSNAGmP1CjDFKM76G
vVzSFFZZZqhudN0pZqNKzk0xBdYntJ4U+xofNuC6jlGlDv1BDl5GzllEKesvif/i
XC5tNFjrgAP7g2kjrZ7BU2tYQmK3DgmplQ8Qb12HZ/bSKBvjo/+HkrWXbYGGQo3O
0sVPhIMj40BBDfQXp7KUyRQ0Bb8l4MLdx/3sJhy+OxSyN30XSt681pIGRqyjlq71
1uhYymnc9tDuYwwXt7jHdqkoR9t5K1bUfuK0mevMgzafbteT3UX/53NeFdxniVLu
9k0LuJRqz+sJborrHmNZoxirfXnJ5dBzKtosdvt4T57zcmo+p+vtync0SJe3fd10
LhMeOzMKGJe5WAVzBnMaz3xNXkVmWfr3hBOrTofpDQ8nuULNARApWuQ6km6ipvOQ
s0hyXcMhXiqbQi7Lz0tncQaOqvoyf2tSBaAqzUrxs2RfaXcWhxjnFYfy09MxuEdI
+oPpfOaFwiQTfXZh8LZM8g9Q3FEV3HcHkdcNa6eIHt0zGtwBQ4Q0GSa9Vjk5Sdba
fAb3/9yU1dn5nGSKSyhuA5F7puv8aderZ8AXswCQWEgqnNRJDb47UU70wEt7Gf8m
6L0x8WkRNJvRBSrkG8f86N/Y5sg+E/yLoF9hOIqJoZnOgGc0/ln/ePMb4kdoiI1n
ut6H1rLxy5Vagb92W4ryZEBBtSlNVODzLu+JC7MxXPK3ZAt2d4Z/HC4bbs9nsTkA
YmL2iqSWBtwiOiIc4vdw1Xy7dUZQzmOfdWdW2CsgEEZVE5MfYMxfTipMNlMnZBVj
wfpQP9POwuVr/xxSmlXW/zM0N2A8spncz19zSWHA+LOA5pM+UD+WqY0XlJEncWR2
ISlE14saRWqarPKgV3rPF80ntJMMqVZWS45vCZ3yD5kppQp+I6KyAojPcu9MLY+8
qGSawradZ0+5Gy22g9/mR+EvQXOrZzaM0ZZ+7euBK/yJQn+QXvsLBahPsnyY4ebn
oTiVrITcJ2IWARaLwfaPmEOycVPSTzqgDUvLnndsXWk/p/PiurVnG9JV9l4GYiNe
9rYIvzOO3/7F07N7GgnLJQdXHAAZw0ySFxy1mUBjZMwcFkDMs70M7djy0nZ7Oe55
Lx6UkBjC2ntfd0w2NUBSKYLFP17a3BVMh+dQRmUbXZ8AWtrPFKgnHRCVOdCXv+xc
2K9Hdhi6Qs2xe/Li66pG/uCHVKzywBNnWLxWigOFMtZCw1AeLCQiHlkAQ9zt6Kgv
z5icc4jZJzPIGPI+FQfwoUd8G5NfkwAwrWfxV9OlkYvhgK/vbDj/4ixPRz7asrE/
i7v6jwMcwflFM3sgds8WuiQBtv1+dYPLqcn/Ptq0iiSs3AZDLvNE1yFaXcYQD4kz
h3kFZnm93MQW2jcXr6fGsUCQoEkUFhIw+dEnnF6Nr5fUBrEke3+oCgB3feCFxC0p
Rzy7GqOnkJWyVqWKa6d+ZalGNQcdhOjNR+5hiGPU7/j6Yw1w2CgrCs+P5NF1bEiD
ZjONktbe0HnLqeE3YLA8KVMFHEqHaFqdawB8tnfwHUOWPxfoeThaTGEhrritMBj9
MMHjetd+gr8NAeMSBRllJRIT29ZbtSER9zTti1RztPSC2NHARkw+7Gds+/TEczxd
X3BSh7F4nipq/4OA6JFe+VVySX8eWNZ0SN9TaW3SF5BQKCl4YY/TsodIMs2+2mJ6
lSwhlngTK7IRgJqtnYN49TUWqPx1hvMINfK/+w9s0EI/x7tgwZF7BJpCkvGk+r+7
HWsNuqKfUQz1h6VhNWFn5xK2vjj9AxpthTqMob+h+RYBgZoeq1gktpj8MCk3l8+G
7/hE5vYSaSw57eayLT+wCVfzw2O7i+3q75xChBljcbodcqWdna2mZM+dnqXOKAqW
4EyKhbJ++ivuq5NJXEbxMYomU2Ag+NurkMx/Dhz9uKp4RTRKoRDAO5dBI9kaDfrX
y01LaIyd407CmZXhWWeUuSIehn/ghDPF/FdoHurbwlRaHJGm6+ZkDoC5X/AMroSU
DnEKyF4lj7fJYPUKHRmbFUjje89EcgyOXQg/o6SuuICzg2AJjTlu+3uUzCj0evsh
85dQzj6EYWO71ynt1K2zmqk7v40GNV8P93wAYtJveeSEbpD/y3y6+zz5vs+MHjuQ
53zlDHlkQHyB0YulzaRfqdE+ZonbWUCtU72BiwfE7KBwPa0qCneX7k3NvHp2Aiwd
5mmw//gzqaPJRwazjOOLMobhOEX5+FnBEZW2MuC0+RncvuAVqrwf2Xyn6FikxHO0
R6EpaVv+vfvYDXNFEgZQMpGBkxc11ptbJOvBp83AnOfD/3qArlski22PgqCr+ymB
qEIWRIHCjqecVrs1FLOiUCWJzxKKNYs0Ce7Qi3xYPbuOSvyQ/LQP0pIt9YaKD0Ho
yf984DOrFBdhDSkP4k3R5cAeQQzk1Ue4UxaM0NfUQirOBT+Yx+T/DZuT1jzWMEug
u1BfPgxR/sj1Noj/CDBMXqNeBQL7njuuDzOFkHpBdJwcdfIt0Xx/ewQ+KF0XPc4p
IL6mXthdTh1JrfbsWYVCRL84cLXSOCmK/bgjmlO8kwAoqGosi0I2mxqEJr2YORlf
X7qSURnrQ5FdeftqYDir3cOXtM60tIq+mXxMo35lkZO70GMtByofGsgaQaRnseV2
PmHKc08EGfDE9w6j0OUb8NkX9SH1JkP1tpk7hZawNSyTHvfJblCpr2FNv9PIPBZp
/MiQq5A5LN8j4SmfDjRtIAAI5pEfT2+Tuc4lcN3d+Zxy7HOMn/wRfpyZan//xr2d
/L2JD2pS+zcSiZjIA8X9CQmbTxM4DeXE31ANI5Jjvv5zPy7MKYKd2m6TPWlqatfn
Q/wyeu8Pwo7bNDJYPPbMjS+sMukIUwmOzfqYDdLfNtw4UNAbHAiwDRqWnuuLQwS2
TLAm9B7i9GX/c373+liIkQK2HKDovUZggwyynNx9xK7dymGTpue9NfiM5274pVhA
mQeTmVinHybTUxSbHe5T+GwwhidfZDS2eJyky31gHkJ3v9GxjZmtrFVF0CQfZ9RW
mcOBgnWfRR8Iz2Y6c1QrOIJnVWb0XOdA7nOrr7GJHA4VLxBtM88y3Vmaut0eAeis
j/vxIonqZUWryu826pZVJo7QJYuBZWguSGprN4Oc9mmIsAca1ZrT5XAvD+Gn56il
1M5TUds8YOlb8M9CbgbJx7+rN9T9UtAedh5Xyevo7JULxNRBM+MTpmH7PHDYrg69
cRc0fKIU2vbGKRtOtQMBHv+acNYKE+/BhUCpUjhXEamCqWRbzauG/bVMEF5vHUHE
wFgMoHNhtb8WDIQ8zXwTT6aRI9Wg+UMjuKC8JN/7qaUyrq7x5GFY91vt0QNdoWaM
tx0S0b2AS10qdkvqwhYz5GQ2bgrdkHIGDIi+6/56m3xOVeGLzorbbT6/hbNd+Xm+
ebEv0jjJ0UbzH4UlMCwUcGW0TRuhih2HUa/iHu3tWWrORWNUBCyQMvz1tIq/jjJG
DO1Fvhex1pYD3G+Ex2QhKf7HHLvxJenWLOrFO/DYfBbzvsrcV+cEzD6HCC4LnjfB
fih0s0/1yT2c9DJ9XZ3skFeIMxp06jcE8esGZ+LIc5B/3W5PWiOqhjfD6XYlXe84
8nohtuyhS+kSXnXU78452r/2h2gb1HJ9/o5X2Vaq/JVFNtsFLe7NsAet6s0CbBFg
HdRY58MPFRPdi89i33l0V8Vu47kfYqFxrnmUDZaY85kBZD74TFYVzefofqUMDA4q
4PeiddwRplB6A6FKZGXio4WxFmLR0zPrugeJWj3msc/PeTWXon8XMX9/O5xSaJ3A
sqnoOYHmfz3oTN93phLnms68dx4yz8XiE5sDOY4j301CUYZ4uvxPN4RqZnmEXyRQ
UH/9Sfp6MV1bFG+tzJNYWq0tFQLbdNHjZbI/fqpaBQrw6dyLoD8kpXb+axCVg2+C
y77Nn8XayRz+nHcc+9aIlfzAQ775hw8tnMn9KGn6f3XB/IVg3P8v5WDXzZG2S4DZ
HJsS9bDMvI4Utwnta5Q9P5Z0VjeDNaqKpgDCzXdOgoZYX3pvb0fJeoy+oU/dd9a3
3KdgCDcPgIUGVV0EW5+PR5CpytXdshFoRQQty7Ku+W5/c6WVKJCgJBPnso1GvPiO
mChJX0T1jibPOu4EUhU5647UZ9KxWk5lSThVx+AbXdiSDUogVBXmc7hG3jYiaD3i
ygNBEOTtBTlK9jqm2WAVbqWOYr/UfHBlerGF0UwMlLNrgGmGEfMDFxLxjFcbLfod
YNU87uZA997a2hUuZK0j9vC0DvtaBnFJuewpku0QkMo6yAFRGNHNFuUCj0EAvBzJ
c+H1Tytwm+GjJQFWQKEtmb1L978n+yO3eufsj/cYvHfLIdTcDQbyXPnyB/vyGWj4
KtzK4RAhqjrj4K9UqdsYz2yOTrTCRDzgqI66LXbO6AK3ECiDe3vsjjX5el4EpqDO
7fxsCEM8zd50TScJ8aXl3k2xsWVP+NU3jisC5gUHy/hmzJ78XFskO7y4sl9AEGNM
Kat2BnFI6khvRiGfu19CB7PgFs0G8rh8ktH3dY9Auc65/P8+3l6m2EwvElEMho2E
1WkdKzUZU9Syk1L+huggX9PCLFfk4nZASPNfZEmn1cLzUak9lqQbS4hyqhu7eWtB
PCgHNo617hgeuvWWJUvkssnuYXH/Rnhzibzcat4F1UzPlGg9/eGHB8HIRBj6boKY
url/iC7lFs7GgBQjCiN9CwZ6i75wy6oUyvddSboavAti9Y3WOZw1XzT9uV3JOtSd
GqMd+qwjT5q1WUKzPOxbPe+3SHxc0HpTpmgODiZqrYEYPKOLgkdsbB4IWez6YoPE
wculFLNpUFPciEX/qrFDKmKy3v+ZaT0GTFr551zS9scBs1coAwEE2/WZnS05gYWU
M9VqhNEgsHMCQihrlFbrb8xiCaM5e/KVNqELXOxU/9OQsJuz8nk4NdOzv3VKw+dK
zh0nLWIUz1GOIg2Dq2XY19XUsL4g+iCvq9tvCUciSvPykNb0DJPBH9AxXLO/W5/l
XOzS7RW/oRm0T38qcXKLpHe+31TUmY1pSjp/NVln2De+hBc31D0GXxxi6ScmDsrz
RQ5VcyaR2zfQOkZg48ZO+W1QpknBOMcQ77TQTna63yHET38HmYLRry3V4OppthZG
2sgRuDbZUNyF1O7w7m0UYFI4yeVjzaoL28ZRCoIxso+35j9yAilDGxDiqtwJd0DD
OUxLN8AFi2t35otSY75heNcaXFvWQjl9qrtFUf1LQSc1LBuPl8IATm0ySp4OjXJ6
GNxEAwfAXd+qI5YQEY3HcJRFEBIyYWP8dD1soQF7gPKlCS8yz0y6F0RHgJOOqp4j
TyXlKMpw8QKrd3d4DgkHCNt+SBrTur4K1HSyTLOQYWm9kVoPKTeDTNKhS1bn/hwh
9+oixYDCS/6XT3MpiMbLX7Fv6kttxAgA8laRRyyX3dm75+lNzr/w88vLH7QxNcRr
SDrABOmmn2pe8NjkLxzn1m4tSOCZ3Bo2AcgegOju5uydfBtW0LJwQRQrI4kMhOqO
AFLu0vf+kAPzjQ0Sy9glTBJz/lTmMdQu0LIsKppTfnQHdc65Z5FsvIYly2MLVivo
uq7DUU0DljnGx6PeIf+MqSDyQZpbTEGYbIpZ0AtzrPbm5RZUEjIgwVhfKL1CEfo+
ZFillzTnjG4v9x7gN6WI5+ZSYGgt7dbnCEtC3FoPSgchdYGQi6dgoNBMqxIY1IGG
4Qah6G3ZNl6wPEfa2fS+DK9hqcu9XdIz89K985l0hJhK47RdDetX+H93ZwKJ4mY7
kOs5IlPbu1KqkWEG+FeIzIt+/FDXXhW4XrZ5WG5SaNqtCcyWPVtTHtTWyr4c4q6W
Fmb2U6ApJPgRQJGASvOyltc+XxxUwwZHbX7Cspsr2eiA2Y9fSzVffPDhi8lZ+PV/
kW+HdcVO6l7ZHPWkYSi0o5763enDr1eWplCvMBPX6mJJqeIR8Yvxv8VpImitk6nl
/SlYeix8omMqh53sCWTo0o5oeaoGV9sl2cSvb/Ov9V0RFKY+K0KN41Yzw+zCTPit
CQ4/mTphtzIdUMbKoHaX5kyIrU4YmRA9QRfS7w57mTMiX2f/gaiKSMes4conYtRf
m+XIvAeJLYgCPqlRWm9SdoUIu5cB1JoDJhSEEYJ9bBSI7Jmw/1gcXUEb2HgkHtsm
Rv2V1iJJ3isu3oWKYiDpdd2CCZEMVWC2XkM3fb/imanFYpyLLtip7pFFoHh0YLgV
as2XGbMJEWZ17QIkntqG4jxguk5fkl7/Iycn81s6jgQmooqdm9wykxGCPAPD7aBH
C4vVWMZelSP1mDValZTpYPpOxnSBpxMv1YC0JEm/FdBR4cSlboqEqbBidyBfUkBc
yeH39zZSjwETvdcA7nrbXmpemvYa5qeM63KGcLhsjQKpjSPei9PHC31ONmMZlb42
Uu/lktYuSCFP2n4txmwi9OvhRNPVofNFKar8wBASYscKp+l9VnbouvMv+e3FGVwB
zzInjtYa2kfbgt+wi1antRokBDtbNZKHNG47hL3rEOecpGbmFRy5CO0pB1HGkCcj
f/sfrIhMuEvRTdws8bZxenCbZg+0ktSGosIud6xHfjIBzil1F5dED7BzT1RyCgom
rRKkv+2kmFslAuX0chpSyVRK+vXf7XakyQkXh82q3PUuIpJ+cwEikM3DMG+9TcqM
SiOYFO74T935nyftnmYDq09ZSykCz9GinhkJfa6MbK6UGVbzVKakYO1k1HXpepoY
B5hSMMWwbNI/I70MJ1O3vgmQ3ybYyVZHKxOAosst3vAHzzlKGe9G7IjIZdMwzPeu
3AtEUT5ewcoWkVE4aMaMimodyeWNC1zZXQj1Da8BjyQ9TBc+pdg/HDOcX0XMqPTp
32RRlp0PktQOlCuAZDhRGBw4VS+bwq6SE20MPIjcGhovKQdgm9pcd8paiRMLrpYD
JChVklN7PAEvP06yLJy6dlz16Gp9vwyraX5h5UzPKPpeD8j/vkwLe8Ccpxx3uSPX
ascyztvsvuB0g0P17kFrl2o43FYDTnNpppE9vJLNOvXiH8Kf84+W7Msg2IjD70N/
TPd/D0UT0aMLBzYFUbvK1mBfY1zlR2vsLbWoIAQY/n37i0ZeAiA0JgxV34m2AwaU
sDAqcStC+XnllSZhYzggOkTjB5r0uEYMChGGX6jESSzP99B5sGzTv8ZX8NmEeJxM
htfDeend20eQHFDf6Px8yTa8IOkC83evmv0IrPH2gFHYYCxYmCJbGHmyWTVpLcxO
A2fRBpvyNRq5RIBSgfS8XE7bWGt9+ldQDhm2tdE5zwz6x+55Nu32spxInI/lDAGp
A9fTFb5/ELt/UhiY872+N6i47qCgq11ELIl/hkdfGlhMIsMd4g923SmSR1Dcd4xw
HPkZTB5Pw3vJqKEWJeHDAelXjUe8SS3p93fa5MUG1dg+LFyf0MEHTFRtVY/ZO+yu
16bPx3e0UcwwnYNETFXUSNLURQSFAronAhwrIitjjysvZyC5luuUnRGPHCIDmBAp
zReYXnrpLwsr4BLKIEF48ypDSDeZjFb9IL+6mEVhLU6SrcFlNeICnsXZfU0Qj3mz
faEgudVT2uv22GyNOTr/mCglTNHryr2m2uGirvPJcpUq1HHbS6zZFl6acG+xVpiN
3O3i3aMVx4/xxu7aCgNFqDQK2MUtEkCdd+3nNgAo0svnjwPxSiBnu62fvh8Q55Kn
9i2jJEGc8Kup0UjRda29sAsr6GWub5xrspXkuafO1fusjK8czOay8minOx3Omb9l
e7l4Ckd6zK9UVeQNj2bAOOhWivLiwRoAnHZnO73TOU6Mp8l98847aEXV01dpbQWM
Oyo0uz6XlHqgMKv7zeV/HlJirkWGA2mN3eiK1dCZnkAELweKR0SARAP7yR3xOdxG
DdTst9sbrf/jeJZweh/UZUpO2xuLjGBmW+hjJ3BnlF3GlFL1n72hNxgv73koxDY/
vv2E9H4pUwaQYYuYPSvtX9NPqso+3KutLhCiXJcY+j+phG4TkgYxk6v3uQ9YkVXx
YUg2JqY6hIxRXty7Gbi0BbURSO/Gen5AU0YL7dtKrUnX+dIOQOPs9JCx22TBXHhO
DdBzUxmtnCgz9ofG07Qq4C/k/G0+Jp1KWFj3grlxBevabvVEM3bEQq8QVjYntDet
AzIwPyBVyZebl1aXFXs7wQ58shaLMFdCXpQr9AUTmYHjhSImog5cACtd+wl2Nwv8
f74/9S6RimbBzeMY932DmlJqJ6O2I5QN7UBydPsdW58wbDSS93WAMtmM1eqxB6MS
lhCv30szceL3N0Vy9L6xD/pP2n8G9C8w3xlEAwhyyyew7Z+AxkXFhCZ+hn1ULVdT
1Un8KeVLzZVWiyuHTopAdLfTOGxZWFaEbfXztyoK7u8tIbIx8zKuFnVnYAtD2amF
Z83gyGOmOcoXv51d2/v3pQO2SBkaZAep9kpuC14dZW8uboz+WxXvTnA2oi8hmFvw
BYWlwcZXqRMhReU1RCsg7F5bnFSmjgfYqDsVfII1mehBMYmsdRRdyphEDHC1KGRP
iyhmRHB92KBKZdkddlwN8oFlnThUVGcYv4ldNLtyOhEXHZTGHCKtmPWjVnxoe25C
Dpn6LxDPMLNNqXh2bWibY2IUeHU5ZoT0rx8Rt8spD5j0BQld32a8pYWoFBPOm+UM
r8sGUCtG+QKCdnLvvkivZZhB+5UMbaFiGo2XBBinSPZCGgqn+KEXcnuS7IWYXPBW
L4i6U11gwlxVySqvB+ho7DzWH4hs0bhZindW6mxDr6pkfx0OZtVb8JVEEsHDM2Dr
UY3/RlZyAZBU63v8aaMSaOVOes/WlB3xV8clqVSSvl/Q7qldmyUas5Ye7VuK45pV
M7Jz56BJV7FUkcvZS8W4BRfyVoKNQdPow+4ag5AWjyIhcIBPdb+yxoeDMeGZY+iB
bfiJdvBHaX4BM8OzX6nd1UU+ReOVLMikuqaheyFmG8bhZ37EA8ie/UiH/c1dY9nD
G3PNyYl6kQnG/1sAp+AoEIRZj1MT+0KamePKKAn8qIz3f86BW8c99igUJo5uow8r
idlFIXHPQiuhqgjztC7b3h5oZAT8LhsoJRKIAsQ5FU8Fojz4RvoRx3XszBCp9Jkq
JVLa8+v+Zu5v0ky7K5HZzujPgj4xG0nbfMhgzw2Gct/M/upF4KMFgm2uec61elPa
Y0D+kKVTxZXBSPE+9ji6q+NnTYD4BsvwE/aXEVQeLAgmaCrmH1M6JriHTdylEKf9
iV8aD1BKGOIbuQBB4NbsoCcUTerGnSZ1fHUCWl12wfALrsnjSTVwjqHX5Wp28lho
+iE9Qb4M8zErxbxL2VhoA+ENj3dbsyh4kp4hRwgupHJbPgMuX8MsKrF+bYDvZUWL
iUJ0pJahaDGwNhnXZcfw3PDKtv/PdJKkHuaWeXqQrA48yvLAsJSZsp0tQZvUIGSW
JJW++sAxtxVWKGqeOkpnlmZzJGBPnh0v6YWQ+xo9JnIMLOYt+gcm53hmESdb/rHD
VkJOzzomoX0ut1J6cUuhj+RZPXdYtjXrrYjRWkkfjpL49SAG6ihPutuj0iWL4ZdI
9w9E9oDBF34F+rUcoWOc0ukUjRPKANTPj+ltXeRirmWg2tWiI3BHQVVgsIJM1Cq5
+TJAXmTSBj3md9MkqPX3GWRemULx76fPvIOLJS68SI0MQQ/gQ0yliklOLH0hmZN0
YtTYcR0xRj5y39TIuezHSNZWS9niD1azYwvekqLjoRCy+PZ+Z37fM/WVZXnAkIhl
N8c782SSh6HK+9RjCHSUvq11LGhPYC6JX3vep8f/dDlOdsZos4iSwva61L6v5f4f
91qfrwQ2/PjOWCjb5Tx0ESGj56YV9AfBk+dfQxl/IRARpzFVyJj8GuGXvQdvwqXP
xH4C9wT2kf9Msq7IUrM1UqZcPatrxo+4e7f1KUivTW0BQcxBUBHVonfbSVrop2lt
/FsGTEPzMXTqOZB3YMMZ+smdXVsAl2c6Tee/wvR6IeYwl+DNbwejjPiQx7jXKGck
XxXqQGdxdJNEC2X96nY0NA8ZJGaiHxXEaLzjOIu00jIddXp4a8BCR7bnvd9H2rxT
BEMInbc3ljDDKnN5sIx4rPmAsFm5Bf3g9pqLGTpgNIgQ8o63EprKzYuM5ccsZL9Z
AFDNlaewf0s9MoZ7y1rypaZ2uyiWOQIRKeYHCFAGj7thekWz7w2XZdMAg2PDl2JT
F+NMLKMzyuEw4Jy/hY56KQZkouB4ospkm+nN4azyq3cv3Xsi6uWkHvametGgMThW
xqP1E8wSsN2CpHljV4xxZf/nxD1OD+krHylaTvNcHXF8XvHHbttDsT+qamp0CENz
8TlEx8P999Bkxcx0I27QxwSanLb6ZoXBU3DQCUmEq/flWZ3m0eWaREM7Np+09Iwv
RkXiqM6rFEu3NZwZrOevb54ObbTlTOUTG54KQTAgQLCQipZ0wPsuqi9wN9omkzs3
ygYrZd/1A3Av445uaRS4NPBEUJuKmHf9Dmwtv1iCv/oDD+xmOniJSByivFycRIsJ
YRSVkygUa3FCn3KMFzKbFDRaAC3vqB7sugsADFjHAOJ6ZULX3GJ7TQJ9KSD0VwyM
kjSVYDvGn40w+eZ15bYKHJAyqq0dtOlFV3u6QOsGJ4Ih7ME6JUr27HYuv23NrSz4
XnLEImdNsp1vCqpWtPRQwSLhfq8kzJzdmFfeMJnRFBSqjM8pdoyW8vxtThgmaxfE
l59Sz2Z29k+tGo/Ry6fu6plz19TyimEf1H3NGK4PvkG0URCa/wDFQ16cA0Ex3bpx
V4ppKRI5PCdLCtDaOFc6XJU1bTFsqtWJUN8gqrblAbkPK54DNGPLq4vyGtNOJxYP
mueVsbdm1254SH6vI8gu21uUxMOYNC7mcH9SbX5E8wwoT//ybxU842FInl8pamDT
lGp7yFTJ3s/KlywraFX3BWLdlJV9A9Qfbnv9rkTBI6wrAyKFjL2Wgy0t3eYnKd8T
4ybLgSzeU6OS0kpc9EJK3xJtuUwQNnhExjhkIWdwVtotu4VT7r5adqp/Ir4T2Z3A
pezyuhRpl+ZvM+7RvkpaCU0/+RFdfObRIHBkyz8ax7j0VuzbKuniQWZsh7sZJLSD
kV8mEJhZnwmi0qRnegT8Ro0+9YEUBO9Julqn9VFZsJZ40POwTcCBWCR/vp9iKxhj
47Xmpw8GnhKjn1N95ymJ7E1O6NSu7iAGvEeGKC5A0Vh2FrRme7c/jy2Pp3GTM9Hg
MSXxjWakPXO0guvxpNF4AxKEP9h1Qy7Q+0wzV+4Q/xk7mN320Sq3j/wM8Ax8uMBC
wCLYiWxovGz4lHPvJW47386k+HjSf4H//FAVInpSQy3iGe/xOxdck+hc5FMtwtLB
YnxP+3XLRmtG1GxFCiiZB9z+XHbvQXMN5ss2P3u0Xhk7KkiULeUZlBVof61G9DAN
asqZeH0Lr3NIvqBLr2k2wFC9hXox3912v8D+9SDkfuU3HltSeU92LMyBjUrsLyyb
v6yuv14ZKdRwE1r3O95zfhb6molzwyTvMvyyG+0Re+5NIscdCUqasmpGScNMaJH7
A0QnE5si1iB3FddGPN2A1TWiOXTeu45DpSJmy+GNo5HR08jBrxsHAke6vjJj19+H
9fPdT9x0ke7UwzAG4nubvugd4F11NjLjA0G28TyyL8FL3BDTVhyNICl30E+dJhMv
TNoikDckB3v26ajWTebxnpuM2R3wj8ZoJAYmESinKk5rM6piXrf0NkzL+hjDa2jo
O+ijcWQF7pdsReuif7QJzXJb+Yr1vpXpPA5cd1XtdyNwpsim2kzLoiHkDPNK+gyU
06i/r26SfLbu4GZZeoYO87MYsHUzR6ReUQcIvdhrOuQvwGs2sIA2KHIfTj0rkVS5
RRwVJJeKrBxuZ9JaK/umWVH9wjnLieW7rLR5EWkFUpX1arwdbaToMf0WTCFrP/B9
bXkWOGy+jBINPbjLmrxvO6S0doXyI8y0eE+dkt/PQdJRfKA/jN+24/WQFHdxRziU
va5Ngkpbw0dPq/qlI47zCBcXi+Bdq5P4aS1AK/EcLVyixNDfSlnXq/pMf6N8cank
Lxhhuwy5H5/Bp0P+RdwYGsOvE48s0UE4zImm49IcJ++41dtrJaIWCEYBu8hPEWmw
bTQQRaqih3OI/XPL4I8Ty/dssYQfKRS6sdR+DGT43J47UpcMxPatOx+DQNgG0eyU
7J6sBS6KmdBJBYunRMFtP08PdghObUKFBqsBF8iuxXNZae4qOgRT9YAmf0SsY5CF
B1dNe13HWdPY8ZnaQ9l8YDQjvz62KlklPGcvFfE+c17ToQ1rr4ujU/odIB+aihzM
sSEfaQim0sj1/vrjVKwHvKtnfmW1I56aUhxap9TjWEKVYu/0RJ0VEm2oxsaUhHOD
Xn68XV/8q0Um50K6CRzZ9MCxBdheDar0jLMMznZXtGBPnpUjJfucGsIaORLMaL05
pAEcADPn2XlqoKR4KkfxY+ia/RUazlzTjWL5FRQj7jGjVyVcpgYUFEb39BUH3YmT
OenD1gg+MPitM2PxM7MD+vUZ05biw0TPUeaJiYvQ0EJvBWFhVP4gUFRFURX2en7p
ocNR4rh4oAfBFq5vBIGiFN50nVxFVok869/w8V4VQgVsOJ83zABFfbuD51hCZ0ZR
6u2sOvLQDNeXvzCHzsAhUzGmnB8+/ivZAhqTcsd2Um9DH/8pL0h5vL4tMqt9zkK/
IdprVIeqtOgpPN+RCj/vQKIY6gQZacgCHpbaUM/XZ+dAsAvqwEoj8Ug1xe14tGyJ
MzkypwjiFAVzSo5CFU9FxeFIjLnORk2FGadQMYRGu2yEc9jrhifsYMqRsvmclCU7
N9U5Zfo/VZV+ACUMMTBLqTHZbxfhIagowvYviEcI3YPnbni1PHGUEC6ALChLaVkH
XxlhvsTIy8VbWNg8K/8vxSfyBxRGx/0f+o9H8JUvWcmTxs+oKyLi6QuLy9NbZmPP
zRX6IUZr+Ijd/ttlz9hmzuj1k13pPexHE3sBTnUyZE4d9PAVzajJBGQU0BocnpuW
jAH+XKddWCJTcTwAY7mNBf9DL6RjOZfT3MHF3ZUBQCWVxbOKyfaP/9Y/abN+joar
1CI7DTmnwxjVyLFkbX7xIPniGRlNCx9IJnAGWxzRJTwDpXg9ifpSSHO9/5YfBAj6
LSSvfTeyvUcKSjbChOiCIL/NQwVFBGLCUiN/D5xDOcFYrAkAXIxoL7+kKzNagzUF
doZO/FmO4brUOQ+DyF8GnQuokaBEQCFZSrcp0Zsc8NE+a9B42JsdktllSr149PUq
oimu7YASV1l+mj3EWcDOZ22u6bWyRg0Y9wqbOoRUNkjhoEOs2prjEI4l0kTKd/YT
flO+oL39jW9rgBQ80rrcwsBI/xOKZgPc8f17kD+H2py7YcyPTONLpBGNjO8esIJ6
KZv8SxS1OsXM5n7Q7EOhwbZXGjlsM8pSoq3bxmDUjW20WbYsaW6k3M4tcqochMKt
oJHM/ZQaAeD94VLeTa8F2x4Q1lFcEn27w//aFrY3WcmGmFDBU56SeeA3DtafCb7t
RbQvE24Tf9g7WEq0Ux9Ab1DcJobSItqVn4xzWYgjkXGUgvtE7DWOjcYwY+AS4Yn4
YXHQ4uYkaj+vBu7m7z3l9ASB6+ERkX5wycziBAhWca71d/vHp8GKMXRGGyzHKl+C
zZr45W528tFwkb2Bddt/spfgy7vHrFjb7wjuRnRp9DeyhxiYbf7+6Fiu+vZ+XQqp
zEKEZp6ocNDxQvFJGlo4Vy33f+LMPLOF+fTZPTx7GOc+E8GEc4KuxYudgxfIQP4h
BpkmLXh7mcDC94Sx8vUG24oak4aIkAk5hPKMsnEYWCAY1H+Qz13qCyJlTz+00TGE
+XHC8xiF2Sf9yhpjw9NFt63nNS9BNQ0ag/MQKTn3Ff6xB4oBklRX5W/3HfdV0159
eIUom3qn/N79jUBbcX7M8mRjHkyqWZDYpanTe2Ba+4auXsrwmpX7xqIOPlVpUKUd
egg9v1+lVk0j8KaUKF4d2Zr4S+IRjfxnvSkSjTYclAB/GZNLtXOi/Vx1ZIYvsi95
a4xlmSv5NU7HvjhR8TzFKhSxZUKmfKV46mcq9WM47E/olFFGK45IXBYvLMhJ6XPw
jw5ojM//ax48nE8jZ9n8j1g+xMaEAL86M+23pWzqvyVdV0HaBjBXTxymCYqy49E4
EvO+ux4Drxhfz+huvgw2ViTh2pO2R0oL/aReOwhR9oqLBC1QzazXOlGKm+Cq7tPF
OwrJ85dK/S3LeUkIOjPJ21WMrh4Rd5OlfX8XndYmHhoj6YKjA1PcPGWgCxvLzNaE
7+Cb3AUen2u5lJxNZ8AAbPOabhdFtmjwz1hciplhjRx8s4JU0nvQrtA+Ax6ntY0b
sYXgPmr7ked9vsl0e0uzWDpNChqfLbuFWHhGmcwJ8mzu4zQ8gZkDs8HF9vVhHSDR
W2Fx5qPKsYXBchpy/u0lXbg3vJpFsiVIXY1zMieY6vKqR8RKhqzyBmQKLeEAh9ug
NSA3ONtNHVGiDtaRKWR0JQhT7HSTH46gmaOMhAKwDszbq6rVrgOuzaAZ0GbGctKC
KXmjsqfHr/1ydGrrpG7S7S3cFTvJd64dBvch+PkeEcF7LopE/5LYusc9+FIf/afk
DD3OPCdejaYoM6O5o7SVQ2Z5Mojs3JfCXZY7AavfqbKuAg/j+luo1kA+s+S3c7GT
jWJ+74BiPJy6K5CA1FsLDCO1DMSWofOLIVsX8b3M9SDX9MW8fHavRZZrXE+liA0R
vo1d+WqnmiEwIYW27EZSatl2QLdSHxuwrWYyRdTU6SwNoH8zSW0EV3/UMrcT3GBN
IG9JXNF05Rsrs2bz81I0c4GcMCVM6E29gO8z617egyZXRnJnhhhR1NvkBFu7yfjH
8TVzU3H2KrQBhKf3ytg1gM4DXUcwUZbe7jhEpfsa/sTEgpBnYMmDEwv2Ik9TUGjM
nequiaPSoZYbaVSsi1OPW88u5zDvWt792foNm5q+87qNp5Y7ykjXDrxZwxuQYUKI
a+TKCLqMD95PHMgvU1fpDqOMubLFtF1O1eB/5FJBRpY7kyq6dZYUpn1L9la4DZIA
nOubXAs522zDFIPbIOF9eugm/U4amE/aprxiEJczjIzPBlOWoG8+dnFT6e94nrk8
0BYgfp9bGhkXWd9GZaREIuGM+X072up72IVDbOi4QDfS9/2MPHIu55YioirPgTUE
/8Ib2cpHXIon+u72puay927KMhHbzqHLSIKsG8734jhPBfWcUexxLTYHUTaXcpMT
uWXds+DiKHkxExiPhra5n2qQhIbIn5vxMw3Fp6E6ii3JR2QpSTtESQjfkX+MHMcH
WGivvxvKHBoHcioEpkRoQUS7M+ApjL5KBG5hWyeL9CyxkdxXYH1zzBGM96vXW0at
x85MwSvbjajw2/wi6/+kVyGHtMUyJ6V6m78suVCv2ybrkq/DBrtIjYvSHqv3eoWx
mLTOB8UoT92tiB+Rx5v3BHT1AltEYb/1nUre9N9Zs8hd/cTFp7JVuNRLRVUAUDGi
dGVHvRoW7hu+woMvDKEHZzTRDepMjGiglJEQ7c7zLazW85tH2IXBGPn/h3FREtO8
rbnxOEuKL4tU9YigxjiFl7WWou3slwXq6LQxebYrjLxVPBTsamj55zMA3U68AhTB
Gm0/SXXG6RpKDlRnwhwiU5IeOPVwyBDw0oHa1uRPsqEsmX9rNNvsTtu1wlnN1jtl
+/uBZZQv9Ii0BH0vSBClg9ogjR3L0e8rvpkRtvOKEMG1aZ5dgQcOLTpmtUhMqpUa
JVHGA2hYzfQUdSY0YyVM2c9gyDUnTqxI/y3OwWrS72aqcg3lhbGnjd+S8KhXJ6TJ
MH9Nf7anvEHr14bfRB3BNYWq/SOnJBbGn21qMFdPsKWRtKWwcJE0JMeIyiC06+cs
Ew6gMnBxMOoW2xloUW8Of0DFvEiUQRp3WvMD/IA/YqTpEiZyvP/jpDLo0dqu7KqF
qUp5DCxlHX+faXByBWr2G7Z1DDfQ8tb1w2WvFyjg5y/sJIdjyv6aR2qCG/00uWRJ
L1Srz7DsZFId4GOFgBV2zRnHbAp3rvc4NMSroEyoPY6s8jBUtt7UAO9imYHr1q5h
5s0xSwrPzjhIw3WZelv2c+jBswQGVLwDsLQyOgJgkZEt7+YppYRxDPVWfE3R/2P1
kbQfxl3pvPc69c9nTfPKgAm7RHI19g0JufwlKygZgecNsYd0z+jnNTLQvf53zR7D
NtHmY0zkS+yW0rb9KSaGBFgHHFgGN2rKg9lBqLY83rOCTYK+YUcuK/CeWjuUlsOE
D6XYbjIFbEDfdvSh7TKmNfiVuUL3CRvC6sEgJhmJ91y9iVRI1RIYAzRnD+7Qrj9V
Y5n4gfnlDYAY/P15Sml3b7vXqG7oGRin4opOsBA4G4aZ+tlZaC7duKck8ndbpU/V
3Kcpb8xgMpEQ7vDACGtuFm6Dc60Bme8WbC3IjKZsnn96NFzQKupnT4cuyDEzlk25
KsyM+5wpYyKTT+R7uyfLRrtZuiIgpktbh0w4J/DWLTsocMHTWuniXm2sSsNQZmtY
6HzkeuLK6v57oSgKZGFCBerPTLsX6Yc3G0KmloOZU++IDM5eDeiPcTwL4lToPqAy
ZaqHJ5OmNvQxj/96J6kCknXs+BL7RxtdqnvzjaIZjJx8CAWbvYLiz/5X4UC55cLF
oxofegG8YAkNaUmhiAjlgb9uQQIOj3ARBI3M8fhQ9AagEl9hrfNzY1jDEgCiU1ql
lfgzEwJVf8sMtZ3Kqyyx2nqvR5WMw55bie467Tx+dSFWX8izTRkW4wdxLuFPpJHs
U684FoyizR1sJyoDkjpZuGxpK7ObzGTyWUZhIi9WG728QiLJxZCt9On3uVq7b1QT
u2KUiuzIjb7PTOcFX0ZtiFXypPaYK/6/1IBuU/NC2DSixDd+mlXXpB2cn0Wdpvmw
FDXBrd5tC0UNx2JzLMPyXW4AAxKEEJZs31id76QZhZ2wbIe4wJ5Xc4pUK7v0K4FZ
0UwEF6TTZx7iK4+3vtOY8rCO+j9O6QdZIP2zodBJAEQGe5Bk2asx2oI0M6VJkXGm
JuydJlXifu3PcdFZeIa81vJo2AeIrQQkRnCG1LHp0/2IsdMYbT9UzLxmJg10lete
RsgSmXBVS+JQ6up7oxI8AcUpjPq1QfFfF+O4zoPn7m2E/CBym2aj1j4VQnIHysbM
AweTeD7E5DghDyM6RoZWBDfzWjjxMHe/OL0RlIcDOfs4ORZdmGJbJaWiXM0tg5IN
rX1OK0kr/roXyQPneDTNWlOOLa26ywFsnpGhMZCahB0WOU6m7Ua+ufZEFr4+4tbe
+dNuCcDMWKgqwY1oCRpSGKX0O4EXzwfZ3EU8ovFH7H8v6V1ovYNFVwSLkdi7E4VL
Wn3UnizgPrwL2b1KQElZxfhVFF4bZ8cWVeLkjeK1fXk159eFVa70y4JFzbgnu7Az
UDuPLpGF6OiHwrQ6uGmN/cvxzFoQ/HBuU9EED2Q6+WhEsSM5q3Sng/axFMSsJ+rg
wpLJJFx8euZbSWrP4BEtLmK+cQjab2+vz4HGx5BHt52f/1MPsfAWE4zNzNNGI/jQ
xJLv7Ck5Piemj3foz4nBm8aRpIQc/Yg/Gv3kZct0vXiyS7NDSMZ5j4awSl5Vq7iK
J4+0vTJJX29twyjAO6COI3H/aWpUc71DFn5PDH9tRrpNjfFSWkLxbRn841DxkFL6
ruHZ7Wp3s6ZFJlypditI+lPWmNIlD9XeY3mOHlop7aSh+3xlhfSXiA5L9Bk54I7V
m9fMQ0AFWhNGX/saRJ46l5Czl4G1/oZBDf6OZr7xodAnO7Z83Zdx2AsyBFRxpSiO
p2aiflat7vDWt3Hy3H4gRPzjh6eGy8gyP1f+oV+iD0uJ9ZbeObUyWPjVF7Y/6LfM
neT+scppH8Xr/HxGUrjFaqAxKY541Vfi564fqSjdOBhizKXf2r1uSnXnN6WsU5K3
yMRd2x4USZtQSZSzIlRFi/m+iawiR6RbEZJ/2y8n041T9ZMEGeXfhjDRUMO+KAid
iQ3aXi0PxDsKX+LYl+emPzWeGaLeJYAwn0uPRVOiydgkASfVUS9AYygTYklLiz/W
8A1NgMXSI2ihPuwhvchlVIOMY5/h2JARt3KFNYPSjgSBqrFITZL8cjJWmb7qw4Il
e6wfJk5qGDoUm9EkyB4GK/7XsiezEdfi+7Q1S8WOcciuTpFLr0xppUSE7eYmtujp
M2r27ZiZ+jmbnDz0vzUc1AU0AtnhBkfBxAxuNM4QeZtUpZpEEJvhMDSKBy9K1ngM
61ttdL0JqVmV+tzjIY3gwNMYfSzZyZuUUwk1CpNMCnmaLH2Rs+5vn7fvtDUiq8a4
brmB7BGqriqNIahirp2gxWidEa+RFXic/nw7koGQUYzt4N3xzoXgx808XAb1p5EO
RLJXSzVWIDtqAGau2GOBnbkBhWBTJaIZSeLdU8nEXukjSt69Lfc5uTomNmXIKFmu
h85WMZyFgGSIWJIjGdAWq8x4dAf6ND1/0kFqPgD6Zs9ZEiTRJe9k7YvFBlAIeafm
jSGC7G+9LJctfdilBW4jqqNdvTcHGa6EXZLSt08p8c3CLaiwj1RyOJYbntNtiE6i
jdaAE0hocWgG5YGPnun9NL5Tfp4zCmFHxcYNXrgF+FWHAJHANou2K+vv8iZVvczP
yCregsbajDffKvf2RIkt+V60bhLXtuv9WMxTa7cHh18JRtI/h+dHSmXpfM3qnBuH
tJqHZap6V42/4R82R1pKWAZ2FBxANhJsT4MBndos9uN0qZUjzAd8xEhhD1LuzIHW
Jer+indJ+hi0pHATM2o91brrhjBzlwO/pO60FsXMH868+ycixL0sdVZB94knPmEo
3Yrk+ardL1wxbPXt+Dbws/86HWyHdbCe2FSK/veOg658OrZxCRhRatX1VfoHU65y
Mts5aY77rtgbsZ4TlG5jD2Dt2rRKkS1mcBDM2GaKMS6hbnKW9WBzl60+rS7Mkh31
pSJTj7VxZ/YPHeuLyEH0ms9tAUcHtbweHjijb1guEYmXUjx9kW6Z3F7DePWfeHu1
nigwnT6C5mubRli+PRLuUE0zJhpdKXzQ1IkWwo9EQwlVqJJnRQ2aOd4+vbfO8iTS
rH4sLZ/atpZWL/lk3pxA+yhZQqoGoqKLDx7/uxZHJ39RGxFurO35dfun5wGFtbUE
HCWJvc/Ej7rA7lLNPXC0JfhjEguYmPCbnDQ6E97qm8vNIqfKLKNhgDc8GoEKiCz2
2zdaKWUs9BzateFZC1nqvdwBMu2+BAqe3matk7LRAOn+xabiUZ/golyD6uX3UNDs
zb4h1JJHn7d27iU4EGX1LVdWO83b3mTUiLNDHk1P5c2g/gDmdn4aU7BwYKQw8CE/
MYZMQknjcXsJ1D3/wred3HAxuKVM6tKGGgac1B5CFhUroQfkANItaVh3iNm9Ip9P
OQNMuDT9ezrbgJuJS7Q/5STmbGqmJwdOKLImMuhgaB0oyJTc1aNRhuL0zkmUQOMH
XttaJr3sdytkIBT5ykOQuFwOITdVPPyfog+zFL71cuRhAq9pjYlQPe+f2Xdnh1yf
oKtbw8twBJcJi1k56SVjkVE+0vEwZrAjdvlmDZgHo6qTLNJeVac8QKQupgTG0S2z
MmBH5uHIQAMeROYCQnkpd3LSCYmD1f/y5CbiRKMsKKHbDWgfYIhST3W2WAiG/J4C
OU3Z1OULfV86k2QzF+b9cxuMKAASoHe7WVuNRlRCdTlaisX30MRcm2vKLgzVagLz
Y3DobcI/Hm2e/UpH+fYqy/bZaf3RZX6x+uHXLAAnoPeuzN+/YIjDiC/HHeOwZlex
MnDDf3myQfss2yjZfG4wfIYM440d7asb+LBDhiSpkCAARNM/JbV2zuneHTkNW+mx
2kG7zYw2Hzlv9ViGOr6PY2s0Uo6d0L4CJiajCQxcneUXk+bWA1xuhK8iTBhNs/Hw
5ehdbDKiCp0jiryDvMTAcPYLdBIdXGP91VkfpqPPzEgCXA1LdIKQqtpxSN0CbfUJ
5bAUUWmHP1ApWrUOYPVV+9G37BmRWqxgkYNBw8lCKHvMYnzG1ah/T5cLvGk4iIu6
VUeSf9U9U8FFhXR3zcz2kZv3Nqn4cweD3++Cz5gn2Sy79xzDrSHGSV8kUIFgG9bh
BGG8nnVdZ38gs22k0hMyG4mCdxQeey0vUwXxBvssG4pINqOnCAX0jIXJtQze2O1P
ZFWrXeQck9wc2rTzJ0lcK3SU503d86bhKi8u91EGW/iaR8i1VyL9Qls92W8Jyi3a
iAu04ZXUHJ36hSYVXCIre3tveNeorOYAiaTeEy2zAnHgFSQa9SovAZ+V2jtyt+Be
jRJrybVT2p4Cj2kCy6fFnNFlXoEFuuHvrlHJeQhXGc+j0ydbxK2jf0JSylok+AMA
t2CxGDjSl9EdquKkBd6vNryeQVbvHMX9EuLB6+2hv+1WG+UxquBuk5Cy9s4id/Sx
kSj7KjzjJ61jbuv/M0LTijo6Z/d3j2mhooKLS7uGs7pe5Ct5PkTOpIwX1ns5eqiO
NVaS+Av2Uh+P444WHzcAVDh5nzMQByTNb5jDhJRp2DNS9A1BSE/IBwlcwv6KPaFJ
rUp+R9LvVjIUGkgrHMjxl0hU+8dC/w4hJ5YnZfL0uQI+zRlZXT6kRhtO43zA+yxp
Du+NPBUJK+nkNfG9qJjbuEqdIqak+/nADLRWne4l92s6/1IOpznJ6SeH7zP//aGJ
Qm0GXIOuN6E3bvDRPNgF8dk3lkQBObHD0HEqoxNswErWhvctutvHXI4jhBtdTm7j
/5eHw5MZbkC+CS9xrVcpLSmpn/N0L6y4wAlfAYW1bqLFLTr0vQ2Oyvq57LnaVMyM
M9SNrr9AbE6hA8iEpm2uuzrulgQmez2rdxrWVswxBJ/gE/VneKYIkXg3/UNOP1lc
6KJL63W08LhF1WhPVK4YL/Kh3y12c4RWivhE4p4BfuzAWWKhLyarbyhcwSvWq6Yr
XNLvSZA5vV0QFrW7qoqOm6GTptYysypo7nQ5pLNKC3EYQgpeb0Or+mTTlpPs7y/f
62q3RbLwRehxdNbl+g7Yizd8A4/RH1z4tduUBephPeu4PrQtuh2uFQUMuPEEYmKq
6n0EYBJFh1qXLW0RAL99GWpgPIC3ueOFbklqeqSiw9zr6Y6SqTuFt58O59+IgNri
Y7QxAlXwmDoNeII3kFOysKnwBt0H3yIWgUtEovb3QKBHtXK/7Z6S9moORK6ClZDN
irkF6ZKUOXoG/RCqizJ462L9Wqn9nC1zGp2oahNB2FgBx6mMrpP7Izm8EVp/LdLY
mgUywNg8xvRJRJIbxLqE1AdNGEfa3sJ3pwr+Nj25fSJkqBvVOcCgX2RMGqXQO2Yq
4SLmyTpqLb3fL8ngM7g7TIB1y8zax84Q2hRISdtsKc8+AvtJ4hJs+b81XcyTJTN7
p4eBKWLOTUPHTRq8HbkLOU0dZune0XaWHAKZYQyN6qBfvEpMdbs3JvOYRoSTMG3L
5D4Sy1fRqMFFILy33hQolDeda3fciik2tMkzSbH5RDmwdc4PadGt4Ie1Nhu+8bVN
X9q8d7XTwILMEgMyW436fRmHVgTCDagKUL9HYRJ71bhmvM/zMPLVM1sOkV7leSfO
CFxW7XbHIOhLNFWNbWkJj/JdiYeq+lAdK95ZoEnJyOuJ6hQkZNRF8rjJPs7ejPax
SGp04/w278Nwqk0p5C4ypeocnUyt9FVQcXdE6rZ5wCjMSvqFZjkaWTsQbUD7iNLN
fI9LlDG3qSeEQHD+FTYsdJwLYrN+xhTqqSwc6r54HNs0ZenEFQONcDREw61Ata7p
xlgonCsKxjUNbCPI4c8dhMVdSX2Z4XtRjmRVyx/E/Ejh6N7WE/88KZBEb+FVI5wV
sDoZw0UaUFsWYD3sWCEHgDKj0jRRiQ1UGWAzcH9CPqjQ2cxtl5W3mi18pYBucXLI
t6br4AzLsxPwd7gB/ZhatOgQj+28jfhc0sb/bc6+amMhdm576fFST9nzy2og21Af
hx+W7ElYduhuQUdB+EsMydk3ICKLVfgFBjL1PpfEjkEWBFhnoMH7JRhuFBeb6ySV
J7+G4RdBWYX6VyRPZtuPsDO9GBEe8VQPIzZ8UDhZcrftvB/PSiYMY3dhrvre32TJ
NpKF7eWbx0ZdISMOCt5+Q12sVkue2T0RbMS9g/CJAcdpzk+W2VeVFNc/F0PHkRb3
GAi2DoZQh5bBldAAYGIYsjXDBs1kXDx9kLYcl3yWnlm0DGXO8WRbvJLwgccUx+uQ
sCBVmkktDkZnjaIINGGPoL+c1n3UsgsqHj9QxG0DY7V4VE3kHqec/UMtl+jKLFHo
ShzN+zUuvErgzQB658ZAkKgQs9nh9b1lvYJn2wsOxx/2H/lQltQtlWHgmQvsDgxv
4WEksPFqmy1w3QK58zeLA2f6PEKgRRUNm62EsEf8mIsXnj2Xyep4zzR686OHSrZj
0rEuGzV2DB0aucTvEC4yJY8E3Wf/LybjiqdAqytxhMi8LgqykiX6cBR1sez3I3Ok
Qncf52qaf2+vbb9N8OMcoXeJYc2DAt9reqbMAx+N6uI6LwpvPkSH0AS6URaenNLl
s3eUjEziOhSDr39+QjIWDswPDir27ewrXghItBqPVjrl1nCNUmH3iIUYLZGDXzs/
/pd70vU0dfih94YgZXR+BGGp0VBbEYWwMTfTNKMdFFM0YCjAXRC8ZtaPs4/crqxE
Oe/1aAzKI4YvA7fV5QpAVY68TfaJFLW8xa3iNNzPhyfKkDj4J5kKxS3kDwOx/eMS
SCrp3da4zmckV9z/Zc8PdXihCXnVA8yBTndggEn3dzlDDy4zC1SsgKT7A5lKodG8
VVoKB7DnMapM6FxnZWausii07tL2q62b6wrQ7/X7fTUMuA2faPOh9Zol2MYbYzR3
k0YP32v4AShebo4LFHZV0SIc7w+O+Ck7Le2B8SPSvMqhfus3etTwMeNspyDsXDTR
Ssl6DfHU/pBx4BfsNw419DTncAvnSciLnafJu7H8wPx9lZO0EeR/IjuWChhMs9/a
skeWWkHkA4cfsFuCJIsM6cxvZl37AfoMVNAQov0AISqoFzVvl269jV4XlaqghR1E
u7YTamXm4i1NZX2Vx9BcNHHP6btnIRSHlkS0p6bJjgost2UClMh3FbVrB/w/LR+q
q6681wNfHw9wi55E++RjiBTqIT25WAy75v3jIFjkzzgh/5mp3C40aozgq+5VC9IS
QJXDcpZJVDt3ZVyUHVC9pGlZKeyGfByxR5HEYNnX3uwSLyd5I3eatFttDTMa/fVl
8OQd4IqExnFw48uiXj7VnIhjych2Bo+wz0MHDrQTmmAZLI22T17uNxadE2ThKcXF
7RgpqOUADIaM0xbBJs6TRmVnKkW1zS/z11b1L6EUwfUpMMZblIgwBxoys71PJIQJ
e1yTWM02+HoCwdZlDQb5cjUb2bIajW2q6pA1vj78M93N5AElPDwKgUr1OYRtkD7o
DmOCb0C6SAz4LYhYvzltxq+dNBdpljPRP1WC3iu712nidlsSQrUOz0SXDm/g58oF
DSQW4XR1Dgew7b0oV3JZ5FJ5MkhkbBraJzjPbQxrSnbemkqMXcLAKoMxboz3ywBQ
pBYx6vtdYFXgfMCnhUYH8kKaDDjphjnqwR80hd7owBM1iydwVY/N3BwFPxtL+wDh
UvUyELw54EamaVPdB932fpM5/Hull2Tu5naRxAbGYtvVHMsh1pTlLdYWfhpYYl5L
+FddcQLMv4DgRpqAs221+jTuFLEFSwJhQqTqPa7EP/yvO9c2dvzFkAiOI5WmmfYQ
BDkalQGeU0KqtHpme+rO8roES5nrOutJur5qU2Y/WrxeZZceT6KXCY7A1QIjAgks
Uyh1MZ9GzAremdKR5SWQSls+v+AwrG2vO1vkofNmqNPZ36laWUcaq7UHAG7+Yvyp
Ei5aa0GPiT+UqomYOAPthFPub6u/lPCTzu8YkvYQbfxs3SjJXRtbDbbaMqDa6zWY
HBGS/q5bRpw10UMy/sMRib6A5szUmARyJ0O8h/C090BrfpV/DFhQ23lFLHdQ4KFv
xGSxqVUS/kV+UNeN+zOybvhXCE8V5mXUTEwuNeuFeQVJ1w91WWgnC3EnvXs1jQAc
4MrpmCuU3DEhdpWxJVvwC0gQL2UmzCTDikzb3W8hZd6rStdGIgssbQQYIqeAhBkK
WSUZepmf/oXKg3nA84KElWH/6n0ebIE1E3FJCQArYMaO8wJWgjABQSZdk/iSPAlo
IyMvAQu8lFfUXMPi26fD9q+D1lNWFehLXTWdLrs9/YDdL6VkSX2b9BvpYZLyr6Pl
l3MMNE6yQ5dRnXM9joSwcGjnoJVx/glQDSaI4+FLj/uSlPKBlVhet87G7Tfo3upf
Y9zl5WHhihTDdm1dx0F8/fDL/o67vJrDsLQvCNcUTXch1xpoYEY3Fxw+FPiMB6x2
7Rn4J6V9ROxXfPSp9K9BTEPROAazPJN/oMEM7jtunMrwfEU8fb5JNKDjJ7X9NejW
APuFYV2ZQBF5na6E9zYx8CkuaC3UAsJvmwcIGCf/X9VLgCuJNb7MoPg7amCMn5oG
K3Eo09U7+DzQIYpkV7Ez0xt7haUWR8iM0EH1nvqlmIY/irePHPUrFbEb3GY7R91Q
2chxeXqLEZUO4rTp7pDtR9H5wLHZ6WlCc6yssB84jpID/+mlBIe+B2HEgeijoTcf
sHAmPid/u02fuGQmZPEytwfkDy83+3uLDSnpjJOVSV0KIQaDKhzAIK7lxEs0lsSq
oPSW+in+2NuGsAfEjuz9HfGxh+xZ/eseq7Y2yK57BnY997vZkFA3lVIRdaCb++99
Aamd49UlX16jN6jgBYgOEelw/NAPb/8IHnSb0EAWJGg8uUx7+5WnfQu9DLTK2PpD
1Jiv9/RhfMXes1bTd0GNa3vIfi4wO6pEwbPUWc7hDGGGK0tcKQ6l01E7bKuwqsmw
K0u/9j3ebs7lbqGus7BKcAFSYeu/FtNTCXsUvkTGsw5HNPO/iDEZtWYE9KK22nuC
+RtgKwKTG9yG6kv6Vbtdx4/4X5kvJ7zD1xKruM3DNPHa030C3adVQjxuG8R9hFHY
N7WV4KBs/5NF7/R66+oAW4E6aKnwP5nsFaQlZ6byFpr7E8uDhwteEnz9nl0yhyEa
72w67ENh2fRuQnNFNDZZPaH35yI0rY85rK0Mi9eYDeifOYYp4UlpGPUyPMAY1xp6
X1YZRNvhjgMgJByEnQW3XXiDDY+OF7Lg+ti25tWzXClbmryiVsWtDEqat2S+ldBW
pWF7k3dtNFIg3wy/oacX0U+xw1v3I/zBZQVT883mTxxsBK0tDDNhGp1QnawqGHx6
hdxerI3ECmEbV4XZj6NA+00N2ZPClxlRxv67AeabGb/RtFL4NjAP3zjney3z0W7Y
MarKIPLvoGYFdu5xPd9ErjvHFTujtZyWSHMyoatH/l3AP9sjgs6OEnXQGLP8/aAC
ovbrKKHDYtthZxQdi3VDc5toXp52/1fA83Gmtbwolm4nQYDMx4S0zR43ns9Fhacg
n+KS+vNWIiKX71RZAcor/m330p8ePlnG38BHcwwzxBwAXQVToODX4rxppw/zR60K
Nq8ROXGiWUnKLRv5IkRa1P7Ouw8XV0FrkPz/KRUUtxX9+SvBpj9qwN9ZTm4HgUFu
0eyvPxxslcF6FFTz/B3ONqo49PTg9ALpmaB9vwfcmOA56ivzt7b0798wWMJcy5Wz
pAXd7sZb26wQLIzO+uSENXCKYiRKmCSKlnGwgQ/wOqfkSxpmSgidwDo2TnokkUtg
uI9V3pZaJPBUIu4MNlZgWSLpDt+oafMIRr+/HPnt2a8zrhuQfFoVNpHyPf2xPN3k
DXx7JevSUIh38rJ6W8OWGFfo/lRz4M2tcmZpw16XxLEsk73uoxwTHGRmJ+MSzIuZ
BeHqrnLHlfHsQJDqMx5Ngl7RuhRxSpscihxFWapKG13LOsavD2s3JjBpAapmLiRd
Zvauwde33NZQnjiBsorrubq3BTXZAgPn/VGLh9gITLkbQ/kWHQoQSeCbPx+Wxtl+
KSEcZPxPuyMRyoAai+mOuF6oB/CiAhDrEGkguhIFFS8jYZ0I/nzlrH8GKjIHnRb9
4pvXPYlM5I3yOjUw3K2EGbxNJXOBrl2ymdXSqDKiSL0T09q8KJtM03g1o51/tc1+
v6G6a87oufwBi7yObMvglNjQzs9KqMq/v7lGxABq+/JI+QwJrlMCbaWWvuVX3dfE
5MBEMVWtn9R//+fDx/yC1A72fGwRjkKNpP4SyS3pt1gI5lJgo5b2Pzj9u1hcCpo9
OGk9hbCnQvpQiq265zrKUWFGyAmrdYqjq+ntAnFJ5ZBG1fiPfkfByyrCv+0s4q6F
MsGzOMr4bFakdpNEJYDJ1myYZQNbyp3tkQ49T4L/3SyAjeg8PYYwMHA93xFqR1Tk
WrtWvGZx77ePV0oE2E44nt3cdrv7bLRmAfcv/35nrhvxsAq3bftVbWifIqL0clFl
mIntEqOXdaUWXln3mVzeI4GgONAJr/oRFWZi+U+7iA0f3DP4rlZrmjo8cl07R9Gf
WXl2pY6No5RsbHuPmITAcbnJPJ5nBkydX4XzGFQ1nae0JRa20E4+Ot1+d0ERoZws
XcQmBz4LJGqPV+azE7gdpNSIb76aDWb5iqSnKN7A+XiIK08OndrMMx2WW/xP0Cil
ii/sN80wU9z1McjkkDkNRxm2k1LE5WiGuNBoMPHAa+PqtQqjiB9fbx+fkauXfNpC
VP6XzpS2s0eDIrCjurbbNfouVO3Tuyx+e1M4JLbQvXJZYGDByqLpPF4n7dDp176G
vckLLBgNwO7IyAq4B7mwT7429x/IO2/LzWtA8YjQv90DvrmsnJrjq+KSQ+8x7R5X
7IAxKbn/tJRvNSLt0PgQFby7vO8IERLQ7Dy4K/pmZsIpzvp7EP9yUYMVJpmzQQle
++YnXmbbxokZtXu77IMY2653tUVvnEuFS4qARmveLV+88bVbMcLTWiqky99b94Gg
JzRJGCEyn5+AS6S/aZ+dbqAuK6REZPwpR/N2fyXAyFQjDGnuCgHlsjFZIfcm3lIl
IUH5gz71r7fGMuIzMtPXTtQNpGLWedSkF7Le9Ot4V3E6cQPPvroscubCwHR4TyJX
GSqipKxfDpNCmYjkS04q0HOJgsat7iGdnSZMxz3Z/gulzjEvUJeWXp3QK0GpGIGm
/xwLwktUeeUomc/GoT/cvpnn5enRt3TwTaTK0lffIQP7gW9Ep+I4HOvsBO+sCM43
5783kG4qWbETQkUkV4myv/pzDIGgcJv+4JY16t5jxu2k3GxPJXv8cPmUjqTXnE9F
66q2R2BDKTYKKwqfPsPWbD50Ung/tp0ZNa61p5lkm3YtknBNqcFempdqpxJKwxlz
gTlVPiVkfIv4FzEi1NUGl+eq1YC+AcuaN1ldd3eUJF4XQ4uVs++dW3amPjRbR1AX
R3U17Z8pOuWZYg+VoMcKI1I4vxgXy3LBhodcMvFdZngLNzSt8tLS0VHrFGzyRnYV
gTHkhkhlM9TR8K8VfaHI066x8MS6ezDUEauvqhh7VXKT30V2LL7ZmIk6JvajNVjK
GFdgOo5IDnaY3x3EwZ5D9iKQO3HvLUaCMmUJBP4fLAbVvycHscNKFX6j51UJ4UV5
8+1bvrMo29z9uh2OU7Teu9H+QCNaW1A5lVQKUe0T75C5kpYoTrh5DS9gYiRHFGya
k54NgbOHRmB8Yam/umTwmsI/D31cYairSu0oA1izGOkIOJ9zx9QtuPBTUvyJAQUd
uKKDEuC5yFxgtXktsnq9h8Enb6jOh1KffzcB0mJ4leehiKmhHpG7yeWmDVHDsdWp
cvqYP3LXJOl4Nex6lUotnCgaBZHjBdutfeACSsjqMXI8BcbHxRR6cw9F0EvaRwE/
9HT3+hUUN8TFSEpCR+LcpKjAm3WkoYzUd5rs1W8REVH/rRGfPpQd63pXlWoT5Mxr
OAg8YFYz2kZqH5rGU0TRY1zov9JdCVGun0w/ehT4yu8Md4SLvlFfOBY8+jl5T9Mk
7VrdqtmVIh8UCyiq8/JOvmjwahrKvhG/NP50zV2bhxfE+SRDtIqXWAjjr8d2+sj0
AucyRK/AyRdjXuZOaYNzfMWAD9SNX9vh8DmrAgLdud+5aRjPFAIsQZt48U04hrVP
sMKU1lA6OAJZvps4rtiK3gRjsyCmAUo8duSoizRRxqdQ2wRLypBE+ltBsxbgtdXp
Ao9JHPs10MIsgQBKOWNMKbBTfo1ecUkVyJ1uFFsd9ciULDqrLuwfRXSQmgCzYz62
MxGh1vzjIn+6bHrXDAF7GhzqYB4Oto5udnLY7dfKqP1c/GGRV80AMTgeoAjzZ0kS
u6oA0124ZLOz9DSf45YoM9D8gBZUQdn1hPHQJCaNUjbcN8mdd2Kh5WewIYeaT7nQ
HrudXCwxoTRhfCiTiH7Rh+cjWDYABhXgIq6lS5JEdBagLG20DlM5rZpdnZTVXOg8
i2kSWdTigd8vH9oIuuM8PFLpe0G5ORm4slSqWVDNUO1h370x0ze3zJdcY+HIY6cU
Eug8nRz/Y2vDeVHWvM+m2nWMxpkTgi9q1ZsC/1G02cXS+0NaQbN/N9YvEAOo/qXs
V0tEwMXl3z5uv/7+rqKAc2JQFABpPwdYWGJleYeCDrUUOWxQSua3kg/wQ1eH3B71
JhUVJhxSW0F7EI3p6ZZT/PeVtd6QJ/L8yKkKDcA+l4UtLT7TU+hUhz2L5t+crxQQ
2mpdeGtCPJLohbsr9FmBUP044wfQBlYihvhK096hP586ieHPb+lSlCrpFo4kQVVt
F3cHtx4tx+Ya8JluohYS7vlBWQEReGuNwbK+eN0UtMyDyDefUCiWtgE7oKNv2irU
q2DaTn2rte/kHYPqhXQBQCVgckioRB20474ZkBKvSy0MHSyeuuUWPNQCc40cm545
77sXZZEN8B4ETMM9ZAoknuywcNmpIbGI/IxxuOAzluLA0ssoWeZE9Z+iNMXs51lu
YiutJnEubzF8zaU5N6BiWPpOMwxG63Z0ru6z5JWEeciKn4qolKMX6tAYPPhTWAHf
+Ev5BZfIiNkRdByUXtyBu3DypeJQ7JIUm1xvxJTOjrmxF1tqicC26bvVdLLepEdL
TpCYv5jZ6/nxclOsq0plEobJV2YNVb1XJxPhMGJEfV72Q7D3SljRh1EBqbUw9Av5
gjtGj+gG/4VWA1/7C3hB33a/Gv45eIYTtb1jV7r+/9uVrcy8jKByOAH80ifUmLyE
9MFy3RsQufcNP7cVPyMTqCDygTExUnE3i1nU34uMlsrRG7dhrBJmgwWu7HafJb9D
08ydR0MpZ+X8n03SrRJD3bh7yOzcXYS7Sphxink5xFRNFeCgT9Ul+2GrtlUw9HVr
qY6I/mjV6q8GlTCemT8Lgu4MT1VoONMNesCPg59sV8vYQhKnKeTUuOE0DTAmrcNu
H4yKAWgl/8I3cCu5j42mCTImFNn4+aplvejfPE0w++8+pBdyjTOaJt3u3bL7pyb6
MbiOs34MiAnPfg6T7gkUpXpXdysqOkmx2Code91sG1gIrOFWJAsmvP9YZDJMCCVA
Ex5sdY5XSH+alxFZQAj3jsGiYBtHX4GAUtXa3d/apBAQJy+GdD6ffzktDR1WjWBG
FW/ipAP90HtbAUCthX4zZZAOYyttUIDmI7xEisXaUg4Dlm1o0/3fx5uso6IPDYSP
Si2IlI4N7Qv5WoA6Emqfh0dTeTdtY+2TBb+6ioCh6Cm0vh3F400olhA8TZFOzDwP
UzR3Ast20StpXW5gjuteJFAfGiXxwXVNuJl9WWFh1uCUbqcF97l+4lKaF3O1a+TL
ZI/5+dPCilbyyYrJWWEdWdgmaTgaA3BpxtF9lfwiBcZRt3QgIvYDHnHjlRSx1ksP
zV6yDwfhlsEcqcI3iHcCco6mGlIUEN/c4bNkpoXpbMVkfrqRzZquUA5HVibNAjFt
N9u2xc9syaywTpZDIEdLZQ/MUV8K9vpK/inurS4ByozNmL3W1IweRO0k3nJqQa+l
Xy3Br9Ue+sRHQpgPW6ugSBaG7Fb0tAppsRq1OQHTmsTUyv54iuekABXbVRq4HAoz
iBHjNVTaGS3fJrQ17K/CjzJk5HEKBtNbDdyk0u2KiLcBVCfZgbEOrrLmJ0+9NvIn
wTwgj7+07NKDEQcNzghuN/hTqkg9av01fNMCDWqnwU2ObP7prKRWJGGFhd8TUWUr
HsoNlGvhAQEPGZqNNWa2vbxaDOwW6XWsBG2mVgQhM1GfuprfAtJl6rK2vmXAOFul
wv2RSwAT6s5h57tpXuyCTCOIoHykM2oZMilfU5sMG1n7tK176CQZ37cp3K3buk8v
exoia3zPH8gktDx8VDHigUi+RfrO1m5cZp7ulM8A5kvQXA9YffoG+vYXw50td5HJ
MrD9LVOZB1NfM2ydMKpaMKL0kufR/K/i9UVy/92jTfAuzMyhlDfXxGbb036Cfi9y
sRthbU6c5dCfMA7lyqM0c4YXvThYRh1c/PIUWVCYLxNXsZCgYZ7uBwI/SNBeKE8/
zsGU5VzwM0VBpD8ssUIgUOO45BeOhV4L+5WtDhBdGojs36Dxw7+bUXScaYd+d0R3
n2PZzUeBtvlCwMB2+wBALgAW6TrXKY1EOJ9UwXyOv22s4OmwqnlCRO6EIle+Fcnd
WwP1xMuWskxmSaC3uOgTDVuqrWHpSwuUvWx54qW4g8aIWTVHXGtWs/8RKqws+Vq6
tpvr6vpN3ZV/tfE0iMsWoqzKdBys9eEyVsb7lKcPluhNObxNTKcaB+TP7W/RZ3bu
2IUl8bnfDpckUVQrBZoewFyqw7L2J+ghU4twQ6ZeBhn0yLBB1ju6EwFbjKgZTSqF
R1sd5yVpP+Y5AsKs7lrA840XJLgcEmhRl/nuDShqHHJzZ0nF0RoDYqxEfGruW+L7
Uul/cv+VjYnafcxLojLrA+wZ6vG+7rKp1XKUojXsrp+witAKBY4pp2ZrWr1Ad2zi
tiPP5o7fcp56oS5Fvlq9mUvf0+wyRVUIaeJCK5X0cA+0Nonc4NJMwt5InmXjwEDC
gSUi9KQqU6NfzEIkUD2FcyvKLCC3lbPbLo0z5mSGMc+j4HR7lf1QOl40ZsiwHAAm
wPaHP46WPmR/lw0GO7ygGUCnZ2kXak0I+XGUYwwstnd/J8JZn1LmRcT9lb/O1TNc
2hy+PWEWuqkkfhMqlyMIL0Nlxg517iV+vvAVILrighIT2xVx+GoP6jYGnwOr1i3f
9qHCk5OO+htJ4LJtPkHobGnYvhTNSmPpFfRD2DBFugzIhrtxTPapNNonDzXzrDQQ
AH0hkaKEJgRS+93LIkebzJ6p8qKaBlFuswiIZ9fuJU5dbq1Dbf3uy0/CuaNhghTU
vw2vCNLrPP6Gh+BHc4LtR7ttZKD/DowKKxAllNveYACc7O1TKZtgA8ec3VWbj//j
SqDQ47RkxK/yccfZgtZDn/gpHg+rLbhamIBu4st1a7RrcFdSBzBs9fTOtU0Okfls
6puGZRdCI4/UecZ740+uvPQmm3FRZcybiIZ8igU5eWrdMuVg9WDypKAE3J7MyEQk
ojeeHW6Ujele6OId/z/h9PrNzJIiYnr+OXV6Z/QF6F5zLhpOQrY2vOrf5HnkxNa8
9BSb10hxRfFHxxzh9ZLg/S2Mjzt7RCqEVxO9/TV5QL5XMivQsg+cbju1QWkn3o56
HkJZ7oDv5znAL4KH7sNn/hCov8AbAic9kzs1puSU6em3+Z5qopyOxL84sPoLeCMe
02ZdXjLEiZTORQd1biuNO1dbGtK+rnMclMcFWxH5v6VnDXH0y8SycPXU8n46mulI
9sMoj14BmX20ECADPANbihhy+HAaPkPL9QVMbizNgdyI4fcxTgBk2/qBX3BbMZVd
m3Zi9JVz3fFQZo73Eg14UPrQbZ9e7APm+Zm3BQwbQEN/sJDCbdoel9mO6ZeRt2ue
sxmX5tuth5YQU4fYJ8FFR1eUCEjBoesSUmv1i8bG9iQkBQVG3uUg8Z3vOq1+4rrj
YJyU4ugb/5DNk+KikU9S9BOObjWT8J3yoqvd0b7IH57gjbAZVI+h8yKrEt1zbHOI
QwlLwOOGIHHowV5uq2juNhnYptaJhsFfJu8jvGYLCVQpCmaFuRhh6N7TlIQt0KBs
1WQbMl3eFj8wJYOGNYjpyjjPDX4WDxJAo89t8/o4p7c3eX05rU2cJx1WErWR8Q60
o6cnOWde3NcDUTpO7mAbEGI+TLAv6U1V6Axpiz4onZZhFz7TmyaJFgxClFhSrytA
4N0Xt9y3seQDKcSrFZuqu6FbbaEZNwmqhVmJDgtCK75UuIdeBPmQ/F2kPQfrRE/g
UQzJKLqwAgL39GvHx5ya7qekES4CL+4BxFSnwnIqNGsiojQb4L9b4i7LIIsD5AeC
u3pT2TKI4gaxsGxIRuucv+5f6noYeTypQt/+5fldNef7Q6HC3eD1j0S/3qWIijOL
nbd8mtyQJuL0dfgR4/Ii958EYLrF6adnEPHCqDZr6ie0FcKeMio7uJfW/KiokNr9
i4GDnUJQexji02JvUt/FWsYkM2c/mhj7SBVIH/mcHkLKnUu/NmJeemNua8PDRDQu
CddU2l0TmKo5QKLoK9ZUIVUyFbg66XQqiOITZaaNhuhQbqUZSao/XLP9r9ghGbw1
w0xWncapmDi+/7bJ7sUKbZ40PuVcmpt8g8Cd1OwNnXKaDrFjEjgw3sL8qgDAFaRL
8CHgbJF2bKGnvu/V4/BjGiFD8M07Zzw3lmNSHt+eN1Ly5huAwlCH9YB6RI1Re0Bh
exUHK6KJwb/TWPejm1WK5ZfZ9ML5aQyFyKjHpovyYU3eq6jSaud9YyDjXOMNV4MC
l0QgjFAQ5yYSODLXLlr+q+0elwuaguIQnctrNoPKRWocOvB2IXbFAbQa5Ze7y5hP
s6OjL6S3CW1pRRIUGSyRP6F7Zb02Kpe8QJ63HlqU1GaDPXfZJRl1IRchE5ktDalt
Lh6eaJySM7+HE+b8vj3ywHs5UyYHk7mpdXqBuvzYleVHSbXYdXsivMKx07VD/IiT
yDc/GWL18BxBSQiiHq1DWaL1YWyf4EOifzsxdVkz/VqN6ILp2MvIkEVql1xRDqS9
mzN+K+bpaG5j1SjCOaKJ/4JB9nP+12Ne8VWcQDWqx5qypS3rP91pvC+c93OnxTmZ
HKHspvAC0pTwvJSAf9909fGnvao7fNgstrarTLkgwXLNgUjGdTBApGUX5LEaZNls
oaSL82bHjfrRQ3BOIcJAikb0MvAHz+wpCMbEAKgT2X50zWPX3jR4aw+Q0NJkhBlt
E/dxwSsNnEYcKAa3XWKYT0m8HyleIOinSB7WMxri3RD3fsAkud+DCthijm+6G7B2
xQCJH7rssD7aZ/5JMufuclgwIloDcx+NN9njOoxtHfKhpQV2o7qvu7cNfHb4h5P9
Oe5KzWx8SGYYbvntsOFVRc/ZEBqJ2Ih9uPVOQGgHyIsEzVHl+/AE+xor04PZ25Ne
6kvpUdPFKWq+ZNAUmSnH88h6qWStXd7qygUxr+rEJ2iDRSchN9e+Ysi4m4P3l3qf
dfAcbfw6Iox/wq4XtC/zbgiM3DAFc80ZBiyD2r8a66WisGlfosVf/70Ovlfa1QKo
CA7wiPkL/nN1JofoJtCmzhlG20Hsm2TL/zLfpKDCcfJ7yAgwIlCToY6oDVa+hDDl
bNPA3Lop0zJ+Y2+LDFsp3UgNlPsRFUr1vPN8RTy7X4N1SQFtKWoGzZLQJAnYgjcm
11RNXeO/BlQUqW2+tlG/nRQeKUd0oyNdNO0LUec+jvHiONCTHOGLnWhyKR3uFP3i
OMxxlc1ZYYFGvADN9gqfXwbLwVc21e2CCQgadlwUJQxVOzQ44A710EGzKHUCxExT
EkEwMu2CH5jTrihieSAVlxBrAdBI/ehQFGuAhTPRGvOMZRAHtMHFrzYBSg5Rnzvp
Z8uWtRhUl/yZReYiETzoX9Q+nEiPMYXbA50siAD1vyCRFXRcbeYQDPI4KPgu97mS
7PS7v6mDnWy/s3ohbxYOD8YdD3Vg5fLIE8F3mg+Tc3djCrtwDaykXGoTsAPu09ns
rMwc8bEkdTnzq+MH9/SMYTbfzfHkrPIrU+Fq4jzAnIGI4yIdiD4pem6wS6O19tEK
ZfD6XNoYVr9ch82cCbMBlbhE8E3yfba26SsyGjaCWszNMPyVppPLwzo0fxP9TUz2
OAD92GetOzEGJDuF45iTVFONP94RhRap3zhSIwLH4R4Frf7I9zgoCotck7S9fIx8
2VKeG5ntAfTyRtgViSZhOwYZCrNwRJ5sSMwhsKsFvuhfeDs1DBgNXvgHHYjSss4L
gRo8HaAxGZiA7JtMiUvJPEEiGMY+VFgZoxeglwTimCyzMVPeRpsMG9/xfJ5jGGCo
TW/nTzgFfQfOMGbRxiflMi0rjYZ+xpgUi8GUpgw2OQh8RzSt/iLJp9AyG6pnIxrJ
aPQS/MVNzLgdUGEiJf0f6TCMEwOF7zEkXtddwNC5Qg4dYZEwvHMwCLXc8wNPJn2c
Qd3MT6PUYb6lAD9oJgyxrTSNUK5LcRUJDAOr2uzs8diYFakK6E7trK4QfQKeGRpy
Bwhry7lj9iiLQiVsquFgYdNQXuQBaG8aIS+Ng54i2zv+yBuUTvm5ZXfBIFIAAaD0
59h/r5u11RquqSPQZs5/Mw7w9Bto3FIvqhNu1JzSUuzMvSrFtodygctouU4QdP3h
sgbvBwXkc/vNhdub51GzFFo14TryoEQEFWo61n8HMwxDsob6AAm86tJGTzXymoCG
tLdrVF0RSxJBC2rUsFXSTDw2QOEG7SCDdHDpL3Nf+T2FX6LAiRKfXL1ruodmNkxv
DFfxKVQBrS7y6Eq+zP7JbFK8UxzCVCRmIuRfDjzuL85O7JQn4QJWY86SvHrsjlCz
RsLDdC/mpXM+o4kWULTv+D05SRipVo9aCD5dIcV7LGfk3PGujERpH/2LGa+FrMf9
+4353plewL4g650T5lI05a8Sfcd3Zruxuy1mj0IZ54JGuDGY8DISNdNjP2NnlVsO
QSeBt0lWqtLX296P5tR9a6khbI7spgFSADbK97N1xPhL/R2QzrXRtxgvQKcL8Lkn
xKUUuZJwkcJfWFYWrpnAQ4r3tohdW+ACAKB+AySv629F6oa28O7SG08vBnTfoq7S
0zEnxTvDFiDqGkoR7ihdse+20crZau/l0fbcSq3LDJHLdftAJHQabTmvh6iAJqm4
2cJxDImdb51lnmAUL5dP6++ZdJpjJEi8dkwqqcC/OEeTXfxMNJW6rwVCrJHpzr9d
EkS4uXwn79dMKawZ3Jj/W74DwGKCLLiAHK5WLL6aKYUY1GhBs+f+CSFE2/9qeD6S
EmYAw4g97j76E0sGPrnoOkOtp8KFgHxGc8jQoCJObcWCINUKN+HXrjC7B+53hNOe
FpYvqnlhFWOeC1KXLi4npWzBn4+eKdg0BXO4PmZOgBNrHjQaVqhvmpI4r+gHra2z
i6ZhLBwbBRAH7QCBwtapgFSDCiAsg8SeAcZcZxPCIi6e7nC+NdE9EZO1mx+k2vdY
WUQvodTPZv80J+ldKUT4XFWtqxXB1ZajPQ6Pf9GZc1bIxqXmf+wD8ukFkWZYMuzh
1/ENeLMRS97xfUfF/DMi1lPyDmnCTPZ0Ei+5RBhY0VEPZD1hKtVnZMO7GPCgS5In
qsM3o8nHRsUG2EYNlwOJdBJKETIKHXKSwUC1s7Nu4sdVn4hMyjWMOOn2DtkYlY78
sboL6jb7pId5QeoTq93WZ4nQMMd2SXFLm2wEFB6t6Ajlf98rTMOsquskR/e7lS78
ES9leKfQKrB/kbgKK6lwhs/uN4esQXNJHLzsvQm4wqjOqO33Q0fF2F6pjZ3Lj6vt
Jsll8Qe2n/grTQClH6K/t1NRqTa0AM+r2eGPE3wMiEhop2vSteHwkrOTnj4vcWxj
zpkrh16jCfMvrsx/1BQ34QiL/BkJBS5xyhua9aniI4amH6lXat0qIbP+7ig20O4w
Nal+mWXDSSbym3KoaX/gQseyW9qvgiTN3636TCtn97n4LqIauFmA0agYfGpKRIOQ
pCBfLqeT/ZZJO3gJAZB+wGcCIgN30R6qw0eNl0mR1yvLy4hoDDeEidmlsBLuFPnQ
5eonTHsTc5Lp59ecVYNefGXaKRSce7zhkwPHBLQ9hgZXUCV4mFL1lwcg8JN3x7Jk
eJKcLu/bV7oK5BZDrWhoABzOCP4QBCj3RQGZ5wlTezbRV42/0x7Y8eFkqAhpIZC3
wkkPAMN98BBvn4WFrAYfwlmCuu6615ifU5Wu/tU3XRFq9T5G4eMetpP0EjE9qF2x
c7scuZUxsBAzF/A36TyUeUer1XcjHwzWme/NWFBW8UVMwtUqXuhInRGo8kfaWAEA
7+BS74HWTFQ5NFwcNMls0MW2KYwmDO9uPRVDyoToLhoQRgHduWmnz3WaLPxYjHr3
6mU615qT4UhG3AbNjNMQd04ZRF3TNAvq18ltZifqiWv7INHnfsJOuYRNdzzzT6T5
p9Et6H5r6DSeVnPD+ox7cHNcSQz4rNgO2VNWNWcQ+TYZnZ6mrk1THxUvqRz411H+
1yxbvacJv084FOqJVB8fgYkbjVr7pzRRa36z2Dh9smgU5iwQMDZsk2av1b3lGXhR
KhYqmaLoU45Yb4cLKACHoKfNbqiTXBrivmY9fyDHOWF40pUdMHscBhuR6hGJrt/B
RyGy2OSJ0s/+MB0iuOnAAMQyQO+Rd0TRBLMNC/4qlGy8e3o245O6j9bTdDivOnvT
/kZGA+MCgEbN/GQo2iyTr008j44uTQrHOO5hLiOVyY8JjlmC6T1XCrlaxZjleljn
OpOUH1Y+rtN+gMOg3fb6cN3Aq6l2ik8gJlG1rHaJMmIWtAGiNhxl9ObJunimyVUE
cwya4Q47UroMZx8REvAqJ0BLPbuYaeWHwyOmcvhY8tMlWVQc5FC1nyMhsIFAblxr
5SYELg8IFQ14DYu7BwegiDe5Np3rWOxRqVisq1nxLm7EgWFz+Mc9Xpdj6Sw+d6Ju
PsGYkoyOVunmhS5LVlEOWb1HeWjRb2HCplhB6uuaJDJjA2unYyw8HoGkMj1wemnL
LSiywLbA838YgyRlfDD+BG47Y8QSkSB1oLcMIiD9D/HTeDVycIoWJbhVipqjssnR
vJc/Yu2x3GeQkBPcPuoR1+KQPGj7kHzfs237yo05KpGcjDNOhltS76kgqNjcJsxo
Wyn8uzVCGRM+sKlVWRqHlTqHtRa5As42tW59Z5vifZK2WW6oroAzbe2OH67IgrkM
DcOORYQs+5k4nXerfzsjepqRQqymz6xxdL133gr8Sgnk8vhHWwWlOpGyH5IWxQ4I
PYc15c1NGCgjZCoQgG7913LO04pfApDsNZ0PZQD/JI04TWY9VnkN6lEAhisANkdY
YMvIQOv0KJ1h0LhQn6XP8bxjf/qAXHg6sElGjtHtuz6x7UdXSN72S+72NyWVDdPc
teqW7mot6OZhgWnrL7S2m/krZ8GaNDgHcc0gR2CFYwZ9ShKwSlgQD4xNf0y0MfYT
W7OojgG9NIkLAlMqVxEqiSAPTbfLGi/slbTOsoqZrA7SDkQ96rryAG5SPVFKqNuJ
zclAGGScUgZkFKDKvS0Rp4qKUTixQc600cBgC7avecfZi/Tt4CrYU924upJq4hNt
0847E1s3KZvWurGPZHRYJYMOICzAF7nIZoO87x3d8RP4qDhjBK41BCvB36wriyWz
NT23w75XGJ15bVOgvKgQkF/Aoxm81YullRL+OhGRMYhgRhbat/QhoA7jbKWdvZ7C
M1bx2PuMF4A8D6QxIsBRjnzNeQ2V6aPwuSYpQ2ZD6P1MzeDCFDiHd+bp0YKqtZ4/
xqsVLjTMRPNQZenbdRqygi8VfmXBzo97Mgmmy91Pc5AgtHWBylT5LWd36FN8vF/+
jdwMS2MJVOx7REVeklftgdWXzQMdLQSFZX0RWFHtTjL7Uj1YEoyTd2UBuDI5Ci4x
KEzFKJPpdcfBFx4Xq8cyVo2XRVNaFRbvKEvKAWn/j78CEc4m+0TSZNx/pDbhpCF6
Obph9iUmn4Zfnww+J/akAlfZZpuixqtxJLfnXHUAnzBQ5xiLMMlj3m4lH5cm8BXk
hCK8Hz52SxXPHEg4bQDoneT+Ty9+qZ+ZwDXb96FJKQK5fkh5af+AdQSicIMNRM/a
2IznBYrIhfJ16K5gBQWS05pTSUbztnJ0TIurT78w238msIF04SGY4f3Dv3Uqe4ld
5ZTGuundqn4FwSa2oRzDQcudReC0S0jV0TLVz3ails6rW4hdRMb/WGWP2ED9uuyM
+igh/+fGa4n9fDJ4eiSYON3/sIQREP5A/lbFGPYGzSI0UIRoU5PGidF1k8tzJ0CP
MWzSX8Q3xLR55GIBbQkcHFzQMMTZGI//6npG4U3tiWXh0silPVneUcdFhFexlX+V
R0GooVAaFYB25MNXRHRL9Rvbm/7A8LEArax/zMAd6d95fuffBe8LX2VWn3pvXl/i
pbNgfurq6Zi1zrbsgFeULC3MGJnXaHCcpN1ZffHH2k7hWQNuFwPy7+Kbb99+pg/x
edFAoeYPXZbRuVAAFadc+IyvrUB2x1tT7/izlABKY057AsWeZnRywZI2/k43NkLc
qJryBIJsnCIVmznmK/ABMRBH5/zDilK9Ho58Y1pLSnn5FnaCZsCjxbFYhqIr0iIf
jRRVkB7Gs2GikItzvJblIGjrmVCi64/9RR9aR+vGUad6TAmsSCsK5j3bp4NcqlGN
yx+/FDkENxuFxJ9IhKpyu0D4FT3UA56YgpOSxt8u93gvSEM1y7Cd26Sr+kDL5u5I
/H0z17eRjrhilWe6m4CcNR8N9EyhKuMYuDrugJA7p32Iu+TiO/oPWNQXcsBwQp5O
sP2xwzIV+bNEW4Zf94WJPk7WP9H9JvuetrH7VSkvy9bWC7MSSd/qRYt5zUm3RLVz
Xpi30w7iRypddf4jCg3EIuumI7GQlGfyWCU+HFTJG4C6cW1dD7Dq9rYOmlaCV1V0
Vb8kl0aQVbpf95Naid6m1miCFWjm1kbbJxRzqDKMMiIQh6nfNypMXIP/BGKokfoO
hURsLEPMlCva/iLpbVTICzhSl76ff4QSVLXcIBV8CezL0U7t0vaC5FfXeymw506h
wNfoFqxNvbGfH4r1ppQcYT0IVY5p8M4Ho6/9iC7J3hmlBYtr6tDdmkWNsDmCXxau
neD1Sd3rbkCcAgbBxpAHBxQFi22WnhhQNnhWO+v+5aLyGBBP4FKfLjzKEfUwsmhV
JPPLU1dEI1S5K9yLbd6djRRewdIsv+/cS6Dnhw51e3xscSI85xnGNNL1zt911AAr
cY8QMOs65MFWHK35f02GTmwTu5/p/mDNdasIJXCIYtXzy3f2fv+CT/XhkLUAxEfQ
e3aHEbKH6P6palPw6/ATxM6xnHlAwMg8KZbVNLCF7BUKYen5W8f5w94IsFbA/2rK
Sornk0b9nbLn3cA4mRxHqfYpPPgMPCgNWYsYxPosAnlDErtXw8cnOFiEyY5Wo6yW
71/loisOl966Bm2DxhQ+wbQbFZpS62Aa8FIorQgfOXDRakvRE0Jzkxx9h2n2r+EF
fBynOGMy6cBYUJGMtgA7aCARUYOZ3W65qqJ1MENy73lqvZth+bWAgYm0tkiGQRBx
Yd2d2GgoA9s0e56wJCnPPFIX1VZz79MAn/1PTtccLnxtBmzgH8EJWC5BPy30JSIc
cMQQ96SpMiTeJ/KA0TgZY2pmEqrfEhaZ1yhwBpNoErZCUrHKRJPpFdFIsctRomlv
qJwTuh6lI90A2LYlPxPpdeVDH4JpbWuoljNYCz/Qe7RGE0DA62o8Yo/i3oDQRluZ
gZKyq+wxHWAK9HgqsMRIBI1eD3WEW5qH79Tuh0vT5xynzNaYvaxz8W5sGUQacnSW
8NdN2fEl6U739P6ooiK2syNqTTXVkTCTDfuRdYkcceHbiTL+rgyS9rkbpzL+7CHA
kvcF6sRClX/VPltfBBO/kGzTS2Dikf62ukoLCDrszLrZMrzu8M/25sFlSQ3gM1co
gUEB6QWE4LK141Oa16zxJGtBVFjH/ug/4UxuZ6XD74GIrDvlXAAQJCfMltiKK59Q
6Xudzn0tKtCkjycevImIMEl+XrgDptfI17TWVy0SvAuiJRRRlWlQDt+m1JrRO0O2
NrOLKWd24JccPKQJ8YbcekXj6D+QWKYZ61ubx/IN7ma/0VwVA1/87fwJmhYlrjYE
q01GET9MVln2HB/M+oAiHHPlMMd+2tQvONdaKlsCMEvrgIwwRDo1IClC5k5jE7pq
mi2PFgH6vj3PjkDUp0scBsg+fPQl98s4OM6WfxTjtPUKPU/knt3rKx23FUbBdjPY
j9YQSkbU0d1FxVQQRa6nwmFbARUUZvEFRqhETRx5Ejs/To4LcOHldlmMxeOi6dVB
MY9CcsEOI78WcBPz0vZhYudOeTOulaulKNnzeqLmlz9EiADiKNxceEX20v52eTp7
ptEjqTKYWbHlwubEtwUNYBDiYi/cDOQRUz0A/4V+QqIYi7I4aw5PjFYwqfHlfzvj
q0vpi17ljx6z+XQkzj/OjwKrihrMQ2tgxpfkUbVGSS7lZj/pd/Tzi1yYKKgjtX62
p/juMs1CtIPEhKONFk0Pwz9sA7Jo4rkGJYNXps7uhcu+LnEKQ1ml8cgpEK1OHtAr
yC9f3nAy9YiS3tvIc08rroAPrME8p/2igaME+9tN4AXClbYkN5wrkEQuhYMy4krx
BYadv8+PvshrmeUkpZci+KA1Lb9VAuIWdXd1lgtWNljarwhubaQPLsGnF3iQIWnl
8ZYqPrc7QfMF0cgg+IoCK5skV4j678hgxHBlx8KrrPkjh3RgysfFwEUYdz8RlD+i
BrvshJpaqTlxT54PYiTzTpSSjvMcypfBz0Koij8YEwv03fjlKMrehviJMM7O2v6b
wSM8UQFBRd8r9M5D5ycFmXgiu1/16XMBprtPu4pMIt9QXPJyhQfw69TQhwhd7FGs
aE4DpzgxJVqpwgpK3jaYL+7HkTqx5t02ROQrt/3V8t44ppW9kBdl1VxoP2C7N+SW
23rGm6kSZhShjNr3LbuqEqY6yPwmTdBnDDdV7gvj6cU+OCjZE1irfN5aslL42WYv
FLWk4Bu1bpvcZnWpmYyEp5auCuLkJieAEolnS895XasX9j8Wnba0RRA+W80+IX5a
TYf5gzbqHv87m/j+Q+0kIxKCx/nSL1/19Kn9+u8yksP8R96mILgOhGSOGv2L7Y+j
yOoNricekDeoKTJxrX8F4CGJbx/CxFmTyCGn/x/6JucouLDoACvEljAMl6PjKWji
G9LDOEV9OF0xnNhDrZyJyTg7D2AmNJY0cPuxAzt3tYxGPKkkhtCbXOzhsAl/Hyfd
kZjiBYh4S6VR1navWS4VEjBaJqHmzLmS9dDeVy27ZScA4UVrpysFC/E7hkURZs7W
TfKubPG0BeAz1VbShIjx3gycFSXhpVEIa8fdrDhE3zbkhquWO6b0MarpIAJzFkQa
2HRUjStCRTM7Wv6V33qybOmlb7RW9eAyY1yayRUAdvUr9pzYBuCxKSK4IQCDRYNt
hpDJ388SNRuznCIQ42aSir0Y0y8aNhhPWKWwhGMoT9pKM07scZyQsOzP11wT17C5
Lj7GaoWICZcs5cwvAL9WlxZLCXrmnaA8aO3TZBYZXPeRgCOJSxjEaqATtiKWGNAD
vqMgGjNlZq5FipEB54qzUjVJR5rB/kh+0Qx8sDNcjdIpjI9yGBhyc8L1RTccQwEU
fAeaZ5wiu1Rc6AsOmhAc9SjTJuZEdV9fAn/Fp6/O6u3y5m1Ar/vhQmloWUsGCtW6
MqdwyQ2BfZEmdfZjyxhUKgnhZ+Lu3iq2TcN4c0no8c8vLdYBuxoQxIM2avkUk7Sf
eX5H39jXEbUArJ0S2bjKUieqoijqT0dGHb8AfJ2Z2YhaJg+d3DN+uvel6vYNcL+I
Ruu8faMHZ/N45Q1gGBmfWURoBCMnXq9BQ1clsWuc+SUcxlDFPfjnZD0m83b6GkTs
kGzYlTEFhJvwEezfRl6LHszEVYEIfxGbE7Wzp/RLFKChK0nuk0D8LvcaGM6PH/96
vgczeeEGK0GUXw/inwDn+IFiEoA0WZd+CyT0wq+t+gUe+1bCkU05+yqBNc2541ja
iMp1NX0oOr5YuW6Sk1c06PCsFgOVWhu/zaI3qh/gY1Vy0/FMnXLgF57Lgl+KV6FW
ju0twMdO8Rjr9K2wSY0+SoCoprwlFUgFcG1VQgNhw5XLbLAluumSr3I7y11ltIPV
Jgm3o7l41LhXVbbEwxJutF16DG30IPhPiL8KO9wf9vWRp3R6diBHLJhNlWjFgUtw
rcUgy3Uipd/dddA5LZzy4X79MNz3BPDXpMiDD94UsFjUS0C+3mZDNds7zrgpq8xK
8EdQJDDcQSV8DY9zU2YD+u4y4iv2SF5i0YBseH3nGtEXYPdi3+Vkre8xANIA14ij
oP2Pnz9Y3kuMy8Ba9mE/ARlfjht29IY5SlCv5BhGN7pmSTkyuwh3UxxcUHPnuzpQ
vHh+OYU5V0IyeELxQT6ZtUS7TJ9CQe62t+g1fXqVEDiHdeDSw7QAcK89zpMLxwYl
65oNlGxdeLETMj/ijpSD5JWT5oJZza0HQoR+v1nESEG3oMSk4g/MN330rpLs1zR7
3LOvQFgCu6k4Epmnpr2uNoMBF3vkGJur+XqbTGnuba/bYMHtpF8paH6dOToS6HCI
fJhxmJRzn3mPJtbFmPqmdG1TlvGxiu63BEmyV2916HjqYwSEMiV4SolQrgHXtWWR
abBDppzRazbSpIpocYlfe9nGg0iichGN2cXQCdrVii817maMwWRzoywXtTqRiPkt
GW+LAdUWbuKZSBWaDCpgsQbeV6Htx9SQwdeziEvhDvR6AINEAXS7o5Ad0BQNqDaj
8HIsa85ha2fgJNxVktGqUuRNTVFCMNlqHAVlw3WQOd9gr2yk1WsoqpNM+hqkdD5T
RYxvquypiZuOyxDQsW0mW/F253Yt7Db0eh9VcB2om6o7hA/RmHNJU7ufR6uV9hAg
+cW+Ne7DR5LChpSIpk3FKGyfKihZ5EMd70+nKxLSbv9L8vA1fKcOfr1fa5rVyt/B
vrr7sqfXJuIExz67c9jZyMDtjxW9JHY9d4AvOq2JQBIC5plXXvf+RimD0TN9XGi1
C1mpJy7DIDPK1odwYHKBKEu5+Ut3lQgicd2e0BbzsYxa/D1yuYnO4pJTdVr8/dGv
Km9wwLYJJut3Zfi6ZkebutMjA6nM8rSpUf6chCHM5hOiojxX9xPIZ3jHTkHHuDdB
fejVOuEdGQmTmoGpt7XwEKWz87JkM0Hw2tphkn/TGcyJpibeNxc9qgI22+BVpobf
FSHG0G00punJdAvZRJr8Pz89+u0BFr4zJJuXhibh9/OrTZeyXLcGGlyrDgGkSnzX
PR/vt5bKf9PH2ifSMcOEQoIfTOvKc32Dc7VqzlEjtPZ1aeIRKgsqM7NTZJGi8DnS
ScJrapU4LK8I79ymC6hlLTW7fJdw2JIsFgFzIun7RcIZIBDiABcMoBjuA1DPX6+R
gWnsWHP03/E0kjlnzkO7VcUYGrnbAug8iVx5QMWTTCFj7HvQGD2V2j8/7ADY/DBf
jIfY7RRWlALY3fMsnUJp98pWKIMRmxrSFPBiW/Yoe1t+lL36QH/9hGbNKGrAo3Rw
3K1JT0+Gr5vJJXBeZDq5qbssfxS1uCMA0/UQNOwKdgbw7g54k+9TStywsulLqA67
0inDrZfzKDMoV0x5oPj3SVaQSVVNz5OV5yTm4szU0HoRE2FeCmCzupjR4yAPieP+
Urzgtn+dmerezW8+1ix5SKOkMyzJpMgIkbx15pPX1QEK24Px4CDCf/23RHgvhw2u
Rspn09ELoLUwO1ycTjTuinOdJ9G/2QYtMdlRtFQ83dbrtkHVyVfHzudbeFVK5gZc
TdEcgf0l6QoufbRO4dbxWhcTsW77jSUu6AvtCmFA19esMqjzrp5sSlr3ddlsk++R
hpCrdM9Z9r7TM6+aZnhGVYww41fQn/GkILACDlo++8G/Iih70DmFaUXwiwkIof0G
Wmi4f9X69M9Jh4xd3RQ5Vf1bOTCev162Zc3/PCpnBWuP+K6hFZ+ZmtFjc9M5Wzjc
eBayqw0X6Z8Aa13tlhZQaVuJul5BYowQhjfQkp9UjnR2p2u3Cfm5ugk5uT7P9SWb
Dcnar+a87kyAy9BeHieJEkkZqccHQCvgx6P9/ExvsTRSUYW1dsaGdJrQTElxDxp6
LKTHTmbqL5KTr6qnlm1hIlNrybDACS8jOL+VIeyOohal8ZDHJRrriJvP3gk8BMv/
D4c4FcNkXC54SMCfLnVWl8YEWalIUZwqrJ/ROyXs1hMTGrajshh+F516F8mMY1DE
+7s+r7M2ly5RqybYc1iH0XULOxCld+plG+TQPfvj4o5GxPZ7/WBueYzdxaZt/JAl
rk8+J+10PmZTBtZBSaMbsqg8FbGDsgiC4cUtxt+KIUYUIu44IAvmDbXtU7FNNis3
+1TjzKZKrMwrd2UIevY/N6AeNOg3JncH9R5C/KjypE1mPhhHcrG31rmcmkR1ZQxS
BXKWMtY9gbudQFor/JzWBvO9LBsW2dXJus1EO5rgPLix/LH27gnUbq2+17/+wWsO
bSW4EDYTMxNl3QTF56uiDuGEllum7+9uZH1OK0oJx+4mbhMRIApaj+ZfHsKlcd2O
rWLkqhaK8xAMlPUNZsEwAKSoV6H8eeTbKMEiNG817BXFoLA3PvIuw194DbwNRPhV
FxiYHtf5roz2M2JMm1HWt+YKjJH7yRw0xsZQL91w5dXbtMRvGB4lUeDg4oKkaccr
+tDZY8AZwgK8na9LyI4dUF3g5Rr13b0O+aBUu3evcczR82mpxu+rIFvvuxFHS3Y1
gdaSXFEBM9BSEEMbf/f+p9IT4GqmOcSO0iX5yc+XCoRAVxID/B2UXzU43hznTGk8
pgnteRAWFnBruXzE9sGAoE2waTOqmtVuUVPEPdwfjCZQ068lcQaCkMrc2stzCfbW
fFN42i0zaMSDC6uehOqnA1nsCvotbMEKBKs3907DVOFGLyhJJCSlcZNojYe15X9g
56Cki6jijaEg++2fjqzAru00G2wsDZI8N+soXosRz98OLFSYng55nyyunRFDTl/h
McSGvYvhzmu7Vm+6BQ1H42qU6NDaBOkh6MWsNuCUltTo91zgxqVlZ4lsROM+JxaC
HdH4DOyVwzLurwD/0txDThaXu3hy6rwwzbCXLnlpeC73fnaIntc2qJ8tcWjYRhqg
Wl12GZbCNOqWOxkMtAORcL1fQeOR48OTwXdedUlGMgGtcZ5C4cCiVf8LPDnRWzGH
rj06nd+iBa92iqfAqGZUuRIndLggtdHthv4Xdv1eCp+qDc2aUhQ3htbWVmE7maFF
fYMDpmEWcNxX1DKAkOMymefVSYoYdoVany9FCZcVDX5N5dfJuBPBcbhzyWsi+Kjf
D/ToF5lqgBL8XPt9fezbW+nl80W2GQBTy4sKQzZ46T15TZTurh+EXfc9DFS0+Rfs
edhFG1/CFeZpVtbJsxzRnlhOVnX7xpsOEdINFtUCKuiZymK+ATcZQTZGg+/BqvF1
M2vd2dt/5Pir48WCV684GnME5AcvubvNOVKv+sz51KxyUA5cfRmum4iah88u3rIM
F4szEoPWlYOul7B2hW8Dwy1tXtcLGFcSU0XKZwH8ch/Or8I+mCjxyTZAWdJcH68V
QB+qTl54abhRvnI4nk0OXw3yrnD0WSh+94seq8qSOsg/hKLRB7e5gEdoOw5Vqiqv
Iow5xSwgZBCmY5uL7RnGexUBbYZ+IGJQ/L+tfV+9CTE5ZQSGFDa4ASo6rD6gx/9w
pKjvorlA9PzAgdwHDQp0kXStAOdg6p1VtA3cHY24a0cTI9aHbOS+ztUPok2mhw18
b+QhMrwUuPB0B6AMI7y9aj3MPdbt+gEqM99YT/3vKgizYVSdglLyFJz87dv05g0Q
7Mt/ySIcRLJvct5CgnESRJKLsYpFj9PZeWf3CxIVVNpEXfqW9/oAHTAyM83xxK6+
aEBLJIPYfW2gPDp+OLHwuNxpBg5cFSzSO8oMMtx+Mfcr41PlzQko4Fmrl9b87fXc
qfeWNenweNuAVgco18zl7j9IHi6o1g3Z6/qYoX1ZxV0ZcVI7aUZHSbqqAvOXf796
Pfbo9UndYmDHkta3TBSd1Pv3mKUfPrNxVKLH0rowpODP2dpAwbx38O0w15pqoAx/
DBhq2ARlgxoQTdgMf38Nu2Gl7VLxIqagtfAVTQ1tgG3GGB5k8Eig954KFyz4Rspv
JQdMwiMDNe5Qc7PRuDakpcIBZZEm6YHfvIA57QsNUQEPi9goQGa/rWY6YjW533vf
x6hMSybTMXswWavHGqiq0Bb+cyK8TUzAkHUeyqsWfSOaqosbFzGc00G3YfMEZGzN
Boo5Axu/lxWpHY5gpbA6+8aePMcKudt9zY/gEgBvj/toe35SkWjvNwspbHKDbpKp
tQ1WkHvXLLCPvM2Fq491nZGNNCUexgMF4T5WFCSywkINabU/v7puoBpIu3tGu7IF
Ge2uqTYn3Wg25c4tMsj7CParHukVOJawAGD6AlSiML4WzHOZV+vsqD1wnVeqAkhJ
nIntYngwdOjJK0MDHlLfAY5QgSbEIrsKCLeMaPk7/Q2Ao+O5GH/IXejp0UnV3+Tq
V6c87IsJ1b18YdRViyOaMsGbTRyzmUtuuku1i1TuhhBsYc6IxrVyTHAoVpQ2+VzY
OPNktk5J4FvuJ9aa/+n4PwukvH3trNiZGfjugx3vM+c/haOjnHnpDQ3AvJ0QXvvr
IEPO3gzxOzHxqAoOs3BFbl7xSqWxexUooel2DZmOI+D7kQMT6+MtNJtAgRBlMvw2
+yy2qiSO0U9Q/fb9vfUfs0tGp8+YVzTjkm6fHaPCkAUHruP4RhrysE1Fr1WkQwbw
NAg8axQL+uYyVcxku/7jxRIYk9aAYoFkbTzz4KKKGk1JQHejQxQEyWBfyugpmbf5
S65wYHj8RWQc/4GQw8HT1kxPNwS6pFJCBmtfZJHeEu7SWbyWWYx0B5vWWoaOGQrB
+xPj24Ayp1y6w6czWLYKACkMzN+qgbUH6vkeTSnaRnF/z5dtLuxszykVWvnubmF+
umIPFihZs3oSQ4VgrQLtK5cUwe0W/JUUuliZ4IWK/TMkJ7z23Fz79z5aJONshvr7
G2DZzQ2AUOioUWr2/to/Hkoq9TV3gK3oScJQb/pxyi4cqhS+kdPdLqDyatYHGMVu
/gNYNbY4FHy5SJYGJmydJnX45BP/6FyPawCAd+Kc5qQQkNQcD2DtL5jXZwf5KKaF
wGiuNlJo/pA2XuMdCAs6DPJEPl+f6YcicyRRciGU26we1pkiiN5169hA8qU3z5vI
dw1odoADXnrKDN93xaANTjsswBXTZoxF8bcf/zIdVLUFiHruvnW0h1mq5VZ0Q+iH
6mVWxnCAJtVgGUKEHgyKjenGM/jOgdB59/bVVxeoq3nwpf2THmViWoJpALRM42nK
PlgUzNGyxvO1nJe44BVs0a2cvkC+fRH5YdO6e+VQZJg75Mz7JcG4OwiURY37mRIB
e5KP5qDG+gys5lHt618uO9q1hlYsnHhO9lWw+ICtxAvoqSiLAcgBVj99fGgTtOTU
WDChoCwf97xC395qkNR9x0Pu6BLXt0i8IEQXetNn9sLKTh6bayemysvkHEbgxHGa
xO0hsC1lwi/2T8XMGhLpN+DTfzs4BaS6vGAULga2QNjU4Qrm8xie1fGGp/i6M5f4
G8Ep3mwqZoiUG5ZOzAM1bk1WH5hHv8h2LAn5nhWyy7tjr/KI7lufQcbUTXfdzyB+
P0HLDXw/qGlibK22W4mNkY+LNgVasFMeRerJ4Io9tvQ8g2tbrritsiOhOcLwD+T8
NUj+a+8MQZozm8sIqbeTYeMcHGRmnmqBdm8ywZSeAO7r4tMtUEDMKEwFqHLVBcWp
3PWaH57oemPEDhGaL0Ffaa8SvMrrFOiC8uV1y4yt4XX+HeaViDw4m5QO08g7Edy/
MsonxtS/9SNLssTrhjusON3i2hS/7ZnbtxfGnTPJitrS0thyzkYjQY6YQJH1vb4e
yFRXGEoo8JX91ocKHd/tXoX7Ot5PStvvJvuX8hGP/mG7n+t5pMYhcCNzQqrFhTGO
m+oMnVxc2TiMLURMw/zqaysyJQvFt9jmu0W6oR0lVDjSAryhrEMtifFkcigSRXTH
oYfI/1jah3oZSkL1t7R+RLzMyGOIzEYQOdl4f9N5GfR3L4szviLhOk5AT75yXdbD
GQv21HeqxjDvWIduic03BnBerj7K37zEsNXaOXNZUYvk/Agx00vk8LCVBjtxDhEU
6pW34CjTuihUqVCaRXgfKt/mqyfRVVPr6HeO8NS6yDVPm94lArHZ6grGGZxbbmF6
8iJpyiNKb5Wt0n6hb37+drMrN1a4wWGPF9zdKJbUI/rcTZrd61/s7axnB0HXDdOb
DjHpNoG7OjlISQ+DhYcbn7dnM/cyff8YCVo1/WTuBfJD3ETmMHLAQbyDBKA7Anzc
igg/dG3d1rOCbX1Qyu67lRy+rpkW506tCnSqKRhJtAAe1UZrNSlz8QB4ZwF4aseF
BGfq9BtoAFVH7DGfGfC06RpFGyLtiEDCmFPZvujbVKaWnCimub5A8Sheo5LZSHR+
/nNNqooBPejOyvr7K54OuHyS2f7AS90d/enIjwoEOnqZUBd8/Z7XOIIZZ/wyRFdD
5+nAzwdv6t2g/JhQQvYzbxV1BlUONLhNDiW8R3tzuiOfH/9LilcZKX6Mk5l/s1bn
NvxUT8UX/cHQdc8jWjh4Op04ItBKrf6GXC6o+V8c6l6fVGdNvVErG+VEICanjMBX
l/tMOAXSLJlIW7v8mwQPNI/43ElpA08phtYllnGJXjHIzLgP7aJvDA5sUzmkEXa4
KPVLlUQ64EMEyqM8ZgRcfUoCr/MFFP/BCw8VIegx8uFyd+zw9I4IWCu2ATiGFL2D
knzzkfqMsJoR8Cbjr0zhUFHghlp23WtpPWGpWUqACVO+8cH3vjZUN0ujeGbfLZTs
wSpAniKD/kyYpPivNS4j3ejDokR8+XPIQqhhIpXZSFi/Xh5r1cw47pQxu6IRSAD9
eB8xrfPjyqeCbltTIVa6LGilNI/1sMBhxWvrLHMhOYVr/HrC7AqGM5xFRwWmNdhb
l7FLKWCZlFJ6R19fm1v+c/7PW1SbzGhthDZIfucU1DzJBUbTG/d5vTC53tRj7UY7
eYcVWvTtvRNcb6tZ8RicBaO6si9FWbfmlyaE2v6KeEUF1IutRl8ebkP0NoDaNA4H
3ZOJ8YtGorOq93812hrsJi2njvGui+W3lWoVfFlXYEzHOXfkFiV0sSQi69nXPMSt
lqMUAY/9AtkMyVIThyn/zrE4hRKmaQvLaSHFFGIqOZLEeyMRA/QlfMHnKyKtzDHD
SwGt+iia1DfMeC9zjcZQuxHJ/pSsjwliy+nhi2q/OkD7dmnm/IcdtbfqpDuSpupu
8XItQDZDkJopr8nSMd3/TD7eLgcXa2K6QerHjzn9SDMbC/+oQnAE20ZommcTt8Nf
iWANBCQbwD3r2/bXaXI5xgyO1M7r1h/Jp/D57RkuvkhZ+0hV76e9/ofHUDgY7Obp
AGefi21nqW69+bKxdZF+UAghwO4pMbOcPXD8MEmjCXdeen1ZPdCtO8U9at8wxAzm
hdKX6qDhQKfq+rSQBBYiAvw5r/Evs85au0K29g4Lmv9fuWmRtggfI6mVAVr3DyW8
mb8qg2msXoXMhwokqXxAQINhYh7dJx+iIsNjI8KAAYQVZzvxLy/ycyrIQKwemoe0
xGjSrxPZhks+dDmTqTeFphzOanIpaWjtFfRaiEnLSVaFWddoYL46u1nxlDz+CLDg
bkBoZ6k1/99fXYyPDLPELLScluKOC+5YrMFoOWW2eQUXE4DQXUTs9KrzRLTX15Oo
YZblOxEqFUJ+pa8NhnCCBIS7hu4d9BTpRtz/oDb8884IxOSnDF97pAkyvjirPgtB
Z8NYHELrRuHT48QmDMbYTPl/bwC6pPNMFZ4qOqv0eWsezCVFsT8so6UNUjge+2Zv
Bx+sRdXYnqgHkVkwAv8E+xSTlYAD/QhBQl4lH4C5D/f6LaNUl1BHOd8YgiUz87Io
Zmx/X0DZZRxdHO1rVEElq1OkLobxB7SD262NDf8PcuLS7tNg0mrI/4wWrPz3UDbB
hBTfbwK6s5ZqQ7ayqt8f+srjDsu0pLBUbZn4dQK/nyEIjGxBE6dQGWnLiAMSbeDz
UZOx14MfgVek4Id6jWLWkQJAHWOdR6ckXZSvm0p6eHSxYaQC2rrTUJw0/15qFwqT
ba07m9CdMFJFPfgUvc6DnIaQX+bDp6d4lI0kgYLDlbOFzz178OhJ/wk7X1JBcx26
55mFR63JZ+fsrI6RgimDhKgLwa0k2Xa0g/2g9AmsDZ/zHcuvYO4AjKJvDLsfiOnc
yZH/IgapokVoA4lPTQhi86LOVNEmWSFfN+IZ7Vc1c5xideSs/uCpngHyRQoOgn/Q
S3H4ZzGN4k0ZlYzsw3r6NS8HHiGFjtA5/TvaSvw89ePZ4LzaFDIyfWkMrqgwO7bW
j+NTyktd1oEDcNCq4HRNu0vk5dPao1/YTh7fkKi6X/bS4VFNgE6DFxinIh+0Jcgs
EDwHkVeQ7CKTWCs3EnY7xkRGXu4FpbmLVIycL7ZYXONy/G+nfs0eAs1tjmAKL1yY
08zfREPhe88cjzZQi6IKbQF458iVPAgefrW8CNL4/rjRa0mNI2Pp4okObCwyuIrn
EQwNN/KbixKY0PricSJ3YpcCMJTvG3sDYXuaWK5YeSuUTr5uoTqFFDXqSOwF9MsB
vCF+HFfuCEbG8CUatnYgbs3i/n45uAAQLL3HQ++nlHINJIP6uEi2WH+3ktp3mjOC
bhzsktRDok6e5l+ke/o2feXvYLj7Ev/B1Tc8zjnTRFD2IPZoFpQg6/7mQXGRLgm7
hEVc+qT8NfvL9lQdYJKQNJIyJN0WH7nfthVnw1l29A+LfS1RW1m5Al2Th3VSg+z7
0muZJBniv7gMy7KtSBv+HCFX6GYjIT40Rwiy7cI6yTCjtaBoLW49zE599gtlr/pD
CLDoDBAG4M0e/Na6/6bJ9pjmWIWpx1wcHuewtJdGVM9jgxAVwfBbjDANtHUo44vi
pXcayT3cwUpH8uwNPzYk5ZfS7rejF9CXNODtsPyY8+UYmQf4XcpTcBtsGX3YMjr+
AQYyAAa1ZkWhltm71e8HbNbpQBCxK8yPKbZwjB4qxuB1Z+2qbRDYOFwFBBqIf2HI
aGIjQjjxK8JZ8ndTbwOZMQU7xP8qICKJxbviMtJrSzzuyJVOyFLGMlZplwznfjo7
6Uxcae8BccuLeTaGYgOzw6pOQayLejfcIltLK+IeqaykN3krMr4nCswsGWWFamRN
NiMNUeilOtU9dH0GbCqhp4+emL//1M5qHcT4tO6PAlxQQ7EQNHwI1qFwfbV5wEGl
4YlUFzdQq9de0DnyoxXZ3nqw/tiFOGwr0dP0uyxHsZGZh7vqdkw61Fho497v8+wW
bD7Oro+lKJqxPHjEMOyudktvpKVi0aPCb57cICRqllnaS/ZKnkoRQVfkg+LAsS1f
NA7zoUzxpPVev2qxO7m+y/PWu7+R59FGHnqq2i2jtw4mbOx4vcyrDCMF67eX9Qrp
iqs9li1wjUz64miwSrk4Qc/bN4Qi99ynSNUJybK0dy1ULHUX64r5koN1f7YNqlgh
FQ5fxPN42baPQ3lFhgbBS93pMZBiOVjVSg7bykl/WtCEsTtCN1a0yZJtHU5bQpew
xjMIfN1wAjfKU0swZ3++yVZVNj73N1yS0SbMH991KZycBPYBDKXiIUDKx8nocLWn
N7hu7ur+djVbIWJsh9mVXeZJ8h9gMuhyaU40Vdz3DoNERoLHGv/CDzxV/07gmz2+
AV1XMLOGTjp0WTpOn4VOG4XGWaGXEhF1xPuRGrS8QOnSXXR8StIfStg0SRTMXbTg
/RaA7hqW+C1ICkcPkXbvMMBNDLlMZcxPVeKka0LQFEkqAMw31paTIAHN+uoOu2EC
mkYv3MIoMn0S/FWFMv3nH/bnoseAhVhL9kHOWPlG7kwh1BOcn5X89R++ebtMkIAT
KYGAP18lHRLOc6SGQnG9zi4vxlyJvibmf17AWJxQsoVr2upobuLLScBc63+F4j/a
7GnRbKuk0MaMQgD7lMuAG0dL8KuZhZHF2DtB6D6veE6KkNkmDRsNM+jzDXuy8F18
c5aYvLnrjZRiO7iQW76faQP575003e8+oPf1xH6fxYguiSe8nXtl4IwabNi1wFBo
wb7tMbDQvmohBocw22hunMd4rXznnMKhkllerD+ezP2HDDKLFDBBmf/l/44rMWhg
64pGjGVB/l1yjTKHNpjsCCRcEnrakSuy6j5UH6y6YFkyXe8kzqefQMjZUl6BrCLt
BuM32o9y8kcyLpDUhgoM6gHtsqgvNNty8Nhe5JGx+WkSaeQubILPLw0nTY0rrSDs
t7Tn8CjNsbXRtH8SGhV/84AlUB9mW+cov7Z0nXTMxjX8StpJ+7CmTfhBaYZQQ0Lp
iOHhVmdOB6br+/YeoOynTNs2Cip34n2XvgShw1iJZ19Unr2awPULShrNawOvsPi5
2hbAk6mUIPE/g5QnnnyYiSSc3gvEGMSCURuaHtE2NnduNckBYH44f6e4yjDb7nl6
wuAnaFBANakc8GXpoZYRGV7uZGm2bKyfm0bw47Gv+lgg6WS4+mRVdeybeK2oFZLF
Uyk2H8YVt3cL7f1Tf+hkAcvC27+PDuEv37DdDFPQPIf7Z0TX0Qrp/0gy3+BjCCnC
wnYgr9CfmNfVsgL0tl6SX5JoQpEAkgR7+Jv59HTWiqe3TK+6LhxRfMti3saGNqx8
XVsQONcfoVCG94+7i9htmDCCwS+4sQ6mummT3b6VbYqB1vxJz95WS0pvxu37+qlI
+otGtQxSUK/sp3KGvFPwFX/JhZuwYH9Twai2CD7LF+1dvm+mIgUTzLsjpn/Xap+v
3Bf7ofRL+fVuoDSptGwGf8yLFNWhxKYMmesJ9+ZiUpr/9B5INlQAip3aF5hYs1mu
tixyITeQcacOsUXE9lSo+wLLKIZzUys/FiUm8LjxZtcOYLuoLDNdT7tmlZqFsFSP
H/lCn2eKlF4nQ6n8lIJdtsvl54TtAHIfbhm7WvcJwYvN203O9NYWF5HWL/vigbnm
62OnnIKXgU2620FsvTrOkhDuhP25ZZlSaUMhmTGm6WV1CtUJM0+Sxdtr4rHN8ETO
LpzlSllr1aB61kjJXrgED8IwBf/3tTYsV2b3ArWuHfNRx1nqCVzsnAixvKSjUMg7
gSXk+Z0qq42b2wcdRABD45Jr4V6S0Q6y9IhYM4EuebfIS8XQYLj7fNfc7ahlL4HU
vSwkfE88fJzsM/Wm8WiqM+SWyVCCmEpG6PQxcvmHCKLYatY2MnuC0P7p4MCaXKv6
MMqraKfEt/z9qtreHhlY9e3JsKRFFvAviQd8kSQFPZFQlgCVJI+C9zB0SjwjtQUZ
U1YDCB53hXEUDjjkezi9DfL7RV4bm1zrWqPEBYBqByXxsP5cOi/980ENy+AdP0HF
8RiuebA99a7wf30kMd39ZYrtoHws2NoAPHp+lWj4ww4PZGoTDb4h7IdLZj1v5bs/
W3dtbQuSO+P3/1gYa3UXwR9sxc691b+iuArnSotIbvMIIeOuyGyfukhV9S+XuNA2
qtmn8u3d/WFdsF8MfTdqHiwdyw0S0TL3SDNrb/PBd0r3yVi65bA7L+o30ovEwPMn
JeYtEZjJREguXAKruWMkcggOSJACCwwcXcH9Qeeyd/ZZyFn4c7WAfpCzHkmrAIDl
5zC/PONxjAtrRi/qMb5sYb3SGM73RUlkwvuKCkXz0h9hvLaipd/diMP9L3o8Yvnr
54N/A+Yhq4n2hNfgbGT6Du5jyqogHsJSUvS7YhWpBSzcwKGRptomsurPVaTEKrGH
pRh2d53FAfuGR5uneWyuNIw0Qifzqo5NhYDr5q9VYC+CEqdRL8qRPQa/W6hmMPF2
JPBDYhasdtNqCFh0p1oprFtF5vMeR4RFs/jbjcnyTTffClf7z73CVldHBTiF0R7J
FkOiv+j9hnrVRv4cZksDfeDlYCazc0nN4NnfWKzb/2cRMx5WeBCRbtpr/QFvrqcB
ucF2NGi2HvqpVaioWgeOz3iKDV7Gfmz0X+/3lq0rKmoUcUhdkpckCCIeDmCg2Bss
/1zMr4YOaPKsTzdYRw6OMjJO/DfXsR99nhHZlpFf5ZwvLxfAC6CNnPria73D/fQR
MU9xTHsV+eNg54Vnq3VIZqv94f1WBDtHC/V+JxuFWOLjVEdkZrom+Uy2V3JnUvwq
uh2kb3WH3MNJqatjre6XL84Wp8U3rf3GdSnUqgrC5sKUfIVy1v2CprJmE2asNyMo
F+PFaXRJTjewGryR/HS0tSK8GmFXHJGJo8Rpb2YN2aADH5EQawin2s08/YNMRZIM
FSZwhnSp0G9/9ihxDv1uBPcpPHabhEj+3HZO6Fj5AkXuIkkoe9FEk0QAKPyM8w9T
OF7oZg+0Nx4O/uRSmAdoDmAE5PEEuaYT/iCkQf0dZEmbvOdIDG0bi+eWQ1wjz6+W
471acyK6nqmY+sickfL6lL4RO393n7PJTOkwFrFPcS7xXhxqtp7f2XuVd6Yqu9x1
E6Vek9aEpg4Ux0naCurWWPEXjo8aKb0gmltHNiBemGnIJE9CtMMuF03xv0Brc+Gt
6hRDAudCmjP55r8HfWnjP70ZA/ZUU3iTH0rGjZTxpaEq/iGA6IUYQ49WdmGWDW0T
Y0ZjkAC03kSnZqnWpv5OTOvLSGmTQmmupzXK+n97evSgi1ZBj7X98WMPfIWkwdAs
L8YfkfwsW0sspxRYQBrbBrMgIRpA7vIuHlsuvCzOt1zg+AItwH5L7Vq0oaPvk0Hn
SDUBC0MygYo8Xpu18P9ZDPmOKTlTk2kkhj3ACQqPqniOxke2DDlvayaexorrI2wa
4UlPK6dUXqO0pL7MOd+k+WFgUufm8ySmEn7li+NNFudzN2vNWLhkG5Sfn4GlAK4r
Q0K3dTCcC8eLKS/m/V6PFLVIRQNp1cZC/h/Z4rYkKIbiA4cYqcygEeJBYOy+pLBe
WfE6tfGEBzApjz4xnTpZmF+rrhT2JnWww76QyGMJcmtDxUkTVB+JHmLQWN6uOUCI
z40djvXGrkRn+G+5wdzo9aLXcV1dmGSSMhJ4v5PELGGOkrJEXs46MnXcjIbR7ERi
IKczctqlE9ZMscrrNwl8VKHhvOp0ZGyZI5qUPQuere+i3dw7Qlbz6GkrAJCYkQWu
sUbzkkF+j7E6w84fJ6Czb0KsYI3MJVkgnTg4x1kGs9LYtbd7tIVHwQenYAXxtxzw
e/0ftawJHedLh5Ck+C1GKtNrs22YVe8WgUIEAKtDWZUJ/Fn4WR+JvtAm4jcIFezh
NbqX8EdJymykJvdiwDuNwfEXHU6ZJEydXy8h6wLS9TEGz1qzlJzh58FQMIVp03kA
2VhyMlGq3gqoiV1dwRBnvp36o9n6lfPOCdttKTRon4kGwL4ab5/btSSxExYxffpI
+RKcz99xzm6lmIlOWazi1zO7gjlG78M4NNmoAmFSTn7fNRlhuKV9YpJWhEFcVgOf
ydFdIXzpOM32nZf7zWFSoaJtIMqbRQ66imUOPK8EeDhVVMYLbV4vK5orVSMTIW4V
qrO/N7Jthy6wh7HSUiCU7jaYZyVLEfVQXiYLg+kjacmdbBLDBT6OENmbPI6cCkAc
cnXU7e8CgJnGE5QrxtBCExRG6HshHu4NJPKyGFNSMWu2Lg0NPGVbPWdMVDAQtAeP
xDC09RwlZwW6IGdt+NDmTFyQhW9k7XvRpglESrZUGN1szvUWq8/meoWTZjr8jffg
/d0sGvi+OIDlg6IPKEkiCFxI/Y5erRuMBbYhc5lzzWwN9rnCX1TnvKr48WYqHoCc
liFakDrdKnyDMeMnJxU4ldntigNtbvik1LIRlm316PAEO3f7iJxo8CbLleGpjLwm
upKlhZyVtiKAeFqArplP9m3nxWciyrBftsCMLDFQiIu4j2YAl63ZqkSRnGGTPRS9
eEh7IZdm383Wk3WK1qqF7Bo7Vkkv3srQeCAacEbRD9g4zlaBSh7MqGikJUMfmuvF
mILgt6vBGbuJcl+kzS8YDqdGDpGK8OrU314W8FVTD10zk6FPMZ2x0h4LGX/XqHgb
ItOUf6+H5vUdn3ocC5ZXN/RC5WbMBbQh29YrwJZ1SOED7dh+zuN7zquj5ECrWSr9
Vl9gtNHOIfdmYrb+T5yGdcwIClDLuM3kWjYMgi+0QDl7QS6asK3nzA7gDDHkWEK1
NR4Z15IU8zBbPfGKo9A0gWqvEuApusYfQ1Z8ywHwNGoQKZBF/4hQ9qtpVnlvAK0o
jAsT5FkynhKKmScSk+n5IaXgweBlxD/jONs3rtOknKx+4vNxk+VBNv+Jim9vjleE
MrvlT5fbaqXLi5JoWk8QLIRu2dOoYZT6REy8+lYlVKbjKB3diKxw+ePyI8d7K/Wf
nm51Ub1WGWgkEtEjt+Lc6OnVZVdPROiSIOe0tFhxDlHWY9jhh3HsAVcrmzlbritS
RpX3eGg0+EqBZL397k/hDw0RDW1Om23zQojJvzPwwN2rgqcSihkDkXNFvujZH+km
zakwzavoJPxIzBH6W5/hyQ0axvHrSm5vnJEVjKYzipu+tMMCnSe+Q0XVZBI222xC
LS6W3TKPP37j/2f6R1T7q3ozjqKBWLBHW3h9v6Q1cyYF9qYRBdzQTLPD3khyz8cX
3ILYfrfbQku7KNQuDY5iqqCG32QZyhKKzUWX/kxDMBzBBvvu2QOhCsaKtLVcTq2Z
GntJyA6VnKOpW9SmCndERY6b2xvcJp9OQAMeNhJmBgYat+4nsfzXpcAo8lp9aLOh
4y0FxI9rVzeyTVz8SXkVNnyOQ3nfrOKgbcaUvjEigCerfaqmbpJh3D/EPXQaDRNd
tZEjmXLP2u+sVls1vtL0F89IEqwFN1Jk1n9fvLPs2okT/0iRBqx/NQrAf3Uk1bE9
hRxF+iKm/SRVQvbcYPPWPxMkctRpzooeO6PcT7dYq1Fi3rcVggeug4wqOPtxaEsj
K8ciSDPiJpJTTNL7Cq8JWBRr8LJp2Yh4HlFkX9t2HSzNIRoIVcH15osYiQovfYMo
l8jX3ndNDqFgWbMmiZTqre5NT2L2UbW7YxaLiTCBA9RMNC/4GOl5Ia3NVhZ412Pp
pawJ5ZJNBm8zHVGcfNGW6PozTclytpw5ad+RwdyXKpiukbAVjfrSBBSItPt58gE8
+9jKWGG10V8KvEmxuZLfebph5xPvIWOPgAtS+r8ED4csvA7QsSUElIjcnJOgwBVS
U0amOz2L5zqodJU5zHWcOYLNwP3OaFDZJUzMsQZoGTH7Ye5KISR94MlaFP1XWDFk
M2fMy+PFlyHrUOJE1UWTFzve8GT76gMNESoGAZ3ShC0XIMTJ1pnRLqe0u4pgIF9o
54Hj62IT4xVvJWc4IZvzbPv+1Ez2CsCalawm8NT233J9lFr13dZhJs5DY/Xxum5W
MCYsO4YgwexNvmiaajXQUeOMgn+2HS0WWI3F05WToBb8dHrlefwGAlTkPIhihYd9
6x6EV6gYxnR8PxW7pDup2mtMFtlw2WGjJsl4dI+cW551W+MCsDCpIlVpvO+ma2s+
YM82pensFi22PZnCnVs1EdzKJq1c8ggCDcfEBJNnxZ6lf6o2Eb3/AI7RgvFrS79u
OygxiZnARr8mvjIX9HMOGfAgscVgPlLCpWNxSV4qmuxGSgqfiqJn+Rb2T8sn5P0q
CRm4kAkOoIqFNZ7Jkl34QjoHG2dGdBwnAfSH8Miz52u01HGUuoLbpKpxpD5F7baS
uF7cplwswvbhGFHQozkrwdKtZVLFkOZfuR0yhoiktsaAdFC47aVX1Q1pcvpFeFo7
AJQY69N2WR4U6l0pPD3gdN7xfiLmP9OEs4MiUX2Atvo70LMbJcg1qiYYGgsoodLc
Ug1KysuwKbqh+lrMVTWp7ofdXAc1eJPo2q21yLQKWY9NCbFKsM49NnKMoZ2+yxj5
1BDfgbyP7kHiEFqIrWqjFfnIC6L5yNcJCSX4eCXxE+xk09HCzLrwOqrmgQVFKtWy
OEXgV7jlGKGoMzY+Se0NWUR0sTzh2SNitizMC6ki/pIMh+4jkI8wGHfVHm820xr6
1LDpnQvw8jEwNMn3az7U+UvPCQhIwEWLvuyVrtc15hvfx7uh6tEV9+OgSfT52ZN3
mx1OtWF+r6KHkprLMCqCT9Kk9gERm9IMWfI8Zqch9sPMNfLIpVOh838OQa44VzER
ZJtGgHs4PuhYEEBdpi9PjatUQFpnQvy2HIJnYGiMzwb13CtpIiCHIthJ1mbid3UE
iKK5amhsT4M/dv/YeqNQ3W0yHpAtsIZk6g47I914C53V5K6YibxSeM47GQlZYZTD
OcEUzOJVyjJJOLrr7zKV226Ug8Hp8Vf3OxgQVYHdEWc9WEQN1V5cq/6kTO7qQQ1f
J1GthfoksM7ye9oEsu/Bh0/8fElRCtuOjax6mHK1Av99PkSPdD+z0pq/0byQqTmP
rUlztUKMsTtCHWEId6cxnrum4p4ZBXWoNGy3w7XB0s9zVNLoh/EbwHxL/FT7AxUT
iOUZEk8XFBXkwRRH/j1As+IBS42tjw6yjS3ABwvWL8PhtgHbIuJOC2PsHu/DJAhp
5xTk6GUIcrlZIxeT0/95dXbCmnKHWfieozrkacVgjfo1BB/emSpveixOs4KyPC1A
yCkoa07IhS3XSUPm/B58FqzPeVoetiAgdkJKPXHkz0ECy+OvumOCS/BOQfYn+aCK
CcmIQq9BGrX2WG6VLKb9jO3pMsCU7c4eWGniPqDwhxvTqHwYNXjKONKmdMzXiHuu
wNt69I16KOlHcyPwEKlA+cjrNkpAvOUQwTSar3/lRdNQkP6n6nNw0mNbD2C3XBfZ
MDca+rK3R2gNkPrEGw/+nL5GPrVoAPudjhGA8Ai/54w0mcTMeuMdtA5QjKWbyZKK
ixIkNqCwsAA8F72u82HHicPMs5DmV4qW8uZUJ//jiaRe8hkvpPFeSmKLMpvu8GJm
moTk/XC0xDA8Kbn2T6Ni0PSJUVQKuaWqN0Tm6KrPZPt2EvY7TOBpLnHiQMn+FTCg
OJPS3Bx5hKOCCCt0Vup14OzbBYd9sSJSLXoB7WS9xWgp/fvbccdbk70ui6CQdTjr
QACpL22Qp97HjlxH9QI9VsceUtzOpPiR4n8oUac4J96PS958MfYPfQvJ2cJNprVr
boGSvEOVdJl/jM15HJriL3J+KrK1QLegZIcA+xP0ZBNlm6WmqDkH+ytEEocrlh33
lxhn53QA3p4qoQpzTHZ2JsDYEAJlB4J6ccUaw0MjI7u3d5opNwcE+Ex+oBSvTuzH
HPP5454NZQmlubIrQ2x8CsSe2/yHS4U3rv6+zAUGNV6Xp6wiAMsQ177rluvZcIAl
WvPIp9rigCWUPfTW9krfCxjlZqHSRWjlgpAXiBuFRd5nhsXD1iibCSbOJYdy0Wl8
j+boQ6EirnFFlAdiOhIMcUOguEoJUc1VAmuq+3p1ej3QGq3mKW2j8G7iIC6O+pF0
eq8DZkkEL0l7l0qNPgvS6BJvhyXe/zQ8mMsq0VuWfVd7YFwvkSAKQpNJMhL9mA9L
+7q9+gUTZhPyLAidEKN7iVyE3fT4nxUBBEZ6frX71R/YamGRRyW7n+gEE1X200gz
4/d3PVVe/tZZGygg1ejHQVxN8p3WdkGLHwE9jJt40HtyRmu1skf9i0JF6tcnI2AP
y3nMyCBE6uESm7wTQ5W6Wk7IEakkiuKScvdv8eYtPjYH1/Vr7FUNp6IlrfKt+USO
da+cH17QC2uPtbYh8OLXv6jkGVg2M215RuoBcqnighTq5b/XfKrL3dVhV6f7qVCs
J2gSJxhaDGVplsjVusg8wJRSJNrsNvGtI+dH2CkyxsPLFZUqMYDU9JUyGiHWm2ap
aK66Q+7oqPFX0il/+xRXjeIstLDZmm+s9+BFSKUMncTq54iEbznRR8CuRMGlU2pn
/WN2Lw/AIhCPBydA1VwD6EONQcTgsIKe7tgnLCNMzTDzYDF0SObg3o9f+Pizvj8j
dE79BHLJa6uMUuP6mW157ZrrufSt5PHe0g5DJIqccDoMAZL44yb28tYP2GWzpAI2
V30WcGMHyubyIBcK8So17W+v7effCD0hybIbBApP1IwnYHlFRV/9PaqBxxC9b3Dt
RxVRdPf1PI3wiKQ3mX/9cOKBpP6/PXre+MkuOR0Sb5kUDbf8G2iJ3BLQ8rYYYBts
UWriDKICbCjrtWofu/ukbevo41970F4SqG0RVBi48MgS+/WXyxSgk40/MxWLtkcZ
AnhHKVCWchRcmYO/VBeqdLQ2+1xzHk5BH0bBf9aJlATIkueLU8vMv2YbTHeGg1WN
LqYXAdP8wRbfMLvtyqYQ28gisYETolUFfTJ08EO1e6wPfIoyf9NpwyUMgLspiIWR
vssTY3caf7degaz5H+UVFXX4fWosTsqfFCqHQhLPEEW653AWbk98uocYBMEj6Bvr
lnrJ18j/LYFAQG/7W8sIyiNLjTihwX/NOMLMOJukC6nrde0l6EEElzVlw0PlQ05K
dKtM1j+0ZEmwKjKNRw2ayo+OBVjiHMm0EahyTYhQSMs4kgj6qjooZ3qdi9nWte4l
nTsrqEtCs2tRZY48Gll9MgNmtvRcu2yoz4hOIWROQ+hIxmYa4KQpptkqhwNNt0Qy
/Ow46a0eObnLu7yHiVhUKzlggzYdxxTAYj0gDDzTZ0wwF1biq/lQvGFiIflYM5N9
2uM1epI+OSyIhLwQFgN2ExHArIUAtjKtJsPK4w+AfOgenx5tMrt+HUl9/RNRDAls
1NMXcPK9zpAVdENTx3eNy9VODmsXdLq7VSVAmBHOfj1A3acnfmT1ieewZbFIzpuc
ZE5ApJcOBDg/+9GvPZiuAFf4doe6F1bHnTgRez8edz+hyLInIHu92uB7mX/UkvzH
KGHVwLMwAkvT1CnC/50qVDah9xN/CGynApTyc7DIlCXYf8oIqBcZXUM7mOj131Q7
dPrkQZlC1/4xVx7ke/c652KtxN5MvuS+Rsg2axLSQcillSemW1hKWvJaqS5xkjhm
aSU1RxxeFG1Q6aKSXukZuKM3CzR6y7HtHlvzVOMjQZOlFqRowTwda/Hc4wThDakb
k3BxZM4j6M9jWD1tjEPAonQKXM12IeUSGUav59hoJMOtg60F0ea0eW8X9fjzGtTO
jvz6DKesC0/UZ8fwOB3LTAFAfjTi3Mlg6ZJ3IoH01DIzaePnCyJsCXeIE+rpa1f8
P7KB+5LhuuxqWDrp8u4Kvo13VIWG/wMRO8F4BECK6j+3zbFH7/FpHFU8VYXVLa9C
N64dmgk4ETncPOJYwt1vc/XuImlgajcV/ET7hfl4NxQPxhE0CBsEfIFJ4ggdP9aT
dafMmy4K00MkYr0Llkc15w/TUowls+gWDM/Lk25l3kEX7S/ZypRsCNK5gP7rCpdS
Uqg4LNiuXC7QwJYbREmilO/cAvBOCCjH+9AcUMX9NIwjOyvLuStnOTGvfcj0c0/e
kivLsbvSBfoG4mt8djBMTzhthOn3jlUfWxZRMlqMLze2y3bRn5Gy2AFuFOZnZnzK
6fJFZEMm44lF6jmoOfm6BeT++PhnVpmGkVF8tkqG0yBO27LZYYfUF1Tw72FBrhK0
Yp1a7fGNcJHR2HC40OGT8adTO17X/GlANQQXXHG+3YiTXRDSN7Lft2LTkNfkcdms
TgX5S0uVlfLaZScwElVofCgl7YGmB/ScCh2DC/srXFYvTgs5BFef3RllRDFvim29
fFmcMFGTHlulhtihw3SA2OWQ6VWuChd31qeISCEAW9O0Vz2hiKh75m/yL60d6ld/
Fe8WbIOZ5siYv8PL/nXOA3thgpV76oQAT0IYIJgj+uRRQHzBtB8Qun94izBR/mzQ
/BrMbyMCg9EahY5CxlRgp1iz9aNuxCY69g0VMNQOK9dVZFEUqERITGriFQkDtNK4
0loZyzQmgZjC2q+1epriAOXxYLfx/ROK28qKIK847haWMqi3dDGSCUvkY/mQCa3Y
PHj8+Xms/lr50N65tuxZd4gGYK4vs9NCtgwok/KCZY3JdBdA0uuyqGLSCzwm6OXT
eJfeQE4am2ol15liI64LQm23Tcq9y31AGopgDXhDDACkC9gH8lffEKClaN7+gADc
k4yrX+CH2zo4Y+9bUG4VQSHupS7MR1MwMaMZK8I5CRC4M1jB6XPM49+mFVLSR1Oz
6syy3i+nnT3FkFDvSaCVc2pUgOVOYbIG0BJIE/lfkLW2QiWtlrHllFriFkrFjExf
5R3JF2PnD1kZAKAZ5TyEarZBakJi/ybAB/CqL0XOI6pCkAKDs8FqBnQaGi9yYkzD
VDdLHbyGVZg/wd4jlNIxe8QXG1Fp5rJ8ppZQgATxBNIbz0HOLr7Bk2ZaZluEcoG3
ZCf8kcWUNIdTiCdU9q+d6jNaVEOXb2nPYRJFRabTe5a4nLV3axL6mZCMoVULwjrE
OMXDnDbgd81SMR3vqMtiI+0E5komJd+6ABfrZuSJ6uSNLysr2hRV0odHwsocw0PF
lR4tKRnPm5CACOxSqpusn3NIpnEIKCN3X54UkNOT0mX9tINdjp+pP7Gjj7gbSs7P
i95+NEkj994cDzF0ttBxBJ9fwym76thW2hdmvnH56zsBOzAyE9oN9wjwPdsMWEIV
Nkdqbu0qJTckrvuO2I/Xql3Eyx++KWc89t9v4iOW6RnXOyRPeCAX5PXEY+4Q6QfQ
8PlTm2BizIZJfCMmFC0R48FVGsesh6aC2apVHIyz2mneZb3cD6Bh6A1ra5VHyCqj
jomEWufhB/LXf8mfMfo2GH9QZB+ycRJvYS5M8CobLIdMz2lnUVHgTBu65mZSy8tm
Pp8+VJkOxmt15yq/GYpFB2tBGaJrtSeJdAtriasL93GB08snIkx4uqueCqs6lCQs
h1Kkz6I69/EGEWoJ9d4t3g7Tz2HethZp7fUqPRrCBPGnM77ZnL47F5/+gThRwso7
p0cKhkFN1C8Ac9W8fuVDD6W/W3e17aEU7YaPF9gm37m0fUZxb1amKSuwhCvMJLuA
H7r3dhMGS9z5ZMPbpdat++ICCCukGs8fU0ZW3pggoLWBRBh5u0XCrGffnpv1VNdV
Jp8vqLnQumqlhLtJu5VmVuKbQX1gTmbmj54P6gDPJozRol8BENunMszk7WIq5J4F
mPsZxCLbJWX7lhxOFX0lK2vagbuCxCVrHCrTfcVkFJrYFOhUw0GOnXX2CUGNlATY
Q1Mzd8PwBhu6kIHfNrurx9x4ZtpNe3eYyUBapQmeRQ1epyS+Dldi45DkboSwjFln
ws5z7WRZCzRexhA/E356Mm6/8bMdi2ettFJQiha3EMmwyDySiUDVMNuj3Q8HSIG5
fUO/R/dts36bcrsg/hxNElrrp2WzLxlRNmYmC+8atVelqS8hrgpPqhlmkm31HDc0
QzWeFdaBnzCty/qeN2QstMoaNnHJrG/jAF1PFCOBrhieNo2clreaXGREWSwl0/aF
EcHKCXs6y1KXC+JZEY3wexr468RJ0WSUz6HtUnVxn3vLutDQFORWkYoH23OreDiH
Bx043h9813yivmBJ1twiQnCAP52HFQE+Drfdn0ygbt7jxkjJ+q81XjHWwyWOUFdU
WQbkJBECNOcnZLkrAArUSxMcb38cIl1+6ZgMw0WYV9yKPsQx+lLSC2WP4PF5L710
2CP+1ac/SH5JrEBRe4P7tctSc0zvPIW7FCAzm1K9QqRNF85Clp3F/yMXitDWiXVs
wnRSkpbKMv1q8USh5KgbrYDLTpU2kqVghR3X4wqdXDOWEKj+KJ2QN7aKPiPCxNLo
8uBsyQOqVphTf+pts3DS9ja7o7duoMk4v1MB+OXuBxmwx8rgiJ26v/nKunG119OA
CQ4LcBLaHGTEGMCIUaWtHQ1KqAP5rqV2xgBTygoRps8yw0cn9DLgMeywx6v0859A
HzgpPiaq9QXDJUkGblj/shMH04OivvsK/nsjOhe6CVbNjZhQ6w4M8Aq4HFUxFyVU
xWspJ95NNFNKt0yzKOAxiJjcK93PGtwSE/x/eAofHC0n4rdn8omi4kuoHUe73rIm
0nIIlmvK/QBztWYrBAIofcoLACUpHG/MBjWaGMhOJ4ZmNcqLYZutiFJYpL/UgRfD
ChBTJLp5o6ILdNBUwHPLiq4ZazzWa/9aVxvVWdVSmJJUSMMy1QvT+GlYsIJ577y9
C5z5iy8qdd39WW3OCRfUxyEnmr/wbCJhR2XBamEl37VS9/QQjx3gFd4IRnmGqzc4
zjK/A77/BD06uERkEDddwweZHA2tJH1Oqf5ASSI3WaOqj7yCrzs5uoj8JcGQXmw7
JYP+vTNCyMbr/3/3964cOqXSDg+MwlDs+Qo3THSivnxSfBhBnk55h/eIlp4VEqsf
lg5pM04bQL90862c38zNRj1UvWiWaYqrLkIAecUoEfNP2aRt0tSwj56pvWmH0Kri
445Pwi2mgsqRpoLAFOSkHNYLZmxbaCrsP/lI29NOka2O9HX7zPgeh758jTmZLbmf
u/Y5XHCNmzevE50OmRda+ZN0Et1sL+I+y32aYqcSqTn1o7Poo1CnEi/2iYld+zyA
rqtHktzSVy04pdM1hgqjFey701DRXUD7N+BiKxUX6AwmkMkcmJ65KfYxaTY6nNKZ
AEK1q93fBwkuAhJZMuoEXAFJdky44ITAvtW385DAuAh1x5Sdz5BkyhJ3zlA8k7Xf
f+6VvXVyfJ8eUUKJal4jnPfnocQu3oTg2Hjup2uUffToPAEW4Dny7KtH/9RTXE47
9+VCLCgrnQoqq2VCfCcv7o5MpcRkJ7Xl7tdOLAJOdU/HmVmz4DrLeBlxQvuD90/w
y0SLVfOOTjlhbTRbnkHK+ReGgiziOJ6OUhl8He288xMNUzAIB5236HnxfoE6huYP
X3f4xFvReqPE7lQ07tuMcmoVsq6RH5eib+YdV2iAR4sSawYJJZOnLDgptD2Wc+CE
Xw4D9rP4wfvzn+HXFzKA+9K8rwLAYhqEdtBGvId0Jh544fUwGU1F24qvOdCvQIKB
Z5o2m2/m/iaGEnsNwzCA2XfTlwXyJ7P5O/W6oDoYko0chgNEwt0O+Jh02RaPfPo5
v++Dpl9TX7yme4VK28t97xrTS48apGnzQ85LTTEl97omD7HN3X047xQ4Gs4aUvyF
DLWRZIZJ3HV3LwROPzNvmcFLYVSbXBpnjZdgZtElvb50vfsl6AXQI6/gjHl7bN8G
8enf/BW42W3pifwuLX+pGfJdxdsGTuAGMTfhOzz0DDeCMP675Uy1nre0f7zfQnQY
tYJffz1g5t5pjhjs4MFEjYsp/2stQmenzDjOrjH15COD4TXCty7yiLMwE9LGN/xV
XVCL4Z3BUERIQBsC7sAo5zCDF1iZ1PS7iTKyWm4RlcG/3tbtn/HojyJDrTYH63WH
F6gDqln75/i5WrKLT69dVQ1kwTwFX4v8t9L+62KLpNIvUqB1VisLzLdv9//K9mrz
QwAfDNr4WJoYKBUqvLCLR9UDlPLIf+FkOv+JHVRvcXqCpNVsirvm+dXM2bIMluDj
nSmea+cicBUAjijgU9XXskb/4wRVvKJLHgD6fY1H09NBcS6FwlYy4NlIcn+Nfee9
xJIHTc8ZudUAL3LNQg0UkFjtwhiX0EtFMx5r8kxyEhIQO3za/aFszwTDesHPDELd
6gCh6VXt3R+Pg04YMcm8SC+OSB6a0pGk1DBR8+Y+wpghRptxqRad/pZbYmELw90G
iguuWykk4bqXg6NXvjin1nZpgiQ2x0iXZomqPOtDsPotAK5cRKqLkwfQrIeYsRzd
FMd8bh93z+nqe8xZ4MXbDzPDYHJUQIAiD4ok/NgJ1d9+k6NZYqpohrrN7shT4Hkc
SFAMvj4UM7jD1eAsnbqVemhqWiGDs7R3u46iqj34ztUioIMA0n/NxozNJoZ0nTV1
fSqURJN1z7AQoOXVuYZ2wTIYU92qyNas4jT54eX+f7FcFpPd8Ax/F7sH0w/TQLaz
Ce7dn47oVm616aKjTZnsh68FaSNBX9FYVt3HtXGgPJQwbgWLV3V6eZgiJ5X33o6d
en9Pfwus/3r31PMasgN9jG9BN1PGX1ifjtR4YevV4KG8R3E9VrGd8lPyhaWsPgj4
rubEGMuTFtXzqTKCNsppu/v17aLtBTj0aQqGGBgOg/GE7aUbrGMlfsKxIyKfIQwU
uqFUz9MHOTOyg1vjhsagLjeBUliCeWo3HOSgJM+7v+OOgIBDKbxaca0PIg/m0Ask
Jlfi5t+sY4hRcEM7j82vMKmUx3cLQb4Ck/hfUcefIek0scVrxBMsmhTUTkFI18BT
bm6CHRnW6i01SYw62ZyAU5b/WiQVympREfHoAP449129vqNxNR9+Fo9ovU+TT6J8
5p86oofxc6OY1C2zIspNxmO2e2OycUgKsQMDWsvShM8C5ommBgqryGlETEbPmSRH
R+8zh/dgBYnDtpoMjjdhJdMOdCBGBZ7t0GyM6cs6QGm0nrNkrwTgcK+PuC2T9O9i
kv7/IDocVj5Ny1jxo4sts4MNfZMS/Xd6VaY7Gh6jH5jatQHKE4BRcPsbTle4JL8g
Kl/rbKT9AIbT4EJUX0Pz0XGa8SD0G94NN/RE1DZiwvtV13la+VyyD5tWBS2Prek+
wmGdgVvISEMn8Lh5+Yek4Pbt0aSStKcVFyQPg/FYq/wBNToe260ZeK+pxJ3xyr1J
X47X4PVuH9Jmoxq6bPGL67EpkdM5i4Ka+kaZEK2u9zv25s3JPuysy3FpNl+u3cd0
KvhpXsGVyLsLLtRBlYpIDZzSdxlMQ3YQUcPfjGCWGWhzLvptzUMaXzsqFgj7KL+R
1tKnAlT/b8oKZT4fzqfuAG8KyDTvvRSrRACCYCIY+Bq78RCvv5mQ8So4mv6xs/+0
LEwXyskRuuVeWdxR3dPfDM7ObFVu/rj3d9I5XCFThyN6AN665kt5e4VKugPd6cmu
mG2dhgJp085NQ2FQ6WA9sgWEZRda5SiZ3NSmHFFRiKbk/B9kZ/2Bp6wLAUaEHXsz
lLKDkWKoWEV6PfncqsY6SHMSaxCwcWvGKFhMSgCbZLzYqhXYmyUGgEBoAi6TYWKx
VK7LHu5vgh3bZdWanzW/pAiGHwmjkTjG/rsaQFuliaNOMtqytm+C0ivR7NkrpeQZ
OPjD8CRaNxfFG332rrrANk+koneq7r46WcFKvf9gkx2Z1XeXhlOO3QBza7DGcK5m
baxkChYG9RdS8ywK7fNJ1CzmEFnfvn3K9oDbFjVzDWbJ6s7CHqg+LnvK1VPtd2Uj
FAgPkcdBPYEZn5SvJg+wXrmA3Jm10gZRmfBSUz5mwyUnUkszH1+bnV6hIxUoshtt
u99284rwCvlpbJTT9FwOquwMnx96yZuFW2iWwdfxS8EX3b9F6D9qXOuAqeCXiv+n
rvT3HBTfmL98v1g9aSfdtlhpWf/GQSnTZ4qtTwA6gb3WkfCK8OS7HZFaDPJb2FcZ
d5YFnFAKd2/BhdPBSZU2IZeCWgeNwMYHdkNFSrBHbakjc0viS619Yl/bCfaXdoP5
BEJgKtFFmfJDlam9RbW3IR6VSoFQcDWhK6l/nT0X+Z3p1Wgq6ey1n5rem0IVyCuo
VXwoX6GxbyTcIcGZ0YP1VZhaeoz7eXgGcuyJm8GNZoL1jQsfo+4yTPS6jO5YCEpi
Qk//VZHZw7Sq2aYHcf3/m+Ld7pXateIDEEvBg7x94Q7qhOH9BMyXZ2wTKnScFy/5
zUh5s6GJISzcCubj6N1/Jlcsx/ayKzvpu8VlyL26HP9tMIFYPXfSYDLryFnNK5Jn
rKi9NGaN0ExeC4CNnOZL1b99M0lJmTL/ImM6Afi4G+5supQ4KKVHj9VgUX35SYBF
E7leSVpekDERskbKVKW0TN6ItPzDq0OptoOX/SV733Jj92lLV08/yWVaNT1SPmmy
mrZClTbd+/AjdLmLGoGd7X3cyCNkmzfUM1KYg48qLh6mQBMEyLHpZnV9if5pV8sH
OV7YPEvjGuUfJdi0wjMWPXXiF6UCfTeVU0pp6gjXySS/gDSk8hoRvRp4QM/TGyNa
ZC5qZJtW4ou+u2QoHzzCJ1FPLzxV31EP8sREFqkDhtBPjLNxkpg/UoO3JGYSV982
MMd5s/00pEMuO/ai5nZjxKIgx5aJNvi99N1ENMH+gPvRLHLvarBOs5IyvwHP3HfR
DWhBN8dFdiLBxUfJ0N9pPVH24WaqaPXbxeO2psd0xT4ujGBhq4oQnAZ1br1gEruy
g+rWod/frSvxOfr8IrSsLcE54oaSpbkaHjG/XwWVz2xn54RLj37g8Gg5w4TPXRU4
lYq79JonotBgB/dXE9ODxmrp4u1t78Mw2Js1ufeqLBhOSbmxncd254Ckpb3IuYsK
Ld4Jy8eHQZOCHv91lTo42KeHH3csZkWmsKwLLQZ2xjslF8FqfMNE7l5j5o8Q1NQk
oADjY+qWwhB4VEW6Szlqmt37UiPBcBtmGlgq6K7aMCgiZ5bDgQoYnEfKp138xpFs
nxSpHy0xfup+xSwW386VYQeqxH6b5MMxVcxjgfAwT9e7fCz+HWzwabm4K97474kM
D9Zgd/rTk4tPCvkUYYHICKtPWOQq3d89TIbDvGJ4XeR4Ud/dTr8rBsj4LBNxp21J
ooAfpjwmn9axnxofsPBfLi1uH71xMA72aNkpjevD73EOtJMTTdHhwpXWUVyCGYOC
JcVroBzxyoT+z+SWQwVPfl5GGESyXKCsaKUjU5QVWVuazlH3acCCAnt5p+bFt5e3
j3VxNMbNDQRH8S4IN66u8dybILwA/7BPZ+Buf5xQDVxG2LRmShO42jsyqOyPt0IY
HrDOiiw3F40zkdAZSaB1dSdNOD6i85Tv9xsnryOUT8piXu+sRtulD73KOPNIdoaO
u4lH9Id+W3lilE8k8CogFBkAqfgdCsJFahz3ligiqzQSU0ZcAs4OMPKEInY0WgUw
YdK0zNgtCVONf2fnUfDsIYDr3anWANFaNL6QqQjx8jMtxcuyx2dggb91ELKmU136
yRYbqLsf6d4wI8qRbBabWaffuvLYvCrkfBjCzGA67Bt/Z9SRJ+llCtJcke4FabW3
3CPNkR5aJ/AI4idblCHF0HijqTB+iV87qR+d8M+Ds+dV6HjV/4SkqxctlzvR/HW2
YN4iphz3szIq7Z4p05HjucFZiZxZmoprZ+Kr34n7DgWB61pqmr2JGETOc3rVqVEC
LGt421LoU+MjZNY4qFU1LLs2jaSCQALPkRFQBfQVKT1kLHecsOgn9z/Xb+R0hzSy
su2J+bKxdBsbe1yHRIAwaFrgu/9qMXxd8xFz246XBvapw/LBbaP/uQz2ON/fSRME
lTWQ1hd4WyyILyv9Yue4bXavkrITgr54KQJffrgI6dRCCIMzhnV1HeNQ+eEAnqbJ
rImo0DE71whzG6jzQQ2lhqcKd4Fzbshp8KBAKCF9CwvCpSKr+aQvkFCyvvSbqDat
FVTG13Ofov6k/sBC/o5PGmzalDKYBDgeYKU7av1jKOg7SX0W98d31NFsb0VxMuMk
hUmLen6WTS4NoaRMbf/KKaWS71elTldwxVoyBzfyVtn/x/xGYnRW7kX3W1VjdKb1
lcWtpY/OMyieQ5RF8Jb8E+/WgaB5g1dfWugZ8Xavdv2L79jRLuP/QU/k5d+j4JOq
0iT1n5VEU/OATig6ed59zvGZKKCpOljVilsvpH+hgvdFkoncgHf331pz5Nltl5uk
8NbbngicDtPFEG4vKfxp2KtrTssZDhDG3KZsXIvmB6Txp6Mh2HNNjrKi7vt69tip
9LMxVcgZcvoYBIDntRpPkryrblBRSDPWHWBuH95DyqyYExRpKwnBZSzp6eW1iTIa
BWocRuq9FDRZvRLm7cAa6bL8puuHEDJVrkCqUPYeDlDZVf/98WqnccSQ47DZqHvT
FVLYRoIYVEfrP4b1phZcn6KKf4dLYVt48iZjfBFg9+RbcI08n0v4ZlJCBX33z2W8
Tln7r2wLH1Meih+rUodNhcb96bZfBB8MYJzs/eLQ2ECOq8DgIqZqP24BAL2iy0PN
YxGlExsIWeH721c3xZZ1AW+f5I8j2xw/fWSev6pS+SUG6rGVj3c60DjOfh3868ON
sVHwv0yWNsENnxjSu2VfDsEIUkwheO3IPHoxKhiXLAKhGX/7L7dFy7hEE5rFV75z
PWm59IWrQkHumfJHiyw+o/hNExUtRK1zyc0/hGSvtZ/Fq2MKAep7V/hI1mHGy8nd
uL3chVud6R8+nMxjMY6YEnN/GPNgS/+CvHZjFHQt/kVbtjZBN53NkRuIl7IQ41Tf
v5qxWsyjm6XDLMmkRhNAHTpTSYHxAsS2IX1nJfHYgJMyqUXItyC0C4GIo8clf7Il
8YKa7k3qUjwecTDDo7sPUZfe2Pegja+f6o9EDNySbep3nHuC5/wyWnxzX55peszU
MuhtWSx7mpqSVuOX3XJRbNtin3HybJKisa3z4/8J34LPRvu52O+sugDbKVMcZFCC
cnAEaip0obQIwyH+osQPmGqJI1knTV1unIJJqjBbbcSE8QjIdYBSNmNM2yRHilfJ
hAp2JFNNcgFP9OKG1iiP8x+oDVGwxficzgG0lfB4+SGqanAe3NNGq69NJ/p1nLID
KB24HbwkW+Va7sZccYeE3drnR+TbYNFc1H8tfzrvGPHL5DABS5+L5j2LN17P0T68
AK1NoMkAsVU8utmKr/mcv+A2ito16rExdP/2I+1INdIO7hpiNQvBhvh93X5OfIUk
orm1tBw22G8bcUx/1yvlHOCSnCCAX1SlPd2FOrWw8NfuZg3KERcruSMCfUHoSXzE
+a/MEzb7cs2PzWTasEvx3hiHTmTQwVrRqq47U+BuAtMMnLNsxb7K7CPcKh2e20Bo
oIGhtz1ACPPcxW/l5893tEMKCKbEAMaqZ3mr8j0zP+Mb1PzoYMIPvbN1hKMz7Tuq
NVtY+VZZzxwpLijWI13SXKgte0m0uIFoyJd+je/EIiN6UB3iJq6KakPrZTSug/6j
GYH/3ZPOs9rprP1k+5vXupEwDI+iJHhIc8Yrq/ylTSwAuq4EIowz5T1tFt/pAOhi
ueKJmXg2qxX8cVyhSY4q1kl8MfrbFR9UcDaMBKY3rra/K9Mdpq2cJrmkkfQ2ODOD
Kb6zUA1S+UurcTkzA7j7xhsmgALKaSg1Wniu/LVrKaKTiO2WfQLliwZOLqzv1hSp
wO0JCwxtsnLrTGgQGM605tTm2eJwiiNItQURSaIqNkzTgIPDXFo9e0b0ddYDDud0
SWTomSOVqFm1t9bkTfEsutzLVO5Mpr73eJviKz3FzsuliUFE3LQyVZD52c2lzpJV
fhnpK0GWYrl2U5vYLH4QTL/r0IXgCR94PoihYVrnN9cyDGehe06DBa0Ol+FCCVgA
YONG5YQje1YjgLszCbxm5UGephg7H7q5xhI2dZ3eoU4iESvwou7POQ5p/Wn44zwR
vzAUc/FJdRTnDfOqKJurs1YF2/gy10ZX0IAY52ObnQVT4oF4OhHPOle4ZHQg53lF
6livUEKkrweikww30BVGvjFxugGe9Dj4E8n2IXoxPKNQsx7ysPrZzvPyJEMUUW/p
aMlBzdSvdLfInD7B27nsww12akjIhetR2BUuSUYRfGJ+pyd344QHW7VIbHBvKNWc
u86NaxSpY4/2VPVyrEslTOOmldDVyuf4P0EmZVT+NF1xrq1m6tRXyMdwIKHXcXeg
S2PZJ+xEg+K+OPDg6mLljSZXVneWahI5qdfm4kfIKTZHEgrIiyBD8uY0Srgqffrw
kGf2VeAOZ0DWlZT8IIM1tYHzAaFYztt+nQzf8I4ke8Gs0JH1utl2sPoy7MHTxPfi
I6rMGmSDwjMcPgiQpJWsbH5WjG495P/C4fmrPBI9XxR79lgEpWtM+m0JDOgYle52
u488CB0uoAPjNKttLcONW9mpwlKyf1WWJSj8MiswV2ZO0Ih/zIxclVzirmQDSl61
rTJL/46HOugJ9O9ez7VcW2zCjliwp0DPOsZLpCoaQZtoZCBCDebGEx4V2ctOBXg5
8Lv+KftjY6JauANWbmKuEl+s2gD0ppjhLxmXpEJHndRdkXASg183wj1S9XjT9C2y
l7RufzmFlpp0ThlIg9Y2BNp7m+UFJm/9BMGpOF6oFxEOA3izR4P+ws7Q3diZdvms
h8H/3WCjLbKfF9SahzdI/wL5uxe312qTkokWRfK8p9qWAn3FnrF+yCAFtGjKR+hw
3aaM2kqeard1kT3B8cs+hc8K2falGZBPnGrXOqR7IfRxntr9ujOEc/lXDfA2RqT3
TRzxCdVp68pcfzlmx7oVx45hD+Q0e4B4yjxZ4RptkL1HAJy0fZMF2IfzR23abOho
uyZMfOupuhnhHSP9pGGNfw3VK4EntJvFxR9AHKcuRYs2tTZRG2I9VJXB/Q6SEJZc
OkHkHbtkPWrnNrsuB1SWy7w2KLY6W5TWQP3R4dV1O19zyoq9Zc7agVOEf80Zref8
Ncfp5z079IdUqPYD8xiy9mOAEomPGNPsPk7FaOaN9fl96QXRuWPjvy1QCWXjGILN
kmmPxIPyzmPoCIDRWl3ovdhCVksVKeInZhbQ72rp+j2d1Q3WJU4C6LKuebVpO5Tx
I4I3u+FCRefMgKUmSzmPrQX9k2jWYezsjtz2y8xAN++5E1EgupxHumtMghM+F/F2
b/jWczQ1N9n+pnAj+z2VC1zuCdtNsHR5hvkbgbTxTrNcM99bQgg1HtVy1Dlsezr1
qIrZcY0d8kuPmRKNxnRD+DmoQT6jsh3e5RemOGsqbPLdhThTNTYZH1d3ncVH0vwu
FhV6T8REGQxWx2DN/vcgrQjluJ8jgj4on8oUO3N4kiXjUl5TP1PG1ERKWo6i4xHP
NYlyYBivpwn2u7VavrmKhUxtJXXA0gE0aVDHpIx49ZBKMnRzJZZWuTrYK1g608OC
j86YwiLmmLyICFeTxG+LQb2jcDBnz+H7TaEcUv0RTobTX30iILFYgSduKjelklH/
0h5vt3O5hCiG+vb4K2CsW2Cwk6yfulbo1gdDIah0HuiivVxuvM3/9ur45I+NwyoA
csu5fazwstM4Axd89Ltc8yKM6gCrq0fjECOAUw+0Kq0bdPY8Cmh7gtBozegZ72gV
V1gOoEWmy2SfOe1+nlTRH6HFBKCwGu3tum0jwssYzzOxO+OZKi4HMgYZGjijPRqO
QSU3r4KQsHVZWbLnNqumE5VOs21/ZVvF0hmRMo8nF+Zfz3XpyDq3PSRXg05ocLjq
qDPM3Mn7E5cW86tBh8m0bPRMxZiU0xfk/xWocg98Fsdrz8msFHWqXv+Ii9M3hFo5
2juHFnVDgpeuBIZzjXQK3BfC2teRnoeApG2UlYOo48BTsk+j4sGXEC1c8xDtCHDF
HvpsxJPwqgAoKSvGrm685QrjWF+ODWsuYEsfQnwfBkE8d4UMg+ypouc1Gjj83x4r
TOl6qaHVoQuwIVOJaNFE4lstd7kHBx8zYZxyUKBrXbTxL+LOMeUmeRC5HxKLTAIK
2nx27oaNOco7fDDuqShLfGP4Pjlh7haTJlsfP8u6f6iL7czFL6BUfKzEQF9LCWqo
XxB0g7p8hDf9j3WVoHMiSG1OL1Y28O49IqJpVzdJdMTejUlbcQJCA/zYNJyIVcwq
oQECw+HiVAUTS1Sq2zHgT4tWJElGAyjEAFsKOyoDiX1j7l4wTXae5Z6k2JpK2wiO
clJ9SbaSDj/AwBhmfey/HayQ+RLdxamfsTdeJJJYY8bMOCRCnsSJuk0RsMPT2usI
WqqQ7ch1qf5PwVWaWfJdF3WwwXlLuVbiscjNl46g9wMn+HnWX9u+s4k9PmF2yNqw
iqNTOL+fGcmT/zlre7onKYrPX/UMBY7nA2Miy+EW04aVFrNz+bmAcb7/9I2qNA7w
g4ZUNn1PZNpyBgPG43/7gxBB76EmhzQprumnvbMSud0ZYg7afbmXj+Rqya0miGCO
nLe9q4j6hyLnshhhB4VSzx6oBYfqcSlPt4+o+v8FXNbMYaM4UKY2HZ4U1y94dHtc
G3SYfjo3NGgGA/ZcB09ztGg0govzKIYUCTnuLfe7GjfkjyAo87hcUK3f4DKLmbnT
2ChGncFXkMCeT9UtUDbRzyfebGuaopT7LHAj1uEn7PvQyY9UnBaKBi9IGUuFNwuS
yRKCObibWaj1k38o/irRe/Tv7sfSqNSU0PiXBvVk3mUOrBOz65jayShnGQz7qJV0
9EHNJGaD0xZPRHL/mbExUZyPLSpHfAWvsgaaX90bYVpS++KCRmqdzRuid/VoB8+i
O1LTkRaFISoQP0/qweSczacWEwvvgoFATs27YZQI+SRAh4jMgBdTjK8BKWQfN5LC
ERsA5fARfBqH7BQGronnC6dXiA2yUw/gKORiB08DodxaPMrLSeb2CfN7xyRghwHe
ObYs1gk8R6i0ANYiLrcZHjuTcfZIUhWi7QMOTfcYtP6Qa3w5LXitzvXHh99AZbzU
CHt0cI8O3ERxqcJO7Xk0Vqi72DKrzQE50eCbtyQwLu7Le90cPB2767k6NN07lwas
GTSd7KQaovBOJ4ZSyIWch6Bmh6Bz0Yc6gZk668WL/qTNeUzRcO7Pa6vmBsdmf8ca
oDEUQ5xKVK3dunRVcEeKC4D1iqmp8Mq4z9pt86n3iWMaNvg07PBXUUgjwiwvBP+I
wPX0VHtP4Szy1g2PNA9AhHi/TazcJHVtmxVvqXC9tSFKM4GIzfWmi87kQDDixCKG
/yLLKHR9S3UTPBQOg55aeP8ec7ToE7Det6VgwyrAipSMxKcq/VnHpj1TEWfVBDyc
U8wAu9RaNQDRyuM3cGLbReZCCmNezpIcHRxHPhI+vveflgx1vwv0/opNupZrEIkj
R8CNrJ5qomcKw7z4yit2LBmipz+R/bHnxNQVD7vnZk0PmRv93REdqHQF/xp01F6g
/PMtP/E5qFLa9dCtKlMGwJ4talDaG/jXleeRqUr96lYtzWAfeWpZVuiNE6ALEWBG
D1OofTwwrJ3N1w7GE1ubjRCsqxLAFPN00iZXTaHq/n627709jiLtEZ6kIXfrau6x
13hEYlKdwZ6FtYz+Dymfs49mpYlUdshblSQyWvbOWKECLzAU4PWjhJ1RaL2Jkw06
tVLNIlftkCfLxScTsIApBwkq9nTR9ZUWpquE+GXJIB9WPkQYWwu6p/duTCNRYsXk
cjQ9+JrSyRz3S0qWfeUywBz8DKSlAE9EQJTLKA88925bwcIpqOInoMqISy7Ahf0Z
0JhuzaOigaZwG/KRgxJUPSYmg36BlUON+qucZBDip1qhZDFZMdTkuwduGT7kIJ5z
pI1z3Fka3Uf5sQio4fkJiw67Ew7UptDBowS4F5Qr7M93S5RqQbSwfYExmWEF/OmE
XuU0iOjNYZKWZfGUbUgjCRXxARwpNkJCVXiH7R/FqhA7U+5vgazW4vA7K7Ru3Bnz
RQh0gHNAA3PD07Qzh/iwViKH/tOTBYNy4is7lsotbt587MHaQx9h2PK+AVc+JLvl
Y4vto2iLgfiLWZrrDZ1s9x/1fzd8aAEX3AAz8HywhEAvl8xTyEP5Twk3lV2DrwEI
fZN5CXe07rQgmfCObW5U2yLq2MOIv8TyfOiAHORA13madgzyfQG17bpDeIeUcD2c
kWhy2xe6oYd+PnxwlcUo1JCkeVPWkQFtzoCJfkpu9OIusvTDGS9KquMZ62VL0tir
Xos7aHGGa/BUJJ6oD27W9uFBq4ySxP/YiDtBpkCMFwJumDtzxjwXZ9VNjpHsKjc9
1oPkJEj7aWL/jWpRPM8+oNl++eQXi0df1TD14l7wxOco/rjMcw6XOW2UDihxPKFJ
3jmaEFgBcvDPhLacuMLPXy1ceNqWWLfQfLOWLPvqb8dGaOCn7RXdsyfTLrvjjVyg
pztWV+0cfPVzAk3mLArK1S07OnmSD5M4m4ZE04/ecZsR1aYsT+pYnEkYhBKyZiEf
G4FEf4RRtc4vu5dTYlxzCS+8AD6qvOTXZftXtvC1H+WwtWm4HDyfdmyVZM4/r3JY
Hkq0hfW+RRQzwiTyg02lYrq2pZ0lfRO9H1e1LyX5WXFmKAAE7+TAv37UAyxEGVrI
HkkmkjBn6a34p+KWAWVEBV16DoPvQxVEtsIfVWn+4jN0t2XQu6vS7whMQDHvM5oR
KlwDug+FYq+S1fgd22fe6mBlhDTrR8bj2fS9B/87xheWLF/BulhT5iqJSufbq2G/
i+MMM2TOUZOgDCkBTXkyyXODPD8FMcGDvdmP9sn/JTMw60U1gt8u7wYyHHs7XmYO
TfOL222t7pyOd8Ggng5SodMiZSTnwZyUDgIFSc6QCVwev/eX8/PNMyf+O2V0EfGr
mOTijQOjnZjSrAy3kgKu72yYCCpcVPQIuozJenfRm8S0XxZUhiKzKzizYg2Hx70I
RwNl16YWSotqsw265ObtokG4CH27WsXRMwqJyXNwhdPQmzCq/0ITEo2dbqFmd5W7
5wkFQRjeW6PESYd6HXwTDSDZfpi/2rgK1FUAWz8a5S8N4Bt9/sg87iELr5HiBVl7
NuaLW9fhSSuU8FTXWdxpaJluy3QPtk0MW8dGrlJgBQ5KmVgc6VYU0ZRzXkNkx0rb
R5z0uj/XBdE7eOwq1mT1jlB5Mgba4IYd7PRSJUZeoOGZNml2Z0NYQssT8BU5D+Dg
CwVhKf5bU9LuAQuZeUNbhbt4HlMbYUzMUYvsIDV4VFJ+R4pdMaXddDC0tG9T04Yj
/3RLh6UYMfn9tLdKm752fpWILvoGhsiR1AL00qou6LejddAKS+bmnCoQm3JQ/RV5
ggOeLj1922kaYymvDip72xUtCAlT774ONDZmS+viJIjAx0iqTRtHhAGzhc74xwkU
bPk2Mybabn7GDeXHW4FpL2M/DAxlJtnq9Jq0Sb/VqIALPF3psT2CSuh6U2iQmw/0
w5pwxUyJsA/UwfO4HazqG0T3WmtnCh/+RcRKZOWSyZLmRDBk9/off670kIBlXz0Q
eIpH2F8mCKIkfhcX4rc7lFTJBRbgzdiBlzt5McjG7sY5HoVjqhUGZM4+tIw+dRHs
XsMDdaowuHjJZ3C0BI9IPB8o7HzXbFm1SVkaUkKGAYJfbLbQ0wJEddp1Zb5cp4VO
biRb1aPGXd6VlwBg3PG6hMA+sCjLHCkbiElPB7we9TBjDVprSe65FMbdoMl6a3dC
eCYPgxYTajKVGaLj7+HJundZunG7O+AnpO8BFFqzw/9t9IjvYacCMhRTJlU5rGWY
DbpWZFMCWkBS+emPiCr0Oz8JmJs1fmNYn8Vc1/+0iXcyg2S7KP5/R8Nx88Zl0uk4
u/aV07FV6TrqZlVTJxq20qkqvjNioXa/U4b8ximEL07YaYKoVc0vcNdT4nnyEXXq
L886q9C0Pk/oeHRYtfwIkjKIakXLUPManKRyh5rjeXY7CbkRqLTUH+TPkZZk7bfm
EvN//resH/LNXsrvNlFlkS5T3Otw4QP74BjVT3Wxd52pqBQDcdmOqqGlTEL6F95V
J5KhB2M9nTwD7QH5p4qc/imk/GdxHTas1BK+zol18jZxSUy/coUpMYknt5WrDXFp
RUd6c03F2rHrJXHEiIg/02WdzWrcS5yj0bxXDeaZphilx00bO3oSzggCN87zRfNb
6411P+LDeAnRijg7poPEGviLTilCeydltZb96/m2k2TVpbmIgfpHTjZaSfkzQ1ck
cFxm40GO5S05veJgL9Go7InHLrDAFdDBWKZXAwX+muzDnCd/HztXurNTt4P4qlnz
qW2N7M3P1A7g8wEMT9uNjCPVFjq3I0nT3843IYO6I5x3JowyvxmsgNnlan+SOy8+
I8PuQgFTMf5agIe2KdGneRFrOjBWp5Fkxqqq3NBfB9Z+MKEnM04A2mZ/iRxEBh24
76l+fhaPbusrZY9yczuHxzXVG+fFiTWi1+dcqg/daIgfrZgSvUUt32uhvRrKbB2g
gvy+WxsC8nFNrjgH/zMjI99Pm5rHsratbVE30yiADTP/lG5G+S4TUlPS7RCXiGQ/
HXLXzjRB1oXE8D9s4ChGvgdUTRC1GcV0RA1hc6xJHkF/g3QWy7f6OpuR9oycy4Ju
LFODBwxs2tqVIkfsaPzSAr1pNVvxQlFiar8I9EQ2mfu6j0g9AogFT0O/nHfd/GKg
SOtlZbLUjXvRH6+G7A+bhggLl3tY30vMQi3gPCDf0DB2aYNlES2WnytfROUzdH1b
Fk46YwSM1K4ceWCQalMq2I5yNUxUf4s+HTWzHlnNnAi5cuMlHW+z8be8QENvsax9
zqJsErpkQoeq9/E/5sM/MJGmQYqRd9aphyNJf03+lAoJapcFQ1BTT12L0N6oCUzS
Z+sbS62Rt9Yft25o6Kup/9+HHSkHFNam1VPIEwrwadO2DFFs0nW+kSyNs8vIxuQW
fVy1B/MNoTmZe+Tgip98WfdUAFGPh8fHtjdujx4B5AppCsBE1MO3N4cRbUGvNbI/
qOy1n2KBA0oGyxr1t/p+obOHlaC4WSBSjws+4tYN5tg3/d7RsX02+Vu4wm+r2qDd
JYEbEsfu4XNhP0qjslwch4Sut8vMB9ML2iWLl4yTAQBwwXbAbrindTL3HZ2YqCmS
xGQVBaSLjunoVUNCOFq8huhbAw6yHuxgcvdmsXo19mtVK2n3yRAKRSanrVhCu15M
aQZ53jalg+8ZvoBoqoupoFrRme5yC6eD/WR9kVt/ju9NNTLd/fR9zAQZbmDPZkwB
N0TEe5mZ6Im9t7HCKIYVrUwsvGAnPK8dUH1dzPN+uR+lwdtV9enhaLuoe2CI5/aH
euqaLMXz/CFhBebR4bBg/oXzUCLDGhZ7kER9Rb6KjC2r1ByVOUG5zMca1zbBnB04
RewWvi0gJEWvC2bci+uMUQ285ht5Pqk3fzDYhjAYWDIbsAh97yPqBacNyutrA69w
wGeyeADRaZceoUKnpM6ANQIg+kFuM3034y8HOx3xxuaJUxM1tTOfO/T4Z9AR2GlO
oyJB4WcFFQQZgUwxM4msRebQ8hZr+Ad7/57wV0+yrEGmveCLlhGsxYETPCrkf3tL
i3B/HyeotXNpiRT9k+r2ejgK4UcEppW9CO5HHa/kjFGcdJiceoIz+FsW7oRD0qPp
wwMdU5ECWiAd7FK3/1CVvcrYPY08M2J0Hz6SlbilRy9qcSQUYPEM7tGXg60HQo/Q
dmCMUnr1owEt4AtO0CMQWb1fTqQAD3sVALYm2fbOq2egXXvaf6ZzQzuPiDy+Q/Zv
hmd7eTi5x6OlQbYldMjca7UfYgSEEen17Se8XvbPpSmpoMXTzBnxM6BmAb1z8zph
9209L02/0dl7xcZI4qBe9JZXc4cvJEuU2r/Ia1Syb4wiT5vwGQNLCc5I99gGOJYb
nYscmUWDiRLd7RrquiXm/InyUgCb+IXXMqK0yCJAh8q0VODc9WTLWWNSUQUYd61o
vg1crZiTGSvzaMpDt7C3vguheRNvgewwIT/wi0uXyYjcgmHC8I0ylycfZHdsEveu
b6813Tlw8Wc8xhl+bLNA8H8gbOS1hoh5Yo8tYAprEt6upOtJfEw9wIeee2f8aolr
qbdIPcpVlozT4P2GQLOvaGYIHx9Vhx99oFl/1+ila0vZeLfXrglXaO1Y2qaNFAba
IwHNWYfkSotarZtdV/GHwSPYoTDM1nQ1peqlzZ2jUXyXQeGtDWxk7QnZgD39nhcy
fp1GU0dhhm2SOR4RZ99ktWz+8uloLKQZmsR99RW8TFk1DzXBkGZH+AOkreZrSaGw
DDd3yE9eUixGgwcHq6kfNc9VsQPPZW/+W69PnmWrrwcrk4tZghc0l02Kh1g46NQP
4AMAzXUKtr43/TaZTZG/b5OLPVXRW49G9MKvYqajONJtYQBkR5jfgj9/pXw6SN1H
6Bsg3XX2KMD2YaugEfrc6Fm8Wlb+lzvilbu2ovNwSgseFg/9t1MsR3GGKTwTTHND
RNbobBjeZZLkcs1PbyhdmsmWPK5faJRrWZK669eo7ui0gsi8JeWjNxSQ7rJ+rntt
9Op6pY38YxsJxVHvux+NUMLXxTjfLNFT58l41pI0c58VOWpzaDKpr3sUeSN92qZ2
qlNSFL8BuopntDmfgMO1WyRZiviVOlv/rl7rqDE5Yi1dNe3OThD/UKbE3ZMiWn4k
9CQ4nNolNnkkKmZbh0CIRLyZHh6CM7KCXcXOeIwedckOZkUWQfRZWa6LoNsldDo7
6ve1eD6ALbh3PUyszcI8iaG6tRV+yNokp+elnpy64iIzyLnzh/UoziUK0VzTQuX5
Dx2YzlA3+jTqWklTR+TDgo0OeFxEaPFUN8ieq7VaUpT0p8VRn8uQZ3C1o16xrtGT
rzpy4mbKJOLeOHi6iL7esK063wheQ0fG9Ensovty3HC0cjhbeffvItJz5zpXkqgc
SAW7jts2GUtNwcXaFNj2R0ydPlH9Ku1Wikt2Ctmzn1a+xd1SGEsV6JJGCj1pP3t0
+taMJxNoeaAeB8t04pCXFYoJsb/7aH8cGvqPht08onmVT0D610eIkpu3irXSzxdw
JSb94J5mM8KG4Od0HCMq9rCLTgPH24gvHX4Sy9gG6ViJB1Dd5+TCViT0FzZneZ5c
yXvlQq9CDhn2/2DEYK4+aPJaqapmCmQQrDFC2dm514VdlvAAbi81l/det61zEJ2k
oGkSZkNenS4ol47poqMXUa8SwhSjt5cVLikXcMof7chuj/XGawlpKeCEES1W0ER3
IO7VgPu5IR9jPH0jD/R3rphjjd0Ii0ycSKHe6vIpNE+i3+QnfBFhnxoJMPG/mMaW
u3yZJ8SQPbI1a72jGxodh+l7t1lSQNpFddSk8BSMunWu9r4v4f+OlA0q7EHUN9RC
3kUWR3dzUstRc+39prGFUPXZahcOewytHLRZlAE2+b9uCQS5dPpfl5qneF1AKDw5
Gqb6cVBSDMrjFT58J0DHxwkP0RdV7NAnw1quVsVCkoOqtAF4ebucHXDE9cN2ZPsN
Yacn4TQxVUXL9kpPLcdNm4PRpR7pQJQqpR5FWgrl2+6wTzPE/Mo404jJ7FJKYBny
25da05OT8I7muP2xqoLuZXR44OZtrSHJo3vKtikr0Kn26erNr0EGLaWCKqRiwKeA
12UbFzAJWrfp3bhXrjV5tEs0BZg7xJcthYDuQJglvxv6xZbbm4Fzcb8BiRTRspLT
1RSMJsq9WRALmipL42bE4ATQTkt8JpBGRKDvYmW/7P9IhEEIgOUPECCKV6s+ut8J
SSzfmxYsGEKEAaP5XILmOX6SAfhZ/1djuLZ4S+4Zui0cp0rNANMWpGPXBJUYnKPO
wnO3tNP6ehk+pSXUAtp8MOOTr9KuaSmV0JBk9wxmA56DQxNHrqjoN5MTWXfGsNvj
OolNuQu8HwRM1FFv+DWZE49SsKwbDVj6zLWItXegsSORQlwWXFdy02aV7gDQsLe+
817G6bIqcCf+6sIzlTjpAOOdb9/wtLD2O92BMa1CxlNSo+qN6q4EHvcIm5zg6y0i
TewsiRedJgttYtEcMcxG5nZ7oLgOIZcsu+pzLHnrWFFj5VLoPd9gBlOCTmJAuDT+
dXHDG5sqAoIZ2l6CAJEhcGvfFqrJTSnorhDhGmIRanOYx8KBSwl3dBDp2m9Zyl2v
IhTXhaQO+d62eKQqVhZLi8s+OVFLwhQtvBYfrXG0VRR2fxJQt2675xmV6l4fWcmY
ZQ7J7VdCUuxfwPfcKvQ5MztCgH6EvVsJuNLl0DRNpMFkL313WKI+LYIxxxLq0g2x
9p7eb0IIhyVatc9MAXaQ38YtR5Ns/snE3Q08fD27FSN+h1yjr+RrcP+/zMra7X7w
ZbTZnwZ8S603fyFlEEctxKihFFhyinr+LpYQA+66FK79THn5Ey56NkN6rsWodLkl
0oGufvEOKN0LLtwNOe+YGJt/tU103y+AORARyMwwModAQv+2QyuwyZmcWsVFlDyU
4WXm++y6p3KdYnEtpV9qY5FMEAY6Xtom+RKqx6smxX/EGpwXRqgnRZpLVtnBXvy9
e4WE5igUi4H0T3b6N1IAEThATIWoD1GSMLpD1zksPDtyOkS8veuV2OfOVyyLRqqM
w2U9G+2BYmwUrTjdfkNPWvlIB7QLw26vNvkT4Dj0GInpTAXC8p4pHIURRyYnIUTU
OiZWWcinUKGSImkuVfYMcT6wphhsW9McRimomrOE1xvKkO7G0GO+hMS58fUh3dvo
AfTwx5p7M5IjvafwtYGn8itbOK0yN2SHgGBUhkShHJCvdhrkrngFyywrOIHjCDoA
qGostEcEVtmd2ndhSpJHssbRv+pugsmV+9GppOrhsAfV3VwAyObovJ7W4ayBPWAY
cxGVuFhDWgDp01DrDy/1f9Y7CO/gHg65/1b2YemESwK7fZyyD4BjtyGlAkQAaDWg
dfzos6ebPr1gvT0RTb49cjZDEeINQAdw18BWExC/WQTBfzCl4VzYUsGcOAsKsmtL
SYZsY2mJMq9OaEKXJXDxhV4wVnO/sKf/Y/yXV1HxHTFdFmjH0LurcDmQhlpfMilE
6PVEwM5Mdyy63BI1LOApgPStUxeR2wz94UUoasG5xI4/I+3qiwuo97dMPqV33aGW
jpuPy0GVA6nXG3qCMlgahqwo53fgAqcXIGkwGXSrUDLetPRgCX95dlxPURA4It9X
jHffszPi0l1K0uIcoHh8kxLzwuyFuYvpxW7mubJ3UZCl2nDdqjIwBcL404u/aw83
IkWD6e9OfjzVv+GuTqaWP+W42NzG5qQaAR/KxD7IailrOjewCkFsQBJfePLny5SX
GhRwIAa70BobbwByL/PyPCEBVY3fCdEoNSrlhaXwGmMexbD0NC6BtX2WtaOzFlnM
GAOtEaAhB8g51CFlUrn0li2Oama881Bg3HreZV2+2jCXOgK3LRJgxxpKCxvRSP3I
T+YN7GR7BKvvO8CTl4chBmb1fYskp673o0LLdBJDzOrV5jVZ8rS3MfNfrv4fnc2o
RuXPE6egDEVCpCZtT3mKjNgUe8a7ydOZK2khicSTTomoHIFn1wIQjy5jPaLTLgmu
GenRbrXX/M/AVdEvPdEk6BwAAK2vE8YSMyizWUbfnJXiGjfrUgdzeoGnNjSbcnU1
jD29mZjaXVP5QhhpNQCCMuKlpHsdTu9JcISyC0H3aYy14kNtnNf9LxKbTg4bTw+8
zOWpeEKQJzomUfoPcIgnaXG8+/7WmZ734OoslDjGO7Yr7HNZS+aFWJkV3UjDDcaU
i8uOrdg5BP/IImZc46zG5xfiiAzsnIYJdvGoP0P8C4cuTyzltCFQB2kM/euQagM9
UH5d9KXJS5rOnTjysZoT7TdVuAKPtFyyNFj+6rDLWGqn1Csla1hfqRJzAiTdUVlI
zrg2P5wqddxBV3W0XteeaLV2Cc5uWbCya7rVV4FCmUXt7cDv4VKcd6DzHKJwjI+G
1jdIcRsbQ1cD9PDE5V7rWh2gEEf0wePFUfdIqcCSHPKAFR6AZ5fEs+QhQdE/N8Dj
dswTmSraiUVDP3bJSNaDf6/m3w6bBRxN//CE+REeZziPQGi/DPi/Z23zm1DC/f9t
u0bLsDgn+b3wpnbHzdQQCNlf3uPwCGfYgzbm3K9Af3vKfmj4Hu+EkNLQJZICGM1d
8BOHHREjr5yTiagyDjDWyw/vRbRj/UcSwj6v0WtqNyt6LxxcZ7zx1rlIy5OJ/Oed
IMvHEaG0A24p/9JyKjV+p7v1E9CzHu3ajxsiiwPlOgkJ1A2uEBZGlW0RxG9Hkp8S
4Ra4DCH582mLwNMhfdhXDpxh6MVq907ANBgMjK6Lo+mzfMf9ZYB6WslvLiUNl9qr
mIDlutDfiFYWA1OWs26mxLTJajUUwkyznjXKy4/kdizh6eq0BjndDK1aUxtLg4vb
t1Ji9USdGgqonJqr4fZuo3HPT0HLo9GYmpWxkkIyDTSp+KKQaYyiwYyEiBbuLbb0
Pp6FqN7+JnJATBS55covAIZV8LA6+Zm4oW7svyDKlScn3HH8yhWTFM5bFLRfM9Ul
wzUh6OEd9nYkE+ZzyfHno+j9XKGYSHFVqr9Vl/Kz2bBUMrVxTkqZ0+TyjIrYtD/M
O3R0gMS2qQug53ZNJw3DJRxxh/GirbkQS86c3tgmO5HON2nQSX7M+TnCOjEpVkLb
Jj/TbhyMknMb6xr1gAzwYB5+TaSaG7bLRxidhKWUOb7jikPScI/gPnxJfEqKo4UQ
i6OeaB9EZepwQmdS5rMf+9ZP+FexaLs8cqfn5Gd57lwUJCxo+IE0ucZpo5Mm1wim
ZhORgMd3CaWo8LuoMMdet1bvoM5LrdPEQjWbOr+FTxFa04mLbj2yH1cdFYAw7ki9
CUnagg1qSyOqCJPDJKqTFE49clndB2Wl52L8xJAcAdCH77m159KevBULs/fOxvlL
yu9JKUGN7XwnFCou404yBxtj9Db2UMubqJx5AjyQC3qAkKSXAMmsD1mHlXIM64+m
KwEwIsgKu2MU8wI3S/bX0g06iK3GDeE2c9fx707/ztzQ327dce6i49zV8BHRba9/
dZNMRgXWgAud4RgiqCgaaHjbgWaqpoYUuQo6+8xCKtNUbIlUFvmRWEhddwKCZLRK
Yjsswv0xAKvlDKie2JXOwJdFtdathIkIJHo4tEWmsOrHgDTwXWmSvXPBmt3+m/zw
GdhOZl9LzjWvJNpHcnuJJoaMNRaPD4ox8FrbOJ2uRSNrIQltV3oNBWPqdWVQFe6E
iQdzyPHdNNwvnFUG55eocvFf+StGSHIw/c5TkOxNopFEbOmZZifXttU7/DL3JTq/
2CyNakUr4hXzcff7u6yA3d5GqrDbLxzjhdmEZY1+M958dyXE5wEw9KzzqrFT+RvX
/Ml/N8cB4bzX84r+R/X8GnCasoWnirHtQgKU6+G6KLaiGBgMudY+wCy3zow4uj9C
ZfRLmtRQzJRIyUqrwAgWuEQIw7pKHCCWPgOsnX2ghWjFGfEE9zJ7ToSR+wnywM6c
CTTd4O1fFLBsgSMD2YbW8124vEw5vtwrtAKRz3Nr2Kf7J5jFIzqK5ni1JnOjsZOx
qTrR8Okta4W1ZEu9PWTTwP3/9/w5dElKqMgcuCzItnKW1Ig6D1qCn6E+8HwQxTNz
PixGSywd8eB5E3Z+MrDuXmfSpQQCAUzIINWqtSWUo8CCUAJKPPFQlfw1CwZm+wvy
WUxIVq27AJoCdyv3Tk8gIX0mYwpK3F90T1fun4dxDNA22dgBzqLpJqYrOAiS20+C
YBBFTqzDCI5ugT7coPnWD6VZ3r+p944utaaizei0s0Exk723UxmodUzqrPyfdUfI
DIveu2mzNNtsjZ7ICmdiYRB5qBZuBypJRa46c/eUgL/rhzXB0pI9vRK3AawpOdgO
kEUIeOExHDuCNjzGRMikQV3E6iPBVQeGjhOMVxFK90Xxy9L9gVR4lsw4VP44wdxe
k0+QYYly1B5jsvchIx0WCr9QDQUvSEmht5pVrN1Eq9iKlugleEWN9JTEgIC/zsC7
Ub55IVG3Dv2/09t83JnAdteIzRmj1u6pCqrZEn0FK+CuaxQvoRtWSu96LMAO41D+
JY9SjfGw+RAlSNNsiwuU5Yn3tKOqCajPPiLGQm3gqKeARlNoaLzGEYcx6NMTRTFX
LKT5ScGfFA3iSnJ3Y+V1G6kpPWKfAS7Ceu5V9hipZxFqzi75wnzkOqQL7jc3PVeP
UqIGux/hnzrnXEGquOVwMFxKdBgV9+38l1Ns5Ppiu4wp4lzHqJegk0lPtn8TGpTz
3QyoHybP6BJ9cZ6kM8x7NUF8ItyJ6eqVkvW9MTqPKR3ijLYdLbpNvjXvaM73yOE8
Y7g0AF9QW/wCzXeMbS97jhSRw7FkUqdjitICe9Z1c531cPBuxAkrcYNwKW/Sxq+y
EDVyYpPzQ3JD/GlRr5OqrAzpoV/4Rkl0LCFNFd1q1uliuUHe86GA5zh+nwEKH1IJ
I1OEFPVwj40lMUmnAyiODuxITYCvmjgg0/4Xmcx0NbqESN5KeY5lkRdFKo8q265J
rYggNIawlzMi/L9hf65Bfm5H9wjYMar/FZ4Yd/nMtrD3xEUiJmITwKW7jwv8k9dS
6XFJKp+oIgbuNndvMZpuZ48HBN70DOn9l14TSIKiq0rfdp7Sn0UB2qQs/73YPSr4
Vb9avwlH0a3knbd/quyzWCTjWUMm/fVvC27nZplkLpq3lMIAXuRqx4aDF2lJRU2p
yyiwHQRjrkgyggR8lZ4Ium7Ko+A2dyL5GHDUaL1iYuSNp0iNPcGqmlNOv8zCIGww
8bWIEJyj/qQyMsyQwT1oYFc7cUPP3hghzAUP3NHB9X2sMutjnSly3MBBEmLB+J/u
e/5K1wgqUX7oea/7SJfDBPacYv6+qj2OAbaKYxYgACO/Na5Obvo5Q82+EBPMsDAq
wUWyX7mkamfPkezwOPuuQWJjgP7VYbGGQy2yunM3Q6p5KcYSRJhxK2Dxrins7sYB
ulycgUN9LUszBUPL8yAXUnskuR8hC9khsY6gZhK3SnEi1zD9S/vOKCIA4RVbmh0U
+ib9kST+aVc5pGtLo59gaS10MpuG2n944uK5To4KBCQdTtsw/1vse+ie5UdLCiNd
L693GYLnhFhWd+p2JhlMT+KdYnGHHRyVJcGa3UgCD9Y0UcAgY68I/XBHSqR8oe5S
nUrO5edgHmiPzwQcg616lLmJw4etig+e+oBNYN33h3J7PGCDqAUZ3A8PQmqE1cxx
c8WUTP+S7xaUnuK5aTw0mF+TuVwzoaAYlIQOKtVMWlG/fnXhsyAiDyAsC5O81Fyx
M3ywP+DM57tDGQtjs6MxTmPozJMJhFhjzOHmE5T090+QtEsYJ+aJnXcuU8gGQqzA
H+gFk43JUuSV5AYLWsBKquRYiBdMHA1NDtmrruoitoESdKFmvOB2iPeOfn5Yrwtd
yD65sedwLl2NEfF2iz2aa9IHXIJ9Dlad4RhQpyS53XCJEQDVF4sWHcu1A2pWR4nx
ftPjl5DdsGWSkbiN90WgCaNBb0Wpn8yFhca/L7SLs1Ugt69odjLT/Xgg/icW8kqE
QUHF57FrgvIw3AiDPsAlOUd3c8ZnfoKGRmCB+peVcqwvltlWO5ap1mzB+AAjPstC
mKS2ae5S4NyoFyeIC27UsBr/B/9k7xd0lMJp4mv2dypBEmMWf+Yyn9ML/iFtQjlu
9bXuEVm+HpkWen8cOlprg3RXial/skJoD9GD8hDc66T4ruVzjBKP/EeIPKXzdSto
0Hf/GbsnJV+2ARf658sXBDv8+D93C94EpWCRdQ9br3150O74pdYnlvXtjle3LHYa
aspEyjlTOFqmg4DEz0Yev4bO0HCBtKKoVLGklzoGbcZggjaFH4iOr9Dn1C369Gqm
JRj697b3/TjcngMHJ5DZL7ASnSL+64KFGQvQOhQU8URFT8DP9cJxRB2zjhwUkQCS
y2+nVPN34P3oc4AFn4nR0GSKwZd9AocCLUaujZ/nQqir4kgmG6353LeDe0kkhGkP
WwiCXSepSPn7xL83cEvzf6JY3QY+E16jqGl1fOjFksI2Uwo/5qB54n4PE6bYQXQ8
PTpODMJv+59DaChr9yJMe6jzawlqJDoszq1HST7t3fxzwzGNZMVDjbYjdP9Y98GL
5U22fpHDYrAth509Oooe/dhdYQM2sUphmhgkHst72hGntwJuPYqELXErzX32xZeI
n0EBf638S64aqLpH+/Al1iCoTSZSCNeEvtKi8uVnll4OoMR0kp8DAysefePp3KVy
4k2GlyRPtYK3UaW/huAjmaOsdE9F9T/cKjSrk9EguEuSGK/o8XpkmwuQLLe/Jruf
eZBIhDSLpJTfwWh5oajwadkL8XkeUDVi7QOIqIA3beCQYKt1BpL/bsF+nRO7Xt8Z
G5vGik3wZvL0ayAeu+iRM17++GDqvIh1i0wtIWKWvwqvZEyaFjAEVjzzK7hAnQov
ua5wktp4GEeLt6vcKWqj5QCQAZ80omtkUaKhJbKQeO41jvrMy04zKSgeIPOj46f6
OwemK5BlBGaFvoq199NbfAm/coa3wT0iKZQIPWUA4Gru+ZWdmjI16RMgQa9LKSfb
AtqbgGkKiUWi/csuiV1ZhKW5EstU015Dfzls9hqKRtZmCN+fWaiIHTB7GFlxeOUJ
oox2nnT21omk3e+a4XPupZkhExXKnssab1S15UuHEbYU6wom0r8ojvKYSuBuNQhh
wf2yzQZ+KWxey7/ZYq8x6K05oKs0EoxWfik1CEQqFGxGKhyOuZe1TMows9pms7+O
sTzrzZwVJTn5Cbn+AnXTScVNRu/y8Crfcgb0RPAb8lOg9xOdbbIkV2ARMjJBKEBa
mP6DgOVfKfCAOtnPzcbyz+ldZxg7tlezrXVwkjipjDSwqq8Oq4oDId8A1JIg33wi
/jHOvi3oXndd5WmMxGc+VPkAT9xChNMvB9qK/+EivGzBCoJSTlTUVlP1ui1yV+nH
pJPqiD2iOPEj/mgKYavI21qLj1/ErA+C+q4S3c83GjM9l8OELPObPPuPpUlmnjgk
9fFbB5r0Cjsr33xrLRE/elUS4X2h2O79Om1ac2BIS4rFn2FtJw+i9v/4IoMiVqWe
Ff30p7354tpHAuYuKPGEEd2nIQnGkCQ9gGVg4RC553FcMeVE9Iv4b0vxbaO2WQ8u
pFT+mb5jnH9LeeldK9Jv5ZHmGtGtDxzCi24Sz8obJzhqjzOX+YumqSQwtqNxCEWo
u7qo/oVoFvwxHxNy/8CZFSpL3a9t/ik6bTe4+x8FJET9ctxp9RwPz0EP2NuuzYTq
xAtmPydD8l1ibvhwVtuYAHvbParTDR6SokYhva+MbnEvtcm7YXrEm/Wup3atwpbv
FgTXGJk8GxU88C53XjeNY0pkKsuiLHszemnDjFkdV6kyzQHMSuVhFsVVcMKA4QEX
+KXmmvWqNveGCmzWYcxNKX47tkfFb6LIJJ0mIXw5Qvnn02r604nmXL/wVep3Qqdb
NOtXVq7S1f3hRRrxYxaUPu9cJLpWBgNY+SEoruxYtXqJf8mpSNh7MG/uZaj2Ahfy
b2C2hKfbBBNP+7aGkTXTJF5b5j9zCqWUHR2QorS3GQ7gZ2uKe646ZIIxe71XhSQi
yZ6jRWKEXfSH8SpocuSMvX15oKNLut7vv6uauEbTYeh1+UUWsSPssq0bB9rFJUFX
IyTdvgr8WMA0WY9GxK7/i9Cs2Tn9k3qAIctSxuSsQ5WA6vhrZcHARdDuDsz5hn7W
BZ/Zjs7kQT/tPr2alCObu8U8vp6zzWr7JHwamRXYXB6pkiT2K90S6kD3bsP7KFdy
jQZHhw3accJh9rITqPzdG2+aC6rhhVXXqqAw0Otd/QBcrF39L4tTOg/YN1RXg1YU
z9GsxQ30C7BQ4ZlWiUUH3/IbG35LaJ5/1wtE8L1VWDur3VC8j9bC+bGygQV3sN6S
c30ZESwn2w0bliHXjzfR1ctcgiWGY4yEMNfQLvS/3FahP00GrjB8uyRr27TL/z7m
lNo2260lfDLw4pjECELz3YLcrmDxXThNQIV1bv8vLapU488zH0AMfaQ7y4RRnhSv
b1r9G8AzkQK5wmKOz3ErrKDRNuDRI2GLr7VyqxjOs8V+eS1LigQW4nFITy1n414K
MnSKSa2LhP9Yhjjk4N4EYoORCAFRrs692bGzqdD5vTY1Ulh/+ASiAm5wSNG6T2Tu
yezJM97UmxSYK2BXxhiBReIDfQiWiWDMjm7GxPdaryisTrzo4lmQXsqos4VCMnFm
tq6GwA7hcdLBvCA+Rmh6uFP+ILPJV/Q9PEfKabWWp0GtuprHJYwoGgTdvWqcKdzH
W8LbKp2evYUfGE79WENSb566a4oWNxJzkVwfXyGD4oSuKsExULclTHsYIq/NoL61
8qjAEQpmcWdUnJ0KnS8/DS+1kqek0I3EcamTF1ith0p0gcQDQZZ16Xq626dbhcZh
A14uz2CJHRTHyOb0j/1dW9gkz0HqorW1GspbKlUE03I1XteXnQ6x+eXm9uHvilBl
6Zhjnotlqru4WjjSN/7eplxdJNMUnn5aqrTaUiNhZkgWOBaUX4UaQMRHIuyqKxPF
Uk/B0IgXO/UN0slqJcck9QXywub++H6LBPrYvzK7B3WxaJL8N/T3pgLnbnJmVS5m
VVb45n7HXLKTzg8VjaR04NMehc3uo2psda28KgaaOhWWnHo6slV2EuVA5WEfRY0z
S0kRIh3glUUsOmjvXNj4GVHSvT/HHW0LAO9L23RCeFgSzygZl43owrENsS778iIc
SykRUsbbE1rsdQ+idIr90EHfL5FRS24uPYicYT6o7WnoozszCWfpUj4HKVKEPETe
idgJhAzoKJx4xbBWBWMqvZPEcnSCAPO2RKJqkDo2h1yo4cSm5QZzk2rdMYBPtNYC
brTAA3tcPqdQ7uggshcnS4x8GyCDJ5E3ioVWcnlRzgZp8tREPNlcVpGXS4st3Ylf
yj/DEnQ6/WXXt8RDsRMjSamFrSWVIvLTztr6629e2o/M/MOfcEOyxx8VOiledkAt
tcdjPOI2mvAJz8rLkp2TNp9azA1DKMF48l1U+rYlNqeWpVPfTBJySJgTBUN0/fcV
gv4DX1D/95FbaWoPOXs2YzwerPJUirNvlhKMMfMNi68V8dgWS0rNbVA61YZROoms
jbmxB8eq92PDVyVq7sAjo/EociRbPB5zrTOfzKk7v+bgP368L8sSfRkJx6fcJl9m
jikF/RXANe9tVgPG3yOA2xFMYbS3G+qJZoeyY4Bmv3p+eFjS5v2g+9SjzLupLv+k
QbdANInbxTU++eBFXIKj41KUNJYP9Azf74oxTl0m0/nOool56fGR1nh9xIaNQj5d
nP6u1bjUSW736S+sPwDMgtWvcLMxKFeyWY55HWSW9z4WPUQg7XiB7uTPTJPx0SuV
d99Z4E1+i89SllASDv/WZzEwoPIRmJWdTi+mFebac+2w1zqweMk6vliJUChBkgVm
ZAqapi3TnUGa07gb0pJ+vj20jvy0cW0fd13iCCYuO2gCHS/mHlgPNfuQtZ5lVve9
C9vu/B/Y9u8DWXjgHh+uoCmmlB6aZSwkzjfIsQWeTBF+fQ62I23SOQZjD+pLRaXo
poQi0ffRgWKONkEW7GrlnGFW72ypbbnczyfPoz2Mhzkxx+Z0mqQwR75KAfHPyG4v
kzzWRq8ZeGvEkTdLnz5pl6M7QhlsryIoAqG4yAKwqP0vfm6fWycD3To/JwN5KT8G
iFCD6yQdclWbfYnOXIg5DserWGLhwkKT04PFUo2OvGtZoCD2DwY0SvjR3h0lkBLw
zbeRnWeRcJbOMi8gthNPQjjfPSvog3QB4r2Hq+XAcP9faLr37meRqRvMD3oaYsCy
14KYuDMRUFW2xARSrWkSHGFqcsFaGCnwga1N97fCla+xS87iYvH56FgkD3C8dZ3C
WgEoWituqnd8RHtePnDLQh8xyKAicyqUO9XPf/cnnz5q4q/3FPClLuaBpZmgoOWi
4mc4Y/nWyE6OelSaEFiw3LiMC+94l5N0lT6jWEx4HQ1Snz8pvg9k8E3WvdrMe3nl
jobCswOOn4CTMWa5ULwUDYrMkjUCgUsiBsvXVeVCZFOUclYP3lTwUh9/N8l7BnjT
xsGkTJOgRCd0M5PWIoynd7axT3zpBpHhKNgLiEOnjxq+g1dzUyf9fSTQ5oOdQAJY
iecVmrjQTTiQrcVQCojFTFRmnic5bgOF0VY4UohsuBIS7F2VVoXJY/mgmBgsLGzB
Sq8c3/cgodu+6fExzN3r1YJbPMxQIpnASeRJzgQdoOSN46Nprxb7Po7C4C3M3Gsh
kRi2722c/USe/F1TpWOh86xZlKHs1gbGwyLRIbPSLlebzG2LgmBaA+3Fin95Zy9p
j+jaVj9H0CkFCGJy5DoMId8uiNNdbCz5PMTQl2X+4yjS+ptcGvJx95tCLQtNlRK+
A32KiMShK59WtISWefaP7PwzD3sJjHs57LuH6i25lRmWUC2e766uoMh4/KqdCCyN
Z6f0brgO58M642e2Qc8Ha7VTxba25NYprflpdtMb8FLfOpxVFg/7znd/bWJ9D4NK
Pt8PTBtn5cqFjf3rS4nQ37gzyPbVGQ9q9tZKbROapLKx2aEmbsgNY5/WQ8TfLJBX
mkqzBc0niKXoYLKR/jDT20vy1CFhHEY5qRfr15UuE9HAGBge8dw+Xlvh1j9V6tLY
gRFp9vlphT4W/YBkqEbrLPBLymE7Ov1fuCIfFAzU21RogIugKgvOXaAn0sN9umWw
il0FYqx1QcLwLuzsUKhY1EowypPhJedgMlGdJaLaPI4tbYT6UX4UI0Yi9G2MQZ1h
Zx4nRgKV2wEdeLCFZdSNIIMQEHCxti2FsTpmCwABvQ2I70RkUrb34kQ/uKmAuVnp
ipHVvKa4d7W+iSc2G1YvXr/v1xeeOl6KP/Ej5qRYeqobzAISafUywqmcVGvwraqL
E1UqeItAHwH3cwr9zFHzfJ4gk07XVdN40fK4dPIGMlWrO0rZTS30xP40rkcdUAZv
5lXdAnrEMyIJY4LHtkxEGDiYLDta1cqQhE9NOXfK09vGcgqDKH+tKJI3mWFC2Eb+
IxDQ/z9icbRla1g0E+YmBJFSjAWR2e6BeiTRKLo8rUsB+90WTHHt/SS5E7rqtq22
Tr5dcdQ4S2AIsrsPCOUiWabCTW6HIpuKLK2Zge8cOa3FK8+oKzMtQTOVjF0En1RC
OPk7sPDCQoDzCpXnRMrB0I75X+lTfCCqXIZ0lkKqJnIvwn+08Hm4BdKuB81j59HG
RDI4B+WLNjNvEAImgVBdOBZ8z2z72T3rfjGX6bw6mks8xJBc3MNPiR8a/WjIRHC0
CYbVoeNqdPtwO+6Yu1IRdY4JLrKn79mSeibUe5R884bH9OsFhwcwQlC/j8THKQO/
julMsO3pQ3aqtmJDaUE4sgIE/EII/IkqLRF/zYmr+uZLr1gsv5Hwix9v/ueaeCn6
ICZqEHuhQ8NbNTLjsbTbdSZendSBFYSl1Q/dzrSviRSvoWsRaqnLZkEXQGs2mXWb
SR4rVpzfU7v15c/XvCkhSODKYluvBvWOhaeheZxfwkmC3jssyHjQdYuy2Qk0d0be
qAPadwYCd6ClepTK2VKiGbE3GMgVQdK5Q0RRw/hqlsWDzb8TyAp6bKktItFd1f0F
/sfK5V1dUdMU/OgFqpApxPOFoajFOSFHQlls07ad471fYEptEH/yV/8lHxrzfcJ0
BYqSeVglh3Ho7wPgQk+E2n/9fyObK4Dn8mb1dXFWTRs7eHY4Y8IHeyKDFjzv+DwN
IsSyPUfVd4vN4uAP1SAR37Rw3E4myaOkhgzqJNUUTt0bNsd4UE+wN6mbf3xvagiq
JvI/KBuLpksvShlBNseAjJSPJtTzF0nKfVREeY+phhMdW7mRIdllTORkLivsyxTd
u73GiIeUwCI0bMvYogpY7j2ep+0ZiWAL12du/jcJM3tVhKxUHD7ieGQGJPdZVvXb
jQmGGwT322xVyUA48KTu3Ds28+uOdcV64qDhHiULnakWyqf1Q8KmWSW8Lu4r+ZXn
k3N2FMGnik0A2nwpaaQho9Qz7FxKKkHmohKcbuSH8j76428nf1C32E3S4HW9Tlg8
LQAJ0cr5olpwmNMifzz633GBslGNLveIm5231krlA+SZ+wI8G2uCeyAKQiHC/99f
PbB0BXoiyiRTPWlSrJ0+aPvf7JtlbaKnzd3n7lUYliFvYK6YBxuAl8j5wo1beOzu
anCyFyMZqagA6XibbgxHJf96/WYBhOADZuAwqAeQuaoWGe6trmcG6QdbUiiGxedC
I8ARw+VCMXnpDV50NmEaBdtcdLSiUcCe+c/mtMNzgsoQgF6UVfU/pbj4CoS7Hb0f
MAhcvXI7d1prjjhp7qAkSccNC4JaD9JTX0cMcYcz7gVuj1WOMsnIOO4CeGSvAzg/
8PUWNFpGWyfMm3MrUxGbbmEMVigN9fStL6F4ERPd5s7quHWUDnHRSBGZ3ojeG0g/
n3n0I3TITxHRxFqVl3qxTLvrSoiBl9vTEY65yYR401MdMCZqAPOhrMxYS02sbcmn
QpnHVKHhKhfdz3app8yK4rTmxjVt/kFJU2eyHFyjvzMWu9yeG+DWRzcmpE/U+Jiu
+Ve/qol4Dj2mZm2TBg3KBKNW0oLsZGt1pZ8rve/zT2vLaOI6vD/jpBYTztsmAnHX
udiszEIK5VPSWA9vtEoiEgaDAlJONcpcpIUAhcMquFLFZybtC5sexUF1mYT9FYdp
5PkBPDBj0aA3UF7U+KjNRfaZw6kA6ECpO+4GbsOvRdVUIATu6SunAvPI2OdOtKWg
Md0fMGGdae8w8hCWRJkq15G4RTlclmcmwPWl9JXUR4GWH1Zj9gQ0MQDazbl8tp8M
yvVg0Z0mbOsQA/NBUZMjn9H8JqRAtHixn8Vlfoo1Yuw3FGZ14nCwGiPzCzLg50AY
bBY7rOc15zr/UA7rVGO/QstZSWnpXl073duisx93VG9NK0H3D/xvc5TOlkfhUFdm
oFAZo6fqtABBDVqfYFIteqxsS6jf5pmSJgYFnbHnqJbn10Vhlb1Y0qeH9LNa36h7
Saww9fsg/7HCNNoJ7PUZPlYNueLCKoNcWe6RrUORFMpYoX2mtiYzOHNevEjj+mZA
/5iRuTdjpFJH6t0fpSCkUaoS1H1+BqXnw1rg86dSTTMKEC2Uwy3o3vROQEjOFwsn
Wubek+ggNfu/EQQDthqu6lBEq0oRGnulDvXautttPcCB+FvU9MOZC399Hb7FWxdA
llrjWQcqnWr1omOQ/wWW8IzvWKqCV+ohCDeFAQRd8kDITpJ+RjtJwfzY4KHEC4M+
GWLysh4mwLFyMX4/NVZn4XxtcDf46QrMDDSjDIXVocbbyiRIuKdYUVBs/lbvdoKU
ReX3uIe4JfLyk2Fv838GzvjD05ej3ajkfOkPyyL4G2h+/rEkW2F1HtGoI6bhzg9U
v/QGPYVtBiz1Gn4X0s+jRfjWn0aKIwDJpLO4hhF9CbUe97Y0UBtuMAT8jkWUkMe1
m+mPHvc0xlkrMgvzzb9kw13jJqmFPce3LhC3a5kabl50ep/OE9gi0+D1NeT1fkXZ
yp3Fl+SI3Qfl71vnMq5qIrarCO/zGVpLny31RTNoexhnVtNbqvPEF1k1OPq/kLkk
q1WTi6/hgHD98YVI4y7Eol18n4wTj4+yNx8D+KAh4o8ysak/FXGhkv7f+tqNnwS1
f0A4xN6QXNrWYEYUK3GCrilwSQjjV1ilmd4ED8k8mmfmrlEMlIDzyGq2d8Thar8P
aNJxNPNW6XYz6Lf0cjAwhROQtSVv1BZeZGYPubOQAtc8nkG2iXtQA+FhN37I7O48
+410VRsZf6quT30VsyxjHIoLmSZPpEA+oBwDBEpq9hPTfE9sP6/19+VNI5/j9WgA
qxAmDz14l8BF1gFu4p2pg8GAAtd0xGRUWwTuzGsi6qtrw8D6d0ZVGGd5i7Hqbh/z
MgIgoDjVqTDgp1VT/ZIeIhwvlHXnGrg7jmfshH16KYxC6mBYlnvb+Dhxn04xez5t
4MBkT/JKrof9/AV9j4uoJJn4JcdcIaHZqMJvaklnLWHsTmf4X9ac4oiJzS7O+y/b
wFpdHH70Tcrcty7RDbLBM0B28iz0rbc9mc6EhG335cQPNnLMRYdZlG8dFj2GdoqZ
DJbsHm1J/dBXHOQb7My0ekubfi2iHaUtHUWlOMw7SDtWcDxO/8BlVozPyFMw+ukW
skm9VeDFwdKZ8nSKfTBKEyUNNqYMTQJSS8vIHDgY+NCZ1S+dcAv8rz87jbMtloxR
ZjEzeb1oau3Ofq9zKyhnYl7Y/ncCOtNvq6KcY5FLs5umb2PVwyI1MdSzastqmfJM
5LibM4XPLEu794V7X+xpBT/gP7JXPh+UUpnalNvs7EQarjyqi1UadyXIQ/pdufdO
hYAk2gNLTUOVhHkhChxPyhia1SqOcofc37GZCicr/CK9jNMy0iVBLq589shR8uo5
yFzab4qHWx8g4OOwyOuspDqRQtx7ExiE2l5XL1yhHelNyPQYd9oB2iUK19BYNpHD
+Ytv57JkMjbSyu1cT8OH7PD535VsgIJ4AkK0woW74yTu26KEwFGmlr5fJKF1I6Mm
wjN8t016k3GraV5Dnf4C473z45iDs719BkCTKVey09SDNBSq1cs686MYnOHYTLRK
8gxEyXkK+pF62CnlHK6WstXTtSProDCUxI42gAs13lgKYY9sF5DZh7xMqqGG6uZe
XDcn6qYeGOFgppfSOtqHJJzAAszwpBsUaLYgx6ZNUiN8Q/L0zUVQ52Ptd+4ajDXz
d8IzTpxUA89Y2COrP2TFaY4UwLeeyZ3dyi1R7/b+pKXa3awI7Jr16DqxwlAR6y4T
PCp16moPp01TVnP2ffnBlPWg5A94N9khpzrT9LD/c+IMcBvjPAkjjptqSXcr6Xwr
E8DC2M8SsZILQm1RyeRj3ZXuGN+bLHi0tIYN/S3XxEH2bfmR2KZXdj3Qp2upbYYi
9f3wSXRFDbSgD12/0xEwcsZXSqXIa+ObRzzYO7URczYpqHlMzbnWcrIO4hntGQD2
sp39RenQquJ47ZSxJCanIUx+vV+Ubl7RKCDsF8WlIDAFRlxy2AnYCF5yn6IVaOx4
fCcUpVxgTr++CYa2oyBGhlMD+We6sMSkxUxXXPggN3/hk3U1HFJr3rKf35oU2zn8
2aW8o846RkAx0OeP/zDUYd4EtuisqMmIZqfRinpxZe2p0wbNxb0b/lIlT9IKjsZf
mvSTN0Ws3FPe87AASLlj6SMDv5Bcvn4pJvMS5qcs7BzVG4wLuqGHRFKnosStsusl
CVhh98MIoNmuARoC7WPQHIBZv7rLMAhnZcjj1wsTLuPUVYIPj3WYhqyIeYXDXtDZ
XKoofwMp1fZ32czyeIcdiTuNebmP+6boeDpEZbCYTpG/0ppFzgGqWtov+e+yBjdw
2hhliPazowSuzW/XSHSHxUlwxVpe8/gajkuEv8y5S8iQBbmmIRJLJhv1p1W40Jv5
LakiODgYW6vwKV0hggp6r8g7Pj9/VouWiUwYqX5DMfQlzGiw5ZP5Si/rkrN5/1h+
g33whcA87ubHPrJ3Bf+gjd2AwPZabWKbEX1Zn13ONp2HH8eFwwUbHbpC/FmzrE1+
fjh3aHmgzrSPKLl92+CnnyGmYObHDJZN4AbNk+ruM0+BFTIRuea0xSizBl8zVdhj
FgIYsq+eTVjDYejMhQIdUhkOYjDp513f8Mo5MttauQUCBlTRskLAdRGjrZD3ZTHv
hjxhsXDAcfzREKZA9vcVYtcSU0CQr2P4vM82Rw1UBrEDcnrlf5rqjyP5azf5LU4v
aRySxn16KjvHpv6GtzTemKmswUnMSscNr3cceBOtqDrWwAyNOxHJUzBaZWE/Qleu
Ed9US53RBwHIH5vRy9a1e441dvZCWapVCqxEdbE9hj5PWT/ASawkYRL4HwpAgAQt
WTeTYnNNA1aRbnVEzrwz7px6016viOULnzqe8iB8988AApZS+hYNaltqTWzdlN3w
9RKrnRAmxlysdpcLHU7CjyKeUiTuobfUF8aoA5ElNnFdKuLJPfLd0fAEAP4Xo75K
fvsZrAc5v/RAhyeW639CX5MoJCPIpSH+aP+1FdXLKiS/d81Xq5AYcNJckqjC6Pr5
8YtAmOPSYGZxbGWiVYzu2tNp0SHZ8eDMmvfQOtl0y7EUmOG8+Vq46Q6PBBz7bKl0
i3P8ZTu+zfl7Ce7i3e+UMHlwLutPvC/2ggonNNL0Rrp06aHLGVn2nIHx5eNU4NQA
ddJVOFIbqPHwAGR/SOtX5cimQpWBrB6ffPgq8YL5zRHJNR8sYyaS/uJBRSIb5Ew8
kAgq0r/k3B675yjdRgrW3qJTaTC62EZ9BPq1yDg5mshtKrWSFc45iijGgfxJIhM+
swdlAh1Jpr9avASp+xwIZgF4d78NH+W9qR07NKupgHZrETJ42eWjPm7xNAKb98zB
CKjbAq9RtWYkfDNG0+ZO0eOVL/HZwpr1x8niY9AUPF0QSrZiN+xBn9sdwHWpzrpf
UbEinCBnLqmjAPpwqW+4ONDN1TLSngZyPdnGUsMtDkZObc2+g3XCpKf2HmMiXqew
4+WZCKc3ACa9bXVQstdO3AJqPTe6OyHCBhOIM+AfYsrulyyqNeqAzbYVnhbgjZae
DxvMVsnQUJHOFk8/zXlczgRG/EDzmwAyUK85DDfy60Fr+99+Z3in33dgZwEQVtOt
TSZ1ZgujsBHeRnGOJiiq7cw1KHCxt2EDU4+ttCWnDeI6nmsgO2+mozE40RKdtNIJ
uagJ/cQ+IPqKbQxE+dLOCcI97aw2MFdYBTvt2vU0lkiTD+GAfUuc0ep/jV+VDBt7
c7GfrZjSsD3YpACs3vUaaT5ZYnMspoUvy1fp9aUMkA3DG9W5KnB7SvWAV4nbu7FF
8DryNQDP9MXZXqqT4biGaXXAC2Dt98zuKiHqAY6aMrAbREQ5mNt/2Cdw9FBY+xLX
gcTvsdqkG6z9D8ePEXzKANMLAw/xMRglzfWRClWaD59J6pYtZQarSodjZAWcywez
El0tVhFxObl2wkElP/QCy/Z4d0NkkD0FbvvU5gQddqkTF5IsY17xi4ZXQxEMV26b
VPqDhXyLOFH8Qe8P0Y6+8qyYcUKYBFOSzrg7dm+bWK91wjfhPld8SKmqpEqrh89X
WahTzlVoa68AdHiZcwu9IRx5vyBcO3Sf1OhgBKdZDDmOM06GC2/O14o9DxbPYD4b
kdHcvoGt/DZpWj5gADTRNhXX9D0fgpJDZsfPtSATr8ZmfkdWftMbHKBtF/4pufnE
38twClmdZliM+mgNxPbLlrRZdnrFsfqot1rSp4e1yfl911W2oByWvbrnP9sjCKCV
2aultc+whMMGk1cWbFGMD10qc6Lj86CeJOdRR9JknALvsays3B97zV/Wb2TIsd8c
7/Beijps8mdw1EY9Abi07VXvvFv3XVoEBFANlG4w0LRgkzgp9NDiPH7H3jbNAk6+
YyJTG5EO67J2VXdu4JlyjpaLD/bBy5sWw2ezcwyD9YwbAVCmPmu1bBol40P8Ff+3
Q1fOvtQ5skuHNC/nj1N5qCoc9g8gc0qJgspnzCwpqYo39AFWcVpl8UbZg902Hbs7
CDLqMDwGYbjbSrCiPrOkbabUkZ4utqfn8J8V1jguRH/fJuAx84bfXCqjKxL4W6Y1
TKWDQ++3LeNYcchkTiR7t1VewLGT8iOHZIaoWF786NFF2jGZCjk6SlMpGkJJfO6/
KOzmRjQwHuwKrRfqYLnlapxfQfSleJz5nRCR7RJJJFhqETMegmZHR8reJXvUdga5
terwjva+yItgXOdGd7tqIUGx1yQA3aS4uam2csv69gLonYyeaEI2o6zDKUIoaDZT
g5MxpSnGUHCxjftLda93rvsQ/xb5L6eY9w9qJCY0s9EMHKKcqTKe1j5m7eXefSu9
HP6F1R2ZzwhZ0KCwfL8CbKyH6ucCNNKkda+Ma7oECPi958U2CslWXINSON4ia5gu
tHDghs9ITyDHBc6P+YTyoB4a5tSUc54fMLI2tyagqwv22rvuVqrg9FLbygQ6zdq4
EVUGCjn3lLVvdI86FsEfHrkNgHe68jtkC7+n1pM05Ede3a325pr/2puQ4SWetjK8
i1sA5DI0M2voqum505IiXCG5KMWgGwCbNxitsRLDnOOKovy7X6W5dPJNhL972P0b
7+Y7I724AJoxpZVhUsBPpLIT3WLox3KggyC/kcOlKHiUxAA8AQlwM+bprdcOow73
OfQyBfMm5PKALp/Ry2kCHZFRwW+aKrxjGIx2e5lAyu2GzC2JPScMeuoJ16ioAOL8
4tooDFjDvUNEjyrJZAo7rX0Kv2qrlfv9LYTl6IpjoyM8y8OGcwYPMSPP7smRVh0t
y38Xxbcxthykf83glUTk3ojMBBT1pg9lQDRrBMSUiBIogWRLaiC8eH4KQY6T99h/
tRMQAYcYSrMJW8jViGG13m3MwnMCpLJh8RQf9sLSFlBQWk5U1U1i3J19IL0Ijmiz
bhO+Rz/Sg7TRBWNrqWF0TGvoZOMJNmBqOR2n7vJstdt/5ZKJRKKvH8aX6IIRA2q8
FUG1tOedBLLSvMLRV+oQOHRp9PJBrB61EpAEEv/FSDDKMlhBStmBUIpdjU+Az2FD
NDM+sWOL0j8xWXdTjoJZw1qwFpUWWOh5kF/ykkxHM5ClmC4a320drv/Ho1PQU8sh
M8qptb9HODSC6kETXy6lOe9jkK1pz+gPAZ6Hd9XXrTMEhs7fEdFIzijuApIwFvAK
tzH9SNayQDXwUqyxHvfP2bUidLnwd7qf7fLB1Caf5HvwGIt2QRdF49h5BLCNTc3w
RKw1W2XbMCIzvEEOPBDjzKifKpyWx+pgBGOqpXqv6QCyPYJYzCT9AKkEzlwCWo0t
xQmNpD4n6h19k7kv5PqIU2c70PFNybDu2LAiqIoKW/neuTr3cNCqVv+1dFuJHYD9
gXkpbfsm8IFhOeRre06IwEmlzrbbT7+lfSJbZ+F0AcZw7oUF2nEDEE7RbXr/tdYh
f6/X7XLIcKjf5ANFq1Oyi3c0FchohWDp+LhyljVdenW5ayb/GNWEFCSKDFBLN8Z4
RJMapVhcZbGXdxH6+TsnslLs2VyqajlPCWzIyJZpjuInQ+zSbZADUdhpOchvnL1F
P/GXqvEG34vQUAYa7wN7KOhiTwHK2Fylg6eS00ubU0FpROwqwduQjh4nYj6imHjh
SItrbr2fIkTN581uo1GAiwy2B0APPiqQaymArrEECYiVkucs0GKpdKhYqgc49hNt
SzIJXOZOFQYMg5rt9GFn+MqhWJocOA/hq/EllarSc4aO0VFfu6I+vvzIhMQkn33S
TiOKmNAJ75bdBZT+rZVRZ3YNlKrDOKyeJwO7hJMPCi9XsgvOvM9ETnM8SdMMbHsL
PJx8ZebGavCqsQa+mYWMwNFygir06hR4hd+EML/mEaS9p3iabxFWr1d1i2/U11Uh
pkKg9toB93h7QXHaDcDhrRKmnLTX/9C3lqRi2Ta/EFosABFt+6lWgLbYcNp5f0RE
NDyksiy44uj3/CSt5+ZSJX991gRm6ha8KUvAxQ+kRS8EEtNBjAmxwG0T58j3twwd
PP4aTU3AKWdteviF3PkUcZ3MiHXKaQn00KaeevtSMI50iEzRBmfj2HdpExcRiFRO
wl51rvfUz4wo+25JofMqayH0Ko1MiDNKGPgapNADQ8EzMKj05TnLm2w77htJm571
bf89Hr5TzRh8oNaU/LyfiMh7wqKMYBOB3+QXyA8n+MzslvYBl1TTZhc9fwnvMAdG
sfAXo3JwMLeqg1ELKghjPqCcKJYyw1YYv+uWzJ+yc3vS0a5qwSrEz9QBOy64JibA
N8YSJXG1RX5bCj/H1rFoiFr0JAGRum1qP9XzzlPBFGP9rhwbDdLgXblEZ0B6rD8U
EcQgyIu57iqEGM7IiRsJ1EJmW4tIinpF+SmC+752lB8Vjduip1PDSSn+W8Agbe9v
2OUoDbBkfpFCwS0DJUGa+nAaWeiC/hulb4v+KQP9aMW/Tf6/A3K5EUD+sl+6llvl
+vF6Uq4YflzBmPFbsDiwoPS6FOetXouURaXpJjpnQR8E7QMCcjwz3eLboOBpyb4v
UBcqZa93yw7Eb+b0Ue0VDnLxlutXqhkRcviUcr7srCtxwtRRZ03waXiwZ3lmODvu
Mt9sIwdbY/mi/6m1QFC/xiSHRrWbmqNjMzYjbSxwlesGmqD0SeKWP6RGDueoclQP
MDMChbSmO7iaTbkMPTg5JSAEkaWgsCtgkDIzpMOojrbh+LTUNPrnezb3kOfkEpgd
wrKhDkNz75Qop4o8SZJ7L4PArQpyK7OIX947jWffhJt5AX5r0k2p5YFvF6SsDpqH
qhQTfFjbwY2aRrMtqAbxIGC2aqYovppkaNPqQQ6YkFVEx/B6lQgPhgrApzsBXw2P
9kSQMCsXpJNFT3qYbSG90x/pTteku61HLZVvDnKllyiKu70OVItdcovYjhi39RtI
f2evRma3W38tqxUqKy7huiTDq0SLpxC7bK9/gibrdzF9gKHYfGSCAvJVcnSjpBah
gJu8AcaW8dz47P2LUOmTw+JMloV0XhNyzn4s1v+S5QmCCdkWQU0mEFT7Cqc2qWB9
Ahd4simWe46tRDC8MXWEFbPn5hysV5K7j3xFMD7sT2c9tQsV03xCdCXVahaLDf02
F4Qp7fqH7KQ1xnZoLPsclSJFxYCWPF7RLagHB7GSgUg6RA/048OInL4CgE4S3hnT
NG+EMuyR2YMibxQA1lqaFCojhR9ube82ZxkUxyC9AQ5f/NPnRuEMcDbLE5wO3wf7
UsoTxp8TxD9swNULhteuHImP81O8WnP9l1uoNhUAEs6M3iPeRCGyrjS6YdUNrsr4
mtn8Zy4F2rGW0/PHDl1ConsJEF1BlV0L07v4loOhOH3ckYgAqnYCZlRd/s8TAAQ0
QUyrnlsQg43XMz3OaHTyQ8rJSLCMfQwVaH1Me5d2Y4UMZFsFnhC4tE1SPtKgNy16
fnHiNOvScXo1cb9QtkPxtiF9FPiPPg78bN2tflBVs28QDezyeow7hHyCQiG3976T
qYgQk9y6+Npe5HjQvO8qXxQjAI0V7o1yhlqqD3KbEdN0ksQHlo82CFYUuhkACnGB
xZZ9p8MbbCSDrjQBItOpJNtx12845xY7nNrgjMLUDNFFJCbQ49rofDkk8JtO075w
nWxnbpV/7lZ+KJndSNjCNqb9m6tIg68bd52077Q0xzw8CPrjfocvdob4Dqnox4sx
DCeRobtqW8SGQybtuICnhO/dXDFPdWSpNlzR6NNAq5qI43XwqqIP99+gUJweICGW
neIfptdUJATAk5WA/htMLhsWCpUKMEnSO31exzwlPQV8+Z4+Jz4yhNlH9aGIv8xK
lXgQt/wz2LmM5yeXet1oRRS3hxzyWFUV8RWrubPt+avA+p4mlgTwLt4oWI+pW8l8
JPEO13WnPczAhL52jClgDJiYY9dLUeYG7zdfspRoWNgICdMuJtV77+cWbuDQI3K/
PViHyMUD9sH7QvanYMvmybbFWH4Rrbwf4C5ryUi5l3Z52rtVldsDYx+ae6K4GjkV
DFJuROCjV86nsGJDXT3WeQWDSSIWNEblmMdG/KNYpIMUqfWeMrTXqZEwKxilGO7u
C7Ya8HM52T1+/GCE10eOzxwfIJlZYJKNFN48zsuv+X1WT9V1xlrOzOtRF/9pGqk3
zzHgytqW/LfaO63ha0nzWJO5k+4BuEQUeq742/ilPhYuYtLkMLh5K0OV+dPMFFN+
Kp+wsK7Nrta+DvdxuGGV7bV8PLvLlT4VnlQ+hQAIy6uZmpYARMzXLFzPcrCJq3Qq
VUlnQpcuA1Y47k/O8HlGELftM3YqgDcSR4VTAvui8saOUltxdmkvOtLmykHSd3d2
ghJmYAk7JrXHRlx+Fgy1UO6gyqVCcFpHWvhQGzdlQwGbPpIu6Rp34T5agFWq+O56
Enao4eoZM2HYH1Mu/HaU9dW7blr7WbLlVNzwOnrxpxtINxiZN9Essfb/Cqa+YuSR
qG7ol+inPtoNOo9SejPT2mFVf9kAxmppSn4PMDPnqlUzdlecO7vVHknjMdNgRANi
4RrIsLBllFHAEEfCgXjrxs/Vu794DAw28KvIqUCihMjDCloHwMNDFXzdNiD6ObtD
5Ry36wdtnnJVHqQ2sM2EUtMQOraNyIL5toYXchVY059rz01X0pU8RpRIC3nE5s6b
zpjLLPhvQcF01RSbzrKK+oDSXsAIycPXpDemBfwWbY/Y6Pa3YUhzJoq2Xcdgc8CK
YFRR2pn9u5HdZhrFznt5mJYNQeRrjPsvyHB3h5ZL0I1FjHW969Tj13LmqYOHNYIo
kc+5p7RCwmGugT8YebtTdanU+3Ot87eGGeH/XmZeJMq4T8ZOSQZtcCyyXfuE4TjL
5PWGXu96NtJMkhHwrRMRZjYK132//ryE5Sl2fA7d17gfhMEJVL/jA6xHA0ag1J9A
ukTzw0E1tWeMgBoHSLu8go/g7V4GkpKhOwgsfYVfjjpDkHgVy+x/5MEeCHJzHHen
M7VgS2SqmSLjb2Ki/uW5zThDBhHXH36GfET+orz89pPdxvM6LrVap+uZ0N49aTDP
311qW1AWydRtuKJjUCvMWkMgUchFXw3dByp4gParnDHfK+jRMDOwQ1X/Zk60T7aB
GFzh7T8cJkZLS2z1ksWoEbk63QeoD0NOy8TMPhTK+JiYC+OimNMTQttE69wuvkct
LJPApUXorxh/OetAMOC1CgV6wvswSCXi5Pgj1E2mBhZLF1AeLe9nE+GuyKnGQWDc
3YLkNb2X/CdWnJDAS8SBuge3ag4t9NcQVHHjaHbLrGxZIeovm82sQSlRVEfWvnzM
k9IraRkaSiQGjJ2ESdZ2G1mNctbR3OajY4K5JV+JQlM5jbY+8STstrFfbXOo8TT4
QKWbV/jX+EBLVnzKKk+R/YrlWELmx7GrmoEd52k4Wt3mazQ/9LBBmoPMFTHzSCzE
9QSv3VQ3dNZzVN32YeuQrvIR70RymqDr6pu8JcBYbsfUzK+yBhDRfE2l9s9wRlYX
Qk8kp7z5Z6U7hcwloFZvme3xp/JjqvHI4XVp+BEYXfPKkYB7V/qKl3PRE9V+cM+Z
yoPXWsdzp90afTsy3yfMzSnRktLwwU+7xzWGw3MMx1Jt3OQWUvnsjff22O+dctd8
Yf3eh6MXFTLQvLd+QVXUvq8p2uR0Tz0bHYsSnoDQS8nTLwoia3c+K0vGIo63FUTq
a+5laI7l7EqE5Y6ktd0USQYCLQemgDHyXmm2WXZ3Y6GRQm3WS11GR8RxiyJnSLaM
mooUhgn8w8T/PhoX3K4a+DcZginoKaEbYvbYlOzu5JljGDMVAh1eYty0N7wdOMJ3
U0l/e0VTAohkWDNLbI6Lg3tLFHQ/cbPgarvaALUO7nHTwVcsD78l3b/ISyQKyTDu
uh0CeQK840vJWFMnCVO7dlVzoIH8F2diWR2g3eycwKlhaYxeKkctLW57H4AO88x6
Er2Jr7gDXihstkK1zxPGz8OMVihMzI9ebI4A9VgMyJuUaBkqPs4KOaWKlJgEnSC6
ciXGF4oinA8WkgpMgT+jMTgzIteDJ1moOzSx8IizkkEao1xymxhAJzfjVC1JP9sE
Qis69wgEc863Ewwp467cCgvTvwbBF39/F6CuAIbaUfkwtBnnTjsr2dnc53EBY38u
Vimkys02Fjf9vcfnQWQCAQ4fYoIpjHX8qfAoMmSJSTYPzX3Lbjy/JI6DcMCWV5H/
cJ7Q9ul01uIFBq4QtQfHKUKRrqwuINoDeheYP+xQIbHNF1tGtAtwWqlHc3e5nyz9
vSRnCIGoh8zMXZM1qy8CgeFo411eNNgfMlir8f5xWd8JZp7VCSp1fc24ewA6KJLc
d+IRIFYDnHvxkVHEn1NNK77IDh1yMLUFe0iWP/8J/PL5AfJkNYvIZaIQFdbyoKfQ
vXVgR3cpuq+5c21oESNW+P0byXvV74WXF7NiFDs8SgO1hxqzH/WdGhfEPXUEMePc
30YPFyWaxVer7IiJkm3G/DiJ+iEvS1VgMmlJuUipXjbbifkoToW8UJtGjoJagyNx
50ezZRog6F+YlLP4XaTUAvL7GqKSNanjC+G38fYmytS4Z+lXNtJ4pGjgg0x2urmC
tnV2/iwlS4I+8YDXqM185pFPUVCGFh4wYbIa4xyznGsMRoj0/6lItY3294S2ElK5
0PccDqrLj+4oWX/gb0qmZ2J4ZFJiTS+J0XV1pqlZgYz/SJ1+nAqZs9GZyrWhZlAf
dH4Y5LklGQWcoNnMzCn/B+mNSbDdsQo0KksL4TPYjabLuB5icX4MjPP7hVYHcZGa
UZLdEGOIRk/k+7hj4H8UTiO4s9YET9jE1XxLrlfQSI/1jMjdbBzivvVtwc8/1FIr
rK7iouTIDTH1WJPQKJ2RF4U+e08ocSBRf2X6PqqdZhOMHBcmGzvExyOWt7tJeU8S
H9uKgDNcpWlkZYsfENj8+cEfUqBFFpHzrD3YHCTfyTbYlKjLagJVb3xqp6FBWJ8l
NYx/SUBDbLvOAM/mhQZGBIlQuz6tYAc851feRp8Ju+GXRjyOVSg6KyCToqsHxkwk
iBwGwMiQxSM/k8zD5UqCZW+C3/lthhd+94tSOqJQrf6GYQ9ukZlC+wrn5ARtJFvp
APXXFlvvLwRG4+Mjb0nJLg/hT3tCCwmtET79RZBzyJePCNiqaik5Jb+5IMwjoUYh
B/5vlThxYLDITaCcVZpQ0/hLpWgwx6z3Q+BwoR0iDAuHjzl9/9165kh1scRDTAS8
EeukQMe66MbjMRDEYSPSoD2UWuuAAY4ixSpYg+PsQMmLg+amKV/B6AUzSxLXq9fd
gTKXdNZw+3kMe0VjYPodwz+nZT05/SBxDOK1FpkmEFn0b8sF5JrbQZ2SvTeHRMiq
Z/lMOVmhkC+sMZHSDoKGXZiIN7+NR7ibWKqUq9mwZFLacmC9KsRixLQxv+c//3MF
bNR78Acuxlw57k+QVkXQU1j+GGZe1O9dX3/xsIKw7IcLshcsWs9FgC0jF9fFCOyI
bHuABQvwYEJtmnq49dt8u9O3uBi5tRDQvr8maZqBMkRiJiMP+Zs4Ybann5pdZRjb
BzMjdDL1idfL5D5qlShI53fV9GXJI5e06d/RZugzRQSOoziad8jOdl2f5SlpdFxw
dTZmVVYzhSnZ9vSx+CjtfpoI8ir6rtFo7irG5SDVaC3nSOInTzVBMhJngq6opy4p
KXkqOAqpn7DHxnbd5g75hvdrk2MvTILiwV+BVfg6blewYqW5vWEU8r3aiyjww7r4
c0cYUnBWbK9eUdjLx64D+vK67y0p3hwC0WqAmOxhzF3ww9WMFBxPOVwitCXu91Od
05A6BrmgnhbLggE/misFK2UovTP3adJcf7vxCF9HwyVkzZToZHi7pBqG3sWAF7Z2
PYOe3rdupfOd5qKNnh3MoLNiV9dh/qxmwhtw5xKW7xbPEOTPByabcjBPOquMieNl
PHgZL8Zic4u+vlRHb5BrL7vfmtdoK5TtOJiViAglOVcPOgfgzKKxZpgTI5BTK6SW
AbjAPerN+b4peSaM0zx0CfxB3LPIYtekgGeTo8OnPNS7n22Vv2XBpfcT2LhPIqqL
Ap5MGZwPupPEJakSTienDg3jczpmry3yhfMcsHvSvWjHyI7Av9A1roo4UKqRK4ve
VRGEmP2s/KzeRbcNPiVTWboKuERK8Anrh43JppIF0+uFkzQvWbfuJZstuCXxPh9x
zJ7M1nKHX5RfgDpYR0nVWWaIbjN3MlwFflISG6SWngBZg9kArjdGabCSEChaqoba
2cC0Vjxq7xctpHOy2rI28zawNd7mEEM/k4PdCPCn+0g3B9TyfS5T8LdNiglpspXh
/ojLBFx29zVxZqvwKcH438mE+hIGt0Xdt+5w5YOFl2rceFzAMzfA/JWHIvE2vtND
j0tJJ209RlNtvYy+2KOoTttwR5HOxO5Gfb7aO0LiDP8Vz1yogMXxhkk0jvYsxXdb
eJky4wGuOSTy0D2eL7+RX48TCuRwc7pCT8Ff00YcmJIN6+2bRxECY9bOl3CclD+e
/fLE5jse384oe6Imnw+GwiaR2FpPxyfhFrAK3U4MRzfAydaNkKdUV7SkY5we97u1
nQpv+jHKJlZUNj7Qq2c++0Z26N6TO7mkRFkijVvKi7r+Wr+ntB0vW+3vDHIIdGgC
c73M3QLK9WsnsafdOs1Mmf6FfqFNwrO4BIvHLNUgKgmmYQInfMBiU9jRHeAQAWq2
0IkqsxwQE7yQiYxU4CxqyrVIRLSxRdWwcZz1qg4qe12KYzYb5pJcjNEO2eAEEDJ+
QU9SJX/INGsjLwDysyfBOl+lHV5NDK5gB7gyOQ/Wg4phn3mOSlZy9VQpxb6x/mXu
INSFMcEMPWvCp66SYJJe11jpYWStxXMatG4XFJ4g0dv/MYeFhAtlSiQR9ve9Puou
2jsrEPZCY30KcLJGEgj6b4V30EEc0Q0CKHA27H6nw5dtehmUW8NDwQYwmjOwsSVv
lrdcR41nfMsvt0/dMRWJS8L5k3sLg+wMMQvzVWtgVuQzAbhlj7C1S3uBoEZ6p+g+
dnCN/M+MWkTRajOf2FRWn4bI1zgOx4ud8FEdMKbJbl0yz4xiOsFt4Fq7QsxJIeeW
qf7NGjL8A1EXWPt7CBLRAMlh0y2HEWk0eSw/Ux1lHyPBFwKEWVy0nN5xmyV7Jz2q
BLPfAUhIvS5yOivEh32/stwUk9Yldx24FNVfCf3NQKVKmghfFob2ncvOxB+0Wr7O
czDDhprMtTBMLiWpAbSR2S3aF6v7DGWypx35w21bILkVBBkKGkSE3XQJ/FSjl0+c
w8XNvOq2obXWy3OvzRvEShVUGgfDdbRzQ/7k8iOdx6nZqEyg2wKl6iU/vXZulB+O
veIXwtPMmQrzFwcktLBirp1oBJDihgARXCjknrnkEHYSdeAy5zum2nC5tUX3R6x+
L7Fmwcvm5RmZpWxE330DTIitlLICwrAkEL3MqZru6y5iU5sZB+a15d11oMfyJdRR
M/TgdzSQRYTrHHlLf0pD2WTBxmu7Xl5t0aPID4OESA8x0zg9i9Kc0lbN/C2ZsPuv
+y9SgEr6aqfZG6YGo19VaO9cOx1UwFqOT5fvymCuzPwr6a8OugDKguPqgFcEv7aS
Zanfgvbcswgw94IMVaqokPm2KvKBtDnTCiKC2ud/KKtDMGaaQfYMIGRPZpGBQ5lO
xRlHCCLnet6aL6rBshaNH+ykmBRCRY7JlnS51p6uINKaeuatNV5uKQfCQtEX0MRp
7khXOytV7bIE9IXMWmXMWMgJVqZVW7Uhi9UmgNJTrmzPuNOGx4c8AQLmLSSgQBaj
WzabvZlKEPXj36kNkA93dlQgMkO5RzmNNn7enPmvUK3AJe7uAKzMY6lpypHwiac5
VCxLDeOvi8eg3CUSRU3uZVy8QWajMGjqnURqAvBNrZHlZSvHaTo6m7OEw8lWzU2+
wUxshp5jevr4RJfb6i8w1cB5QFrj3cn+bamLEEdvg9+oArJOmd9Ao/mXDqA2aheo
UDdwAkiUB/6WPQk3e3F7mZrhh24eU4U27prKZ4kqDFasAm2uUZEPUt7wwhwgMV9J
JFi06dEjdwR9QEmcCHRkq7u0jyU2yNe0CB/xXVKKho8V4NXa/BxwTt6bq6W1HCNe
JIPIuh7SXVjmcIhLh06KhXl/OhxFioy6lQv9X92zKXAOVUAZMSr/GiNqPUS3Uozk
xNZks83VddQx7nDTe09SYHOvOoBno84zjJ0ghGGEbEeajatg7K336DPn2kmXf6Vj
+rh3WEG1nArrJOJAFKGb4J+iIva0L2ChCXpxwlEu3EQ+Jk9Aj/bd0o7gccs/kGWc
hDm9ix/aNXZTOfduccW6lfFIY9R3YhvyvMuJwF2hqrxMupFG6xuNGVwtjxXcwiMy
AFr3g725atuz9IRLbQAjnh0q4Y5x5BMTbdFgCuEtL7SrBNabhKp/J8llnx0Tvo+j
t01PyxqIioe9z5VCUINVGQM4/IKbjmXZBsQTqGmYo6tMVU0qsgZI0SwzTp9PhLH8
YzGR+Zh4t6EHnXkDHUE1wX6wWBvT+nd5Wy/hlaeGM4+4RxnPkzhJzzxEaj/qo2BT
1KvBnnoAPAXrXdsqWEMFHuvsTuGJHpidZyUFysjYyftYiCXFPkc12UmhWAoxag84
OJruI8+Vy5wiRcb3mpviVN9oenioLgpvMM6Nn8MMDCtAojFZFNjoKYqgRnUyTzBK
IZPiCD0f6jnX5wMnhxP2zNdgOg2xo1l3koiK/hxZJexzJCnT0rBHbVAP5KMjyhxb
tnSOmyM/RuRVNPu1hR+W35Lpdrt3qo/dYviT+bes6E7FvKHXMNAP/O4qxf91Hj7p
hAtXsKwOI4B/3Bdr/O10+zkik5IRB98k9lu5BK3EMWg36kTrl6WhLvPLxlLOZIxr
blpxmNjMWiYbYHKVdAi8efrNZPiBrlj+1d7RTSEnHkswa4/3I/ZZ8c9YCrW6LDc4
rhbjYESy1ViQ76A7EtCYDPgtpeUQLxOdLYjYhbMouQQwOiZOF7f9cN5oaAJmRxvB
V2+PB7q3crDDQcwl0owteRKjt2PzrbYmSiHDVNUxBLZnEDQi0M1sC9f7w4teP/IS
89Rj78nQDOmM+YotNtB3Pi0KapoPyHCv28Ih/7ppqsRWdO6fqvVwhHTR6ZWzZ0n3
3h0kMAROvnZFB2Tk2PC0kUegt4GB1J4UMn4P+eMOTm4U/+uB/5dTBYJzczM0AMpz
sO/gRPPK+eqhucLJ/jxkW/CvJvHEF+9MnjpIcTn/iWZPqFmSC5NRacbeKvp7gp+t
6gvvhSejhjJ19nfUHY7oIU2ydfU3OmifCgkZzppXlhUFLMRMvH5piH2SaPqt/fET
8L6CDCyNe5EwSJ3MNbIX2VDf+/RDHDfXmoW4n5p+vIfkKOjf/TUWrcVi8SLmQDeg
znvAa+K9UCBULeZeGzxkLSxvCSi+7AmLN43crtsVNurls9h8abhvMzgvl2+3AcPk
1DSO3yT7R7egifaSWTN7yjfjBN9XlRJvd7OR6SVAJmhbaAwAXKHk2/vg3J43pI9c
r+V69evcQp1Qrul4k+wCDtQcXaZUalx/krUTKQ0Iwo/kXryQRByd1nmK3LP32oo2
GDTbdeSdUDyb7HTErNFXZfiedfHurhd1nwb0g3xcajSiGS21PrIQej9vaaklvnX7
SExwv0E7MH4fR0BX3/x7XBzyZ8hkKA91UQ2/TE1TLqlnEUoKtrN9LNywVHZaU9+6
UA+auF1mHbcgO+vTU0iboAxf2WRN1+fh0Pn019kKvM+aaMUidDG4W6FfvnJXGHqT
vKRKGGLAFqQ0k9Y7h0KV6S5SRFJ6kLB7/kbJg1DKKLo60UreN0s7Sfb2m5VAadZJ
mQH3u2vL20+W+Ryglb6Alv8ory5JD8Nts31d9Sd6v0c64xmcieBnUtHRIFrVgvqU
IRQloZlHna0/QWG9cYu8AwladU8QQ6chYNU36WjnB0fPvOEoWco7c2rUjcvMIC0D
3YX62DylsE4PPAVNrcdVmF4R+apI1mrQHOhVrfG5DB5H+y/26YJI8o3A6gF63Ynn
jaM+R4MXpR+ZKQMOIOozgHXYKhQwBq0Ix+dU0UYRFo/Et6Sj5eOu815t0Uu4Fgmq
wwg+vCa3WouI0OWkYK0CxEdHqvqVVk5tzUIEARsp/qoLBh8dqKTNE83IqVBqnxBj
D4DYmC7XL8UMiMRcWmom7L2Tc8Zp6qOwpYK6OdPoJ4qcIf0C4fG5bjLEiTtEFpzf
LX0ebLwlIZwcEqpDmI1TJtnlPXfomUy7a8M9t0WjFGxHNRS7zZcHKkLWCtaHE6is
5eTpZPGlq7ThXFzmD7lVVPdE0WT12hyTRQZzWBkWwAxzBRgGWpFphYUDSVCR0LDx
w6QqIEgDcUJ6CDHGWqY2p+Qd8AAplJxerPHsXpi1egBrG3kkyhUIdHLO0jnbVBWY
8a2AROh/QV0m0jPoeHv1dYeAjbILnfAttGHqeIkuvtj7p6lyhGIns4VzGWJ4jh33
U02pqGkK3NIBG3DAl52XGKsIMP4IlV/hPGI9rnIhnOG13HP5TKV5lvpRh+lJxYEh
eLp8G/czaCaQeCeeSLMTpcm0p6SmS7vixtvasFIjoRzmkkITFJ2sKN+sH8MoXxVo
TEIwEzqC6aTBBGIc8cZ6DQjNm/VI4tFvOAIB8noilKyhHnVE8wc3D71VPKjt1sQT
cv3p8zXcJUl7cbdoL46rHPCtGbc/EelAvs3lH25qYbDjlqN6Oby5SjlFpnVWjxVy
OuggE2kP+ybQKprSKThuchDjBVjUUBctPWuz/cJf6o239rO0KKphhOin36AKiV4w
QguslH9AR4KE3tUvXRmEpJkyAV70z7pBEmRRq2H3XDfpFLkIWoEw4lEh73E+YmfR
LCDMo5A9APpRgoemP5HaMs68hTGZxmfwhIuw02HzpDHQt+4sjre1vsTejsPi6GT5
qcrbqiQztTRS/K7THEOM2Vl1dTTLK3rT+9bjNwZlF0sFhcQnrR1qc1H4fUhW08bE
yatxuKMBUucU27Oey+O2m5CM8q04SZB/18HXvqwRLAD4fiKOMB2mltQ1HMOzwc5U
6aswQgdPtzBId4/FYXWWdot4YBS9u/pur4CXbv/LEafA1PKMcty9KU6x7xo1GTb9
s/vl3sVKfLJ9mEEWuovqaa0ht0kXdcxn+M7z/KQJSYy7m7t3v/XhgOFiHzinjtaQ
LrWvkpirRnxpt75AIP8bFKTxLgOsjGFHzL9GrOPrgZFfv0ZlJ/DCmA9gBmvcitL5
vKbdpy9GSZlXzKZG860syDc72yioD86WAjgjppspiM43OimVPeN/DsTJExDXXWyy
fcxr24RlOBmj7oy4qszo+YiiomE4Zr/qjzCkVdMoiwYaS0XB1AJZSfCldKZe5JGa
Um/C9cbWZIOkOqYtaZH+4H6AAjFs5DOrVLKRb+Erj1rRjS+Txg7eKnuC8fP8vwTl
oWoOnYyWPJY0JHuS52ANrm4lOuur++dny6/cMEeyzSh+mrXDNWHRg+6AEIbox0QK
PFDR7RE2kiJzkhdP9vFoBStlF/gbIvlSo16dSXV7wuIdrV9wkihSLSlhVSCSVklX
/WOELm2bnjpFFKm8xzg1klxTO2O0C9haZEh5M/tpMP0wQBGsnA8DnKho5u7tN280
+2Z8gHQqMeH+ERbV5kkCJcM7gqqFpQrY9ekvDwVst9Jn7TCOjzp4tZ0JM5nw7RO1
ls1CelE+QNOs/TqRgwpLMV1JhBrVbhHIsWa+lZFU/oav19oAToBDJ1W9B+wOE2qe
jlpxUbYZQmVfVbpIHHTEz9XQT/iT84RwkJ/HVNXtHlDZpxq5+t6qtB0JXzJYV9yX
SXg7/9Qxk+OAi/+C5A0fPNOT+vLghLpZjzGfWOXcs9nQoc8BQ1qFuQo9HNjDzEP8
ZSD6UOMlY8pbIKHY9ZgRyaPMZdfLoRnVGkR9hyzy6BPUqddnKuXfSWRr7JzL2ibN
0aQaKZMVHarXaD/gTbvkSTCK5d58h9a3Cho5QwW7zkM8oLohRqY7aODf270z7mpM
oamJFMDzNFfUIZ5WdrvFOQxa84EXH4xkITw9oBGraw3JwbNoeYyyjam3SpjK7Jnq
nXqHxsaJnhoc4O6p0yRAFuRsqMQGnYbDw5mmKmRDsjGqU9SA8izX5FrCL4aYZwDa
4la8hKO446sqPVSvbpdqSoPOPTSLpRiKO4e6DLTBMyzDeB1YSmOwLqj2xA4abBxY
E5aMkPqzCJgw1Zpt4rmuhiRhQkd3Il9E2ACUvjsL+YOhDszvRN26W2t/1G/5reZ6
I8ZD8PnhKEATHdxluDxkEoGXkKCKbm2WXdW9ApnZ+yQVo7ctuqpSaUFf7xEbwYbx
+G864HK+T/DVYEP9/FvL9l4MgxAxKq6cIbYHqif8lKJWs+IG2U/lnZ/rb+5vzK4/
O5Gv2nTAoTvN1LZZE4X+RTJA9lQNpz3eVMeSIbd1au+dvwnCflfixcQ0qUggjqpn
w09RzBDtGgLYA87RrSQhLrzCxE+Nna17sdt7HUc/W1huWR9ZVaMspoXXqjQ11xgT
7WDsDThLTUw4Tl/4mN4gkRPZOLIbYsmX7StKirb3DPuch8U/nm1WAzw+sqiktEGS
x/OY0hIQPAORnpjLjxJNHN7ktDyKIivoVC79JzIDwi4kF6x7l9FCsopRbGgNRewE
3xvJOAPl4/+4JmDgaazt0AdLPE1WWUlYwwDZh08egtZl5eLK3XwvVx1osAmLjUfS
FeAaay5hDArW89gwJtZbL/9NVbg8n2GPHSlLD4lkz16A0Bq8aaL0Fmj6vqLeUpqm
MxgyP2PEzHQSKn24B5pp0I1wOUjEZf5A3jRJwbCoNUWB3g0G+uEjwQPv/lFMfyBK
RR4MWzC2WlboTFguo4bVWpghQ5A07eDco/FOMDjQjHdIt5Mk1z5N4Vz8CFaChBv/
xSNpZK1tS+k/+JzPuOiMm9bXZmyXPIi2bkZTOp7ObdFHIyGf98ElOnkeW6/fDgn9
0Tlxy8LWNudB8v1voHbq9sqqEJGxCrvXJrlkreQVvZDri1AeVJ8qyIRM06FppNQP
81xrooG1iRrBBeqisZIYr1fN4/oMSzNmvXaM54hxf2OG0frIbpiIkhqyBffd13g1
P1nmZvHSl4eqNeslf5HWdvBIKDHf/4uzNg/MyzVAd9k5w00/OrYqxO99r34bAV/c
zWcu6QGvcaOI7UxfgW8rzgnAgUgKd1bGr6TMKROpcBZw1mz7D0nxFwmJuceJyTYW
yHJKLWfM2o7VCqkuTiedcppdbHrZqhGxRfKoYfuLqfX0g2hkpUkX6WpYHtLl2EMt
PHJFUS5sJAct/J2Ku/WWrF4acJhFaQEFS4NZyuOym7Of3KgYTNM09L1jjTQYtdTA
rQWCyjJn0D8uGbLY2LgJOXaloQAFTpN9mYRQkrFDHXznQVfaqgAaQDWGmI4+V/u1
sr6wEj44UR9R+ZNOY7eQYN+PSPUJjiTdzg3EVHIgiviw1m4BFZI1zyMwppvV3b29
IIqpmP1QbLarbTMVb2EFVCgIFkK1zqqHxY5ugiFdkcybgbRiGEVluSei1WabaCjy
W3cwYBEqVrmqHFZUEPxkvS8WxDS9uRBwhTP5v5stXjcPrgp9X5XOaZRy9dUh5yq+
Ej5xhOi8dkYLiKGANti7YgjdxkCIRQGNCkTNjj4J+mXPz0/b9DmjcBgC/H6YZ7Tc
e/H+a9zUSB8FgJSaPqp1CtnBlz+h3ZHtYv9mH6dtWfR6qHB3blrf3y3BbaJZXGBY
srs1UuadWJs0opDKJZ4tKlGPQNAhzvaSCu8b6AhaehOV0Aol71eulG4lCLAZNsLj
+/kEVCOjIHM9mQSOPEkrq70f8iV/UZf3Lc72sqTOk2q+pwxM/7cavhzDWTxpMVxQ
wlVryjZxXO7Hk4qgSCGwaEXkyB/hFeObATCjLgRyv4CLCMK4xFBeQZGqeBWdcHqZ
qX1/GieTznNOyxpblRHr+jxxXmjpiwN719/JXV/o5l3cPSQgjeau8s3s21R6x1h4
sScN7rFXkm11WJuIuMHQNbaUH9V97orpmXKTlWuCPc+aDQ7QuYejQ3lXuPAUtXBm
ogc7yeI1p+BFZikBzC5O5B9vG3Yz3PaX3+UwH/5S4ovBXjHdRLGlCqP8y056j+pf
QaBkjDFLJkZP7JayUJVdcf3byGRe9QZDsyfjm8A5bohQvDWZvmIY9VNo9wqR+9h0
Xb9hQfphAMSofv7Wlo0NKR1vBKeSB/dxk/ReBYra75wuqsv/libVT/g5XvS6xr1R
NXAMDC5KOOn2fR4cOgZVLL4ArL+mrec+y1KiSO8ge+cSCTODPnD/GmMvkUlisDHo
dBZBog+FCWxoV2nbS3teBvZef4lvYF4BwARJS2nfK0JNm5XiyqqltG1sUTALqKz/
0Z+mQ31k9p1VoyzMAQEaDARzo26ZTLXdJ7J0idb9sj9uNVnCKiQ2O+DuJZb8iPfD
JzU29wXMr42ZMNUrjaBfAejBl5R1PzZNeDV77oAxSDKKtop6356ISJxT5hIYEOsJ
UCPiCCR1kLaJ+arUd2LWbD/m+Oxrl/en2CGgWMY0ymvv3rBX8memxz7PKgfHkgu8
Xg0zD9YGZjB6Gl22cbN/0xGDFDCOHBCJDqI9BUkR2mv9fgX2iieWtAuEAjo4YTak
CuX9EWROJJ9FwyVyObjJKrwYlu3A5d48Y5IDAe7GkzTz3NNjJkd7lD1i9SUj/Qfu
Do283s+cyeMgjX6clml6Jcl3e9sDy9/sxQjpOaK9VWzDy7x79ibeNZUWclKE3Alc
FzdSyILAQxVg8pkm5BWIywxUgssNHOSXfDvV+QLukW695Sw9EwpBJI7UrpscCEdY
Hsy7BTa2FRloBPHbbUV1GTVld1vpNp0X2DyFq4VnkcqApTSU0C/APIDqmEIuSytY
W/ltCYwNP2v3laDDT4I3xXtJE34PugtVYnAGJqW+OA7GQPDhEomxpI9t5nMz6sWB
bwwBqfJGf3rhpGufyVJ5g+w2ezN3sPzjf5OPJtSmvha3S2RnJ+VHqhlvK2eE9X8a
idvNz3ivrJZhuVJQvIsNg9j6vR0q0/rUQtQQv9bZxMmuPOWmayM6YTDdXkAv1q64
8GER/9m6aN2TWvQmYsjaij5mXuEyrLWjC3PU6VmIO/SBNnjc6xLNtpuk/zYCwNQE
zNO7yXe2PTBmKLuKn/i6y4neVXyTQfrzUww3oCGJwNRIeVVJxcbLMXxZbHJxJA6+
X0i7brczK3fcnRonSQKb4KYHdgsLv+9EQUofa2nyxGqaKPY8GWv1Ojbiw2HcMtCc
5xwjmmG+OP/n1m9G9ZjJbFpQNAB0i7fg37ct93MHDIRSl+/2lCg7Vx6vfTyUVS4i
9CwjkvGY/ALvSdvdc0XKXFgG5OMJ8T6wRErr2VPZKxRRHKrt/dPx6XDHbxYgBD4F
XqW8XCsUPc8WSosivHUNOiOs9bXlTG2Gl7yN6z7ejd0pSvbLxrVuMe4ll2W1ji9s
Wi8q2xhKglbVKPJuP8qD90krBKbbEYjkX/h5Be9bRZsxp2x9coXEgIKPPoJbzdax
0rwIFTFuswO6Olx+PwXAJRmwEuQWYnfNFDSB2wFMh6YJ8sZry26CcqcKun4UnapA
NbWzYBjbdH9ywcutTgP4F2gUbWXMlDbzudQ1vTtuXvuEmTpLpsfSuB+3G6T7UvWU
Ig2YtbHGUoLuWpJ94sbD8uogrNLZmBVHxUXXvQNSo4HG4dJAJRWnQ7lGYioCaalk
vuBxl9F0RboqsoxAB5qUqkIGOmbo7qyZ2BzS0VUi0lZCWo73KKDaAtXQDrK8qS25
WPceQg2WrX1nZt6cxvaR++rr70rlbFSw5F6pQ6q9Dt9tQSBElqWR12yZ5mnQcmQj
UHJ15Ir837lj31JjFAR5T9aCw8UAbRFSWDURDbh9Y8OMqUsHqsfTTYeSM0kqEc67
OU5xwWwDkHUAZ0Sv8C9c89FD9xCSG4opbkLcQOHSW6Eyay3fgGejErGhyXSQ4dPy
05XwBq8ELtM4USEfYZGRLr9RP5XWcTBhuHiJQNf2PkQduyua2NhfaU1ctZ9aknZL
3/xP0mwH8Z3DK3RwzpOMeCxH1Vb1zossvKfALxdQuSrNJ0kLS/RXGM/IXKzPLCzr
d153dYyQAIHc8vw2hBRDdqQvRotdnMOKQ1hEivglx/mdmEWYvP4NH9VoW+JXJQ5v
pFOHIMlVM5CTvej/Fku7RW89AtCvD+Lvq1AEjNHmplIVwIJZytv4r5gmRtPtXAXO
Z9pnS4bwn0XAZw01607mDf2Cpz/s4pMd9bYWBHBQ9iXg4AmBVY2cgDRSXmZCHuvh
OFtZfDh6VZfx49aWawX28IxmswhSmgA5BRgpE+GFvF0QRfRbAOjJ2oJ+oZkcP/Np
9PYtHxrb1liUGSLwMStrIqMWerL7Vjsz0WFsQ+Ic8dKHAzKSfCPS8pzcJQRhUyic
dQ0kV3fo74O/GBAqkBtZHxHhjHm5drcYq8yqV4wUhSOM8fSFo7p0fFxYcVZ7c0MV
sHkB2NhvGANl3qmqPqjcyddTFWgSYBEcTRb5F024EWsC0nn8wfK2jUvmbsJ5rGxM
v8kBETM8sCgq2f67njGHQgnRAcofh8hRSPdee0EYGpn+VEtuzxn8n8G0LT0FGyni
zAkEb5o3tul3ZXCWIQd4RvDNMVO4DWT6VuI4FAyC4jrE+CMCx4IL4gtSFL8DEPrN
mgdcWmerHG1Qm8isih2WGA21VwDRUPzq0PkgtAQ+180ajqOQMvgolQQJlPlccYiA
RPhIV9U7+y7l6fvWtJkBARkM/Zf74emPpr6xpP+MsmZDebywlTFAup+Tp7w9iyOm
T/nexDXwWkQCkCNNRD5VPrnyzp/Wf3zVV7vMRK0MZkWZBDw+52SnsAX+OGABZEoW
t8CayK5OKs6ZYxo2SzZkOGGuHfkwDD+J3SPmkNUNVq3hvXhIKpQsFDdU+BtNB4BM
/HJbr9YgkHJ/lvY8EWfP2D2BKsW/wunPqU86l4aZhc/4BJetF11WVOK1HmNvEy3T
9ZeruKaeAz5NP1GDNpzuZtqDtj5pNPB9qW5BRlAygX9aepBxQ9yQBvWVqy4zLsYA
vD+/2DJv/rZ+/lIBE4CLwyI6mxXU7UFLHQzS8lxPSf2wDE6cz9PpgvQ2074litSz
LnJAp3boYckIoNlCggsKXeX5VVfVb6Cim526U1fhp90/EbyiigJvn3EzfLbITK7s
2HYRkKnrasy9RXjJ9tbNvqglL0nNuQ86zuH43A77UqGwIJ7jH8pgZGj1QD2Z/PPJ
j7QMQ3LMrKjK6rPuypxTEr2sWp1kTrjsQEnw0BTsEtw/UITjUV06uaC245oXlHsb
xk3XC+84s1xzqrOGAHh7lFjDdt8HFA0BETK7uW0lSmLmZUoC09CY+XG8MfHcuOa9
BlcqYXgDZxZVe3rBet277bHswaMdLnYOeH+Il97S+WDlH/Rqd5ZQk1HKGzifZQwj
w7pbOMbiX9Wnu7csTRfx1sQWzDK5KeFV/X1pgYTurflejZy2JPuuLF289sY5yITe
nz+5zmO/qe++q1pJCiKNLN8XOjgrkYFQuhUbS2OTSDflo02HQhWZ8kVIyqX6wVZd
IdjpA5rZUBjGsOmibosrHsb41BTVCFNT92doBNzq/fkFQBcokiLqHFFdSoq5BzWn
/ijDPuxkuRxAl9iJPqZtA6dAv+Wkf0PtfSoX1s8A5PqtF/clsPnkKkesMjG+aknO
22Ijtxkur5hDTS3yTBZT0HM9mfYzphf1TgprR7fYWlkTNL9KgLzWa8fCoDRSJ2b+
begpymocvFa4byUlLUyjObb1L8UhLWXje8kSlF+5XnPDrPAhay6Sb/u/wjRUpkkP
8DmjZQvoYJzVUPVpyb8Aup/DgMAtBpndeUXufXGMEPbHqSSNY6ubZOjdQqlFArEr
A74gPyH2Ofnd7VaFfMEWD4lh9KpTj91IIDUb1IJlV0Y/o3OQoKGHKDBRjiNCjy6t
LXEPSgYR9xAMxRR53/RMJbYr4QLx2B6mzu4aI9dqR/F7lZKbTxCN9idKEqPiHBTZ
TkA5px4hLE3OM9tWlMkGTrUyzBxVufn19muVExatNtnUdxn6+UfU5or23gHJ9YEw
ypG77yTlng01kCKO7lDxnHbFegUMh+nt5GdoZqNXf2eb6E0Y+F2Hjkyh4ZLkgQNx
WjWkW4wWB7w+I2WTuKyV71NS5V9IwzJzcBQfelW+QXUF3lcVn2hpsRTrDSwGDO1v
wEgviumD3Nsk4hn/TX6deVJ8tAE+CUQ9WUz1an1C3MO80AHlUnDZ3Inz4Mtekods
rrCeaqNlhaA5d828cS3ZIugoVQI+CyifypIy2n31PsrejuhwHKia2qIwCUZiV0cN
ymKCDpv+W7saINUvKpKj299wzYtg5eP94jdW8S/qxQW/bxYKUIqpMwjsWvyXUPDF
TbIxTq27+wf1m/PO55pd7jJlORm06nS19mVFaM4lW+fhYE1yIgNFjKIdUsccKX1A
UbAKh/kubbjj+VxPDrvK4SnZR2vH/ymQ0eFpo7Byj1i7COV8s21qxU6KWbnB9rq1
byHsc8KJv1IJFpS3tvaDFpZAu1zo2p/Kkeanslr+KQwK1O8snJ4yWhmf8dZSvSpc
95RNYN+RBZnZjuHmfP8kXXUwY3R/U2Pv8LzjrPziJynI4c3MA7SpDItLRqKuLkp5
hr/0G87EAgsIHRHYixellbvQBum3LIa8vfF9IkGjitZJZiKnWZOnMit2eQbf1VJ2
qupXaWr5fGGWcpn9fEj8CVPwppbWrFfRujq2OOcehWm2oM2fMkwsfTuINjvudde/
JYyzyvqdzl3/C+xCWMHIYSzM0yDUMUmv4hzYTMb2zCCczeStP5itpFUqI27ebHT7
pQ//qHtgujj7vipxr/PQQWoKHk2uSjxJWhamnCfgSq1ZwdVfwacu0VoxsQJ3ChKY
exERY+4+iJbmnS7dwES0TjK8dBktotKCL1NQRThnBJYrBi6x8wWXEqdmikDqqLIR
5wSDNYUGDnMtd45fF+Prp83mMW+kbQ8ljz1b24Te81Di+SILn/5ch1xfCv3nSF3b
kou1WnPixx6vL/BvIwOR5i0axDkDDJ+vjLxlusB/gn8NnoX/IEKKYQc0nLI1sbxB
E7432lETFc6Ff7npQ8PJDprDwMk8tlbrMxCyIi37NJurOl0gbgm7neyhs6gMaNgV
970sD925xE14TN4CDBmHYUE2CuxhtyiMH3rn8yaczfqbVQbX8B2tfDOvIf/oOZ7Z
cBRv6+kM91JGnK/9KnGQ6CiwG6gFF78iiqmo6Gf3qK15XOPUmHTlRvFyihVA+R7Z
jNfdjqYGnBtTZcBBGzIoz8PmK/Ra0SitoCxbdllgVn42yRzXK+ZaQP+qcXtCFzWr
2EY8DUmPzVT4yJ1iUQEhm/JGSo0TRB9tzyWHNk2yO9y3TRaB68JzxisvhhmXgant
jtjPZzFmbHIMrYu1PoaYKrgQnKy0EtaWufKFIjdtHlUIC6QrunboZvIRk1/0bH0n
wG40jSOTzETXoA3HUxipPNEQa3+peSllbGh3E0QZuwzITrTxEVZQKMo70KZiSWPU
IAgVYeBHgCAOoi2X2s0Y2ENk5A8vOTSPsEo74Gvl+Hqt8BTL5HjMwdqOcJhbK+Lk
QFgx/Qvdx+zKtv7K5W+mvkInh0G51by8ZHmIjdh+fyzYLgvNBt+F/VhXqvj6osVe
2SvkwCf/0HWCPFr7Uaa9ETZbG04Y8WJgiKtQgRvMP8UxzYJaxDXzeIt38q5JEXJm
HEQbYdE9KcPveaZdkkK9yKfQcq2Gm+GMzluM8OBgz/McWSg5EIN7K+8UrPRXqVL3
rBKtebfbpFVQ5AT58vtXKGSro0Qxip+4lB9EaxhP7bYWCUXKC/UWOHBX6Rn0SvjI
OV4Dp0AzlXfHlHeqP0m78HadDVIWxK4jwRRSkbTeLxB2mD3lFB5CZXvEd7NL/Z5M
YGuJUtHk+mAst+L2qQMGGNWCbkcoI0N9VHeLKoQl+lMZjZ/UyjOvkL6Bc2vlKMYT
QPFKEk7mxQs5/+9d3JHW5psZQb9Br9ZG38k28CfTiihhjoK+EvJ1eJRaTFYWgfzG
C7nMnwNRhpNSJDqjZ2SjZZ9Ss9+612QXlqAo3md8gO0XYY1tVjM5Y5lxhCtGVJVQ
9rGjrZBeuGXX/EEp3zx6/ValCoJFJb/LjFxnOUtVn9wmduuwGZSuRKqoqH4DHB+4
6XdnZVcZR699/PFqoOiAf0ANNF08oYkHfSS3p2UGzpa7BweGevIA1IfsosYqw4Pp
QhGHhLINkzOFAADwhdKMVfIvqn7JkErJDopt6GnK0g8sIE/u9sBHjmwYXIy0pck5
Wr6++dH2yUnpuKXNRzl8FYVChu70IBUYVsEcuHIroG8+AmcFTzxIaVOrPWNIGM4V
y0c5hG02XxgwFQDr9e/TdRzGR6Iypj1B492fvbk2oN0W34Omqe5zbIY5QLFMaWh5
Arvp8yiJ1wmnTra5T2zqLpspxSXjsQK/Klb/28ObHbk6MxBmWnSfpKLqtnMQ+f2A
GbbZPNDIvkxERMglqYUyjHdsFmhppQQQol3LTzANQwcKggMp2lrCh7/ifUyAvVHJ
PYC7Q8Qx/qiV6oUFh0qWbyTN8op92+bmb3xnJBJAc18wobyGwtOmnP3zlk+pxYUQ
x2DwxLdchMwAJ/MPGU183K8QTi8Y/hGfWtArTCdaX5d5NlkKO/Q/wVfvlKXy99qD
ubjCoR9no5tz1JOjAU+vsj41JZyktN+8utEfOMmOP0DGwJYSfxutg/d41X0+PQps
cc56cxAHcKgqw8KMoO7oBQWKaQdrHFawyO4crrupw4+t1UIsgLaE1nJ/AsQ7nIkY
9L5NaGUux4TbCRZ1ZB+B96ZaZgxafWdbOrTMrrepxQrERYJltyc7ayg/oqCMAU00
KN5eB5qe48zekKegMzz647dklqb1adfLcchYxL0+4KO8V0nCF5rFceszxjW04Rff
+lLiCPpHSgV77eKSF1JhliPS1lQfXZ2K7fFfxz8KCgd0FlhPApSvdpZca5oXhl69
q8qqpke8ibBNowquwDGHdIbkzgyQLQSEXXw/HakkckJkdGaoMKNp8Wgesr+Pn8Ew
To6q9bq+px3NKVZjY6oNMtzNT83QUghYVh6XTSTgdRcmE7IRiGmmYZ/kSRkJi9CC
XacUtUd0HLePaVO8uh3zbqPj9fc+/Y2jDXL6DEiXvqhsVxIreBBhsl8T9pctCu0o
yFv1LWefkEf+A65S6yNkw7WIpcH1yPxJb5y9zW+L99RzTZ6SpR5gZ+MbI57fHU/b
Oe/IqWgSuNSYkEt/gk8XioQeZFfLcs4loBQFBDwe5tC7HL7spnftb4KZsgL3RYr0
aCrCu/PNA/FOWdejES1sQ+ZchCw6mXy3AoIX/1jHCZDkhCByXonoqUfDfup2hs4P
w4fnaFjhySCqo+L4r+3eZXDn/5ea+OkwRx0qUOuSA6/R9yWMsm0txO39jgSZrmi+
p7N3P7KPLHYly1Og9amP90KgQaPJwTsvQwFXzTJLyoi6EAzfKp4wu3Fep9LJoyeH
9MFZcANyp6jbtW5F9TEIdFeuioTtgmjk4FVSpVwqWG0S89APRu+u3Ltivoe8MH3C
gUe8/SIlXBP6ryQTnpS4wwNhFosz94d3KUczKuuK1+LNSevujeUNN9Vh4NJiz6iK
DnriaOf0k6MlPW6Sypnpeq9of243FYV1hqf4IVLshImY/SmKuc7VTT3Ir0CplhwM
S+prPpdle5qLkzK3FiWwjv97Vvl5uzjgMGIR2t5W9GninQ3mu/Rp3U+drQcHaggp
Gb58P3DzJ2eR5zXf0ehNGBhBE/inYlcrMiUS4xqZipk9/6wz+Aefg1hrBUDO4sLP
5GQx4t+FoVwRXHUdEOvCO4ocswEFPEUKjZfvGnJqKS/fid/wqi7iuISQXWitSZhr
m86lmAgnErDBtE6WLUbhXl8aniacGwXsvSck8QckHWgR1jUVmC7tETVazipmC6gI
hSjrp8aZg/S6a4+1piZF8oA/rrHwVz3+R/UVruJ8RQz5PujNLJeLtVSl71/IYVNr
smIfvPviQe6YjrV6BsLU7++BAz4JZx7ZngE37O3HeCWP7hg7JamvSmks2OH9k/QQ
GoRN7NriDmc9GKLgy2j6bJrWhxrW+N5FFnEyVB/w0skPW3ImENCyY78k0IwlXT+S
9rGBpADZob4dj2q/9Ln+Z9g+hpL77krBpwQTP1i1CXoMip+Uym9iORoIDp1YCA/m
sZw5n/5ltwyxb7oQtd5WeAwfPG5hFMlrOVM2kp8USWSvFXjBkFAkgtDPWmRnGJ4z
SWYS+ch96RTvVfzLb6eqaZCdXeTL7dEPFk/1D6qEVdOy45O3Oz8fYuOvLeVcZf6Q
MAi3ojrniurrMHEyMVDxtMDebS9/KNOf7rrIx8GaIEq31XXxGIPFH0CoB06b0QV/
WgIkOMIfIBhclEUrOCc7rrvNdCuj8eqJzZQBK793mQD9sQWnOLIX86Cdvx2xjf80
TP3idb1Gi8N6lHS5PjYd/H0fFF6MHsUyPn/ZqURpAbJwXZttn+7gxY8aS4L8JEq9
wy+ehhLuUTnT6CddbVbsuwr4YeRKxTTYSAH81YlARKEMECYnWQuROyjV4MdKOhYH
RyvfYhcYITX8NFJrn+kUYYnJKMXpEgukML/54+zPRcDx1wl8maVsLnWLlKnLPI8C
UAAUiQsx813EFWkue3zz4+pvTm7PKSWuiCALvtladEP/JG5akVHRots+o0C+AFhG
yYcd3XvwNSzThHYpTEodDNeZjS79YWw3suUZyhOB5h5ZjzjG6+7cW+1X69KytO/5
S51ZbAfWxWLx31bBS6K9dw6Yq1Dyp3I6Ien6vzjO3i8IMsVq4e+pq52R2sh/pnMw
yJKSYHNnYVkDJjEl7MAx+LKW5PwYIz0NIUnA4KzvwxJEOAeyL4ykTcQL48OTZES6
Tty4tNpueG2yVf/ungHWwy48w1fNIApiX17McmQCQRx9f+G+YHw38SJVXoFbUTrd
tIJ+TMZFbp0mHfNUWSapWlFUwQfyTHZgJTm0HJSoAjPy316eFC9yz48O5KDDMYS2
8fS3lpW9hKLcF9lEUNDlWa4vep0BpdQRWcUpU8kNY3WweFPEVxppcQCGAcK5J9Sx
V8N/75kjPX8HnxB7HzqYNE1PzBvb1X98lvxH243156GoOuAaeIuEjUBn7/70pLa1
Y/oL2nCEJaomPiKlTYXn/GfW/IwMbaecVhgBxnXRK5+zjZfmCwlIFrpLoOWyzu0d
QwOC1Uqi8PUqNN+ZmhmWYH2DxHVZOwvz9MOIX3cJWDIz9zSbpMnDSujEVk9jvTO/
C5BeswFZsoEhLOUFCEfTyG7cwTrmpej7R8UzKcrm79okn+HxokTD6FDqCqmiKop3
xi8h5xW+7deVu7arTxCGg2dghCYaqcHtqc+dm5rTOM2cmZY62DWlx0ZIMsgQ0dzF
MG2sMMIvUG1hPC1XcVqrSxgyBb45mv2Xi/j8GCZ0ebJX+kx4bmkNfU0aSurdy9si
ny5J56d1waiPT3FYDxaVyW8kf9xSV9HgYQraWeexc4iFmgHWB9dc9N0oX9S6SHch
LpcMKyuXM//8mD1TvCdUuWogfAy9pyIF8pb3oDWy7oVDhZySI7n1HvcbQriG3V2t
I0Wk3qP61PDT2RTPOaKOvw1cGpn2yv4q1HaY99bgnNFXrbURjIPdHze251T3g3c6
Ov2mTD5gOq0QdD0PUez3Hmqm6MaQYVuRoTwrDCyJ1tOCU6oFlrKaBMyTuJMupJ3E
SSG59entOXcxz6M6ktXv4ypFustnHezkRdIQPfIlhmn4WRD7IZLpKOhx0WZ7ATgN
UFhheijeNziUpY61fvNNTgJ3cPBm9hzTGWgzg9I0aEZS2FMzcSpgtXy9xhLleT/X
3D39Eyu6VLT69ET2sNeRqO1egaosRsNE6yoNJLhQxVFrzP5AkSwUK5AzT1C930jG
z+xvj+s7X6favJldE/aDlHzdyQy+YjjoIc60GbffDDJVsq7SZD6vVxk2sjBKY06+
ZzJ6kDpgaExVA7ILGhfDFDbVtS3Yw4WQFaVvgK2+XGBODuP3TJgorWaR1xbS5vL3
OLgsXvR74r48B3rP56xErj1kLlZ1oKhy+jqu+qIbgOnnXFkekKG1p2y2cIRyf06V
itx4quolAG46dZkEAR6ZGjYBG/IVyvOb8ar3wfB28kt1Sf50CmOWaCivAyt44rKe
/LJL73lA1hVU7JnLKDW9Oawd/OAgaXyWqcPQCQ9xtIa6LZJnJzXMmoqW9w69JSwS
rng0qbjAUNfFNfeIIX7pD/ExUvmXZbG8jInS/OqBEAFKNRcGk5N7jqLGdEu4RarO
XHNzkGTse5+EWZltwuM3DhAR6mBqSd4OPo7ixjk2+qs0tMUNWGtHI00QAB5mLTR+
c7oAGPJceFePgodIueG6TocVejlW17K4XKRq084rOzJYUeKuoQjqhwEDe3aaK9nO
DcP50Z7toZpobqsXrxFXt81pLF7coabmXk87e1v7o3LrE+LceJWGu3kYXA1lF7Mm
RiLpsLqWwMW2gE/Ra/aT1JKPseZvmntTRyViCL9ILyb+qHoqSkQroy55HZcM9Qfi
Soc86wJd1por1PSww/yH45X7YT36XOGvGgNp+6M3I2TBFIaWFH9c3cyHwvKnaeZz
VqaWUc76QM56Tr5lJnFKTQn11mU1bfhzR4AXgeNKjBZewNTTCzfz2+N7mqPCMVDS
DDh5IEV30CxZDZDfEtGtv2vn2GkYKIn2I/bIwCHTTkKydAiBBJFmOEebnLthj3eH
F5D1Ro/o2iyJvawqZcquC0dH5+Qp1J4TxiGqOcMrX/AI9PMWr7BVtgYTAxb24cvS
qzEyS0FK+8naN04hRcAEyUI9ej1g21GiKLirF1U8+TQjbCsCrRkMAybZhRrI1rfZ
sIyULcUqIIRmxfjPWIGHf6iBy+L7pgI8Lqngl5eU25gD0Jju6aJoNvMlDRUXd0m0
9e4YKJHBh1FNAQea34jw3ditPf4vHa5KxyNnBe/avLwBp3H+4RgGPLHPbdOC4SLk
n3HZlzGvbYIq80/dNHGrqZpeCApL8roG+thfUJVxHsba4oYSxEbFkRYAV7wwaePv
Q46NHwMIjzVkGThZ2Ozxxas8JOIpL2XdBgKZGX8tWUe67uiGpGB+U1egbA4PTH0a
AdhalsgtSy5uny/Pplv/ofrdUUzJNPU+ArY6egDNUXevsaEyqUvwasuzf9QwsqgE
/4AkOJYMH7/FT2h7GMoOoVLIaE5OV2SRIFOseEiZ6p9o+twQL4HSfGMB08EjCR3E
GfUnT6pAig0cpbhasFY8QwNxbV9Z6n/5BnJL4TTsRiShp6gZJ4spzs94Mhbktvf8
SiBDnaJBkhK6ssas+H2H+fwD3rDH3Kfku9wmx/xrDaqdT1Sdvef7UpK3TqtfKXNb
uO8wevJ5LokFK6bjLbw9XPxFN+g2RwDZ/RHYNOzreTb2vJK/POT+waH0qBuOfSOz
NS9oswaC1Hrlpayr7DlR7vGOfpnVFnvambdMNbbwFZsPVh5p05aWfYqBd3L652of
fwIJKpE0Qb96PHUAjfWn4fn54ijZ15rmU18bw0sYiqQ4mUBu58mbhDrcYXuXr0zd
aNjJM/Og9wDV3oQElLNhtQWmblU+WNqe7I2r9sZRhOqMnZ79O2cOVMBRqeXA9sHO
g6rngIrLibfLTd5xocAtHXiFKtFFSukO29NbGQWYWQjSRa+ylk4Wui7WnLHGmyg0
SwkQFYRZIBDgoeO49FRss+7KeOAloO31uASxF15MA7m/5It7YCVf/dqy8bcVlkYt
sLabjyK5y/0Noj93yFRIw7EfmZXHDEfJ1kb5pVoGnAici2N0dFldviiAsDsx8Jeq
oK5BrUCqbW2ZTFoACkR+20iUF8Vu5HML1AUzsTksGP5wd1iLAkkDkZ9JKz6zzyIN
MYHPJmCKrikwyiBmcFiGo6Fs+4m/NzoehOop+jcXBbJ5cRvoErtTYUY6BxBLtv1i
STAFVruETgZhiDI9Bwjvpzar3dEl4xESxnaSdvqnHUxKzkkoxUkO2IGro1/E08sE
UUSBINliNtCJR7ipzSM+BSs/SIk6jCPJTfyOFcBJMwgIUXOZH3s6aYbatcz+5iCx
vi9fFT9juf123fst75e1sbPfZ8sPeXFOQmYK/0QSLomdIVGt8JSLjLJkLjKpyxmX
VYMJp1+gXh7tk8agdTpSRJTZz1eUST7F0j1EssWoTx4oUzcQOWYMgINkg538XWsB
14YG1VwtK13/LzNz206Pvbb6F3+HdGUUWqW8JMMixdw5BbIPQmIq9cHa48OWyZJL
030WiwDdMIl0gkYauHgjzteSz7ciuH7Sse8j4yEfoccHpCt843VQC5WRMp+KQ+Zj
sOpSZp0blufDdUpJwQ8/8mCQV72TkQ/P27xFoR+r+rZQjDMBRGsLXb2AH+rt3ZaG
rOPGiljekcjgEvT1a2u0gWZjJmEzagTds/+zoCc0Z59sfkRoA+kdGAKR89Gj8MWB
wARLi6e/8IEuBnfWNTVj7r7zo2lCSghLTrza6P8TbI171DcF/MfsJXq771HopHXr
Thgi6DKjmoFT8kWLQl9V3AhWKzgwQqcmO+Fg1X9RI25BOKYZ8mXX2A1IDRYG6jIJ
3eNtkOhQvctVWbd/XZ+HP4YJJiH07b93LwmoSbVHRlnoXPfLGT5ggGEGGklrsOr4
lK4/Dstvbkk++xlPQwkm1QUsuJX4PiJrTHKn1caeN8cxcXQ8aJoiAs4XqmsP9/zu
X98SDQXCrF1sF9eoGeT1XzRhwB5kBU9E7feHz47zo+zFGZu9BYlqMgZxWJ1gjDoz
y+pnU5si2GJPz50C4OPYYpPGkKRDnmPpC/scvUkdBZOh9phZG7PYlY60+yQ+HCcP
KKSiCRe/wHOno11YJbkxe+S8+ch3Hm1+Y0mpTsI1HvRDAXxbVVFwEalpx4PqZMNC
7IJbfoRV3+PWVsQ5DmheKEMTrn4WJHId3iZf70S7okWW4vayXBNJxnKhBsl+nrBj
8XX7DHbBWt4FP0yOnCENJqfZdTv3Sd0lYxHlomFJ27KOMNuJsX8Q+zC7eGG9QCcl
s35IaTML0xIL6CibECL66VJEA9CgxKcfjGgdYgJKdKFmT6nOX0USuEIp9ch2Uxdh
lKMt7+/gklwWsc3OcxiyL/ybY5+wIh2n157w+IL49DmXjV5fE5MmKeqsTJen2xOA
sMF7ACc+1mHt2zUEPXjsRBntlPDsk5dd/DWLDFDwdWtM/qD5wHWvIEJBbSGFj154
zB9mwds/COLqfzW7lddVzxj/tHy9A5j/CRXN8+P9OJgpa/lpJDIG1sTMd/ltfNgd
StFQ2vrA0jblsBlEwY8KC8yuHYWVnjuazTkwxvclcOmCKD+l1s6Ris3XlVc9bRyJ
Wzu39zG779tHOZlG25xT+mhg/VTwgnHmq9ulGrdYpcZGo4bEvMzae9/5Ptfplr9S
/R4CTYw9ruTkiOwm9wHklx6pnmEmAo4ru2eip6cX6xtcgR3a6IQ0eVSrfPLKMqTo
46EEIa77Sb6/5Rnfp4psNlyq8IasW3Xao5ZAvky26Q2d2p/sqmq2hyhW3rnp0XBe
jM/Hso9Myo6zd4pnmlzqZjPg3PpfyoBM5jG7ZZ8se80cxDXCLX3hp7PcPpwXbvkr
azZ5519+/3MPOhhwe/FQw7bVjFP+UvSvQJPz0fqySYj6bvKoLJA8DXxBp2u1RZNo
d/bSN7o0EP2X1pLLShzc3W2gLcdI0I/VZWQa66R3q3nw8hZq12H62YXLzxdmSV+f
XiLVHjJQA98yJ/wq5FGOPamDncsqAcBTKq2cu3cD0Qxuef+YE0Fn82dz6KOcPlkp
Hl/yCltk4al5uH+Iysa7ZlLnX6VFYD0PY+iqe6PWFMTfbjT1W8svlvRvVzrdel0b
XuNxNCayTooLAZLmGlinY+BQUMwyP0gzd5qbW1J+6CXWoI+7ltXbXbFaKRb/c5+O
nhvaz4SnFadQo/LpWEnSqI4d1psFeGRpq9ygX2tTkjAsbz59eLPWxWLNXRnAH0Yk
agEmwV8SSO9zcKVQy9DI0yeC12HD5XbzCk7kvzM1f4xN1rB44y0BsEh/kkC3dG/n
PhhRXrEkjxvA6DjRwoosmQ4TpxIdwCc/7vAKGperz5E11ikG7PUMlg1u4N9Co5uD
eMzQZs+EaOfmMqBbd2OsmbctrTLaQZK40Hebf3rU3ocDGbarMct9upWsgwqwC3nF
sLq1f6R3Xwp3Hf4wDS6bgoeXyi8rMavA3vDTjm6ED+s+v3y0UUBsph0WYFd8z4fg
UMaX9hqdYHT3/6L4/OSCfZh05Bw/efQoXYGkrjwSTMDNNQi7t/ZGwP08Fcdb39MJ
tzT6X+ljnzDMuLkPcqlDhiWmV7IAzyfKJNeOXx1a4Dgahsha4HBbL88zYnoMzeJ8
I+Ul2SL2og0XXLmrf/aUbrCgBApNEBwnjMilnmo2xnr7/4g4DaPToxhR54Xukff7
NLbca1w/rTbNC/Gn8hYfhvuoxYzL8qCsnTMZk8eJG92RGHNJLVUfFHjHoSZJTsNa
AfVcIvipa46Lf+aMF0eeRWJkdbMebuQsG65NzrBw9a+ptsAdoGrC15k+nmh2Ekma
1JYumjJjbBwb0Mm0PhCJOfnmXMKBCXzqh5FcvL/SnrXK6EADLPrNgxXfCZESc7Fi
Z1h4pdLznoIWsjocI5vp4X5sBpeKteUQGMPTmcilUTW1tyj2LmFTgReWUUMIqUSI
ID1qXdhYbQqR+XBnC+M9cUfKtRY4PA/jxnBnNWeElEYQRo5FWpBHL1/8HqCr/AAY
KUBS7WCrcxa4i5jiV+JAy/2OPjVafnzcSsIBWoVwbdRl1vwg2jutjFCzdCNzThIh
9RXe44th0E6SmfKumTS8YnMWmdS5rU+Yrn6VUv3tG6VZZUdiZsPOj9A/FUMz1epY
9D8oKte+1C2AxOtcNYjpBl4WUCjY9PJL1SRW9m+ymAMHzXjNQbCwyI9I2aQx8Rz3
xRqJ4o0qd+XCcd/m9AkOOT8vhmacWJRyWL6Krsf1D1FY/xdu/8Jpi1tGKcuJhTwW
B0Uk0OZb3Sbk/csCEqA9D6giKcLRb7vwiheczjh2NAVnx2yr4m8sNfw2U/HrANb8
cbRob6kutLhcU/ybbVR3/zYoa3b/B9+Xu4IK8git1TRtgCkBPWP67XhFGax7ncsg
0lsCrkerHrFM8Vk5FG3py3Jby5MGy1YdrjyLh8X9385iZyCGk179Ry49xkHfq5Lg
dW3h9H9sCbPKbdFXUkbihdCbIoGYpZPs77UicXvCP8T7+DBZXBmupCbHDw2Ft0lx
0wpmrQ5BiXEoAsaXdbs1xsfwLNHGRVkpHWBirGO1KJH+B6QgyYR7PFBJ3d0SMFS7
1HrAXf321uPqRIo8QrXhLO5PeeytZ+P4cg6PgIjP3bRieEMmLHZKf2lvIWpswAgq
4gzhQlcn3yWFwN1LJcN5xNux5gYKgKILdKe+v4KPoU41pCqWdcTlLS8FvlXbHO8/
ugiAjwm8C8UHyFT4hmUxk7hmt1YhFGgxO1A6DUb7Ck0pnR6jj3CO+FIIaZWhEEve
2ajHrCSKZgIuzeCD37Okpy7fQVVC8HADdH4wJZBgI2t0cwcqRonkOeJm0Xp6/3G+
QzmtQCU5FXbASVu9astW/TbHrbKWFrUwM7fQPnr5Ip8qqkcRBN0tR1pDfCD6dotr
qyC6S/9d/mECnrNt00OYnUFMa+EQq196fqjL9hfP/QpyuJjHnGHfoauXdPn0m/B8
fVExU8tE/3LzTXtgcDPSLmpaHTaLUDaYw8Tv9ylhMNbHGr35ePaIhwXQqz7oj3PF
D2LohcJqkDxRIBR4sR3XaL1idecdZx1gHzYlNQAZoNU0DWR8KBmPTFO32irgo9Ek
0tJPt+0MUp9vD2V5NR1tE45bEknfFeR1B3N1NEIAYI3ReUNXzpkelSmLgJK/+jlp
BaWC0B77jVO1L7TCPOCjBTnuguAhFBNrQssGNyjeVVAcxOiqdILCIoYl2AZuSEzb
rDlHmZde70BJ/cFwwJ9LZawa3FeM+xAep1aaZsouNqlnVjtknRqGB0lgBAS8YEfh
DlLnu4+1BotQvFXFlVK4hPtkbR58VG1IpP4tX6FugiY4jxAQXCgb5BySDaMXirxI
7FdHyLZ4/icAOAf8eERMolsvHRp1sWkSmiIRssUfZvhg6RiYHNdJ0oS69F+XX8LR
C6O8KoLv91u3er8ax9L5aSkUzO+swyzuacJYUqtPj/Px1zi6zlKzp0c6Y+KPmNa4
kv+eXm2vHMpxdnQi9gZ8bqyovOyvl7HIYc+NyqXPIQin9xcMucHFaDnDCQkdPdz4
fX1CM29oL8vouT890/BOdyehkmUWSeoJcuk6rEED2WI+lUDRjWPOdItpFr7iA4z8
Wrz/sB9M3Ehfg82+ZKSSYiuLtcup8kh2owbdVn1TEudh81GXe50MiVIE10VQhEH7
re5YMqLbZJkKboPMP7iX5HpMAztGXZz/qNjxu0k7RyOnl1JO8xgPzEA4PzhqSKyj
jTAIPsRcf1GRU/cGF6DL/fkxkJUc/JqQOvoNY3h+yaAo0ROUNVxinrOH8CyGGkAU
QX7xJEyH+llBKHD61c/CB8/FkAjqaekBe/e50lXob8pc0NSFmdURcVUD7U6zbqxY
aloNlFoXAn6++D6VXAH1tJZUDK0ioQ6KouTBRir3YAL+eU2uIFeb2PGCC/6t50zC
FEwjOnGyixqSer6/rqtalqdRyjmxxOq7MuCcO3Ea9LNrE6R3vAQRqqrUvPQci1QK
CrwfpBF6/sfsBelb+GIrFQ+knG7hfnprkb5lcv1qz6MOhQbaR8ljO/3PnO9vvtYI
ETEEAEISThY6PV9IbUCIW7/uwsBLauajfb7YeClqPL19zYidggarbpj2Rd7i6X8A
7NnvyMqkVIC2iC5NDvfFFjCwkEkLxt1dnjrrQddVU99bwHgjQ07etpO+/+Zfm162
FW+qLr1eopfJxCL4v0clqEWB8El1nTGEoafIFQAnLauGrq9DtQOV6Sdkjmdj5Uv/
MGUVZG8e/EFOJUsCFPmSQgT7gk5az4LpGwZaXjWsDApn4dEINTKe69GvSck6ngnZ
6nzJhOZOK4e26/sLGyEKfRrIGJNuqWK3bHtO4fIy+oxaTq6FNjJn20k/b5hf3NR/
wYfp48HBMkORPQhsmrbTyKGSphg5E5mSQufD586/oQadsXj1OE5j1PgXdJM5xFLC
MAFNBJ8pn8rss5ouL94NqyOh6A9emh+2EOhdTAZhoXMa+sudNXeHwF6RkYFSpUbr
b1aWD22V1sgUzWd/NUvII/cBqtQcZkElDLbs00zCpmvdXMcNAUMvvYjAvfYSPiI3
DscH+0Zq8hplGkVV+TlcfXx+/GEkncKqd8B1iqJDOnk5JC6fdpG3I3ZZ7ky9u2cD
5vbiD13pC2Q+lmF50eJA4H5exzYZpgOz7R8Eeec74z7NlhDLgpS3GiXAsaGY3m2f
WphjV8H2Wv6IW/6wWCLs5vm+kymCVYXHXVV+BeKK4xVtzyP3oAfy61wGbx4Eydtm
AL+WicBOdbfVf3Fz5Y2jjWHroLzcTyYIZE2kOuSb2Pj6rq29JM/6cQuA5nCrUygc
9Ddxo1gK7TGnnYl/qR8pAFl37LKfJHwhubFNEri5bdYgECa8TwB+2QyCabKKZks5
7b10avE3EJcP+fBl59GMvNErH2rkx1/w3yrkPtr0KHDpqJ8p8TZBrDZXXsC1khbo
7Ys3aAFK8ICBgja2yD2AHFJkkpN7ULWX6RdMuiP4KarMkdavKr2bWpwh9ia5VnC7
JFoqqjUpR14wtMrLNJmb4N9KUgfkD+B+xvEsvFK8HK1ohuDqWRgWzZvS0eGNmNxL
QgV4rbcjOoKJryaUwfeF9IAl1w6uc8Hx46YxrmU+jCc2pQz/IPbOMf1gNRN+zsxy
fziyq1dUztwBhbkh/oeHC5pSpZ1Yrbde0gQfIOWDMIuXAL9M17uzMwUUdZGfLYlb
dq8Zc025hMvUP6K4oKhwlQdCwUc6xpiVapqqqfUH5mZ0K84kYxct3VKxWdiRbp38
MrBTXfaId3pu0KyVwfPbK5Z60jYOJWJzue5qSfgHqGQjIL/6EW9aDI99i6KzB0Xs
/7K/qohK5KvvvuFeFth8PHmL0cZs7VXXbj9B0zqzFgXHR62Ee0PW211wEb60Cv/4
x/JTwpob/3KveN7OmCZ7giJI49qct1nepixDJP5LijnRtaoztcIDBOmjZyyBYT1I
uBAhjCCsGviQETb3PRaSjrARCPKbtYovG2DYWxT5XTi4ht9383PiT446bk6UViNh
ePwxAbxk2Ms44LletGmV4XGphniGx7dKK8h9nGht00hqSRjX94GFbhxL2zXudH5j
LEz6G/TfdmPbpDzsul35fEou2hBeT39tZeWfMx2os24QNjDLMCGx7ucAXVvXVtU1
QI0sdFTOl2aS8607AfNxY88op45jbOuDn8x7F1Huf4Tu/yb44kSAZun7I0HZU0Xb
3xbxeG+tTqFofmLJ/2yammejOwQ1QegG2d1X4zOEJWPcxLvXqcdP32r7kg8kv3sY
Ll1mmH7O9VYsViTTNdAHzNK1K8K+WOz3fDtNccUZd2RlN4NKbnsVs7377FnJiCcu
ykZTBkXazFLC64L/49dys2XiCoO95X6O/tsbpB7UlN43xqE75/583hmaJjOrveyx
XI3wMgVtXRJQsZJ9c4xEC+AA2Ga2vYrtVnfQC/uDQMB9UK5AI0VyBFFkghpSRSZJ
+YjiJL3R31pVhqahAZbS3NjSBiZGPyLkC6ETjDa0CorwqZAwyifhsrR87Tlo3LLQ
X2dIUCXnv4AjW3NlkJBRbhiKhYiJZ//a6DekM4LKPVRZGkpOw7soFPkKEIlBWqrZ
Ucdrv4NrDuBvv3T/ohQFpCOvITbyzh0yDZVqEbbCrFy9BsbKiOPrKttNkwJ19Rwm
GyCVXobrdPRzREHh90vBcaCk6yhYJbDJSPC7BlbyU5OdpXG0kk/lWzw6rSGad2Z3
m/rYRFVvmjIklbPIQmPlq/vZ6q8kvMLxeAd/W6NBcGvO2wuCQO6jd7+cIiTfsx+W
vHyeFffGHuHzlXHr9BrCOVYEXhN6rehdqOJl/Y2h+uf6ieuFBJWSy0JXXnIQkoli
wkZo9yjUClMlXc7qGXW/XE1wbRvyWT3gScTpX2MlkhDpq/9whcUgGcA1q2EV5k84
wU/q4MJWSvATFZL55mIHVqGvK28J97J7HxWgJpW9iNjH/M21p42Os0LGUcpOGiPW
ZKa1DOVIZBjLEnVGzAdQEcLCw8o8c6u7pUapko/HhFrtWxkrh009786t1bJGfC6z
Kv99QA67Q99I0fNQas3vxREvV/+w3oHA/QgZ4akhpUgpZ22qfSur6RXlOoknaXYg
YrKgTxZ6/85w7lnkFr0vVrsr/queajTCK9eqINnsrIE/VED5xWllcQuHh2UGTQ4F
8Emc8Gu4FldqP6gqzw6wQlEPLtWiJSuS3PSGiCJA2T/NnGj4AurgBoL1deBQqVEZ
Ev8OR0nKycBQtskc01QFTxKkm9Bp9HgbctvkxfmC/XH0gmjoRTFTqrA03A7he/bk
fQvg/cqLAOP7m5CnS/Mw5pxDEdDtHPfcx42ondFUde3YoTYtKRaqPE0CmCx71vq4
92pBnLSTEcHWJGoBUpLRFs9pBDXdmhXCtpUSxKELCnCfF+P9kE8fEekMZHyvvdKa
ZxGJ+D5LUgWYGssVUsKzY9ZiC3bhYwjPtdEFfZrcgrlf/F/blir3CSxv7iOnnfxo
WtchqfCj96DdftLJfXUHSluT9jABLjjZCvmAW8JDRFZu1QSl82v4MCahJHJmuTxL
2sQyWeGjcGQtS4SrtV4LSPNKvMl86Rn07yd1UuuushsfEhNvLEX8nLZ+pGarcgmr
lSHN1XVc9bBm7SYgKrY0kF38zdiSDYOTelVQExcg+MMioPsfoX0pO4NfIqgvYHjR
rSBiBrRuvnvMZwpDpzD6h1Pbv26zZFyIAk7XkyStk9Icez7PiGtO3B41g1I7HLhy
I5mJyc0I7E7JefFiyFdB2+zqUjgfe7gFq/1hTPTtbqYOHKIgGnmrms7innHi7fMe
acYKp8o8P84P0uSwCejeCc8VhiOJ63GaOMhKmFWy6Vs5NtyXRCHUes9p1nWtOOBB
RyAdz/wGjzzrFkPj1v23AfqXsWowKcZV+yjx58E9pAErwCIAwEkRijQSakpkuuPd
GXCPY7tck+CGXMrkHD2xjSG7Xbf/91GOAg4RAexb58auwm0gI2jBYzZOrthe2fsL
YRyY34+MelFpLLsZQveAKDNQdlxXWKwpbxa2bd7R7jrRW+D0lASEdlER+KKDo6UF
TUjQgAUl7F/jEYHMiaJmxd5GzjRF9o8AaW0PoTNrXoTPezpuUnk1MP07z9W1djA9
BoSuH/+dlt/4ToI2u7K21IUDGbiSq9/DWWP/GJsme/Z49zOcAd8CAD6wosWubvjF
9tAQHHenK5Ux9n8ICQVVPjYQgjglgp6yVymPaf0ivKYCTZZ9k6oY4aujScJj+KHm
e63/wxoSe/79Wijf+vNgFa5Ye7QCQyAg29wBwhiIn9dg5rl09TRfhS44ZuWrrsYW
CRi6InZG1V2fhrZet5zmz6jyhCUmMvyCXLgjuJhGfQQkzTwOm0DBFCCPLJ/0fCSB
2i4wa+OnctIa+76Z1jjFw87BM0DTfHtDmiIAm4ZDH7igXD/YkRvdymX5PP5HWclj
fw1HzrwA3FejyqriZ5d1rOKoekMWjJinWZzVttuBZUIUbsFcwf9x+PJbuKl/bvmJ
Y3tLYSxqnnSdQfpm3TmeYmjnQm++xJ/l40sns6ooLdlcIKVLE/zgtNFwvIcvLEZB
gGod4+jiBKKZ4QErslVIrXOIgkJNYG+xfyGl0Y3HQJ9URpjUdvcdq4Vy8s265NOu
LtZOOLZz4Bd0BT4+eg3YRWO7XGCBHYY6H+lK9EdEC7oAgR8ixrQBhfTD408GTbmI
Epln5xpiAqoqWrOTmBpEmeU/v8+nRQ4p1vnGqnKdC3dYWf+TmnfiAKrw/m++9vDv
Ff8IHgkdYoI592XpTM96mTauI2Y0dbgisao4j//2fLGzXIB9Y2E2QsAshmMn3Vr+
VCxj+Ame77I4j26YRk1UzreJDm+7/RxORA/SdhC4Z2BfcJPzc6K4/bOm6Fl92FQu
3kYLykm8HLgkmWz0iXknkPrgpofMzIoHt+r5UJmOnX3R0N9+KvKwW2I23vTEPpUg
8hJFyTbFUwJKrvYr2EkK1F5FuhoPEUBrya8uQeMRGZ30GD8XEiVkJIobzzHv+BLy
kMyLvxgD0BUyz+dadGOUC0iqKvnfRgpTXzeuBMKOlQuCh9JJCeHAwWrMENy6DZXZ
G+6d22i1QCSTWJrxa8BmYSI7XxmqSY5cnc0zd+64F++wMdzgi8RwdLRkrULCZbfK
jfSBg+vZDhmGuIr4TIfC2Mtfla66anyWr38PwC/9Sasx2hA2wpUGXTl4ML8zGf+n
+wHfpJX9PslWlvIiQhSHHaq42RfLFXouv8wJdpbiY+h7hHvSo0HE+ZN2op5q3L1k
GMT5nb5Nuu2HkOOu50pgo8SNTERmdscW7RhOQgrQs/P12bEn0mKiN83BDxmZfGri
DuprAPOr386HxWxVw1bJ1nrTyH9FLFV67QcIczOly2qYQJ1llBbOKnyRlHrfNxDA
hij1mAHeFbRozY+j670dMV/sRuLhSMWUCVeSz5nJ1nuaaQPEn9Jvpwzi9KY9Y1yT
skTVN//2CovY4usVCqwSqsvs0WWCG3OtNw/CGpvu+DM8Oizia2KVD1maeIihH38N
WMpu0lldSpnAVvQG5lguajwdtxDvLEJ/s33LpgSQT0Cn/0rbuKm+P9/kz4u3a5qZ
XILSMvQpty8+Rwx903xHXDigNrVs+q9kP9+98OGWXejZU9hf7sxmYXrUKYBJfm8n
jk1W87VC8mBFyv6vIQlp6Gn2EEFGjK1ZkauGz+glm8EbBwdr++ALwWcLBN4pXjLW
nWrC6u2Exu1pAK917gTZUdYahNmb4nkwqYGFpWpDvcH7iODNCYvQ7OiBUupQRmNg
o5zrqBOf0Choqbc4RMBTTxwAMTH7MncwlBTjtOdxsXZRpOZW3XCs2uvh972I4Ltt
Hy4FpR+K1lbMd5SRt/RRqARxG98osUCdS3eb6SelAXVfiRPUjQ16nde/zMwJB5+M
A3bmyTOaUORR2Uc2+dVA/nmaZDoZl4+V+6nTr+VPDKdoP2jsrlQ6AaPtvgji4tF1
RYD8EykYIMVgC1uTCkMvVn9udZJZYFsz5TgHQTk0abPTcD9Ak2Zqnt3PSc6D3leB
0kva/hitIMntXNiH5Q8OvvV/nEh0NaxkYe3JxCATP7TmtgW3B3ftPYlJYkBdH2pE
UVtiD++SnWJZXCc5fvZoAjlOMmy6U9y9h9mHNDjB7yKZxNNCBQG9dhuNaaYxZuWi
JB2aN5kQuu5Jl8/jWnxG8RXLpq3v3X4dsNdhhunw96wLcoUA6pwMYX1W7oLjEHT+
teCo4aBlRL3AmMvfSJ1h6ocTf/QJPBelc6YVEj0/PCeg3Hl2fIawi19B+hMo0PKa
HUyopO2Tv14mdH7U97qiTYMb38ky2QaN+phgzVgarCwb1Z2nddixZOSlsu6+hpTG
sN1gHdFjNJyh+RNVsVeHEtM1mopK0QMZ3VEcbFpFNSz62vWxIdKdMKBNKDVoBACn
8LFLODPWpVqGXYVQyLN2ws15kTu0d3HVbZNN24tVfYtUpkvExMoma/XKmLxhZCD0
vnu+ThTXWVCGZz5ETptvnC95SAz6jhajO2Dqy2Q+mcOLD9srQHN4pcrUbYaT+Bc9
9kzlBR7lzVQoONUgiH9/ScWMB1FEPhHB58CMgdBwqE9USmXD+EQOppjjOiPvtXl4
2Ft6fRlDCaAutqHnHkencR73iNUUUxZxcnPdDw9wAtAKPhmHnUVD/g5MaRWu7HCR
4KlnNQR6gHqehCN5HT9D1u12WqeBRapxCSBPuBv4INaIkItv8Mi3s94R45BGjyDY
kNoQ9Qj+F9E+wEnVmt4REH3PhpgKJ0lNTJjdaLiq8n5/uxCGI1gXbumns/YfeAW3
lS8X4SI2ny1NGsl1gGJY5Q5ckuBJVLid5sH9IFcP6ZkAeK0Q3qU/ZMQna7364Op2
wqXdsLRI1FLpFHiWxaUeO46BjBguKgihEZnVGdbkyunbLZ9T7nf+mhl0rw94auJ2
pcm9K44Qjwv43NB+bm+dM4cEBY/XVDfjTOdWUKGo7NwpvSpbadjFm26sre7KXw4j
8ontsaH8c5IiXlq2qXFm3dJzlUz0w58RoQixnS6MURrxfVTiapNYHATJuT5XrVAx
uaqbVFvEcpiTP6NXmWhjKO453tH3Iofq92XJtD1WCgZVPEJU8HnXo07EmX8ut1pX
Ed7yIarOhe5+mSXZAI8I+oW27sGRAuM6Sx3ca+YhnIssNR1iUkooJQe09UtnQO4U
xFE5gnVqJYM0OqYCLVvTXfo/72NAoOvVCsE0eKomjimzPS4pzZSrD2/Ytn7rB+E5
C7D4O76fAOVKhZ4j5gG8WgIHy45L05ZTxZ8tHaoYqRx8sRkCi9CG5he/iGuOB0fY
XbyaMfVHD2BUkOG2VqseDC41xZLXs1F/WCUVtRhOL+wW+HarBa12pNOPCsj2K71R
2EqsLLiFnUEr7GfUeoe90bGiUM294+Y259Myb/Hzge7cjfclKufBan7c7YGO1QQX
Yg4CXSxaPHoDyh1rJY2C8iVNlJCeDK76fgvatn87/Oj6MRMyoEQMJ9ltBFQa5a+3
nvYMveuaXbobWFATEme1VxdXlFUv6tsDw4Je9mpxZ8PELIBoVX1bIrS5R3/Vh5Yy
OfXF0b+qFboFrW1k8ExVAMVoYuqh1GY20LkrqJ0OUG8HL5apI6qfKC8ePQ+qBt89
6bHSREciDsIcewV5BLv479CwlVoyiphYDI5W96AtRFb4lXXcJ6LpaDslJK74Trs/
MV7dpKbZgs5kRnDUNC+0GBNKhtRYKxg/QqFhiFOnUDLdtqYFRY0z8frg5K5NpF2D
hLBpdr9jWJYcxdh1rHQopr15WaUBX0Coq/NwbOvUvj+tBi+OgjnMbO3iul7W1Ye2
R9UQSaw66E6MQcxuOB6/mNiP8iLTLzj9vUP14Cjdlu6ZKkICEQNNhjM8wBUPEcav
42cAAOu3fPlCHsq0WY4bZCXc1ZcAlradn04eaWJR/gh3/KNXAJbedAOSnCX5oPlN
cEnXsrLvuuDNjHztZ3t/eDSUk3N/nfV+jQgALTgUqJF4l+WlUSlUeJ05MLw7PxAA
kO6Pe06vZ8jiuy4bRVMEESTkT46//gYfOnIte37BYxz6Dx2rPZieOs7DFP8JK6YA
QlVBrbVO2KPGmUEBylwWj9QzA/HDUCPo3UygSq09NPCt4GVSsMzHz9EIKJYe8ou1
Y+RLZ9XUjyOqoTmjAyj5Anx+ljDcPadIqLvqFCS1h+i51KizNed2aufzqo18CfFo
t89MKhL0dDqwYNr9acMCNxjbx2tdmx4QYZsjq/qECC2SFtRtSROOspataL/wwkQB
RbmGH7tKPVEgp6+8NroxPgV/aj5Gi+HBdH/6BzZUOnZ92U6qZCPequcaCG+qPBSw
L/doCq6/WSA26/nqe7la558OgaH/iO9MCOVjJMZIqlieqH1YPw1I6UfGMj9GZA2M
eWzKl08SrvNJotGQsKe+DNf4wNWNm+c0+otec4WLzKqJ3sVlhE86mX+yyuE2g+FB
NE8dk8PyEOh9ay0MNrzqBUV/wkpokLyu3TrU27ZnEBTMJC9KHr1MMfp2eeNAirUg
ImCxJfUPuEia6HAjcr9nBDEQBj8NAxQKAKWYpf+JwsqNmNeFz5oqW5priIGwXU3U
ykCmPJCKGJ4tUm2cM/IseaveOK6KcuAlkw7taMJgWHtniNYJU1NnvsxusQZf/EyB
SWFHUo5nTax3R4U03wpvq5sFnRxYPuROy3i+fvf5KF98lJCWpr6VxP6q+y9Nk1X/
B/f/i4uuv+Jb2ydAtx+Aq/up4p9PuF6sAd9pOnDje2zup1tYBsvSVE09Udsocx+V
plvqZaXFBiSrgyHyI6ZFTsXabVa4kLMOaamNbot3RWvmJAaLJ/EapReM0IMvVS7O
AMVAoxCvq6w298TyULeXlL4sA4c6ZGweUdj6fKqvCApRvwSeIjqMZ9JWjfMSuwX4
0mrQYNPHeIhtfQVosEopkIyxz+XoWutFND9EmndJCLfec9o19YtLy0rK9hg2QK9b
1amhEb0dBLXPx7LGc6dtywvR/zPXVRFNZqW2h9OKyvsM1PUj8N2zyGXuoO+XjQAo
zGwnTf310SdL8BjlczLKpM+9vGtFhqby2aJkp0hcIWqxwB4coUTusTcQVeqsbHx0
ux4YCaP9MvI9tCInW5hiN4tGvN3EwxEC8+mJGReMsMQjFXeIdNzzKemwmaPjEkfT
cNF9Bvg7BWW9vovQ+awfx077tywAHjI2XzO+W/ikvP4roV5oS6D30tMpndvDkPGg
J0RZ6hB7x2yuEOLNK8HBesCrME0yhUnUUuFGw1XFWK2LjpV5/bbSABCSiiTX+x6i
gSllxbz2cpjV16+GyzKovMdU3jJgkYBeBR9sxXVT+qPLUzyzcw2fdeJsBzzKH+3b
HqiqqIgt5bpt2qasJpwtlFRIOvL6K9aW24tJpNF6/8b5zmkIsN4erVzKAQhAQS8p
nFwITnpdcwBL1+FWTl/YWZJCkbRZ+w3O1qqa7cB4/3wUXCZOjSMlgmDXxAVMNEqF
LMN/fgoA5JZlBL05SRQlcSAfULq+ZlL7UdJdOI9TEbT7+spHFFWcw4Rd2EQDSbn0
o98rRmPA8h5to6EFF78fZSUrB7I1mmTpJA9Ft+iyyY5hqgiS3GgyHdVpIux0ffgB
vzNdvctlV28RNSBKlnNdpXGJzs7S9bDBrz310AdURG98IXIKkYAT9ki/jh5KYfrI
8D7QSmmeV+5zM9dtO/xY7NVaQFrOLosc4UfkwuTw62BWsTlfa15xSqbFxCyD3cp0
OuReRyOUe8Hwvv4s6n/0uAY48Hpug4aP+IPVaK1RVB84gnsHBLj3UDUMx+9rNM/6
DhOonVq8pQopAv9YM5Bw6mSJlPt2eaztHqxrxnyayVZ275Xhg38C7p7TktgJjcfp
mcq19MGaq9lAImr12rxtzHE/EF1tSCHpOtfKqU1tahtXd4KOBLILdPThmzY7EmB1
Rs4M9cfv3+1HanGK8POAMD7jixScHMxHlGXAj5nUFXb20s5YoFjdaSvGFWDCKTD4
aRt/NiDYrhxjuy9A0UoTdSA91JRj2+eh+k+fP67FaXJkEXMpyjTePLoRHhTZkMRo
ofpb8I0BMgSQCblPDPaaS6jw7dkvdRyyYsYV3mGH+CzYLJOpOBHrVe4h70vNYoO9
zCQTv29KuJUp2WQjzCmndHzEFpxG9/LLsLKJlLo18kaDqUxH1Df4sWXX53IttP06
tS8jBbYOX54GEr5Mx64in4hV7bky5o93QBTeSaQaqZwWFQ802F2Hg280MrzrdH74
EYKRNi0niMNkULWd9/qN9At7V1vnPHZLAav6Tcr2g5N13hxPrfnHJsu8Vz1Y75Vz
vMaa8vaRNkstcFjJfn/3wjDNCxxnBg/8qabefu4VKs+vv6Kr9LSrZ+/QGdSFSqrl
/kAi3REnx+CVLIazJ24IyfiT4ApkJ2jBlaWg/ZOlCXQSL2dIdej/+y4SMiAXdIBx
/VbJ5bD54QUsfar7dqNvR1+aSzk6LWRUR5lKqy8Lw4WXnTgJV/A95ZzL4UG9mYcS
wD88hSccvvAdmW+5hXtldKg+cgD7g93TqQCrkVfebDChlwssCp5dYsFxwzFZrMvV
Tp4szACKKS3/aSzp+8hU4t+KeDnJsRwqy3w3tGhPDt5+/px60go9x/pF0hKReviK
e4XuogsPFWs2JtvP+7lAuDEs4GefuPH7KiVNTy5O1pMW+sxIaXkM2E8A6zOI8CDo
BRMuTPjzbxm0QTnmOXYdTnyaEPHjRoEC+A5Co/Jg6SlPqyOQiOf15zj9QAqqpXEP
93jpQjYu0ih+AOR1ty99BZMOE81teGFeExS/3cTkcOWiton6ici+4RcL3cGqmfLb
CZc/LXO5Vmqkr/REWmzipS1C0n64U2SzFAZINQOXaGp6zrc/akoCsK1eHJvVV5Ti
7M4czs14dhDkKOi1GOxk/ir60cA6f7QRDs5mwr6+Ml7zYr/jPL00S15uGkwq3wbD
SQiz+iDIWt82wri5j6zQnHT734/h22NzggSg9C/hwTPza2s7Rc19kccUUfKZM/GS
lQnxJ6N0V5gxKBHwMyJayE2Iv2SN1l0M9t0QgwCsjokhCMypDv0y5zTDme+yHV/6
4skUZeHYVg1eTWx2+N3l+NwbSuPxTImBQBzcJtTOw5eyZmTx6sbh8BuHhiFfokp1
MV/1p+wlfrRGvAFrEMXnh3BvxxXdTtOY0i6Qef0wMt98l7oMHDZEaR8fTP0wQ0O/
V1zwOWAsyk4dcFOPEx/uzej3voFNiwAqO3ZcsSxfpzwTrNXEkIPLG75duA0LlDlb
/pxaLAP/e2Qa3VVevEINteiTEuMn2QKq3obgIFmaB/Vils+nAWrm//OMhVDON8bI
Paekz7FQ/LQ6OuNVwFB/d3382xY8p3M5OHzTjFpgqq666nA06bFKn7CAmADz9Nxt
7lCgryDLZKCpdwT4hkR3Esc8xxELjYY+cOlNQ/xUvJhw8RfDwciLyMTNEZ3p+Bsz
CrtFK6JfRftynDQQCPUeF0dvq+fUHMWn736i/jk7ay69V0tfSQxvU16VxHNOvlCu
ARNW2c4ElMsUTA1QO4kwcUIhzuJELleJd2G++8oXYUHxpZrFUX40bPGw6gWJjTgm
cKjOenb9wff4/ksTHLuK/kfJhgvqHHcQNe70g/lIp2IO8JUryXfq0os8ValyvZcd
oetEyTLLet7oNlWTbFdz1g5bM4KwFnu/tmKdGRF1D45fPVvFOFzEQCoZY2MJpU+s
ciJxC16hqmWqyYl+IpfMC/yWzeIT3Ct6osC52G/gwLOSWx84jxH0l/1TVLRjFI5r
BpwAc1G5J50BLf7egOLekM/MiYV9ydlEMjYvVLdgBS/xhGlc1BVYhM9t3ndP4tKL
zBslFuEaiwhy/wCaC0UltPJXXu4f+4PMMdYWw2PRIc6uu1FA3txBRvSAS0hUuBmz
4c+Rr623B3Yv98O6R8+bWbTWdPkbCjVSNtSHjqHVenB+eP8k9WL0rixp8lHnX4g3
b5Zq8nxFAUTxS3ivBfB8bkw7YV7PVTy7cLQqhOH/KZvRXE+TK6NV/Qed5JQI/xey
tS6McQKkYRDuP9QWp+0Ri6lFOuSTALg1xd+Jb/Ramc5V59EYpknKboCk/cc6DS+8
vEcip3woupKJ2ExkIqqTe7iodAG6l2fbcwehwtLz7MZ9E+v4gzvFffcKol7HVyeh
hu0njBRVjWUYFA+WlZpn7bRi7P2SVXx5ob64SY6W4lapx3PT0WQnQVGcU1jH99NI
Bwf8ldSAd6ozVIDxSuWpy8sWEEd28zUytoZf930HAPQUyQBcnwxTNil7BpjFztL0
Cw5aAirW/YdNuVyAx8MCsQ5TNu2I3ThViRjuPWb/uxASLdqawgJAJJlvas1Mmad+
kB4vTQLmXyvsuaExX9JUR7zlD1W7v+uw1P0Xf2Ju2CdMwEI1yXLBR4hDGmIwdlvh
ZY0T+MmePnCSSQBft3db739bKAg06Bu6g4Rske40KZzt787od9trGw/C5bQ/pSVx
qI7IHdm232F3l2hSjAmzifDj93/pydkGm9oTMyAB7qNy92uN2eYy8dXaNJ9qB8XJ
6gM+B+p6EX24bdaf1i1aiuOGhPyCnjc5TfdZSEBbFqvN+6fil1h4HVrswVkxxXJB
4GZxorVy04W4kkt8LdHgw25U3U93mIND11auBeK+B8vTNLa49YGchuXohpBwbQy7
R/DUbPI1gdLshWjh0pNfZS4I/rYwB+Y4BoOE10up/lbZ5UCBm5bJ5b3H4lke4fyu
+MYjhYpiovi0+sHGXJgJjGpVxsPWefFCdzTI/OJLH8EUZNjWW7TdR8/KuCDQq897
2TfwmBi4caJFTUKldqFlDEYvj0FyOGHG2I5T6D3QWv+eXsvNG56qdvVA8Q6zPlzm
DrSjQBAHb03cwjheMDAefuO1h/r3MuLaY7h+Tl7ytVJGEkIfx2GysRjpl51b9orG
tuMtlVhVEHieUtG/voPUcMADTrYRC5Jjbi/vKmOonwvPe34u8buqQ0Wium99WkSC
x2UAIuqT4ljPQCGrvyXMPeY7E9/vyjKj8KoQ25ucWt6i1GHnLAiTP9dcZ6rf67sF
WGhrVqUAzC3m2tg8OEXWeH3Sy4yMiLv7wiFmMHBErQYz988381jeVy0FW5Fsq0bL
Zn3T2vzfqggscTH1MZ5q8G4pVzfpUk3Li3IlS/s2iUUzXWiITFuL4IfaEhFDialf
eq/EcPrlm0VZwFODGJnPIrYEhBNznDUmpe1TwRvrWxKZ8wCWIxNL3mkyjxtJzjjg
OHo1lalZyNfOPrJ/IoD1PuBok0jwymunl4cBmLTaVilApiaeu8geOSvSPRAN92VW
Lsec9fzAOuuFqStwSy8CgALIQtFXAdhn3pWuIwhn5P/T3xxucWR6oTuNmVjupsnl
mBONxYWVS2JRJ4KKZzv5rJa7TGUQL49aOzPgAefjY2ZMcWjeqYdse9nOBNLEDd3+
9QwLVVQPy0tpQtoZorzfwjDpnw8cG/SAUmyzPX3SJEBpLphH+BSmxplL/KVJum9n
lCMOYtgt2h4PWlIsjUGoWugYRt+fYpNSU3U6IwTvk5+F/gO9Fk7zcNWpQ9TuVYG6
GeqoXNGjRG1lpTwwAnIMZsijpH5sOJHR81+L/ekhW12UIpwi3tvSJpnsGW6qo4+W
tvp8js95Y08v3g8QX/IryNE3mayhPJrcT25Rn//4PZb1wDb/wr+SqFVuGCIx1VBq
huzYWOkHLHY8o2wiq2NhbMRZhByl/B5cXm7B1YeIjAe9gYS3YlVDIK/kkr8f8tDf
HVgI4dSOyL5gvOrHrLgeoJ6ALfqGe0ZN8BlPjgDpFZW9icxW9bda0oygB7WW5Zeo
eD72yTzNUMyjrUUzruVt4twG+epJCF/TmGNCtXb1W3fHJ/5VjqxCmjsM/jZ2k5G1
q679GUFC6Sgm/QdUltabdnMVH4WBCFPZzDhwrSv8VxGT0MMSsOnewpTJm3zS+DYS
H6J0H5PC23ebDHk2arRkssUout0et/N+om0rX4P02rTqtZYL+63Q48RM8jIasbK7
xJUo0k7NY1eegYh+rN8ln9XVs5OzjLWPomG+5sEwgcAe6wSXtUb6zx5lLYm1S0op
/mfxt+COhMGUCpHnIonOGJHKdtdDB4J0qzvlpUXOY407SReEZvpksQ4kOBMmRdGH
nq+jxSuC74w6mkPbJOk/qcehH/UdxAUO+fXKmroeKQPggyIImbqBVAtD/f2DndLu
6dCimIP4d6MjTdaDej9gg2irEfwpzzpbTs1n/BJqf0+l/4Shn2S2lUTF7GeaOsU2
J4PZJmR9ioWdQgmAsbWaesBZxhtR+lmB6X3a2wdA1CZeTnrn7rM7chv2swOK5Qub
1/uySEXKVKtL+pgZDOBxmtWmLc7uLvxqoJe0LjRqoBsKyeq1ZiExYonlMEfLfsnj
RWWiSR0c6gxXAi38KTgF0uMURiareZIM92s354Np9GbYjcGftqTo56VoTjxEh3j3
kuH776MQd31gvXgAHX+r+hKzEMKN0DCym7yuj+bKjKwUclV5qhIoQrhD5SPZ2MWA
IryESwXBXtMGGDzBVvTiyrS3pQV61M0bDf/yD9oFd0LPKRWjplU0LfTH4dOols7S
zItKvL05yGIgVent5nZ4rnHFoR1nGBWPLRaRWm/0vWJ5tvBKfTRFw9369Ka6Z8pg
HSh8YFmesqGF0FgGSaO61UsAgfhVc/c4Q+70RxjystGJljVBZy9wgT40yEe9UqfJ
63kba7LeQSHLvf0yDW0TWjLxknVDJeOXeBEgUzdMTs9EYYrb1WfgA47aoHefh+IU
t4MUOG8ZrE9wZNz4Sn+DIiXDf1WVW0kma7Ge3XPIg0iggToe5QnrZr+/QiWin5gT
GF0b+wi3kbcO6VSOHDw9ht9x8F3dyDt+uiS6vdcPzUFyGmY7/gdyyBR9wXxJF7LA
N4AEtna5JXB/TCnNcKhbNhp5Eb/kfaMnZYI/rxK2u/7fuTc6RUyP93szJFvPAoO7
S/QPztmAuIaj7OnOpM6AFIB0oiptpTHA2DenMIGSczfRwTLLNDDVxMDbi6918+Ke
7uDBQcFNWjA+XquhATd58KAr2TNUyejBrE8bfXJzteb0+QtxJ7XgclmWGxFZqJhQ
0iB11OJfHjoFroU1Z0JNRHuI85yQR2L7hkk4BM+TyEk+Wrxq/qjZtbB5PzQB5e25
RibY8vrnau9kHnv3YziWp9w90nIld9xA1mWIF2VLgfOYA1zgIECqRlAEz/mTkWzI
LHkdCvpLceMtJ/Yi9H4XkcWTofvMtmnfSihaJGxDrv0OBzm7XN+vubeLfFy+XN7f
PbFYQGZlVMGMa4seUfbxuFvJaU7wdgNseNK+rgq0xO4ZFG/Wm/ws1vJyOLqDjldw
1+aFezTCK+rDgLCLkc8hVJTYpk/Y2JrxZ0ylg0SRUCpSYnsOB3VrGFwWc6LUHhUa
ri+PgTOwtRjRk9z/vBGhqRYDn9thpzJ1HQLGz1r7vUKZw/e75Af84WJfZmPz4wy7
7rUFDqTOt4x8hPNUm2rQSGZewJlXOYtFTg4L1q3qPi4sqLp7tyoFznNXEIWS54Iv
cmisuTFwC9qdHRPzumA3o/ezA4j4g0rnrh7G2HJEGyuVhLoug1CyuL/xJ+CUxi7y
PKQOeq+IFCbJ8ipCVHEoIvlfB9gEmabXKg5QLvam5MMHPhBuHU7Qx8wgu/BqZbNn
q1uEVFQUfBxy96IxmZG8jc/tD3cb+3EY+WnbZdxi4L74eSlyI/8a7jLmiHpUyRuo
AiPh4GNwyIllwrtvwKTCi81CJsDQPj83CW/UqxMT6nLqnqYQLFIvhM5Fho9Slwg7
UD/c/ZP7cp4wSF3piBDleRlpgtzwrHk2OxGv9AxSqi8ZDzNlQQJrEgu9s/6Zb8OF
LwWTXrTVLluJi34VYFonvnhJZBpuTBgGMloz57X3K7CWi9KNkaN4LR7FGcasB2HT
O8yaZRVWHfwESD/3FpR2yO8HQGP5rZWjCcaWOHQuBDRrEIyTH8wtTfqA4X5yrVBQ
irexvZgx+gcxwe3HuGHOHKikZ5RNSl2gnG5av3OjHSPM0zL5S/QeCt2j2nSkFC0s
ys7FhzunAQafORyc5ywXU4j9Ktx7tK81WTP7EscgvQtIMMO0mdwPwk/qbf8e/4d3
SyiALcOLKnl6jaF/ttCfqf+0TjIiI1ItOxzrgtPanpNee0smwxHHj6ZyWwj+NhTv
qotNqZr6X9v7RG9EcSKxR70wBAJBb0a23OGMhl8T4izbVTXoxp8+Ii1fFnDs18Zh
9wWbvPl18EHcRef8CDafxr0OE2RIymLH8wm+70JGyED+/keiTf66+yw01EM5X939
y51NKBZG48PiDnoZCBrNUgE5VJpji6NNunt6C1vbREwJiCUzoS4MWw84xdvaM3ZA
lnXGJe3VbFAehgi4aTT6jGaKED4RWHarvxm/s7nSrIDtqDiDHd4pgSGkFKhAqfZL
btDrJ2Nl6k0CQDIj24dH53uE3PSprZ1cqxAjVufO5je6/Wbt/Vk53+5DS1rr8PHE
qlMpMdjvedVqj5UYhpV5mwlxosHWJNoO1MvOxicDn97zDE8jCZv24nXRKFMoGHxD
yiQoftM5mF+uf524SRr+MXBxH24YZGcDocSrcN8tolx4vt0RJvln+i29wOJ2Ybeh
BiaztyaoLANSH9FmSdZfVI/pzUw7/QiZEzHUw7km5BNe23gK0poTXRediyDdY6+9
zRRIIVOKk5HPToCI5vIjQ3XvROy0yly1yvy+xivuttYU75F0MiIjxjAQZncVcHwd
l6mjr/zNtH33gTU17PIg/UQCnyjBOuKB1hkurXRRmUy0sBxKLxAcpKOojNVXzEtM
CdykS6G5KutPDylcL6sdgctaoMyYDJnxKAXzQVlvXkh6ItH9nVqtf7T/WGJEVujn
B7lrG3OkmGr2StpoSGQXvYZfwiCa+HrmomUsBBbtSTHitcs/0aRM1rPxfKN9MHxw
LttXvfr+gmFwteor3ZG8dviJjA7QPHXBTCWA7iHRIz5Sf86dAEtBueuJU59QFI3c
8KSCPU4/sn666LSot24id/dS/GNlf/J5esn9rieiWJc1d/saG8tU7gbhG08jAeHE
TwfEdRG0P0ujV/BgziwT6Kezz76VTUb55I7UgYJUZ34uIn5HvUHMfg3zWCBMBmEx
QxtP6dOd/CuZ8m1FSE8KJqKCXNt22TBfPkJQKwhroqv7MDC4HIBRxT2QuMvETS9K
WmWQAGZSZ+04bE/92lzQRisJQ40adBzHg6lVIfWPlrHSKCsIz1xMrl5rsvf2DoB9
Z8xuoy2KgaFY3BUwYpWuPqu9JEGCX9rSRGwPXw7mkPhdaEB5mZYYcaOW6xl1IhXy
xsnODR1n6fsqce2wvfUO8YsrwHGQTmc/BIbTDJ5T6MZAJmHN8Ww+u9GlTMJDC90C
KMoTCL1l7aGBa3TqsHVFEH1xWmaLUZ5IQPblABWi5RkK7XwtHZIlenyeC6rZZSMc
56ZMYK9DfH7ci99pluRW7uCZjXzR5ahUjRyruSMziG+MvpiVv9vVrIPpQ8cjkj0t
9ddz3fpC599GwJS8QyIJ7oGzbd5m1c29v9cWNOy7K+WZ+U9mleoW/de5Ao0HOCrA
C9akEDKnQVwHStloeAHvLZRrDNuXNHB/x6zCk1fMYs1CfDYdnR6M7h0aAz23PiqE
QgIzwWbpAo0DgnE3koMaBUQpKikx6wbgjy7wJxomdm91ql+w+VHExfunktKo68jK
JSTPTUsXMMHb4QGvcEr4ET/iqIbqclGTJ4WaVlaXe2qLse8xdN0AT+6BzkfctwmQ
6s3Nkf0lX6a9lWKQ+eLiJoyRqFh+X3uHFUpTJHQTboqS47iBKLbLkGblZjr/lj8M
ItOBNQBzXVGGyb5B9ND8cfk0+1gqdzgFChmT/gHSOdr2hLZByI87ofG/EOKyaCu1
/g4GodJmoI0NWi9XzktN8DzvwNLc6EdgYWhgUXhGTjQUvLLAP+dzpAgS3u5OZqaS
kKi6hjsgPcVHBtNxGUMJr7+waWT46VzbbKsN6HaqiHBxwyCC7h6Lrdnllaor2Dyq
2K3ng7/Prjp2s3bY/T8PIMGhtlHlrvKQJa7XffLHg93er/gFfix3+mdzjGXmBXdU
sL55qfIsZ76khdqt1unjb15rG1snQqSTx5H3rdePkti7bblWxwb8etiumdmjGsxt
7piwN2RnWZNTKO9O7Z4Sft/coEB0X0ZhHjInT42ueUxPkL7wnZhbfSxkgDteU/Nk
L6xMawAREu/vtzbRWYVRdTba4mnolJSD/fi/sqmQFZQ0L6bC0SY+kFoI9dVpq0fo
FKWjV9JoJCGJ6TuyPG48zVwZcSv7C6ZRtnvyLE9Z5HBfGhHcaLVkZbhXpN0MU/ZD
WqcWtL4YxApLZqc5DQ3p2gLoMsvin/Carh34WsUtEYlSqCbgbhP38sUfXIkU8usq
AXedNOSKXfH0KPTVysljUAfg5FRzBQnYPU6GISfzBJTwerRdo1ad7BNavKjdV/fC
dxrXy6GUXqtaumhxxQLEXePMraq0XTzLUQc1v1ENz1g9lY9eIuscBKWPJjgBuNGr
f7APMKpnXYhsGjxC3YAP/hBzyuZXqrrIo6md+R3lTuKr3E7afCDIhK09bLNjsbzU
V6Fniaj86hL2dMgL1ZtuHLzU2Es2U7+OvTUjmTYuygNhAOpDqZwo40sUSDIR5oId
xE/mj8TE54l4ril5B3CMBT8WYaaVuMhp63veZIBfJeI8yEuS7cItsClnP813k9Ww
fEy6mKFL99tmtpk4dFFz6Gj6+0HWdScxKb5J/BPi4X+7nu3yOq/zU/xvwPGRwcOF
WsMrfhAG7qJlBR8GclWoBFJ/DBlNXN4h8xDrLCxgQwueyFKNfW7/sdx2fXmSaqbr
ayVPJvVBjHtIdtN0uOyp1iI8KwxIlnyNtF74h6y1Dda1s/47FLwbsX6sjBcI81TQ
2m7GT4HBWDmBMtTyzaJOPdSkEqeCt94L0jHRECpuda2Ue/iPXYGAD5qAXT6oU/xx
c555BpUgc9Z74u0wQsvaTlCH2nwAL+4gbK5nVnT9wx5SRxXbsegrJiKKRhg/uCA/
azRrx4A8N/yL4h6CWosx85nbLasRAqmg0e9NtHavldqRgE3dpMV0LJu0pvc5xM1b
fzCvQKnWDcr6o4gx1QpHPg0cCeW+YoousPieTIbmmlJ9EzXL05h2H665O2FXFTX2
MVUERvGBn0ZICR1u7C8GtMidLU8nT5mYzo6J83wAmkdcbxqCT8KxstOL3+ZjqQVO
GeNX5WmEzQR6k0pOryoB1T4nEI2P7CMtO4mstpLFR/jBpbzFu9KHAievUP/qxpgq
LCvIy9MkWAV8ij4cTAapn8cBt1J65Z2JzmOR05TyeYB4Y6GA8o+TQhllVB0Eqt6w
O5eduYm6mFtquThXIzXpnV/tqCm6ZtBYSWAZHji6NWyqTKodkkh2WyFu3C5/+VzR
Birsvi4VxHVCsagFVQQZWck+ISJgzIPC2aBpv69LTpvx+SFecN1+ylBXks9TtSJX
4kD0nJ43a9Jdnza8fTqdTCWOOQXEO7R7v0syBB9VAdgzUgIxTI5WBIiIWsHDdVbY
zVHWqKrXO8k/AAFkPlqyLRQ627Ctavv8Aa/FUyoD//QjjOd49jniW+EtxyKGotmI
YFJUUTHOKFKhv6UBYgQGaleOWh68oylcYqfqxUOs3cCdymbCgWGFD/gYzU2unSMG
nP0q1uI9V+fqfbrNyv4/ohDmt7wBD9jLKqzXI7u7kKSg0bSMQ9tRhEH4rDUyQB4B
5onABWVM9+3DXIgP4kyUP1Tlx5Ga9j1cOzsdlS56g/tyrYBlFMpjEX4dd93VREkC
6d5JK3OkVozVlRKGgSrLqWp/uZiapy6B/AXmc1YBqdTJq0kXQh6Z63IShpBK/fM5
owSWhSwrTY9SwwpANEf3dAk7/H7OPBN4m2kVD5ny88VZnNVJjfrExczWeCogvMwb
W3Pw/zkV6MhfJlnScqfdFFTXJM9Qm+S/LchUMlJwQTYhSZZDQudceF2aqO3l5Ld2
5lqC9Jpc0sGjl+TXi4jQx7NCWXiEFG15MNaqeqJLv/EbyTHAD5oLx926xFu/qgu5
qOSCXXdO0rXnPAYL0Q5n1XjbukokrRDmGgRhARXoanKyABlbKcxZ9tnMxRuLgbpC
yVe9MGJWFT5g5ZLqg/wYwT4xbjcoh56GU9g4OoMdx0ciFPeFRCoPAKIopBuOoyru
BJ8yhfjaShuvTaIe+95MWV5RfMqHpXWqabBiaYUeFR8LPR9PGbBmH/+Y4F7B5MjN
o97STFBMIJPsRBcosleHQcPc8JyzfiBcEXKWG97DN13W4r8H2qXNGCamffKpylcE
VknE7xnqLx2Z7VcSPQrybp3+mdk8n6qKXKdMSMvVoXs583Y39tqK3rMLYLT0XzCK
/q129pY58TgC1LdP5YzV/J/aeeUkHIZaZfR4bgpCWw4xmWVgTqgwyoLaD/UWQ3QR
hHs9KSQIUwJHRZa64irtPd+Vb5+uYpHgKiM8tsHO/GVaUR0p2IqbOfSGCONwIM+a
xaeuAfWdxJv4S/KtiT3tBxJ8OrVLlutwj0q76Ud40HgcX9L8AL7Fp3S6Dv1SdyWJ
pYsq6HDQjzLnH00lqksEKbbSGN829pGCIHXaD79IFrRSd+aVlihV5AHGMOEK7bWi
KIXTKj+5rwwZDPE/iAPXLb/bSegiozbqSdQc0RCpvv7lG13a+rYae9cI6rc+tdPL
laz/3vIXe/pRXSIZrT0lJUmWRWCzwrrNQKECyO3UEesJ9QnrhP7rT6fJekIOXq/p
HF8zTsXZ+NBnY5BOZKHqmT9Sn74y2n5+c5xGlT18psXErfpvsHQUg9Umdo4RHxCH
CiHyt5+yJKK+TYmxPMPhDt0voSNAzykJygIpAqnx4MEZ99UgGOkWLfh6X8m8rlfK
T/BU2dZt7JNNlo+i9Onrqx0O0C5mXJrrVaBPd0Gpe7mnajdtzk3ob9jhsSxfJ9K5
Knwp3PV2gfZBGq2rSQbF0jTXhmmBcsKenMJ6l/+W9j52C/ytDTl98P455lBjvy2t
xWqIloAaW8vE5lfxeeRj0YEpg+jQfb102gspGzQmrvV57t7+hJ4AAGjZBSjicYz+
XJR9PsHOQ82aTYVfanccIKXFWciOpHk4pfqvPZX2c0xXFROpjjGW56Wt7LlUSTUd
uPRZ95AIQl9Xnb7IjBhtZrM2zZxBoS3wUdeCHVHMaidab/RWttuWuFPOkJk0KQQA
39opPHcfK/pcBIlGU2SCL5vJY1Bajr5Fag+pw/MPd9nEKrxRG+n/ETQMgNdVp2ml
rt/ZuBNXaSItD25LFJbQIE3AsMjyPMIGZSsLNMvS/QDOODB6Ov7seug/n2jjIq6s
Cf6UF68aDOse4Qms0gmGjkQAFrZFq2b8Bn2XMvhFxnQQhMBF0mmLZfBe8hTtAayZ
GSr6vag1+aOw8+Xmuc/bMfCUncK6+f6lueWjgYGgeZ9Eg9vGoymKwpanHk18jSEI
1LekzVUzKH8uGI1NvmZoej4zE6FT1aGiVMQYO/q07C6/LrGR7xsF/az7UKLg0/cE
fp56CnH4wR0XH81ZnqgPzjDHIppg5MCPAt74TMDo7Gvm2+OKt7ZOS4w4wpBBFIWo
FQ01b+Lq0s5JvuXEUC9axbtHT892Ri18ILOg+xykMnYr3XrQeJ+RobF9m8jPJG9N
y06B9II35xF8wO7KMJg3yTXAsw+jGgQteaSgLvESwNc0Dw7+VyMb/4v08ioTxGGT
aPhMyzBjEOWW0aPNX0CxEIuQ0PCnHpadomlImFsMBAhxc2KhNDvwDs8iduAhZCfm
rla88x2F5NJL1gPAJqHon6+kPn/gzYZ8q+vg3hQU9fdegxqoytnqFUoAehAqzW+R
wq7l8jBGtPktzYnJ2xSgEQn8hgyN5SxeLgYTwi+qD8OH46KlHwNZnkj8BCi62FxA
91UWJ7PU1kjlJEUj/1xz7+QtDhbcW/xcIDEbJE5xn2q31rTxDWeiVY+2VEKRnczk
aXsf4Bxaqxe26b6G6Ik1ZXUf2emEPPUBYN0W9Ig326y5QJyhY4S0WveMuNIWOi0Q
mqXTTuF5CEoBWoaAKtSitDMvHc0POY6L4cPNHfbL12iSJmhmq2NJyKsBgmQy4+sP
NBZpd6FdnZameHRS0XXjEAcf2xLfksS3AcCaQTX78fe7te/MuGWIkCdsNejg37WX
+WpwHxGsB0rtLhu+IMczzM6bSpondrnh69AE2p2JWVyt7/YBenvrRoVE+59tbKFo
Vy0RQdKUUvCFy8dR7VppTDEhBfFRr1susLk6kwf5fCBSUUboQrJtdl974484m9wk
IXXnO+UZCHQAzDZdPWcKF+jgrbC88Uxm78WCvg97OJBvhcEud/SJfBRp56tPU0/V
HUqIMZNJD+Ez/9PN/97gXavTl6fMWZYp6cEXmqs5T0dKodKrzhwUY6xvud+P7vye
rFvHp3MUY1JtiB3AtGu+2AcOfvWqlQQX3D2R6WDX2O8HVHYNxkDeqIl1y/8wq4NE
NFJY6QUyH2nPKD/wMACjHAxmzo2ZZzoli/+BzCqPj1/UlAJu/LCFcgZIdjWV0i5B
6ZQ2FP+tX/a+Z3T0v/I/Ht2XH5OHq3L3tdehJ5Ti4bRiMq4zidtJ/D80KTmhEUB6
Fp9XnYCNRh6HbBnAvbfPz31evKtnXALhBhxrLomataMmRB8IImkeExEDul/JYfj5
GR1bmSbL0VUEeGJ1OuTkS2ga4NkoTPaZy84aRAAkH7ZGRHTH/G7ve9+mGZTFEZP4
QHak/s+SmDh33Z341EgiM/oXWxaqbrSlfqpyX+CARpjSoM5vQhr+/7dmmQoo9udZ
Ori2OjN/sB8ALtK25vKdRl2HBg2L+3PyjHX6G/KjuwZoU0sTe9Da9b+bFhV5qWjI
JfwfiswF4k9oRajuUOCCfELYf1DIfue7i9K3b2Fyq7nDZmakuo45JX1AKIdcYs0L
j/Orkc0vqxv8Pry+P6wtpFKXuqCIl4TqMBk1PWQK/o8r0F6VzqDirMGVYLn4Ahtz
hqyV5uMMq0/jYoTeArGPX/pH5EsHynvImDPIn9yCHOtO2IQ6APySzgH1y7CLnEI5
VyfSCXoR4rIfBHZdKRLLRgEWkqnu5j2GNhxiVrxKLbifqcMs4wqYnHyKXZnQEbsi
Rkyp8E947uLLQHY30KYYR1yHm40MBEYlngvhXoigB6CADgbkesd2u8ChBztGAlak
LbXyE5S4RTQCw7Ia8FikLchkHGFHdV3MskTBgAODqtJG7YBwANftpWtLt9agP9gS
K/ip8spdEWr6iOmCTh+iw+rOfbvcUEr2rFFmWC4nYXT6J4j8h+dqtmpVtwyyeBKR
htUnLkbLJ6vgqt/rVY00UDWrtqZUvc4/Iqw48pCIBP0t/QSigUu7m3jizPXaqjoa
gB8v1YksiHEPbtDkZuBqigDqwjQDQ18ORDXJY/3NR5mEyBB5N0wSCGlS5dS/t5mg
z4Xvvk9AIE4pHSxqJVPLsNkaLJqqeC5NOkEbMJ6CsrZTrDMBtnGIeg1ILvOpmkkC
1NK72KFGREm/4Hr/6tBNeeOPd7YApCr7sU2bpD4qsDLGMLAzjWhvRI600Bam4OCS
TAMn+kCfbvTr0oHRi5bBTASgFF6pPNLuOQhmUAXF3BgiTBxfXLTdVCOvDgAO9YeH
/KqsOqhIAsKBdd6OgQradBv4E01ysvKKmVF6E46isjnKKy73gIqaSxzwbxzdh7F1
aCQ91h8aJ0wrBW9OXtZtxuGgWpcHZpszaqCXMh0IOUO7EbtFGH6PYQqr/mdeEZhE
MTVnu1UkbQuJ4wS4dE/Q7a56LzNnBj6ZBGpbV7iMYp/Gxx91tIk6COYTdkHrkgDh
OJOQwfacZAhMVetfGSJIh7JIBXiRCan0yJ2Z9UEtIGYW/5lrNFb0xmsiO2306yPP
rHrVTR55jKf83kB1ufwKnLjf2jKbQgT48VjOZdDM7O60eapvAo1P7oYlennHBBil
gLN66IBHzck8+sZP8MvcwQ0CMHdfjIyoN5WjXfrryHVVqhgWCBsb1JOQrUbhYLfo
t7dehoEfH0zX3vs3lcLbuXRQtedPZhcp78abAR2LU432krZc7EQDe/05Cf3Lpe2W
q4NEeuHS+c/IA4ErIWHHvqh9413h4VflWItqEcq+6cPH6OZkr5Kj5aREM7Vz7sKp
YZz8ZAFoKdtdQuO8RfQfqrH3ce5h+2s0wxsSHf0yDqL06Gk4S6yTDX063O99dz35
o9MCPM1fncqmTitlGjKOXJaOAF5h36MUr0nimUmUq4LFFJijGiNSsCxAS6Cs7gUd
nOafmAm3gioiEIzqcPh0hfIWpdkK09C8Qfb7Y5z/hA2NMK6UX1/H2dHEEynS9VUH
ajp+ae6cSA5LqPgapVJoVziGu2jPu2hWSt6qttPtxzeHAEMw2kUtH1+Xfsh5sSGp
unyied9SCIONgbjnaibccqgXVnxQ7VF1adRWkfpLUfL9F4klTrL5oR0UMIQq7Dyg
U4UvhpqgWl0lgcNADRdfxY5Vrg2yf1R3U3qGnT1C9zOTB+UJjOhn2tIAWldOqw2V
9hOmzrs+EFJEMQAXjdtiylouEuXJBc8XyDFYHsBgvSbfVi+mmctjpxJV3K6BR+WF
yUG/rOeMFRJQd2IWDW5n2vn6i1uZ29FcwWzSAoIi0hwUFfQU+0acv7bGGvy+QyBs
mNWELUlBgestR72nGHRomp9yveSxpjNQN7k15AsTMhwtlBEpPG5bbNIFNmEImVFL
c2/i6TwopBjJs4tuFBrrg+HZKgoP7h1AAMZ45eZNrdBixCd75pxf4uLXoXihS2nB
G+An+6UI7vYRAYCOig0skVktKV+iBmrBcUz96azHV8or8v4LHNmJIc2u7Q1M8lk2
mVw4e73VvQpUX8w68aJxq0uhG1Xfm5/1J1BiIzLES4KHYBn1q76yciTalv2yqDIQ
BAW3ZdoFWw4fo6qbdEtDLy+DrkIdBb8Q9spYo+dgi2mVrunGuZb2ekGkA35iUZiY
TzCsGTb6PkbGQYDpGeO5OTqtr7/WoEbMElbepJFtlrvQZzJqV//GDfUKp+LlsUHU
oGwXq2Z37m58Fsg2Mc8WZQIzVmX5qbmAby6Idg2bN91EwxfGkeM8IytPFqjP0GNq
OPb0SZBN8meDRbFzM3Ix4rUEDM25R3KXcvl+Z9LPQxpgXsbPSbdmSj39DkgqwCe9
XJiJ/sCTYDCsQ2R9QnseMb2lPX+qMEMq3lZyp7w9dI/HLAx5W+r9sksGM5qg7ErQ
IKPPXeLxLEAcSE76VjifPJwy1QLxX9sFdihupuPkrgTaKpkh44CVtQD7vK7waqjq
i6oBJ8QIqpzABbT8B4qMUXXJita1D6KiQppwdR0zne1eW6VkfH1bzIAs1fAGCFp6
cKQ0SAMw4e6i1bzER8sbLEeubga5A1z2uRPjqQgy6OVt41IqOamRUdrBmhw5lKu6
vt2hfDsWivl40lN3JRz8YTSa2kBVScjtxfj4iFjzl28YEuq9B4MpsvaqnpAT5IG+
xvSdOnA1TqsjObjqEgPUabmCwn9aPfy1+AYZ+C3RaCEFOP21MLGQ1wqjK7f/qtAS
om93WbYONZGjRb9Ttqe78smnuIejXtd14iOHcU+WRCR8lr5CroDgiq1v2i4a8KaI
RZy0HeOabgFGdCNiboIHTy56DPhv68RkIu2OQBf9sQbAyKh7eJfOu/qqiEtnRW3N
uooWojHXpP6mMoOT0OkrXP4lHLgjpWifrngqmirpZsKYWl+5IyHSMk61Ix2y/m0M
0Ecie+jXNwGJIdkXoUi5+fW0LhSFcr58YchWb+wb8ebAXmwHBq5afJPAFJMSbjOG
6OJkBR4K2hKk/CAHEcbqRZvZbdvgbVQjXYJyuethnXGuDu4dekH5AWTnaD/ddb8x
uNm4w8nnHHs+iOhMIUOPDRRddpwhYiDg7C0RRDaqBLPMwNo87+DusB4ajTVLV9ad
GMI1M7ZxMItsNn6UBTZOJVMWECk3pLQ5aGAFC1LucvhkgaOjCkcyNxa8q9hMUe37
SaFMxGn+E5fY3hzYJKk0tCfoLA5SPG3M+5Z5wcaDnkztieIxO/ktEi23/cH7bhcB
4JR/DvU6vYmZeEgcJOGSw4cQ/DPYgcLTkQJcDehQJGj70XvP7LPJ0V9SdIc1F8Af
4sllKsATYjL8wlcziTvhzUWcpmIIjLB4LO1ZhrExn8NGGg/ReGd39E6y7PlQbi1J
YOgsD0amMnH5BRs0tECulbZX7VjOibMc1duFXArGigKqS0pFOJIlbmVXxYgmX8TR
0/OvsEpoojxMXtoYW8AF2Ai9XdWkaTj++dr1uMveh7ltcbmi8NNpgUDJaY899dwG
+RPFB6TpbUnXTFAbPrOBEjA18vvEBAHdJ06r4RZ3PM/Wz/wU3IEkTSVcZtGWR8YG
0tmmsYEuV5qlrgqZdnYIwj204qbPrwJJDT2MggH+pgaSXEotFkwd/JJeAAQ62y4E
cxmh/DwcAbh+2qxTRm9/uJugjNoBUaWjzCE+qmk/3b4+d7WNKxIFEfhmUTQmxfyy
YntWYp5qf4jGA1GTq2C/sqJ3A3X+xAxNazN+uLJM3vo4UrKV+HSIKPOW3iIx3N3M
R7WkjLTzqBioFD3ZcLB8rDhBGEIf7RATj5W1SATB/AKRye68AMvSwf9EOyrdfMk6
Ttt0KNQlevkB0HILtvRsGeGQYZ5OBkL6dYaVzuEMpCavv7olqyBd3nnGAyuWU109
3cVaD9jKbXnCavg9LtLKQjFX9cfkwFVasmt3nhgmhHQGpXHJhSK67iCvx3ZM8Qay
OQgbY+3bx6tHO9QkN9W5G3Rf8Jtdq41ET89A2bqnofWep5a+C/2R/0ZSUd8fd/y/
6W9RJypgCcF0rrG8sQBFlS/P4IZFFjDomdIDY9L4Flzp3dk2SjtWsVioJiZPimPD
wsPIPJBC2aVhflsRripNS0g+q6MJqzzTgXxiufu5Z/32oirj2lC1u/cez2dCFPzC
WS6E3oqOgai0qlzons307Gk9wGU1vuteWitkZUxYID7I0+f0VrPyMOpkz1XD01Kx
6uJecJWnraMpqWXz+DTdU8lLpItNiCrniy84C8WwpZtLx/AqjJLvyA2Op3RXgX3n
c3r0wQZNhEosm5/M6OJ/J9O+B7506XXmde5Ut69INIrXtAuErYW0lnKWZ1MdEamP
GfQoRIVDXDPZS3O7qS3fI2s1P/p51F3BRW8uO8p973WzhCmIZE5tKnmgMZ8/wZOs
PXAmxaOvB2VLsRRUcVSwdDVsbllMj3sPYa5B4ZDk51LqWkYZcC4bXv2+A9jRaUQ1
+3gTxOxcP/H1N2WtsmTe//q0mk1jm0XTDXAWwcmtiR++bRnGzZkts6r9Txurf+FO
vxCjvG1amDvdN3yvRpCNL+aFGsOJXR/ckR0lmZOWdzMG3Y9YOLVQ/DZiQjaL21QU
wG53fZT8FFbkgZyyk7Rr/8TAX7B2gBp14w3jZKtZTOIxZYNRP+3omSzv2b+EHKhb
FU1lNPAviIC8dg8z2473HvWzTSNkeLRU97Q4rTnhY0QzzAkMPg2OG+lC+WNviFyB
XeIp6Ty/P5nduNtfjGrwLk4/kILscoRotbFJIxX4Tzm1aufcN8UdaWOyuhTdew4a
qG4xVcRo2P0OrMDMkYem9khgy4xM/P+FT3QQ3/l27DZotgQNmkt/DuP5Hqh3Eed4
XGJc/Wz3AcHuLXNB1+lTmLcbXuqqfQhcJQGRy8DMIba8tMGsrf3jPJR/vFUp1r13
aPg/ASJUrHJKUBHdFU07lbrRP9vZ9Lg9QvwOcBiubI/JV9D9fIAAwYU/MaHZg/Aq
koesy/vU2gvdHwdn7wfFlnnHdyusD5yu4ky478Ie2i6+5NnpJvPbmnQMo416bMLS
4j2mco2y3aLhdslg7gkuBNrHTXVrpvofRaDLIg8JyRlmRrG3VCfGcukFuTYPCsKh
t67vFmPbR0SWuTrLbUmV8lc+lpekEQQRiE/UwvmB+8+ehcyBQ6j4PoNf7BTuYFEf
L6B2m7IN/QfPcXUIkZAtPP/b97YOMGrO+at+AMiyLHbCACWOoCdBggxL0if941hs
h29xPis2yyKJLCFj2LeguxBE2orxLiUCiJcIKhEKvIu7Og/VC58lL+pFx7QMbIpS
Yc18tMPUiHyKM9bg1X4tAN1YJrgWAqOcSGWdUnL/spr6TXj1biFCVS3QRUpbjDy+
X44umfByRcPOqPlIsWotsV9Zjhwm+NPocDj4Fn+BK7/AZfwLzRBZQYmmPEu0xjji
i8q9XXakr2nslCxmx4xi7IJfI5TVT8IIjYloLenlv0O/1ksDM9J20tE9wOmpHE6G
qnGxogUiLCYlSg9IQDb6n1ieG0K/ePnDR3QscUUn/Kpi8awtoZWmqqTZDec0VtZC
O355gcpdDa+p1QkmA7DyqYsDM+7MIhtBiPgsvkbCNI0PiU51KmuOcEBwicaLa4e4
LZJDWJB6xsQBrz3HtQB6ZHKqELgFUwfVq2yJEFg7pmOvt+BWpWN1PaKsjW8S+gU0
KypbgOPzPa6iNvfLX0uhSbiunUVqD6+PTbYd6C5zU8IQcjqP6aQoWPq/aybi7zWe
kzIEOVoY0x67iAvj4grs+xDQT5XusEIzylwZa/RWUnXdItnKQR3DPVTEkq+a3dnv
/0uCqzypMRybJ/5LSzfoJs1CT9wmaKcC9nnwwoZmPOi5HWrlEpGEv0wtdwlA9ELR
gtF0BliTZqiWhmyCGXFuyCAAigzfW9fP3JwB+pPfcbqyJ7AhR9AwUGczcwI2ZiiE
p8ie/CxxEgi9WJM+ZVhZuzK+uc1XlzhbELIH86pC286ZI+68vX0timepT8WhqRiO
rxFYVN1lpGVAYH5DZf6hREkCQTXeMpaMhsIJ5QqrYTzx6ngiwKFPoMfp0BfLsH92
hkjrI7drXfPH+2wSqzAlMfmxONRekTeHML3lzR5VqpL9tD43f/S/J9hgBR08KIli
DzA/AnDHoBnNY9QQZDx/rKHiI2xjYN4e8NbKKnj3IZi1V8EyzwU1Srd3cesZu1jQ
Cysjo8SsaMi2qo0zcv8CbQqmd/XUjuSGpinHeQE9g/yJ4dnYz9xJSbrrxhS9lsYr
cwvUPh2OEzIfdAjF/mHv4PEeKhDD+tWTggK+kc/xurkJRBvJ2rpc52KF8N1PHTiP
LNj79iXlCLDWzStMYdH7biSSL61uRiUIqdr2OXSFdZPYubLotyjjqwjopr3o8rHe
DYEBLLtvq3hDNKncWEe/yerM29w8RpNcAl4lShm7fjme6s9cCLdWLhe3SWnyVX9B
FMb9lIg4TooP+F7A/Pn3BOLxS4BSBDn+TRzyxbZbGSQ0hsRl98ZnbVGK79ztTwMU
1EIQKW4XXhZbpEwa6kW7Ku863eT5me47/GQkkk3BJKjLUOXTZ+eIUyWT7pH81xPx
+fWMxgIPNp5+o4UFRDNH3byWtd3nBpI4DrhNdA7mfHUbOW3al48KiNFC/tsl/40c
uMW3xQUgOOWO81l767A234yLBMTik9UGduVygrokwALjO+LOnmHITUkFDsfd+K2L
dOhNJl9+Xz55NWlkjwbuxF84kWxs3E8AjB8tBnrZhNkHyHp+VTVIsl9vw8YehQ/2
kWheG1lPefAjwYyFdkmrcGSGZ4sw9gPPv5FW+EGJXxweOMjdmubQyUj9kQKdlofS
wJv2pr17urlzLOzsBqVgHhGTECLrRr+Zq7UN4LTovgrKMaXEO7zNGHtcVFxvs0+t
A08mrkXJSN/5oPNihk8RTGsMN3s30gOSg/vKlJLNZZC6noAGSunnA4oLvFZkau69
OqeHXlIponX5OFL20x48q/IGz1ofAxvgxuXElJvyZCuyR8ratsIFnIfbbfQ3kcJg
SEYlDSfYwd2wvCfUdAyxZlektGksg5FHVic0aydazME210QtXI2XVllcPnipp8Z3
4fzZI+/bBiPLRWrnlKubtnD+cxVRqcUJtrRpjgJbrLiZI6m/qBDI9bHXP4ehDMff
QP0GN0lNpklaW83jW2Xm9qWwt+6gII73deFxjvPeP6ToQo1u6WJucZcJyBk4u3W2
BCbFVH3PBfCuykZIJTMMU8WiWYY31yshRg7+4BVswQ4rVL7lIgFBIXf3MJwYxQfn
qvi/0UgSq8dqPEhillTMm4H2r3UDJOkDbgz1HpgKs/V6eBNdHORAVbzsNxmcI/tb
I15TlJEbFLEcVReYezPsA4rOuscPI0J3ZZGPYn3yVo6uZAsgY8tBugxAMoqPz2lg
nTEGwC+alr9naGcghfOPwvkx1lgg2GysTtupk7iRusVy2t0Uxl7vaNH+VI5I85J/
PPqbBinRjjF1dEyDrSQ9Rx4+9G6Z+UangKfr2r3sH3SqPfPIJgKr6cwG6eFRizsa
hD6XHb8u9oAloxRNdHYUx2wLy9JlcvKprjAlh24X34CUvjkjCsBk9wshrs8cHELh
5BpRrd/fIDZg+cmoBLmB4N2PmpzesyGIBEz3Ug/ehxukzsInWNydYK8WH9E/+ZOm
n0SVicM+bapGLx9/Hoq+Q3UXAbm9yDZDxZSrbbiVzOVKMG+/atcbCjjgocmWTHf1
vuR6FyfWgQgtg7bGMcHVW3G8p8kZgGMAvJievkZKkbqLnjdFicgItk/vTibUbxTb
48jCjHQitgKD0hP9pW/NNrq3wgkD4W0R4074+tPTt51ueZ+4yWgNl33KbcMpsqgy
Y+raizyaQaVXQCFyDxA7WRPY0RMTQQEgdcXM+T9biKrbF68iBQbxAPSCQ2epVqt+
PHrrQWK4DdrCrAVhvLos8aitubP8VCxs5g32VSqRkkVmIgQtHFv17eCAPw/eZsMV
kKgn336blRuOKQp+cG/Z1T7XjWFUWkJLCDE4Zl7iWSAFDcip8fL/10Hcs1WBwKC9
lbvWmue2RyYXzBWDU30SLW1DN28W0e5thcRhzMt47zjcGGb3sYDhszn1mSmuWxI3
6Az6pHU7NmCuBkZG0+ZpISVfNNASO8zLTf1x3i+7lhDI066RCwM0klOwZYFTwxba
DPu857H+67rVnsZe1NfpfEp5gI6HMZX6UU/OftupR7Baqv2ikAWGE7/p+OY6nKRw
qvWs2rpQgnv0yiYDqUbBaqsh7yV3SgCo67cIQBL30Y0BRUbw9ejvaXzyfI7IbJwx
RGyGJ9KQSC1skpUCzVRFM+hLE8fQMOYXi6tk2+viFt45ekWcHxa+nVCA24zsOPWF
BSxNILaIDR4hKVJsMIAvTVxWBHD1J6oXswziozp4GLUVv+hO63BwiBvf9IB2Wj3Q
AksgrDvdR1AZDb0RvbKYKN2cD8ZHOuD5a7K2VVPQSaMhZDBT3/InjNAUj0IAHA9Q
KnHTB1wct7hMwXERTCNadH9Rw05fCg1IU2PbF3Iz+kfMskBtZ5hSJK9ZNb4fZe1c
Nuuj9FA1cUDwaI658+wMQ5GPzXc5Kco8bQrF8gGzBYGGf1hNYVXseDERpd8ZOL7G
GbqWqp+y3zoiuxCv5l1S/hHJ+rpSZMY2m/vRQ1Mu8t9qWKxted3mzaFU2Vfewjbn
0y2btCNYMDhdMyNHUZwdX3eKs4N4hytWTTwz2uppPucdoFzRmeVxKUQ0ogyMnfFT
4ZjV5o4hdW/fueP5tHUr/QuoXqxMwP+A9/anBlAace/AnrPR7uLNfqGiF4HOFnDm
T/FMJFB0fRYzBil2HZLyKFV9MPH1fquHfDcFYkLe7bMLuepGarulk+MkkuWLtSOn
0t1rca/eKaLy33L05hfd1NEETkg4alO0zkci1C50w24D6DldJnYsl846U9qJ9dXp
3Z3T2vx9UXGarM/2V4iNQfIG2bLVhM9EkSp4WEuyheJx4GzUm+S6EkQ8u4EZgLTx
qxd70eviEG2iBC0gHC0ZIzOQmbSc4A75FeF4TyX4408hWMh0RH8pilWX7C5FFQmh
ys0W6td4tOm61pHXNTInJ8inGZv+jZUTAeWYQqtFMAnOjgBcZOrnANWjLRoe4bDy
uIWGmrc/LKuvwHzyZZ81avRCB20w55yDr/Bnm8TTXdarQxQ72hPMtO193Emc8GW9
aNxiwWKJGswV45IN90MmuxYWbgMfn2owXNeK5SRwHx+sdOpRg26iyXvgctoJFpwV
VPrDO8QqzQsxRag+a7wujfXvKHDWIdeFYq8g2mHGfv/0u14jdwEnbmULMRlQeo/w
4IZ8psmU7WnAsF6h17D8nTlb/E389kblx1XL18x5L3+ZodKqefIkEm5EhLpA8Ztl
YLYq4zhkBsUCUc+ohovyV8BXaoVy1eANQ6eR0sqxHFdfSp4kIQk/uDX18M6yi7+f
0e4Bg+DgCS9407ACIcM7J6DDwAsu6WLqAh6yet9QNqz095pFB+UApO7gnZvZxuuC
7ovXAf0JZ0gxkIh9egnLkkguXzRkx8S8VlwMI3b6r2XC7ibrjk7qFY0aH/9zHmql
SONaqCotZQQbdLj+HG+6fTPZ30sW/WZFeCKR7M412SIhZt/LNEVkFdZ1qjLoBMoZ
x2HZNK/oK7tuIa5VZVbUFFdIUliDLhsN/QbJFgqvkoEd9OcMm37N4XQWmx5NqTtY
JSBcYJcKdQhi0lQaaq5j3sMpMpoTYPqOrFKH43P6j0Xhl57rsHUKUceG2/mF4kaz
tmu5TySv+/aW4vpMxUvEQLXLRkMErDOWmBNBF7Xm+f3QvuJgna5EL94P7FP/yNgF
YagFpbBNAUmQq51XqxiBQSHYjEKNJEKOODAfQ9jQpmVn0MueiTGhckiO4Wp2dpp+
afVXEE4UNvS/plevQy0sV1JRS0ciVXTJ9oTm2HqCIwRZuWmB1BK4pb224rJlBNpp
w5aU/c1vQemYD/CV5sdjRmj0mr8iqcpW42fIv05ol0EQ5TAk49Bs/L8Ha0I+Gvkl
s/5M++9f0e+nhjbPRd6ARnWr7ATe3er0Lpma3ylBIHsJwp+WlExAzPxgzqTVx9Ak
IwjC3+ShUDEsW6V/VmKLQ+v7qJAr9Kmy0VqmYf2za1iG7TCeSbOIm95AON9mQVm5
k/aCF0gWv6q3QRs23LnzCSQsyyiUPK+H/PZQdh2V0dfbCjQrhrgH8iZQ5FqK9Ecz
hgXgd7++IOSZvFQjmq81zAPfJHDDz/BfzzOgzQC/VW3OXRU8H4xML2r3hY7+ferz
Gc8biV2dzjo+6s2xXS6nSSfqMUFQuean9xifCFmkS7WhjDn5IssO/M18oR8leojY
jR0NuyMHgM4ZMyBvVrSCrJ5pQvThKlSxVzMm9VFC4toMB3lcHCQW+5neVtWAoh1V
yZSqyLdSYeWB5b853O3fPXQEsvRVRMG4PHpzjyfPpak9H7i6hGM72+QDwRWBJgad
woUz/pzZBTdCrAO47ZDx12w+5SOE8m66NGiIepvZJQdN1r1hMddkaBjDLH5eZfAn
yKvhtVFt8b+JcOA8gb2RFAa4dyo1fWOIjt2BHJhvUT0gjhW/sJUlWReNo8n8gHuw
xIt1kaW11OQpHkuNcg2mE6WZhWnACYkLv0/RlNDsCrfg4tPeQbMMUZxVPczx1c27
gLJcOdnFCJJASclEjXQotIzIWfH0AGYU7k7p9DVuVdS/3yrpkfVr8Rzorc5c6YSH
qdYDHcfoDMjtXXbN9+q0MZlch76j+S/wwpfTQDWoYEKMztw+ACG9XohFefaLdAaI
YQQjBh9UVG95JYMCl8FcM51dhXNWDnJDVPWaYHwKBbwkjhsgrSWKrlXjTuM/naqU
7S0Fu0Hrov+TT4eG5vSyoL3Z9+h82mc6b41BjBQevFYqT9bdbq3N4oGSqaXzQI4u
15XQhw2SRKFrwdtSUjEC0d12/Ut4nu2DzUAIz5d3D58Tv/L3hen5I/At/XUXc+AH
a5rAUWMQtcxok3mDIy+tzL014k78PvDyZggBBpaQz+vW+6spVYQVaPJ8qro2+t2b
l890QQqIW5wSRdFNXwaLMfuhdhjxEWJDcswZPUIZ6vSnfE7ThY4PYabzCWNFNSja
CJWlXIUBDhl9Fmoo0mvgn8huW+fYePyfwuVJen7ElFNdBzb6RC6cQ3Tn4IuTpQeU
+rDHoVAnXTuWa3dTDnsQKd34dU22cZH9scaABIbgGdW2zf38+V/dW+Z8EXwM80ib
otnVYXK0VKMWpMxHb1V0PUBSZUuJXCHE10MwHZ/prDinWrfTs5C0bXjYGwOhGsAG
AYfYWuNWxfEG5zC8B7I0cZyseQ02Efix5iO5McQPSqLlMmubk+LDIlWczeD6Oc2K
kEDx8tzwrm/939cloMEktFGQY3WR5ENGLz9/HHxDZEcFbLoNDFAAXUs9H79i8tre
Bq6G/HoMi2YmHX1XWnYxYUAZoOeTUFRz4bFP1+tHaoRLFzZt5c6pGflx2bOGxF6v
y97qMvRyxCCnSEO5BOLGe8LC+sdx5/9I3KzJm3w/coDx4GiOyAzuxLv3mPSCziTb
+HfLK29hD2DFWw3T7XoTsYfMPKqY4X9B7ZyRZ+EHauxCKqpFGagE+jtDPdJfSq4k
V7G15n5E785EgQt6WpoawI0L97r8C5u2mEC8Y2BwEPYE8tlenwLY3w7ZPQL22Tw/
D5rap4sMmKMq1CYXuqRJI+0mAD42vD+EUjf4JyZlWkOeAMWwqMz1wAvc3mTAhXbd
RCtnjdBFhso6yczB5r+JIv14v5iEsiIs+gzJfcOt7BnzSQvtOWJ+Pt135BiTN9A0
VCsY+zMIIWsJ6Nohda/QiADMBS8rzPSIP25+vYijEX60nWmXpDE0ZVo2JhMifuaL
J/mosAz4RH3s5bx2nwL6PE0WzAYdEOspIvvFFYIcsG9nvQM4wTwxo4krDUPYln7m
CIrfml5TsQmmDqctnoXLEJLIt1+D0rzRvTplp5U/VVTl6k0bOCkuTpuktjwxaS9M
UJo1wZ9+fvwHgXBrxYtUXSY0AP8EgmmtDSJwRfI8ngzeANadRY5codIWH3h99qGo
NTq16aVP63aDu62hDC5Z1ZYz+5a4auDXSvbXFcpL56wvBipLqQzzh0bKeQChHIPm
mfgckRvpeknT0stBK1W8ta+DSKG72puNZWdFvjjyTSwciknotIdGLcaTCaNMJiKl
0vUegn5iQe3oXX0/JE2jQXoN+eeIdENYOlzImrIeK2fhp54davfZ1EWOuMpGWqHp
uoLqxbQ8RIEBc/NNwHH0255km9Y8g/Vq+tM3F9hd6CVUJG9d+3gne24AhD3igo0O
A7uQqPyvyT7w0LPM/uizU8tAfQZu4wcI+abVWsNctq6kYChM4rk8XibJlUIK0PY7
wrF7Ur17l14mcUP2HUWIXVScMfgFi+x3CnU6Gfq5mRDAGUQxrnyLhpSqI9ARQ15r
ecv8LCn1ilm3G98leBd+q9XX8x/ZL10GehcBs+zsRgI811sEWpswhBcQMhCn7AR8
UZTAL8Uuqh26HufTOq8vIydhfMWL8tuDpFigYGCRpNwyN+GXQA0od0LQfjh0+qTY
s7xGikkwEzpO1oTW7BoRYmAtUX5ydfWGqdvKCuu/lQ0haruIOTpYsS+eOQ/pqn+h
k873hiynpMevHHS1a6qyoPkOJz9ETgxGYxHXD/oYdCDo+cOl4OdXejCCzA0i76uB
mf7/eKi4yhsM/DJvwCR4Mn9NbYoI8ZFHqN6GShWiRzrXOpDni4UO9RpSM1Cp1KW2
CZ8pS1K4JQyMkDWz37d4ps5lJiszrBcW7Z9BWk9ep/LhFlYsR0qOYnGbrzIV9qiM
GzqzOK53m7dTp8N0T3T0UnfQEt20M+6eX1JHDPtKmLOKMZecRdhnDjDcdFLsnAYe
7wu0Dj3B0QKL67IWif0h4KWWP1i7GEWlFwcenJ9TFzK+D+kuayyLXaWwtFt/zaSN
4Z28eKCEN23bnJkaH4G2iBixVOZkEI23Q1RDv1t1NF3gBv5qZwtjExA0NrmzmCVq
saVO8flgTRakaLozA4FAkFFGHBKudDT4nQX2AjtFO9yPe/QsulMX2mH2zh48r7bl
ZBJhBt8z1yFO+QDHtylbp2IKImScYU7uo43BhiI3IwOBhz3hzRjQYQOsOLHlJPVc
IqT5jCNO4cAa1LmblVNYiPHqCWa+KI192X0Cuh52Cf3TTFtFg2blpsS9WMIG/TzR
nJQU2HI8q8QJi7az7DvFyCVaobk1PE0b6N8l4XO53x+Kfu2pCJPjDM9XAaQMiic/
mXBY2LcT1AqdwhXro7Ae/1m6byqdf4RnhHcdlcLQlKRpyVo/FL01kJs8wcOozfZG
sVz/rl5e0lRctzFjIBvHDEV9ZMtnlpU375QdoYCJLPSBgZAJIoB1Zgitxc34yLed
j3VMqAQkA+9EH/i91Sn6rKMDqV/Y1sIJRQOmb8BN/aiPiID8EKHG7j8cDxQiLiz5
DXOy8naQFT8ageryGO5SQXIM2ZJXt3pPDS0N1/qdf/MlN8SiTbqsnBqB6KrAPEEr
Q0qrm0bZOUbNvds/jf/tpgn8J8C+uPeEka+KGF4H4ctJCSevMwSlhOxAoPoHdwl6
O74CzsIfl7ODPu2uXdPsFbZ4uqwXBc9SD6q2FOFAPzTXsEQWCHfcP20IZ4YE2XiS
1PUdebPUQtZ+nhb04Nw0FgGZ7VLSdT9+LC+zn/8vzAH7YI0EAd0ZfA30arox3lYQ
tDkqiHSf/2qfrkspmQzwq2O+grVvQVXcU8Zeh4p7z7T39TpGsVjdU8hvssFVHR5f
5PSx5DE3UGlbLwt2JgHHx2zGJCWXBig5tL8I1jB+al/HQ89u8iQ/wLrS2E2xSxXc
TFBDZsbjZTZCRlbSzogGndjyBL1CYiJ3QCniLNtMlYR9hm3FFRg+QZjWu6PfP84M
YFXuki932wXj4Rs0wNgwbX1dYMVvCR2+Hgjt5ktuKXc7fmAtMsNgCOCYGW9D4+RY
LTbZS9UWPZ8zjcYR3LYm1bCZMsgBPz+rmYe2ngEQQAp0QGgRR7tj30UTuxyS6zxb
RztYWduc52Hl0+xDxcG2/XAmbNwCpYCABKwbUl6rcOVQ5L6M9Cy7s7rdnZ3o6+ab
MNH8zt+beSkguKbTTjrjPE30vi0mVLZ2hLThBS9CIZCGXru/hB5BpS3RIyLb0JZW
hRWDDlJb85AU6jwAu3ZntBy7T5fToicBbhQfEaWA1a9tejru1so2jweXGo01o+LW
UFOLeQLaXk7YLcubkKhf6Pn8pD2dCE9wobEgO4wL48U1D1eszGO7YsDMSvut5pb8
HXgADqPevfTKjhP5QpBd37kz/l2zqfma7PmdQSgZdLJMsLWw1dJ0aHwi8VVYwZ3C
Um89ZUiPHdmBAUJL8x14vI0Bc17V4PT6z18ymHUGRDAePwVbLlHhDkDf/tuOWw5r
x+tY8oYOhVAaAnnXG6UrPFm5VfUPwAE5f0RWV1UpugmKanhPFR92zogHrcSlo9a9
a3eOQgPjGaGrWPR+leOEugcjuU4MX3q3+cjCjLUwawPg3zY7hqx4AqFF2lHqki85
14oZKiB8HvUT9dsou0zex2oWSd3huPoJEqabr0M9cC6Bh0cTQQX3tPbVr8cl7/+y
d+6q3d5ibz1Bh2NBGNCmh7QqMH6b84AiR5sbyyKfrUvvmY8iRKVEWMxhPmaFQfaL
KzTojunpiuVk8FJGNpVBUHgZMbXrIZUbbQpPjj4ZaKtp7UQ7tBZzKq6LB258glKc
oD7YYOCrzqrnJ8V4rW4d951mHQoiiQPkc3Ntv03CIUplcaGmEmDpv5GkZ+QARduh
NhrYmbPRaH5pm5U9vRVTNpe+q86hjpgBAJgnMPSl6xeprCNMT7U/weSIOxAGxYvu
odsa3qZMaZLIpaCM46VmRDkQdPZZwkxgH0pom2Nmme7Eg1QCnUcIdGnrGECWwqdy
bL++gmHn+l0kViHtLWCHZzACIot7oKgsDnpKPexHtTqq2Xw4gbcMP7JKohGZMQ8w
s9OR2U3kLZ2Pgxkn+qnXjOme7enApeJSBaZ57eufIi2wuxW0DOXDoSrlW+MqhGGd
+E9bDqPWVHTOrTf+uUj2xVWgUBMri0dUg8JbKCLmW3c3V/z48H3IMQ8YGHGudrYx
ApYEQwZkznUG+QY+DiIzS9GU4lc0EWMVPJmAS1hlBLGRe4sKZgaG7WIHFefIAlIM
7mKm1c9ZpjXR41I9Nr+dSL+RgbwQQnAv3CoIlO/IOwfWelcRrixX28eCuQ8zas3r
htWD+Z6r9sSxjGsEs7VKezVaotClO7CjGzufeqITAeK+q0gNTCJiu7jHyqjmZWgB
nDVxC7Udl1I9haXMh2R//vPYgHJ/st7++ovGw0Gfkqj98DUuN+6Zjl/s6Nlf2ZPZ
WIoiPYkIcXJwrcK4mpnmsbk9I6oEnLWE0R9tMsbPzyqNqGNPuLVuCuPKYeMXKUz9
o2V+l+vN7raeEcNVG6AT8hSrGt9uZdUYX381yYEXhK1G5WTtqjppWbsqMP69rHaq
80ct/gexC8PlAyUrrMjcNP/xTJvOyGA3mfBhnAwFiaYVJraiN9p8orIQ0cwdFBaj
y8qoRRNVV8QfBp6jIyFtQDqhpVZ0LkPETTz+Eiuz5pd64h5CReGBHoeVKeHISyB5
Md1hw/uZyqJyzXLm/nZJnFccoEXi0pYK7oWvGXLFC48u+3jujtb5eywaVOupRo6w
FMVEEj6qUPyD77KUkqJngzue7Jz4TBTeWyHDpToTkciPWlEn1e9g3N0wj7UuMXcg
Qadi2n6+yGy4Iv6lE9FXRkWGe+BoZLGfh4b82D8ZpRa5jevXDcc1ayu/kQqnmFxK
JNovDfMANEWzYnv9d258jiM5YIFR8+9tp/NuebuxBxTZ7tRRdNXz36k1VFF9xrrE
uAYE1nmVYdCI+mst1YCi9VGEYx6YCduVu8eF9lRTk8nDTeiGcg2BWzL+JgsTA6e+
T0khfpwHSMCmMqJZb/FMEdQZM20b7kO9aNq4STyJc+TsELFTVZ3F21OUo3AVk+C1
hyhNU4SvsGwbYOqUDLs1B1deE5B35cBDij6R1HLLdSBi0ZEc1oQx/NCe1Ck9S4p5
cMerv2yfQZ+Ur2m0MtbVg+X/weFlmMBZqsuuDKms1z1aQi/60PNtSYDbUlTd099P
dasoiVE2FKxEDrDfZ27tBodI9iI6Ukn7J2hw/Zt24xP9B9ul9tDKf4FdC9GHDHFi
9V1MweOEU0bKVXx1W+n4/Go8aBOuBlJOomgzEEj30DIjWmxKhq0daK44UVvd+oO6
sAXHLNyo7d3MBRdSq6uNzxq/We/xK9DcHT4btxRmwJ+IRUzpJYb1Wd6JCPADBF2H
BCF+clJ093C6662BAP9wUyGRB3bn2Ro80I66PhdbagKkNaJLVploNo/of5DSpnU5
ifXlKivF6rQe4PLJkjda9WsQZX6Rx95/P5wd19lc6thsZXtCt3VZ0d9ukPKGX3x+
9X4JB9xBjRAqhsie6ri6OSg+BULOaaPHj/Qp8MKPKWfLqNqkSK+q4oTFGYD+1C3g
e25iiKc6pAiPq4ldUo4Qeo92IKNXZw8Ej+xtDabHeEyBAsNnZ7zUvaJOoL6M179P
yTUiSYzhkbeLsMMiokvrcuff0kiN1FJ03C0dUVYeRYbERf2AVjvYc6uUI7gEqWBW
RFNsgy4D8akstNkfXxSwWmywQg4pCZ9y7GODyhKk82+dZnMcrLddB4A22I7tM85i
3l3q2fsgoC+cadyHTjajH4kUD8xh+ITSz+ylqWCNoyvIcnNtMeEmUSNyXlqtjd6D
idPt2JJn/NRcNF+Drikfp9MppCtM0QkbhngxhHFel2C48+a/65bDFpBZmAiX8YIU
7S7a/bty366vWOWtWuw9HztYBAr0wVER4P6Nh+fgSB0505LGuqY92qJZdus5x8X+
MzHNTqSbvMBLLlknR9gRGpOvCyce4igyOEdGzcotL7bwqhx+LhM8wt1vf92KDEbs
cIpVj6HkAsT+mPJGQvgYgAsxJyNWOD32b3C+JosA4vmzARJ99ekJFKWJ3CBv6Bqs
ryN2jzq/m17G7VLFKke+WJToYytbi1D7VqhInyLRWy3m0hqbE3uxRX8lsCQxC7fg
b/D6bXXzmru8sWp1JvHttbFGeJ9nX7WRRDcS2hgBCIoybqmj36V9MWTVPiUMJRUx
6y4Zx3oEk5vvqC/+bHGgU+PinyFyewINJ1DZgaEzNV2cXG0Ps6qqft0+A8UC2Y7c
I7sXGGw5T48OVu84CVJso9wDj6P9sjftAD4pA/0Oa29bgjOD6O+HnTr4X+lbk5CQ
ar50Bvdx8ksnkVyb/TdeL2STn9Gas+BckkcyQNGFuCImyTQkH6HnyvI+Jq3XnH+j
6MvYMtrG+mjTTP/VYhQPiI65AxNIVItalBkBw0cCn1c5b4EFhvzxAGMK5SdLcVbw
NSIYmMAXfytoY/51sURC5V+VOYN7G68tOPWlM4Ax44PhAUqzIUMiZI8z/KQjMCtV
DKRlYLtmn+u4z1w794goHtk5WqOK2WYCQlb67kVrUspSYtf7Ys6BLKa8rCQMT/pj
7/N8+9HSO9scalkMBgKgboQluliXE04314BxiwFEIMZu917EAcYIv5KPerkXKsXE
qmrUSyYyq32b6x39mYQ3IPNtj+kPiDPkZiWMLZPgQic/46W0JElvER1GMaQXE2Se
YKtNUphe1M/ac4aUnZozF/HvTrm3ZDKp+mJFXB7z1NQOOj0jXcy+cTK2JuDN2fZq
5mXQ1TolA/FXGOBBDuoT9NJO2eRFQUWNOpGWaEWlzmefpi2XYQ+bQBfB4Hnryljz
v4Gb0qYktw137dFY7Jum2edC35tcHW9HEUJyx1R5V5DAnzJSpROKtLAxTCWHNahM
uOK28Xnj5c8g451Mz85SZcXo7HuoPLCVmT8ff4jqkLqPKlaNQMq75mJpMf0sAW/y
sVZjTstNmpkvtYWTb5ow6u/S+8pgIrWPvcN8Ewb1SiVAjE7lNZPUmU8+7RD18TsG
2k2knwGu1gZqvuT2bqZlV3vdYPNVjsEHmHiVYA3tevPpWv3bEXCnnXssUbF/gsfY
Si4CuGFZIyhEpDw2H10sgxhoz5i2jHPFNUT5d3KvC1aCo+sqRgzQkSgHJEcUs/Al
XYirNVWVYGag8JPpoY7l/x8WNqUGDt8Y7CBepQB3cKukGwWwH53FMrfCQ47uVVA1
iP7oKa73ICtU92dI/+Sh/e4/MenFw1fH67LOwKSAjIE3GkTl4q8RJkIhdOd+U1xx
TrsNbluMygo2chy1jOZ7Vo2LoJRRYJA7OV6yUrzaVIYxKQJfXpuakgmcjgLN9hjR
2ox61sFIM6fYuJ7tW/11tr1LoZN8qZvOYlyV2cRaWSw0HsbqD+t5AH3EC5zAE+Hb
Pb0mO1pWLqrApwuF0xTCp0quOBC3ByfFzRtP4k9B4A/l1QxnNQCnkyYmEmN7ulI2
8SoLYoQxb0fVDZBDDsh9ueGbYxOiz2Rce+RAkkS3gIQJcCPnaiKiB0U7F6ymow++
GAe534boCc28sjdqCPT3xPnex3eKp8C7xEkMA+IFOtX5o+amk2Dxy2KL+3mpe1OH
up2v5NLfpFig/iBaqurXVL835Wpz0IS+lFve/z9YOOuosZtwSuB3mJCp3KnKpi7N
xPODzHKYe/1dha/tzIiRrAAjJ/E3oKB9m5UZhRplWhFqN4vNH8Tmy7+xEPJSm++G
Yx5nURMjidIDqU8T0BEEP8WGvcTxZptGjYEMd1cyMSdPHQdS4TL2vQiza2wRukTv
VczIkknIhZqB8B1IHzmIrZWQJqbM1aoCAhU5oSILthhbAJH0zZ3broyVfzVNpxtt
1rk9mX6HffcePf+gA4R7TexOHUY85vRqn2+NCu5Ul8AGX9RySPpzTOG9g7c9qOJ4
GoGPyMUDKjaxgKBNin1E350wgknJvqndHa3GhpQ54eU3T9fy8PLt8COuDTDnipPs
wyC9s/QlDI0zNyNnMl8l5k1qr0BagY/2Fn4FG9ChjniHExwopTcEbea4JAhwF/lI
TB6WKlfYAv3o72gaf6FR9NeS5qA2BU3lLWrSkpBn1EovH0VfccT7g15SFzB208EP
YmZHgQrtD4RwjB3op1Za2tGQYc1upja8ggv9wN4eO65IntC896Yffy0vubLjgud+
TWwcwFd/C1R7Lgj64x1buSJGhX2QJnms38uWk/v2+2bS2n+SqfwL5EP4O/rT63Wr
r02iRysjkLF5lDcV/gn+4vaAW+VWjPFKvn6xRT7wDEnn49Fxl/xWBncD1785nHY5
2R69G8W72dFjLIzF9wh1D8b0RQYAkeWd7SO4xgHM974degdIo3ZquuUG1oJ1TGJO
JSlkVC1XLOiHe+RBLxOEhg6wlKYuP0lCAqLy1kCGJxNvxv+U+T2Z+BF5Zp3zR/P3
jhAAJGB3Ovy+la6VK9zppfluZTGtj3d79MBsMcrxAZXp0wS+8X6Ud5eRAsH+haSs
XoYDW+gWvOTLiTC/35ve7V0P7DnW2uyZPMdskcrUwujUn2829tvwyDCHNb51QRQM
gm2yP5PUoX7ThPGOlOI8jdhemQW9TJyO5u5fePG+7ox6C2ch6wy+fGQml0sddpIT
Nt8o6G/syZxtoCKp6MN9gdSSqnxivybNLnJSm3hUAv1mc7K4gbTPf8mWn2hLw1Qx
pI6uJwX0F6iJbzVweQfMW6re6R1ZQCLPXiqOEF4mx57+8nUkCVEzbatdhGQWKcAv
L0E6ySNR93NqGDG667hZP/LetPtClhKK766/utXaeqAdQwMOCMyq+k72TPK3WYqL
7VsvLJPPSmaDa3rrHUoPDswuTWx1zgCVckNiet++c+s0EGg12GzZQvUsrJpXZuya
jgSx3wrMNrPAuolcJXAM81p+1dvrGuzPC3ZicvIe3fEXUDfBRfbSHgQjlLswVnkj
tF5CHZpDyIFP3xdox9JdDjJDR/iliYRoWUfdSa5/Cr2mHB8p4/Nf2w7LASRSybqO
E5tbhF/zqJl3Te+rrgx5qZEsBcoM/c70mhkfVS/KapOb6GZEpimgrvT7+omFAbYN
FDmBufU/EWEKwhL6NQu5wo2F0tIxoB3a794GUHk4gyCMvD7QTdT3CuPH1M+puUQ5
XwbeaehK3BBppBNATp7Q3Q3617XWOyOsoomMyvPSRp6LrGjp/PLcqqyzghYabyy8
maLEplGSdgt6h+DuVxAhz91m/+z537GNtyER2JegenORtQcg8do8JA97yRO4VIWS
LDtm+HTyAGwcNcFoJc8BfRMBnBGhwKBGpCed0Q6GG8CCgLbp3o5KCwAJmxLRBmHl
k3qWfAf4i/2KJIEet70xMnzFM3kueEMvpW81ZvjScwRTK15FImHJ26DT+gpxEId1
uPiHC4LUOLbIlzhhGljRlu2j4Rx6rbeszCKWXdm8eTSzcbUe7QmvvD+nrsnWsw6k
NzZxJ08l2bw0R6vTx10sCW65QqqrdsUoGwWs/Q9uLvIpLLpmE8eEUoYpGyMHZbqM
b1TaHRe1KPkcMUCXZoGAffEqQnDWmF0UnfNtDfw4Us7FAjdPqmvWoIDegCZSg6Ml
XIq4LPAsLzJPtdfAdSFbxby92z+GqnH/UhP7K80VBoaUqNoVBFx+bz2XVsCfZ26O
tmPI94df/lYn7PU5HjyvjEQY7HmY4ktIgOEvTFq5TlrjSzWhYK56qrQ8Wnyoh5dq
c8e91ZJFqacdAJt5lTR77c5byHfdR2Up/ki3mP5r3m4wNmSDuIvBNILU0pRwJ5i3
irMmGI8bzTa1e7F69lR/siTmIec8YT1ogY23hhHM5ytPR3EwAlWgKxJqHOyAY4qy
7mVVRpibVQ+LeabZia7QE1LItA6vJWiCiPpmgNYLxAPvAqOKrriabIVT3+nAiIaY
jdEXYjpHOlKCxyCpgKEv6NyLVxYRepzEFMdrLj+cbyGq4Mm7+WyrfZY+ZxZv8DjE
2+xAQmmBxTVmaiowowy6mWKo4G7m3PN+JM3GiH0zPn+HpZ7Yj5pFOar2BP4geUBu
BHirgS9yONoI5FgScuPrKbVVBcllbRG1Yu4l8VKSFdI19HxWVIbUHzSFD2tyKupA
4dEzraD0hgHiZFmyR8Azvc9rSyKiKYh6S653g+cC1Oj4RrDlxrGlMz1vU2fR252Y
UTogHPBn1SXkmmvRQ3UGi6wtb6mC+RZLke0ZlvWGloSnrrzRuKo6HPzoTZi37KCy
WJXp0YnwMOX0eJ+z/op5pVA7I70tTFD0FeqGnhB+wAR+7EgQWVL3QYC6+vRBldtU
BrmotUJDA3AP+RzHZ+oQb2xBUAZkJD1Vd4fHx+xovucvKxwoLamAYnO434qYXp5q
jpomtaCrhCzuIan+HB1iSwIQ3B9acPxyxsB4LXCN10vLabxz9QV4AqxE/aoGA8Ea
pKA5FUCXtKT/N3JP4/iIYysr9Hs41tgxKtZ9RUg5t06XLWmgpogaRHedzg/nml5X
vWzHnFC4KXB0LgMbGQFqVDDLaEGWZ+ecGsDLVZdmXqYD0ecVHp0HAzfbKWkvG0Bt
8dkJtzY3qUcN4YZGRWaK7D7k5f/Syy99qLnGMAzE6jlkDJ7xLolYTLY0RcGIFyw0
8K9k568J2Mlfq3GmvOeqwBx8RRzppjPIht553wQ4eMqt9m2fQeN2aqlcTOaZVFQJ
no0k2HT9ZL777AeUTH0F2kIzJPTP6RiFBsZhu+gIVrHtGtYXi7E/pTkBaX73UjqN
KNcp4TuJVEWgDxIrWNu/i9qHBD6bKtq3Canqv9MZZPe/UPmjgsL213OLfhKfyY3y
frmx7qc7LPsGJzxlma/xXhu6ESTRAG0k9X1jeGBFU5JcRL3bXVw3DDb0g0g+3GGu
9BP9raj/Dm5ipo2/sRHwI+jJ6I8cbtW/iew2nB/9wm6/5yKFjyaapdqJeRkLETyi
BKWUKdT2D4mluS34YFjj6CshkGVisKg8kW91A05kuQuvQnmGuFEyNN5NdEouteEx
srQbCx/D9VDOIWXvF2Z21gvVCctwiRtKV9wrZLMNP/Na1/cv+yd1LZXLvUS9zRvI
1exc8oCdskbq1Bn9cA2R1bQYxigao9p61zJxXjR11uoGpGzJhU+sDZTp/y48QZPe
ivCT7AAwrhSw/3n5JkHRihWcK1nYwWcRIuGrFSJHPVrbZSibUGWemlBPO0i02Kha
N1ViT1zPOaqZxk/BDQHjsLrDPsrE3bf88ynbheSi8lRtpD1Y+rnJH9vDkH2E+X5C
4qwo6cLOxoOurD3RLTl5n/SqBD+WU2gr9iuAXB8YQtuibGnVPpl6a0GEtU/1qCil
+KBn19Xw04IqS1KkUkHlyDHBd6POQrBKYRY27tBHh6WN/sWAhYJgu6mW2Wolk/y3
pRJyePoqooKxhqUlgXFbv+zA+Zl8rIcxPR3e0QBBBsOJfWpSTNOyUSnNbgOt/IPJ
PifrrIDAG6TonfbhUGkKiltoXsGQO5dtWrdqN9CclQIi92s/Tv92+8wpz6HxlgW/
ThMFt+kGY+urWH0AWS7UJ8JL1AP967pES5Fmhe/s6+I1wDmhMI58UDIOFWZAPCUC
GNhp90jEvar4i5V4LJcgdRqsaYVfOoB6wwWQwM2FjbVTLf0TkFaBqScKJccFjFDR
tgGCd+Gx5cn+W6EbmchdDP8uxpv00m+nWiNRwAyp4vKtvuZd4J1ow3snDvFqHR1f
h8GZAx9qwdOF1oH9633qUf7omE25WhjUOemdoI2kHqPiBOrtDYKNdGI+ls6KiQtC
IdNrSAhTZ6nsjVfrmMiYmUg73QOeUteiToen3peCfpwoMuWkyzSB622xNytqDqR+
Uk38FljQWALhLSKaWASRZ4nWyNwiy0v9nUJiO7lGpv8spzmi5KeVW0eWfM+Q16Wb
P5boaZfP6BlmMNjs1802kqwwDnbw+koTwLWsaFy0t6k8irvsMRELwWS/XqIuwj88
9N29JnSNYFiS2/3KOvKRr6ShNK4EVKQZIJ25IVeiCqaQ+C9T2F2Snjy4REqdX2rC
nbDwPh+5GzGeOTVoc+zYOTZwuqLw9ykdthSzAUTo+XK89HlNbgq0Hxfr7ydB1VEh
K+GK9ecPFsLfCB42JGs6U6cFuXVa0wu6ZGet340hF/Efxgfdsv1iIymryJfIhZrY
i/KnKeHi6SiiBvKb5WtxQrnMqFMvLgBmrfeqGk9rdXeDy6vqBY3zax6E9YzwmWLe
w7eexMA5A61tyIH+Aqq/d6ykg4T3FKCcx5fhyt+4DWrc0HnRtG/TqBh4fEBhxzW3
Yw4XPErdecpWihtcNhUK4zn5Aum+m/j+Y3Pu7Q500R93uXuykhiZANOqGjW7t+oQ
bFxooREccBoGZ93tT02KXPgERQzxYXJxlJRj0Ep9kdSnhlkmPRN3DPivci2D06cY
Qmm0tXO16+8Y7swB8EqZu+dCbeVoiiOULYBEC9V+WNoUrmj+RYsV/lW4n7uerq4i
6FkqsuYahLG2bdEKNHp+4OJvWKvccvmi+uoCwOGxyNl2VKW2snegZpEBtB4Nvg21
46ZiSXzx3jH+EyndF/DvJlbJk9/msnxHow2I9h2HaAOs8fZfMl6+LtoJAmXLcATc
Nw5U4UbYne+EYGp3SlUBQl9M5Avfj0sl5OHZfL52RcCtSc1VpMHxG0Npv314v3L7
VUGry/1pMnf8jdlIG97R+N5CFvuAFQAdf71sVDmo6bozq88Ix7F8jiwn4i0WV44h
bjwG4dkoXF7gyd3FRX3z/UHZhDhYO9iv38bf3EITuvC/cozg+geDPXwKFrt+qUXY
keBZlMS5DMkadAQBJWHuFttg+JDT39RRKdoXeI7VGm3VrLQtVDlMSMrVva+7ahxF
8JX1iaDWKtg5AVrxSm1esYGi2N+WdU0Sj+4MFR8A8l7CBZQz1NY+/uixZ9OMUOgU
dXpHCYyp7bXtRv52ce0NWVJ9JA7/JJkqQiYy/9XDPU0JbQNZHc05afnsqkwXlWH5
yoZ1SHgG/atXDjPEyaFcaAPR3v9/WnsXEye6dC3F0+7K2ar7GBaO2F5tMRLY5CzD
JC8Tjfm48KiyfTIHmyWxvVLY3BZhFaJOsA/JNznLH3ifknD1fGZh7ev/+3dPwyZu
aJc1eYgTsXb4urYDAPhMQn1poHptY0KRY6O6E6vudZM7riSuv+QWuAVIm/k1IEUr
88v3XPjSzcp/9OxVYNkEYMWL3PYSE0Uc0RtNGRy9XrdBBaEZcVhtULjiMcSPlE7z
xHj0wE+PMFjNLGxLX4j6Zof6lR+egzyacOpMyYaBNA2ReT9ipPOjhEbZ63z1AZ6W
ZkCPtQ7oZOnRAOYcYVoXMRApFwxB39Z+/rvvZgqWXCjDxU3Pp56xxIiglgI86I/b
0nAloE5u8deDsRslsPRw8nJDFm0haX2tR+zTesXc9a98LstNgv+paT5+ixtLBV0U
9rqgUj031DttvQWIVBfhSxNmf2jWH8By02tKdi9yQtcIsr2CuuK2VEg7bW+C0glU
NlJjmxvEcJz1YPAc9Gtvy0Q6jxGa+h/6PHKxxiTag/N3LPM2EpyvKFOGS4nAopRO
GvrIWm6FAWt3rYQzXXyNm8vjc8tGDrNFzCZpEqMsroT+IhI2U7YnNX0Ide3oQzDx
4NcT66TULtm9W7GBRGwxOkgP1FtXf7u76KpGLxdgwLgXJJuPfThzDZV0P2qttdY6
7MWBOP3hw32/ZNRXENVmwOIp/iR8OfSK5sfaQK/ZHVUHrpNpmb6Wn3dIeUexdF5J
NT2I4RNHPvGgHNrrkLIBGkx6s2MLL73fzq00G6mNqSDuBy7glpIIsT7ssDLf1BY1
mO582kCb+WVR0DOhsOFKs6Z92WFvAkqMJrsh2s76fUyb2BtCzSJNK+xqMpLBIvJf
qst6Z2r39guqofIpe0swzToja3T2GpapKbCUIn9DivVpQXN4ihPharYtVuiRvMyw
q6etw+jA4MoJmY/VjPLMNtwS7w3s+YrW0dtk8fe25EoDiW1/3dy2G6G84OVSPMSx
2oSW4gLoik6uVtjS3I2oCPtSlJz+lLQr7NyNoC/h2Tdijg07lNbPBefds18nrNJM
YzGKVIdDbWJj/OURvvFxcvqRsWlr/vEbKUco9y+RsuUPov9BveI6LIhultHQ6ACB
5Wh0BK6Vpk81HwUXgO4Ea0zjzRge9NnWx0QGLvxaDXwK78arflXmCLXHUYVvMMU7
LX1BJyYj3P4P92P5wmemdJVN0FUj6LYpScZ89ZRas++bqEKL8H7OriC2w6O1iD0R
yPqGLpWvCDYAeXYlmZNhrvMMKFTqCuFjZWmjKb8kwFwd6EZ6/AE64mqVAx4TOEU8
aJGdNeZlQDEKCMMSUWxRlHf5d05gTg5QuOsxBNauz1YAqS0SIppoUoSZTKqdYKz8
FcHbyi8iP6Bk0/9nKIQ50gN6+O4MKq8j/4r++hL/7n+6tKcj7ITVKwezTXQavARS
sFQbTOa6paolXd85FhV1ugChhjVht7LKkebthy7kL2hqDn/bgJbmK52h3bAp1HZR
uVxAFOa25HOVKTexUQr7IR/xDZD8V0X2onF38jwEDlmzYSjf1HA53T+2cPPol2QW
x5HgD8EOWspN7xzQMzdG//XpEN7PjN1LGx1OlWr2yOiiZFdxWV9CGGY+nINAYGPC
ZulE8dTySYHU8+uCsCY1LMa6pAIKuJg2qEbjD1x7EDzD5kg0raR94lL4LmaFxz6E
nC+Yy4sVBuptIKbp+8MnrNUM9dgd8T+0po07xBJJOmkp3dD7d7aQL0PTuT7gmP3H
l9CFDlUpovajeVip/nURMesLLVLwXKD7YL9e0z3qcshCQvLSMVa4aLGhFIwr58sO
sUNTY+Lt2vaD+KJqlSoOLT+1cQOBFPx9B0xaZMGn6+hMobv0BlsrHYS/jhqaxgWZ
CfaS9t+XxO65/964aA2nsZB/vJ6rGAxL2Uay1PaYj0QM9mCHpv0wqeVfS5x7Quby
GUM1P4dX0tQNh3HQyb6CCd37PH9jNvB7PCO0IraIAghoQBlKGylCO6IRzRPAuXXx
uSM5SSbSeKX6zboO2ynPOhhjldZzDgkhggPtCt106yORf309iPdllwmgDFb4KB8p
jR3HskZKIJ2UKA1j4jWbtvTP7WLeJPscszatcDQP12Zlg1l8HM3Wqymchl4qFhIz
zavbhOXCLdHx/IGeNx44PO8Tq8H5/8ApVUTY9pVlNjTvT41L9h5bMC9b4b7RsiCb
uLHZj9oc7zRMzn7pWYeGs+9RdYJwTJIba2PqUsu/HXsqvBBMCoVrlTUsWrhPwrnW
Stf4BtQHQybJi7Zu7LLjy24/nyn9+Cq94uQxQph7RyS3jfo72t1Oxu9o+Q/iTPXZ
tZlZBmztlXYf4grqGdrUtgCXf3FiOBIswE1w0fjT65ITbbAcXmAVfAefaeVUt5H3
D1S0cMjEMpk+q79I/VO8gFfhGknWfRnyYnfadMdsQPX1/XZyp2GJFceSrVlH6lZa
x8w7mP6cP7Juwi166quVp4cOzy2yEwM+OgWiPmUEGrdslD1KPlvlj/DXyjJzt+iG
QzJdpAhJ5O+YodrjiYiUiv7WmX+tVli9QAY9dj0A4fqzWqtmWAEH9fEveL4Nw0fJ
XUVISIpv2sVdVRwUNnWE7M7olVfj8nAFYJvgdC69ytncB4m394H2fDDA5Dq+gWxt
HO6dkC5REJQNoBMm2Npkot/G6m8q/SzBQnFIJwEu9rCyMUzK4tY1iremJbiF30/+
HPBvuE5l8EsGuk0CtiTjH3a9PA4mPCrxSa4glk2iwnqMExnL3AcDpdHvnnr98N0M
jH5hnhc2sLNzY8YyYpugpxjyWQpay+90PHi3sndm4raAmdQpk74/yF24M3HHWXiD
0UWiOq1QR+L61tIsq3Wr8t4meaU7TGVJwblTJi8jUe12L4Zt/luokC/gLmpjMu29
mdqX8QTZcUYY9VWhT1aFR3i2/VxeCGziYUn4YG7myPqUmxIHy4RFXokwkY5hU43B
XP1BljDb6qu/IleTQnzWYWrsOpzbVbWtVqY0UiTqRhfg6P7wJbxYtPYX2fximjXD
gMBqYGfdxvw+CDixlV6TBsAAN0tpjWPa0NbJpGundYt0Bkxr7LU/rP67WNq68hRn
VtEAn70/AF3TnxR25MnRd7NhZjX2VsJ5Gs8dQ2Jd2axHzqw29gE0TcrP+oA/cchd
7wUj7yG2tx2M9ZmrQ7LWEX/6xDUNxC5CF9rYuGB2l26R5JV3xwY/8RUJz6Ft1wMj
2AOisKT5JZaZDSYt9h06Aoclz2kc++5GYd047ZkPvOKNFAROk2Hn+EIGIWQjvU9J
ctlmKf3NmTJDuVtqHzuxfeZNoLglFjVmgGkisZiBFRSVevDYg3ccRZ7OKEb3C2vS
B5cGChI7SVqVRDSuElzp4OusOXEx7HLse4pSLOP187+2n3gUlzUOdr6zWjuC8AkQ
FEHOcfZlr12lNrQsMieT/GvzMU3bcBqb4NfzngKdQzUQOxvoabpbRWdJrSspJgSJ
nNuZ0LdnMvZtwt189HyZ9SKlFgj2cXsndEgdHR+RKVUjM1fzEvZhUTnG2LhQxVa8
+smKCRT2118ApdZCQhkMYn6W3j0MhF1hwg9HOxtXqLsWHsoCqWKkvOnhK8v8OQ4j
5Td2KrCwAenlLkf2McpSg4kBxK8cDSnThzizVyoOekASGr08SU4tidtA+BX5t/iC
c5PNiJ16dqnEY+CN4liZDvjuqNELOCeKyZ4fWqSXeFvil4gKFSTjKhGHrhf9OICk
b4ukt0xFtKv6n7OC5mN/Vgf2OCoOZkNKXlLNMU1gPDzo2WgMKHpgVEFtLHSy0/J7
ch0sOBWmmXZdXCDTZm2HaEpHxNTeISFKgZ+93dg9hYWXEiezrGJWPA6vs9jIjxqn
xrzjg2IE4auVaIdYLyVS34UqCTpWQXTii0h5ZNjJVW39TR3NEP/R8FI+4iNhdNpy
fGftsfPP/pll+OGMI8zOzy62wj+Fsd7suSnSkc3GY9PBl8nO/h1i98NnY/JEDNxr
RIn9X/Bu2gF5Mu5hm4TILtjrTbewDUbvd4+RHf3V4j9+sIIoDMQi/VIq9k1ZWarb
6HtxOfHRuK/gllosBx0rnN2ZbDQ7X9iPwh1mjEWY5/dg35rLCf2W494CYy2Fiogw
sr7FQTBSuNyqUiLd4WYaM61J9SllFGkqAOxUVTsKIiZywW5Qb5fEVEIp9hjhe8St
9RjjarMplbKBjx5X7DyGMuuLHUrZkfRSPyiGRYY8qQ223oZOJC+c2/gB6FLrhYiX
cgIINDFHwxATNm7h5cqnrnGsG1+LXI2DG6aLBSELqnzDFzLWk0JYWtir4wGb+DBv
fstcHq7k1e0VhkbMoCQ11HqHi71bJ+XRKSMAw3bOTCi7QX5KfmL42EEmwVdauTi1
jftm8o6lKQnBLXG0R6hta7tk+kTNk5mIahg9xZir9jdB+48nuH7m/P36Zo/vgLIX
sT+RBgJNDsCCiPjBKMizFYpXrBtTN0AuCwJp8DAJSy154WRcp4ah2kgYlJvqjM3Q
s3keJ0XuVDfpoJFnrE4J8DVneTWsejacUZWAe/0nHkRMHCHsXdukO7D/hzPYPSxG
hCt0+0HgLe9JwlLn1zAcWtIIYSPorrdA7+8/7kEKtH9cZQEwnRiBXsZRNICFVLQd
U+CcbgBqE/QUuOYkUQVYUTdPdGzBwp7pBH6EbrGDbiQg2FtX2D/GbP6FW9It/NpS
huMh3r2AGjzb1hHtof8GlnhWgMyKvCyoWOvHFTvY3WcqWWHM8Dhsut4CoV1aO2rR
wsK+Fok93l4fvFns7I58r/yNvOjEIn8wqRoXVXapW+jNB1DLxJnr30KX8Jy9L7x2
M5RU1BEgc49wp76pVS5S6FgRHwaCebqRc6gln/yiSGSTGZvuZjb3qTuvtfeyVdzR
38P965wnlCR4IYVUnNPMv+Zw6AScA+4fSc3vRxUAtIWIscJAXNdSOYpj3GuT2V7r
YE+4bv2MjJtVQH+SwgmsNiqnv+FMeQjK/kzR25tBwTH4QaFNMHYgfrz3OlucCOrX
BKxh5Gl0Gv/5WBOou0Qfsp7Vc6fi2bl0KURywLsGbNB7xz+Nd52aAsV/62qNeVCJ
T+VsBHqJx0pL+qK++r8SZtoMDgFwyl4atay0ASpgy48wdL3WgosJhHm6s7ji+sMl
wgQaiLBHu8zEDYIE4yR5z+q2kyS/59B7xBQ3edn0vY2sOi2cu6Ct6dp3NpC8TmVF
h6FxjHOzxwIAmYoSJz0DjmEF3yI88WqI8uLWkf9lbLeqN5ldAuFbSiO6vN4WsI0P
BQg6pRmZDxo/OGJh2+PB+voI5GRuMhcWrkvOVJ2mJbs16LV5Xcr0IF10CHKm7/iW
Ev3boapjYZxyqakFExgNxgSoBuAl2hcfR/29LHbpcEsrpwUzfKXRKBex9+oRAcdj
5fIg7+TJHy1Gwbu0Xg49XmcbR9CrnL+J6B8Fe8D2/KD0t2JGtXGwlbRrPKb01MTc
Da4T/Yat0MUce2UeW9vz7ndFOm7Rr2wMPM97D117kZwvpw7/QF/fqFYymf2ahSoC
Ywbv3Ibm/x9wjzpgw9DohgUh5afst4PK6j22Zuacv+q7JZzqWjxXqrNryq7aZfeP
gsLYPXftmYD72SP76MvCnFw8DNpcpD8EPYVYIyBnh5xq8sDKdRZ7cFdmBhBRnEgg
YODvlwts092MqfUIDtxm8KWj4ZmCcmuOTBOY8SHM3CMrWxgX6QMPP3n/a3eBnzvz
OMkTc1bx7Qq6zlqIg2HN4a9QFUcA76glZcZPguRPO6T2rR2VJhZ/K+Kw3UZMdCr5
AYfjQz1NS8uAmLkKMH73BhfDZAQi3qpo+jEBUoPcssW+ZLfuXArW4P9OuLXvhBB3
slAUfjtKpZUm+hXh826naWDJA6NEQeyqRjaKWzZgmcQtUK8vcJL1h3/glfy+YwIF
tJgHhmXC6eG0Iy8UynZ4trkbrRuppvjLAWevVyFdqzKmU27q3qNymS26UY+Rd422
er2dWRAAD5bfupsaD5eQliBQNLwvUSdXv66IJ8qJlyx91z8MTvKDNy2IDDc1KpSW
KafMg7y28j+Bmg+ToEWfNMswwRot1K/XounlEc1TnDTXHGByONruQIvnjzS/T3MK
2E27//nTKCMpulFEhkur7uYITVXsUBIXBGOpXC6xrfXNcg+zYNnkcED0BQ/jCe0N
7009YGO2OeTLOF0t4BuPk27iOgZDZ0KXtShbF5VBRrfecwGzkpdRiuuAheb8RQv0
w0WShNzp6xGUkKhbkRRCa8CkY2XQqEdWwti+27cIO4LF9pmKxeC8/DmNY4MY9L6X
OBkEIcx4RWa9rSHHln/xP6OvLQmZDE1WI+NfapATd8qfv7Ht6+wybmWuJS3EIXEj
ira4F3MciKI8ZgqoHeSgGEA3mvGEWBxJzs5kPI3cA8Kk7HWX4kHT5DY8DjSkleOE
/jW82mIZMYzX/l8nvIjhBYgy2zEaUeaSx5JoVTSuRTzcsBRZKUYCHkdSYbNf0v8g
3nWAXn71f/j/VOnM2K85cOkUDbSQHiyE2eXNDxjioQfmLw8n6aIkdz7nnaBaqBJO
SY9ePXyy91ANqarsKZD/ySbQXo8rXUzpoXU+cGIQ3Lfo3Z0nkGWo5Bvej3yCm+dr
YZfG8Bm8Uxr8BfaDpiY2J4guQmycVrycHbpLnl5mAI5NwdejxLXUMSFxDbpiZx08
6BSm9sYUtWynmece/OpHgATo6tWRnZNJrmDzjnGDA+hzv2hEUiB3T99rtCU/ilfF
KmzcJwkcKS336VNl2wXTFqV5Rqr+HhBcWboojFJRXkhrExou9TmDQbDX6gPPYXJ1
NjdgZSiYLqYlZGMm54786rL7/WKk0MwnebWmtNLNzGYcStnWHuJIQbxA4UKeL4VZ
yXrHtXC5pKLLkH091rZdzOlO00s3hNdnIJDFVasEFZWVzsHIcxLlv8l33cR1flBt
oECqFT4LkxGfLjowagUYi1O6KhpCL+c8ddVN5B2NnA6b3Pz1TpvHdQSVkdHM8x5C
h12IjNqrLMFxv5SzmNnHrJ9NsWcJijzUyjnN39pdHtEyIM3/R7WPAK2L4J0pr9yy
95c2WDQYxl/WX0v2eZeAxB03s14CTMzU/I1CQ+WVdTiQxbvumNYKBxwTn/OB5Vkn
GZymOhevHMiBzRyPg8zx1vBljK47BTumn7qNO4hTsaHmqzOE9Fq8H4Er5VX1ajoH
ofvO2iAj91QyBzM/ZWBjofCY2i5sTZupnb2g69kQvyGc9xZSe4N91mgxajEO7zpQ
OTloenPRX7HVof4kXE1ii43DbAOEtxcsQsL8dI39dRfXnxysySeRgNBtQvz2PO1e
VExb5EJXgEeee95drmVXk9aAwfoTzbVcmMBXp8dr2PIU7frUmnZXBreZ2fCkVo8x
Ix4u5nWE5IoIG6wyDqnyZrZt83ziO4eIEjMeasRK6MDKCwfCXItlzSHoVlyAw5GO
uAbnBDMIv2VHNQ094lnbhZgOBrWBH5GRnj4fB7vyX7A4nIBh9sxdx0P4wmEXsY3M
t/m92nVG8xI5cTf5T2Ya48boHK+iseSrRRlJpPZhTzQv4IeWeDCSLmfTyyCcDbGx
fzf+hRFAqFrLwrKeQ1Brlp7hSbA+kEjduPXzNWuLGhk2mTPu+Zi0Wp5cyu0JiGOr
uzonttiTvLj2oQQWjgkI7ZKTdwjmZe1w8dSPZn6480VwAwTsCX7m2XhPuVSVgDvo
mzkal1IeA+pXucR9Ialnb0rvjE+AQR3JW0JZts46wKmCS/qWbq+upiZRUq5Snm0o
mh7PMKHOP+eeefI/xiXroupymB0Nn4kJBuno9xlnzb/JGzjJexgkUk+4HqBfKGuP
9KmdA8o82cX8MocnfM+KU3IlzfFPcyAtZMQqqgbA/QGz0xTyZSlpfy4nqvpjLfh4
/r/KUfuhf8AEEYMcVgy8/tWBsO1DFX9B0p/vkBszPC4BRc7b1dL+GAzgtYg+31lq
p9T8ctZ6s1FbtoWZHExFDGjTvoWAhATr+8IYcvqjh3LZcOo6WE3KRR+tfCc7eLdh
IFBASir/xi3eMbrYLWRMliAf06ZAzIuFTe8f/Iise9+d1SIfu00jJsTb8R8Pes7i
6eYYRe2N5PLqLrXgTged4roy2QpZAGvaJ5xxvdQ4xHQBlCR0ncQnx9hbbzf6tuTl
h0MoMGZDx9FtHCC0Nfj4BHEjCiuOwLJJob+nvvlZCf3vBohVpT7cdxtz8I2Dsilw
79npaKuFaOxsHh+T3bzAmVMdE+N37GLm9CxIHMBawi+u+e/Prn9aUHNoBBDBzsHm
qNVMEyM+ciGKteMSK91EdJHu3YKvIXv+CFrTA/gGimqH9pPt1Cbq8R619D0T2hNA
oJu2phLS6X7f/NbzGXHyMYWZcq/pTAgTVtSir5VWHJFmHr1tolGI7gacw5pQtavi
2efoimD++wgGDx4LM6G1dpukRUOmlpAOQdkcEunDHDPhh/erEFAkXbndKY/gTFa0
voMuOMGN8riloyGvDd9fhxUFgtbtyd0sjT0gekDXQPhNo7PRbWsoFCrH6dfYdrkI
Zl2iXVNUnZE7ivBlfn9/JY6m4B/u5iRCAdehKqIH3v5fxfQ7WiBStUIrwbvmD3O0
Oowo+iHGEVJX0t4UfFaCMjO6a0akDxgIGh2p/McNtb9gZ1juOqQ4oyqzyXVN8ynX
BhK8up2PQJh+1R7cIgiohmGelq5YwzleKucDC0fT9wflCUaRRQ+JxDIGLbnfrmqC
FJUannP162EFYmxs0w5lL3s1XLFYqArePKvDccsZiTHSETLi+rKvOwQbcCzhXxL+
VE6Tk+YPAY49axr4VHskF3q/KAScyb88OVsuMRJsiEjKzaR00Pq4ua6F1PMJYo9x
3iaY11oIDKZN/DZKOFjlVtV+auswKo5uJnO1hzHeLU/b7mvvS6Ss+ic1Y4anTrMa
VQebesyFeTz2aTamOKb9Qg36wLX9cWoOfVryl7NuqdvkUda3rarYkbreBLRYTqZc
NPz+T7Ll6JZuUW7z6xxqU6zyspRvBKubwHaGbcwdJ6aEm7Lz1H8TbzVKSiTNW4hs
VtrRAP4oEsI5BwkGxdUIw5dj7SfslIqiWl1Rgi6shPQS+yHuwByFuQq2bkf7vJ6G
W53Smz2qxjnGTUIDVBka5pOCIW0BewGxB5ao5jsnzCs4dJHcrd+qQVzgDPMpwP4A
FtzTFjlzh4/XTfjaEQzNiMgmS5/TK2opzYsWVrYpsEEv00mec64tHx7m+Y6yLSxC
E1gpk/Q+XviDeOCpXDla3DhTTGNDzsIY1uobOLuemDbSCBrH3AZ7MPeao8nWIEKe
dDwosO7qvFwGWQsyG5+Un4r2IcKR57b1xD8q1tu12UULVoy2qyzjYxUgm//YGkog
jL3MOcnwri8XWzL/KaitDyDXGg9vCX4t6aRpRs23okpISD3JiryKP3CbVqp/2N0h
Fp3ajPoI644pM85N7FxARDgskb1PbCP3v8ibt8UrF/adSQMJ5MZZZaP/2lA2UTJL
xMiacclkqC9bGyGtcYq3eyGNfahdeqvSDRJGS0mkUOcqkY8SsPIzS879CV5YmzmO
ux0SyhmWrVmQsuLopiMA4BG6tbieYQ+dvKXYloRDIVOyjVSMOxgD3Fv2eksl9IH5
XrRALeqUAtYauZHM1OOlXm72r053O6MYYywORFrlt/tMKvkQhy994JAkOeWzBo3m
fEk3ZCKomwaX/Yxyo/Cg04RwSbrSJbwt9HX6wECITREs3A7WNb8BAaiUpqrBA+Nv
YMecKU/xXomuwqAKvZAWr5J+BOTe+mA4amKIYPfRFJPUrAEosIFvCzxi4Xen5zcc
H8ilFpvPyQILS8OzOltQ8791lurH/uoE9iCofVmPhaL6MHQaU1482mS101UPLsYC
DxIIzrRlnTjqHmjV5j+miliqiBsewqQuAd7tLC6822iq+HtJ84d19YzpE8Uupllz
nuCiCK3rHBye77eRMnmQDCjdHPSWg/HFq+CEvXFPtTvyURPbdc8ssNOzVZgbjxfp
wpk3dNGKbfinniDGxtey38b8w2L8cF99v+sFuoRJUAsyN5I3hTRDl+4ibXJtyQko
nf+dxw2IKLIxAwXo17+T7pMKoobFE/wWIcQmGyNer5TAsEH+ME00YIxG3j3ObziH
gXDRaXWN2Ll+n/knOlXpQhW3TCZ+jKwTwNHala1LLCeN8v+ihVCPs5vrD1Eb04bX
ydZIVm68Cw5T9jo75CwuOUf/wgOJIvGrgp4hfA27qD1fNR8GgcbIJFNH0z+/Rnoy
EB6GnRLsuaL2L2jTEq6iWTkmEQOixDMhyeXsfrRlyfaQVqOsiR6Lfi2WeT3lkp3E
Wkdlk7Gihh4REFul6pkxr0wxOHa0bJfzbNT6sk8ujzpJQJmRat12MaLdaQ3/rvBC
x4gDh4cSCgyzfNAwUhhUyfcThEKOsWRFKgWidYszYa2BQJ55uC7D3D4fC5kEF8hb
rMO3fXQy9kAzPl3csL6mQkYL/spXj4vLfZjMAte0s1Zt5RljzB9fXCSKTZfL6dsh
OUplqTTqgsaElMZOqTU8cXSN/wg3qtbgBy+f+WyAJq39mczYD3qJT3gIsZmAOBV7
9PgQZjF0+GYIJIdAZoLWleRhIcodAPYaJzy9/AHX5Ayku7wQDFfC57YCmyAbEAKP
mp6QqkQYgkDbMKFJuFUSamWkd/aDnBpqC4+aWyfDP9aS7YusQhgdwLJg7jhZu/3t
TH6gEFeFfFVLkog3yWvkJNgw6vmJhaZzfh86TxRzXVxmyANn3pCu53sPyaoTS8aC
szJS1IhTC6H8UUDAWJdrQJYQULXCzrQeBG0bjSPxZ+il/NbjO1HFm9CuebPKNFUO
Z0NrT4DtnPfUvp4zO2hiXsdrw6nsq7FT13Vc+roasCZpip4rxHzUmfoZx512XjiU
6wdqbEgePVxJT5YhTeJGvHEs7pgAk7Tg1EyZaIGQU6mcPgUTrPLsuwZ4xzJwY3tZ
rn0VwgzpyL9ZO8ZI/Mzgcn6HdYyEpQD8jaOyCrLPh2i+/L/S/EKC+sbSNxJMTtD3
+IaDNdkrw7NgfNPIH+T3706Aa2hkoNSvbnnBI3vFZA1EecXya2pBHb7iqrzQ7m0m
58nZ1krhET0tQZlaSFHRJSwAelo6JYo/fgLg9ltYB91FUYxt6amc5TSpddQkBauY
ldFBJrWg/Nx7UnvIEMnAsfGfhJKkbHyqi9tcbUfaFDsCDRftoho9trd9c1o24Fe6
4FULOO6JgPYeZhfnPdh7grrYmBmozTs6yOHv6MWkXXZBwlyiRiS++voWeCkFErVs
rcVkJrdKyIX3HHhf7HLoQ+XDQAL4z5Yuh3fDD5aLnyb5KeHjqze1NXvSujWb8RQV
ifqUdl59jaDBCKrAhM9YnaXodyfvLG5hKBQd5IHISJjq4jQeRY5GlnnWvK0GFN3r
s0hEN3QAs+xE/d5tsBgDWc9eNpts0I4YB9YfC2OIg7C220+wwEeY0+putDBGhLyG
XFSeGBEB66r1krUMj39ZDaSbN6h3triMnQpJR7icvk+eXzjsTu7GGmrWOiLg7TTA
E8zTJVkZiwcwCjg14gwFSf+5pLJWaKxpQC34hCj/xw20Oe4ptiosNtO2VLnmzsi7
HpXLB/2Doqs1JWf8ARmp+FUfGS1UWo7HPVeVrCz22IflcnrnPDBpNDs7MAgv6VeH
E4nbWgeLh4Y6QsRYdoOQCXWP/zezPyOJskdqwNJJENGXRNyUfrgyVaaJwizhBk+E
KI+tF60Nc39z6kIydgkdGWYcKa+91aGgisUr2qJyUiTPqifXqPzUz6QKWoAnoT+p
l6BRZ8/zCZIWtfblVlDruhYatoH6h8iwyTgQtsF0hj8Dnh8fzF1trX5F31bhHdZ0
vBT+mzCpA7UQMRqvNItT4BuauJ3wt3DT+pNdSTE5CPmQuaxA0dJX4aemeHO6JdwN
lEMMBUY7wnwxj4cVeBXAziZZPQcUrea1eHBqiaZU4JM+Otzdm82UjGcYcSiRrIN7
60QhDLqwLHybo5boBD6PN/tnZTnGpMJWCUQTBWj2mfyEMTFH4DNIVmH4IINf2B/g
VaAvwQm5atSdNUATufbrmo9jqDxFiVNh6WaFiHWjlMvtmwFj3kUKXmc95PARwlME
EhPnUzsw0kMImpJT/6ObTb0Uu9lgDizKrDaRb9BpzamRF4RI7TuLCU/LxQ3YdgL7
VWJEzv2MkUv3VQl5jayb/L6g5+Ak4AqRPUL2hWzobIXqLqG7PhTUHhwbVwgDZVuv
4P8hxu0UsU6M/lwNeqJqHHdKGPZpIP92cOO2Igdwr9LJxBCx7MrgJjOiJyuA/QLs
Wj/R5fFCAHLuvvoF/WAiajc4m21XsSTENJ+y8kqIA0NB1RFlmvxc1z82vhA58isU
NRJKYkIp16T/OaN0F4xKXLq0jc7G71GceEv43jjE+PA2349Mx/Z+5yZF1ra0pISI
nnoXcwFx6rFr+4zLxjL9f9MDffWPqppmAqLABpNyqqRadvcc62t/4nfmAYanNP8X
s35n8azoh9Lg7C6DqG75IGE95ukHfF78KjQCX3UjiJ/0dlckM78/lSBPSt9Uc2jC
rqwSEHFWPA4J+yGsB0mte+D5RDJBAR1LDSRu59+qruy/+/xNh2QNsXZYMvLVzRek
ZoMnJPLUxQlnKLMaECZuyUx56hbeW/RCEgfZnZe04O2d7EoyYCefIYWHxiQxhlo2
pptguADYKdRqQC9K/d6hVZsYV1pYzU+FqzvIHZUlUi9Fi8qzIktmocg+EV+PDYc6
ho6/YSuM/DvvVDd8lzzqp8s+62vOZAYDT68Zlw2cVO5WDSfF84q00Hdi8QNDvFe+
YhZzGcHGqGvzwE9ZFpZCrAS4nqsRZC5dL1sZSLFNgV6n2kowUGsrLUmgMLtgaYo0
DdTwTpKJjvcn7CvPHsZGmf2m5VdUGYmA0CsJA0wFIYYh6QWdfcAhG2q9UY2g366z
ZzuOa7M3lAtdLGyFohqjMcQUBH7hKt+2ewuAD1szQF9zmo8S3ItX6dW89ydbLoF0
nEyAxPq6pi12zMm3nRw8U1GHZEs1oUStcZ0tzyIoRdLPKxz604ha599pIYmPhjpa
g5h2tAVGn6TInH1IxA6Ruw3IHZzJ5MjBTAWZmV0sWZK7KOGsAovg2wq7z6oWqjRD
0AjWE7ArEe/Ym+fpyHzL/VZpBONnBM7nrm22+4guIiIx3i+9EPR/OulNbq+yZDQ8
Hksf4I1IP5/mQW4Dx1/5yjsKVnvjPw6tYRpweHwX9G8OuIY9fzKcOXlLWCeiaTLX
g33ZanPPUOyl4pAxnDDROCSbN1ECQlvQn/dK0+Qj+rKYuHNCQfXzYG59T6mjPqqX
aJ7it0/R911gflCUy+NPbEPs3P31FV4MBdNgkeHf6VuiN3QtAuPVx592mAbmeJON
WlbmTANYsE6BU9o/UtDwduTv39EQBUnfGEpjZ1NxkYfQ96QqknO2ONg4mel340/a
IT7o+oH/bN1zp9MkY/WnRF3Yk8sYRorieznEWyyXrhzI13GQH8ElQuWP9wXVviig
/GwVPUM+YkZKFB8D8UE171LNxw2rGTW0rxs6Pm+oI7QuGHdCwUIn299m9renBBYB
hFrAgAf2iaeK6FL4ZWJ3R4s0iyZg8ZhxnTVkimICMHxy7rdD1UW/5KBvUySigxjU
DwmzIkUfpf2vxTeFNhYmwQn7PFcBML4B7ag4/brGutxCzlnfeZKnMCoYCxVOz38Z
Jn8m0/u+RvB8wYexV4RP9RhpVJ0H1Df4X5F9l6B/17ZA0lZdKaHCwclqLSWc+iFd
9HtaBUvPbkP0KKGo30wki3cgNfo8F1uaQQWlbuRZa5YVpCxyr7uJdHR151qnEOsy
pWuq6QJ+C6QzWmKnBeFuiYbMTPa00uABy7J4CMkScIGThjVlHYlmeh0XzKO2VoIF
YRyk8k4x1DmPxOGvQDKNL5mXgYKDjVaS2JiIQlwkEzbzKRkz6+LZByZCK4Qg4gdm
tQq5bL7fTvCuDjxRz4ftIfKefwW68SONCSE9mMJaM8bYEJGYFHDzcMpbNdBmLmJS
93AebBqNMihVT0W8J17Euv3b3ndYjwKQrIBETBJh06Ap4jy5W8fQVO9p1oxkjtYN
/ZFC1DPUHhX7AH3K+Kx5cSV0MGjFPs2bvH+CkJovvZK9hOshrq04KseaP2ZKTcN+
FIuq1rdU7hLkSrs7cPcs1kHb23xqciUC43kE2Rx9303lCQIedbJHi26NH4RnF3zm
PM5hJw5Rd3OWCuEFF//nECE8dr+FXRDbNsttGBS8BsOVBmrGkFwZkpDqk9Kqtmh0
4xXOI2Yvs8uiZNzZlMwc/2tSrTGc6NnGg46Ytec/62HORE0/TgHzxDGCcG0OvcTW
5vk9JvsdW80Rew2bXxhTz35LalPpk8KOHtxcHHPNnGlH1761lAxXouekBul8QHH2
aDHsYuK8b5NYHLNF48KPCX81ntoDX7QWSQpPUD+Qz+L2v1YSPZTGHGz0TUkdpkTJ
1L8wabUb3iGANxGQLDi7tXm50azkg3Ky+T0vWZLvBSoKtTHhD7vOmV+wSGCyVv3r
rXXpFc4zJwYSonEO1jt0awotLHzWhpiiJVINDBjSoYMMLudC6QbJbG4zd+dXXWoy
F4Xvc/X2o8+N0SIMeryb3hnwOvU87J1W82ZKOJJkggptibbsrPX+WRM3kwssT26q
PhI+j0pfejUvf8qsFfdwnoCCojdrv+cioTdnI/cUfF5Pb14nmF3xBjyhLCkTfa13
30mzDbGtNNtQRfTC5agBHuMnsHd0Mah4oWn+2oMgrdVBktl1idFktyBUEZM9mJsE
VRGGPlezp2StW5+q1aheSuodGF2Lxz5G0N77vppAnfcRJAswVcb/JXw2u47WPOpF
R7WZdRLKGaCnb6DmVVl9pMt0qetPpyXrs9Usu51hLuRFFjxrSjHok3Pq8pWQHrUI
u7fvnjatwtXhfnRttIeMhhc5cxdMKfDnjfHWB/HGnx0eQjwHrMMii3+z3yiNKBC0
uW1rYY9muF9eCMtgZaQM3h4MUljfdreuSIyDiJkgMYv9xJeFIWjcN/1QcXlNuNJb
6Ztj+iiWc/wVSJzbt+VYeg/1g3LfnTg/lXl5yJqmlntyD0euabADcGoRsuUwZyik
3SQ/3ol695VlQ0d8frC0mJ8CeZuW6nhsA/9eJSgEte9eODwFA1jiLigdlkANclEM
E87YPjuo1hZGFZAG/0NQSHGULt8V2Mpm5Pw9W5UTQLwUytTBhi+ZmHQWEgrvtD6T
2rrXwP2d3PoUSXzs9Cd5vqfyNvO5U+uWVY5xtAm5NBJ2TZyvFEAUmgEcofq+csZM
AacQX1HcopatVziunM3l0dfJUF/5BqutIh7ISwvtciYxPNfvg+mwDNCd5+7D5aKP
s9OH6ZJBTV5v46SoKHBbtEQqbPLe3SOQrxSynPUqoA8br3Izw0aoh90MtvoTIeZW
lUiAbSfaCQb9jMcJ+mCk5gmlzS0Y2ol2mCBMiax4vaZVr78LGCMmY+jtEokQHb2N
fIGfoTnW5Uxnss+MdTTK/Q0izmCuChbC+a6CO6AcghFaqKNfq3T2x5og7sQNF8i6
PRvQi7SM/WbViHLcgP/FzLaG4OleWy8XdrJUk3WTj8yAhrb/4uAv9+nlRxDjcaCw
+McxYGTLz5fgheM3B1m2V9kxVgDi+/C697PwMwqHag6Bz+YJn+x/O47O/wTUAb79
2NN4SDdu3RUHWvV6+WDFJ6lm8fgv2HEu0joSv5wF9WSgV+2CMNK6SfueG0rIdpYG
v+U9ArLfCzwQA8uW27VXCofjL5OgdJjRVI66AUP7oKcUP8YeOwmfw7ieTcXdagvU
NoStGUjDza/6kQDKYkL4vydZHIpU6BdiGa4+vzAaaxEP1ZSx2ZWUmx5Dp4x0YRLQ
hv9kq/t3vxT9g5IWZiy4+U4L+RcY1q6gALuSV5wXk3rQISsv+Fg3qx2wsTM0XrNa
E0SvYa+sETO1m5PpIHCd72H0Qd84kfp9WHE4B2al9u8nSNrxeNYFvBscPWL2P+is
oWvMn3BSphy6RCsJHAu3r2jeeE6JvjaAyaLSXAXsbRhkL1QoDMzLtV4mCB1Ydw/v
7T+o5SCmYz9S8L6hR66k3p3cZZduq9PIni/X+MZKaS92vgdW6rxtDWCGdVge5lbU
s2pave+mrmZZJhmXjBqjxH+lI5jzObAia/Fp6lL2PBVb0YDimWzUvWnrw8uJJK7B
vnK19fJ0ZWkk9aqZ/WbQjHeQM018kiIuqIgrI/OVWbaAC9kuNfQSdvF7uHcdWwok
Rjz+CUuW2nLbX8kn0XLzFgMgAy2KMxrxT2RNm1lMUXI+ZDNdcHskirbnueK2rVm/
zPSlJVp/qXrzhYBhCSMTdX1yRIosgzN/woByTwjR36WNGiQHrCnSYX5BqkvZPUfB
YCLWvg7cTai4VqK1F6PeDv/w8qnjCfMAxCcLrztuYQ2C859Un6Gd28XDasjmdG/7
Bb/ROVrH6DsJt9MNm2wLXmoBf9n5lJdbt7bX76cLeu8Mwc8yPuQcVDnnJKi/aLWw
ukaBkde3H2IOA9EHVWFYZiTLFoGUdPqhSTMJEOQb1s2jBNKv2a7YQvhbMv04nwK2
S/4Xzhc9JnAb880P5jmUT+UiVTDQT7514qHwOZVyaVawCbMb2MtuRIOWyGQqw2o5
c6EGkOcxqHI4q+GjtjQVI3zXDu7oR5n1GKDFZHqXRmFnKUWem3CTfsoqOhSUL3Jh
5nygJywYOGPOm0r0a42z9lwI9raEqfHaRym5u/4Xvzl1FKZZ56WqYeBrQuxXHejj
N4V/rbCgcVz3xHNHOiIAU943Q8zbIJXitGDii6Nmv62QlmoNTHmnPamtrJ5Q70Mk
eu5tsQ3vZ9S8Jss/a8Bua7MR0wDbP/HBkjBaLATsQpbRjgUZ6Q3QE1EsJu9oEjvV
u8yeHRAtOmJrOzqylWlLhCVGTjLS4k3uZsL3pD74DP3+AhQd6Phj/LwvyhRd2Xlq
uo1rc1EA74eRGN2Ee/1mr0J7FgGdArZPv1U2yo2+w0/NhGYpDLJn4OulTjb2aXvO
QynlDMZb2PQwiyQ0NLOBir64YDyVRZSBPc9a2OwWRUD8rXrEfWXVaKHK8iX0YoZ2
jtZGtI5e6mkGFx5yCFqvV4mscwv+0dU/6qD+0Lh2sC/3shV8pH+g+Jg1wiyc8DJB
M2AyG77SosP2Ges5BIHj4QnVxwbCmOxJcfWeUaBHzl1YAXgaekByU5enLri0fShZ
qKvPujgoRlkZbc6RvrFvtkjcnsC+iAyKpWaJMZuCOFaB1juOYCqn/0+4MwdiCQXA
YhF2nQqxNVCssewDlHf0QZCKz1F+8WvzVdRc/PoYFNTEKVnT75Kglj6kkV+9P12g
TbKLmHDj9wuW+dJRzyISKXiryrxCm+YHEcyIeE8WC8bBxKj56RoFy4QH/DkPqBjG
APqmtcsU+7WzGe4do2esHctSc1FfDI3pnUYbxFqQNqHKjj8ZtZ2IhB4/TL0wOxKI
m0wE+pYPeidodY8PM93c1cV6RPgDrViHB/FnGfjlAu092ipbabJ3rT+YQGX79aT5
Nu1Msl82eW735vyP0nPasWNFvxrtJ6b6VOJHJ+UEt9DXQ1+hQhOsO0Q4PJhuQhfR
ZvksqJgaFYWdy48Ses/Z2SFozsHMamtY2X/dHx9YIwaf2KrTf1HZ5wbSqvkg5TFY
q7b8acYMKLuuZi9UEuT8pEdsNQQvYA65l3i4FwZlTd7fIQcg4v/N2ONLcjbGH7Tf
763LXhQSVed/tDv3wXBEKpEduDrN+1Mxwr0LNzojqYJ0y33GGSwnRQA1EwDFHJsY
BKVEVrzuR7VjlrJ+A8iyFQT8rIZqjv7Tdl85GDpiyxYozePRTY04+6qwGWiqpHJN
uoxPR+ccDKnmFSJAfH46/4NzG36Pkt09itPAgld1eIdsqph+8P2DHhjektl2YcFv
KNFfbYVSK1EJ3SuJPucBgHFipUaC+vWJbbbTrh+1kKSar2tIJQWS/pag6cNNihHq
7m6xKHvt+DtRG+47FPY25ITkYPvUBBIyf5VcwGR5ENu3aQuJg1CTyiB4Vy1ISb5R
4JJVMeT9oSh2no7+w+eCG47lyEVCLEYt+OVrr3OnAQQSjHX6y2xRGicT88kHkqmZ
0ZpacTbrWvPbva4Zhpm8kCJkFMcVJsyLXDxT0364Fc/Gn8mDY+eREVxisymo7xJN
ZdP7beG1WGwtjeC2zTBuLwNGsFw5CLdW2Ch+RnulGjiKcO1aGzS/BuhppAGPdi17
fbmw9CJIxZXGU5nxmAr2uY8U3bPMWFUr32ZvzPVV/Ty9kl6x/Gt4vQzhxnqXEv3T
EB7W0DlVpA8Cz+s1aSDp1cN7y9hFdejKUOa4TcajqIl24/q+m1gorWtynlSpPLBS
snnRVJxv1ZWb+UJxcB3XjXvBI29v63TJv+E+7E5QuMAZ72sxBUUostiz0iwgIlrj
Okgv3vgPdGY29iqC0HFg16xclbV7YxLaBKPiK96LrlYSHKwWgU+dJCs5Nt1tFA4f
6QRmi6+79v/uJfz4TdnItnhVnxztU+0oDkLGd53kl1IJlKldOHVPOCR6hdI49mhV
+5olbmdIE76doSO6D5pzSjZI5VwgJGt65vCNXkVYqPwBT6SntHRAX9BO3ba+KHB+
mC8yb7lN/Ao2mtq3tt3AmiFCOh4aRo4pgpWNXnKQVIKK3eCCcAhcdYIFYW9Yb4Xb
/JGhKgHWd48Pjmt7Vo4wxsB2XIeQZ0rXLtKCN7dhp5DPd5RyDG5RAsBX9eMPbi4B
dUunFhPBknXi7XCYWa2BD0MOLmPkFFR5k18VBZo26Ar9mNEseIRvCLO7fTe3iyii
PIsn+MaNBGPIAkUFsPGXft4opqZn3lDVKRcbkVXYrCVxyspv7NbfrkeiCvJ2kRaB
7FB+yjgyep3ZIfnZGqdM5qv9NEk5mqTi4vzL0/XubtQ5GdQGWTT9IeCvABCiJ20d
2fJv+N9aCP3XnXhUW5mKQ1l8zZtSgnyaW3fJJU6qEt29ovIyQw5pe6KC/jvhA5/E
m24ANPIhs4vUfM7PFMe1c3ctng8UemNXcBPHwdWKIlAfpIkFHhrJxVVRdD9DOvkY
Ex13qmsrpSsBrbGeo4TI+jZ/I1N9dklq235rO8fa4jrBwI3SRr0E92lSEaoTobyo
Trc+YSq2+jXfWycT/0UKKd9jaz5Lh4FXaPGHt9Zy/YwEMH5NAyqt0Wn8QNYxkkb2
ZTcgbiYU6NKU/M93G4nso7igKHwnP5zinmWkAu/nD1+iHYGfdcb0aE2buKKjeQdr
mcxak3jY2eZhHm5rCeGAg14TQIiI8Dcyef9kpsZ+K8sC6573rED8ydLTASyxv2+i
haFR0LDZTmY7n3aOqYCOkdGvycg69X42aPxxhB0h7fIuRWR87xrziOvfYSVch4IN
2uQEF382dfk4ee2mqxgrEYxS6IizgM7ZmgrJV9V79bAAfFZ0nxrws8ufm0w22HEy
QB+DjkCIML513/gQsmx2SnL//0DvTU9QxvD4GgofvfKXhiOc4vBa17ZREPjMx2S+
sYHTjM5Sdvw3HUZyAnSDBgkw8I7Qjv2ipV7mbfo3GWb6c5TItbZ70drevFmFYWE2
1kVpoD8XqFfEux2eNV+Et0jga1PGhRfhvKiT3zUriXAqlWjKZxaOkCvJj6L7INid
VnO6flT+4xd61JDTtTn9WuPUM4V6lGVABGC7nBfJ2QaO8J27RpKkxwwzDpxH4UJl
Kuubuq97Fu/vPrnt6LkfZpDDONlTO5Am94nOcFm+NJjePZ8Cu7oLM90uuOEXxlzY
2PVj6gBiws9VJ10v6UOvnJHeAh+QC8E/tn4GuGH6SGO2BgBAo6N2Nokd33YqAl22
AxUJnt1XWuEQU+HN4veJm8VygdfflRnPpXenxMGQvBuf/q0wjnFenX/QQh+qLcqJ
0HEOtUt23lEEJCqgtMTELd2YKRYFmSNZX+lt83Ble2SqZhqhCartepd0Js5/s1t+
iLcrDcsg92fOkr6mK+n68sXbntF4f5Bs17WwDf1PrXfSL4rPs0mXfOxHtQI70gv5
JpjwYklITueE1GO0ISrjKhO7jBRgbGXhWlfxRXw72CdY64tmbqKNyYoPqtVNyEoI
+4u3tqDWmX9mhpBdI/K/21IY8fz9cThJFb5POiwDfYHlFayOjqCe/MXk9rWvd1eh
tNcAzZ1avcVwqD8aRTA8Yl6hwN5nhyT0/LuCHiSJ9frou+S4k1Jap2hmapA0wvWd
dZq428oJARp0kdzRp1mOjfSkDvpKi8jZWjMsBANh/hYBlud1vLCSZgOkxFg6lHgF
9lSTnt8s6hQA1sM2vbBLXYKHw08OOM3DEgEa61UROsPzTCs6YQdsSGVIYKsLexZ2
cepnEW2puB4pc0y+hBoAhEe7t7723RC8UYgLzfQD/26yPtAfNalVQkJw7/r+vB1v
7VcSMy4x9fFU7enku3hKUd2mPZpaNOkjG+zOXpGbWWQ0shDJmNVD2xTmGGIsbaT4
pyb4DpttlGYyDxNirvuy4XYsAwSso+YQZgek/d3FXcvuqclK88mc7QO2tnwaFhSr
hVqwUeVbXPKG7HsGFNyQOkk1KWi0t5i+acFLe6pDpqBjsklidQhUAPVMXCGSjQCS
2lcVQoTPMohnSlXrKsH5W6JW6V7Ohz+tL2t2dCx6/xPWlUvAAT4YE+hKaF2tTsrY
MhmYjykrf2AQqy9YejRCUzd6Tr/t6AB4IGXRVuB7URc5mPECPYXe3ei//E6tpyo3
9ZjNnVNgCEvJjlvPzyaharFOYLLVHzpGR7mlCccQCmlJGFAk/bl+/PtXGYYvm5b+
l+ze6EVeUx8xmJ11g4wF4u6eIu6HP6uwWtY6PeMA9kOAygNwQmuExQk659HkcoRL
Bz1T319aiqgbhQ9y4WinxVaDGod22T5ozhnZVWdDBTB8hjY0r53hx9XTTdEmN3SO
ShUWP3tdVqSIkbvW7Y3MvuZziBYXtSHXds3Lyp138C3nr7Zl9bZGN9APdTojyDuT
VigvTTkHspxmrJKc6NG9tK/4QzB7QQT8/pw7MUyDclvzf/fdx+gZQR0ARxyvUxBm
WQYAeq3YbeUKVbhkzVHOy4mMhxJOl1u3OFTYYaq12H6a3VkQrdE5bQektzZElf/S
CVvPRPZZ13IZa0MSeTdoPqBPN9OYzZaO2uQTrSt2U31NBrjoJ39+XSwtkS4HBqsG
UUtgH4Qg8QS5HEW9VjhyiLS25Wmr6o0Lh1BqIDLNP0IyIv75nn/NZoV/Omp4JhPT
mP1PvNm6bmdlP+2mg4+vgkus0GTtVArGbwIxrbDiqlQIeakosOtXI8lbaApOmldD
2Dl5eLLdDA052ayB5vIL+ihgsgGf0RcPFBY8BnQN0GfojFFteamxdlkN3bozB4Jr
tBo+uZoQAR5rYhP42KARq+jBh+1bmtfh60bIcw56g8MFpkP+bPNoPKZmI0VqVkJF
bcxSmNHiF7/NJKscZBM3dsDXtKTeuepI8FyyQq7MAdtNxB2IAmsn3r9GVCMNn5eG
y7zj3pKMNSoAnBJ6YMMkRBEpMG/sYgbcrdq722HKfK3pCPTYNM3wFnVZSwktqv2G
mHCR+bmIMgl0ka/zuoEBjmlGjEuscLQ1CpjK8bCW6OAZcNp1j4bctAD5/g0D7VT0
ZkwsVIl4oCM7A4GRDUxRjQ2am+ByyuQjwNwmMfvfdsoOxgR6A+x3srOVPrMarVKT
iu1TbWrHUsuNmi4NiLzp8rXw2T9+fCLfFnI2CjrGxvSMFTPU38AWRcJ6dVg8HI3u
wnf9RF8wAI4xQrvmnLg+9vHd4R66oU2elPq3bFV+VdEutBCEKiBu86w4jcGrWIrS
fVVH4kDO3h6y6SQQExrcW6/TWElaBq6+5oqYuccFj3OSAFc2yvi4Bmzrzrt0qjLD
BQcu+zg30D+djL1/5JUr1OPM/KkiY0SdFq9h2wqCjdQ+j7R12zcmQz1p+8Ry6gWK
FqNCkQYsulFYCj3sCOdKdR9UdDq/OQ8uzg1A0uMHErBQlqxRHBCUfKtiFdbJk8Kv
vKaYuYR5dqOAfox5XP1RRfWxh9tzZjTm7I9msV+BM6hNLoO1eKL0BqCOdIg3RDsw
2jq8eJAy+smHcQMRFFFKYIgh/EZylAe8B5PZKmO/3iORQQxmJuj0kEP6NE+u4XgL
uNFQTMl/4JoRfG4fMWV8TiFqq1l/4CXljctDrRTzxf8YQMl3S7p5A+x1Fqt7llzG
Iqt/GDKkVi7u56gb9W5CDCiOkYHWXqI3ovTUzEw3axxjpkbXiZsqr1sPSlkpJOmP
YuQ5tqVtDmWXW/aMiVCgwJylrn9tzkWQAV3l/XUZ303ybwnk1xc9sSRZl/aH0mxb
ih+q6QME3sav3G5wWN7XTTArcKSZwGpzV5GEzuTOx4285sOT8IVxUti5xoPHbNhU
fw/Fo2kbbFe0nKVHVp18y9JLFp3shgUqJJXzzmNKADOp/QaeLlOBEZYveyl8dOn/
7k5INK+ZOPQEsmuAw5q9rgV/KvW//qsu8JaxjMiw0nOPe8pIX+KCSCZ0EkD8zRhB
mOUTh1q21UR18oZZ+Su/QsLbAGWYKsNLK/ebZyopYIkO26wXtydTU018t5+4i6Ma
YtTbPWKuZxtpHsqvz7lW/1+7pV7ZjIo5K0U0Jn6ATovoqboYepReaLt9IKcvBQLe
L05pNoPvDtCeeo93jWoySgdCyZDDNdCJHMK2MdRaBt2KUNeiyHCxD07YsiPfUfWr
vZ502TaSryInO/b0IcHVyD+RYfMqYdWGkc//tTridPDuhKnKmgvm9M4rhak/H93a
+JW4Sdf/PnO6FO3ZA/bZud/0Gkr5/lRrxcIZl0MhJZp2JcBOkKBYrAHGVTmnCl3o
o/trnuKayUD19otcNv6rWGUeVZPadlAYc1LA65sXVxnOCaJT3dwaxxV/StGGg3Tc
wjkQXyGevSXDocSpq7OZ5lYVT+I3xN9izKT4YM4QVN2oBbTl8EFRW2j3Yu0HAW8F
ZHIrY/P0xHVCndG3IJYXV4c7yNaH2QOzvsaIKUdteifTJN896VHzdn/Gv1deNebB
HwiJJKdlnMaLB+4vE7jSNga9fSQ3jtMgSslb5qmkPSuYQPpOqomc1CFVTBeb3cFQ
nUrwgL79eTyEFVZcbXC/E/EwTPZKP3p1GATlPJtNdfmYtIjdV/zKzNGdezzqxQA1
AdF4FR8MrxsOXRpDm6USaZElUJFsf3+UTUBkc2/yw3H1yGhyaf/qYChVt77M3D3b
KQuGy7JCLzTAr2dEkg5KWoQDFLhkG53bY3pVeeqWEOjEfaHRATw1J8jVtWzioXap
oJZKwd15pHhk4d6+suZhMXSGsAZ6AwTeFaZaq8/xCSadCvf9KprosBF5SK7qVNN4
bqXuBxXenuvlutH83Kh3b/H86egMBnD8wDlY3uGTshwLyHReDGKrDaXse+k4h+SS
0+osNqPpb5RPDhcydEqzcSZ0m+HkfqF5yNaUami2lI0fvSA1v3pjOQuGRDyzYCSv
PD2lN/N4XLxL0LTnsRWfYDW2usRrWbbjmHabE10+iuiG3Mb904COG0snjyDe0QwX
YWzVZ/AnGgm3Sqlnif52NGuk7H7K5wzAkhGGU6gbmkicuQZ7cYdPjsmYaTV5KQn+
JVTr2DE/0uP2xT88excqjmGgxOiHeK7fmKSWWRrqym0n8ivCMi1XhwYihuDzycvS
kWu23XDuf2K92n6w2q0lCbp15zUqs+ktEwb1ihv4P2RjWwcUuMiUR1RUMeaAkImk
Exv+yPurZIMUNUop9YQbncGEuNJBT/qvdPg0qRHht5Wz3ymFPh/+G8hH1PK4pyn9
9XlBarg4w5pZ//OV4UVNL17rD+0NuSX7NXSiadpBmUESeSHOd0KWrRZXutfYgTsl
c8XSra0VgvAv6+AYPDgrIu45fIiph47Ib9d0fGpWpLqLjW7BjE6Op0obOXVsQwhN
PCBUwydhMhT/DnT+ujwx9I35SsPHBtu6L6doQXdKwG1oGq+EcQp91+ADfsVVOplS
7N7mOIVsgN32ihHKu7i5C3NOxbhOxu7EfqCALAjccfDKch1cJjZBCes391CtQYC6
t/NeRJfDJA7IEB3uhkJBMz9znOmXpTdoBae/2kOUjlTdyhOkC+43jXtwaI7L9KQw
zeR4dRq5kcMTyWCHSMOmYkiKyEeZsf4RcGKXJL4tHWFXoGnBLK25YiCzuD6bgCBX
aVxEWQ5yqOt9TOIUpRa/6lufXWzBgBYIql4K0OHVyur4oV7gU+X0klotKu+J1iyK
TN1IH1MX99XULJONYXn8SsFHiG2wlfvmA92XdD/1OnI6x+wiUF3xBJPTWk8JzIgf
rULIKCoCIrcwOQHQBwj7xmnNpXQJrx7+063Rs/wkMalq+ncf6ssWmu54vnZGvVbj
ACSyy0PIthNLi4jWxXhVF8Lw+++KcOKxTYit5jO/Om8B56PstqhhihElGMmaMBYB
/6oPuiorepd2RRhb1sbTulB/zmGHZLSAIOYZed7KtgB6vPfCbF9KjBKOp+p57UOn
d007prBptsnBj3BNcXV+y7+isO1tgH2cCF9fySys3wUA26pjytJkU2v4wsH5AvVP
BuxrapA/di2XcOZt7xmb47uqfiqa9CC2doB3L5/pCIbDoDYUFJ5iqELcA51G2aew
Izw8Kk5YF4U34S//Oz6J645IJ2HpuSaeFgM7eqs6y7I/6smLqoFeeVJngQwYI2kb
LD2s/ijn7z4AJubRP1z8zkVFjUt9+3f0XfVlA3FCDoHfQecbxsJiJd1Y0cZS+n3m
H/4hQDWqIVHYo0mf+SBIYT7zCKeqB27qv5XJnv33DPq3z+/FOpM101oGUEqW5etV
TvnfEXGFQtvbRakQA77X1rcM3Pv3ILC5ZzVoWGhHuJoy1YuPrxqXGuBKtagP6XJE
4V1J8/utz21nw6nQs14pMYp311r1YdtnlSJBUSOR0AglRHZ6vXC+vuy/wbxC0+SC
ycv2XLhDVAlXEhu2DeLlMhhB5Ca5BBjwOg6WjBQT6k8aCTNAlLh+zJhVr8NnEl7j
CrRtdGAyJVoTN8eccSninEF4XdmMPaCErvZytwV22S3b68whEjSs7bUf8AGknUqh
daXqYBTMMDmH29yxP7MvQe0B4LQ3r/CN73YECk5ChHhjstT85/3gEgOgqdBYwhqB
CUEW6y3lW8V6rp00uO5uuKO/aqnLdfR2WiDaif8jYnj/QxdUdbSVSt9wSJEDoBQA
2Q4j4TkFe8WqxFOwUKzyThLEZI9c4YxM+AyEMmdvU66J9boDijEgPDZxcP0XKqNs
4kTlbCbWQi8jJ7um9+YUD5+dzAHiCuLMVxdj5Bq96bU39CXXg32BF8RX4eHr9Thc
+SL7049MnejmryMsYukdjAraircCePZDqSEy/Td/KF9EAoDEALU28kNJ56Cw+o+x
sAKT0cz3DikxEXAvR4JOxPpJSuKepqZshgyUiBKqG+xbhVzqF9RUmmMGNy+L2p5C
XBjQrlem99RWo5mCNcOhkBJVo8zfWZmsc7PfDt4dTbmyi3TjP+Tj+4D+X9vrbTQr
wKxF2QRa5xxtyjnm/s9O5Fg7MWG+6MZszrfkAqoPT3hJftSL5athvG8c1FvR1GbP
GG6CJ57ZvKY+TwxN7OkXWIepz65GouKb+jd0VBmI5f1nsHzQq96hFrF25hIqP5Lc
53L64y9gbM8n6LBmYezzdtVowFls+lKcHN3hqDbemMsQ+UvFLeWy966aAaXtFmzX
sZK4mFkgw/3wINM7+AsO/mH6cFezkQTacfvdP4wkzeqbWKMpSfPJfVfUMJlLxe6h
98JSYALiKf9rmRh90LLQCBdAogtrxQYzI6AXNkn0dLaiU6hdmrpLYPVVyoOeB573
SOlTnnO0bEPvxObgyC/wREuXcB0tStAy1Yrr/CJkh9KY/xIvbQAIP/pxNL+maJwe
PKuQPV0jHNHFRwAT6NEmzsAdZ+IwOpftEFpUz4/tI+KGvApJmoHjUAHeOaT3hJp1
2HZ+sXIhY9NeFZVdRiPcVDFfV0ZB+ux5W3vHAptffMUqbcl2+VQi8Gm4s+j3lPh+
actUyMg5bea85T0wsHy08vUnmb09uoruPketCLMsGwyQu1kG72NPmhTl6q707F7y
MVcXPrfgP2rA8uCOw+xd11kJfLu9DJDtZwPn8u5l10ble0TDIFp4HLzRDQ90a8Th
CWR2p3kQHOXZaVFOYclvuWgwMsLB5o/F0sE3uX7bn+NqLWBt96/GktjOwOifeEJu
NuAXc7G55WVEja0qdwXJoe1kNTWOgFnIOSM9j1b9YdOmIIUWrdcNqM4wFrpTtKFd
aJWyO0OFJBfL7z1OHLUA4ZIUEC3Y3e4QpX8AN0vx9nC29wmn5znKxzce2qgRw9U5
j3/CBWyoNfIbDylcGxg+FNJz4FM2EPuFr3bGNy8kXgSlo8JeT4Kf+eswGGfww74E
b6KlB3PqNBoBxO/6YeSgn/OU5oTvfCdqZ4KEKAF+BxmDu7G/BjxZkUmFFgAdSCUR
xJXye3GHVLu61Ql7r14zPYUhJ/SMVX2tVgI2xYWErLyWoXCr2bBj1RcEIz4PEn+b
qZ7GneK7/H7IjCaAiw9s4DhEX8spDKg6peUus+RXSbbl3YVfKMkJLumXBNk8EdZZ
oZR9AVhSfIS72Esn3jgH7B+aXYb2m+G5m9N4KySexI0Da6CxSBh52dqp44ZYXpOc
NLNFsB19kPCUAdLTddYSJRH3qxvyXuNVy0F4M1H1Ay4ErztZGu4OfZRT3rQgzI6w
6jdrAeLnEgMCETZf4H7DmxoExs62GVe/pgGnVAHy3WQZHvgJXGF7LMeU/Gjh3UYK
2AKwZQL9bi/dyddR/itPCIGX4L17KEoCyJfFcURw5qYesbiRZhDXZ4NH9GoNOiA6
W6yCWI1z0G3wDHQwpufgRFR4NY4yrAL8Vr7wFb33SQEbatOd3Xgk9xd4uCc5V2Ms
XIdAHNhDo/afWb+Bah8msJ037bX3ADOdvFt3l8eLBLEXba9w+tGO3v9TA3vJQStu
5OiYCFKSa2+GWJvJWDMIcuj+hrjsVI7VGd4b5g77EstoAs2mIeKh8fow5qndPNHH
L2Eo9MLobTZufs2vMSoE5Jp0e4gllfJoCUVdfuTjegzGtIffTBXY0//ZEOPqICLI
dWu1HWw8GLl8JuxU7mdDHmgBfDaY6qvpwBUeoUApf/J/lOv1tfh1Ltv2VshwEIeq
GeQQFIagJPe9O06RFIJGOazML7i3DENhMU5TACisui7rWAnYvuBT64Ht0uLVFovm
W51QMScLlkDKpr3Rf3vs+aSwh2ppGcXPpxBCcZT7//8rQtOt2yKesoULsM2noUbC
ymUqy8t1a2RrbgnokbL89mZ+Yard8dyK+a2uu4BHzK0++lFes6xEWGHtrstg2Dv3
6S5tGhSwK0i1Z14+YniagV1vFsoTgYTh5ZgWL2IkX13ltIDMJdMyllKJrNLO8eZ3
bUd8UUbUTmKvY6mQQ2YITCJNp4kTItM58Aj0/F3JLNhxG6f6SedfbzHse5vDxy+W
UqVy7U1WaHkb5+CR8mZ8Dpr8kJcuRqa739XD+IBJ5clQlwLpvLetE5hBQVvBe01n
T/2E/JAIdeMeOGc71A9Y+1nLpEXuQimqz8N/wHn/USItoVUjxX07yN01NIUanYMr
2ZPmtE9S+EFkAqsCj4N19EEw8rIHENyTtpy/2gRhzsnZNyO9Lr3bVDR7NPVHbGAu
nrxwJFgt2CtFBpWTupHPxuCkH0fbtIPrJSSXbcbeJCbUs4PB6hiQJXg5mxp9SvYe
4lMIkXUoGI1I/PjwBF8Qb6/5ePdn6QTaWqJwpyivP+XEqV0ZSXbvr2AKKJgWa+IW
3UWHWRWbQ/A6wG6mvE9BrSzAmDuoQHPRCrIQ/EnJvMfGnXnOGtfS74Q5aNxj58n6
KjBGXb00ETZEQ0q2j/lCKuVDMdYAK/4+aWyFjLF0dANh7NvqcvX5oJKuASeKrnp1
PJrX+wVd+eJQUHZzqM2nSjJFTKXeaODjxShVj4Nuvl7HU0PIXV+UeEk9q/lUm7U7
c/hv2tJ0e0qdIopQgJcEBMVbxWiNX51TlRK0DX6kpa2ekZsTfmFLqAydfOafmWMs
U4S9oOLHNdli0JTEHcs7KaSqX2O2p1Ipm0zscud4rsOHdhINVARjcqQWTs9Zoaxe
hZRSXVCH7hDz/c9OCLk5K5Rz/ALowg18mDXLahv8W4vMMBT9hfARa/kUnYXSxJtl
bbgKgvlAo+YX597WuJlDCgFGGLTsHeJFq9g6wpeOWMO2StY8n+5f9htIgZMEY0d+
alY5VxeVBkpql27F6nrNeofQHMKx9ekmM/7gEuIsgsEtozpen8Mko75WpRTF/Nti
1EyOAD84CmRf09UQqxb2hhY+on43B5qgKbHXVE3fRpacgnLEicTxl1Tu3w4se8VQ
9P8I0taEhxhwdzgv1yqJ5SmLOZt+B3HhX2SIxYZgJ/4msr6Co5J+hjvmrS1RtJzT
3gcWiGOg51dMwywHuHNO7hbiIr7d+B/38jX15zazLv+SRYc2YYK8XiMVrTXhdknb
CWiOdkjMTHMo50PsytBS3rgOT0uV8/er/FAO4sQyfnwgaijrLbABX6lqwMLfFfbO
sROBfCo1QgnecuzsHFn5+HXBGQldownf4vsZo5QExan+RQvq9bWvWXn/HELUr2nZ
wKb0P7+Uiypd+aUzJAPspTpBOWEnKXfXvJTbTHfF6tswjVpX68/agl0lKiQyWpYj
dZqe4HsG0Ha84dLL+GWwS8qgW5Ae2j5NS0jmZDL2/ykW4wghRVFG6IKyu0qpSU+N
OLwy9d9ohrS33yx3F6LYMqpc5g4gp8Hq1qUf2nprOY9M4KioPwb5mOvu9FvT2Mnf
Kfo4hupJB8asBCiL5+aSTEhuGh9DYzQeRAZkRbQKJH5lL4//E7cO2tYJgUYKxfgb
+vzoMx2h1Gopbffp8dOBJYhhoDTv64ZJSZFuVBgSMuXfON2kXZ+L0ZY8ritsxiPK
JVc46Hy1JSkhfVPsNhTmU+WYBe2dRT6aYBXADVY0wikYYeMyomMj3HpdqQkbgcsa
fC13lcLPbxYgPONwK9GXvqBg3YklHTOydHnspTUj81BeW86wSm/4cG46SESPiEqy
raewMD5/Y5zpy5lB3DXPjR6v+1Yd5Q6vlTjJj/szmffh2NDqE5GHGqveorgkA/Mf
UlPhIQY084w3b9pxAZ9/XY1O6we5ybp2+aKxJe0fiPjjgv77r8Q1MjaQAf/UVUQM
KIg6uYe5wE1OGZ61h/WDXyxiCznNZvsimKq3VOIMRRGpoIQ36/KGo7VEqKxy68G6
R1i7EB+7Ep0KeiQS+DrHdoIiHRAha2XdAe7WeAnXjgp2kddB7O1SNiAM6yq2LMUu
A3npslXa+LJxIhxTD5pWyb2gt1vaUuU7RwQX0CxAOpRmImiGkr2uwyz13VbNbamf
MibfvIvwVDWOXD+qk+BQB8lRtfGGt3EDacYReTb+QlZJvJ4ZxPuhJahZjfbkEODj
QkFe0WXmXmhBsOWxDuWdB2lULtt33q5YQMtc7UJhp0qYhm27422VvIG2n4m058+A
GVeIIfDYvwkH7/O8A4JU5CuWQV3qapLpzU9lOJKxAsfoDrJa56F7+bt67ZCwlNuU
FEpzYcsJQA3HYURbVQ4isUDDABWee6M++fFhPTM9G5PvHybnRuneV1IuVwnu1GBk
U0KgsvoKA/FG0gFdODIFhZhyKLo7zYiAnieIwEzGhy5wkH8/KeD/8NGE+c9Jwj4U
EBcitFzv5Gy3b8+FC8JOTxWZCVT8JHEfvSDrtIT1llTiP/T8fEDqT9U0HsyoG6/C
It1t7eYnyS/5SigVBbVNgbwhVXiDe6GR7A10n1mXAAujfzvcEWfjNIT0JFvoWwkD
x/HBEdV0vUez0mLkQbpMs70crnE61h6XKZUd44wRmD5TqrakGFMYPY/XJ6qHRX5l
bmYH3LzdyKcDev19skhGSmSVfGA9JEt2rT5xk4u44N7n2FZ9rf26lCbIMd40K3yo
Qyb8PKVg6EZdeO3F5mTGfsCH3GFw1Yt1VXA31AB6q3nxgiztgrNAyhuiMlxiyT/h
xyUfzSV8AcMjJWE0b5597qvxfyT5/DXS1gFRrWOAe8Fqdhu99uBhL1DIg9t89RpI
/pz6H745P60U3zEXx4w9youQ7qcdfpyKNRUYCKDhfGelWtKUeBhFwq520r/rN/85
2RTUCXLR9YWOTcyxkQrYZduyrX06I88K+2a0p3x4JRqji0kRScN2w4Hmj2SEPGYl
uOLxH7gI49FzEt9FkoV/XIXiHrRp6PPEVRfMnAkSyTMiVebsLvAzCs9eeZ3pB+y+
fZO9SyFzhGgXOSXr49gG2LeKu/7rr8ETfc7D1wMltlAR+m8/9IT2Z0o50iN3W/a0
54lx8pqSSe/+6/Pl9razWKBElKzZBAM1+PFG1tZeZOeQccx/kCQvHdk+B1wdgk3E
HBTGsRdGShUtxuhRd1BgtFSkXpzyx/z1xMblkg2UDsYxDzlZjC5Tm6xqD14bJGnF
/7Rbk7Ra/sc2Fp8XrgdxfdVgdxEYALLDaZbF+QEMr5f/lhLogAb6/BrksRBvCckY
sf80MLRw96fxp/0bFk8yNCmwvnej5dBBoCIRpC33ln/1SJ6c65LloO4P4qC1jyl6
VcaSEU6IPMU9eceR2MmYJy40mH1Bsalp5fDpyQqF6VAj1k/rNUdW1PkQB5Kr+yHT
wCynZl5YZ0ibu3wE/qyqobIi/to1n4NBJlheiSE5u190EDyR4eAfucMF4Hbh2ucc
G2yhQTTz6l5QFsICVv14L4k4QrbNLwiwXKR+29glvBv8YQLrkEVUuJHiXFyA0UUw
gVyBoRTnVonSXEYRevlsHyJhK/McaGITnR470p43GtmiiU+Dl16UmCL7Aa38ou0/
m48DlJ97aQx93xiyjo7RRkS3zHNEXgQQpMYQlefrBbpwcwqMSPqYEqCIpGBrSPWF
QtLGwXHN1EXH4SBFrxjp48ZPD4Bb88peE/3vLbYjHJ0ZQt88TqiBOYdu8DJo+Hfi
x6HQ9UZgBDY1VDMqLjRiokxd0x3RVGmRioLQYytw+mAAMW00ytObwQQOnNVY6tZQ
1qRmJchV9NNFtYt7oeW4ifs4K4jQL2jQAY3MH/oSVBmILRMicD7GS5TE2q5HekRV
UPwirb1MRr/UuXB3DrbsKGk/JaxgI7Y4R9IPiPZA+nZL7N0fBI5ZxkbhNaBKC5QW
CO4TE8vzfiA7avx3rgRq+lEhpM5P7uhcPgsCmBwkjRJ02F2m/4jX0nETcL062Lg9
9bUnFGc6c38tX3+R1zxvCsizFKDfaVTWz424HJCoHVcdlMvYb12JmUdGFlMMvnhw
FYFLyVHw74xGjwYKT66CdnVebRqeu74CmOx9ruhATa4a404KNytQgVjsVtSO4cGa
BEvhUGJKtXZ5i5pf06AYNluQxILCd+qn8OuN0KUNuvL0Cio0uif3hitbGE5brr27
m6MQzkHB5U7uFsCLLxCN2VDn5UF/3FzbZzxMl+bn2ESOItYtpvVKWENWEG6DP5BX
259EjvAn1hXatgN44WyKiUa34iyjIUHoybu2wp65RMeh8gJcMVwHRKOMO9KxRgES
D8tT0J7/LS8KjOtqYRPdMXI8e/t9rux/XcChYntYzWqwbpwMxjH58kgEAyRFiGzV
zLZkpSzEUYvEZzRv+oQ/XvafVaeN8kHIDlhFDl9K5ME98R1hZNpy6bY9q7PkKWer
Y+RKi1kGrCQQbgadbgV3mOt+S49fzo1R4XsLv4Wq4HBxUIiEzX9V3CyL76bQpia1
tWd+0h4lI+teRx2l6vgzRqzqnNoCAZP3ekjGxyQuyAfrFVYL4EcnJ5g7uz4hetCg
lw+Nt5/j9vn6eovI65s5qVYUEJF8Rn4tBgY3/I0T95dXOI78kFoMoCCqZGpZn3U7
veCQmUjI0h5hjfAmkjeadkeZifmqVUAFjK3+RFSIH7gWBfxGyYipJEF0tZN9GXIo
lWJbqV4YXOnjKfGfP5U9MPFjmm/s4ZxS/aoRKa61q48Mg7Eb0C+OzmZt04kJ5H/g
jAjEwxCkAQ6YEqZ3L7Q9nMTYGSwJmm8nExICOy2M2d6sKt19k45B1pTCLML091u2
QCwIFAjfTHy4OmJuUogwnyPfkHqzgRHZsL+UVq9YTuDltw9dYvBe+T4+M+k4l7n9
KzRx9vLLYVYlMzFalxPBZamTUrWM+Io7hlK0rG5zLTKDoiq1LYri044/Wbi3xVyR
G88dfIO39b5qzqomPxgSA7dtzbWRhQAFXChQGuA/0g/xarBcQUlKCTx3nA146QNm
+NPMBGvioXXCumC3mGJNpAL2dfxacMuhFtaU3m1yv4E9xLZVzXtjeE6usG4efjNv
cpIwPRVJPNHQfdEAyNEfZx1wiOCU5+uKv4LHDNkBGkjMcGZUmCeCNYS4i2SYpjca
UuAZyNQyTAGaOkIfBcWnPnvYJtjwiCtK6m4FHJ8PDmp08uFV+14vFaz0v37WjKNI
ZZrZkn5D+nDWBnm0msCjyvzJrjP0sDXWdnxDEw698dYYKAoSdABsYQW01fzKqhbM
xtL15C7xVEasyIYbKhTyKTY+gx41M/SlXLxImuGI+7how9QoRi1EZhBVIaSHaV69
71QdqUpES7IGmFUNDOcIwMQQGvs9Ms+Xbqt8PxWvChYIW0EwkJOaWa39ty13Kn5B
sb1rb6CxtcSzmn2fj2vSPV9defwKPb4tElHsIzoMHtF/3sFDyJl7ol/i0UTEWa/g
Qz2uBe1mmoQYWRu2BHx5V84n/WyjuwPk82YNVkAXXH2zs5jR6UuNzgUGdRRCEMkO
LSBsY7LcdhQuNziaSjJhoqQjx4D5U8EPquGx87rqHdKQypCAshO7P2RnE3pWA5By
QXURtzqJyVnuYJGng5oeW0rXc2/CXObKpwteKpbNyQcektV1xNtMjAht7odcWTHp
6WrKMI9mZ+CbVjVvw9fQ2EYgh9i8gQIujTh/CdxKUzzYohRGZ03UGtZY8dlQF5fB
vyymP2q95o4o6+vMlpsxMMq3XDUmzpKl/RMYEbtTSMJpOZzXDLdHhvGUgEa+lWcY
zCm4OhSUX3wkZGi4WiP+wBDEw3sLn+479Y/np1t0RwfVNoiY9+WAGWzaYcYHtLtF
gv3kQCf3YQ+das4UkCqXlzLAuTy/kymy5NujYxopzw/sxgiIdU1vjnp60Kx2STpf
1G/SO1Q4CeGy4Rd2RvEB2w05fSXudR+5p5rnj34hZRTb+DX0ab2lEzPSpWLaMzp2
UuinJx5ZKJkXcgkSsfzMf9d6p3ECYfa5kYtYffFS31m3FlElX/C6aBXG98Kc4jaJ
vQbfNeGXD4F/8Hf0rvP4JsEPq7ASKbVvExvCE44pziuLwuJhgoM6DaA6hdL944Rk
i+YB5xFntZtfWuj3K2gLMWv/vkYIDEIMIt/G5gXA8qzgMYQj3kNv0/XahwJueWdT
8TRf66UN+YYEiYYXNz/h743/quHYTwzsatOakUOWghkn/JlbE6BGPgxoya2c70Rz
sJYs1wYM7dK3QXO5roaoQt9vZHjDrkGEIS2p11HYRZc06dBG7SoyluE517K35flb
UvPOwceQNkCVQ/tnXMvbrtRCYm4ePX5eiFCEIEBEW+aU+yP4E+o3wTukYeqvaRkN
QodmsjJShW2eFduwPUj46dg/tDhANrzMQHefsB6CBh+h3KjkS4sIPnndIuhSrdiD
MsutBl07/2K1LPTocCGKNYQs38yIYgwAeNGygA090Y8uT6lgbYl891SWT8+Wtulm
NKJ55B9GxWFeo+Sj0LB0e07Lq3sa4/15cdsZkJNghmiRhuL2SGY9OV4YHUiCTmyz
czdBjOMCcEscWPB0GUcrLuiZh2BrQ3hhOtitkA8BQvXStCP25nUKAKb7KL6Hwz/X
KnIxkSgTj4KvSMweNCpMjCX8iF3kZ8rrUqivaWGE1QN5vE30Y5JNX4MOf5AvFcPw
TIb92aYlcSRCZyyqUGp0VmnJUq51VuxkGX4Z3mh2NJJtBaRVs7Ron+/UZaMk8CPh
h80cuZuHB9RmUTqr3ZsbDOAJQJICXiyChRYWqu2Lw5itnA93ygTeCC1/APPRLRau
fAhgOJYs/BvA/z58gAuHCdBFpAg9mmIL4hZy8v9Cw9nRaNkDTU4PYJahWA5YOfbS
hEtBdEKptfE8HB/dppX2GDushtuFxFJSJhUJgVpKg08XvVrJXueWIw/VMUeNMTYT
49DTYvKkzeaz0/70udNTowFTmgGJw3cUGpRaaQFmfrq4/9iKAso/0XfEPGsllLfJ
kIM7vqrXN8D5CQGby3mCA9Y/QBVaDjSE8LkuXKoXvn1OoWViCYd3frrzvQbPw76S
ItvcdQ82ZDH/4X5SWNGrZ87FQpyfzLZObCH2kyEvbRCOnHtIt2Vxmc+UDY0TnPtc
9EcU+Evd8tB36mKh3qqkzt9Lu5H91OiHJrd8pchJ+ydtGU6TtXnMQwWC4Mc6IYS/
hL516WEh4ZIRP02VwgfXxZsDZwGx1cu4LdeOR5VlVvBwfUUeGy4EpUw3ZLG6UVQk
QrJTJrB2rtMbAkKn7zkmPNvtctfx+u8fcYRUnUCo0eTdmQuTkaaPwJkKQ5k6dlRE
Tb1gD6iOBDt4P/3xQNLq2RJ1pcLlr5DH4HAJwe2D09NAQ54AAJZme37Mok9Rr7Rs
I3zReskZgP2sOMtQq5EdYPRvLVlOPraWdvi+ivQxe9MOjLv/fT/D/fdKaCJFbUzN
mfoomBh38L6R20CJIDYeFbP9wTRX1d01DzKpA1NRrpjdRpUxcL5dWE945/A0BLuY
qoq6DLUzOHOA0f3erV4Pc0YnTRruqqO+7kjuxTY/LtbpfT4tyDvIM1luAxZBEkak
fn405ovN60sLq5/j0loUR5cu5wlv5sLAz9EZ6CVNI16e01NsFC2FvPAwkExaS38A
ZOxdSls96xEcHnRI32cxynSf2w7GPWbLmFLmX3FRU83nbwRsLQGLy9YzIX9ZS5Np
/9Gg590itNwH43+t/2W6zKFYdACSaEvl2BvOivGB2xL23X97CzhYiXciQi2a8SVq
OwIO97WOK4cEurZ5BS1zpQtiux4n4m0Ml0V9NhmDybzZcNOTeJC60QewmBqyQQyK
OeoZl51Bv2Ydi3TfpvXBwG8bKDQAsBVBpQQ7yHg1xC3XRyeqOFxaXIPM8Wdd9Bw3
+PHtKOkuVOxdPIxWZxdR2aL1eQQULzB64/WOoIhpzeh1WdOKMPzRJVd0amsZbHoz
JlV2CHxf/7wgYG6hOOsPOFpw878IE4WQdUlQWG+HBzVwrOlr4HgVuK67pOG3oqdu
8TkX86hFzeqp/6KXYVau9EMDY8iaTN1Ujauo3iVqHEYk+XfXaqEEPf34SJMhIOGA
szGAfs1us11L28bt4jkCOITLDwtXEuN17ZVpUpcn15h00Lz8Mu5M3DW08z2G93qG
r02AeDl/J12rV0ohY0mbveGIlzoWQibqayiuBP1grxbt8rU20kYn5u7eXav186nq
XgHk8/iq1Om2Do22/3K5ow4fcr/PFZCFFQVi+XH51/QigzOpkGtNT8LUFoHg8d7y
aII5HO9+CpC9M1ZOm3dsBZAYfsx4wJ1Q2iSnJcFvzng6GiF6te/X4yCTNkNkU5am
dE8PzpNtCyuP698Lt3zVIJbcVEXrxN3zhJYeUVPGvoXOZNZzl2H8+JPklMBUlpXV
/dtT/yvcTgkCSwFH5ixLPg5EzC9ZuygT/pCvKnQgDP933vBYjVrzMqiFwHZfUaFL
6negBWanUqgIY4vtT3ceLbRXx11GHpQDbObud3ywBi3pEp3O8ioIdbLg/BnOhbKU
gaxo6j0oThQSV8cxTVxuwmTim/jCrAVc+GEVdx/GqLiC/aAvY/+EI7orVIKRvLcV
TwShi2lvmKJfnAtrx/uQ3icQq9ypR2AFispMM7oCBE68TSRBx5HnXz9PamvY2/pg
0CfOUwY0GNUh079/cGdTfhwhStXekMK/n0K3JjH6y4DRuwdWbrE5NAR0cyFQuHGP
g2P8nmwiOPXPJrQlaGjb26kC94g6FYIX1bUtMKhylZpkekySxe8ee46ADzr5MSD+
+48MZSvrQzWqOQ3Q4I6O7X/DePhSTR8NPmLIdpGYeAju+J1ZP/jMf0kzrzZNI3Re
UacEfctDUC2UnX5N7upwCBBw8zvQp0zzUPiGrp/9ez7BB9pC+Az229LIt8IeQXzX
pBrmI2stnMFmxwuycGRYiDNTthVM4LDSqXvpOljZ4YlOi9TxpAheXDv3l9SJoB7l
WKs9033ncmBUIYKo1NyBFgdLELtGKjte9L1wcaDB5sudsQINRv4CaIkvlDLO25dT
aNDp3C1/W2Jq85oCzOVeJbOTIoOwZobFHKD8+BmjHC3hl5Fa66GSmD8Pp5ph9+6b
6FSG3ooYPSuqfIdQTVYV5qKbNDDF55z2GT2hz4R1JfcMdENd7Ap6NKmDNk1xrvbw
lTWgijJJyRJbl3BQ64LCsVeNa8odVLdoCgnOAgZnGNfL4IMOAwzH78hyZ10Q9zrx
STahXwcqHTncQL6Y9zoxQ8ZiJ1FUTB32o9+vvOb+W/lsXtkCvmPHui6GtxJGEkxD
EnzmMAsjB++IShzj2yTfJ8oZzRHftEfSFo8QWCfFJY8y4nIHdfzBGWvXQjzmi/KC
EToRyAt2S5ueDpdyIw5VFMYaMbuBjvZGrbdd3P8KmNNHkd6nzCRC61FKjwwS3UVO
ae/lA4xhWRn2ddWnqCbMNZ2XRbEGPO7m0bemz9ch/ESarTNc0+HK9+mfNi4N1RWK
XXEVvmaiDkBLPHUdqNnBQVHtV5itR/JUzYYsUItOo++uKnSI25Q6mg9assVLNFi1
8TEIs8OlNT/E7MwU7pdaWiOlf/pgnc2uNwlGCnHfStJ7KEeqjBcIPh1fVxEAJ+IP
9IbwX7VYV+oXR1hgxEf1w04pQIDsT3NvZ5PmNXpvtqS55ZonUoxREJRhTx9fDF0V
Ih3JNCCLsqfc2MtrmW2GGyuY+5WbmiwkS2ue0Q7zJd6kCKDAlOA8HmQ+a553d6YK
lUsLnrUN4vs2wDBt7Jq/M22xUYzO60mfkXMWmpsKCh/t6cd5urJEkF5SD+xwOXfW
Q7uxI8PLD5lFL7LHrc2E5FSN6OogGsGrV13nCEbhZsMzqB+58mlkACWtHk2M4CEL
3Y0tmDkXpdFHT9W4/pkKom9MNxKVZLcStis4AtX3ANYVkQvmU0qi+vjrpONp5WQ8
3iXs1AAIdwNOCNgBOCVe5OcX4bdGmOIfB/NgoewdVX/sOzc2b78nYg8foqAi4SS+
pahfp3viGmOuIrwzOivCA+0oC6BUB8JrEhP2f29rb7aiKIbe9GGHg620BkNwyJtL
Pi4avgjkb99WpQNAgtDAYgbwE0KliQTt+gUJWI0q4M5DiTgVup7XSu2X+z8gKLD/
VvcDSZXueC4JtYDciAqWT8YySNMsdIJynISIqF9TGrjoGU3RqCB9af57imKiJDV/
X0NPq+Sswnc1nIyDOjQwcjW6duD6AImFu0HXkgmLQra2iPdpUlrXHxOO3vKKOGsH
oOA9BVu9sRin7bp+dJLqcqen99K90DfFctuBopWzOFUQvDG6MQSy+dB4dZ1qkUlD
TBchlra5qfd3U9Pk9CRW9bFPp2igvcOa4+cNvyUPVkGlmgGP0BEoQGyIEYhcNsR5
7pOsbq6iK+Xn/Xis2KsvQYxkkCBq7beO+soy2RdpLi4ry9PVl2pCyXjIZgSjlIop
tU8evtrcjU774/7kB6TKsI6XS4kODirMg7ACbWyBTyHqNPEMu4wtUhvfZpz3+981
sGCaYTAMxAu704GyRwoC+puAxPvoDo+BqUJzp4TIVjbf3ciHTU2tmtEdAkAc9yQ1
qMSLNV8zU4/qZPON2v7tB/m29IF3m7Rnu9mqwBEOvG8LaLaLQDO2wP/ef951T+W4
RFztKV9OPBaAU54Y/AmiWmvP9yuv/pu3zNWmOprepD+BISYgLowJURBjo/JX6URi
a5jN3bpnpJymkMTAMkzgpWdSbDQKnxxGWgpMD1fYiHHniHB30Kl7aRZAJkFuOyJn
uYf7jkSM1Oj4FeLmgSkv96FL/RQOqvmXKJvB4qwCYHIJJ8we6NAnXL/fJCeeRw07
Fmvuh6iIm8Mj22507KUcI/ortIvci/MgszY7b7aAXvFy1Peg5mRKFdubS3OwEamt
V7cVlz24d7N7BWjC3qaNZS1heEYXOEAe0GuPCEZj9aZAhnR0iHvfh6esqkTQc/1+
PRd2DFXQK/il/Tj5RCLJw+0z6reUr0YY7tCbpL8btsmD/42UxXLvgfUhD01X+CIb
MCbT3O1/RqsY+4j5E4U3UA67QuPUVaQHJb2igLc4an/LWS6/YTvwIk5coXafPBKw
AxtsgRIdcZJUT3EohvAPW2f4jM2WcQuunhwMoLieA5NkUrXFqdWasKwozAPo0mMH
KwOExo3yV+DF1dJMCi3wXxaM49M9rm8im5ApEXFCA4/LXRuxbaQx3Us1YhigRAlr
4ipIV4pR54aCVIDD6RD6c8sQPHuJd7Kqs9y80XnDN30V7LwbtiiBa+sZ2KuCTjf9
GOPgBxLkM2Myz+XXAAtpZzX9VzM3E+fWLHctLTionmzqm6tP1Uis8HKpX5qKTeAk
93twr9Csrka9dZqstsDuIALjnnTndoCxbVZ3webRPsyKRG4FpdopgonzspwxXDEH
rc/cqTYpQrfwm6X4YUKkvp/4byT0YnPlpidRnxtQBKrLYmoDW+lxTKgkKh8mk0xt
2Igqfa/fhsV4JKadSsrsAdc9ar2gzxprJv2AmTStCWKo/D6L77wC5jEfQo9UJGt6
3iX2gSxACf4R2bNj5VZOp5b+l3tycqOUK7T+ZPu7WE7SHoUkZEhSStK86MKnWP/I
CxBPpS1N2hEwXVrR0l31rUHa5Kbv6OhVX/ZYYB+FF/cmxCeZnA08f616ekobL870
l+fyeu03SW6RTck766W+IrG113d6i8OAP4yz4k6siCPjFLRHnPRqE4YELb1FVgJb
mDY60s77VO9oT+uO3PxowWjWa/sK0e2MendrF5AtkLyvweydEslQuokAESPVmmN7
wU+wevaKZVcY6GnR4lMKb+USW/5m1Ckmun0g+Xt5yTT+SqLzTKlYoBAfKzcFFFuW
uk2i0e6bHQmWfPluvdlSAH7X7wsfpvtDKg+XZ7UuTbPlZYF6iMH9Av40+PZiby7T
9XjHWf6WmmB6USNYN+gWn4DbPx9AnhNyEKcgIbqxiEKmotAh8V4r0tvQrk4R/Ui4
GqW7AOAAChC8PRnGrfavPPqcCg4KCZ9Gt/Y1CW7qXjG/UfjzJYcn+UxdCrgEuCF7
m/ka8PsT9CPMxlpjsZ0XYcDd0VMVSH4QqlwTKYG9NKil+HabE1ogKr7Jkhtf9zVs
DIYkoi7HoQE7vaCKfVscTa+r0AkvuIipdDlw/2GnDqtBKdZSIBeH0mcj/Ch1OG0P
x6qtsqYIKFTpJY3dsgoqPrhADB4Au4d4hP99Roc2hmc4c4w9Yd2YoUuyKCcFrQeZ
K83KrzfM23qIQakqQ3P/G5iMakam3hfIaCnngOS9vqe3/1shW542e5uB7GOTZc8a
Vg2OIxn/o8L1UWNIIGaBVofSNKzr+qRufxxk7UU7/3bLTgiWYZBxOibBBDwvlHre
0A1K2e+Wl6ehaqyiNqVAxzw6xgyzMq9uPHOfe4AGMmp/02PJESMzaS9HbGfCDrcN
LoAcJlnqGWSGAv1uOsYr2z0gPce5Vkh3VwN3RKR4g851if+kZGKjYh0NY35yfvIb
tSE1ZPlmVAvG1eK2KAxUD7A2J5eB1WKyy9Udnz0PDWcYwSTTzVATxJ84Qht8MY42
osIESsYSSR7h2XCXMChfXFdpqsr9nDFwz+uQO4xd+vOoBr/J6CVNZdUawMRhPZU6
ZD5Gn77zFOPtt3AykHL57DGbXZU8YjxMYns0M/BlIc0fAWsRdefgUXDf5qKGYbz4
KxTN+TSccyM14MckHtMjRs0DTY5smnthVt2DTH9PZNIeA8k5L6mpxHXbyieWThm8
dLq7MRiPR8J7vROqrHnCpPHSP2sLlKmvjVew5mZVDRNbyep7cNl8GMKkJZ41HefB
0Nt3n9rTQsk0u8wuP94yoJ8akvE2bh4hYt7fTjYRmqqbirfDBZzYQEs3IfqSSC/L
6LUXw7Dvu7cSCV9IOsJQK4dcuHQAjtSuaL/h8kZUeR639c++Qat7MJ05IIN+qS+7
emjv/x7zaaH5wR7Fjnn61dO2rR0qoGnG/z33PMxhAdeicRDqWEVRnQQ9qsiqoll3
dtvcV4TOgVDQPvATc9fwkYMDROe9EC/igAjcx8m6HPHaRUZfPfp4+C7OJGxmIJth
HHoIveKJulq3pN5MpMztjz20SspN1cjdXBPC4h7tlXQvwwBa0EclVANadpMsNcNh
YaylwOazD7BlXpY/ODkza7bA1dFCR7jOXQ2cqgg+YsBhRNUmq7zyTMWuYxEUwP14
tMR2BUYZMsexJZ7us5jpLryvVDlC38ecIeXtomIKW9/IcYMPzkSk37jp3WfCmXR2
3fAtoD6SgvOHnETUC3EWGe7W2jW4oM8Z1/r3bK5LI0a65ZcYhuFu7av5ictwEMDI
E0jnUB3GHZo/cieq/IhdgOENw+fkzIK4YanPixOCPp4WTVROyHKCSNXxIx6Jniyq
VOSI+EIplw2uc7PwhWo0da9DwfjbIW5mpk39/3EGxYrz6zzvoSErhmK9BIoMKs5q
zRONs6BKO/RCAFWyKORn15oXAPmnRkwGpohL/u29lD7mU7Uwi+xAJ6DtgpnJjPsE
lEaAeWX6oyR3Zc2U5QgoutMegTw8qmtTVb+zjxSvSHvtZNkb3F7tbd+3EkhlmTgv
k2Rg2Dwa5TEm5IKLjbWhLDWOS68+b1W0vHJV8SrsSWKTIq3rH2H9FFDnfc/v+7fO
niDoHRyBb0u7VxGyCc+uW+NmSJeNU6k35rU67VnEDRoPTy2ofWBsWY6dslFKc0OL
4SHTPMM5rEW+hZEI/ZpcB4ueh9vec3lVxKngtKCbIWueY0wma6W185YVrEs4Ho1K
UW8hYjOVCLnN0gynWu2ZiMynLzIhfUCqIQ1fuMzvh1trOelqTBOtOk16689ZKMrr
0MxfxQXIxoR5anAC3ol0PXDRgRqD+0muxoxCGwEaKN19odFywEwCxHJkZthGXC9J
fvwNlyAO8wAo/FcMe66bbh3H4hKWjAwIxxEULTDf+wtag3qHpUHvSorcJ/xXXI2r
5UpXmEiWN9bff//d/WbPznBkRzB5WDKY4sKWZmLWqz7qtKT6cIR+2wWFWAulTsd4
sovYMrEuy76C1aJvWuI4wtxQRG+BiGBv7cLdc1DDpBjayGW9nhLzrQXq9isuLRCk
TvKDfgePBZEMe78fGlvKWcDIMAy7SJxyJZ5yHdyZhjIti4nbwQgpHMZKJtCfI0N5
7Jz6TkxfUXXbmrJ09AQQKJgoEBtQlVa0URiWMqOduD4yL/eP6OexFUsCGIqihnlV
oL1gL9sMcbIhtu9KUcDCVWwxhX9tBiJ9aloHfmaBNfDb7YKYNIrKO4Km/OgfKnWE
f+472Ynbri4dA1KtgaHYTyejSiUVLAI7xwGEEOSJb5IHqFW0XHG1HbGenjx3YPPz
Ssec3NHvWYYqXgl7y6mzzHafv5LNFM3aRTzRNtcC4g9woxfZCMsR6c0iX9VHkNrL
nK+5QuCYmVWWggIxnh+S5TxXonLiv3ddmbQKP1tinzVIgExchHydp51/KbXESIUA
HLUwoaNzKqaJks/wTfsP7OxJqvwE+YOQ54loBwHZg1zU0uOOXr0b70BvvsfuiY7B
dJWzD0qFIwYyh7OZvrjNK8dbjELCUmmHSgUM0JvfMVZOZQc2ov8kn1hlw0myp/N2
pRc1LVoqvZ8JEupANVpO1ko7aaPPPzaeL3IAyALQ2pt3BWjENH4kqGjmnueRCp38
7AiUs+6hvUcpSKibG4hTST/QFl9ZT7uA7hcgFZ3EKOmc6a6O95RIgUn1TitmXjUI
YuDEuTl5MuGDnpxesw33FHipQfuiDHEc5+BGRxi0KFJv+RtNb3a377N/GC6reEL9
7JwEYZjCecGJjvG4BovuMXBQSAy7XuajBV9o4Y7pt46SM/YZHSYRHOtr29+G0gcr
2OfhunnqWOg+MOnDsEDgXT8/ehgD/xOjwfxxyHe+1N/e92R05gr1dwr8K9KuiTyl
iHcVhFmLXkSXp1xfDxrEQaPmteE6KpC9WS1FYBCbe/8H5B+k2m93iV0ui6HGVVEf
FuWwMZf9eeKV5mx7TGNzXRN80gcz2QLD7zidIQ/0XwQdjXG9X5VJ4J9AZ6CBAMyR
z20+fxRKhJmxxZTU9qAeZBKIUNzgkdoOQSq4r9FSFbOkdKRCf09PNldXLNsmJfbS
X3Virog7QS+4g8uq0/3VEBGsqBujtbFVA+zS9UPtknxDAV+XZ65R3PqUoB+oRKMC
trzPHCMbX8APgqTSoD5xVG6DH1g25epTQ+KivNlB5q08iGVhZY/Qia32rFy5GM85
H1EtZ79v8+Si0oWz6OloHz8DbSBOWjCtWIcorHaoHIGJf8guuujcV07zrnNAmyu9
hOXLRgrAlMnKsnzo87uR+WcMFEq8LPAPtKglTyqoq2Dk1GHsK6iEwRqQSk08GdCg
TvpoS6ZbE6gadGINbhfvkrmQvFzR5+WQHVkk2mXsbYX9d8Am8TQf7ryXrGmQMsaG
qVvSEEi0EJ5D6RfHnHUk71hQmale6tV5cSXW8vMcW5JFgUhUYWn6kU0CV5THe+vb
oemDT4WRlp0kT2MTdyOoKlEB1KoFHz1PCHH+dap5sO74iVSGJL/f4lO4PHneqDz2
c4ojcUj+QCQDN4vqL8/a0fB44p045DxZag/hBTnynDym5La3N/DgLJIHkhzSqR0z
4F2okRv0Ed2AShFhMeOyyAc6vburP2QvsgzwdW0kFDlhG6h3n9ToHolHCRlvpG9a
UmDzWV8qA7in+0eMXzxWW25Z8uMmXUOAIt8kygiajs8fyecvUhHESrEo4GHwo941
MGL+IrEsbMXvpX1NK7elBGParKEG04t1j9wOeogZZyOK8JI0eSnovdoUwan9tmQR
92ueKUcdoe9X5IVoQKOPOFd8wqkKsQKJ7KZKLm7djM4bKdq6AYGcaADcirPSn7Xw
WayzIZvsEvEsmB4Cz3YawCTG05O2BaWENaZD65UY1A5TSyJBQsR5zaMORNr53L21
7VLQmyXc/T8sN5CG3sBm5OxeU/vJPOvJd/7bvQwamNfBxUM+bCc8pg2BdpOj4m4A
exYq+JKERf67F3OkyTa5bvoiOOcV92pdFFsevb59iqyNfz7kdp+gbTmvbdkQUPuY
Xbkh6FVxF04nsEOK5sOpwZqncIAOtiwkPU+rLcYAG1a8nfHlJB8pX6X5dWd/sOVi
QPh6H1E1xWzsonF9JiF/QGmE/Z9V5i3qlblxYKDQLvgBbqtwJKYm/LTogMC0eY+Y
zcveGDRgqheVeSFRN7yJnwR/LkkSjDfgLULwr0bpsnuZZNORlOKt6JL08wbmNAjw
9+xgKHWr9SNO66lZ5IDe2wpP1pzff3uH0f/WC/V7MZrOeVsqL1qgGTFppuS2PUro
jwthbXMficuPXBcKHuyhAc65H7dzlivOVgc3Pxtd+8lglh2VJY401in5Wliu9zrO
sWzp+aZYnF4wPnFkmoIN95jWN2xx4n7Tfj3gIZPRl1UfdKka1HoiXa9CmhQWT2o4
/DpBiPk/C8uztGR6HeT1N4ceSI8PCMfcpsupvw6ZoW4gHU3rwbP8ZecEM0sqmAfs
H+mfkTkD4firHq+SyiHIq2TgATb95WJU+qj2VkD5u+Oe1TOc3DcuiJNnxVtf0fhl
4zJWAyzUoCuSZXacEPzhAfgWVUyjN/QkjM5DUhSEVGAcjPRblwyLSTvRf7rtAIbJ
XbvVMCwhF0ENwTKyj191wBCgIyY5xf/S8e/S9dqPMjvYafXKg1Rr2GNqVEeSWqps
R1ntoQxZn/JP1oj+5pOjfKJ9P+q4cp7FlnDpSPfSZjsYw4NZ1M1zEPh5U/r5ZVyk
AGaklMRfYtg1gYxtxLMNyDXCdx+h89xXd3AO95XIRBuxog4fSRKK3+QGxb3NbxbI
HSNjwPFUiGjgq7P9OBrGzTLWxqQPKToUWiO2IMNVPq8T2mxM595HAHIqmeHKWntV
IfUBrTW9tXoHv5aQijKXxtFXS4JS6OoWH5hHmFviGMEp4HGhoaPx7tqpn8aRoGu2
ti4QfU2LjeslB8PDA0n4F7rlIZe+wZzS6kiKMEo1Ix9ch3pozp8zXnrtpq/d+KR5
qrtCCMM1lE9hY/Cp7zKAnTxNehPzRl7twpULrjtY4Nen9eS64hCvmwAOZYnosadu
1smXdI1btkKy+HkZu3dYEYY8xahwNLOq7mawgdKiK7Ct0ILocaUq8kICNVhA+QIi
7f3OgkrbdqDVOsrE4uHGRI9M7qVmWjQKYHKPVCkE5a8kEy5bQ/PHzrjkh2DWOFdB
vQglIql6cOMFEsy1h5glHX9lI22xO/Un9MTSz7UmPGWCOcewKv61GypBuqzJtvtH
TVZbm78N5VLeLkakTQD3fSs2I1LyRv6vPKCpBFX0H1GD1ao4G7heZ0jyI4UrMytk
5dBLroc1dlf+wqC5gjyfsjKOH9enLYgWlCQU7DQP0H4+q2FUT4hP0z7defsk00jM
DmDGL7VDY/jfc9oIQ3jXDk7k9pXrPQ1EFpNQBeZELbvdhTZ76sHcXaTFS5i72gSa
/lTjDv3lqXydYke6+JfbUYGhUDrgi0bTw2rfoDGY4gUVP5l74RhBy5ZNw12xN802
OrS/QqTzPuXCGCFnSyeg33mxnLgwKcswwNAylK+F9RX3OlgokR9RBMCa8wDKdgNt
E2X/brQzLoWYcHj49Nth66pnnhNGldmY0xZzZKpX9S58RlCMN6C2mMRfqRYR4dh+
pQqy+c1DIFcZSotnCTK/BMALZSZlJ7SOGL/Jefff/NMDbOuaO8Mtyd6uESMk3e5z
Y0+e3QSs26CWfz0ErcTnZtMEODhqVHPF4ROseoKngcD/YCBABXaPg4cPaue2btLl
ck2S6YalM7wT5RgqZgoT7wEGJsu8DX2V0aGZqjgMLVQZw58jzjKc1dw1VT6GDhKY
xjINDwswZtH4MrX/OGmyelNuR9nZrf+C0f7ucd536FEG/d5KWZYtXQl6Zi6nx9v9
EZ4uEyZfv0Xyh1WKsFJQwpEUSAwrOgw3zhPDd6VpiWmwWKPg9vmU/crCrFV9BWQk
O/5dy76V51KhyjzVgnpEZLk5L+OrDFFeFeOFiQ84VOsQrADgDGp3utboihrVvK18
PBqD2uD9kLUBM0PXpMFEpMEQ7iJe9OkIuwvNazkeXKoaK/EkGGFNNv1v4TN3Uhh5
s4iC/VlkfM4XPXMc9mCgiklak80h8o/1YVNrPvRrdgu9wo2QS+g7aWX8CnzpC65m
jCbzSf2kG3LO9iinNX9fB1NVq6ELSJfO8QK6UJtAdx9p1B7wPm5xX1YvUSQVzvQ+
WH82lPoNFSCCYX7AUtUZ9qo5/lqUGVywRbY+fUnnw+lQ8HkBYwOsbNKXxxYOardd
i1JupOJJuvglWGQWFhDXI4zu/OFbqdQaxJwnRduXWgbyC+V6IYQws2EpC4Hc6Iof
MBhWKF20BODRJxvniPhHM6Y19w6VzTIdb6M5LuY/qDtwLtaZDB65LfZHuAV5DB7w
VUUC02oJYmMqEKZlttj153DAt2BWK6LeYLCr7lWSi1aisTpn6hbdJbH8Ukmul7eN
G0cX4Yr04+fgW2JHzPRBBTcD6LvwI3pjK54vwznitVfvGRbjJkQWq28gxpuDf+dr
kq8t31sbaCmoCyCdOkU+2XOBwNXenQfGmnrI9OjI8+PQczo6OLgsfq7YutRI6qlC
EzBO0RHJBDZTafkuagCnS6SqgrB1rEL/PRiq5mAWpF0wHSA0vevQcOQKcI+1ouQi
TCLwIPJrUrKOQs9UxluFEK2ZneBdyjwB3fPTGENC4f0sSAy9jisB0/FYZ3GoN5gj
UXwClXsq0OqAyGlFCrZtOg4VbMhH6dWPXUoIYbwwiBZEUPLPc023249xZ1sQFKPV
/kXMsode0HHZdXKAVuam4ax5IxEE8mAT4GCtAnOgVKGDRW9NnSKIw6HFUAhawHbl
IRtQjZOr7kY5wS2q96EvEXbQ7RZ+0Sgy8JknbY8t7QYpjb7legP1FcEcfVDqJAjr
pNp0QGPOwix8ArmwjIFopL3bDyHFfU9cvhey6B5xBJ3xfI96Fyak52UJutZGpLi5
tDixxSSiJQKRz179wYeVhs3nyqAV98vmQ7tq6j8g+IpsWdrHnYgDINCPDfVETCyE
WyW5//RZeew2tDwWzlSRZPzu6FS1SAz58kTRaZIMWNOm7Oc5K42WF2/3GwwEVSj9
iSNZiPWVe2UJHBvA6C6WTjiCldXV1y+E8uHZF2bDvEBDIMBXyUISpaSN0/xOA4hv
Yqu7OfLT9C4fV68qIifgTPq1BJvfRiamJBBAGuDrC75Vk2G/HGZIASY1rRh2oraQ
g9YQGEhqDPP34rER5VvwYdyfNL+Fj4pAd5yfQJViwm1rgnb1UOOrux8yYPH65+PL
GIzaxOEEpKI7TPSmnMtpPTRKlwNuwUXMYh34I6R/U3MGjgRUCPiZmkCkIQg3Sl4v
fQj7OopT6IeAfIiE8WuO5t8npPuWOinf9Z7oCr+Bdd3GFBMg3iqNemickdSFjCdc
6BmwhgYpZIofUDfccRtBlyMsqfi+TQQVxWBJ1iAbBXzF8l4/fgFK5Qe3pGSt3hSz
7mN38Y8vPioPfB3smApuTz/w7CfELRP/IIIhtktB2c8dfz/IhQKwsdnORKx3ZTzy
HynFtxsPrmrxl4mSnqr3I3WYGdJfo9eYp3PW22VyJ/fM8FGj8BFmjkTToXpQFfB3
x2mqvnThlVBCh9QQSeHPCrpM0oo5lO6BlSKqMImpp7hSqvqeyI5jTlTwcfF3NP2S
uJOoJqSHbVaWgiekzS8Itls7yKy6Bh9Zu3Qe1UwL9O5gEOQkhZg9zaD2fS04cDPa
uf9E7WSmA4+FGNTchOKtPKdyWBPflk05wgHGV/Ys2DC/X2Zw5LKoWBt31RtGWTHY
ztyR7XonqvrE8mOPF+zTd+yR2eNMuL02A4BFn5XDuhVcnfsijLUWf9UJURYCMGLC
LagOlujT02huYLP9UNTFUTfvvB4hwpZ0TjdAbozSUoHZ5T85O2hSyGtzOvy3oM2r
yee6GZn5USNhdOXLumq/0hr3YBsfIJy4mbzPKh7Lx7NVx19xpYnwDq98dyZvZS2h
598Ma0prXnkAG8t7dNcuAEzkgWzVfYzz6FznKcYC3PY2KhPpq/VSqnbWpfqajROr
Kii7ziK9Nq9eh9SXcpB/HPw9rpXIYehaimYcVs0GYQt/+KzOd4yVitzHSX+rWNUm
cOuZzYaKzqtYpmeKYl50olxu8pOkO0lstFP3zSAvyXigcbO7d+M9lja4RqQ8eiUo
453A+UIMhOwE3k53IGa/hABi4fP9KSjcymSHpfT/pX7xnsOleE7Lx+JZ+efUebeL
hOVld0pdl0t+YwprRZcj/ixemXIjmq+VDy0ghRJYEsSfyhOGUDlDX41dQCwyNOqM
+M40xHOVYcIQxcI5UrcutbVMu6xHsz76Ndqwtj19dsZGz2ib8/3svwpW89XGkY0A
6F9gBe+5oEoj0UP1UT48+f0VgbSLGautl302O+914W+9VB5W/rehPBDCijHFuMcp
5aMDTtIGZK8LsfYGofRJDC2XIhWGKjpClNeKClV638mLyC+x40/fHnGhgham+re3
UcN3RZRZmwQosd4JGVX78p6Fi/nCQPd+pw3rsALQwYpUGsx2rkA3bwUXpQ6kL8Jt
eR1smBHiNjzqQwsknimTFCRmENTozsFx5kvSXJm2p2hEv4wrCauoTxsJn3Rp4TFZ
liEe56fTD1jvr/I31EC0qC+M8TjCxJEzz5KxtyglTB2xHt5KyPTvWYxCyMGR82Bv
8ZiFlRjUEyT9L2tcl0C75yJRmcUoWE5SOlnCRzbenm97ev+K6Qi8Ax4pOVGDFTPj
S6geTdmC5VlhgIb4mYdtGrquiSn0XFQiFivDCWiCsrtXN/wnJvy5ey+0ZMzyKyuZ
j6DAjOYAgCGtO/BahFkt0q4120rEiuQNNW1vGvMZpljmJW7DPkOJtMZK4a3q0j0G
LndGO9XKp7e1WQWiMnOGtXeFQcR5YW4lSZJtlx1sm7aaIyeC3I6Z2CGgJByU6QLV
svQ6aYIT3ePz6HTLZEyUrlxXjInXmakTU7f77I7knjCcJYpYkUqKv/vWYu3pW7x5
a+8hJykMwWtsCq6HH97Kr/vNiLm8KezimmMy1sGyPIlfG6u6wt7+DrYr5hh34/by
9NvmKrUlAIRmw7p19EVE2EIXd7qkYVRX/nany2eEasfgh0n4VzvqU00KsdTRIIun
S1X9udSD5n0fqCTso1uXrIqDoSWKpWHxe6H0RaFFlHu91p7HW61ruWarLKwHQLhw
Vu2cZsN/MZPwxeZDv8vsLpiLeCc3pgIwFAnIWIiDLqzINkz633VC6he/mV/uzVZ4
k0/S5gw+7z2OAHSCT1k43w+AX7mIluXAx5ZzOQA5BSmJRV+iRqns+61eqhKFrP2v
wohBo1BSUmyNNGyrOr4rxGLWd6Ty9to1rZhl+NnVApI88msrB08esnZpCOxmmUsS
/CqX6Qx3OxTEiyEjMnIhm5sHoQ7xQYwinNn78LT/ZQ+VTmypSHaNMAqa2ihaeOU2
AOpQS8I6SAAv6d5aJ4e4JJhBZjl3c5bPnJycM9bhYrIK+vkjNXaQDInYBbvNm+RU
aBic7uIGlpcWohuoSul3jtA+v87Ly5zmUqE5ks6MNY3AihPr5IXtfItRUkb4ciUg
FWcP/g7xCErsWORdJuNKaFg7cK1j3//S6259O1bbYilAwh7AO8Pp9kHJlMWxKgg9
fWtODI/IuOx/+vrdLSdVhQqAFKS89gAII8Raa+DSHCsE6ELJqQmX/ZsouRANA00g
F+6n+bscKxcpb30NlOCra1Owky/KmSGYyDnCAyV7tNfelIuq3+6B2bfctGiIS3kI
O0Xd7tyESB5GKVnSjByzCnoDVyy66xXVq6C+IX2LmkJgiml5WCJ7AYNTU0tDI9mh
6G3lVBMgbGoO0MQIyFA6E7bX2hE3CpP4ni6WKL0BFV8+0fXFseJ2OFj/Vwl2j6qm
cYzdXQ+fvEaWTcWiovIakyH2lubxvb5f3pccL9bMlZ4/zoB/4urjENB0muumuJND
oA0ZxZ4+2DLX9UO88jauDfwS2w+mTjBNEXlANMQ4Ryaq4C+pQpUo9Wx8sJZSVlcw
MtCkS13UVB5diPSgMNV596OMYw56hw7CEsRyK+grFRhI9oTI0ECAA0sZE5aG1JnA
kti5/urEG7M1MwV7z2Et3FQ40W7fdUEoLdlb5UX4jheAKFu2g+bKA5RxiheeGWAU
a9xtwAXqh8vDP79S15vZnwuOOVTtZJD+Kvb2s5A/5WHom5o+A/mQY6TReuMPSGSK
cGNuZxsBTo6/S5f7iMS3vYaGjOqvPqlR2r5JK+0ZKL3AsdKUMSaEjwfYsLy6Iovn
MINndqbNJKModo7A6QWzKp+ZIgvB//5rETRXdQYzQRra6bQCKdyPwjlWJHUlyTBq
xnVjnHfOJL3sTeNAf7C+0pxb9RGR/qMWcz+ajEytrSXjCpWA9lbuYb/v8MQBSF6e
s2l85TrT0bLZcwJWtHF9CE6RAYK9/SrbRC9JXBeEDBUkMMXW7lxVoiEbGbfIsuQV
QehO380Q6WoiTDTGAopVlvQ6ssW1NaEGAu4mUem6Yoom0ZnSXoBLHpVf16BgxPlM
LE1/YTNXJ0/C3MRoFWF0uW2cXmZtxH6/hdSvXsxZsaNIG0ffU/1aNj2qMpwPSFLj
JhSjez2vwK/fp1ER7+aQqT08nV1x2k0pyZl3po+cpOfDs8iE19fNURHBlPPSq93E
kQ7yoq+SJ1X3dLmeOljevO+btS1SC2BRu+QfBch+w1NZm/EWYb+yZ5BecXjz70Ao
u7VmveMl9Ayh3yA7wS+2YLyyo8nXjM0SpFo5a7IztalxdHyq0N6AC4oUxknw+c2D
zd7dUDOW4GBKtjPg1+9pG0m1NANZUDrChoaP2b4dvBqQAKwAQ1ztMauwp/kwlK+k
4fdtOuS7Zo7H3ObE306ut3k9qO2G3gbeVlgvASsQ55MKn1pwaOivhFBBEGwwAk+Q
gJ8AOc+/njzNz32w6fNWUDaQYx2k+lAEq7pWuOmFaXF15ZCNYQvflpfZioqGFBgM
LY8uvPAqcfWQrbsg0Esl7wlgpttiw2SJcxtKJFF45SmZ5zcUYss5x7Iwe5Y8dgJv
BSIVtfu+e386KSGUy8cS1vg3/MY0E2vvcm1wh8TnQ20Ydk3oQqCV/t9Pn7NRBhKq
tVhaJDRkb+9ajLqfgsk2dbQXzttyYedL7ntrvYs2c224NiHXgSr3NZFTxgxzV9bk
m7GCNQRV8UeArzuMNdhoCu6hDx/G1/GWctHn9yeeASptCgOD7sfpHYKhPBKD7i/N
x+3Z2/25SoGAsq2OreHFWTzDZd0a18u2MiyJ/7yTQSUsH/lohnRyY7ZG2tan3Hgs
7rTf7fPm67fdILdoE+rEMCCQRaATrMRMiljrS0VuZbT9uaIFmLG1mCKJxZcdX4vG
rNiY9wvVQqNf2qEXczaoTm0KO65jaUHEzKGzTlqPm0gUxFLVorr6Cp9biAG7zFgf
XmNsyGjv+YwG+QB0Wyp5eU3ag559H4beaoGZuc8US001YJNzeMqsYfNr6gAcUegQ
eoZ/2TcG/PseQWl7CYZrNehNiZnhH4Js6UyUcmfxfzwjHk6GAkqfpkUvCJAxy5K5
d1mR9Gt+TYPtP5bhhBuJ4NjG6VpnOch4KA2B4X7QARfD2SW7TLkECQVyML3TCJFR
/tg6bTTaGqlkBYHxpRfGKR0kMiaU6dY1lXdV9FT7+JMIDv2EKXf6tqW/RdIZwvHn
qTTIlr1IY7wPBpOjYcQWha5tK9vZgw7iZyVbmWUQ62TsWQItyK3NT5GjAnfDRPjI
ut9L5h/cd2bFWVK568FWh63qFr2l3LQtr+298Ucy4Nkf1R/GoXw/XnKdEbE7DPcC
Viw6J+n08j9CMR7o43ICs13sM2xQ/KEBBw5PGnd11umy0O8xyEpZYrtdO2YfMOfb
1lNE1/Z36vORaUnagD4Nwrjdj3oU+4SJSbNPp0xaANwaqVPW+3vONutyMuOPrGcV
hGmD25pyJ+Y45K0mZXFQyRez5/c12xVQAUZBN0j3zK9DRx8VskBZXYh44b4twEBo
yNx/51TYdZfJ5F7bc678N97CPdqrQeQHp5vtdsNybfbBDlvjplF1AvTdLryHHoZz
1XMU5hjgfPpe6+AD431KlDxqAq76W68QwKtbFWphANI+928hViXRhxDVCzsuVZF5
OTPSvbghM2iAMtMKk1zkKexVPlRoBgaRFNYA+Xa4LbK4mYSSd6lgSpUEb5v8PE7k
i/JzYbNj7GDzB4uj4dOMI+CntqJxXQJCnSMVdWQ/MPuGvCcyNXavISK8h0QIr5ko
uDGPeCrPfIUI4dIUolAqA1WThyejxehdyJth88qS7PvU/Ehg0bRl7jgOnZh59sJr
tGNdnPhXpzFDAgjyzskPkeG9Ns56Oz6rG4gS85+/pCkshS9BRFQRt9PFsb6TcR55
r7fsPvJWsVTwvgqo82fzhdsE6lcBf2GaW89tdbQX96ksd86naDFZ4Hla9qmC7/oM
T8HTYfufnBmID4GLrLRAMp7DIrhqWucQB6BBkvdZ0sMEH9ZbOC/eakj+/XjZioJL
SVDTbwTI12YNalwoAQE+ue7+CPO9ULJnjij8eli329lItXXvhEaekh9l4XuEiHIN
6tO9v702ieo3JJbkQxgme3H7LoXDGprZGHg9QPVxEy0IsY7V55kkPFBI0zqkwO8A
4X+OrMpKqJZyu2R3Tj9o03ME3wYfFfK/lHlFy0lpxsUjF6u6QSLXJuYP79QcE+wd
x0DNm1+Z64DycsrNKfr4UbJQsLvMve6+cK7hcwbMS7M64aGO70mE1xyoWRSYuouW
H1HdPbDDfF+mg5jmSzsKg4Axevv8TVhrIj1grx+pH/nvojTjh+c2H9+8dbEnKrI1
+mqy5LZCDklnTYkkRhcVojFo6Fo6u3jsQAbdepr47NUnbj90BuH2bV4iY/uO3n1G
qtX2nvVx/TKZHRHc0pjkU9lzr6DTZLtUEAceYMNwgSQAKZNzRKcrke/90fmXg36u
ACQokv8WWYTNGVRVv2EbSrxuG2xNBQrjg8RSpDZUZg0uSBZF82TWAzophKqsJxuX
7AnlyxMdIfPvzcv71NDdjGiyuGjbZp7Z+SqXX6zRpzYWRlubLUbIqxa0p/Sak2Mq
qVQpaFXR8nKyPrEfmF/pguGTeEC51uDmSEfifbKZAV2ceuin4vLaRyht7ux9KRwC
bQL0VV4hO5+p0r4PCg6/oBOzpcTzggQnUVOPZ5rJ1FkiKjpQU+xA9wHfVAseoXdC
NQXj/b4ZEu780JFOB1O4WpKU4h61KBBc2hLq3XGVvpyiMGjwnFmcPeUU/i6XZiEo
2TaWcvW9k2/n8j5d0E1WrYfS5zbYRzYoguFx0PzXkCR0mVx/do0C60tcBOGMN98i
dvgDiEec7TTGPUiv3z3gK/c1A7UQVn/psDr1x1EctaFqzkilzdIELnVR1BCsX9LY
JoYoXcGuvgvUaEy8kcrDzXPjJvDNrPMaNJzhaEyA4XvA495Lg+5L+LbMKiLe8FVA
uW2bNsgo+0ZBg+beCHSokUQHV57jVhde95PROghlWoQTHeG+lUs08IfNMN+HBRuV
H5JZ4THhF03L2Us7N5Y/dRc2YGupZwJYRYSlPWhgOMOzxd/GCdXDoEcUtesueS5p
aOI/i5j5TTjLtrdKbA4MWY1FMknK0Dmmipje7SULMuXXEPgIL0AuKZMY2cVfxTvh
dJui/Tx9nex/46gk0qL5Pu7wQ3Js3mw8LjMb8PBfxMTKX32RvWUWPXv6mxM9J0UC
W4g9TlsfDhWsOO1dirwZXQKL2pLt+1ggZ/7iu4svoeQTQHBc4I+OE0BgQJFY5nnF
/yPyhY6o1MQY9race7m1V+fpzkPNVPdVLOLfLrxHdHgpm1MzdikCvr/ClFbj4ENr
Uq73W4+lkpN/yCifamquy13KKYB6fr3IUJEXlSxhU70d7yZg68H1OIOHWFbmioLz
KgHryE8nHGYqC9NSCqYHxjaYiXASh/Aox6gLfB6uTKB0pdqESN7lkqjPbyEpSXsr
h95XSIi/jA+X2Sr5BAPYwx/RrmURP5dHF/+1XjQxegQeNaEci54UcrCmglcE8ZTq
xstzGZFdJhfNTVGnP7M5/h42nxQBqN5u0TGRhnlAtqSC0LpVYoDEgXQZ2605Hs5K
8NlArEWfEBbLOv3Y6J3cUlsh9t/8N4Y/Kt0tQI7tJuY/KUF45mQYL14DnLMWhxOU
9ubYMB2Xsm/tx4QqaLxf0M/Z73Vh43/uBRXvmuupOm4V5pKA1Rhhz0fLTjDmj2ky
8t0DF2Xbjkh/Fl/OZB4KR8bMhbl0yJ0Q6CPUVJaCU3Nu7oda+h8sDpRFGq3kKorh
6oWeTLygzqxonCZpgFE/QVZVJ97+hRlGq5j00CGV27FNeLD0RLuamRHbmZ2qvenG
4tKh5mM1jh1772oF5v2HtJZwW+6wBHAUI1sIlA6rC24yZafkCAAsZvkxWvKXve2Z
zGifZwTow//99f0rjtE96vuGznj/gxGQ+MG35/4LFPLTm6y56JI/AwVoveqlD84w
c8ULHA9bdL1h53DgoTA6yHScnMTs4vzulfl+TvkgMdQaa2MIQWuhrLeA49c8AZEy
/nZWt9son+nSn3MnAQR/Lqq61UmYjhOs8dZ/TIeA4JhecshTR9xKkMIh7ieP6Izk
4OKVa3buxOYkuLhtuelSf598Cbo6K6e8Vc9rkrml5TE+ngqTkm4khwxuaueaFGrh
mC0MF719TgnzO6ZiUzItoM8t9kwRoIoNyKBvYLkySkKcICFew9RzpP/3zLMC+hdY
nBJYwkYA8RbzCfovMsySX5Z+4O2QN+17UG4xxnJr9EoAeImGdyWV1pUF9UxUbsqY
OlPv5NO4u3yP8LnOu1NBfWHoGdyep1IM+PxxziDfYgcYwaDamRH5hhPIqeCnnnEN
NAFcevJLxPEggnjU1VXgIqEAFQ/rqwmFPMKFvu/sWLLW2Is3gwpTkuDq3VL/kZZg
58aujnNMrN0fkO/cpgrvKjHeTPe54XzNdkShJSAsXitOltLDscShuc/cX3TUTvK5
14qiZ78FjBSmDqrS12ejM2EpWUe6OhFi1b/mompegvcrR5c9d5RhQoYsjvujbdJ1
zem83j217HiyLkaYNGzCkwRrSCaesNnD2ZEKoiwKApKAV5JpqrZv6vuhmIC+BK+O
ru/Hudc78MyEYmNqTRAYypguyyihy3Ka4RsejlvVvztFb9baKvNB7s0VdCP/r+9d
NwT6691YAvGJhVOcMOsugIwp3W4R6I1I3aPzuik1/JHkQxPWQFTvhsms4XeAi84r
ZGMOHY2qjOPBUSD8PwFea9wtIPZHHB9zJHAnrs6kb5RLChGpcSfurNk8iN55qeFc
N4nNfewwXoOwXLCN47mR4/BhK8dPMWh/RBANI9fIP0eFMsgNS6oe4bGirEruZQrn
dHQcGXbOy/NuF6+s1pBmE92CkY7K7H8lsnBKXd+jjaxY6WPlvNSGtr484nnW084Q
tNYFAngiJNONmh3qQz34O/GSPzzbmR+rEvRV5hlskFLng3RdLZnPCEtHiEa6ImWQ
XMiCK4kkppVo7E69a6IN3mSIdiUTCjt2RODwyXKQs24DiiKSAr7KDHfB4uGvEdAg
Y+yFCpHm1KKfSPKWLWtb4XDIA5MlhhsztHw+FIw4Na5ECJOu2xDBFrSogEhLGaX6
4334lontHsqS1qldNGLiFxTPqU47cdeUAE3IXnlwao5/xh0l5RUdCm3KNV/2TXMJ
klozvU9IlEoi5Gdoyq+Csn0xgfU/tccaGGb2u0t4+a6fpS1/D1UwSVxNP0ZcpUb8
r+JaBlSxG2N3HtJ8MMpJTsft8/Cf5Z6HOBenss0Aj7SpQUJXS5V3fh1VPRCYik0c
UV17MiI/r+7zj8BUZiohUs7o4bnEqnZGjr5PILWCZsytTaPVAPHeKwP8vbfR3Mw7
bH9PvmCj8ffTXkYWK17O/ehEit5+nw7K1fvmYn0UwwHC1FEYNCvWs4PnQWfkRx0P
cCIgJrd9U9L0fAhy8DeFKeUW7ONNIMWY21UKHHO0/cjiJaT+p1MYFSFWS/Q8xOpH
Gz8dNtUt3qrM9oGKQNz2pYh25gQnnLfFIu7Lsrewxl9YJpf2OXONLvbKWgDnPop9
Uyd646QHVh9Ou9cNt60fokq39CDOLhFX2YUcmd9dL8mpz8RKqGa59QUZEOKyXOTB
wJlGL7USnFRb4k73oqv3azvw1rSpuaQLANhcoxrTm7NlY7/usx1AX9cEfDJcfzZM
XAN3pKLp+DP1ZQZJeFNoqCfBaAafvDWWoPHmQkF8z1QiBA0GhZfbGuAC0BROtTFH
0dycXImVWuX35dzEUvG4w0mLR7IVi8zKtVCEWv4/EjOuWlwPdHWbLA21AIj1LZlw
Fxio7t0Zhz9S3W2KRsxzsf2hyp+ikVQNKgnyyt513a2b6+qoJggOO54n0C8gHGCw
PCQI/B/D8WtJDnEd1bhGkvoKtYM1nCqsP4hsDrSj2PgB//YsZqA3wxd+NJbgWWIa
Lnf2n0bzHUEJCXunBm+hWrbfqGIxvrWxGlZqGP9k/0Uc610HerWJtJ+vBumpOOP5
Cma7dPk3zdz7LPd+YFkpnwGnJ45pEN/wcSPolWFRyd7sm4VltcU2coHMNCSDY48N
8iV3Ud+Azv1F+E58Zo6TINfZEk7KvFxN+yFpirkMKiDmvEiZVIdQm/k0V7QJVWqX
5uAXHrXCVP/EoMgBUNu5O5w4q62ge3xUwney0IjxYmYtwLjgZ7/jrUB7Y5OKnXXn
i5SGt+IpYvtFGPPZ8EDeCt9l+P7OTPnKvVC14iTiBaNwvIbhIRI0O6cdH1An+pa3
FosCZofSycFe5fDe657NO3f6CeyVkgk8C8iYd+hjzuNSdjvJTkABKj8g9K1bSfeX
A75IXIT01Legx0YgbqkG/5skEx6TN1bFQV/4YpZOeIqSRusESAzJ4DNkizojDa7X
xNv4N+yZuFGKemKxfXf0iNrisYkTecPOnkpv6ySq7tPy/BRxhViDG2IgwxHqzUXE
OkLftoqWlHs7+d0WTos0o/kQbCpVLsDvFrkdG7e7oUQJW1z6+SxIyp2MVYXxS0fz
ba/GRa3baeSNcilKjRszMzwFLNS+mqGQm8BlZRguDnLCNY1sLJmFn6bjvLoqPePK
VvMRZg6xvqDvoZu4Jj9Sbg4upXqeey+vk3jm4IF7rLOcp78nESiA3s7LCzhnp8Y6
dPycbxc+M1kYyvFL6WU1bnSRbhCWh+6jI8Yg+C5Y72XyyhW7F/GhpxG+WTGLZpzC
3z7XW9iB7UCo4cMF7UXE51bHCaDepz9XO+MMCm5ncRBOYbteXQPznjjwiNf0qCQW
lJb2+7HdWSFaU1qJiOBKwNgBigyyMhNODoXltE6YU8aSuO3Cj2cyGq9zh9fABax7
pTpD1sUMG1A5ZR0pFP1e7sdcUfvx1HNakxWKjifRel+vsoXnPyXjqSWxP/XIUDOH
DSKxVP7JJxZa80QnXEM1/LrK39DOoW3hQl3GW24P0wiJNxqFDY7uhqWRxA8zLXuz
VUG7cjVbSzv6RIaVKldPfJs5oik1PBUWIXMZ9xlDW2QHv52PV+rZHRxBvqQlPtsX
bBmHC1c7UgF6zzAAC0mE8v3gjRaOyVGsiNjCCtbFNMG3zj7ITVTtlhdJCJKj0Rnk
PouLaGj/7ngkOpndTiyF4kNhI3CUNP8yIxdnfAZcKpmFW3SSuEAInKVsgLvuizy4
dnl0J+8Qe2te5CKJqhIwqFGvtv0Sye7bzveGmcMTO5WYIcSjI64Ha9kO3APzemWD
aYefMekESD6jrho3XgAVu+hOWxYdXcYlvk3HttXNam9SG5iKO7cpOMOBR7/pdjcO
znQ/uXuq9tFaUJ8OFAkaVRN9GHuAXcVxik1HoC6KM+ZaNwpgGkw3yrcGgGAWHofK
n2pdonp5YaCF3R+qC/z7u4pcG55Qd8tvDYO4do6b8Yt9O2AR6IsxPKQNoYe/Lm77
Jd37c8jXxkt8Axy4Mh6P8KpXkSbAQ/B9LvZko+EnByFEdP1l1lu9h64ln8dL/vUT
4CirEsHEoX+b4ZnWga+7EigV8LWvGtsjp0wh/Mm0WusoGOqDSkPtM4sFNmUehL9m
hpk2sm7gQqWequLn+BCToDrhns0EtF8bljeQ5P5S4CvXstDpCs0F8E9s3VMzRBPt
6gol4f3k98E2t9RyWi7GJvUNWBo+KpJ9xfkwKiyqQkhgRwoJW8VntcKeoj6syj7H
HY9tWkv0SVgcXG5BX3r/p76MV06toiOHd/MVqO0N9p/ewo6nRv1GFP/PjIPRuKor
0ygWoNqDdwl3jYove5FnH8A/YVf8HAOOQ3hBmFI0mGDQKqJmuH6gOSZJ36y7nASz
iksgGHFJXX5IsE/38QMfmWK/1pP+4XlFqS2Nol2QqRiMc9F5vhSClFOroVoj/shh
sZRRQLZAI1UwKVxU+t1Z/hKPrTGH+8zfniQrfVY12xKqALcZ1aXrZSJ9k0FpFdrq
HvuYm9Byl++apmYkF0/3csx1QYFpdRlWfaJby9lofR4PI935Mo+JRD0rq/GbGRd+
93xs3qN91iCVNeIbD/X+hHAxwaYyp197i7yvrk+lW2oMoljowvBbBN4DucS66FLb
Ev75HmYn5NxekS8asCubmwSJA0f6QE2ivPD2voRgFgZ3ivAyMn1Y52YtQZU/cJ5i
9hZ2r9EzwJYExl0iTaQcEmBYlOkH1viSeeEs9HMWZ2EkJcxE2U1vMLsM1kSLw1nF
8gjVVZ1gFh3ua0O69MqMaTXs4BVIugTulISw44k1xbXg4I2m93V443dYryS1rexp
58BxNr8yGzL/nTiqrW/29pyJAkSQDLbJDI5QwS6LjxkrssLON51H2FhZCV1cwL+E
khf4FA9VSAXI5v5b1cHGH6KODoXLeeDbMwGkz5azRV2XEXaX4FjhUMj1YayFHZVR
t5lhkwgDKkoiDbmmS187xy/0OFMobzrzFhdoyFIlI5dGoowH3hmoMSlvLvJziSRw
O1jj0H4b2vAKdp6kOyf8W+k+/RQFkjnqf4YWHXHrJMB3kuqZpoLuBMl3jrzvljKk
+xEE71IodiKMrDDmWlL8af3+mcV5jVGFIJq9P0ruS9qe3EqdFqTX5vubCBR5qyYb
veus/fvDLyXbkuRWvPPawONPHxWGE9TDHIArD6VI7bZr5Gp8cijmhmUkm/Xpp648
KsyZ7K7+hQ1rBrqM07irrJnYl2n/yMpWV/UGIvgzTbC65pa0DKoDBRLxDcsT8J4v
TucxB3HaavDuOFyxpt3VRlMMYuaUHEmdnX1FEUrfaxnJESqN77FBfPcPdSat6EkM
26UZsJfaoJ0kzQ8P5Ipp313iref7MlEzfqnRB5ERggBeNhhMBJ6is5QhQ7S6vXjX
Bf61iD/McoOAtR6D66Le1ug58y/3dBL7k/1HIOzLvcvqzgcrgZpN5m8ioHX4IdbE
CDKnAZ4xAaqr5mUzoyhuf9ehPpnpk7SsOhR2X1eLZ7ST49TmIiRrPgurlVHW0Ikf
lA0J7ajwXJ8SpSdz60iVcwzWE9EikSq278Ghbms88HoGXFd3UWe7MEN0jTA55ZE6
o//JdC74XB65A/fnRQF7lA10mhXDb/WHvN6/Zov0Az/G5//citTK+dQ/bjDiYAoc
jQhg0YJTPz5wF3bnMw5vZeJEwXn4+CKPISQe6h1aJeT7y4gdETfELSgIMuHsVcDY
9i0C3ActoBjq0XZN/9DFn6Yt89Rjul8VwHxBJBzNErqGEvQ0RJDupgSsq7sW6a3Y
nOIfQ+md1pm+EPu7/FHKswBEfqOYAAV46dgXvA9dfR8X/4FRzvZTcx8YXkXjfv2W
8LS69LojcOhmgAtgCEnJJcoByt8ELJqz9sp94gHkKTGGh2D3LViw1u4bCmCDC/oj
XIzQc6SkhweAp9FEp/SRGtTyhx0/1I0njGMAwuQZvRezdqnWVZVOA8O6N/szM9d5
8t7QNd/3XGNWTuXcdQQ2gkNwAiGnS4Y60bFRb8jlM3VGEvZRTl5AIJI5q5O8xiOL
0BndRNg2uXmz8mkStk7DSDnxufRq6RJDSJrZuIQyttd7cKnltIv4myl+R7+AJdVw
Hw1hrqMxpyo34w3WBQtpM8xfGgpGAFLLSzXvgqiidDw9gtA9aAsGbtmkJ/a2It5Q
JdSkLhUpUsSrnGzeoVTVI4abDojaRJGKP4K8AEd1y0UNA5zXmCBBaBj2GjWsvthO
m3saBZT3be4uldngaDjj32Ocu3aqqO8cHGA+k68xuO7eDp03XunrH52Y7hzYVFsB
/MUxAcrTnolJCtd8DyQEdLjUvjb9nHzE9QQbZu6BrmhcYxxUVJ20fTt51cxdKSJp
aTMn/V4Zn2+fcIY7VgVZE7OvVujAmurWgUcQhxULATVKu0a8Wg248WVF9D7BN/Yk
kMJwTSVZ/rlHGAgN9+sU5PodZkVCLFciSvmgvBXMF8S6Z86fI3iKvpKYkOOwkcMG
Aab2Sj1RYDJfDPdvcUWc5tFw3QmKuTL50zecjtSiXhDaABUrFuAcbRz3PxvRwZGY
tl6BlfkQmVOJq78PaqpzithTUYzKyYvgWIzoPkhBlUBemENyusTbg/mPkuXXdWiw
A3r40dP/6/kQdR+pYx6AhjbdmyjWoBDPIX0pu13jVWOhjTo41R5EGysWuv6ijiJC
l1uU+K/BoLEbY9jbuvmBjwVP2kyvTa/S94ForUhE+dBowZ6MuHeWGzNWVfZI0oSX
SpKo/JSOgOlaM8NWlh0yaR6F0e36lf8NIykrSXgb2sRhWXy8y/7iJAchD23M2fGR
5eBYDhVUHrVmD5z//xftlGKkv+kpCLU3K8TyuXI+IQzaDdsj8AFNt/vKot7ahbDO
b5r43zJHWOAaLUT6ZkrUSpsy/gyupCf5B18ptKc6Mik9Le3VyRmw9tYX0cShmg5A
CdHAOsX3+5CcKnqmEo4FPbaGgkaZ9T9D8kmFmf9FmBe/9fbEiFA8QwwBwm2yGtww
Ge31oGcJNWl983LqPPzB/OaeqtVlgPtiMEp11bMawsHTCkodofxDsczRueNDF89L
YGYCCeaI26marsvPIKQ9/c2FfhhxbGtObJytMeerhWVQqpiyrAE06+xTEZt4hkKG
it6RYf6r7QqukexP2NdecHQ2LLL6yzWd/b/oFuunXRpmzw0+55bId0dAF81ciTWu
LlrRmZyQGpZ7z0PypDiwnfHsSerc4Q6sy/oPmF3T8lACriH2A1u+mIIp+Pbp4kE9
su8vEzHmmigVCrtSjRbmXpo+pFS08CYKPn1Ih9vs7KjoNkvPtIgN8Gz3ejsAsTTg
4YPvyN1bWDvw+kcdtbs5fOLB1Z/ICcysYFEuwr9YESMTAOOQZzuNz2hLc60kvhi4
1pKmc9tWaOr1NmsujweSNDnPM0LLIuaMdeC2lSgbuQDXNuv00yexlH+6Wj5cgYkS
Ah2W3SRDeSCpR1rkDTjGFDReJJmzwPxUrWqzMdUEkX32ag8RESxCSRKqhmbZViZ6
tQxm5JPAhxAmI1UWlsMj+7awYa9QkZlN/m6BqLu4PwG3OaYiQhKm7pmK0oXibNUX
y7zJOIp2XztXNu2iS8+zb3MO4NxYsKoVeDdIPpHTRtO+rBMBDiwY7QhLjR724D0L
S7lvAR4nufgudxZJlTXdrpHIbNRnEfZi0TguZCXlqqHdJKwIER9q/3//GC6Bqmzy
PgIJAFjdXhiI9KQXxnwFfcztNkuCzojrRIV2qkmm17DIobLFzFzcu087N4Bk/fBw
XQdLBYqGluG+VvQ9So22m6Bl7szaM3nfeImKYvyT3ioQHOftvjWT71Q/L0kPZm1H
dhp7lwLVyN0cHvZLPcuCifvgumcTQoi5/H/LKEDgXyH8ovWVa5DJn54iVC/n5Yts
dJsgOaYszdx2ZlixvaMcd5CyD7sxJ45hV/nJPC0FRHPObdr6h0Zn7lWugrqtk6R6
HVmMMn6g6nQfpTUUXwN8tZPlj0bKkn9kDLeBbu/Om7yqgtJfy5GWTSmsECiJbISD
BOwd4dTn9Rlns3rfa7JxbOTMFnNUKtyq08KtICzFGV4uiwQMI1+Npc7wFseEKz6J
qlXA1FN2tv3GxpN37/RiyBI0LHHtsdSHr/FTT4qNyvYvW8br4mTQGo7/QYpr5TnF
FuT8KsFDLX41wbVa427FcaJgiyXnTipcyrQwGzHXfRDUE+bue6j9a+VKMfcvesxJ
1YNzRLUoCzxN/yu0oGYyKyVB3/CX2ZiFSEcp/5pN313KnlIclPZXs3Dynh8c+9TT
p1JMAyIph9LT/2/Z0XnR9WgnpjHRL5grdVWFmOYBiEegi70cG/5jF7BJvvuzhn4D
Czv2CFy8GO4nyOu/os6ngoPBj76QB63YQK6KjF3aU9Xfmvpc2oqzv/yzoUC/7haB
74r0FnE0RRKteDwwTVCuoM3x3GyMIA36X4ndoF3CM2Lr9V0uRl0jcnOKzZUm8oWW
Wd8/OZgKWIHDLA95eomTknjIfMyDBHJOq15DMspFTCx8ycZLSLRbnmFTJgPc9guU
hkebG2JTzwrSXW+ruJ/oZzkaiGK44LpdkLtZopJbIH50/udLj0C1urtm2suvX0K4
XpjjgHLwM2e5/O3LM3k5zL6DvRh/gTZv3jDLcetZpQtqo9BeDalpEmavB9Fy6tkC
e+09aWj6wcPKj1vG4NdRf8PWm6yKzyksIYHgtC17CMe8tJPkMdJ5HmAh5H12SDL4
HHxDpaRLC/s9YTi7uitW+KWQK4bA4J3EJBRjhiXgGeM7yJsvQ8xoBCYX/sGMP/8m
IX161ZYORBH/gbhPyjDyZzxS1fR5scEmxSk2vuNlGPnCj899mWnx9R4sqxpoIvq9
O9poVCekHvbXTV5hPwUn6m5wVVC/NtJMR/3dolmM9zTb0UXP6tGesCQU4euuYGDD
HLJojK2sWJkWI/hgOJu3A54JzkvdvBlyJ1TYmg8QLr3gqCrdPXiSGG9ixuMk45Km
F+bPJw5w/0jmClPh4Xo8w4TUbtyDMwEfhPWXQ3bj8Nh9vYdwZHKBM5lOI3q+REDL
5LNz45YUAVVHCvo7DvnqUITsLieXlVs8jXaTGMFAioUyF0ZYl9JUPInZGJhV7J+/
oR2CyhZXofNs2y1kC4mNERAkg5GviTbPcMcX/q72WPZJZflIKoAgBfUtEoYT81iK
WIr/vB3yZqwqUNZcQ/XFpAZNoJCZg5EcaGJeerjxbrf4TP4TiPmNqTASwL94HE9Z
fKKTlO9BSzjvmmNEZ/Uk6dVmKDOmyJAWd/CpiocdU4sU3rS/n1gX6xXcyWXHSXS+
QP6YkH2CgFLtkiAhVXsPGpgRIIftK3wP3XXVvEyJxXPryWJRm/CFgS65LlWCWRCc
QcqmVD1kIRmJQRSzIK9v7wdSXq9c1rzI+FrZ1L4XYeCx0xQFiwqzbPDUca0G0RJY
fhU5yPXBJZ4cnw0LhJNsL2cRs+X9pywIKLC8J1upoRL/LvFgM1Iyd3Zkdc0VCk1D
GCty/m7YzI6PmcZ01azHiG3NmghlLGHZvoRdXisibJSATES51otaUJieHxJ1U1Hd
Wd9jdyb2XZBfxpbCD/zLPfzz6MApoVSrDiNbrTacAPfMKbwhkJUuvnCIqIlZpVws
yv+UYVJoWxqTceTeG9p0hc62B8wNeOqKxNXABcV1iTG6FEA+kiupKqEn1zP2kzLt
YvBhrzQ6bugV5gvy0Mg2+fDEXGj+efflzHoYgvZ/moPf9QtT+AwFBRcq79QPwAUO
dbgVwYbVPOUWM3TFhxQeJpJWsMPynORUBmFvAK/Q4WXfpn7AiHOIiVB4hjFZdjME
nQhUw931uHeYLbs1yhSrf9OZacv/U3RY5CTM6qCPXPoS5vT0+zG5DHhP23aeVdEr
8nfMWreBQTqvRNl9INGDnM/qn5seG8mapfNaMtgc3WP8GhHn5hGdjy9Wbs09gC1R
jEJdLWiCTzRzzvGuItIoBhg4uLzz+NhkL+dZr7q0Wxl899GXugPb7n8+W+z3RZSv
XaVU2jWlO7+Gc9yObbpsIOoWqBZIGqe9DvSWlNwSz9YK53PDQUE8D811TkXWXYq1
Ykau0/fe9wiOBOd9iQZGFu1qV5M49Ii8ap+2CuCrzamihikJ3OEZK8UeGF5wj3FM
BuGkuxM1KMWMPGTt43zHO66Df8z1kclnMFgZgZ89dEshpCaVj9T9ZcVYiV++0sey
GhRBqngH2Z9pqo0P/cOf1EPK62J5JQPwq5yhZcutbZLUf1pe6OdtCxjACTgSTKSG
gZv99uMAXeqsdZ5J6ZM5UaRbZfBTlRVWY2eTRsa75AGBfaG7KNlOCOkBCWKmLruw
3SRchoHIIJGwTnL69/vNtVlSn9FLUs6BygKVTgNgLT0b66Urf3mPnCWQozudn7Fc
jQUDW47yKQnsjdg9aZH73xq4jHMZLjretnfEF5/oTPmJ6UciD8eCCN/FBHmNLCMx
Jrs1/auRMqy2jLkM74efQTNulyX/WLhJfxvG79y57h1ZmteLp4qw0XNJYpcysiqp
0dF+wlMOFeimxdUjVku9XArm9yfeMpTIaLpNuH2jIZ37OOTUOqENyeuPU3Wyh6Eu
OpRAji5+MFrZKKs5k9G/X8vd3kFcsUXjF8rl2WBmOOJ8UQ2clQr1wPGA8tJr0doS
6cIQ3I6E0Ro5n5ycBsMzrXiiAzoRfh5W33N59RFWCSTm+ZZHkl+ENoubDU53fk3g
PSz5CEvyPV1tfQZZ0PfXIWh0H8feQTUdM0I6+9qcMQrY1SRqbWujVtnrCRcqNLwY
ySD18qEflng7jV3km2lrql38ubPyburGduM+UothPJoli9jyJ7fH2NThPNA2HUnn
Hg7p7sA+sXU6kJPj5HRiiPh+6mDnExc2+XL2T2Nce3x0polQojvVim6p48zFMo68
SFE2QqXtWCxhY2s0+NRovDhITZV3lzczADI6x4yb1D4ObVqCduwer3Rb3NcasWRI
m9bU2Kaxbm83JkM5XT8rmmd1gbchCFMbV+TDO2GpkE4Lre0VzG5s1+ZsMCCZJnEM
G5acWFvV9RbhMdsyPKHfAZp0Tt0orE8S34eb+pH1ELrBTEl9NUFPBloi7Comnfjd
QGhOOcbjQOM9SGQMIeqVZn9irxMveSxwyxIEjWu58VvcAcg0IKzfrSk4GFUGlpC1
BjcNzJASqqjURgUsT2+UKvvkJFGI1tqr2DpaUCkafwGi/QIMTgNCzZmHz+z/3PrZ
4EbisVg2kqSNvdP83u+rHXtlnEgjXiaXvzqY2rd2Zyc7q3l4insCiiLUv7glLTOe
UqpPLAjmlOXKmzk7Am5FKBw8EdVhQHbGf+AGbA1UbTLFiAYfvITVpNAIZ2YJTQzO
8MrHwnGzHWw8y+seTzLM2bKZNuAWcLWESlwCe+rL2O1NZugR3XNr0gezvGSYJjip
Pd++ZRI+VvWpBcjac0W1jDEUCXyyhAUjkGKD04yTuRi/bp4tk1TGvJgkEmITidAw
Ae8+I8z/Cw7jLafroH+Taf1WrykGP0xkFh8YG1OIOoO1l8P34+wC9XK7JXAd1gHc
cANGSx+0nagMUol64XBHOXlS9LgToQXhHewMjo16ahOvDOesCU+6yiXP7rapd6hI
B7cLFHvbdaUUFEb+omvgWZvVZK/k7Bi4vl+EkNQhOOexkcfY3mst5rzTA7zbTDeS
eTm2mijspmer6dWXEGnZjfGIOOl/2mst2Dy/c5kVbw/63wzum1tR3XCE8OteMEvT
/WFRWESD+YMs3uc7hO7XjWbrFUE7y+u6G1LBAnv5BtAInAH5LzzqDfCepEUWFZQE
03QuFFSjWC4nGVJSgJJKfJL9FKxuv0NgtS/R61suJOjepSS60FVxqEUaSd+ogNiz
KQfG7/j4RgcRPRcxssb+8lvUXW4jmYXm5PYrJ5GsAnl5S0PenaX6VHSw5ghQzFuH
YnAOChryGYyNIaDIbMHN34E/lRlP2Skh+qqwwf8vBrcpiYTSXHooFYPNKKZ9GIgI
oJSDPpoX/eJz7q4RqryWJVeDD0w3TMJ2vIYjGs71eKwRXySU4Xn/y5rNFYwEkZAh
Lktp2jiY0jbJs2dY/zGzu20it93gpjT0dkOjouA882XZ+LDbmrghqfqJRXKZXOcT
2H/WlOZ6vpiuqozIQtJAZQedT9JciY5ICtV9ImYGzy3pYuNNHo+gLgGAjZ0hGRKN
nQy+Dro85IS8OzLsejiUZ3iePq0/8n24B9hOqdmNPAKZb0+8Lo9ioP8o2k7tLPnT
XWum79DsXGv6p4ttq14ymLdW4YA6h7zVfRVgK2nOiSHwAWsjCCsNKZIoxa7ItWuL
Q9Nx9/ELDmM/Fnf4a2zI5GvPdXwlL9LvSE9bSgXcL/GJJi3qBxtAC8OGcCBaXz4P
ByzCZNrEUcEqTl72VjREHzuFQAwNcSfEDMc1XnJM4xvvUfqschF3gHRDkWdQpgt9
QQF12yH0cI5GoSelG7x2wKFeOw6Fywb6lg65sjePW5YwOiqQJSUVE/wdtk9Q1pJ7
59h9Z0jPijx61z9Dp3Z9S+FxsWTqnVLvnmG/O8gGmM6A7fqL11ndoMr9cDOinlra
Dv38mkYyDDyjKebKpniPniqXg+u2+V97CswTYOXleOGGwvB5JFMnWNJ6KnXk040Z
tz4OX+7Btg2rEazgW0Y1RxruPZdzX9CMyPm66SzaovLOu3rvxM7tUMmT6RZru/b/
Ng4qcckn6cEU/5MPeAZ3o4q9drBEDnR+KIPOH/dSynrG1AQ41wHkzyoLq4UwU1aR
6k7Sf5l7ec4YbKhPJXg3xSMv/k6KdkATaW0gF08/j5hZ1gsLU6cGmM6zoVQNrZDx
QScTomZhu98qGQGcj1UHEaXzeoc7R2PHePcx0YVy9XoQ7ekPq56GlOn6Ka2YM+DI
iZhPnCPq0o1feygKo7zsQLPSH1oCKaDA/JFUNUOGD34fsUt19adI3b1JTo45hWRA
fMplWSi6byDmNUWDF/b2Vh6gdVW7vn2iw9Vu0EE6I0fkx42szvCXd6EIK2Avnq21
/DI2dL3X0nG9XCX7yPgqXKUvf6c30hlUFy4bpAL9Ax1fG/VwzKY54Zf/QmHBaHEJ
FV9ML2UEcsggA5GnXPP5UCyKJOaqYwd9FzRuO537C2dScIxEvBbrlEHbzbkcT3+B
p0/2Tx8NoLJ++evSpkEdhcUi8/R1xoL26I0fv/UJejvA4qvng/iCbLGZJTh2hL9Y
1oNaZCWVOwDIMeOtOB28WEtgTxKKdq1Xazl2rkLc45jmQghnQYoBjMlZ3Wo9YZ72
Hj3cOx1/t5EGEe5+yJaeBwM5v/aG/+v4rQ3QYTK92JjFH4IAu1+/cnctPEXXB9I7
V3GVys+Cj92rfxryPjI3sWLAl4IWu1ZBiwnC4TLd6G+jQoZmQ0QSvHpKWqIL84Zi
OfSMcsBNkVJPFNORliNJVdoXdZfRMV6Ft9ndlBzOEWqvdy6DQRriqtU2XXfzc9Te
UbCDBWm+kxO6ArNXJBftLkyszuhTGPAwjLnanrPzBtJL+svnJZCpblT2VoULoVtm
EMqcpWhULoffPrR1QsZOL1M3fxqqVjWwMFNpzjgn/jn7rcn4H5fCLByXl0S41z9d
WVCgnBfL7Zt1aFZ1VOPQyX7MgJPynscp+0eZa9MHE0qHnTbGOdrv2AxuAaUX6FTn
J9vVc0CgleRBc0mVOEqfkfo2Fe0S7odTczB3yAehO/Zu14Rjpmafk8zGvNxguWVI
Ma1PZEYMRw0YWh0aCrPaskuKi9+UAm77wateirftqMeLh5/ZaXPknh3CNB9Z90tZ
gbO0mUVACPk3jnaWb2A5U/T35jz+pOqMJPlEuytTllOqJynATxut+UETknJm6SuU
xI7pJNVH1190Z3mTDXx4aDmQk/hwqbn1ZIDBn2G6IUjiicOhaViVI+wlIsxkiwgh
z9/DlhCSpcuXL0RIRNNmDWjjjDUBAli8egWipZcLHGrsB3pj/fuMFnVwpa2GZESa
z/5EA0w1W88lLhAZIsxl3CzA/tzJOPzhw8yIA/9bjH//LzIZhvAtnPzZJ/Ue0OVa
Q8csWjt5JfEarkc+LLT5FOtt10SIkwP0O4bMh2HGTp5N+i03WAn6sllZWiga3pVO
I+S76O9VHGZgakrUG1osR5nxmMNxUz5NDIFqMbNm0qwlfwCSsxktpza2WpZvokoU
xbi6c1b5XdM2fOZFNNUPHeYNmv2l2qgl3+THjITF6QtcKDNIGGK0uUC4gkCwD0HM
XR/7kNHT6gv7RkAOB2CqeRJh3/cZuS4w6GTK9ZJEYs0Mk3PYTpCGV+y2AQLRRxKQ
ihtuZA6syLEjdOqSS9kVfyK3VMHqvhxqE3lJJ+IohWtbD4tVWbv9N60tZMgiM0pG
AYTQMGAAe7omRL6NsTu4TthSP0afYPiFpBinuHOHewC5Z+qyg3yL5QtdQh8Jjvs1
0wgoaTojaX1X0fM8uVhstl5C87EJe1Nm3xyzQ8XqlTQ/5rLxGG16KQS1MdgjolU1
Hw93ZK9ipP+E/ExKWrG+Adsqg4ACA5145RGvJjanhfC6hrD1Rznh27r9MqaxbUnN
Y590u88YsFmYj+We7W0ekJj69oy1Byqmjxw44GgyTq0rW5uye7+9H6/nPAD09mDe
QpBCe0TPD/M5P7WCQMFDohlJcEJEwOC2PEEJxdNmW//+FqywtWkG8xLLwxeZzXr0
mur3F7ROrjWJZx3LbOArPnQsZFQtAGaHhKA4ARdutpaFJbk7xn7vAOhCFvgdPeDZ
KiHPu3TOCSeuffT7Bsq6MW9HAS0qcZWTGUYJfYMsV73z3vQZNYYSbsz6CpPIKMrQ
cuDnl/EfI1i/sM6k34ign0bj94BfxvfrS1TgOS3mIsVX2HS/BFpa5CtgTHycR/iB
7cywd287FvAShREKwQJMLAKhFz9aZZcpNtd3DvavW10vWv3B2V2UczOUQa7gsa14
u+9FFzXrj3dQPps0+gBqYIhNf4aiMzO/Wll2ygon6lM8bgj+n3LR4t7q8K8+kUv7
mT/QUdAwPvUDLf8lplev8Up1NMxW5lMfgdC/Klo8loHi0/oTXIKkEMc6CqGwhhbi
L8raGrPjZuDi+PcA/SMKQeUS5EGBIn7Nq8lJhTDWdVQU/HMzK4b3EaTWCwXW+O8e
MWEXimhdOrif5iyI2qwOVwBcu5+4gwDQveW+/ZUvBDL8YneJVatOu31nVZHm8vC6
NUkvyHy2fY3yJoshNcyL3uquz+p6nSjhXBPaVDRUJeW+zg/I7KBsPIi41R0O8nQn
4hbCLJ5JAoXlQBd6rf0hLqNXPLbkl/J8zVbV7aYDIjlvF5Y38q7wAFNCzd/NB2ir
JQ1KIDhYebAGBJO8ms1eMzGvG0dyNWMcxxmlZ9YWKUEUizZV/p+rHrRFRgG3iGFm
tt1nck4vz0ntlogf6Ng5C/Bi+3u8/0Ffo+TNC5S1rgJlbw5XXsku/q0/GX+DXebx
2lfRNl9QWsKIUXtumtSzEM8pPGUBzbfsRnRVi6tIMV9J3tnrA6Ze0rDzuCVcXFz0
PyeGwqgzm0IRdMK6X1n0fzSFmzT3kchM1bZuuhAPZyPkTTD8JvWvCMECpPmpcFx6
FUay+gkro9RHllMrr04G/nOOSzIqQMpTL/Iwt3vtzq4ty93Mz89Vug/AFfxLfJv/
sHMJxACp3584mIsQUKzNJEhn00qWb88tv1hBxFs9G6P6NvbJKtsIo9S2RxVefLqp
bh4xXyRJm4Bwr4ZGKGkWxbfGXkLssWsq3CKrSpMR5UhupzplLq/75nLLrC+W0aNM
bx34fCLw50S0ZrLEH5E/BFwYRmmWhk3fisyX65Nq1aFc9KPyqpD0GpLZc4pyQM+3
Im1QTuvhar/RK3PYNJllCgFV5mwLNKuWdzV6gBjHECXYC+DluDFKz8/n1+UsOrCl
9Vp4xx44YqKRyvhIUe1cvOkTYilr54VHKGk/PKJfmSDnnLvHjFyj8t3IJXKBnCwx
9JFQj1qKpKWjYYuD6AwmQu92JROX7mAvzZrZtMspI9mU/rBpA552BnABY5JpPECB
J+f+rRLS4OdWejl6VdUnRav1wEs8BlUsP99F66VDP4MtAGLqFJ5yjE1eYmL+l6cL
JZkjd7Etn8+y1AfDyqK5KP8toO/XyFRcFOPdsztfCb0o5+BiTzp0/xz+z8w26v3s
Ml5pkb5YgmBbt2wx8zyImHibpRX4IFMVEA6UHR2Q3V6RZwROp99vwVesToVWTQC2
b4uqwR15xN9UeZPQZWGVpTAnMxj/GFoxHrpEJsg1QgAVJcIeGDQnVCSl1BFq2abM
2ld/GUSobQu3oqSdA0AvS6fKrrP8aD94tDzyDgYzP6fbMmTzvl5G7LHtOXyNsBsF
M86zsFgF2UQocd7Hhdqm+JVQXWoyV1l2mH+8HIS2sFD3Ytrqm8tu//M73kfHz6Fz
MgcSGF5ixMJjwXIjhzbxX4EmISJNZc46NPMnMtJw+5ZkQoCfIXPT6LA0ZZLSikVM
axMC6MD9hznoWT57x1iPSYojC30vcw/DXfoS8I2jVw+dwPhgEU7D3h2kMeJvlZam
D4uF2xkVYzc+GA695O6XGaUKel1zl9arJ3qh4GwJlcX9SI/eNXKhmMaAQU9+ZzPt
YRBRU4E9TEQNLX1cIQ5ZXtbyViucQtocissB77gF9hrlxHs5eKPFShRNXH0IqmLM
Q38Qxs5sMpsr0BqHqR99OKfiyHokjusDk5KW2mVPVvVVqBWBJtux8oqtW7qETpuW
mfjt2X/pxJl4+T+yG4vtbJtYvVMqo00+P3dQUK4y8lTLHLJsNP9nVoTQ7CjVaH7e
gbmhEYmbM0RsKxBRScD8VLm0lOf0FNOLF2+MhktPmxVDuxOC35Ct0PSHbXLSukQu
TbbLUxVNcG/W8HYclZCzaN30k2hJWX/xWq3KUje4TE8RK/ve+lGw78V91RUyZQkU
99VRKnWdbPLFt0ROgwYH8nsC473XBSE2oir08elMFwz58s8DzqkNEs3qHWOpOJ9B
aWcMk5zpWIBWtHGyaBkwpDOHOqQ9xOYKNNwxrI6b87YJ6XI+Ao6rTUc2ZGZKIsZO
5uL9JxM0UDgthITHQcwTr5YU14soMf86JvgVr/n8uJ0QhlXv9iUMNLmgNSrZiRmO
eZlo6Y72d2IdLhQJ7YyDhI37WPLLqlhD9sW278T2oX+9nt29r1laNXPMdhFEDBso
ErkTT/jE8b+JBEOvgjg3UB3LkokJFitsuRcPsl06CRrEBob3qCEgyVW5PYljUBON
66QZIumMXcDGt6eP+VHeQAaJ2G4HymDtfiHWeEQp1ftijozOBb9Mgajh9bg936Yz
rkrcMF11pLM7+HjJka6NwoN7oeyndY+rpo8KFgTB8507+/xALfC2j2IIhF9UX610
0pIe6gvpReA7g7ao2Xn16SGhxWu3h0z+sWNMASILiKbFVb1+FI3zn+KRzsOTz36d
5zn/6WJk+83t3ZCFoAEApQe2/w31d/rURiyV799dLpyqBgWylsChrPv8ZP0AhZhI
ejtCqgfmgJ4INwj+LSoGnP6hQWV36EH3BoS9KQBMurwfc7a09/wRkv+iDv/HLDvQ
MtSVvE0mrwVsDZWRopXVRi3q1Ix7vPtsh9+Lp0GQOXiWlsbFUWmKeMG5v5Gyt4Xn
3wPrCmByhFcPc+8pNd/+VE8612FmZLK3kNYHrv94sq2M3AZuk3QoAAe7gEXybL+j
4GHdlxPtVhy9FE9W9cJIL+ur7Hi1yGA+qjwAM5jBwY3Z2WfcVSEO4dZqDcqoO3Gb
KX8H+wLORG4CBqYEUIl8p3w5F1VO1ogr5bk1SgxlhVAOEz3FUMwbft73iqI0NMMt
MaJA+7mHKIC1pouctxRcuaNWSwIfYTlSUmNNFxq3iK6kj73V+XA9wsmM4GQOeeeX
aw1mqeESem1ABgwkHhVAAN7WgiL3OgSNlW4NND4DqvpPB+jkG29g18VXUkSdRVoZ
NLEHy62Kp7zDquIdIJlNDnFANbCmpun9etyMfAC5EHuYmGrlPA5GuZrVK7ws03U+
UrGaHFBENzDlPdO5rjfRlkCjJhZUFyjQsfzOEEKjdtsegOr1ykfjN679+CUOvc7q
iXdj6+X9BHA0IvwVbZ+Dj7hJPpwY/EIipU5rcXHKO6VReH9538MH/17PvobD1gzf
9WaQ2jJG+fMSESv/TGiLuRWNNlPk6nhODMPqCLj+G2oSTyD+NnE5IWHoECcLbZp9
HZdbEKr4/pb6N23We/T94lFIV/dj1HoeiavxQSrooytiCNdKjcw9aI9vC2NsfVr8
ZSvmIotwQYantQqtU2q8XW1xQyna7rddGf+CbcocN9gOUCcb2L+RvCw5jBAjC0nl
R5xgfbE/jMo7aySvYZQVlutmHYylVn8RWX6QBNq6K2vnYP5eKPf2xsEu44Cd0V01
UX9sn9zyBVam/Md/rfZzFywCRBGhX2AKx8MIE11J8ejZtXyB+Ae882K76PWekVkb
nNHwsnddfrfs8vlVzyqSb+0VC4n1L4jP5g4tGxzYu3Tr4WDG++KYe6OewoL0Pbgt
PnZRzeen+CRCF4UQwPGToBTqBsoxXIrU9tAs/Wx5oK7aymekS/5CbYacNWWePuwu
DXX67ERflPArfx46m9CdFvcBtOmvPrS/aUIf6wbn6LlKUAQvdYiod0kaNgRqWkGR
GocQyha9W9f4N+XjObnmQ3UKxPu6RXtdxryi2s2xqqBXNUAIjgEcwywIrwviSsI8
tkU9dhln6w/Dh6Zg3OTlPCINd+zNeAur8ItqZmtwgilcFvuc7oSsO9S0vlpcN6FR
nNVzNRKLWSj+KMdUVPny6jMcnnbDfoEBPkvH1B/fICluoxxhEhcd+btIVaK6BSKV
6W0qjhXwUtPhxWUqZmMWS3fxVKDvNGzVA+Aam17V5XWXQp4a3Oh4GGVYFPKGBx3n
XCi0L/qzcUcn6EKV37CKpBYI9WKZseMSic1LFS2PaomgmhbzQlihw+EW2pj//foW
+dE1tz0cH5Atvf2tzvezUXIWbj9aLsX5/1wtR+J2G6m6QHIQTTToM7N0VWbfmLS5
ktgVD8IBPH75urQAMH5z1JtFvyR/rK97tpgf4kmn8pYDSNRDcqXYJEWf4HJfkwNk
gL45DYQpiwMnWMSSb0ooxycnHZ2v36mAF8dlDX2ZUrpt9sExwphJSCE+18gJ7uNC
csDyt8h5NMQVduOMEgihnv/42HTZDgzkOQdQhrEFUc1qAb8jdjSMqDT3kShhsBKM
7j04V035BAsPS0w8nHVJ7l9ooYqw18WxTI8qi7ffByP6BH88YxefBwk2rq0l8XsM
D53vTigwVgA6hJm9WU6SP9OVgAhjsE1QutDcThM6C3xgR15EHKnpbphm97Oab7yZ
38SlqTeF5vJjKZsT7NzaVqHvoOEwdiuW36tY71BPCW8VIC9wqNkul5kRtTtMGh+E
3/BfRgLvgTG1EjsZJaSPW3LwZRviDn0fYIPoIUxvr8id1blPHebNkncZkbccJX1R
gVRycc1BeQ8INqyLKeX3XT2H9W9Iam+UZCzzU29j4zaazMxTm5yAPQiWLKZxDI1N
q9nMW+030PdiEqw1uL5+qXW2vNpRJGOlZR2v4trg17GiOU3oC4NtqRLBvazCzqnN
qeiYASQJIbDPWglPxZvNi2LtBWX+tL6cxr3FwSKxlg1teYQoA6NCCTt1D4gk8F3O
+IDs3xI/PQsrf/DdBXNhjLWN0jBdLbPf2drocO9t+aShOLMeI8D4Ich3ODFHGgvv
Mauh2nO/FVpeEiASdu5qS6m4JKcjPaNmCfZ8PlqADfiyGquxg4aMEQ0uUVd86Fha
b2sBPtjGpLwHgR8sTVfwzMT1ZrC/Tn5C8ZHkqC6iTNHEIhSfyqGG0TTu/ipK+6vQ
G10yGGtEy/Hc4lhyrN+n6jIuR6oAYmoadp4lsohjfwPdN6lvRWcIAjclC5HOoxEg
XgXGekqjFsKsuQCzsb/lCzzHMNf96Nm2dqGWnKbJtaqNtmdpbmO38I5MMO1nuZQd
dGDu/p6TL3rWgDmP1EBHeLpZ2QPq0u/3yOpUal+x7L8Gf/tcS3siJJ0Cf1x9kwlJ
wZjBO8MfzuEFqh+NCWjropvJ1Hs6g9yMFwVxzDxfudFu7gX59mqmC/wyW22xzZ8C
m9YRWyATFJYNuwddBa0h3ExgmAhuvc0QbP17VNgXVJu3oi973eJxoBp78i/k77SG
ST9tkhOcSm6/cBIcn2LPhrJr3R8ouQvW/i3tNItO22owcP6Mu4mcvIaDeIcquFqq
+9J22RrlldXDEBcLACiO5/4d0YdOIRinp3HL9d6j/5oKf/mR5wkO0C8FawhkwSBe
MsdZ51pgDbzp/LFd0qoUP1bZ/5eiTX4cihNiw3woK899SGJZe5HH6C+fh0VuJ4sG
rKq6L5Y/zDCx7omvOOwGKFzrJZ9xUuHhFsfspX3o0iCMzRtUeMl3vFWLku7IpDPF
91z7szsChyEVgxqYwcjXNqXRY2k41vnWuVTTz58xIcYrauN9ybmCTM1ssm7bMZgP
Qm/zBwKMaWT4Su2ZfSIxpaZNfanN+bx/TxYsuoDgnh7/kts+LfoeJaBRlYnwFpsI
DsngwWH4oZIo1d/R35R/tba86iVQ+lWJVOu5yD1tHXpA0KRXGOB2aqkT2Fu1hCa9
UQg/a5SZGV0boPov0tnhU4ZaaYEo61HqfxULwlodUwRg0U/QAe2qyVvBUuubjmo+
FobfhMFwpW/CBSd3zLIUSiKCkebue7H2Dx1ourUx9f5dcj1Y8m31QNh/0iz1fA4R
ejotuo8m4dhL/T5ct3JYum329fsfKgV07pzXMyXVSau0+JFFwxsaEyQ/0XccHAYM
plGnixQiGHqqn2C4a++yjAfNDviwhR64OiwOHMn8ZxbxbeykG2cxuEmFatA8ZUi6
RmMiuwSHAeZzeH5l4Qhaz+uxEUsDYsfk5H6lMEkcaIqGP/bq2jlvoflYvpgSNwEa
6OIHbcHiviYUW+ufFmNOYn4GJ2eS7aQnw11kY9a45vctguaTJ8eyGIoz0VYDuxFN
EKZLbjqy/kWBlmELdCVZk83UrdQ4amDv5w3CBc3KgV0vJI5cXdCAdpTRKQbDrYDO
3AnP7eHcb1Q5uDvicweL4YnwEyv7QqUeeaQz2nhIcPfOyo/VGjOjh2TcubO5iiy1
QNpVWZGEFVm+schGmjFHyO4c76B76bReVuDEU96qwG6Ufl0wVV6n1iVjDhrG/WSx
AbKTmjPJ5N/qZ/U5V7ursLVG2gDaCtjTzEtiWKRKkdknD+kFrmLVfct3+ROsyyti
J8bZTGPqZBEwC1AMUwTgiMDl+ZDHDq6lkNPkS+FfyqaK2ho4oU/lBq0sEUH6DA8r
cxmAWQ3mN2Cr6enyLnGyAwcBa771MyvYN34IHyHtKhtS6zTuV4sbNtg8Q1oM1W5c
FxO3Z1FxXX6etkZvLolgh/a2ZTIu1Tl/PA6Rp0uD6+QoiEP+MvfHevr5SsjAhhPu
vgj7eRETr3UfHVkqLFTQV1HeNYpvo5SzX2yz9jIcK0D6edjFih3WFRZwAiJr/xTx
XZmh+O3Gkk4Vgf/WinNRSbohlbFK2B7abCfpBkHw5zJsNePiVwZEoVfBjdBmN8S1
nsKmHeSoxo9xC0KeKe8GWsr568mv+HTZVLiCS2qUbP5EqzvDhbRCShD4QAkAJfPm
TaQ/B0N4oYQz3MLiWCih7PnsGYdKMlDz9wCR9ZRNrnC5DZEaYlQKWlxvOCMCRquX
gPtJvwwsiJCL+QFmCaPV4UAHSawQ645t9H6EZc7mt6GypetmF8///gqozD2hQGNs
QZncynQirRaqKmQ9vSxUoiVfoykDyta1N7v6GQwD4YB8n/Zl+UXJavV4VS2OzlWU
U+jDpkS31YTFPq7BAj4x24Dml6mT1E6SI0AT1Z4hxcQpV86snKUpmSY9PBWiKzDJ
UrTfuTRnVEkfJoE+t0z/trl4LamAP7aVsMo2UD5ztx+byQ57xO1/oh5FRKQoZ6n4
31f9Hfyd/Dgh36CPPGABTTEOpqTHLjN5Cm+di9DD3uVeg4cgrCNAx4Cpn8d/scQk
zbXsKsYseOqIVKy2QLfbWVHRhgPt11hyCF7j4Zyu15AneXNkNwRbNSjB1n3gHbPa
BiH7Xk4EAvwJX8dOtFXlYoFWfJZ2c0zC6dyzfmQ8ULhQFRli5Vfa9HWdxxPHJdmf
S+gfE/ZseWmUV9UeALd+8VsMN9be9bK6o/l2cT94Wfd0HRKg26SkHHgC8vW/lvn0
ufUuF8havT89BV/HzQ3nnG3rUexsw/BO3CV4hciqblJyD71Ql1K/6xBbKb5ljfR1
XD2HBkA+92ro0cfTZjemPygGXsKkByEr8IA1fI3rd6kanEMCVpG9ptU5Y75gFe9p
8IwjwZZ3lHmAdGIV3+MQMcQe4C6nBO6LNBDiWURdGj9ldNgD5t0N6ncz7oLov8Yz
A1JqKtobgQXHPif3vuaBzWRfXz4KEQpem8qz3oBcVDd3LuAdzqD5/CfjTJQlpxZ0
UkoCRDO/ho3oEAkJvTE9qFFkCwjWw0HJ9vHPLCJYM9S66u6lhG7ZMAHgaPb5cPTm
s61AIw8nF85t/tdX+3DuWD/eHucmKEgQubq15XGcBEhQ0Q1Nn2dh8GcovfPZAwIJ
HojY0Ixg4W9GJZ6v9FdjPWQH6eRxfriLfyP3J2UkdwVjmLCFtYasfG8p7TGYy4aD
7DzDOSr+lfoOWzZ/rRV7+q5DOz5Sogrd/YZpUDkQ+W5S5/Za4sIWtAHRm/BBeICc
L/URA3jKPPjTdEybj35Yu2fUT6eai6DflZ4kzIeAZ3o1vZEcrnTRPnUpr1Y648eH
5tViD+/eEKcIhsKcEctkulbBbBSJHzuDqJhXRxMomz0Q5xgnGmarf92aLj7WxNXs
K2bVaCZGrclnZezlpuTLh1waRTRBaMj/1tOKYjphwTdTpnZm6Mn2GWAIycykSces
zrdgyyrSspzrnJrNFD2NnAQtTWEk/loSw4+j6jwodxRnpuuhRl/IBd6Fm5jQ09Sy
Mb5J1arA7UW5DX5ic8bah2SY6uOXjKhuM/zibDySBxJQ/fCfEeNBuVBDWFr2lBjO
DWLSuO22IHShIS+vdB2m790iM1iNsoPszYjq+a+t78r0XsDlqCfSRcVuJSguexaP
nmJU4i9D7UeDp4XJPSRcrXjRZXad0lVJddx/fOtvaIG246u3frb7gBf22qSDf1bo
XwXq+axg2jnt74KpenOMzgbNH+WdGsG+vECyeJ19JwbQhl8+U8nSdK1yiDX08c6r
rmJ6DV6eQCdJKl3p3oA5PaLrXL7UNAC3rwwxcranViLToFwUizX+ReXRREB83r4X
wtdXfflEl/vgUBVJ/8f+9O/wz7RJEyhD4TW0e2XX7y+Ac8Qc7vQi0X4Jh6luUtJ9
7mcey48ACWeYvS42j8Yh9k5TlzAep8BD9rj0E9aYR/ybU6olla2dLHFYBZLj7Wzj
Uwh9LiAI1FFs30rJKLyIPejYP9Vtt67CwaK6kNAaH6ipVGrSird1h/QwURmK/9vr
sIUxWA5zepO4XBkq4mM097e9pb1edk2/Kuy83kcCg7DjVKSjkuvMu0DHkQVZZsVB
AHA1MrLz2lc/JlruMtZlRlKZ9+9x8qI28Zd4vP9eA1VF/m/tIxqcPJOppUImtN57
V8dz2MWXyABXwSsmItVBq8zsO2vvs75OGsH3AzFtzGqBBxkcm2K4OpEVL5fWaNzY
G08dc54p8LO5ikNfqyDawSXRGBYvNnA6uCa65A3djMlMWZMfsad28Rq3mX7v0J64
l+XJq1XcWvQlEKfrYeLCs3q9kywC3LBBBYrl0zeDqG7TUsHNFtVq/fQ7nMFyqJUi
ptUsS0HeXR3L8rc0iQcqlR/wCOBxQligMRW84YVAw1RVsjMGr8xwg7N0zwhRsG1S
4vluJqb3SQpkZSMpa1NuL42Sep7a/p1rH7mKZp1rYmc0h+G8wtSQfw6t5GM3oV1O
z+wBNBKsYe3kkx9wVRKRYMj62SGW3MyKbKv2Pbd7E0xZKLcgpig4p88whirRkjvc
CdGPfKYcO5VpES0XDmykvcJYNPQQe9RU3mAzcx2h96LruJUFjvZqZAG/tVFCdxKg
HeJmGdNx7BPujodj0QFyAS1xM0EOjuUHN31ixw5U9zjmxdkcEDNAPvrC/2y42+lK
M5fOgc4c40BpkicMda8KzjG9tDEoGQyJG7CABIkav/+8zodZkjKzOyCIPphkdMUD
wrjOXTVHVkb8gqdboJ7SrIvg4kK/FlTZDw2sVe8n5nf+msOGLLdQ7j2QzhIm0+Xj
pmgp4oQH/dS7PQFW6mlxiIdU3PTu4Gl0p7D6qY0qeY/zk9E3wgp8nYBLX/mZrbYZ
fK0qxg7SA5QcgZ95Ibw62LKwyHBSfnrKNyV5slApE5x8zJnsWBO8I27hHoolAgYN
LvIcVms8gDpUaJqoTF/Aucvc53KHDNgFpYsx9JqMhNPYWa+S/awHL73q7xPnoSW5
ffjelNo4vo7Xmf3kBvfBQEQqqStFj8YKVsDD88oiLwDbYaI0yPHGv4yIZC5ZlOus
P8sL8MRuqOBtS/D74UmMUwt5fXtRGVzohTA3fdztrXh3Kax4m7g7vezacN9I09Ct
EzCqGH1YqYh2LrNr6OPv1rgr18GsWAYo+CAQ5/kn1rzW9qEIeSq31VepBvE6X3/x
8wMv39MHbjZOUawQfSpQIEOWC8HGVB5j+YGRdwWQXyyYlQJ73wC29Hi7nrpIo3k7
ScqxkfZNJeXTzB1xLbk9Rt7iqwS5kOJMp8aUWdb8yOuWWkjpg3GpjhNPT9dJuO1W
O+Mjj1eiQWXhYSt6NmkrmEoT8u5miSg1P3ie9nl2MnkQV/ueR5iIuCsrziWipdBQ
FKKFOHP0m1toMtLug5i/6GfxPVhR2S1cUNN9Hz3DjS9QQEGED4FLkNSVQ+tExLMU
59ieoSC4KH+tVEl6eWc1Cng5fJtc3WmZalt5bv6sAvxYYtcwBuvO/PLF9dt0Z2jq
OIrAco4lsUApL8aKK00ih4Sh3B+BHPfAimHkYapcetaGvEJ03o6pQs+ID65SUHjz
eNRNk7WchoQyx76KLqRfpxhsiY2SqFwaLcWTgANdy4OpRqkVWsCXqTxThuTFiteg
LQcff3kWySCXUeTle9ruM2Y/T/chycVShsAm1kRdN9CCAKrZsPkZ3+iiyQSS4hl5
Y8wr6ZR2bv3r1NaYpiua6nw/R+KTIhQhENw5hCfTCG0cKL6TXc3pUOhjvu/6yILi
i4nETviy62dvKSxi3k6oBPxUZ/K1mCdAe9+VAf+L3kfdI+digdpvcQo5tfloUl7m
isQzE3jGgJfbL9BjDGjX+xchHmfz3qTThwBomTvJifdzdfweTn+MgIPk/NR0kEd6
Y6M56F9JoDQySL4CDjeZcdPtKMze5MkNnZ9GVRLADJFU3WPbrNpn5oWv/eYo/lsK
dAgpbjroHAHfs7F5nuWz3Be/ovzcHhBm79t47cCAND6rS77qt0EztZsof011U7Pj
3SpQBPpqQBTwLOmIY1LxGqsoLqUL2+kLAmxxyMyJvcS+/7P21ltnZXx/KaX21qx2
Iizq2EHVJXp8TtF9XDlribbWkiuil9JzkDnaxi7PL6MQClqImPLyvN4s80Q4ulqK
P26effSfxOrd2TtHiU9QocnHpBkta7xrVvlASNyY/7ncuXL940bUz8yVFeEljgHf
qesUTeIVga42Ke1Z1ccetISQVHv7HKf6oP3Pk42osBHQpxTBVT7llVUIf/8YHfEZ
EL9edy19T9ZR3IfBdX55fZctugZW5uFTgkGuakjkbX1tqAkyixSJ7Z5fy1ZpeBDi
fxCZ3kKaPd12vquQRMTLJTbkLdMMp06xRo82jKCvN6tGCt4XImhJf+wFZhlwKEln
cQlRUtZ/OWDmW44g7lfHIzewZi1FeaznShqTdA+K+8ktHmjn+LY6NAOd+uxujOWA
90HNDLVFGR7YUM0nui/lgZDbCd03X7aIiq3Q/ijwZPWxlTnwcdHyMqkU41xxp5CY
5ArST4Q4+BGT1xbXNz77srZHmL38m9TR1voJ6cG2RNtKOWhv3N0qJ1ihIAMR15p4
4cMYmQtSfOjuIv/P7QOWjacsbQIHIFyw0QFFXJHHMEmRaYmlxZnwAv9J2wnTXeJx
dQ5HcQ2sowKhpWknSqCc7GuDo/7ob+P91wtbSRfPWdySOGfimc89LGTnFlv1mKyp
K2bQVhDhdaiBmwDw242wEITxylbjPov6e5moUkAhbw+CNBAwRkGm9yPp463hpuYG
apqtTqbO5In0UCwlAQM9Ua458PWaaqVtU3NiUbYuBuEZoFgPP0hyticixMh33CCy
WWHZ3/WuKOCFb/Zs+zvVWAsruW5T50QoMF/uKQ5Iw4b4cyWhZNXlij7vZbKk86Kz
17av0+Ie93xGW+7XJqGGKkOdef+eMEux2a7YJzzsvzCzPD7H64PSicX5GS5XVt4i
W9QnhIJYxySutaCiFhdTiHM8Y+9uFO4aTBvi87PKgVOwrPK8XFyWZSHcWXh93z4B
bAPMgGC5JvZ6P8n3DoGCRSwwmMeIObBnp0DeitO+XoVzhX/te3mntNAexkvNfBEP
4AI5jdXaaxdS8IPBHPz+oZHi2AToL/qCKh4jjyucRdSmGuglfedPlThS7oDgPnRh
xpqZbuIWFI0kDZoawZjAxCjbq4zMZ1QcV3oi/wcYfBKzkwkHmpfE0SrMU01QWuFX
dp0HkwZZp9obO2yK9WUunmoOz4U9dDCp0UMcpdcVRNUqsHtkvsLaj+e54qx7Bow3
EUCDfLMvWIUBAeO0CymQEgHzA8rdjL0eXU0Gz1hKlW7m5L1+Qjm8hsgb7ZjpLqHA
8mPUAdfaZim09n1IZlHXNMPsvIcG2FXJmmaxdJRsSXDocynBMEWhXD1fyJ6LMrYz
SS2lTGhNOAUUD2C+EMgQNpPc2OdhpKbePZlDVlfss5YWuaaclGGs3ByjsL14lyCH
Y/7t8+/sAKxSit2IyB8ggqrirUhm9FrLj9MfE1ffAATKnzJZzkWGNRbYo+2RvIvF
HjlZCXZyvxG5SsB+wH0Y1Gb5WdEU7XRq4/nozzGHdQZInzNOqnWmrTlfNnWeetY0
bhssr0jKteVlmNdsgnSHdWuHzu5bm6sdPna0uc69nFqIKkab4Mu04GocjmDG6XFx
KoA8teUDoWNn/QEMUUDiWh28S7L58kmimWAuLOTQ5sd7lA+uCn1t/eB3aHGd0Qur
PmOBk+vmKKDhqt2jf9KR7GpBKs1BTM9yn4jbE0WSQjVmvGRGauT1wlUFGLdoR0mA
0fqQyrZfI4u29A0otlxiXblWq/mKo29c66+1zFFqwHqbxkHisS0NGdbsqDwYyFdm
pYTvwT1xdiZWANxcaRyZwDDRdI29+PJD2TSb9wFoUD/kQunbFM4ph1bg27vH4FG0
gHOe6GFVSFqysOkoIlqVymVwaxhujnGST3SHHjsajKBDaq1d8nYNEew6wPX0iH8P
UUSUg2kJ7mYsJs93+akxgXz++9U6lMsxBRAvK/NipHJbQGRmrnl5Q56aAnuynR9f
Tm4INiRy538+MnILRvH1e7ern/Fx++SOy2ej+9C+tb8MAHzLqVdpNn4sBGk2ID0O
HYRizIxQkw8OWVYXY5SKj8QHyYvNniVJhw7f8JPPbzVeHA6tFlGuZT66ydzq0AW3
Tf3U1G69Yi6YSeHHi8dskTe6xXWTGRDlxfp2RRdJijoclbpcFS6HlA1SgbIkV+Gs
aLisoxXpiH5Gy5nFpX0plzsEKpPYiB6Q6EK6Kq73Nu6RCqLRjawu6K/Oiap+oPiW
vcRwRNdNk0n0ZgifNVvngPdKmfci8jdMvVq8JkT/tuwaeYkjV3yel/vbfY3CslPd
vBHfmgRa9OomeK+ptYSjztXhEFK0QCratCZkJAD/ej1mIVFca0tR08hsrAJ3VTDj
INvCpyXRk5qBcGDw+i2sCf3UpulklYf/11pYzk0w4SF2nEXs9FxOcFTwb1qRXwDy
UiGZMeCxdu/QhPapZfPYIBFPiydUjlOydCkdLH79sYMezJsEWkcWQdSfKYQPHQy2
oe8/nd914xcrbNy9bt7wyHJr4HcEuw5U1nExH8BUV1vbgtGsgwZxzkPYaUylTsA0
Cp9qtMZ7+0G4XSvjyB6Ofj6DUxjA6PA1UzeFXC4bKdjsVXUPcW0wx6oS8aokjI9c
xLH1Ww/hZmMqSmgFycG3RdFgAoVzFq5Kv02Gaus0OTwkCVD2GTX32dNUCDimcQ3k
j3HlB8c3GJzUBie4VoiDWznNuXgQS0OE0LT85fc9DR+vFea9gucV0hFbBlb6c0Fw
LPmQOwT6VUbrKhUF27vpAwr67jGQxt/Xz8y0IHjwz1Pq/Dgsl2ULAsGISWPiWzyD
Iji3QmkE20TMdSFyZcHkPLulG8tcBpssJG7i4eF7vfCZusMKWQLpmsq+GCGz/5b4
/EcnMyD62z/kz78eFNicChyrQ8WHCORX+oAyfjhYJiTx1jZ6qa0bSNf6JKFbIX2i
YpzLhgsOMzaW0/H3lB/APPTpbDPBCHfTZlYmEv3J1VuDxZmFEuK1HMn4JFrW8OHc
HPcmTplrx/RZfo3/Q0MkrN5Wxz0trYumEclIVxK1hWGrjiql24He/jiAEJzycctl
zKcCMlzp8d0UEMhbi+Wt4sicj/BPTtVfBrC7E+up8zMIl8Nz9BPe9mzbXD1B9crX
1ZzJxeRwt8juovVATLvXXULlXnNNaB/5N34vqI1TWc61gnUkJnW17hcjePjZSgJF
C1kjEwLdQiD//KXb1uOynCCbcsb35nPXDl+o62BM16YKZbPmJhS83ybJLdMpmsDP
F5Jo/4lBtrtfspEk4IUMzGcX8X0jXk9MLWHwrDw7XDT3sZUkDB46PZwUxrekvABY
BCfUqdPlAvisj2ZZUUYREraRYTyLVGgF/NW4pJx3NYdqSqMUxPbG+KUNuQdR4UpR
0nK4k1+I0UnTEF6vuZ8m+PQItBx8NHN13nxnue50N3c7pcsa/qlFbY1YyxS5iJr7
n7ddAFWQHJSFCQw3tJjXgFtH1nOxHAb9Kyrm98lNs4vLQCdeAGNbTbIBXbnYp1Qf
6AuAJTYL7asyk2+5A6qhL6sEv1f9u+YRoYDwg44iz3j9Wq7KHMMRxyE2vHQ+7mDv
Cwu0bhdI/9ACAg82XI0xoSgKjIJmXV3FpcGPLtdsif+JOUtpl/RKDgJPkl4pvgnc
YLKDkZJsBLeCB8I7pQaZfSsLaK0PsrUMLTPbnLyOwWpy53EgZ1L4yzeUa/Y5orkf
wFnHxMyEOcVcbnaVEu1niN/jp5qF8jb2pydJi9ctLj+v0mElgmNAMz8m1f+eF3AD
2eAoWrdUnwl43/vmce7ghDBy4/Dcx7IQLLE3VarGxD028fXsZ1Or60lomH52aLc1
Jb8d05+TGZU2JdzeBjR2NGH+ugExUI734splykEyvjSyZfmHAXw1T7EJz/9sBy+Q
qSnsShKDi1nkAbsUVJvSFjoNEOkgOEm3550tgevMFYym88BYuK/BmOqU8yIPaDpR
BQ5MAgdjQEnQ4qMEBPa6YeEnmA/ruGs/hxU9V2sOEqt9ft8XbDf1hLaiwa85r3H6
C87J6dNMXla272PLIFjUGgNtCJiCILlwyz7IBT3sT4KCD/gMJeALSQdWWSP4d/S6
1EAhtRFvbwH1ZZogX0K5yJYdPIcPsLwtMzE/9QhP0hU0VEioD/6CppTMOd3T0gXA
/e5BKwd+VVv7QpZkFaH+T6350ErmKw50Sfw95Y4BcwCtCdpblVBRzjkVj7lnpli6
j7nPNop9hVb0GIejThEE3y8vhLBGeN/gx4elWxgurNTQO+DZauQQBcW5zmLDV7dN
lfyhpYBgFHeJgB7mdVU4rVlWfCGrUbeFC0RqpwwzgmzaSlb/90eM83PpiJvdiiHb
eyc1BnUZdb+WZIdfL1FX+TEhHVSjopzu/iqZOAf1O/QomA7oPbPdggIj+j2hLo32
bvtVd3JlRWt7NdtKuZF/t17rKiWmeOy5EhzliYpIWqgHhm5uZdfoM73cyHvforbK
lkit24WsDejnXgCL7N1vF3rBMiWSMOAsNKXTdBue+gbk94xpRABJrvH1oRykgyqO
6OyttnGTNavpZDRHUVBm+fMbBPnaJJQQpvMdBzG6/wDAM0eC436wJuh1ZHiSB6Jj
G9IOYgGPa3y0L2ilZ4f+wOGOdIp0KeBlSdp24p/5VLQUFTBGV1qkBq0+V7zh81Pt
44027AUFukw9b2R8aHz8rf1LsTL2WEqgn2+2rWYtgZQTl3g89/0l15/yKQYhNvtd
mOB6O+6bYGS+S6osoIzqopxGmM4JU/XYjrJqBa/RojzvBHWvrY9RohksCmriSdL9
7PptMAHdc8uSVd64XgFUD4aGQ0Yd4vnw6a8cyzTDvNTbfTG8WLijW+8utG+mbruf
aKkswD+nj2Wb+z2jb0ykxX0YEzJQ1Z8vqVkaa9phvnP6sh5dRJfo3n71jx951su6
LoIr/9q7YcgkQ+swk0RJPFZaggAVHlBJBiK04iuD4ajjY3p483fAGfZq9IFG5hFU
YGI+9PJvJ6C+wURI3eyJl3dg4zYTDusMJPgQDivMcs//yIA/fplYyCY82ZGdCCmI
NJKZgsz483MS7+2mo4XMU01523kh5JsfOo/vLiKqVNseuzsk0k2K0nHrwUkyRu8O
Tg2rKnWKTKRHI1CWqQLXgIzI/4wZolWd5QCPNUHjmCwIjyBGuhPp1qW1opCRaFRE
KnfHj45+7TB7ewPuLjFNGCcd4S0N8ChtRH2jemfjvFFn/pDVlOoza/qukw9BSOij
Xac9yEYvk348kktow9KI8bWc1gXNtHaMIlhjdP8NnIV/oesV8yBYNHV+obo7LVjY
wlnyRvPYa2s4H0wZmZyjutnBqy6TlqZSsmOjGRndbTm5F4UdJu6xu2b8YpiV4tF7
RHXef0zSB0P1G6EIFV3cwQAO6zuvmAuNblVsqB+5yDYC1Ho+f3/l3aTCG2+544z2
bRB3rbXO8jMY3ga3Xrii5+A2LTYk74zYFzvMr5r3BQQBBGVNqaXHvngQlLizoMMi
gOcwQYx4eNHcLjNJFcYUZoZyR0yNBsWWzYwE1SqdFbcx+rBrKhczWugyQGE1hFIv
bhAeWESqh/0/Ctq+htJOrLRcAC2cEoIh/KoJFy1WyCd4XAob9aXRxcy9WdPAYgUj
Hh12tpXQ/8q5hRUzzcKkuMIwfo5IE3EIVKYVKkxhddEP3KPXSWEl+mQzzOCF2Zkv
XvRoWd3drRbNXzbD3TwiSxLZdhq0D6beBRmOgMd+K+y9WRYE9zpc+pHIzXuEliYy
Voksbpt3ySnDNrf8qKKDVsW0gDK1FVGUs0876WVqbOSW8taaQyzgswoWHBz0IBqc
NHmhFTQCsUTUKVzveXQuiXH9fQYQdREtzDUGEsmv1CWvfxyqj4DVnyl2DBUJ4Mh5
rpB2iM8idGwTwxaWvZG6Pl3URKXx7s7ZP9MPCUaTPWyCGkPzHu/SvMBpfwaJiGYn
URS9ml8EZQ+ztXWLlFePZ7yr6S6/xuW2v4h1tK+2/euvntcK6BdssFuoSoqn/XkT
j+qefA0IMfBUU9xfTvD16j05rdvE1Fhr3Z7Xq5HN3lMBLod5FkRP2GHlNHE6ZRAa
NF6FbEEOKSaYrRDHxW491ccrsEhoim/gx691pDYWb994kiaQqmKYqIh+e0Zhox6N
k8C6eBnnhFcGEQdq/y5wFqu2uG1/ELIEhbpU2s0JPn4bDecaxbYeDhIbnaunsYG3
oQ42ZdsRIIO120Y4Ucltf3pgcSTEkqSnU+i4+iz7/3e8YGVBGJTefAprD/P0kJn3
TGvb3WSj/ATmI1++bOUhcQZG0cOATwz2VAY7Hi+XknfdSxx4mbJ6fMsV9LsgPrIi
97rNs2BSxkB9YzHC0gmn8NH1kMsU5ydsiS3gIs4n/ENrPzHPj5bH0iApgoINln0a
lpMn2njVARXg7Kk/5sx4LxCW98TUm3UbB6UFivHAbEncpnbK0TqBC4LCSxWqpDKP
l3u0BVg8rNRO6wKSL3rLUPimPleuAsC/9fPk8ovqwKlYiXhouWCZH7mKkpYBgl3i
icsKYlzy2c4/zJ5J1TLJBgcFonDZnphKh0VPLFcbaNl0lltnfdS1O28EyvIfse18
q9+smTf9bRW0ReZr4iueqd//nf3+BXLV/JT4YqyNgN226B+vomOoy7cVuBlQ0MdT
M0773HwdM6WcrhxWU/rlT03lWuOFpwGv6H1Y3a+o5LvxkKBW2E/j5mGyw/9zlSkk
zCbkKMwD/wI4yB5pF8i4wVF/Mv+lEMBTYPAlPIyLc9s/+MTUUjB/OyY04IL7P0+I
UMfY42ZHrhtbyGjyPMasiSjgqmYR1jH4/zXEUoNGc7RbfQcXAZfNUjfSw1rrGUSB
GCoDMku63fD2IZHL2jTePanriVAkkRU4q09xAfd7WjQFHgl3+90sWjkGUTtgHQND
iM4RIqdyKckuVCB5mJBjk5k+WP7e1FGKsi6WzihOqKbV0anc/gMSBynEW+FSQPZq
RcwyXfWcFL63JvK0UqlajQdtACMWpZ+yWv6N1KzbRzSkdwl0ybJgyNxberDflQsQ
3ew/ItlNEV3mBzAfnkZRaRJUbN8MjTCjgc6AHWZecqf4kAhXAs+cNz5uGRdt+yrW
PrGm/aaF+0eY7n5qG7cLBbUUU5Yj9fdxvCMjU0WFx5Wq6jmUJWg9DgEmZLdnUD/w
LPmqUyTKlrvC9wWrnxp1ygwrwdLQo/RXGoTORdAoJpCLX2g7B+eIJiXvT4qJkFxW
CewZ2/zDRgdy2LKTrxKIcDDeCxIcjMhk8WLtMtFlVOiuqT1KU3+eweeBwU+gxTs8
aCaZVrMDnE3DPoeQehQXN77zR9ZJtKg3fN61lvGC4q2LG+dxPmV/KI4Em1cSGnvn
KfvdldsUt3MMMT1quVRlFYc8DCb1RBGRKX+SsVqmGbuqmr0Wwm4waYASf/8O6OnK
4q+lfc2OI/uztJ0YUl4pOXVYZm/jGZzCoWzv5Z/HuZV2jA41OjC6sAVr6jsqewip
ARqN1llT5dHGGLJDYr3Rk605vhoWu1iyl/J9aWIlxtDVQIGgac0GpQ7ui5w0y8VK
fwzFwFkDVv/LQ4f9LItaG5SAkMgbGUcjLrlfmxXkjADDR/oTouL4U23JdvZr8LGu
u9dKuWdzJq97PAwGYPb7CMDz5wZIT6wZ+m/zbQMTnsT5gItpqF5tK5SbVEBi711q
Kh96pjFvbzSMaFfo9FMykld5R2QCDJmI5MQylVZsMTqv0V/Fk9Lm/4zr8FHN2pXW
cW3wLPqeGQvIBl8XByRyG59Z7h+j6maVVFiSZ6L2eyh492+TJhRnFlCYB+nXKzxi
6izQ3UIGwbKv8ddjdz28OL8NBK1b6hlh2Tt236S3JqedrfqWhf5sjiZOOBc12Sdx
1LRPU2e8dxKrgTRizSH/g35TaRH5i1LjbYnHI639zjUm1XZtNHZy+So4Nz5nj3We
hphB1S0ahdpStlGQsgS3N8tRMQmarPT5ho0gAM7nxXijeIB3wzASDat2gkPngVmT
0ceBAxoA5N5RK81AMwB2gmbW0K7qwph8LXUQ9XDtgMI9vSlL5dtifEOXl4Qg1PMN
0s/wa9NuwCmGMjwRv6LzyYhBEzj6oyMjjEH4zGj78bkOnhqX5pMsKLT9PCrEiZLQ
ZmcTnBRGf/8tWPCxhmARS2LhP1yCtiRqiKvTYyPc6VP1Girs8Akk3J0byGsl4EQk
Xp/Rga0sQbYl1fSpnBZ4Kt5B8lRj6izABY1h2hhes/lsabbvsyZE+dxCPrIzUlET
On3Uikh5n03rs4J+LH7pwiUnA3XZP+DC3cDzwcR6TJicc6J4aAEpMbm8pxBjI61x
Tm2jPtR3e09CS9WMyI72fnYhGuzXwBdBnLOiJMGNit0mto9e+KU/p1m8zS834hbv
T4PUUdwqnMCFfTH18lBZRw+QdO9vkvO4g5fORCzoSTyyy202bKcCKXAIf7OOrtbG
B5zGVqB8+b3WIc0/flBkG+5P7KEH3nx4joy6ZD++Z/u58wdh3NqgiqcvOWeC1OxK
rkR6FsmZkVVMga7IFscKPjtJZ2yNheY/HZLGVAovhicaaEpKOMPei4w3opmgTj8P
SdDrNuNw48Z4jkvjuWVIHpNZqeRkA2PdFVvrKJ8YFWuLOfV5PvKRKVsmomrW4ar0
mS+de3nqBkPJ/uQ5wjv2YKkQUXvG2WRDEF8fOiH1WpXP2am31AWgdqSo+NonnqO4
7M1CaJNTmUTbX+ifCv7+QasmamFBLwhAramDiewW73VVsN0a7GCMs9lNUwHmTbov
PG1M7ST7vLRFDVnW0DADuOEEnKcbX9Z3Nh9DJsV5ctZn0iKzq78VHn692v6hl/FE
5sUwNHgqO+e0QirISx/9bo01j/cgXctz8p7BRyfmRa6owxQlWt5zTEIGH9rYfBZl
nnk1S36p4h8JHtGThnUu2hOcDMa5b0NGEU1am4l5w8ABeT3q9PqzhVmrdc2Ov/4Z
53oKpiRz8yWE8cNynQUi0DzPAj4lz11knB3O/MXJ7bYwerkc+uBgm2OUkWC+dkYZ
7MZP2ybj9yohoaRgaUZ6KJxvf2KSyRUQjDKcLA6qEIphoQXRqfHG+c3hg/YFdTnf
aMxGz2eDW6k7+WVDDLIkiAD8Mv6o4QW+uiAW+ynfIOFZ6VPAi5G62A0i1szZP3cn
dUjf4K+bQ2LcAiK0k/DHH4jsfLkth7MjhjRIq++BNyiCe9nTEzJpy5hHCB8K/Mb+
xEtM23MgQFxPnXRqCsyw2v/XONcbW0QJ9WJRMsEV7yRl8prnmA6sXlHFki9pBIUU
oeuLuDxXHTlBTL9uB9Y11VxtzRdGtP0AwvCVznNE0rHiwn4dTUiWT89R6kyLRq6q
FruSQarNwact8NDXV4jZp2sAvmDTN3v9p9dBJv8XvCDKddcX9X3H0rgMqs02xtN0
lHWHMtdzeJs75/HD9TAhuC3ilqWOQ2WULHHwAkdrMpNw9vnihvz763kk4Xsozsne
jcekv7/Mta6dngXpB4oFGN/1EO2iYM87PlalQBwhXntqqfbFxHdfQ+arzVEoDity
SNKQK1vCt5qNt5Ss1Y1M8YYAWxvad85NrBnQ0T6/gZ2ME+TOErTRHngxDV8dI7MT
YANfgNKxH/AON27Rv/Y8EQAZQViv+hF9bkCEwAdMflQwfSvWP7sSZlk/30BljLaO
DAHc4lAiXK6zl4Xx/qYJfvwxHuxvAZCVmREHvUQZkzm4OD01OpFL+yeMNWRbuf/o
w9444Va3+GtY8kJr6XwMzGXGVeehMFE57ySObXpPz9+ZnvFXd5wzm1Ms50k1HONC
RzD4bz2SCZ8YDI0WoqJseMezp6IJYB/NsCtgBt1ijU2ck6QXBdj5f5X9nbYZ9vaa
A/LR7LD4SM3NEgiOwBxiLE/GcuvGakOhyGESzrB7WLst5mrKRMfsNMIqR5I+MmoM
tMdSyqJz7G1JMYcLO8ApJcSsLu/WY5eaElxaziGmhyvXu+APKm1Zdfzzliqx3s4f
x2wYJcvCBnSN0jWB815EK9DjcmptjGmCJ3UYG4owwrOVs3xDCpEiODAuS4kJhm4Q
fl0Jg2NylqRSWVhRBChXRGo3kbvNky7dV7KTcsMszcyel550el0Se+OgpYxdm2Fg
P7UBdAMIw+42BEbfXmeXk3u+nDWzG+lYodTcx8nbVXxcwKCJVKjIaG5Z9uMvvVhZ
KGmt0MrvCKvVOMZNqq6AMIlLymeHPBi9Su2wj0j/QHIQm202GOFgVWOK0wPPC3E7
hBaCWzTE8gZwxJbYjSc0UhZ7PGWJbsNk4Wj8eQ0S1OxFyCaTfXYqVOj1LleWxH0s
o6jIpoLxhM1Rifd8QFdVQYa1SPYGyBXVfENAL808LlqBJprmgAbfMXXsi2mtRGgs
VhjXkzQEvHUnzwMdt1Q6GDtF0hk2J+tj85XjFi0QMFDJrgDiA+3hMoksqjnhenGr
se2tTIznffhOD/wnkk1gyLY849Az7ePS/nnR0EZZgdZsgjFW8S8rMW2DbBG3zi+N
yUwOlc86HLpxMGJAUr3GRxKHHbATYyCQU0Gozh7t0XojxeOKVPFsWm3pxbUcC2yc
RbJcUyehTfcVOmZwIya/DdomtRWiWTL6v1B4d+9daXh4g1nNjNkQ3y8vW95Bd064
SOB8dr8CmNYBzvvqU1MsABDndusAx9c7JA4izkGy6tSF4A4xkQynoghwIAjruLPt
1K880ay2c3T1UtD4BlpcSRDNsZ35FVcS1MMr+PVOfeFD7/zzuKzSBYpCRhkjXr52
REo+XHp2P/ET14q19I2qkWKYFSYYdjHqeEizUqn8iAp9FFYNuswn/SCmLOm07WP8
H2nVqQclfXoYX6L6LtC+L5UAVfDiI+rfJfH13B2Sor1h1/7eXyitvYB751F8Ds8n
Pq1GT0Ydzwb6SVVEJ3RqerZUcj0vAynkQVcYA+OMEKwhhJqEnyqedS1jQexW4WQK
K6IWAxDHN7NHUNcgDM9Hl9B+TzAX2ka1j4P/dI51pLJrXXiazSnovqt2M+Nrsrxc
TlxZ86x6pCe2l9l0dwFyYqGIp9Y12aekEs5UlPUPqZ61Evq5m/db++O4VC80deNF
FQSJ1KGtOG6rLLvsNRu7EO9I0HlPV6eb0B0GfUeBnPNuxS2XPD16UiTruoBcbxO/
K9ZfATM/mSgDZUynPDdCT2K8B/DFdrcheS9Mhcgfb7CBt76I2+jCEWru8r5dWwZ/
1IhkABnUhHEHKNDDaGT9EcjcWoXJSpV9OQoz9x+UMUYhr1si06eZ8IaQYxwEtqYl
Coh+c3HIIPZbEH8FdtDTj9N9e/JGTV+GwNGgnQdLhpFBpyds7WpBwa0km6w/Bs+D
vT2yKAQMuzFcS0eYUTziVm1Ft6MaGRWyBRMPlZ73RDBHax6lsp/mfMx1xOEVP1Bb
eDsXCCPZxOyUrFDCUJdJWSMjcfrHjAxUPa1uaX1OfEZrI0XcDa2UJDZWelKL6JCu
+yRNDFiqCXkJta++PS2Z/VP7ZNY7/3TeIT7pX5YZ9cxww057F3YXWn4T5+c7rdWE
dOwmb73qipRy9gnj/7WSqCScGcT2wyV0qmiLd0R/3zGLlxK/kph0i8B0VBHUEIbZ
cRZr6/85o8est9bsx4wRNksPt0Q5jTUlS+eO+nv6YUnvB14K8JzD9oJqbp139ipc
a5LGwzZsX2x4eiVjgXYBhsOFXk/zOwhIgcharnusyxpQslCVCeOp9dOmj2u1x95J
u3Sls1GEVzY6RFI2VzSIA+o5qkwaDQ1MdOUaC0IpMpoex/nfN5lsYjXuGrbOAeZE
f3kiWRbYff11f4wmamPSKMDKUDWBgqRMzrqXz3m3UsU5E+CiNGH53IFvu5cSw5me
2CRt6KC8pyjZJ+aHZs78e9b3EkY5O1LYxh5A+bqD7PtCc7SjoqU3f0h5xUMByyo2
+RNxFMLNjbC4BSnCo3Mbc4/yMhypXHqVSNePQS4wry0Jk2IeUbHzdhLIG9Qsoqba
iP1OSBLCQnnv0edEQB+rqF8Fytn4xCEIahYlN52yVC9pEOGXpfvteQLMMeG4V7IC
Z/eimaa30a/vkIYjsq0f/w/TNi1I9cgaYn+xG5PDYIoCMRCuHfJ+kOhAYPe3a2N2
4Z9Xh4w+hmRhdvwshv+O90tx4j/JSFvF7mnCSMKnEiPM0lRrYRr5Q634MkhL+m80
tlYTJHraWuV0/dMttO/Vn9e73NGMP0rpCxMvEYwxLnBC3+lbKxtHTJbM/AbrYEHS
OiQRuuU8ghIgEVzrQ/ILp+sqHD/RE2eQ0x2FBSLsdns/IdKLtHGQFI9ilr+rRH40
JUyars3035WmT7BRRtOId8Ld/LSB8L0WtAgBxnbkhIxaduy2VeVU6UwJJsfA6F8g
Vvj+cRBX/lyNV+7FFBlIppaEmhoPXJpXiBqdMfZ1qTlXzO1spYcD5eeH1vKBFKK8
Cb9NeWrUW1sU9eifqcaXX2+1Wu6s5zVkq8VTC1Y6Z1oK8mp9VkBJ7Tq4HXaZDwo9
sBjqAxQNMVUzHYHMyn5XdkDrDQRYeSAGAWhFonhy/36Fiy/X/FstXf66C2zMcCCS
4WI6rHqF7WVvKwkwUs0xWF4m3G9C0fBVXRujKVdY7q9fxJGHnez6BvTAyC8wU2X4
X/1DZuAaWT33Klc17GxwAmCpbjhHSYqkq1gN1kZQt9IpAIkXO1Pq1J9WEHTYfpSD
C+Ee5PNXiT/5/RhUzg3hTkcu91lCdHsKRc93JH1xRW2izbY5xK1d1M3MI+OEOP7J
AEw96lwgg/muIBON5F6uycXSp8rVXHp3B9vUw/iEs6z1enn4ZI/Ay43W+bs+DzYS
ZcptvvVQ/OwmxR9aipvnX2Iguec/gqe8SmnXCEUTuvwjgw+3CKxLsTa7MRJAIAJ2
s9Kx3XlAPzx8j35hbwp64unypO4aa4Y34bEEUEPilJL5C1qfHcoBQNP3YOxQNkdy
UdSVwkIhYPcMq48qOl+hyksALRtuM2fND0lKejLwgFDl+keA/vPOyGa54LdxGIZB
PBgBt1/CQ/JKO3F+V93pHdDzf8IZaRO74TdedhALvaGzDRJLPq81aXJieRPFPx54
Sh5sip3AeE85tYKMgFKdXXSc40kLYOTVfL5osyVw99alP1yFtG91w1ZKXixLthTf
uQFN9nrNbVnz4uyFmiBEGdmvPi9hrJvHg2qTtjQ7K3D8Yu19hJiw6drqk4WZY/ZB
F96su+ZghiihI5fyZAF9SyP1xdybLl/XWv8dFnZq4kIeRU3YRiYMgQgRVmB22ICl
i6/qlycYOhi8s5GMIusM5QkPASn20iHwcYPWQCsHKwRzgq7RV7KpwXcp/Jys+bXp
dWuERKmuJzP4nnjJDnHoRnKYGLis5+c33BkX074SzWUaOsH4onUHjhMUdKIAK/Am
zEsfLrvUd8mChn/W99Kszv1UicxgzIzXdUEpydR19/dbmmMsbo1TQiOkG00Sbdzo
HF5kiAeUJs6Les4sozOFHCJSUQVGUPB/6CQZwMFzTRImw7c2qwc1zwE7eAhB5kaQ
El8UWMx/D6DpBMTEDPRUZydsRKVbhWyVt84zVqFrdAiJ7w4S18vyl/NjgugU3K2A
cNxEZIzQXHEo2y7g/zxt3Kl5w9AcFLiE7z7c8o5Cj0eYJPcIgIVF5JOYIjEdQefJ
4uWGUdqMeOvZFdtxH867cvMAzDmOxNn0PYLNVENaaYCPyMc8/D3MjgZnh3cEuAKZ
h7XoyUcuLWVu1tE46qqGVPcVRgarYe5xxj4mK2rRIPPOLp1m7YYHSFxCOokWs40l
TpgSqZavOpmjtMWVNhGzugx+ghYBeJiYDBSFpp2zpQyIeZQY4k6u35SMgA8wZC3J
a6ozgOBB6F6iAuVVarzsFTGN3NZgGJm/CTjPt2cZPoeNmgQsFwY5Sd0Jo0t+K2V6
K4N60PFGy4TmV1IyXHmqVgo2LNqrbvkTJgBBZUY6sIN5Y0d8TXT8iYJr5eTbmMfI
SOXaClw9hCNw1lSxObu86FICtA09XVO5AmM0kamE+AtH+uzhoqY30oqPomCPNeXH
SdYFgPfpms7vHSwoa7nvy3c1Tf66GA/KcWkOE3eTvlxCVuDpWVmOYwPRsmxzrGQn
uWihPg3VG4UKWgUxBAWCJR3kplgx4faTBsDb0ab6qET/S1n4DQ6jAZm01Xn9s0dm
Y3p8+2IxYBDx8tWpoiQvKRUIdHc2WAM34qrqALqZ+xJt6c84ItYLsWoUQ+aeqI0L
88nWtxRoMez6wLty20VZ3uS6xHfeyQwQBJUs+BfhXhWeJJZ1EmgsriT6qxDI2LzY
JV6dhkSIvFQDuSj8Fk9+Zo1hhfLIQugr9uZb1PQCC7bZrx1qbGgxJf3TbUT/9RqF
STxVP8oAz8+KBb7yEL0Z2y9IhHG4g2HlLElABOncunS2wLgRUSjI062yGsaTiWjZ
Zsnb643jLPyFZjL7/gpRdbcKqRaXVmjrSUsyNB1PymvGmX2QTjcWtMVwj1J50QKF
yAtQrRM8EVYkChWbbvKOreEi/L1EFb3vuKJlhHfyWJ5VHKNQHgVfSdgOAFwh4Eo6
HB6Ew1orsdPbGPw3Qy1FyKPJ9a/5DUxgqidlDoUg4duYGczalOQs8QV2HJTerWzk
tv1B8Yr9MoV+ZxofWtxE+XUsf2BKGxPokIQg7l4+5ptBYNsHMXxYJzF7+R3hk58n
ujM7dIT3Yf9iNAXPCniiZWzo1ajzwR2um0GrrjkmjL2Z/kT7uKjqkC7L4KCuBCau
PJH3GN1l9JZMMRFa5VgYYgWmzKuLd6F8H4fInNrJlDE2sYG2cKE3Seyz8d8cSvry
fwDarIMjY6yTpBVpdHyF/QkUCONpfPCeyk4WE7FIu9ZtDjIJ7gkbM6r/xjtpyKlX
nf87HlbXx2gpNFiNopiljrj4W/iJJJGN21sQdrjaCkgmrZqmzKzfTHy5DQPUnEeF
RX8Sam9VbEjWmr2fmMqbBBhNGV0Ho38fAe5nK3l3LwkJcB3Lg+c+1fI0ea8OYr8P
BhTJ21yZBEZ6FlPMLhBGHBzChPuF5INyrMIrn09myGTmuPT5TzzIyQcS6O208YtT
opZb0m0yjFFZlU8Bzufhiero6SpZNDBskN3Hh831SRkSRE4/HBubDQYGx0YdGiK6
xb+1iFVFgFNLUxE2Ii4oow1KaqMFJ0m9XxR2l32ensiKE43ZFkKUlBXROOESn8G2
TKB0SYgtfAvH/iB5dmfCYlB5JXN1k/yOFX6rSKWDwZk9s9wIE6My1B8VKkaob9ly
VkX0557Lz3KlXDk/aPZJsmYNpR3yltcZyHz8Dm2OHi3CrV6X9iRiUCUYYORKsHTb
zRN3G0bazr3BUNHtsUno3pYSB+zURnHKgJiB1dZtM0jfLeBI53QTLQBpKIB4FK9J
+RBu8H9/QaTrySqrVgxwquNU6liEAaJSHkrXJ/icBWDrvJNR6duHE0r7vHkSUPaa
adhYjkMF/yJgunH6ZlVA4beH4Ux6LTLcTjwkEcVQsN+QD5n20j4C/4mlhPLUZzoP
ca7EW9c1ZfmJT9ototTlWy32zmOaThXwdn5J83jS3G0/Be3zBfO6wSUKF6v1tG2O
iYYHumpDuqR4BNXulInvJYNLauqgTpAMaMT/uldga1hLEh/C2O1UwEWf1PjqcmKO
PuuZjGJUCuHbi+ldDnSDc2GcsswX3ztioNW0k39BAzwK/TAS5KkhwiyDDUtGCQcM
PgUl+0uBgWwLnTdlQ1Z2dPW5sc7vWxug+IQGngm0i6MFeLgoVz17G7ZFzkBBI0+D
0fbl7az1bphxzT7+XzaKiqzgdD5sGDxyRq0t6O4XexHJ2UdeCl4lGEW48wM7W1DL
N7tXmAR+qANwrs/pUaTh0Dgpcm1TR04deqTTj76rwopnhTie6Jb3xvJbPnf0mNeC
47OsEJk5CP+ncwqoKGMsPcCzhKuiuIPMz3ZQJUz/qjzWxVPxd0exQCV/0exh4v+f
lN5+YyRr8+3m/grPXlQwzAk85ap4t0z2zc0bArT8tQLhV47C3RSp29Wf/fZZJJk8
O5sl/HLcCJzyEyOi1nu8c1y3jTYPlj0b3IQqbdek61NT5sQOfvuBycC9s0Ooft41
6rZKh27EYqNCRIBejhQJHCOj9FRLaq5f1pXOWimnyJlgzM/QLMT5foXyJwY2pbFR
kpKjF+9qBt1l5rRrGQ1S4LhDdJK90uJkj8Leus0y4cELDlnUliO2T/D3thJeAOXU
K7aQZJqZF92O669iBc0di1kXjKMaBseRCnSxfsTIKEksOrqH3GO33B22lZfH2c/b
HWkoTGG7wZ14ppVEg7Ius/dgvwFVVL2gLHbcThmBjcP85ZKgB4rpUusMk+bBtD3y
axJ0Zq3Z3EHCQaI9SEmumyLaP7e8Ivs/mlz49rBap9SB5o8jcEPwYSs05+PHFi7e
U/DohYXdXJqMfKu9Ow4PBG5uX2zY8y6gI2C8b5KFD7EBbTcNG74hpp7kgXFmMKnq
oAbA87qQtav3GW3/74C5BplS9UrMwwu1DlEjElyCY2Vlyv9Ay3Y30W4pmf+QPFa8
mgCaU8AwCBvO+hiDgnGOnlU+QZ1b2Nzi1bafR2RuQcE3wJ8rhSaoS6jBSczUrgCz
i/eXIwNySIwy2FrvWRnMQRFTwILyPpbb7WWE7V12t2MhOzt4qs83QXerFrvIEMGN
UPGrHKsjZfjqC+XFQKGWL0QOS8DT4tj6abRe1BFn7n2Jqk1LCAnfV6WrqNxdpFno
dIa/pLVp/HccrtJm/kVyK9X8qiTYrq6xLxqOa2aUaDR+Wljo80ZgLvUGveC8j7sK
gmi6whcfRqQN0NCOsKl6EBCU0qjWwvS73aA16nRo+EqdKiKR/qsq82j3JfppLyYd
p4oJx1DF5eBcXrb1wwf+Yw3BlomMtTAPClF+RcpNovE3mWYdIh9or9rN4w1Ec8yS
/3hKMhWQbF0b/xF0xocpjnQignOSjCP3r8tnIa0KJ3ZbaOPTuyn5Vtm7nDBcHH/F
oZ+wMSKb23yUv1xpwVvvbrgmRDGZ+hwAsWYZllHDdArbxiJP/NTu9OUeSu9wvrXT
HIQ6W3gdZA2wcGZq4vv1/g3L2Kbmd4t12no2+qrZFc1LvqsPr4WLQG1guNWo3SlT
jiq0/cKnVotnbCFeVoGtA1ktecQnuF7sE9DELpkKSKIjRWUsvxQr0UaD+YeHcGEq
CxTsXkhHcYYRzRpFTyyC3hZO22Yw918yE2QR3LHNKBCwlMCD7VohNxYr25+VGYHF
gGikq53cyteXiE7CAZ7uauU5uflkaAlPVU9hq3ACzwI4HofzZ2OAhH7a6K8RNJrv
8Bo4zuTqK5KRIhzePbNPvgt7fUR95O/ai3HhC8B7fCbVq7yncS0nL/vb9Ybo5rJF
g5UYjwcVa6WU6/nBNTYqfMMsusdlDPJCLhqtJnfcRD+dj3IsjMxdYt9/jdcaxWkG
kfiZNyMQhRuoRucW7f7fSvGioQP9H4bDVyCY8Vxtg8Q/RUFe81tWTRvwvZKAgTs2
NnFuuvjmjuIXUOCE7Sbc3XboaBisErKQ4rbZNz6Dsj92vuEGN6lmkToAz/7RshuH
k5HFmN6SRR06vAFs8AKW3XLOYlzyGe4FJ+ho4D0dWsD/bNW9ir26m1O3uWttpo+K
KaiCHIFa5ZOwYw1vuxC2HA79UUU/g3nvKlN+HI5/YFR7LTNd++IfxHx3SLv+HkLb
cbpYwWv6fcI9Z/sJAO0sYn3rnl+ZPQHLTUrh9cwTlV7ej5qwwBD52Z9ZsSbL6jsG
FdKnWCSrtKXqmtgZQ6CJQbufFJDbmp+I66lbFo1vb2/Xlv4WCmKA1vPKgVgrGQac
jHjuCf39ayh9usd2QyxObv739t0H4RKKOsjXyaaUJRY0QOu0UhmEalQv/kBtOt0H
XhaoWC+02b3FVhEvVsxN8RntHNV6QO+f+QGya3iFewlWqe41K6NeLxhE2qhwW5XT
D1U3reWWvkI1usf8C1mrJ/0sTtI0nBLU+ezrCS68PdsMsZkLuwg2FYxqFLRK6r+9
/3h3p2vHOB10O9xRvsLwLslw7T+kFWr/DfmbY+TyvcEm6ty1GfSCLxFRkllHwDLc
PIHWdb1XBg5xCsgxixgO2inMr9l/f3U/G5RvhkarGT2GVtdRwkw19mrMI/41H7CC
dxcwv69P1RxpkQsZ7zVZvQRw9p2cGYw0S3PPgzA5rq9QxC+tNaHCYuMAfXtsuio+
irpoiVv8adi6xKybnqrnzdH0hPnaYw4ymAAvH0ZmtQCfe+p8KrR8CFyu0Lp0Slh0
oma536VmuUuwIIaJSH7vJqTQKiHKQnh7lve5qly9XGuiGvxwjLplMObELX1dEKz6
bAuYB9c3EUtbEg0KhLYUsVBoQ7syb6n1KaAWygrQxnnTJ5ChqLpxVIr+7jBrxsbz
xX0Rkvqv6fx7Y8TH5mhoUfgs1RIfjg/ua20c7YPeYKsE5TV5nyvIwMXohd6VDUsk
sj6er4Ow+5bcrSpXTV2TUP+Y/XoBdHrwLiLDrBiFzj/BvkH+7zdldIvvJeYUtyeb
zwemLWGptnzeCfXJ4dbdbLiqxUTUiCHrx/53MWS/Jj5jyPYchWev2hG1ghGdJysU
ZWSXKAxt5EwXxMRoLakobQiDiQ/iqJQyRQgfH5nNcOFYZHuEGc/0PgO+PfOZXxN+
K94qJp9jJJD9Zpr9zsbGmJwrpcFML1mD788XN0zLG69u+3XeiS/00JaDO/D4lJME
x1crmKyiC3y3nC8zcXgk2WzimMlLTBGsx7BK4727A8HXHvJksSSTaR+upfKOAlSY
TyV3Ofwb2Q04MsavGUGq8AQGTbXYGkZ58g33q+2WM73lqi5tJgofak2b3fCbWpPE
Q8eTCqOeZ0KTbmh7EJTo8BQIoaFIL9vixesIY3unWPhE1rjV7mtBbrBp8C33Cc1R
qF7JNJ5lL/+J9Un0uAZyIyIBStF8hb2bHnPfLNbprcPzEC8VAq4YVBwC8qYwRnvt
aoYgbdw2TT/UPVCYzFwaSt4FrRPyXQnr+GuRvg3H667CDTV2XBovdq4Cdz66KOGn
NvuZKSgdSqnfiJBEQ2hrqUxaC7JyVTMExTryOnPBUkO5fmOueM7ZXogSyRAFompQ
MD3jjWGjF3SgehphmOkQFug77ox1iUmAbnCd+Pl7O2JYjp45tE8Yv6ans4Pv2oMe
U5w9XiJtZo5/v2LAcz5eOwHjDIenhiwxfDwzJaWL0TyjnJ6g+Paqr/ak+w9YEqJb
oLg31dOZf7pcXwGq3z1qraJDMOcAJyxeMHhBI8X56SaTluHaoz8pB+5Wf8KvAybJ
w15/wMF1poiN5ycGvZNfBUrqnpGBvbBFrrU+08RtDGp9HeHELhO+XLDusXNwatKi
Wqfr7Wm3Nm2WnGFa39bBN7FzjPPelxkFMDWoO/xQpY3OYU8Pms+d+CjqJyhIQsRw
8PpMwrv1BXKOolLVTvE4vPuKiRv2ipscByHKL8cCJrbXOaq+S+dBXCQWcUu/A2dk
27kLecTyUqpEqxPwBDh8/gU4S7vkgfl5FWfCZBrxP1HsXsBwGaE8ablxyVFdLdmt
utcgVlgxau4LQzMts2189Cr1VCl7dLb+jK2cp6tsRGgPR6B32tRcPiRfVziEGZms
J4tVEe7xQ/vPnqOt9N8W5RSBxv8MKITqElJWRllH2tkBgXjKd1ITi4DD01xzIRss
71wibQQTlyUMftlX033FvWCxTcHRk3+N33KOoYOjNqXyR3VYmfpFMnFSVtaCmPZK
HxS3okcN/6oQM0oTgaX4v+54QliynF+2qbZjg4jtLfvFfmCF9DLZJPrrdnSnLaTN
srxYtpoUdp9Om7hDooSD9TBC9nT7vJRb6KJfWxMxJlT+AMvw4oq+W5uXuN4GMIU5
3OTUqh14vZ8osuhvsfOAE6RmGMsK9I0Ppu+oZhpb9DdwEuuZqXEQnTx1bVN2yMv3
q+ax4NpmGsEaW5PqlLuDZ0vS0/8APRUe6yrK5cHu4BF2Brxhue9jpwQtmVAuymIl
UlEtvxAKQzuqLS9HdtiQBt3re4SypSmUSbKVNJL2fkQltDR9J+XQFFHd9lr6G04m
tt3taMOOpr5CIsOBrfgv3lE0SKOX6YWm/r6KSclD8rp7oiMS2Ud6uzx1tbJlLd4K
rZKrMx1zU4g+2PR697oDRpBPCdgy4Vyjsjyc3Z3TcULamfVRuMvCI3XjVuiINav9
fwL/Y7b/l+ji9AOmjFK8iFhBIlVCcyo9cWrntOKBqmTqM0P+o4BJbP81cuKTmWBY
8nAhU0D8tVoTRXl9vhNS7X08c/yBVB5OepeVUMoCYtYbRX9WuiXenplXpCb3Up1l
zOGoBufpSCDcIiKM09CqRs5pkAtzxnTtOvIx2Fv/suP/q65RPZzeX/3JPKq5x41L
fXqKYqIE6lix8BWmVXJEby73F3GWM3hZVpUD2pCR9QgNo2hFDgacTZcoAkPMDE7n
T+QnZcGnZqnNIfN8zALM1uWaskOxjQE7UJ6IcBbNqUm58iLcc6qco4u6Cnwd05od
4N6qEYhhHqY58G1eXgZ/576E6xhNzPO1/8Qo/lNC8x6uGKUFpD+Llmzc4oDynpuQ
/T/rBOLeC6bGIgZMl6iB7krYBZgCnp00Ejhm7zNQD9BocwdX77cSnAsJlYXVRs2e
aXMS3bJtLhjfndben+cTJCvKtLxJRsX3ZL8MWyoUm6RGvwjU/wG2j/Nh2aNVf8k5
FGProgHY7rZNP0fXtfXLnEvSPPH6D94Qi9WOMu+NNT0FOncIp69IzzWgl7EpaFVL
5HX4MyS8ss8c0deUoDuU+Jor0XhVH1bcqXp9ZXXSZLRaXNQGrpvhRnlIiEuDCPDL
P6ohSky30nGT25HLIV633nLcdm0tBM4pF7fxFuF62IUtxOPSGLvYNlCe2+vttVN6
ZZVy6KxlGFMpoakb5JiSSYqnfCenpCp/ObqwW7kE1abAizY17fCgDMECe217VAG2
1MeQMoVLaFdwbREI44AMfQw0Yibp9tS1s8mpJfkyfWhQXAc/qEsLl6Cg9+jP8Gbf
2gWreuXTy5BQP//3jV60ce9ULeR2XmFC2H8vkf95u51E03tTc+KE4qJvRNBy+1if
/57z/txNKQlq6jBWOX7/VqIixEi8g0FiwSG8gBQeUfpeeggOfMMxvg1gMjikf9SV
2Y29UwQJfBNYBEhfq2C/iCz5qJg8taJRsGl1fCmKhUicr3eQ3GqYobP68DWVOHCC
owm7ST5kNNhPQGQsxVaA0tFOUhSN2QCSj/5HNy90KNr0rrvoky71m3tCCo+DJCu1
v5GuEMjI6QYjBNTp64OEzr5OxiRzZJKM4vS3dLK4FdIbrxu9lLFT8RobSDDtk5Qp
K9uY56jpVsEeUN7S32ONUd/UF1V0zDKDm2ztlUOep5UMUDCdOfbFoIlFlda3o3dK
aB7oOm3O+ti/7xFfBygU0DOwqT1cGYQ874u7MZpPheoFKpkQnEtbS0A8rny1jqCg
zz/PMNQrR3epCiQhNKHATE6YOM+zZDaqds081LMxrOMPYNwflh1XrUkDqoU7lfDp
4fENlEKVayH/9B0lEa/Bklj+aHPnVnibtQKd03+aIxl789IEEDOEj8F4C2g5QEAU
39ceG9JJRdMYrhKNz9iVFQfW+8lk0HwmNAWdAaqhHBFhIHpjCg75jqe1I6vHp+a1
NrE0La0eMecv66qgk7OyKOuP8NLjAkeLWDnEBl5NCFyGJK+WPxdYxFdV/3SZJzsN
hytPXqnNoT6SFMKS90Uq6iQEmXTnuBOcsEYkRK7QwsgALrXyHgZCx90Cr+k+lpUO
AOjoupi4MtoSYBhIrF4RNKM3tBaw9cseEs/qqzHBXKMSXeTmX3Am1GhurtcNuaWM
psisESZkO5vUr2fIvfyNUv1x0+UngtUa6TPxt5MNTPltOor6KwddWE88nTmhakCe
CJtyERGusI4O971INl3umrYleS4/cr0U9hMmiZ97/HDOKK0xtxkL+kYMhY2SfF+y
6fqVPUoxOx3MpFLTZuGmSQJUU/ny6tP7A1oRDCg5tJUFSs3tStvnCSMV835ko33F
7th0/Mc5t7MAFjNY+MUmPqaq0LpPVYqxxragHnVgXvTIxZCp22/kJRP3j9/e/uQV
hVbc/I5A7KNhiB9clfVOm6k43qHGEYxco+fUla9fk+L+J5BhY+ZFonR9A06+2uGR
XrmRbxAjVKLJ2+jnYRtHE4X5g5HFE2j2nDbL0/DQuFNAwDwSvcSurwOr03N3YYAV
vAOmfDvNaKHLig8qnq1FOv2mJ4TiRoyJyC0wCfVoSSKm7+06scmV5FPT0MLI1tGo
CixMulCY6PsLvJUwWmlQGYeSmS7ahO9WsnsbD+4RB+KM7xqJXi/Fx4sJUVi3tvf/
Tr/heXOE27FDI/psO3oAU3HKB2exv5wixpJr4chOumjk7nY2cca6D6SOxv+x9mTB
YUtwnVDDoQlXaBjGG6JkCg7SqJ01SlMah+a5Evnmwc32It3CRU9aEeEbjkR2DuCC
Hbemdk3pYh0F0LrNU6kWyzt5XmWagIJiDaK0TQ4XWBLO1SJRxzmxkhIhkZz+anLm
zT2Xp1gqLL9OFVmlUsNOwkUrc/ZJ4BchQrEQ5AlNhCfbgJvNRYoASeYabqVnr/Ic
u2UqzPgWkCO6DsvbjYK5i3yURRSDRuUJRk7txTd7mLiq65lkphGBIXRUmubjV5tp
NLhhuryYCIr2rlgXGZCWm0oIT1CIyU9NEgrKZ2xFE9Re959iOfkRk4Sdh6/EBMhp
ZPkLa3Q6ugt3XgVk50X36A1SmWHaG7qkhnZgm9+oWHMo8jh76WFeBRDrTg9PuOv3
elsNnjA8XPVvFd6T/Z1Vis8nkLV6U3Lj3ebrdmL/6IE3a6nDTiFo4JoEmg4Jov8+
cMizvVUmGQ+k181VNqbcCX27mpASyxtz7sYEV4I+cm04f63lhsqD1tx4LutWEzBF
l1EQzXa2Ou67qC4o9xThgqFRMdokb5rVsVky8S8kwIBq3EjdXrEP5fBufWPnJHXW
D6tsyFIwFI+2YKCdgxfJKLiHwXRetUW96q13mq5I4AQCClvBKF3G5XLiW40y9UIO
EbcS2vjSzm0AsRNM0SZfDNkGqTU8KDutmmtT6s/wP7Lqj2WYiaB7SUxBxgkCDY8/
zCn2DD1Pu0gEJclop0kNdjxmP+AKU4OjV09kq8NmXDbJ47gPRhs1ZUD0zsWpM3Ku
AS6nRtygdgsSNqAiWu2li+bMgKQWjK6nesbfcjWqL5PTi74pmc/l10ws4j5SD+ZW
6mYl7NI73kdEknRCMxNds+AUb3ZNtDmY+PY6kiJa74I174Ogb5ZdpmjwGpNDefPf
MZ6j8s3xGygMNFBNj6SPIMnmkjfj2akcL1dpKNPGwZVhlGXbQobvUxwEIDXfWhHI
c2gcPG+Uoj0Rd/uRLh4gGG2Pee+QVvbzL+UUN/6N1xrX9TpcLHWIDrvkAJzn4Ar2
hYWoR+LwKWpV9/swjH53Th6AGivoR9gsma8kT46AuyWG7gK5QZIiJLAKzFfoGnfq
+QK3hW/Q/az8xyEOlqLB7SFHFIEmOYlIpLQgMp74/SjaEhG4CvGwjg/GC0WiEsdK
a/mN+6BeVV2RiVIrYoFHzDw8H3QyN1otYU+d3mSxY/8a7HcXsTukHdJKBsRY8ahj
q3AH9xKviHQ9xIfogW/CuxlzuCO3mPombXBAfgcJxk1I7KF7NoQd2uaCU1pX044h
0eXA2rXwi2MDV3ln1oNHJGwvCht9S+geRdox2QVtZIE7xd4aYkvh7FecRFqgcNjC
sD6WdGHsb+PnKUC2U6Sr4W566s6Cu/R59L3nQUSQttPjyKf2+TeXifRia+trR+UX
SiDJi5BQwiZGJWh9h4ng1pNGvspMCGRlpfa1if/e6pGeH/hATt0v5IC/7+RMLmco
8nTEO39TtepnDD/msTxH8WhZ1IwwFdUigWL7Qdp6NBKMG6a9xRcTdLzvxeIP0ktm
N16OBfBK0ypF3bN9fFTAqFoOE40Xsxqetax2msG/0PBXJOpRsYjZ4vpw4fW/aU8H
RLB4PFWTBEhss8ENbe7lDXg16ld8g/n6rN+W8JYQP8pdNX6KCx5lU+xXPSY0eWNS
b0wPwDIhkF07TfjvVBrPZ1qAL2V+u+XkltiCzdXKEWPPGH08KbZlnErmB1yuB2YC
0ababZBwCvq2JcSHfjq0SmfR18jB4ho3Xr1Xib60YFZ4nc8h8DKceMRKgpxP1N3w
4k0BiD1ETmrt52EPdFIH5qu7SiOUhGRpfjTmFZC5/44DvpDUAC8gG9/R4b2/KMFU
4wF/ant1MW1qjNMUvJYcvnOpQ0tysterjmNKy8D48tZHCKkrXj4zXszdCVoWKtSY
cwX/90Zza314Rdd06RY63o8OVdW/U1hnLvIxOevWPUbK1Jjh3XUaQzVEO+k6TAmn
aBi0Ai8RpT0lQu16aYTYwyWNCs5ahk6yghaiW9CRnspHz5onLm7Mf/SAFkFV+aXf
u5S+TFSiYG4wOVIbcT3OjMFfyNMwQyKFCpODA7K+i0JASXasqlJwz3yP7V3abO9F
VW8Wn7U1/vvyc52qaCnP1aQZKNjLJ5bF+E/S3uIJ4sE4fGUMcw+/sLQk8elSzdYX
nx39bRqr4UPvxrrD+UxyVDxLLvhYA/2NAe0JX2ftANGbthNzo7bfUqoDdVd5PENl
YXFGosJTgzwLd9y4T8jgsuLOoWgFhVl6Rw1vd6HmD/vdlbnmLa+sSQqHWaKZUOn5
gLJSH3icxs4Tyb3uCX8cl1oc15D55XzYGMZN8EiRVLfm2x8EJBpnvfKo3xitCc+c
4L+mc81bEcHg/fBOLC9rcFCZNP4Pm44l97CCoHa8875t/XrrP1GUK5dP/PCAoFht
A0p2YLHkkr5VQDb/SXnYvEYmMQEJ1/GLIalG8BsEI3F3QN/W2eKAdJsj3G+irqBH
ebyZgMST+UJt8wNmk8O6Yw8JeMQU9zUakT70AcaADD2CZuTEZe99ucULLLekcU2Q
ccGQUXr17HPhxEonzsxGPwbykNG8Lmm6CtSHNiA5WCqNDHzpNlplRZK9/pfMdUSR
TGER722SgqvC7eTC9X5NMYbGYqgPAR6PII4dIhKu2LjiDyLcGuyCpGmNzdxDtR6/
Jc3z5ME0/S/L1N6kGDDTg//UrxT/9Hy+ZR+xNHGUlRwPdEkUucewhbBMUx2wFZaR
FDhaeSmMDm8xHIMtU0JXP1YHB1CjCdzFisda4FUB1ugZ79mcc+NefYN+AalxH5DF
10ekdi11n+Tb6ymrH1+PBuXu8RCUp2SOlmi6LQ3OuGGw/ycx4qttNZTKXgAV5Qvs
F6nZRgvQzdiph/jjYQDygQGQlb8RZ+MCqigei5pYWPisvKctRZy+0452waOL2t5u
/7R34bh9k2xaV8kY0h6+MXwydt4eIl7rjIyN05/HbWt0WYPmVhi17JiLmShI//bd
AX0YXRRBM5mn4smufSC/kotiAwJ3JqS/QWUNdgXHgPL45H/aS2PyDRJktmn4YH6W
lnzcqP9Uzu0IvL/2Yf4W+GgtCAd12fgN8ajv2AfDwCFqBmsqRyCAGKrNSnOl1jGL
rYelO6bmnk4TA4PTa5i7VuuShyG34Z9AvMcB/D2FoP7zHSYCUrWUX2xErZgnYXgp
w+Om/jaxbmtfoV3MYsF1+gsaPOwlGdTktVLMUbu0IWS4qfbhlZPLSRvDeCHpHOLG
bGU7NItbak7QtXqSGM5xCsXn0nE0r1XEtDQOQqW+rBDTtQPuomDOxVXOGu5gqDew
uJu6g2WPWw5QOyh3Ol++O3bzzq70571RWTB1SFVKS7Hqx14dTFfXNjCbGOGX9Rx+
xSaHbt4erMNT/5jVr248G2sMVeebplZRuKxqoDt87dEXQKvvlS/QWOCl5uNtIQK1
AKgvog6g/jF0X6U8nxq4gaaZTHEz/qdHtxNZr8BxJwuNgaH5gZX42ax9C/Fr9r+1
38YV+g3VNXi6b2A0jBc1VUQcmSdgLgwO8Zd2tRwImULSeQCES6CokBV61SI7Jm2A
U06ZwBOcqSaFVoK1nlrw7HIiEddgBlXSFnDS+pjysIL1P/wJg7jLCvcwNQcAL1jl
75TpaRRfH9HkdYJgef76NkC9rKgV5b9qtQsSD4U2j5iYu/9Wh76R7vLHrHVgt7k4
LYODvgHeLxnoBGrwaGMtGmtf7Exyoniu8yWpUTTiQXztGvZ8NUX+gI6ftDmds/6j
EThqBX57PiNsVaqoQha3CwqlB3kG3k3XxY+79Zvgas9hme2X4Hhm3R2T/VA/+08W
LOk4borNgpYGfc24cHog3fwnLATkk6oV/pxgMa7NPvueAzJlU0mmStgOCBS6jUH/
glPOCzuoV88JSDdaL47wEDyliwximItdQ+f9tcL3sOkMgGLlQ92kJ5RttLJHfpTd
WiTJGdATXK/PRhmpgc3AjAb7OYjswb1aumvuemL6eW8RhTnA2RGqH1/R9M15hEFM
x1XHf5Uh6UKkBH5LT5QWCcJ4T39lvaP3mD/HlLDX6EppcJf0MTWkUiyJSs+jQw1P
H2TMeENpdo2IEZrePXC344txh9VN1LSyqqqGvYwKqxYnuUecnw6mnBcwtvRm7TKY
BUq4RrmM47bVygbtfogdiqzxFBjzHukU3kXXFGUbx6Yq5CoLAuTEorELgPaxPjno
6WLfIo8MQ+kd9Y+G+tL9CS3n4dHAxp/rOjKiagTo403E6UoZ59hvmaQSN42m2HVe
44UBS3VvXaRBVJPxygCobeeY41b9dEMICA2zmpy4JEwL4egEURNSlGwnSrI0zaDI
TUOlk/8vbahilnpzyMhe+qzhw+ppbIEc7d8CFL0ClcFYoKPCnQr5IOLhd3MAzHhb
IV73MjAoTiO1RAduESSJazmwGyyEFz0fvyyRgSN8oaGeMuB16Q3tzufKC1dSpIFX
dOhYqnBVNmL95kVV/fqNE5mTpnP9hp6Cs4TlwoVpjCyAM7L9J1xVboiSEx5HXC7l
gwYyhzuTv3kJoQrOhKj+kfaNShzODrhDjyQTbfUHh1/XI6Rin0upDZg35VpZKDRh
PGRfvmZh2LUQ2pFancLa4tCKSiTEEvpwxl3I+9++YFrweM0cfrANq56+MsqOvxnx
0lusSFyL4JxtXi70VfS7doQDxX8NpY7H/kY3eaiHAim/+xtjk2JhhNhKTI58rPU9
q5rqcrEbbeSs5J1riLOThOKP26waS7Kvv2pt0GkXp/smaIqZf3jJdA/j3XWE7dlM
nWyWfKaIVRpa1RPEf6dKabPZaV3bNpzloTJFIe9z2uqj23vlIvhgBFzoggf9Gkeg
gWZr99eC8/2pL60Gso5rguxNe9NW3vsp1gIYaIAKUmwMJhyt/Pj5CVP+vwhcIwU4
IGNEFswMXEppaKCNVannf0QSiNrO4O6jT/QmWJcos0SLUoDYVyopVV2tH76fStzP
5Jga9GECUoquM4azn2OAphMg9w3rwcAQV0uw75/WiFcBTCcbCEZDCFKfUVQfEwXb
9WuFTjNx7NMlOKydywX3k03OPeYelUcrcbcdqAv2sOeELownP0X9/lg9ljGg2+QW
KlEoVvSPVfvvUG5vDFzHa2T5pnLiuD3CgXwgsUgFrAMBnyCGTsZFImPG58F1Qo/P
y/vjStz8Av3BghvpihjuWaN8G7/NRBJhn7dIRnhvDOWS4IFK2zlK76hwPRrkkl1s
DyN9P6hOLytTkkkIhWMU4ptwr685x6WBc1nDbaaRhGXCZ+1RBCuAO5n0DoJ+gGlo
HJXVNdJYmRQCD0yK70tjKdX+HLXs+Bhy6R5xy/jC5nRyL4JdjoRFw8qlpek/R+yc
dGw+08RvpLglSwA4hrBVhEcvacsML1O3o69RJ2O3Cz5wgN9mUOCJ6Kaa+z2Uteru
EQivx10JEFlL5a96Ro3cVss1QdSNf2M0Z8chwFVyLlZjXOZdc6dcKytC3RxGjrTc
whvD6uUPRtnj23pl6vkO4MmL9U9lyZU3i2Z6ejk+wxnMQhjeSE7Scs7zE86/gkeA
X1OhLIvQAOj/FfZkhlBkHnz6y7zi2/UdKT9x4riJ9UqPpYapA0jguqKoTjH88bX1
cD3K4ajvaGbu23jJijrCvEbS1fDNlQV3HO1MyDLtc20SCZnA8s92jQRyRuw6N+ca
8bN7Lpn6GEh736RUeIX5+RoyCtpbtbz1XIGIsl23ljRTRUecW8wDjmJAlyLq2pxL
p2c++FU6sK/t80qiPSY2BLuYkq1UQ6GHPkPuVAns5zeDr82/RzB3c8bftSbhB97y
IudgfdFDOv5ryfYjJhkLphFCAL2nQn7GXZGjaOwtSLaj0hnDUyUlL0rXWKnUPKFW
DfcQnmcIZex8Yq0olapNU8O3xeZo6IlCL60cboCVdgL7qJUZRjyYcBwjlsrtVHij
4y9v6UGKJV6iPE0Rt51fHUlnt+sdYKw0J6yjDlXyzsYKBa3jc1hfL70B/9Dze1dl
kxkIjItcQgtAu82s+ugllOrYSxZrvr/bEj9c0e/WLlUTxkBkFrLzntoO2QY8ccpc
sdBQW1zXVmrhC3pUy7VXZ6JuU99Y1KFEgu7D1Sl8cMSOfCQYbVGCyXtctQXiA+TR
4bBCrArPHo1foM7PhYvCRtlr59oLR6YXH/bQfdfvgD9mGCNjEHTpk/lLadwjhIDU
yAa6wuwARpJ0itUs2NtaRwCrW1OcrcOeuWyzQDz04A0VrXqXUWNl5h3Oe9UkpOn2
S/GB/c6pMWR6vz8QT2n4hsu+wGmnwCu/RZCbCSlH6vy9mdRyLxuSxdtx5GjVEDB/
CSxwEiZIyzYjgrVwDxZyMC0El2vj906BhqtBjmUyWSLyqWUJkpbdAc3E6WKvTeEd
lA2qS1XOAFCJ3Ms75eZuzVJPeMilgzkRFgqnoyVCije5cMOcEb71iyaa0xKI5zMB
AxgE3Qqdhh0/Q7k7PJF0tjbHrUKqs7nxZ0FrhbMtOIbIPTOw4fmctnoLlixCjQlB
nrFGQUorZmXYhUZLpln8IFJkQwThFmy0edPFD1t7hsABQjwgkSynG7chVu57Yyak
Cls5SLKUl1SOeiy3yu63NN7s1Ce9R002hJ0lBaIKDyLTp8ezj5bN6fBh/YbcAbDF
5txHzBNVByjRm7/oSgQFSiTJ2D0xzJQEuqChSzFm394yUgZ+B95X9lgL4t/GSXZW
B3pAZBNRjagy4Zz9XTaaVpOxqEc7wm1uQT23g+6ue5cUNXgGXRkvvj4bDcEODr2T
CX/y/u1iKdfY5H3gWyF3Mmzq4Y8RU2xWcpSVeRITdPpKF2oCXAsTxzRAOHTCx4F8
MPe5MY/tOq0K+zup9qIWj7HNL9wFtfayWxpL3HcKxwRKmyc3n2NWj6ljJtKvCL0H
D9/uNtSALgw4KJrfZZiExjA59YpP6+n3uYPtbwyiYdHyWlwZLm0CrXP16T+O2cJq
E7sts2vFQT3Hh1ok0+wIo7braXvJ8GPOjhjq+xowDglBHeezK799CY091dCZdfhi
aXiJUtWVfd5+WyFnb/Phve9/xSV/tCQbeJ0dsS56GTP4oS6nHCenGXCXaI4oM6yR
uwxpSTmbGK7I2dqPHgoUddU2ASMI1+TgBKLcmENSQ8KlQ98xRj9dfGr8USPlzccV
BjpDogDQLBxuvzHntEfFn6ol+dK5rdl43tQZmCeFuL3lUmSCHDc4A0+xJbmU+FeV
hBBPTe9yPWHBDaXnKtxYrBjLM72cG7vnhv6QUyMY+GOHeeJHwmA24wE6/tz3StMu
yBz6zAG3fKMK1QVleEAY/CgukMaxB4FkjNi0f7d00Pl+8XhuRzI+fpOwy3Y/hR7p
ND7r0cOh12tFIAU9W8X2jh6XAa/OUB/PiT+GO7XfCxXrR4AxAFumDdz3asrhVOuv
/cT0Uh3aeCl0IwwzbyoWLJcHoVSVa7ZWTdXfO4+TmdJ6JWPybEfOny0y8isdfKzv
98NN9F2wZlOFlaHWM4LNFeQsO6N9+0y9HOLf2KRtSslTWd2Ul7DgkC/LL0RDxTAQ
ra/8Afov2UPyVNbDEGWuzPkTGFQ2NQWEt04tHeY+EOrvOMyhBERHyjbZmp2ML/eO
f4PR39ZfMQz5cWntHvKxmlIsOTEabmB/Ovg5Hbfg6wOU89EX2GaK7eJHXIDOPD2Y
tte1KcFYCN2ioV3K5JdXig58yE91p1Uw19b5OBY8uQ5Rj1wdEAFxYsbP4bFj9eti
pVa8oi6rKjH+lFgBgAeyhQiLT+C6hNi50rndut/M5/72GO7Dl6Sr/pePmZX0s3V3
gr2PF1KOLjEZWO49c+J4yBwkqMdNQKqX0fZjQWFh8PiNEhrQDpmUHkLiZGlBsQF6
VTVmrRtw5S8CgkwGNia5p41TapCySWDMsKtQEwjArpfyAj8h6n5qpQqdIdXExKMH
958pSwD+5tPN7e4vfBkmw62azTfFv1n5IxFGMj1thC1Xyt/jdao9qxyl6yUEqum1
xCd2ERbkwl+hTfMrPn9BiBNvc/hUPAXJEt0gW085IQyke2IZpywpc0JET+wzmxHO
pwo8GUEClUirBIEOJ41NOb8iAVREBs8iRhLMDniDfqrhr+ex68fs1kPclgsVovLC
uKosQF9FXXHpdrxpICwk42bXzcw0TeaR9UBHWydzE5CM8Kf3WDV5DWuHhtAamg1h
hOVJfVm7TbVJ485cPZLyOFSGo68aNCb2Z7ggklsHT2uIw4MyOYoY3tmIvyxnIpcz
2Kxv1Y/Axh8YSrnn6tq9JIx2fP+viA8iUKuhHCTo4s5rTQdnApjR0XT4DR79K5b9
KZ/dhqhy7JxgMY1LXvWKsPyg7L2UfoQnFpH1aVeDQCbbrVJL6nwB1JNXCFBm8mvy
f5koocYH5QIskzi0XiURjemncAu9m4xw5vBd6/c2YhS+yKPXBto6Kd2hNZseHoZ6
krkHf5srD/OxfxJy0SPToUMwE7ovLIPBLa3crY26+jjTt2+IeDfRvIY6YwghM8VV
T6ah3QOnbooTHVZqJLgbxYK7IwtxO+SzKeKc58N1S8LwblfsctULCfv1f7mEZxHZ
fKceSNESRvjZ4LLD6C7Tev2pfY/jSc4YA1Nb1EXlSjDyWziULbJdGFTJFw0x+R9c
ZtJv+8hVjnX6oQH+qi4SHoDTDP84jvgt0183WMfOiLFc83MsfYa+Ccwy5jNBEZsa
i/nBUGuv511bY82HtjJ7/tLiLGgMGAopTec1KHXIrDIt08vmn02GROTfAtCbGFnW
1PuqCg0jW4npQHPNThQe9B2C7y5NjheUsfozYxeTTod6T2QDawnJk4Ra1swu3/Ct
dQt+ZQO8gzhvx4lMXYtttkbaDpH0nDmIjlRxMYwSczVi6CU9PeCz8WpjNfP2KJDV
65AmZyyjlLLNZDGygkC0aF0qDgisSSWtddYPCefP52PLyq6YsNFUHN0rlriBexkl
8OgdG54ZJpBjNO/wkjJBjk8zs6dk6puy+JqjDQwzoVjvW4flfZdyaPv7Pmj79s2i
JvWQ19RaIkB1tvH44CPfhujAQojbgTpDDZDAdXv82BPHo4g40ILfbt6HaUMLobMh
w3bWlhHMxXADOmY29N0L6/gLgvk37//7zPB3uWjFURQAe6ulZJkYBR6PWKnPxMLb
y8QeF99x9DMDbNtIxeubXoQWqCF6EWe3hOsFskF36WYh8iC0PFs1ra2wKjvrG8Qf
PVTGB6zKUilJoC3lkKyNMS9sjk7qCAzeVafqTFC4Q9IxXB5IlBtrTpSc9RhfdfbM
yyDgvbi4EnBlmF6YK24tYtdoHkvh5jaCCx0FeFKOk5MDPWgXhBQDwwnnBaY7ZmHM
WHQrQcvnDs0tgnf6cfCCEIGEfUi41HuIZIBuq0GI2ohAxKDVBdzTtvygj6SdAY52
0ao3lgHhQYkopMwzPap15TIUbQ5iwplcoUNTylMqsMrFFhnDXP9LnjE5DxdanZ/X
mV2ZKStjuk26D9HSaOZvFFQTgo8n2x/ShdQEUeLnb1qn8k33v/+TMEzOG3P7qtUP
5KbP7WP+hxyRdUoji4fXiOWP1zhLDGZxgGVolGNX2B5uUxrkYWBl6f2JgenmnJLl
ZGxy1EKt53h5wO2lxWGgI4aHYwBWTxze9Z/YGIo+CE5XzOCQKWaQmfM0P4rFKpnd
nAJ/KCaMPCReVD6Bvuyj2O8ew23ALf3BoGzZzNwgHjAp376mK1jPivLg1aYlwjAr
tE87k52IpXo9oe87F64NRHHabx3P+mjuAzxvLLHxLjLF3qhnIs3KsCI4nkvrIlhi
ycnqZ8swc9hjpIgDglmKz4y859XYKxj9wwWhF7xbXuO7DVnfZqeDUVHaImYGlgJC
DJHRERQif3Lb61SBpaNoyxFSz27HeOb1DUIQVKJ4YNSsn009v7v5hNgFU04e1gcj
ayhnwEJWCB75z898nIPgBlDq95OBe4G+AY6ebx4BZ0DbF6zPgW6+/LH1W2LnNhoL
xJrkJmOklxm9BLWBeSVkTOg7mjYl3/or0CAedLIrwmOyFj7VOMG8+c/LtQRjl5XP
rFakEbf97FSd5NZY8CU7I/vKcdaZneR9BWi/gS7aBX4fkJwZlRvPYCI0q8RY47XK
L3M8/wDBxNJGIXIT4JICP5ZYqvUHHtHRp13FJrdyqrL+xhsBQ8i7/GGjBO1SYIcz
LP23rjDStixj8+LS7RG1kaU3iwVuY2kJMaCavqL5GebCAZZ9NmOtm8/rF+mNdN+7
M1q5irxR2gsC/PXhMpx8NPYPOwRCwIPiUSUukgYaZPN/hvi1HBfH4BVSoR+wqnGV
nKywKJDow8y+UUIXSo9WQFd7mIvHFdlW5V9WihbjV5zQkZA0OXwWD7B2zxEHRVWS
kd1N9PiXTLhy3nAKK3fvyIpG71qdNc97jD/t33avzUKm9FAyBF9VO5wWClx55i6b
fef/yKz4fod1rg6pcWy7pW1x8amkdQzEhNWVxbMjYoL52Bt01m393c2Sywoutonf
6yvs92a8YNXOCkYaNXn8HIdVe9H+uRx54lnjO/hjRXms8qNLI8tJcSM7oBHgsvEV
XwTBTaRuA/8xi433uIyQzOyi4HSRGBeRRf99ttBkPxNQiJZjO4wnZuSXTZcrD/Ou
gDWbJRFg/wZO68mLbLglobs1vWjG/qS4cE6TWGpMru6ggXO39i7ev74/3lYApEJX
GvFg9As/iyOEXRYPFU+lDv9ZXGXImR2tcW8YwRDfBSw/Cnic6jLXaMJxu4ZeNn6V
8s3N20Vgm5J/Dbft/keAIl5RJfOddy240jtmdo2VUjBHr428QJ8bXzZCTNQ3+uZk
JDGSOX9Rof5OCAePEUAKekbm/SvIRHhaPE6DzeF1ZtolwPAeFmHenF7BjwvYsdiK
t9B6wa+sNi8CnCUEFTrJXGovsTtJhnCc6mphA/HiFadiHracNDRKetSnuSdZ6Ciw
vFachN47o8hWARE/+AxqlK4sqBhNfqAeS/BkLjkkv0D2hWCI1uQ6VqoVcwgCbLCR
3e6bVMoBqa83XxbuPAq2UJzLbtkRcYb/+P81uw6U4ftLMT4Aa7xs+y6xOGCKPA5r
qibBtQylnt0nGCn6VlgZYoRIkXVyM1OqN3ha3qutzIkRTWMIf6To8O57s5MCxB2L
FbJJLE2VklXXcV6Rs7RgrA5qLyhIkHJrzVExtfGeNx6DiTYO6kFw6Y+UZGIrQ9Ff
hZIJMuLcZ4j/GKZK+rvM4KbHOhby0fWtluxP2QQ19bqmqNOziWnYxS2XipnzxwSo
XzRSTVT7ty0vOQ6PtTX6OXHCI7VvaPi07SeOtyU5G12/qOY0WeiTkOXfS2wsBwdY
MJhO24Z2SpZd+X02h0fcpgka43up46OQLxOoTf9bNzNl+fbz6KZ5S2y8N7jkBbCA
yWAfRk4AkH3ijClsNsymM5zM+rziHAcarP4aKhhfKV2veR/GijW6ftb3H2P8gaHo
zV7ZFDPcM3fNxkvr/6Kc9qgDGYOiQe2Or4l0IJavjqo/HF+mw+AtyLbINDvagekY
BQHyV3W/4+NfLbGUUaCLv2tqhQhY0hAxkpIrNPXB+6lQFRFyMlzwRNQaCDlC5vb+
rUw3KuiYu3ojWDh7QnuPElBnDJdqE6D7Cp+DKswAZXzh0YZLL5+t4Ub7nV6kEWPy
wI7sBKNrSOs1aZ+EGHYi5sfjx6Ui06zIJDmsTbJO/N7vyAa2+hytWwZkpv6zqTUp
KWdwmnv28lzMuPl3TcKsyrzL4kxVJHo6Pz46SOha2NBozlvl6RMKDffxnVQmmE8O
FVwNdtfz8/VjCCaObBwf1FDVPbmKM03hC9UDPy3lAatzd1J485xYztDO/G9RjElD
ZpvT4onnwu+pb5A/KHtGqid76J+AVwNDJmab+zC6bI4sCLJV/0Ekrot/jrP1/xhG
kjDgAQJPza4d3+ns1BV1JV2ZnCedB7bYH3hiSRNjlNgViDzAk+Soi9Sc8rlC86Uz
d8Lxhc0Tc/uyC90TzXDXocWCGY/SlEqSy0RrJekRZw8qT7LnKeVl8cbWKKC3IZ/+
2zzUU+B9t9VfpwoE5Ke6nq1nLrhbmT8GgQV6+zf8jGMRezUbCmP+XR6Ca1fNVG/C
NMOcl/XX+Ns8kPluXAyjXoSgpoK9wwCdNd6HXrAgLrd8nMmZ9p9RW141EWYY91r9
1vrifnPBQQjUYMTYwPlrhqLPW67MP7hNoi8bWiy2m1PyRsXYL3zOqlLQVj7oiJAY
Tw58lE5t/h0/t8zlZ8fNgWj5N7IMJDG1Lrm5VzCOh5tPvuUc2/7uYjEIsrujFSnc
jzTFvA5vRlT+AKhHGoEdtfdk+MIBXO5TUevNOi3PxLqIivQLEKHq3pp07A78ba1Q
ZUk4UjUN2PfVtrReXl+tCdAXMllSlr2MZAy6qOq8L/Y8NdhXpLtS8YrJY9KNLwsC
/jCbEClnD7gc3wu5JsEQoZNKwcHWTVQpe8lhjRF3+apL0KoMEn+c+9lGEZT5Jh9m
2LXbhnLO+K0lzKPz6O2ThLvzvpYY5PEkib4f1tc1zq1i5cqSNGycFjPX4Ufzvwir
oQlXhAY3dmIWjm3PDPJSqMpMSgKFX3Cr0vktTqh5J7RlFm2cJcn0X3BYgcarFMHF
r9O2l3Hs5ETLO4KqyeFxMmBeTOUc9wGcopRxA43EtwwpkhI1w/5KAn4h83LCWhDZ
s5tPDmO0PI+gB/CXzFDLQXYh438+nIlVb4LGt6G79nZcPwvozbgg5oHzGN6H9kfI
BOjqUwlgk3tK3h3h97yxxE5DrT6/8R9BoAiCICRneSYEHYyzdCNXtPmVZ94/7tKc
l3MBkTQvChZjMG7A3Smi2wybXsxmDWyuGQUfi3euUGhnL/mtF7YA6oeHi090MRPu
XN+TVLvwpVxMbkpxMc6BJY1UvpxKG67rzXfpqKSvcmWM46kPGJIbiOBFfYhucI8D
y3LLaWXH4xKJoGBsgf/HRLatOlh4f+monPPyv8jPV+FTRyaU9KmF681BVa/PXpq/
Nusu3BwVJ5cXnUbOM45ktb6FkKOaTaiyaBzm4dHzH9H3Ws8b1bv1SA3qU9q27l/I
9ZVVmmLZJFERW00VOh5wDqLXuxaImqBjg0Sy3+fOwzEyyLyQCq1KWPPU6DaY3Z9b
Wj/sNxVBCDOd6FZ28QQ7Z2bZJ2TN+V1ZX2/aUvYPW5Q5k7KI95zkU/zXoxjH7+4/
Y6dUN81msAwk8SG7qHLc0ozF10aEjv37IeizEq3l59rh4E0BD+1Vd+GSEHuPbbHO
UTOqIap1yYtMnL9mcWfKANweEmnUWIqE4FGyiohWo9D+dTUGjUjnhMEZCHsvp56G
ylJslDgiMtRfIEywIcod7M6opZgaV3wcMH2RRoVubSkpq3Gm84bWMsZ1sjRK6rfS
eUkpXw3qxFFuKiyuAeTwKotLtYtX1GkLxt61V0EQZi87N4GR9afmYKzwd5CG87Fa
sg1mEa+rrH0fSNnydtTf/kfQTPfiGMaHFyvY56q+ytKHz8k39GlsvbLVisvqhDk4
x+PdayBVnx6uzc5KH1P2b71ST8tu2uRm21q+CYbl2+YvOpe+umibPV0SJHtGXPWU
QAJGeJxhT1n4Py4gXGLaGwpDfgGFU+SaCZySIH9vdXmMbJWT+alIHI1Sgo8W4CgW
ZpdL8YC4cB0V+InRQedg/tDAPE0hBcnuPj5JjtPTyNyDLDxAMuboMeEoH2NhvPD3
2/35AMMXsdU7TCw2BFisVJ2xU0egkxE+K5vqkSATWj+7MBSiGA9ZFvq+a2bQuNVA
Km0rfpt+XVUiBLHtK97pUaYGQkUhFJlkf5oBLHnoowsSydZbac1X2bS/CcBE9tBl
4s4MEdJKmplL/4QtwP+yAgKRBrWf76M8i7oiCk224Oot1oNcN2+za3AMRE1sQyYf
PKMEwWaHraqsiGu1wYDaAlSV7CpkBvRmkOld8w8RLkBusYeNz2Z6bZAApOxj9otK
eYpsadrabTxWRVyCZflrmYxKvnI41wbmLRjTXkwUOhBfMLa++T5YPyMHmrrjNFeF
HkKRSyBntIxBGOv/9bkBPMjVhFi0Gvm4TSwxEQQMGYLAFLplzCGxLX8V1RioP+i/
DfDjLrEi0qzVtZsYx5seJxKRdfIIJttBUyLGJpGCWJNufZgRA+TR++A1LhhIN5UM
/5lUtl0XjFThbo63DnW/OhL4JfUSVmeUCYx+mFUExsUlRihwmSifd/tGZRtMhATn
+GqsSCxgvgGP5hCmVnB3xy22D2BbQrxy7GvoZsXtf8g0feT/23/m9UGm/us560X9
qT+kz1Lvgim14/NFqmekI0AxKkIFXbjfWuUxBn8ClNGEI6SV15Px8dA0ZRsrzlWl
GK3vzqq03vL1PVQ4bdcqD6rj+TQ0+PGeqG11FbG5IJyCsWHzyWc8pzVtfJyd64Pi
4TVAYNDVRM1xbdEcdtIqk87BUnIWPzD2GDfYnRL/c4hl5F7E8gNW5XUR0c4TclZB
uzC4ys70h9e0N/kfz12LNELV0VW5JRMPsmkMLaHCC7ddXTBzTPsmHOKb9oaeM96D
S97iwjEjWpIkeu4O9p5zKM3VcOpSMJ5OX7pCg6R5YQaDc5PBYqGhg8oj9lpEP2eC
Vfx9Gp5FOK4MFMjwG14LaCt8ueo7zIZ2RxKZFCAsu5MOInSv8VSvY8n7bET4m+Ob
76IRiFdtiw+W8L0XmyGltFaeENwFhXSVRAMo+DebZ4ky3+Eft/DwTq9+IaLneQrl
gWj4CR54FxlGvnY0BJ50Lu8bDB0T5WvwUIPS62NI4dsBk79NRv0I845DaCH2Y8Hk
7GDBA/CwJat/LIKd2hGJ+FzxQDlTVSOvJP1IdoJJB03+/Izo/j5czKdI1SbhxTSy
V4pDFA9VZVjrC6bGl9ztfDXhdujLtwCrl/X9rkgmhL9FyxfxeuU0A3BP5H8RTtYk
NFJvXsT4uq8DvoQyWVm9CIP0luqN9JOIVu1BPqfnEcx8R7dIKalEdKFgNfGwDYO5
hKl6nV2+sne4rt44gMXF6332iAIRp3MQh1Wfukdgo0B9DC2wJAIRld8h8q3JiwT9
JxB55lxVeySUf/Y+Ilx0AOVMsR7cyrHL1tI+PLKe9PIQMTArPZF2ip8WNUl7qhYG
1hgnAAmumJWK8JpfToKdfllOZTZB1FPY8qhJrBOdxLEVQHhNm1cUzO9cQ9QrGPrP
abd+EAASBV8QET9XR929SKyFjOFuLBoXjaPnsF1ztAeZhshNE0oqGZ9mzDnmUm0F
6E41BmCe4hfHvshie8VNDGFwwsrUh98KbVam71iKGe1yZ8JyLj3kSTLvwO20i/bB
M3z5kHlFrz/+5sPrlhEj6FF63jp6WBlLCoqKHQpET1goJFWXrXiAERwPMLsZfIKx
ykqzy9fEH8ycT0mc0/e18XpSZAT0XOf6GIwN5svgpoDWDAevyg42Jn2XsRDdVANa
PIYXtpdmZpX4qzdSrcMxbb6p1NbHNn747llPppyuXE7n9Kb638UWOQFKWVIzLx46
eeJwItYJoqVnYDQSvKo+qId/bGHU8HwUSvxedCa021hlQKk/i6cAR98YIIEO7jfg
76kO2VR02ZOyCuJoJzUTegoZJn0QbJOqppxq91bk2i6bKGE40XZ556/LallYkNeh
1/IdSKlivDRu6B/M68mqvkNiw0t723LWV4Hu5BGHsTGoW+rVgfmmx5mrTWrOoeKV
5aR18wK+HpDJXrywAJ3/DxBOyRgf37hE4cwaYiEGqgmDP1mFs/TNLQvmZ/tkNgNr
clyR2FLYJnDf60KNRB6kX0B2+kzWebkLt8E1KQ1PypenETuLbPG2Bp54w5Z21e2n
9/1KdNxcF81pKob673tgh9lkw4b77U66v20/U7nON6NxVV5Y3peecXj+CnEQPAdC
1mT5w5t94rD+1GQTP1CsP1eUB+DAVEu8i/9sd3OUvCmEgubFCglxqLUMQHMPjZEK
M7BwImM89+V+pfrictW9YCdLXJj/9xSarXa017aAGjmdNB9hVVDin2ii+MFks5WG
yHXOyuwKg7+JFZ4GCyDVWJyfdqJoTFTkrohVJvONYa2x02joJjw1X6bhOytvIpmv
ibwozh/fM+iy6KK/UwOCBuFF250diwoWxEamprPuGJf3RtXwMQgO0A//1kiVXt0S
TGFIIU8z4qw9+e3//dGdBvLiaOPS070wPo1T19ArnkRuyVyjpMjGrAIdcL6O4lZy
iWw1YbwkKgCiGLqrGsH1ICi/i3lhCuRSKt4SJYfIecMcCwOKirwS6ICHhCbtNFPQ
Pg1YMqzVhhEzVIOg876MzEi0xIAAa5AZk91OBC7gpcj68E0UU/4LkqRwegjOFS6C
DPHnGwFGQPNZL+MSlni8mv6yQh+4jc51SZLRz0pbF0ahDLUN2fVqStEdYNCRI/xx
nQaqGCzYPNAcM0lNRYHeLfoPNg55LPyr68f390l/W1oyvp2x58+/jtnC+Koiysy7
IA0P5kQxI/NCBGlzeujkrunT5worNw0OMP0LiVBC9Upg2yqW4lKVmxGnN0/e68VY
+scXKoZ3Q/XpITJV8JIR1qn48U4m5P4PjQ55GLsqRBSXvA5pP4fjI4av+91Jyy4e
aCyuM73X6IIvo2qF6aF0x3yBOrquqbpDJr9qT8CPsCkW2rniWqvuJoTtuBH0+161
4NtbOsTgi619HR7hN4szGFcOspYUS4GfWN2S7loi+ZfU+l7N6Vp6Q8rFz94//ZLG
93JzvbEXGjxxPKEEFy2ob/DBcinidV5ZQsgw6QGe+iaFsOIdoEYSNQP5xPKb3fA5
C/VUNhQ3K0T3yi08aWzvVlj9711Jgew08zHvB8zvlrbNVdUDgLkHkHJAwofUI2Td
v4HWIAAGGAb9oqphprdnxTltXKzICvAfgjMz/Hd0zBG63+dm0ifar2zI5Dn+bZ/Y
hQqw+ltASFrh8tcKhXVjzUYum2ZWSVwFOqDxPe5stNB9gFyXOgCrqhtRL5ZvrmAM
s5nQf3mUa+a3aWLliEooRdNhlWlKALXGhUKv6Dn2LReupfcMgl9ehNi0vIMK1L8s
JGntqN8JfNp3Io+P0cR0gwNpLS4/bESYNV4r6EtWQaB0wptdVaWY2XaSxyyTtzII
QeaYQnBg/iLpG2ddiaPMDG4x0Fxy5aubKBAITiB8gTnb3kg3tzAGfIaMp9d+klCu
tqekzbVelomsp4EMVTrav2SeZfwKJbjrgl455aUC1w7wdBlMU4u+lEDwbowQFBZ2
o+xIfhX/AaCTumBjHQYzVPvTvUXcCnop2zfTmk1FSNla9pgzaKu6MXXb6GGUt8C+
ktOxakHtpzcnJ8Vhmm3o5ngwwWRFAJGIFCDqU2QVSjZPt5Ya1cBfwxr6Xu6WrkcO
8oDJVCRjgFIw9ZkFfoVBVxPC4p3fwS2DbcQQnPMEcvfVeUIoOuFQFHeKDKB79HpL
hi9cDsRHVlEt2bHSvKCMNSOQzYMibbhJfTfsAOVZ71wPoZCY2oMtH9/1LkMrRehW
iYuRtI4wCOC9pee5Sx79s9zl2FT5N+D6eL4qHwbsOn2lo5wt7ManHnbIW/UuO66p
T3pJPTXIVcxokcKDuPraLnV8Kj9uqDkg+GrNfero0nYzghRygf+EAoZri0yhjNrN
z45/YtUJUYkIEnWODIdDfrPy6PG/wWp/XaGIFNwXPtjtZ1ryLdVuJO7mF7Xlx4Cq
T+AUdDNRy7QJqa1Pm+fMv/MhQSSDfZubFdu2LMnMwGBIR4eVCxMrZyTaTE1SMSxB
o+EIXWHl7qFNEtymIjK4qC7IjvMzS6Xn7cjdcNOovycyZUKeGwkgtkXO4Xduhhwn
kHMqnCMmsJgGoNt0/A4sTDdUHSkok+LMqcPG/lAxdsTu8b1FewqGy60DZjyvWVVZ
0PQxmBf47rBppPaC8CAzE5lgCFP7TiQ1OtFoirRxLv1P8Leh0BWFLVNJuQ2GYgO/
Jjxv7S7c8XDQsWY5Q8SQPz/dTgR7bopbDyL03DaIopOQml3HEU0471HWzqHO8Gqz
nq54JRHVox6Zjy18b/exP8fmJdB541bgRi8+t5r4IXfv4rOrwmtt6f4F9HVkXF35
oLz164rbQnRTmWu5zUJhJPIPaW8yfBmC1N1TR4fMHQANrK3Gnh1kvrGb/oV/38fe
EBEa0cQIXdo35lms8UAa/mEWY+/p+j/WMvKdU4WtZKaf6wKUu0z755aYEyuJlmdH
ela+iESWOu3hHJL/yHOpo/3UNbu7Al925Lja9Vp+9+1iPjht2iCTGb6ZR9/V2qgq
hvA08DDqVtL9psIG+gwW2jHu/6tCY4vyn7OFfvaVqzM+4ErY9PEXoqCKOWN+iqih
s5Isrqr28LVRHH+SYODKLwVLc20xTcPYqKXzUZiZUneCVcGhtTTr2B6pLVeXcQ2i
ikg0lYEfazqG5vbADozl8/mAzKHgA0fSVTNWx0qNvxryfODETY0xCpdpiKjTqgJz
115heS/wkchqqr6NYz9Snym/Qw7EwbO0tlsEleT8sV9j5UgHN5P5XsWehkRtafnm
AKYSTTvLhL8rIjIV3ri/z4Q+Z8QyVKyExeoesShRtLUh5Fg2qKRuo8ow/yWiXIzB
Rcq2Hzvj3DkxY2eDCXmZxovP9S2jptc4MGCm66hsLsf9vvCjZxorEF1JwGZl5WzY
qnWEYJGNoZwDa5heKM0N9fClhrdxDgcsKOUdqybZczY85/u+uY2O6KgXcnq3I5FR
6LBtmjn2d/nw0wdHUGSQOWZHK/BbJZIm19Cj0ge7IcEZelHgIxFATXT/76rswiJz
ZsBt02WxGaU/NhB2Fwp/PUhB1wSZNn3OO8ayrGGtq7KHezxgbZdoqn67KHWX8stn
RQCGl93+kPm86zAx8yhcbP0HxdloI1EAxLrKKuYKOF5kQJwACXFvN5MUNDmweP+Z
wVu6oMqU4/E6TXmCMI0RWdszAN20TB2/tjIvNFmknycrfHwr2qqrMzKArUa5C/Yd
/R1c+Y8N+ade+jkQEYX5a2nqXE6k0H9Z4mYMFfRzIQXcqLSj5GEDKT3oEGVumTTL
iupSp/xqaw5rDBpS8nTDpz9y5kNf4i0Ugmf5dSoccqUwI7UKJA7VhY5q2ij/Qy8I
iSbkodjJkCyCa4aTCCEJwjhcuNYJfztCeXhM41axwTHc6TUMVprvB8Xja/RFzzOw
Vn+iLxtIk3dJjc5seEfdOVuQC0l9bqEBjew8sEiByZhr3vq2mvWREUYO8eaKpa/n
YrnpOEvaflXdCEgbAFAI/xki67gR8Bq3a2cAJX+UFc9ILtsvNUiQdRBOGKqEYJUe
3Uu9G1X1k8FBZMogNhHRUkG84YUBy8ud2mA5jj5TEbd87JeXEahP7OFNdwaPDDGY
2XljQLQPgV+0hIPZ2mL9s+XItuChpnEbEDpahcO1slHJNxxlZV6QfzF3eVQneSKB
fFMJxF6OG8XZkuOBhwg35co0Rub1FzNMpnlRnaXjMgQ292BUPUdg0sMhngdvbfGR
e9cLOBIC/MVp+Jho8U3EDLNWkMRdI81KaDwMSbcc0AkmkhsoVJWJpPf3QUoQ7BYa
Vs7W1knoWZRdVjMs/iR4pKCF4FasotXkI+xj+bPhVvETqInyZqbyNLJG6Dw59ooN
6dQ3CXGH2FqAm33d5FkgVxajqojBLRCvqdeCgCpWVT1WQJ5IPXcLV7RWrEqEtDyt
zku1j5W+Ha1JYmLH01wXvZIA7NPt1CIjNUyUVS2dHE+YD50wyfgO/p/fNj84o8I9
+UXw8HDE7C/nbwf/0bbw1JWV6ZO13LqJSNeEIFIqgzpQuNOdmeocy8E1tdlc+ky3
o0ZJthomfe6YbP0OeGlldijO9KdWBytRQlbbEU1yZfh6rAcz+eeye8QZ50VB52JF
1hKEImtkx7+H6ghz1crlQxUbvQcCGka7sQ22kM41whk6m6cnGCcboxiaUob9KjWQ
BAnfdPoRpIxwhui+/GKFglWTGWsTKwnvhN1t5isNFvVnYyHq8q1aXBEgK1F422Mt
XIMSRqiQNoR1Pkc6rvsEdK3mcR443uUEYzsugVUeo+ZtzLlQElBa2VLA/L+dFkOS
nJsNqdXz8VrjxQDTrtDIQfffwFiWw8yZ39W4jCTZIOHe24yjOvXl/1E+tQQh+sGB
RM4tqCJ/3dCS+YDQXMD8QQF9joSEi0w4vO/A04A00c7zj/RrCgJcgwxpcGUe1t6P
0YeiWRWdRmI2UkGj1wKm9uyPZblQ/vcjaTKhKvuKvPcogiO/MaL1Z1AszTNi9Lzg
5/NM5DMfUnJxS04y8KYNmOUHFuWqrAjJQHkqD/ARAAZ6wTG16YyLnB5NCstEtqkE
T3zxpY2i8ocHiylumd7QCb9SVe1AATmBFbkbyh07s9bTSZuYUKzFWcRocDzTYneV
ehRBUIWejcfe6SMsxc339nh8t+ThcxtnCNnaHYz5qC1SjQlE6JlN7F+amO1/gHo+
/PGuxpPiE4qvYtOlFFa53H2TxCejZMcMs22Nd2RZ9tyOJuhUlEssq6sVmwzgmcRr
fmn3OMygBebOYLbhb6cRsak9DwC+FlGgTGc643Egu6K2yi/4YWe2vbyDQATn7NFm
B7QCzvBl8KAhFkgOT6e+AMbfSSbN8c0g8Z0U0KMFBMMx2aWQiQJ1iYN7V/AFY2NQ
+0KYurKGNdWOxYu0lUAya25lKxV4oiPfiN6JdmMaf/yeuDDdzOup3csBajFZgfV/
2cXiQOfkekUBONv4OmqLWNbhG1bahKfMw/TMiRLw0ZIzASzbuVwPvd4wLQ49sg+5
WapBryHvJbcv805Yg0v/F3d9Kc+wV+A6MDskPBBGxHc/4kzB8QVNPZ8zdL6gHmz+
EBuRPmGOOqyesxu9BXbuJtnRLjvpQsFM51TuZahOsmQLJKH7o0r5olI3MdSWR3Jw
XCx4hottx+/dLImQjvZxCN+f8xMSq7vmtb+gkvrPSXLFxjABMIuYFgjUP4cAh0cX
G0l3uKLZFNLKfT0ycBnBB7NBo9AB3S8cdUdcfNbvyUD6RPFnoZe1gCRV/mhm9ZFT
JVSA5S4mLtcPtBrj8foidVxPAZP9eHWrJ1bJxSyymgF6Pl7I9s2Uwn2JWH9+b6PU
bt8N2TAnrmdh2kBqw+vtZqn473qFO9u27UbbsULMiATlFd+LK7RTI9Xh7ITVIPip
NKELbMdfr044OFOhlfrp+njCdDYBeMOM8C1oWMVCZK988buW+E6SBzx6Y+5N5myi
MfcRR+OyB/JrREjsMPvJmzfDmW4zhGUuDaKHMwVx3WDip6TBg05wIHpuUisa2fbH
nIxCD+Q5bwyWqJSdy1dslx6kRbqGqxqF+x97K6D78V9k/scqVsbh5KRKVysHL+K3
G1i0hBmNBMeJk0bP+1Yz7CVStLHc9GbAbwaYcUes+f2XTTo452Kh5Lxm6fha1jdv
kqQUwHgv2qgEpwiSS/kwsKrxw41Df5HRRNIKUCkBnMwkPRyJuGWbYgn7HXO+MYtS
xYcc+A/OGBOnzowfMD+Dsv6AVCHJU6df3AdKwqfVkrDovl4mdUahgkFM5h2G/YHP
/EJqNxeha0CJFdOwfKE93obzb3xphELt0+LFaxFoSuZXmbL4YJDPQnzGF0OpNPR4
9Pm2BmpQ0+wg08c40WO6nchLrtpm1jWUa3nJDVltIk7KlOlTA3GhG/3IYClAXgBU
fZvHjbvGyK1tFpykUQPFJqWAse8e3VjGrjRAUNs9erREX3SH759jzZFd5tY4Ltl5
LX55qGL5LSurQFwt1RENsLcXfjNdUgo8gRtnI6oQt/RdGTp4tKxwZhndwz6UAaQF
Y08oNegE9CV5sW0Sj87J9COlu9evbSk4kcGBoWsarPkhY2QrskrycqhvHwzSvwWu
oaaLv36Nn/8ozqhjIRjLFQHtpjHuI5U0WSNQ0WvLer+fnq6r68dPqG+Zw73rDOmw
E/RTw+HQnC59wMrBNGRYAXr443bOQOA9Hp5kD8YQsLOaPOG7OY9ESHV9hHQ4FGXK
hZa5ksAqM7+varvKmf3WYGfHQiT2YlI3MWopfmNL1Za0pRVeHI9b8etwlsVLC9V8
yI5pROBO0WwWTfUdA/qYh1t5gDrSiOE2yVk/lacOtdo5aLSuoY+6R4Su8LMHEFxe
JccuSGHmHffKyLev1EJnMCb/3DOAVaqC+3kNVtWFYKSaZPTCmpvLE13j78dasl5F
bgi/atQNeA97DqMpAW6+1/RLpSLwSzpiwa9xKE41ySqBMLfwMVa/UV/gUeOKQfFg
QuwSQLwJVA9hicbcQQO82VLOmKYFrNXAQQCpNjF2dkN/PqF26LiOBOrcD1sMrTbP
DLweIjCFWDdSOULWEapakodP1OfEG0rfZmF3lKnuuO9v2/bt7x7iXfajYF7hVfqe
6IQZgrnIc1Wu05W8qJZGifnuDjshcG0woMXABWoxKC4Cm0cUlS/ndm15Xhp1+RPr
Zm3rRfiYTewkQmVMgwmvstfMSAY8Oi9W1uk8d0jJtsMJeo1esmsfXl0k1fGONE6z
RGHmNsOw5KaXnUjpTw6i0p3RS2XZhpml93avv/VGDj+yAq8s2UQth8O+2wvlFntO
TgWOZO9ExlvrbrZMXoAZaxAvrshHN7D+ffuOSHg/AO5Gpd90hYX3zGTWCkXEuWfg
Ug3+ZUvdkfurfNZVDwvGsRCYj9WuWPIqGsmyodQncojRWUSY7qrDBxhRS+wqD3CI
jEmjPdc7f2Csy4c4HcI0xO35J45DT2TvmxzplxZrhGRdO3Bi1p0mJQenF1lIAm4+
CydymouC2TipB10PqtY0Co4PpVpAfCnDlzLfhFkwCO4H2U6+D6I3hT3DsHR5eqtK
nOlb9tPjhETX7EanC2mHsdlJOuvGE39R1tMopLV/z5lBCbIqlI1Fw4abWL+JUooc
WCHNSNEsy7684Ca+Poh0atXDuhEv7oZn7iiM8/74vgNFOJOYylSc5UIDixS861Bf
miDKfdBihPk+u8TCM3iW6MT9gnXlO9fqFPA/M2oKg6dsTKyXz3LJQyOAIt7oXqqa
5mUq8OVXAZFMK4QBUPWdcZyq7KETlphjq74K6rO2TQfcWQZ1xp/P1zOgaI3qHTiK
hY2pa8BZ5l/dGLuP+XzaMqdODaDP9Tt7o78cVy0pArlVaezv0IWvdtG8APgWOWAh
6M4XO0p8V0ijTyTXvRIcMhRKD4LwXin3YnJlT9ON8dXzIb9zgSQu5uQ/WXVUWQeA
fnZdtT6PHeUicdelWuu2uHxLRZppeM8mtDHDyajRpmDXO1c57iIDVI9cQhu51b6c
R6XcAflSVo5udWdPgxYi1i9H5g0zVso+q8lAef8dUVekf0m6BA3WicKwiggs3pDw
0C2VGrPEdAP1XOVME/c4UWtQQ139Pc+Apktxgah1W6x6ZGO90q9N9+mWUPWJULiR
4JUB/6i22xI1LogqMspVgYPgpWc2Xach78aPXUKbgihX9RdB/fYqYitPl/vFF+8h
Hm0iDYuzXVc6pbmRE4UAyE2Dqz8y/frklcFg5s1UAJkfA+9ywJmHcGG8/veH5BS7
7ruj9aXwTF50hIO94lbiMnKccjpAKJEUMRxXW1Adk66AzMkHW43nJvVD8xzSEYxe
mPVh0HaMgXB+sziBMEsnWT0xDA3Y1IPxOGAo1HaV/iUSpxGDXH47EijyxL3O37vX
7gaWlORTWO88X0uyXkbj9YIKaThGpEt0G+n059qY9V7HayTE1LbS6Zmbys2Olm6M
rz+n1+CV43lPQbgN6OlsW9ovC1VavepR4gq8/mvctx10OfM5KzCPzzzmKYK+fzRV
ixf//zY4A0UesLIvjqpJbLY6RxERZ0jK50ZHtZdwgGTgAYv5Mwpiy1/y6soQWYRH
3FzIoax7rLz56ekxtEJ2UnTwdgLK4uC+8y2NJ/cNK1xufalubUfEtsU8MW3q4y04
M/xLzeCA4Pb8xVqKYCXjhISD5qGFCJd2zQd9rFov9GfwdlA5vyWrANMHJMoP6BCp
7OXZOAjuGe3XNj2wsYoWlPZBA2Fdr19znhSRUhB1lVIDuvuhqT4Eu+qAYf4cZDUw
AB7qc+ZFfJe69+zh7th86dTM1ZdJvR1yonIcZAu09YBV0lk1UyQtQKrEqCE6wI0y
nJLp+fy3Dfqpumd925t6z6ni+YuFqkwWgox4GFIdz2EHTEWj4jAzQ+222D5+dQrT
ME7bTuGsdoXt1BxPVZhy8l0aeu35i4It7qStcN0MixLsnv9VcW3sRY3Cyg0tp4+J
FLHk5IwHLhdcSY4U4r2Hd5/6vviPYVKSEOIT67QZFik/3ODhL7D/RrE2JOkMfAfb
CyV0kYl3w5aE08KPXfJc/iNguB3hu2ab6dJxC90L6OZc1CnQ0Gt8iB8bwAIEkerH
GODtZ7kDNMeyjYOIFG/kmGXowpRyuBMbIhRLGhivEivbJbD5OGAf1Qgx9B/CTaHE
IuiF1Gp1lwIVXtd0dnXdR5gUgi98BVHO6uCOfZryZ4FCqXCKIkPP3/5ZrNGq8GPz
hkdBtZYCbgzafTWsYbu6fmKlq4uDLifBWOmsp0qnOWAMVUj/oo4Nbj0BvsSdb+XP
6UTvrtNghOPWY+7Y08SG2gEyWhzld6nnydLUZOacUE1agdCnoTLUZtkymOgHciok
wE+/L+XRDX5h3BnFHyQfwuHXFbvm9q271jQa2RYfEBqIkVGzlPnAbZrUc33+f9TS
fPcBnWM6v1N6+T7Qz3rYdfcNZCrsYVZwz3AE1XnQAKIlQflbiH6IVxwMGECgzIKz
MFaV0Wl8e5jMQFqFdrb+3vh7WtVJWbvJgvWA9TMvf1bhvEMoT/lR0VEcME6d5LAo
lR8psNxjHFibTglJBe/g8t+08iUzqXHDxtABTIu6+l0uxY4YiA8LXvKbU0RBLigD
KDMMKDsXH/CB9vXN0M8z0uf3wPK10SSD+ybtidFa2Xhms88chawKCY50GIv6/jfr
q/qmcQNBfNM+kWnakCP4uwc3a5v9wAMWOvNxAfSfbq/VbF4YMP8jklZV8Q+dxMho
paFf/o/197/Wr4HNbLzhosi5ITg3ERfnJ+uJnwAKcQvgWIm/ghhOJgszR3JPXW+5
5goyPqhalMPV7OLK2UNkhTXKB8X4pq6DHfmJp3B2g5dwPTV4sxIEUTDatQrngTxg
6YUyP9PKWAPhnnHsyrJef+D8p60/6da6hapbU77xWWhu7Iy1jBLp8GqqMbjg8T0c
TtoiqporBx2DUf3Iz/dqqRX9Sng24jirVSF2meTnJFyeG2ppwHJRbQrO185dMYHM
HGBuIfJJKBZdu2v270RSPQiCzFgEeqDX/NvzTithX9hgZsw+eJcT1QxHrgQUKaMd
7maN9LPOBHgAZMqDTI1mby84oYWSeft59w/Sj4dYhHsFyS2XRrr9zq/dpm/HPdwY
n34G2ffCKeEyWcAEhhPb0npwa3y8uNwKtebZ+6kPqALWdDyqRcCrxY2LOwYlb1qV
TwquCpbmOgUs+8XrXpOApSXf3BQeTK6Z8y2FQv86YaZFhtsRLcVc81PcXYCD/2Z2
3YPPfIPsQLeTXJBFHmzCx3+TUa715cNrmJYsnmrpYyldmUlkqCa5DaanWWbV26Ei
9OCQr7/7uWsX3MDWz9v2iHpBakAqnnrqMfIc+wx6A73UqmZtEDKWc8ik/zFtTuhg
QNB4B9inJaEa/Ovqr88c0sp+cMi03AUn53RK6Ffv9lUgIeApRDEGrwcj12oBJzWD
7lHqmTAD+wNqGNXjWVne+irs2vkI5Jh49xpR4/1rWMA+eoE09LWoM4fLhNcYy+xe
zJgrFObC1NMO2MjCKhuCY3+4iH9d+7bIK+dzAjBqlC5Oh7tUz35+vzZewL/HT0dp
uuAm3oJ/srS1uuFEJRJcgHLnxmyla1uDtGKOW62xYZ7BPVh7EoU31ORm2n7vXIeR
d66D+8IW/3Gz32h82uvvyxwz6+sx3L4x9ln0CBx8WA5iIs/KmjVCoJa4ynwrgDsC
JzfQRcTrjWNYLvDynEYaA7DS05dGHhhBrdyFny8BHVTfgKGUUy6bZTwxfl/8XUxZ
EB4E0MSBiC8k5bIpxDppBZagJnTUJ7b1cpCQlj2yl7ludoRaJqufUQrxKNiakOf+
SXqWuRqgnMJJ/wsGNi6cpZZp+NPMAdZq4pAKPzuiqudmhXQpxVZaONeQAcg8WLnj
KsRO1UxcpgdbCiHpd6T1M+eF/Imr+q/TV3OwGkVTRz3xHxFHOCMBrMFaQcpYDxW8
t//9oomGmoXzIjo5kt4F0ImqsWf2kTzuDN6elcpPrV4GprNxwlhJI4nwB3kZcHxW
/YXBHuSeLCSmmdSYj8ZSUbv3KstdgOMKnZRlQgosD78f3UsxLLS8r1qAGIp/SSae
I/JGmUZFcxc4PL7M/l13Mob8A0pokOpM06EBPD+sfZrzA6THMjbCx+PlWy1GkvCH
txAQ521ONsJEIXet3jap2w6REzmN0m5Z4OBROk2po6vX9WpbFHtdeTSE+rKtISeq
TSgttWNJqSyGZeocvc5l7YEqZXF5U9P9dUm3Jolj6/4tXLHF+gaJqIftvCEzpZR+
qAbSsWgsLac8LuiIbRA65BQWuUCPnL8MSCxwgl/aCVqj/JEzReLBHWC7GgM9M5dz
Q6B9AC6GHwwcVIJMnZeWBNrwePvWyWl0dfNTKuHBvnj+H7nHWvTYOBuHKODItELV
5nB41JDT8N4rUhb0BD8U30wgcc8zoExnWQTHwR7Uv9PveeFuy3h/EPHioSOZSXU4
/aW9ewQDqjM3VBMHDvJZh7GKnfBQPvHbX8YokdZf9SyE2W48CwqKr9jQRryvAVSu
jfNBqC/mlz1t9w3LyAUX3vmQw512xIue8LqcCwwIgfnv6NPdlTYPC36aGPuMfVnF
Y7CsVQqfrQwpohk8z7Q0yaw1PtNJj8xsk8T7Z+lwtoaxrkSRPZgni/I5Je52Fw77
vh8zremnm0y4p9HE32DBmYi5u5h0MNBUhK/CjWQUQ1MTjLBL6JT3HN1Rb/CvM8DQ
a97hLChSi5gdxI9WBMsyYz/rKbIM5MXpahEqcPCVR9nIvXO/284WnjBQFPcBgv5Z
x561Ej0zFZyLP/JLdv7VPrDcCz/75ClbvQr4UndjCHYX4g+pASwrvL5RtTYzVvXO
vOYTslwW/MMizGO/aQm80Luh2Xa7hskhH7U30FhDSU/VNtH4003H+rMj0XhiPZ5F
aZT6JnQg/KJ8qNwvt6AxYDLkAj0l1Xi0AtYFysWdjCl40oZfLQnW4E5uzmFQu+yG
yeaoMlPg/BQl6/XI+M42/+K1yBmMPIAuNfQdirAKzgGGzisWJ7VCbEk888l/yMGw
jWf0b7AiiwqOnG6ysV6erp1Y2Y+eJqASByato60oR4LcShm/3jeFHPCJVKKF1zr9
g+gGOTgwICMOSahZu6BgbFWu1bvlEtMvANBZu85+9DSeyCpD8UggvPz//IIfUVvp
z3OVk0RuqwejfwqktSPH+ZQwUZ+RoK/b3rQUk15TuqSTeuEpM5MHadyScNcvOaet
fsAtRz2uWT37PfmYYujUo8iqz9oKlP1XZhKnJbtAIr4NiSpVXPX2reAHdtZlNCuK
z2pTf/T/wAbUmyKMF3DgvM1K6mYlHzdMmLW4Gt8NTrgKxY8YtQwc01MmHgx50s1x
k8l6G9kJrqR1orj2ZV7keXgAg713yjuUxx8njp+yIryensP4PTW/J3B+qjbpVIP5
rrNsFk/LyiYBprWNQKiArKM2OAyBvkpPaCznwteG0uaG91nny6l5IFkhPuDpKIIl
vQYGT1u10Eg48V+cJCNmzZAR7nrjlywvoLkHvLKHFuF/tSetna2Z+Xln/wXjgBFp
LI0FnF/x7ZjCxiZhjbvyilqZZ8nxgwGIySUl3Sp0FSp4P7F/I7mtfWOa3D+7g0+6
N9wBfsIKFNyUyedKd3hSiNumfa7H9OKexgFRUeNwObocxvuCAM43DpKBItgXIs7I
bVe2m0vTttO8lS/KEgCYlwhsq/AG41qw4RMbXCK4zzjFqEYUiDdQAjhxj1XAxrQQ
DczHwgdSQz7aUDuN/4ZYjp0qP3t/9Sxu1umCqGIp3BLdIctHuHudnMktaKLmAO54
iHHysaxF7wOPmANnMR1Kw1N3QXLBXS+gsegR81toCZEq6uQOjP4ANgsIdb833Log
0xja3a0Qkx23omFz8jBiaVwlPfyGy+7ExQ5N9ae3bCAj04E1wcE8dDsXtcBi/Ia1
YQsCCVEd3WjLiUMtx4jvU6X7phRdz2fx0IrRDFpn5NU348VB1b4DrLexIEB73fEn
FaEDxUNjv1kVs07fqtMwvsJU+vTJ4iRyWZd+MxzLCVqYz5XnIYxyRXTM7OV3bWr8
JmFKkw2EUC0ljiir0evanK9uzgMbCAuTilxivWKPHz/oCYvM2vFE3lsM5UH3cc4v
HFlbMRpyr/3BspQG41eEm+OdTN+6ncA4gRNIfqliggAqBtfKbruU3EGu9R0UZAPa
r3Xyty4IL5mcN+APst+5GOPm8VBxpl5D9/xoAdgNrOk3yTUTWDZeq7EtZ0CPiz7k
wnAQGWTkx0C1xLeaQTpuEfxun2WlTIacNHOnPnXjyXcEYVoR0OfUPfBW0oh60sOs
gQNCQO7NwAFnx9UhoiT/Z5CSNthxgy2+ri5IHDfCXieeCZoumK/I0QXhlBCuCcGK
FtzgjNaK9UwNaxCxjlsOwBvl8ilbZu8JScQ+ov8EWmbcgSM0xH6bsb/sk6rm8ZpF
AyLj7mFfuDqYUI/Gr0fbvTTp9jLwFM8xb/DYi8eugNcA1EFeY79rCBzXC85O7To0
vJx0aCUodE3/olngT6NApAv1lgzraL8zbxD6kOP5vEb56yOm+LkfOWb0yHDHN7rO
IMlW5lBDIzQSmIG/2IXaMDinflCD4a/KkhFob+TPSWXCEmx9qCxb9prYF8g4l98x
lAoO/+hHd3XZ8yAGiRtZoqv1Q7eU7N8VNxeBCB8k0tb1ImWp2dfxAz70u2fyaYI3
o+6f6koyrwNkoSpQ+stPfZATDkqSbOJsLx/HgbUOyd56tT6UJIWYqEaS41xIfkTc
CjwZ0HiFntTiirQBqyLyF/u/1r5QGV1axguoO967tkc0Oa4njDSiX4wFCLgwcXd4
Wfktk4go4y1nASnA2wb/K8ZoZ9yCmHXnlzCCbaYTd1U3egpHhANpCqueoFlbraN6
QJQNiHJlCUkKrQ6rsibAvHYQNmW0s0vShv0+0J+fIHKxTgANPkBdrHotWGDEP1io
db1GSHSzQc7yt/JL91lOGBSsfld037OqJzrWYtwMb/HJ6d8WPDDDZQQSbkB4ii/2
o+blupkcFBnlLr4EQlM+rES0hI7g87TbNirsQuN7d9xLLFPGw3jIUlj35XjnTTlq
KcA+vWpRc55qCMlE4K2bjSACtr5omqkwPhAayFkH63k1r0RKsJBK1jjACXTAY4uq
dY66wti47q6XcojunXwbJRfXxlme3x3MBRmOGnpMeK0PyIrT6Bu/fF/tPL4WCGEZ
I3n93WwtWoyTthOG+hbrHhkOnmjKi6nFDQQcjZPVwF6TFLWLSQ2QWWuN+IM+5l0/
7O4LPl+qe1zVOl5qBaL2JYYNrR3/wTCSjcHwKb37okJIj/aDk1GfLCU7h0GVI5zH
brOWcNrTa3QWnUYOJ9/WZ4JntMeNz8KsLSRt++gq7+LRf3E6GL7cpvdXAgEieZIZ
w9JT4f2Narn0boQeL/d9nMjbJgS6n4CkqLNnJrQpfz4/hZeGcoOaqZZzMbITJxT9
vtRhWj8L9ZrHUKKOEimKL2RAEm1FCZetuQ6c9fkhRgI7FM7ZMjIsyAndSrX/AqU8
/jicnvQHXJ+uFJPUkPVpSQOAN5RSPpxSAyjw5Ykzf6D9KjkRRj2HvoOzbM5zCVMy
7SeZO6sREeCOgvPbgFTzSnPjtMkIxWwJfNvoOmIjHSDkj954de07LfeQyjhmv95O
rqQl6QzeypKAE2mtU8sUWFnc//nfc3PZs+VeIszJW2zM3yh80As8feU70h8t2bXD
qnGBoZWuDPTzANoyaF3Hm22N+9HDoAZvmjxsV+CIGdsYpSRNOHeWhHXRC0CFT7ok
uyAus3paNWFgUcYVqYUEhJn6kpchDy3eJ+aHwG6GIUbpjM2L+X8T7jejzX11uDy+
1zQ1PIazDHE56erpoikXTMGPX0LtNyvmJA6bDWujuE/RteJwx3eh0cYvzKQtHoP4
d8AAxTa+dRoAqH5bOeCumjF9RY/lrKGSfs/lgL0+MRbObvUV1Z9BAuGZUJvv07h5
IQnm7bI6iVH2Akubj6GQy3yQnV5TYNJTFCLZ2g5EFhUeRZQt5vH5xReedd289e/e
qZPBeLsfPdxIbKPzMXJwQhTAsCn4jARvCD+P+GFoZKC9RMNBESaspEvKEbFM2ZPK
GGxiRnNshyOMqDcu9KBLw7XXa3s3GFWbggKrQiSJ337SwQKRimdqad+HYSDrP34s
+hW1w8Mb7ahUGfb6CYREqSldfhxS+vY8xXO3X2c/3kgwjeYFq24EF8QaKanWhNQn
oBCrJIkEpivCUQ1PZeNjKEAdSDRDHND08eTaldJabfNgYD2TI2vwwcdHlsabknOq
Z8cCG9QE40fIUe9jPz19jBcGKiVqRNMnwMTAQzIcN9szab8nXfYldU5qkXLmu3hU
8FQjrBXoE4qiPON9z9n+xBVb53uDmHyHv9YdyLQPPJ1V/nKQ6FBYoc+fGEEt+EZo
8E2+i3z0V1CtsCSZfv18iPWx+bk6trx+AOV7Emx7z8z5ayapeCVLkXwWN5H6DzF8
nHox0G/+RTzW66zeJeBs7JuhVfAKuzCxkoM78TlejeeDBvSZGNHB/X1mUHe6Mbym
itGxhIPHqdUcEWI8cmd+Ft6OvuBt9eEXHoGUYmjOIkvg0EJJS+/aBeez4Bdph+Jq
CJaiyvPvsIKG+oSXNbnXEF46pOM0z/1UanGFoKxpc1whQmTVK6Q5RjZ3BIBwNX69
hOjW4mn1qnOnw8OYce0F4Oht2xwIEqidBDv0jPhT68npuSuCI3cKQ/9DtH1pZJCy
49qBMAgjYzQUyasrf0MB1y08bYFODxVHxbIfD/F9X9BtTX+4bZbu/d61Bv/HD4tF
CP0XTUi8RTfkpjd0OCnCDGheQ4F30nxWitQDNSyeSIouD5lEu2t/MT6fx2cTqfWm
S5E+F1sVKm74TBnkDxoM0Xakgp10u7IU0vxpvawDjg7B8EqthpfDLCd8Fksi8Z2y
VuJwPirgx8KrdSAofxRzCZn4mB3wrbHCcETbpyMC6L8zP/6IEpNLlpik04KcS/Tq
P2dWa1sLnkAIntpf++kR65VEtVR5w2D8P0lPSKftyR8swAod+hBxgeAX2nsEK3N7
0gdPG8Ucj9N7mLNIZNJYY+/oMB12GJOSa3Wu4Zw6RbLQ+Otr1jpEKb1fC17YSule
oH0yXl7iWfTt6NZ7AAcvdR+ikMTTtPEqgLxvQ3IsGgxMivySqKP57jBRsgjeSpNc
pzmpq0zA288ncKVylVR6bdlIiUqewavIylhqeenFJklPDLFrWOAO4Lcswi0k4Wz6
/8nuq0uVQOouiIdcjZhVTlhdQ/oKQTgs0nVDLZvzugY3RB1VEKiTSqVulNQVlQdL
ddTSm/FbI/80lKA/weuSukiXXvO2+PWZszUb5KdqvRlmNnRRXC34zRdcXxGxpDJp
IRi0+B2yQL+OdJKsQC3XmnmtKKfsta7kIlO6LJNZyPfQQVbj5oWaAuVo6XbVjikN
2uoRaqcxrubqQjWSIHaMTbwsASRNfUQZ02xjxoLe4VwVA0EK50hdCZJAuKOAbDbb
HKymfx2osgZtoXiEX7JGjlSq9rAFLcAzLmv1wXclWGff7b4aMM67Cba8O55moCHC
I0iVCSK9HKHrJ+M5bm1ZPQE82jy8QmowVdz6STDr2fEudhKQPKUUqZfD1m1Y+Nrb
DqoKh48ZM1aLWPUfkVgjwtf3mCaMFHZuX2IE7LMPk6n197RiC3JHoILpMSAlSUAV
sdac0diS9kaRqxaiMAJLP2lUksoBYiRLNrcn6BrlZlb0XqTUZjR4y5awLC8fJpYC
+JMMuyacDY/a7GPcltoR1YS155FIs5GkqQ4aFpJJ3+aMVvEzG7UG3lSW/im/XvRc
Y0rdFFmzZV33AoW8AFc7gKsSw925VHaT7TO1WQkNS5BWEJkfvf/lU5U3F68kQhXw
XizT73IUCPfavdohHt2FpLexfASNYpYUeaZMWxKXHhxzyILJ94S7cCWCvPzaQ8h9
HBxnui2al5KG42t+dTjDPQPO00Q0SCCCxIYTXgTgXUZm7BoJzrNkzdFChflTVzgO
FvxmkyP1l7atdeSDQk9jLQwS+GaAA+SjRZ1zlf8IZm4mr9+8vezzVfKNUmUt9UR7
lE9fTFyXBhcmEzo/S9fplggDDhTATbgfKB3+4cHw1egSRtEixO11zxD+FJCwe/jQ
yTo1UkADRTTFx3Z9yb63cU1cDwYqtmp4xCPYiyhLyPNH1ke+wb+mcj/wqRgUS36Z
dsmP4DfENWXb7fmYVXKWs0HrgRvbpGTF3Ma7lXkBjpWaWp2EgxtD4AXkRWbL3Giq
AsjRb+VvVPd8undtQWaDUZNyfLS4PKl6WsTbwCF2SFICCxyU5X3E0EJ7cE01GOpi
DYWAFLvmoI8Q967bGKfTLsx4h66qWzUmKZUg9OmUfV9tWqVZJPuns7UZ2CDoXqCK
rDFmMs/j/qy/DbtKzgN4bVmbnn6WH0ZNZNIk/UNr+eZ/6skyYkd3/wQPkhI1bN3Y
POTv4rC2Jwj1Ey0U0Ggeh1wiIlvSbF7mJxK0H/E+hhA0XWwGJbk8aiPdsff+S4O2
H/Pvj/SrQfy210HnNaF5twEEF2JJSk8uvhKgx5KOv8wx2LBm8/2rHMduJKlyelDE
Jo8KSnkJE89NhIKPm8qXj1keR8YSwHXmGFuYbIKg1dChuRJzm9gLTHD7PtihajWC
p4aHnr3e3qPDtgzw6qKIr7sI47Noz6T3myKEqoxXhNvyfUQ4a0cIX1fwlMeYDhfX
+kFNagzJefa8r3AhfQvpOuvKFzn3PKkGiV3qk+0TtfMcAYJgYLyIHcZGKazgsslV
RdfitdL2SR7siN41U40IiNLaHFpAZLhHJbTWCAt0VcBxHj0PWb/1U2MnpRZC8xQv
Gg39SzLVD1eaEIMdxhNZZ9sbd0NLonW+Kz9yLeuOAtcv+MiW7FZjVrsf3S7j8Wr2
ehAXMyMOHT+7Qmn4/Awp+DAPbD8KDjCIQn5EJV1bXSOHBXkkWz9mfbpmzK5KSuhF
DLWA2Rv49Zw0N756U54IYkFG1TAqbLvCAt5w/SQhUb6xTYAZmYygZl1UHILD+Pi8
zh/bg678XjYQzun1y/QJf445WQxBLG1YuJ2Bj0qpYjuWVf2XWwZJ8XIPt3mk6yJI
jhY4oaFtFE6zE2ZPNvy3ccdAdltnep50r4mdKFZZKOoDpv4hGb4bu86ob+fHLAb2
z+28S/8ca5psF3BvxszKsqC5m8L9AN7VbqB1/szcCPcXmMHv3QzaCSjxS4iDQOj0
d85WDFSPgeQTGARPCxv5QMJpU6H0W7GUulVqu6c0FOVAVuF6aW6eHOi39ef7xLGL
oH5v8Nxf/h4wXZbKBtBCVR17iLIFbSB7gJBCdbQ3+9DwJhsyN+WLnHULp3oddyeS
zHyre+nOUAiSzLpueIMnbeN9AYcr2SsXddbqZn+F7VH3w99x2T5U5Ze7gFslowt0
y/I1losXUD0R8l2JgQR+7rmKBF5X4UW3MAPt2QZ7ovH3dw3DtSc5/ZbUiV6nFe7H
eW7RyzAtmB0r9sGKSjn3o6DLns39V4rQ8BcSXzjaezycjubhgCTeMJFDkyOK3BXv
A32EDKOXpSX6DB19ZoJj5hiMlim4fWoFmb2kq0oscX8dqtAaaNMi5YSEhm3WaD2l
/N92dp43s+M47l9wXOvlvdBwTwmyRAU+nZAs4vwoyaQAPFab5CTERd45CwSUxDWA
Ax+7lERK8MtvTYAnUlUiYJw12Z62VQ+7tuYpYLNk8r0A6SbT1tfvSsgCOWa6rnvH
F+9Ft3BRE1XVe3lvpG14S8kgG13Ymk5SRonaeVeQfIyQJJ6n5PrxeThJcRTwbsC7
mOBoaJ0THe8JDMx9CisL6gzKFznaHvrpta0q5gqEHavnRMEnFFvCQ0uLp7llVAoX
fhnkwUSL6fvciRVpkwNBbqdUIn9vGdbP3BmF8D7MjE5j9cP5lGi+wK+j5PWXhCTl
Tm2mNxmcRfZPM27t3Ul1bQtxLEeGaYDAgTsjff2gz9e6MtK9mVbAGKD/IlivGFaJ
6N0GJPxQS0gTPfuH6+GfA0TY7B/Lumv6KHthTSkMp696W2Orzi79o7oGY5okwe0R
uo2zMinsIvts5P05th9iREDpt86nipzR/7hCiyKlAerJBju+O1SjHDW4EJ2Tp+O2
dhAEQsTvvqIdBn0RPw6NpCpZVqdmsw/lC/W/8Kgi7sATBDDayeu7ZgX5YVKSg1p4
YSJUPogtnzbUbN77EdyXTxxTc3S0DmWF0nRE09wPqwuOMkmlwmkone1tSgVy6Eqr
Ivb7cr6UzOe/KzHQhTxTLR8fkr2qI5z7ZcMedIUfJlJZmb8WfHG0ClaWOgdI7nqI
DLqniQkaZyr4C5g0G6jrtxOiRXr3abYwsDRHcgKxz42Ig0DR/UJnDPE/3zdChMdn
cXt0NnNBIQCJmUAIZKv3VHPlPmchfCjxF3Jn3P+uBbUot68JEI2X+3PJOLCoFw5t
RIo/RnacDsOwisNZF94g15gQPL1GPLWO/4YLmFwvWUbQxveQ3ZCqcxm+kYfGVstn
DQ0uQ6ZifjI1AZfeN/ZZ6y5nfiHahSm1WET8udGg5C10HkhXtqZDHpDVEdPToRnk
ulqu7f/UyaIQu6TxdPkZX7AOCJCmiltzpGIrGTBkmO6Pw2Ud2oOtQGRtsNkOT3AW
396ZX/rCd8vIUzQ3xASgENyyhdoubkSqPNyawTerDgJRTBbIYgQaK6FyMYqAymYM
FFDe2l/pQ2V3QrdRCsg095C6GyUMke7HPbI4YJXeWruv7SkYEzXeAKdxHFUGwUjh
5XLiCn3LF6N/eEHBDV0suIxQAav0TTC+O6FRTSpXyFg439R6pJUdfPL5d502pUth
GdPi7WP8LCO3FZ/80ZFyaKMF0i9lamTjCwLwnAyQeU4yI8BGWBHmboj8GdasNw1c
CsYWJyGTY6pRiA8XiYP3of4ARB1tZAt78eEo+H+An4dpRrnSqKNkxlmvkDjIRB6w
hDCbjagSjvrMW9+tCNr7XCXUib6LX3lA5zV2rbDf6MvoOpc7GBO8AB3DBVPZpvC/
EXk5XgsXO2jLnR4rCklA6akpGB6Pp2tWCJWBn50LbvcYuzYjxBiGHBXtGmX/Yk9A
u3eiYKf2zBzFcocdmwDukvAdaegCieXFlPo+Q7Vm0NutzcfVeQJO+eCiXOAh4Pz6
Mdwjv1TGs2sC0asROcQhv2W2tXA6EtVDRvFXRDbFc1j5WBDvrBdv+681zIdAB8rA
gJccQ6XCxqIqLj7QtLn8EDLuikDoDAzuxBemH7VBtX05zD8muQ1Fj8WpLvZ+4BoG
Y7BuuovDR2HMLJeeOWtGeeKx1oJnzhbJnJRcBjSgsWRv1/xnOKX7MZlbrcMSPi0+
iS2ul6XZbSVufZy87eOSdqlP6Ggu9pUIVcLYjx1tuqrX5In2yTG/K4d4g91S6lxP
1sAXzinOZqrvYlQbL4u/tYel8gAB8UO9wbR4J54lKAe8/izIfB2w51T6ChOk7t+w
/2e5rcEEPLjg5xyX3ZT9oyLN8i1Uita6tGvi2RHR7KdB7ebLf+LEsMxa6N41q106
LGxe/1kZtUuOT5v8M989oEybGvLcRp3fLJCZMNzsXTZoflK7n8RW+cWuCUOsP7qF
0mwHYR4O/vY+2tkFQ8zDB8cQ2Ourvjt6MQKHNytlYLZGqEpvbA3lWmtvVK1qlyIb
AsWgc/I4ffYPy9Whg/eJKyN8S6aWsKDZwfZF8B0w62o6ea/VxORmuguj3aPyRVj2
4kyxaSBXD1Iye8YiGFcBXiEfDLzympd1TiDYSD7HYLu16Bv93h5A8DhARid2lhqG
PVNoN/OnoB07o+MjCPuaKsWu4ms8TvP8eEZKUyBG+BMpmXZxS9pfZVe+Hx/elf0P
HaYWpSSoo6G5+fT3YFBSSVUU6hycpdiddEC1PV1qEa0etq7RWZdWmDqLYNqQr3H8
HGP5RkFS1n8Z5xEfZ19WkH4jYrSqxoH96jbNkgcibTyPOXuQHByQdj3aZPciMDU/
eAInLtpQT/DZHjLXlPuNThE0fyO8BSrT4cE4m3LSIBLAqzpn+pLVra+epQKx+nHQ
roLw/rUqqlmfK8Xy9XeTs38jm9Nh027TgpKdPca/i9zcwQIDRT2r2soLUhHNgx84
5e/brEYnHe89lqU7nWrxhxqRzRsgtYxrnej8rVorlu2CRDG9Oiek69KhsHKVt5Za
4w2OPfD4yY3HQt+ZZXMGN3tSUl8273zQZFX4d14io8WNTBvmxiMUtUmrMjAPSyYx
uBvthUEUEDhUk+VvgOA+rL0mz/D86r6sHUZlUNfY16FS72nd02dlXNw1Ljb6sKtO
z91qAb1JQG2k6InBY1jjuvD6xwrDmua7qzCihk3dVb2JDR//BdUvZFQ3eBK5NSC9
vnu5iwTb3XmRiahvxiU0RA0Q5KZMU9EaQGkoMiTvjtMpAkVq6gS3UVSDxLdy29De
kYVZct7lKsoyxTYN1rLQFSmDY+0QULrn+L3n4eCDPRC3IJIDIoSexfDZybo3bTw4
PbJpBuhBjSQ/SoaCA1Du8w0Jh23lq4e4o0/0tLLbZoAvvX8VQiSc4egn6hFrKdZp
cTrFEj7i2nad0PLGsRwtWxkYVDts9nWPE7ITe6SILoFqrlkKXSbxGsrLQEWabkHB
RcHsizpC068oyBuKB2X2PN0/i5lJAfEjBAeS3DWkD4aEx35LM5P0xCM+8n7OZfHV
M+wJDo9lXugkD5t8dgWyFTiuMBwn6NEfA9FUZR/yOq2AkjH1j4T1y7Yg4NYhWWmi
cLVB+YQaIEXc9hgeZusgK6XrAPV8BVnIWdJ1aYB/616DSsK4KamG6tNAGO7m+h13
Uv26as7sy6iVKdgYylrPrePEjCRFwc8gW2FBMASclzCggdNb1Qv2yx0Uji6iJsMu
doAlBTsy44oW8V6QRBwCRVX180ZkoGejSVVAzvzwVEQVwu/NxxqSKJ8ze341GxEZ
Pba3IsXy1+uCD4/nc1y3C1d+2xKLTEpxOo/KP4P3nJOHyMT28UhiRS18NCUPYJ/o
bjC8qh9z4o5rYoWDrGrMCFseOjEAK8OY6lUGj+SkHwtMax1zEQaIqYKRSfrD6gM2
m9kemmY1Welt8Pv2EuMRICWfb6ckng+ay73sMQLzgivrNah3Bw8MqvmvAV9I8Su1
en5DAg2tg4hUnVTNBsxtLHX78sWGFy12T9QobDm1vNujOt6T9xwgr3DceqTkEwmB
Q+PSF5T+YWgOPdToX3q44gNrhA9P4JfnqW8P+Lth8XnM1nBsue1FAQMo1g6DFmZH
Zme6stzFdxBgcPXGUBgWReI+fGvOjAVospCY8mRlkYw0STPaTGp5edbcHIBHTjQe
DCVmT0NQ+yGmgA9Hfinol9pDbAJlg39OwYQDuktsaE7hUgvtKT2ZMJd03A9AufOr
UNLBo2j/fW5pYBxwQonK71nfyVpGwSy80wHB+yoztz+EZUvx/tpK7GUfOxT6XROC
AEBAYQe64ELkTwnvbFKqYkUTgCBhvP/tOVSymkXCH7iL4KHzCzyzQMecMr1YMfGr
ku4XmDsjzplHu9qeRJ4yZUjHGEmgcsqfsx1BFP0093agLeaXN5EWKdn301ROV2HT
m6OtC3hF79xOe06l9FmYZbQMYhzmOMUTpAeFwap3Dku+j80Uv0EHwDVFRfWtdNAe
RvRmAVxe3ZaUndxlX+Ofx6XNSpjciYdbaYtaQeDNcw6hkZrjxuW/BnxtMplJCQaa
cIk1Sw6fz30larIrKCksHfCi1fl8duLP3dlPBrYrfPAAiwcyY5PcQBV6YdCHsopU
VbB2C3r0AxyEDVRrXl0ymSwo3INTqRjk/sIiJ+TIe5fpqkSezljlyAt0Oo9tKw6I
sFyc5EOGU+i25w29TZJKtEzLVseN5rqGqiP9bBborkl0goR2lRH1ylz/TNEtK7Tv
avXFYcFbq3Evk9+pF7qWtkajaFd3VfiStepKOELRgXgus3LK4upbEWkGB1gkgL6V
dOM2DXO9umDdmH5+9Kc18gNsolWJS0CqO+/8tlewALMb49FADTzMoqqpEFbYquD1
k5XclrymoKx4kQEEnHpWlKT0j5eVgOgMiORgTZi1vus2m7PP2MhrRx8/24Z2xX2C
iagLeDO49yXD6N+PqlQ4geuvpkYTPTVQid7DZQMx98I6p8C4+Peoa1vg8L49qzeu
Kkjf/lknAqpzXuz90V1rCujICoAxpq5KbJQShMcbE5sB7CQc3pXWRwLrMoghNCa+
ZAQZLKPhu8ZGd64dTrQOB4yiPRLgsaIpH1TVujjUyFjC6frXkYh46VLoqnHpD5U0
s1iyEjU/8YJLDzZ1JsiyiZlHNXMm02rYhpipfBknX96Ys3nOHqL65qf10del4iRa
DZv5pq+8UDMuy0MhV2jtG3BCNWavBALEIIjuR3fqFX7xaC3uKrgT9oirl5UlIt5Y
/w1Y3COgmS2/r+Kka8/We54uoOoAYcgNwdYbGseNGYpJEJz1H5YEH9im4eiq2tcw
5NR9ofdlWNu/CsTylqWQrSFjQ7X2+VgHLWx82lZZtvu5T/hI4antdMuYB/TFYDBO
eyq8+21y/gemJr9a8NhYOdaDp1Tl2LqhlancJE5qkzWtuuuH6or9uZb2DQm5WENP
p4Fiv91/4tJcm34mOX0ChxpfMNenvTo8wEzETQGsb2Itv7pYl6aPtOIYTFKPAYWH
C6m+JGqEbhuHlIvxUVQm44CyuMt6ZXcFgoyecMBL/8pHAgsBXd2iHt84sZaKx98N
pKGQxpNOZva2THExQpK4/TjFFUFAV5LtcUxNe7aJs/XRkQAxDJMZFuoORLklWse2
9s7i0n6v5AsHKQahnHu+530TySujClm1ivLBZER4K0YT+1wN5pf/hdrBJVRTE1Bk
YLaFQ3zYjcDmfHt/yrYrGPPLdBL6p5sYVGt8zVJpW1bTXz4mUlHqvjJpvax8aVrR
zYK8D8u4Yctg6zT9pXFE3Gz4jos+zQw6L9vtXl61NaW09Y9z1wHRjKsYvourJcH3
WHfboocN5lVVqXWRYWP87J8x4b1Co5F6m54403qrWUdE0dVgYElBoeknM7JJpcdF
03nI8UN8a/OZfEzhOIJDvzFdVBNe6m0r+2+fnmreSlLc4v3OyBiP6cWW7HIPpwUj
1gvZNPBjK9AGUqhbFgPdcy/M2qDBTRjW9Lp9zVvebfzpjHCQAQZVhyEY5Oe0LPnB
BCdA2orjhPuSwkF3LxYJIrYrM6sk/MWIbTDdpyYAYBRBKjZxivGyQpTs9dKhkl1P
ASW22jhK7wQ15F6BF/zPDx8hfqHWHcOFHnGpdTANJ4MGP5hmeNgnYimWyVbCXf4C
pV6BMlEmHT8SXdiHcVMbFXqfPuiqVxQZQqzP/+CXOhaCkTym2cjOtg5Uhdt5kdSK
oPpS2CqkpzKTJMHU27zs9PjPFBFhI6EgagvzQknqyamgvzr6OFtAGxs7WrkmIuL7
wp2isJ15FMsTj7Ao99KZy84niLx4d13saLzuZX9JCbrSs0tXU8WnylSUtNgS2nVg
m3czrbWRiXIzRfWBp3ZI7dcuo1zw8ubt840cwbkHQTH7MYuzltln39+Z9H44EaT9
HyqJwsrmTD94KJoQKcrV6ElQfqMFnEZM3NrjDVX0MudQeLZ56mgBE9JR+kE4FIxd
gEXAaPBfu0Zw1kVuVwAU6PtMqsCoAIdDmMftm7CaDaiPbjt/cTlroPEB7scnj5u+
aMOjvEi486+lBcoL8Uaq5R/DihmYORDhWl0QmTWfwzSeEC1CnZ5/Cm5obglKRuv8
iIC3iOKYEhlVWsQzkX6PTVTAbMUeTQoBBWg+BXsyfY18RQ11aKg13pOBd5se22dD
Kve0fjgRosJ7/S6+GQN1Aj6E7TTLJ0X2QK7KcMcvAJdWEkwSVrr5WxUHH46N2UqJ
DG1M/WcYU53s3uJeIitatKdBDsy4z4yeoQMPNVqTej2VWkW9SbEkvpfoxb1p1VTC
D/npYl0/k0E8u/N9v9p9fepMrNo9xCCaXQfCBsfGrPwSKSvAFi/1S9fJH6Sr+TL2
YaaLAOioIrV9dxL/7H27Mh5FwNIZvWaj1mMJ0KR7aFkYZpjOpLyfpJDu73pR+0cM
71wXrf1HBVgCBXFoan/eLr7i3q3CtM6W0y2d4EuDhU7A8AVEV5ufiiax3HY3Qhof
LQEyYu1dsTfCt7oTc5QMUzzyT3kXDH7jOvhkRIKEGlf+InN/3AOjVtztsdbKQ6/S
xZ1pv6QmrSsAAHjCelYVxIuvt5G7vwgu3E+iHOBjJmGmCMnWzyiFkUXqa2c72/iA
2ZtC7tFvbCldhZQ3QJmWbBZpt7SnkAKJTFCLdc6tZR5HatMv7Y4LL+DPZqbZ6NyC
lVelFeOXseL9n1u40+2Bh1vOYWeAvDSdGMOidDx7LiqMw1uMuhuR6JoQ7a9T0k9j
WdgOq/MNTQ4YtmgIFew+BEyNiHTR252xUzWq8PKJW/i+DyVPMz2qbqxsrtVmcgyE
CZwLBGmZRUHXfUgDpvHZGbhO+faCOdlu7G0JwL9Y/oM6+ujSRrJcRjAC8f7jrnXw
jt6zHGvvGoiAe0egFV/Gk15ifsBhjj6ySFhqqVaC2Ks1jEX7TveK5Fwuu5Jn5j9v
AiICJTgB9GGLEgbbwjK/mbFmiKH18YvU/JfJx0avuJZOSqPGDe3dWnQO6s9eWJTA
hfZee1H9mAswZ4C25cEHb5qqWXg9f0xpQH0lNt9oaKV64/DmBkJq+eXgUmqOfw1Q
l7BIoCkXDIsaVuRxbSI9fXfsDFUY+vbbVRt8paL45FvO14oC4WfgrgU8zoP28/bA
xS5NoLPkLqUh7Cl+VkiGhrf/ctbTMf9viuC/0Rjn2ELxAJeJjWcpmGjbSAAvH0Y1
bzmQn612DOuC2oamYyqmaEVWMIsTqAA3qKc848hx1P3EYKTdHsRAkq+NOomyuE99
Baj70UfS5jp9WZEXr1CGKmPMTV88nPVy2vhfvnmNi0S+509j3ynN7fLCO/6lh8uT
NfUp/8Avpo6+UHgT8jqxapOxG2frOIlDPrYYnd5NI2NCyx6DNA/WCgNGfSIjl4zD
ddClDg2DbfsoaIldMwLsroFRavtgMA3YzAGrUiIIjNwAy0zVZsNiDAj86kkFouAp
T3U6r1MlBpHKx34aY+AO5Ecs1AwatSz+kl60kfx3V4z4i2sxs6Q8zuyTtZsoaOw0
fKHBfheYZ95J6zknzSUKd7iJ1iTW5KERVMMEbTJtEZECDiLNse7CXhxd4a6J4yUb
ObbwJbpNfIksuQNXehJn6nS1jEvNAiXyD09O8nAKu5bw1g3EGmBbiEOUCTRqYjpl
8ZI2EO4/YuFyTqWbyTEPMRBA4/tG5/t0xBGYSnFPPSMEH5VLK/7aCs7Hi9Dq3Mjz
Fw+Jl1DwLT6dddU9oceiUziKd1C97L2ZSpBNFolbTwEdEWvvljK94yaKaxoSuCgV
qv9t1JD0zcT1Pm54IA9cv5QYQdmvuXY81BTI4M5NDIcqvvUAZjfdVpTapUVpxE1I
yYJXiH/Wd/X94xgoIAitELRxqPZKjxlp2T2Tdvc0H1/GQcIFCs7LGPSxdw/niRrO
xQLm5v0voMZ0la93EOfA39MPCGnvsrfmQmjocl8aKSLuuUfC9nvqJuW9QzlGLFnq
7SoWrqCO/3rQkuYKWXK0VfZKcR64x2Ac1x4iq5efzja4+Y75/xM3PKoftC8o4oj/
Ofnuy7bxtHKBfl2TOcEYcIFPFDBDYkSDNeAt8S9jrYJV0ld8BuDUeOX7lQ7n9RYZ
jF+m2d/KeYV/w2X82RvgctGos2TzGCUQWpSHcx4J3aV7QS6t0fBu6ewPCrA5hWks
VpoW/gQCM1oNm+dsLlV+JUPKthtYC+02476gh8hNIVXVwY5cqjl4OPFAS4/V1D1r
XZHb2IyCPyH2h+j5/O+7uuJi7QYTQTzDBBLfwpVlXttJjpBD+Kw4b29KRL/DhbCa
fGszvyuyDKl1PKPt18V5I3cCXywIh4wilN/+SnlriIaMwmYZ8gz6IHUFqxSWoWID
VjtZomiix+toKNR3lz4qL3KLfHFH5/WfKSFqEdnpVkh/JUno2XLMkk+6XV83jH6K
yzDT70GKHjBE5FG2pDTM6UC08WzBokIffIZ+oF8RaTqsoBzIY10O5wB6jPtbd0/m
gie0g4IZgj/6DvifJz1KM6xnwiQ3b/T0dqC06bSafsLk+7NKvqzLLtp7XtjWCrtU
Lh7lsJQnlylqF7eYNyZDRBdnTMfuQUz3dVTjzGB+O8494fWqUpTPktkfoXpfcWQL
6bXKfoWAeUh6jlUj0NHQhOLJonH9VMpAXLNaJXULmCq+ABo3GxasRCyUbHXMLHq9
iVpIrUcGS+8Hllw/Gt9kED6rpjI2seRGSTJS/XrNRK2HK0oSwEonajxHsrIJkYuD
Ch9E/kPOVi5lTR+7waivH3QMBUSSam3DNdS9jTJY3D1GHlOZx5nXHfN8+7MtzeUW
pGb+fO0RCPFwiL+HWWD7gnEO2JiK0YpTlIfIdHUZDbG302/nubQd4+rvBcVzr3pL
kgf6ksr6C6sBvjpcmh+Zm0bMF9XZ8+FUloWAG60JLM5B2skrBeRvc9V8WMZ++BCs
6TsTHO5/u8GO/eHBaN6tp2iBNLIHzv3VXMbQ87SQOxTmIVoCSHoLPXXjEV/23b7L
0OBIzOc7LYRccBw60krBi78kgwI8ub2ZPYKylvpPHEANAMVr4GzKj1p0/W+F9Oa0
GEbtekRJ7QgT7T155RtLdedsEA7WOK44Rj35yev+BI28/EpiG4qc9jDN/2Y+AgJw
Bmrq6DTxI7ZvUdqYEH/lKDS0Q3RHt/keUvIDgo74YhwJExH5dKXUAD6peNeULv3b
gDpQigydC5WBX5V2MuqO7CB+1WCyFfg2enRv/MQBWlxMjz7VZosRTzrbAgYR+i8U
TORA3UX2FdptI+/cg+/NkOmZ+aB5NTQKXSwAfqnYCpjs/DL0qLf5QYA08Psaj+7O
hd3t0NEpJcBkE64dkp73hCCLblCas1vPaNa0TwCzMzmI1zg8+kHSKgw2M7wfg0zX
ipUE3agWtvAuRb6BRNDEn5vbeRv6uZyPXYxzn0Ukc/dJt75MQaf7h42WU7/edIaw
xrXvCHka+tJ+g+bXucqp+sBO3en3zZq7hswbyyOeKo3V7e7ao1SV+JH+5MylJoCn
/yNccoToQHCVAx/BpoFJN7uhVEPpRyiAAr7WQeDIaedTO/LjoXPTYr8MCmhCGwJp
2E+GYxE5p6nA1sfi/qxJQK3Lgvk8XFFvCWr2K4D25hsX3wARNwtEYeQA/lnuhWbE
6bMcz3y4D59AGtkvDFcLIymU5452GZsvQNkV1ORA7oQqbPYFuTZUd6OpAhSMipYI
9DTkyPRM59f54MMZvAflQnSw9o4+QpoFdbvGnciSKW8x65jVRB4tDUbz/gOW1V/G
+WPwUtWMUvcX5XOmTi3V4xF5jeW9qSErTOCbNMwTJm6yOmWpnrCe2NGW6DILwbEV
eRWB2FknW2dJ8I+X/Jr9zo9U3iPa+8lkiVDzXvNpn7UtLvIgUIUyyV5vdMbTvt4e
LdFFB+UYvBkVuBVb1KXYQlLWU5yDog7d223GlqYj0SduRq4n5Bx5Vyfb+5UHn1tf
YCgCxuytd/+Pct5R2br0uSwtV0LIHcpDrlYODfIrmXba+r0hws2jgyhlEolpKEDs
kk/LndufCMVVQObEEtj4cl8rsS7sMzEHmsK18hyIUk8OhV8BvM0qHR4E10IZ23Jm
ea2w1Z++i4f7AwjBQlfL4pr0BoP6W4NaHY6EX++VVhq/338zqr8LnpTbgONJbdDw
9/TUFTdTQsGphLJ/gTiy8JWE6+9J8zMRd58Umbbd7c4j0DVjMoTD3CcZOJWQuPu5
1E4s9YvUVkDHi6hfh01XMZLWW0S2DbyGB0lDAtZkjpqs/fiNP/JsJ70+MGjLWRNr
k+K03wu4dcmxFkUbiDvU7GdA+GvvvoMcBHuGnV2fgD8QEyUsWbrPEXxnwJccmhIy
cD/j6+em2lNYyEfZsPacz35iEOHyeqs6Rqxu6XefOFSC82YVILI7Gsaq7OfQt9Li
3+cHuML+uXbea13ZV5UL+/bD9oYhg0iTfjTOMObCg2voUeRI0RpndhLmBYF10XNw
9gid3rbdCTebzz+mdbShLyf2s10NR1zon73YkpwC/lajT0u6vf9X8Gg7KsS/UC/t
G9PszVCi8s8CUzC4MLDzdg+WSRVqFvn4OQrIKU/IfQ+Gz8CrsoEmOEkNG8t38myn
pyaUsXmk/Ei8ihwLQhhyRLuhnzQ9Czvbv4Y/wqgHDxdUJW/xCsGRvqIq7SOS7Mfj
h0cM9KIopF3rxEuFHAFTXqwKRPwuoeTXEllWRHPC3kXYTyMlb1TIr+u7hBzQbYQv
7Rmw2U6SqiLxZ+VmhB9gf0zrF2JTMooUfInQToZ0sMrTpWSHCL/BEhYeVDU6I6Cg
DWX6yjJJoKCcZS29PiuEVriSaP+qY3MPvgsJt/3u9/S9WUqZQmWiU/lJUB0seKXJ
9JNFil1S7mdUEHh+cUfdezpVP/MRj2JqBVM2GZOc6/e36u/1RSgfkwDCfJNeVrjj
5vi3o1th5Vxuv1bWCSw88V0eWNAj/U9dUtZLOEeaWiIkogoo8ZFKBdAYWOD7otEN
qlsTbo4YRIJQq2oLNSJ0mlmmvd1Hgggjw0pTDjvJ1mgLB2cAKIapfd0a82lkHLUD
qQmXyQx9rEJEdZD21bC3zWL6qgr82rTOBlV8mHg3jzPIL9hwvsjPwnrShglq2e1l
RCFBm9nllAHpP1/W0iHM94kr6KNK6wa6fK8JqxXEWTk1sj5Ut37WgGsIAhhus01d
W4cQ1NgWxnvR8fI1rluuQQss5jEj+ltX/1emy3h81yQEkZ+hEIoXA5zXIk9Faair
GDBF3xD7lwBucvdfH//cGC7SmKcT4N8FKk6SMt8+ugqQRyngKES6Q4D2oB+awxp1
2FAci4TigBdfDQjAxYolGSZyyKGB/OAtBqqA0C/1hF6g9LSpFgStUcADEd5OA6gu
U3XlK3Vhqw48ySx41KUQTrdlF9RYxpR7vcgZ1QvanAVZekrq8q+CNmsgf5IskBHo
+NBHlEnxF6lSc1nAUzs7UKJ5deFnrr/NRJh9W3j/kbYeYPdrdzwKRjQ7uOgRvBDo
lKy+/te+1Vd+IR0dRST8VMRUF+CuROs9O3ZWoM8PWGCoCxTT3D88qHT1YXECnvD6
tSyrgpJ7i1hJ+dkH2N3/Qt0nDJSdE7Luh9MGq/d8xcqopXcHUG9fTIpuZZGEQUpA
d9Vp15aAlRbU6spxXRhnWxIoWU5XMs59X3dMRTUaAmylNrh0qfc+HgOdZ7IDh7pr
8rdiJsU54w9oXcZsrKmhlTCBwi9+v42yC+Zeeo6H9jLaPf/fYVs26jFs4jL4mpI6
g3QhzIa2GyBTEuMYgHAXdEUBPPwMH2onZAKjzvIYRRIb0++d/tDasB+cxHcaLp+k
z84C7TX/lCvq/MJ4EJWTN8vhssmfEEgcF3s9fnqUNl6FbIC9AW2bpChGMdrA3C/+
PjU4E0M8dX5m+1Wnukn1hhiF7sfzXTvZE3JYe5AQjlFJzr7fkpMTNdqUtPigBEyS
/qQirq7Yq0qI2FuuDYb5h5FfKr8jFg0stovFbsOUoeaQEfy8lwai5AHv7dZYccG5
81u5Vs7b5k5q8T3KUjK8KXJloINdeLCevUZckmP4YzirzC/xvHG3KQMjtFfG5Tmi
l6ZOWihmodIvLAQEKoDSupQTmyz2FBOpXn9yK+THPpHmpTrSGIisvzLgT25fF82P
DL9DePbVnfn+mvbQDOjIhiIAKM+zFjhzxQzYmzGQuoCt5GwknR0sciNRIf0p1aX1
Lxmd8UvB5rFVyl1rw0uCW10it37W4fyVXxvuthtxrzO82Fd/egEX54eTXklZW0CL
A7dr3K2eTxdL4Huz61h31pKLpm3Gi+5OXHqmWDy7dqu9PborV/bOuNUQVwbvH1Rk
1cYqQKLROTXfbAZ06x+1qujEFqkpqDDd0q1rBpZ8N8pqTN5mqxc2HXl0MeDpoIjf
NdnAH8FBaPfs1Me/47wdIQbU5NnfZEzk7q/s02/rd0nFQQMB5YscpQKcDNOYwB3Y
UlahMnLn4FAx/0MdSoJ3+HLvtuPe80UrVvPkjJ8Jg7zN4vyILLQHourafScB7sdM
gpplO79PTGRltkcLVp+VyvJViQ2Lr2036Z2ycqH2hzT+tzByYlxe99POIIgQf84c
9gGyaqlRHkpnqsX2mmzu1fHDxuT0Iqz94HDbHyv08Bfi3IdYyl0kANawGnBe/emx
IIZwR0KhIYHWLxG5Uz9J/SJh7sE3ytpv63aVCtWAg0VQ3Ag4eFAmq8IyfJoogLSX
/nymvK9f9r9ygLFZe58oXQL5tMDko2nCI085H37OMZ8hRcNZ31p6+u4OnPzj1xbJ
B6Pa1Y+LCs8oMfp0Ruusj29/9ywhAYklGcdbBwv5CJaTEz6sIhkdgbYpmIkx53T1
ZYa+KbMHX2AqqDhOz0AYiKc/YrnsPi21WQ+lEJs9OM2oXA4JT4J+IWIX1M08J94Q
Uf/FczXJBMkuZHhsqgdNqtfr4Y4Vb7DKIquT++wMiS17xv74kpkHgstJR5dLIZ0J
U3FZG4QVUDs1aYwxUjFq75ZJrW8RU6+MxAZFEfnKAPjTy7eSydR4tRWBRwwQh4YN
ckQQY1kRqPVAT7MAaZBdfnohQCiiyS1KN/hMR/awmRFOQ/TmeRakRwLer4zfjpKz
FhoKFOk3+eOSdzSmWGPI3jEsq/jFj30ZDT6YNGv4KI3UW0qGUiUgB8mM0wfCsrEJ
F4SG/RsrVZ+kRJPsacFd8Finp1sCs8mCV1s6WwaFBgDDdVL8q04uBYemeIeSNN30
gusPl/e6AtevKuVVoGZDR78CWZ2K4MjchY/8OVnAUUtSjH1IxeLvR2dcZ/+DQowg
jtjSHTTPLvewsrWBNqOAdbVSfatJYnseqeYPgSLA/TGSNYYFq/oz19XtZbbwuIWp
37YJguG6Hs4Xxs6JqYzAF4AoDJnWN8rqxwyTt9/Bm8hspDTiWNldxibPS/rVoIsx
5OiM1SS+IfZ7O+uwhsDi/4hJCK2XZUu68ZBC2twBIy7iQAbW970VHxMGkaSmgIpA
NP7QlMVKqyOIDMo/OCt9kf0pU/ByUkyXD34RIExeCvSoT65l3E6Ts8ESG8FVYcHx
L87CCmugesQnFRbCbwPrIweSbR86l16WxYY79u3yYgXNs9LbkCUHn47elYuc2BBE
bFx0/eBTM9FGIJwn6D7ZqyBmtugg72ymgvwq0sBFPCz2JbWSwolh8pBx9Qb20CLB
m4bii9IQn91gZYlugKoOWSw2XzYOUEPZblfBrIFeBUllc9OebUMRMmcpGuY1JU06
HCVDXHImWk8gIvNmeoKJXg+jQNZ+IxVrD/qL3XRC3STd+mR5/cVmxTGGbONqtSsz
uqKpGyfhF1OxCGk+ajZP8HtMA1xOfs4d4Fe+1hXNP9Mu1ONnsh4fD7pPtANbNVV/
gKqC6uP88yIvEq3h0vfGS0tN3RczFUcm7xqVZeHTg4JPoyI5QRHmrYYVY3zIub0C
fhfgUI0am8KsBfwAMtqKkd4gDc3U+GZy8hAN2loy0fakCxXwqlVy45zKVqGSHA1m
2nFxWbNEhXG8AwP+4v7+VFTmGP8KGjkLKA2hIXbZQslahBHKd2jWwj6xDMKgGqxV
Y7y2Zzh2UTKaRuGrbsI3Bq5IIsGj4B3ZE9xQ+XDgu6MZQV8Cg57gWExJ+sXclWIP
qOTvK8aV4xcGcEd0JVrnnFNES6tI0V+FNvzAYjNeHyJfADuVj1D3KHQ3o9zgZ5VV
l3mU81yri0idhQ/vGT7AnJXTjl7q5XsZPOlpIz/hDviMwMMRLOBf8f/yUKk7oJKI
6AbkmRnkth9NRDIFm9PA7Vq987JmUiRpXybkyd+EAXrZxwLrTe0KZBK9DfFBVy8w
HTaFK06/VZsmhtppPejEGhEwPoSJsugcRxGLy4GaYvc/j+EOBm3B4NJr7PcCuYcb
Fxv5fUhcfLlYlKm3WV5csZOryBgV9ZnELDkx77RuLbL316X9omCm0hVq7rzhgfYg
oQORg0+wf4wUOduP/896lNtsn3ziynKutg6zlcbItszVKb268NM/XCWfUjL8g+e7
CVBniAejDGLxl9ev5g0z9vFL4zB4zqAhntLhHOIedSndVchn0iNNJXzQzZMlvjac
odiWf60BHbbA6+kN0fn4MuwhWBbhE6msuk3BVGhfgt0N2oBNP15x/ObmtFKjXCA4
3gPYXZw7aVPvf3b2ML7LqTwqnpOW4Wc+edBEqJKiq9SlbbVxtLzEyMkKNYsNM6v7
9yDxwSl+l71SkEaUVdyaSRSM7r0Lw8Mmp/IqpJVbtYofjR8lxisTHIP1KzXbuD+H
1k21mlfjlZhcBMzKdXqtN9vmoEvcHAv8Ue1fBq4QrppxXk31KE+JuUZAN29r0iV4
NW/a6zNh2deG7m+L4+9kyc7drZjbFfx8X9X8d7/iXuhBd8x+70WMSCTm7tz1tZAP
mmOILPhyOR1w3PYBODo/Z2Fi8H3/v3fsDzxjLOdy84Jd4u5H8hdlINOB2lDn6cCU
GqmVI9Fs3AAjATylYOLDvPe8xJh1ydJr1mJuEj10QY0brgkhskoiiueZB3C4tBB3
8CrRqAyXGRkzKjxZN6OVC10PE85rSBGOZVwxcHhZ13sBfLJKXVNBQKzQCY1FBzRp
XM+rgbgZfzWE368ZN8RDDTGJGbd48CoFhpWsMVZihpI1ZDYo1h8Oy1hbuCLesLLh
TfRx4GXeUhuQOAgFM6wFnv1c/+EmhgSvCgDm2CKuf5R27cZFSb3FioJrdF4UA4Up
oWNhYBb4NWfyGR1iylO0U19l4xyLPPzEI+WiegtC3RdXbmLMA9wr5iKJ5oPLidhw
tPoWjUebo1nhWYe+OD7A7aTKKqjC89/RVx8f/Y+usXBrK9uxy8H0g1c3mK1wzRPt
wR+0JcTMZa0LgKqRifDes040S1/+91te7vrIZ5panYBGhQkxXwQczGlLY1q1LFuv
7pAYYj1YRBlNUcngiS6DvYvB2m9wh6FiwGgF2cLeX9q5DP5kstAbrRkzQetsX2dM
4H3LRUaL+aXv1c16gEoCwQX38zjt/6zJHEoIR4IqODjs4x/b2tzjTjUjgPIXOeqP
aC1K5spYVcHJQ+GFyx2abCySgz874QpKyyieYhG2g2TJGnD6wEJp66YI/f7QPjzD
v11FcdREOukfBS+vIcxttGpa8qwvmBnbW+GlnotCFXfixzE3azL8zBO3KASpMB9g
Olm0PWEXj270wIcyeI+bku51qTvAM7Axtgm1IjtX0Qd8BAcA1Ufp1cJjTvYB8jV6
IDK5im+gnsr8k/vTkj03LvTy2OGrLn+0uoY6caTx/dx9RckX4KkvIhM2vVaJqT/p
sCcDUyd8kedHsWJfKQjVv3Ijlkjc958u6MMs/lVccxFi5EFKGhTa4XatZfCTWWAL
b6+xJhIr9YkNqZlDGMilMyvZWo2228vSeOw48tV5Q0vk56TdKsRxOEum+nJkxVvb
PHjUo6KZjLCw6J/9giBTq4BSuYo1xLDTewJRue9+1weNnZ9VNaiEkkSKqZ/UW9xv
kNSS/54nCrkqw9DYI2IYa2NTCCZXhkEYLS2WdASJOXgB8YCH2MGcgrNEOIsuPMSr
BxMC6dnfkTam9js+lCHwOyEmma+DVCTlMyQU0WnoTPiEFNpDf+VBY4WSGiaaBqUh
/wmC1OKsGJcknnLSx2m6C5fVqWihEGLM/E08X0EIvW9+nW6hdFLD9WD7xtkSSywE
dudgoW7h6t1ExqAcjjpBfDD1xeuJ23vtJOrqAqN0WWueG/sfcHtWbcnU85LrZjw9
ElkGNJnLxyOnSsLfReh45iUT/OJ900/IgUy2w+l67wCOAIAvFqufN9VBeOmgUvxs
5nTRsBTtn1uI5h4K0BNAsKsHTKDt7FszTRK7MrCcoK9RTd+fGmGUTQFk2SP4qXtY
ZDpr8FLEY/UzfpjqhRcl/HuPCAKTs5ZhWaKsW+NUTW367BXsLK8q5xmyiXCevQDw
ZAZjY0vwtGP88U6nq4WZ2kThJ2cS88wz38zIg/HdVZJ+ZWy9ftmzq1NoWq/uYWAT
4LxdmvYR7gTmXUV4u5DIEh/NcZeaJJGh9B5GIKUghTzeZOWPqDbSXGRjOi6LpKaM
cwxOwiBn/SMIh9YoalqPU9D6BjIS2pk7KMhAGJbD63XPOMLel4S5DXgfYtUTweF7
K/hLoIhFlFDhr+yhH79a+a3Dkb1g4T09uAwGgRd6onIhJIwMQ1tt+UIdcA2u1cUB
U4smZqeCDRWIlthXRQHLsNUCf9OGd15E5Zdjy4xGApiM+udw9Sx2wG684YLJ1nFF
9K2wksKAuKG6V390wVsu2SkyIt+NSOku5S9NtUEij6C1RoRi6JUkbfZh9OhTuXGv
w8I6bujAULKHLQA3fmQizdUfwAp8gnhou0F+Jqdyvz0h8HloFTINyWQp1QhqYuzA
ACrJC/QLgO2cSc1AUsTSRBPdzU4hrwEoJTqdHyTri7gZ7ka7gQ4BI91I+S9UsbM4
LNFTiS69kG58ZpuN5ts6ryV3P1g/yiXTZl7ZjgaYbubL5W2ZWLrSZ1YpT0K42EN2
59RFpcG+hQ0epBbQq+Juj0h7KDJfAJkHsErlt/kMUPyrbbTJ5Q5KqjPHYY/sRl5l
IWR0NI0l6P8YQvqZsDM4HeagjCPHyLa5H4s/y56V84J/BZFGU5sYFzKp6SNRBWN4
YoxCEYtNfn7OPLyi5KvXwMJ1dO/ae6Ir4o5z0kfD/QTSUedOtXT40jZbVNRxq533
nSw1eEsY8KctzhJe2ubveXAu/HBP5pfHlDiypHYi02t4y0HSbFGX4NtYjRMFqTJm
+TlyblKfOPsDi0QWSvdREzaffDd4lg1y/BxO/YlWwCgJ/XXCv+XX7gmK+i6webyY
dx1uklYxvZlvRx/gIkNjK5ui4Cz/cB3v8VItig/8ABWHBYhXLcAl5ueRXButS38Y
DcDnCLIv+Mb5NuPift5xQYLeOkoaqQ6JEzA2PSWEZLMTNXO7az0jbELfUP6ocd0n
QXRBJkYk+FYy/Ix7F/fW2A1GRgO5kox6L/D31WILuabAYBARXT6vjTUWCEQe5P2Z
088R6e9C8Gh06pE7XD9rLIxb9Bi002jp1njc3N8uaL0IbiVBHFZWUO0Ti+NL0AMh
N8kyaRcWb2uRdfvs/U39OFa3FKkeTu1W6VrfiBVEuFhhsF7Z7XiZtjWuJH1nxf6o
+aqTAePhKhLpRl5NWp+IM6Ve3yTz2b+Qf4Zwru1eju0/uLA6fcS2KO7Cq/OUyGJR
AsWQQ2I62V6lBd+wECb+3mfV7taVjVZVJfVhIBZPMgCUH9nLCDnU0usrurVzdEH/
kXXNYQgamD5g9aB2fjQfr35Ffq0uY2FQED5fUUPXxyHkwWDUAi6nabVZ6B2HOu2k
7b9pjW/VSWqUxhN9b9vOPC6mUS7sPY5F4Id6p1fSIdPHe8opmTOJ5FhvmAR+syvk
HpgTHt0jwwEAZfqAo55DnE0kwoTf6ALNBsU2VtQmFWIh9Rv9d1afzevD7LjQUa3W
l7oX9mPHqdCZtMCcV5gQTlZRdOI2fUA7098JmKlTZP1v2I+6pVxY3JON0/7NzSIE
kQZ7H/7l6BuyQ6HLR6qYMGskAGF9qjUi3TsKi8JCxPkPVrIqP060xjCNPeXBVlsT
WXB+7pvgrDRKKzWs9D/bHNEXru+RDtLzR3IVWjGpvF19oNTCPJSzHT8rz4ZlVhUU
tanvTFfev7QMgXmKDy8oGIuc/A3baJPVeDc6A+ftlmXL5GGnb7VE/RmMbVLIJE8P
eDiAF1sX7aDFfTKXShcpTzFWMGhZjIWmT+SPJUUj7w/vh/tkjsUvISOkejufbOt8
jaJuO8TBHupbAPG4mB8ixKyXS5rwblaRnjUsDelNs0hJn9EbWp6kOZNnpG1fMJmD
VkL9TUO85+8sY0Q6r5apti8tq9c+BjMO541yfyeo3No3FrawRO8mn/cHuwrqbVKF
ZsuPkuypJXPodXAIB+UA4bcOu1xbnZw1T3O9RaVZgNPENm5ATK+dNIlk3esm93K0
25goC9s0dU9wrKB3CeGJjR+o+mnPtt0W/PaVxSHekCbFhMV9BdY3i2RhiligPtSo
UcGBLDz4eG0mLI1MdUzx40j+twG0FCwrgJoPIiWup0OFEqP8AQUJchkFF+wOwxfS
gsNFjWKOFDO/djpp2b5LJ0pl5Ige4f1gXjzkwI3V1K+jgMrBisfmo2bhbY4DGEiw
Y9iYy8a8qevXVwiInwvqUNN97jom902y8JcVUUhJG8nJxrEqCNmWJViBfqVCbQUL
uCU43KoBrupM6rvz20MdupYZcLcJ7sNHn1am6r+tt+oQq4JkvPpP+anyNTtq17D9
u9KAC5FrqVOhp0T9jnUzGqk1mYXiw3+0A/ipWaTywdDHzvZdP1kGUoYy8KiHy719
qiCGKM1ua/fRHlA78kRXwBYvtE8VCGgxPbvqwEqnvNAfgjv2m6yg2YQjsZVLrlRq
ijm4W6Jt7HBIuj9+2fP0vv/IhN27hhKhm3kxbqQtqfHmuNvJeDjFqxpHWrmtwaeB
SbPsyeBZXWa5ThkjwQ1nH4WCASawpSzVnPph8bqkHPociXPxVOTLBDBaUA8XaQbW
RaIYFJ3MQjdL4YNf/j7qXp0ztNgL4wDFRg9/yWGYpQhDxFQZQMSlWjTRwju/9Iab
iiB+pQEtkzZw9Rxr/H2AcLonMupJ0z9yaipM3tAO+nZyMtSmsJsSQggJ3E/npN/i
pdMVK9aiKIup3W2hVRH5gHoIAf0/4FAitxlXg6Gd9vL/UoTukZzmGjoYQDb7irqS
Nor5QQROeEsW19q5pUwWKhynPKLs5QjkNNl0Ke6OQi2QqUpoMIMAWTcetJ4g6gbM
IxhZTJxyRYHAQCk269QJEjKQ/XqWG6g32MPfDnc9N9147vQndq6zc4v1LHXxAq37
vWX4N+fldS9gAqXBgvW08IMA6Jh+4BgSQ5PzNNo8nsHrtZZwN2fSybgm9SmlxjLK
+mTMM08FUPNwpKIaTnTCAWdIaYjpoqIO60u4iwkMYbHyt/nYlpkokr+oS3TaTdYE
XwQjVQOawVz6NLIUunzwxw07K4PNWGZwHm3Woj0geCPagfmuJynsSDxN5UHidrcm
ZIudv4jIj3HmXP1wF99v9PQ1nY56BKDEs2YLB+B2YyF3g98A5/In/tMP6cxr6n0q
D4o1MXe1ViDxdEhmEHuJcYD96Iss9khI/rTOrgSnXmmx+qUbUeXGDu/PTIdb0Zhk
tKAxkcGF7mvsQne0Oa0ebwv15bCZ+6R593TvlskxhL4j52667C+7sYNmFjezLeKa
xzqIqnRGAuiJ0s87zg2tBjMw8IsNFhv7YSH6GqgIeSyPux7RhiXfIjjfSOmq9Yrc
VbHRv7QCtAG5Cq3lKNrQm/E0VI4euZS2moIfTQ5/FXdsHlu2ZXCHb3tfxNvbzef1
zsnGmdxb2j+lJTCsCNDSMO3fn3ixVKHkTpq2iowxHiz54KyoApoO8kTeinlcYdIu
co2wuYIea66eMi5yADXgNeNXnWX90IeU7LJYYhoeGeooriPx6+fyZRH88lNQaG7P
4gdFx7cRSJ+8h0OHkv+zZ+ShHVub7QR1kiwzMGxX5nB+qhtjG9OmnRrO1HqiCtP3
yEnCU5icoL9qWgP3iqJbbBh1QDOVIbO7ZQrsJfU+JjQNMgW0QusVlQ5dSj57tKIt
RMycKw5xMAobPf48WoKUZDx7auut8rceXJG9Ee3tymM3ZeDNlmXGYM6HdtheLl8C
M63ESyvswgJbrqQqMU7IcSGh7oI+bARe1LBN2DZFKhHB7H7uqqrv1nxAOmomUX9s
HOETHZzGhc43qF0mjul1fP4aVjCMEok/xQHNumzwJ8K+2uoIhpjQ7TLtut9EX9+p
W3rnu/zHFB2iKUtLAldiPBwkei0P3iWrI97+/2W03Vhs2ral/aNvLNVboa7MELtM
obEdIi0ltjxKFBA04GJjn3ichd+PYUzIrysO8gRZ43RcDLhXcj/MZ2wbik7XGx2O
wwIce+7zafnQwG2sUpIxWTnoyOLaypU3EeE8oXLt7pQegqJEjjLpngfSmlX1TOWh
uF2i+gKDM4sC+jTkvwzYkIlvK5MCtxYb0kJEL2gVZSdH/F+UZW32PQdm8My8jDx7
INt7DmCuxnAJB+QKOnGnQfrMlTC4s+8N7YfoDy4lVvYDUeUTQwoxVFVI4sYLA00k
zmViD0FZVoB6tYBjoSG/ZKfcIUexlnQb/ufzNp8y+ufv8PKasRwbOymlZ2XogUBd
48qN2wRXcrwTKPcheaWJq9t70u0d7GvlBNgGR9j8R5DyQr5MWZmOYsESpu3YS52R
CZyCePRu3jU2CrNfjl3wvh65pvYWg3r8j2ieIcmawg0UWQ2pzldl/Xd90BDVNdlp
9DMpti31zkBO7HjAh9sl5HCIPKPI5JaZshNQTFRGJ0nw9MLDmzurizGqExOQPYPm
ljCAe0phGOHWHk23P+PQsWOJaZLBed1EhZasnEZd3RW1WbwyF36v0P+fwl0UfVCR
7UsQ77vFucB62bQ8NL5ZyNYsc57SVyEV0/DJPv1Hacr1uQBMEc2GJcKpxnBuHGj0
Ym91Tg7+M6PIr7jkNAdtE9KFNOCX4T1pux8Ovpp1DuIwd2Ie7PXks8GcC3na4//5
B7qHMMW4HECR41xnnWeNAF9iOIuB5zdr/gZ3oaau+JHLz0MfArH+mvc/m5Q4GEw6
v1xu7wx8vbzmlNEVbsUBmneg8iIY5G8f9AS09v1403G83PThUz0ZAAbcHW+r660K
Gc8FJPDcxdyzgpXNB5sM5zpRYplu3gU8aOT1gm1Z//QxF2/LW6sSL4IqPSyD3KJw
FCpUjzutIfxbDDakXvpUxuKN2mPCTNR+WrLvwidXjzVLFY1HYw2wVaOqq/Uie4wS
gyadGRDjT56yBH42jPtaXrqA0DxbfoVZE1TbXcbLzkv9bmlUcNeCDhUoVD5SbMPX
2orH9VIa7XMt6YLXTpinZuB2N8Z1LGyTQXKnRHXvTYWV1QDvppLrGzeL41yqi4KV
0M9bRjp6xG0gFOL88mjfXYuj3BrWQ1OI0ljmvdkbbWj3ksRf+O4HCTHc5dwwwXr7
v1MKOKNEGnnQ+klAP9UB/muMTJOcBedFprVQt1M9M5eYJjKGKsPZESRrUMzy/Nol
508jyVHKwy1nOPB7Xt8UjbuMjOeEjbB6EVlG563wPdbjFeWBDfogAuDcS4sRFQWF
RbXf9eZuQv9aSTHvPnNSVSsSXk82cwGZjOgaRpigGecUqwzgFYCl8xAXX+RO5PAa
iQbsoWPw0b+hSwczOBIRFqyvp/2iM597xtHqwMJal5IErQdNjYSdHXEGCWs8A1pY
ZPh5aLrsfKnL9xEtrAq/fXnWiufYL3dlqCdx2ZO5rlSRVreX9+KfBATmJLn8x6mH
0/ThU69UCiViXTV96A8jUULrFawA/5YcAC63CvEm4sRoPhh5MHTw/b6THKAN63aa
dpIkUaA+DrLxUgI0YIELbStLdO/qR4pMSM7cycOJLfCjPCHw/Ztw9ZRMm7oY/Dfm
1GZEQlLuGze1BL9BXsAhZvMeQUnV6+ejW+ZozewdcjYMozoAONyMLjwcLAqK4ORy
d1a8IcFBZK5L0sNX815T7RHYU0jvEmAHlTiBN8CaeHKUsstA2T3Gh1iM3r6mFMC0
uE4BUoR2ww2S4A+ImMS+JYH0Y9LiWTcacWLpLWS0JfCvv+qrCf2j/7NDaVm2blsT
T9RUvGQ4IWhCm5OuOB9lu8GQIWKncAHEu2K1olZP2IMsLqEqAXFb0EbPNze04bWL
zKthp8mlZdg+4V+nJaVSAC+Rw8xGugJ3gK1EdBB2UCnlI6Z4vi3s3JMZAHjEx/we
re4OsISluk/3dcNqtayHccZRa4QipymRyBfjB96MkwQz1QfZsxT8TFIBPJZ7TtN/
MWYUmwVbTn1mhFD5zKR0A/eSaP5KHSjBF+I1tyJ1k/uUDZqgrIN6ExbLC6Jdc6IL
krb/CYo+7A/G7dSl3g9y5SKZlakI5fo1hwpawoS58qKl/IQSXTrpMXwipJE4fFs5
MSYxPdAqpITxm/qw3QcVzTRxetnVirFWfoOyC8EdkrcGSeTrV5IYpZf5MPVOgDRJ
bTDYC5fnvFrX3HHp4WnuuuRjlPgw0hhUbMhITT9/BrcReO17/JGuhGOE1o91aDg0
DJmfrv3MwHxSwIpMA1OB5mD4wQZx6z+yU4TXlcvH9YTZVgImbynMT8K4E8TguUp1
Ey4NFSt18GLv2bd/fH7Lc9HhhAt4YpxdNVCr8YNlm/Wlcele+kW0t2EzbKnhxiRx
mOYmFyI25XqDVMx9EvtZWNGvKXsRNvwN55mcAM+P9ojw80lXW9JYM9xkEVGo5sOE
HZa8zeXAV0j+RZxoLC0J2oGqJ/bfx9q2qtCrwDfiq+e2vRzRap2a1W/X1HdRuyGm
1+sSar+4M8mqFhiLO9pXoIdm05t1tmsRvhn+ZCN17BodFM6iWR3K8EUMCOc4Ueva
z7KO9gHmado5qzcn+cthsXRViL51xqMfvO7Rn3RiRx/xu3qocaG4g7VbMgCRbN6g
OnjfKMBjO4puQ1t879qFwfoV0KZ5EbW6HyymNOjb3yQLD4Yu4YawWIx/HCevLEcy
cK68fKlZwcDrI8xqtOqw5q6G0fQ/4PIR+nGGwda8VUhhtv+uIHUdvolmuwpDIs8r
VlaPdn4y2HLmYVvx1eEQY2wPAsJsukv4sTW+r3M1KU+LieF63cWSwLvca4w2HIPv
VqVgvjExFSmhP4X0rND9Nzv9BnLYaFIxfglXgmGLcBJ1AaqXttosw7HXdZhengnb
UOqufI5FbHhOK5pvWbmWlHtcrKvnSg1rue58MtQ/JHWd55uugqscG77ztIhUD6NO
lp5BWt3dVae775m+wTmxAeDVxasVfmXBs4Flh8N7RMeg3WAU4r0fi7pWXtvYtzr6
uMEvanP6mnQI/WI44lpwTuYuRxhGyXZu1HHIuhAnBEQBsUPutjeFhe70XyT5H7zw
SbvMDvllz+06oVeDndm20wjXVcWWvL2a4qcQ+bV+lA4w5SHRylez2PmKi2Gcgo7F
TtjdGq4NaEXfMPpqhj9OBbntJ0xv5M4qNdhOtxJFhiCoTMehP+toXcliwUu6ew4v
Fgeyzp4Y/WEwyrLmD90LJ+ua19Jq4BLlFa3rExu23VI2C9SCYCI8FPDjjwHcctvG
1ugbyiSRPdzgmJdEWB2RjGfi0MADQZmcWwpS6DyO2KIdq8icgnDmxLAWdpzIkGIN
YKJIFe8QHGzlDm1vBmm2Wdbq1tkD0bHBhX4wvpFVAC7mfkyT9lyxehewW7BDgaJR
14rZa/NmkCh8Xaefx0zgs6GRZJt9qIoEDG6ouWsw5hqmaug+Z+abfq99AyCm+hZl
Ua4x3wcFPkC0Du0gjJ1v+SzBph1f6VLeXpp2B0+Nn/rTL2YNpDJSjtbKk4P2QZ+I
JLkE0NQoF2wfAvwVhZOIBPo9C9XME9gvOwWu+KKVaV2Z9rwI0LKhGWaySZ3gUQEM
A4TIe6Pl7Rk4d2eTlDjPrWrJGDvJnpvt0qK3UJjNI6vt/kKNr0sRoS3oKkiel556
10xFB8poEw0QnV+n5WCL/9eCXSbCFiKj4MswEg3jF3QveQ6ongt0+VvhjRJ2pWHO
+mDC8oO9sv79dCqu7ML9oUowCU7w68+hyaauOAaLP5LISUmr0Gd5+igophq8/43D
RvA6wZDJVJ8Cg1XySUcgk6i9aY0TpKuKICykS1osi+zxeG1fCFl7JUf4ZLSTEhO8
2v3NkWEPvF2bsdsL1WzoYXSVDPPhMWz9FkSOvFtRtwXnk/uUMhYj7+yEeThAYpKU
jdPFMnEYAZ3j7XY5vbYmPksh9Jbf0Arn1OdQETdvdemwCKTujD71U8mbAm/ThtHi
jsgw+KluV0IwgtcEXBlpY5YnuZnG2sjjSib8eNHGRXSLwi0bLu+KGdAB97EU6h4v
DO9OZOsalQP2qW1LAVbLkM7DgLf13Z95l4JU6AosbL6eHDEChJ8QUO5Rudit0ZBw
VMEKJpjeRo315lzMd4vuBG28fgM3CkKMm5YtG+YI+Y7gc60S2v1bW3qIbWN3FUko
DxafsXpJRrRN/tuBVIR6mFYVUE2Kg7CW8Hi5d6seDfbfTiPCznP+9OptU5XC3ou5
XwmQ3W0W40JZq5m/0aOofS1PCdYtlo+neWUziTmy7hOpe2fLFvyrlZgXhLAM+ylm
zwR0H3knnPurK2rNYmny3PwboUkzxcbaNfYdM6XOpg6IcQMjUjyP3GOTXG1f00zv
QD9FH/KRYgA9TYoC41n2wsaOdWhc4p17bzABtUNQnIpFEmLIsvhYaDumcSaToDmN
gRDYHnL1v/vm7sIgyCfg0vmYQFYDO3Qrpyrv/RlDir+9jZCDz9ZDmtoR8DNQe1Xw
cb3rvEOFXn8BB5uxGuw8zHxffQRL26sF1GM9GziBKHgI6VAJWRDJMNnpFbVnv+q7
33l8xMrK7mX5SnGp1mieNWn1vePexrZ2ia+sKylmqB3bhBLSCEJQ8ShcpcYmsxCR
Gx8l2PkzNPt8Yw49mdLUQ3swUrv6LSP0HIT9OMw9dic5E8XF8HM/2oHtIKSf3MFQ
asJ1glDjcE447175pK+n/+0tO8BkQyunWYw+VyGYHtCU7WwTvjTZWMhbWhH9IV7l
wdoxVw9HkzgNFW6KzWTJZuwMK0N8qoxDU/Ly2K1SJc7XQVzy5EmuwEJmrqo0stfu
+krjyF834kJ9WOmEmUYUNNHJx8GEQvYla8J3hlHqRV4y02ABs+DPHy7i2glRDUx0
SszWIM1iKVMJRmEk1NVhcrd87ZdkrF6y8EvmBb1++s1SIMuQq2CdWNJG8UQaqZHZ
KsCpnMn0+L2usblW3BX9EZOtL6oMinfRCaP6X46+izvUndv6XNpV71VZRKGnSvhb
K/Fc/a1MPjP0vQ0p1+Ybg0qzlgSAsn0f9WKV84kWhSLWrmRYcXQPFWmlb/Dco8tk
jBWzjCaDBub2hgNSFhkThuxst1azR2lJDe14v0Kir00gT+MbQ6hH07BkEw6Bccys
w/+oEKIDONMvCHJQQvzO30o4N++yTM911vxK0sXo6+7a/ltq9eLQ8Gi0K4XQJXTC
5+Lq51uSZBAUB21Mwm3NjP8fTR9isFtCInhVrWb9jAmUkgfEJzH4LyYeW3YwvSd5
8JkHXM1KBdEVJ7aKBp04iC3X4r68msiAdQXdlGNftTXDVu7iDjmrX0W1tE2CxxC5
iT41bZHLiZIOIYrd6VYaMahJRKOZUx+yWlCr8OLMSBJKnY6CesSwCnD3bEqMHOEK
SBPUzWXxc8SuHWZIOYNUrV4b8Wgr1dVH503m/Z+s3vERUKO8XRd8oAICaaxM6rm2
4NYvJiJ+G/uSwZFk4aO2ALJOxtQSDQLs+pN98HSIPcWOjDgnDapjqj6EU7R+u6br
/2E2Js0FF+Gx1c6KIecUNpxrwHiAOMbqv8m3VmYGfuraD6mLHgG7Y9ylJMNyYEM1
adj8/04qxEBvJHWasI+ilGSnQBPhmDxfZlfYkZlQ8wWMijlg0XCL4MhncBjvNfFl
YHvx8nEmLArCz4uMhUU4cfHYZKq+b9dH5uZkrW/yRAbxCsqCo93aPRnqJgLjCdv0
5KjpIPiJ4JhwWSTzrH0z70N4klvS3kHhYJEtVPB4KqTidB7gMOYxPY0s7kWLiL2V
65p16OqHERARy2IEZRU+djdf1PkkqkNpvJMlNe4ri/ttyOT4MEmQFlrs1rdxSZoC
18TrO4Zh2B9afwI4QMbF5HX3R/AaJ77wLJ72wi1yiqKtMibSZ+8ZHat+u32aCSkO
eCtN2wZKOHiBYV9epTFg7srPPoZgs+kwOSysE+QgsACM4iGlXm+WulyqQkFdFuMN
/+910aPtFXHyqYUWNj6xYYIIb8tVRvFr75h3ao4bfEmYRtgLVh6Bk65xtPM+l01y
G8x5FuLygZvLVKF9EbssLjUKAaxVlDCfb2n4axvPUB0h07MuwwTbXmKKwrMzOGCn
r+8/GLeD0JXAQh9DNpr/4T2r94qaUmBNIZ8wNZyP/Ar600+HXjO4JQ48AKJ2mCMH
TuJ0F1JvNZFhnd1yJl4vgxR4h8/LSQuIcGuCt8O8Zgf3MbZ1Ry8ZHNIhYzKiRCo1
C9oLPvOxDqhy7F8Q/KWKAcOTNcNg2eZsOPWy+wYsG3tQwmxukGi87M+qZ5VCQYV3
V1wj2KPGGN5yI/K80CTny0zU71WEs0BMk2SRu0JzsyCbdu+9EsvfOxY+92W0jUIX
MAvCc4Ds321Hq5W5JFZRziyG9pddTsxL3tFXK/qDMMdQAyRNGMSv9ESGAGFU4Nz6
8Ea7dx+AebOPVig87keMsx9fy9lnsMBvtlHR5QhJLS46sOMtdb50oBpesnbxX4ws
F02VxxLDd46mxqxHqbb1mQTbZtKJF9V912Gx8fpELxItgjIg/00MUkF1LiAWckyc
DsgfjqducDNnmB0/Z5y5CONV14aTlMqUkz9Rfij9/d1+s5mcAexlCmrAl0IVp5dk
Bf/DA5qmZu4wHWsAVv9D+wS1yagY5Pv9NGCOU7uh5cc6Onp7wGljRJY29tJBn/hu
XX1Np8qVlcFLvOhtYyLIbaLKa0x1aQD1W4jmS6t5FDR1wfH0//7rOM9TKC4wgjy5
oPmu0lNiNcPbo/PrS81fDkQhDs9gHGv40fN8gagZWAgvYfzRXun/PW3vSBBT5HWW
DOGKqviwvmM5ZnePYSYCNRamTCAahXToZH00y4Ws9zvRO+nQH82m49A4FP7EoAj5
jvrIBOe/eMglFEklNfKxbJQgywJOfwAK6HsW2VKl7m4HETpQJMTtjKC/hi9knnHN
+YV1gNkrogZKFaCEuQToC5DF/JPpquuRQr6I/B1GKMKyKBATUcBxxQ6JivV0myHU
hKZdRDBv0mYwTpG3+LBnL/8sLYrtdFgkyu6ftwB8QUu7U2YqOEyfTusH1EXKcA1g
6gpYkFW4me4RED3k77ulH7XsxovmqCxivYGp0rgIqw/Ir8qACZu/E9YIbsx431Jl
Sb9F8yTaAklWO1gUvP6gwnyWXSwqz068CSVJyrESfKlL1uKYi5Y1s/zYos2ywba7
5gYWU7lbsFBEFDLlADFp+x1YWp2/eBckMMUY/nMcyXDNYgCDxSlgEnXbm9qs+XGV
ooVFkvH8y4QZA41pr1/ult1rrYl2sB6EBzyZwsYEZD617fVJlIREoRzMaJfG61/9
szEXnwQEU9vLIhQWO5fq2nH7lmMV6wlWRbXVoG1xFJBos8cI2754bRZyxkLQNMmW
GJyezfzSxtOHJMzW4dEzoOpOnFrMVjgX4RVTJsOQMF2oaAvT5RbBjCUxYbUf6L13
VO2tK1W/cZMCI5bcWL8JSFb0HDdIj4PbnbhSfqNqwXoXOEu1aTvnjeDx3MOnF07E
xL9kJzIswH4W6Z77Mwg9Aeo3bM0Tk2/MHwZHSJzGR9uJd6aMllsPe97Q1HDi26PQ
rkWGOBksmhG53Z18A2wSkMBLZCwwSNX2LwrYUGk6DrX2wNbPZJf9HyjJ4oKy7RPm
UvhRmzpQoZ5e9PAFl8AmnCRfzUhO+HEYQMGEEx49CVHdvF4sXNeg6vVp1Q8KYjAi
56p1n1i2c/jxmXtVUEL1SCju8EbxB9T/pvaRfO9QrjfDN0Zyun7dCuov/ToL/CR5
oaykk7rhqQoYk+tpu1oDrZ5CE2778UBYVqPCadGTQF+cBypuTG62Pq9mf+6eYs1B
mZZbyCDkxisig0B3SJ/XjMySJazD0nxfk5CBQFpJHxozdQBr7ead87tnnEbCkAKQ
P99/0xwQ3VzBNjxnVoBMhiIpa8CYYo0xGgF4+FjjsTmvKHA0BpYcbzqZ81LKBdM6
LDQR1g94oIZxHJwZqBWXenf0Lhf2b5Y06pWHK6wJ6ylXSb0v38orMbZDXj2aXuOx
viSTDpKbk+IO7V3r5W3reeHU+8lXP+c8JT8vbSU0VYLtW+PQdpyYq8mRrOY2Z9pQ
RtU3usF4MLNAyAkkglrte+I0ghaZtR1tZkrU4WZP4/jJhiz/+xxtQw9b54NqgQ7N
IpJwqu8buEQqHlWobHPvJmseksErKk9ql3EmeKIFuwfaXYNbSyh/zyboGce+RmjO
ZRsKvqz2ofjQr1CRaU/TJEgFxmnwzh/g1eVRxOuTboNKc2YNMqQs6IjKYT5RhUCQ
OS+eSeAZKCaVoLxmUedDUyL2gwwcTfPXECEBpHRr8IG2dOVTlhgmM2lvguW6dC9v
7Tj2AX1O48CwQnNPQ1xZlGe8AXr6v7XHko0teLqjTWp0fkOO7v2J+ittnG2HHcEr
YciLTn6W7hbI96tFGSsl8H+XllKKPJ8n9ZmeV+0aWtmYKLHjT4oEvTmrScJGxVbh
Oikrfll3VOUJa0CXYV63+TRFP9/YxFBPk0D8fGSlEFPK95HTdSTvw3JLQWnleF+N
qTK+u/siB/c61hKE75MhbyuOyfzJWo3XE0Bsj251UVvqB//QAmQirWM2F5uNM0h6
dNl2FxMpCgJrJ9Lbq/dXu3m7c4f0eSxdE1aG6NZ5M37ycDok0ib9iDd0/1Jc4eMd
MSuhRUeu8fLUFl5F9n7u9zAt7Xz1isWzIrA2NgHyiUKU3I8Nt4ffJR9CPdAZubtS
T7APLU4JVhCYxjWqDshdbkuh0BrSleVPJIwF67Xa416ENZFfIVJ33uXTbz541nC3
mFAVZMHTX0eO7nWlqN38OmX0A65fPM4+zr4xZMt5cJSU3wc/MrsuyX5iOMW0JPG0
zC918BzRGbmBG5DH7ySld7n9tPgNqMwjG8AR+sIj2BiyXXC6fnJ+albnhrMEXacE
+DowmhfIU7oCHnOIyl3MthiCuTbXugMnR6E8G6Lc3a0TfCH4Z5Niokqeu+HxnVUu
VSZ9b6h3FQ4wvDrhzUZ4yAysGRtRNOkxMum8CswUUoXJheCiv9P0tlIBMHuE7zyN
k9ScOOMkEjwqQcrXsO7Ry1vbS7jeX/mEzUUpqjAHHX+6icZUvr45hGPjvdLEKvaD
nY7TfqhjxguVg9fM4sr38NqBS0ajr09VuI+25dEbTiZSw2aKtpwUyzf4fUffsDeA
sOLy5vie5ytBa4mGjukUkKNC0E0OmnkC0DifBHjS3XeIjxojG3IbiGU7f9nTHLIK
Ea2jyfelCLjzT/R1XcdxsR0oQcyLCLxvQRxh+/tZIMU5r+YHGW+E5yzLEovGYdnW
Xfol6ONWzmbU84bv5cG0p0n6MB+mK/DFpA4UiMQevmDRG7zSM/EIZgpM3N03tFwZ
/BZc+dUK8SgiHXRcebXSLU3I6ZrZtRcMN66GG3X3s+qgEN+Y8R5SgdKXD64TT91x
7KAPtZEDfj0gKH/9JtWgBuH0n7ovm/udGQlVpMW9QtMR3oMMtRY0uC6oqeJTKNDg
+BUabQJNwD7z1Zj+3JsW/zlAMbdMEPGsSv2EdT2WETXCZPFH04QQynWegjVNxdeB
y2g/CPQswEi+XiSU6H6zrrzRkECGADD8VZBoTb3ctyj4yveCxL3r74VY1Sitmr2X
9EfDef2bXDfGV9dTS3IjR2GBUz8ZnfAl6l7LgBxq8R1lyB6FQJp2a7r8uLi5Ctzj
TmyG9fFw1aYeW/GeGUYW72oiikPJC+gcvPAjWTmtIvwPv//QQ4pcUqwhSCGB1uGC
CE2q0IAZeSmdRFdD3fmqe+XvMhUCaGCsUKiNjUpx8FGDW3UMwR0rR3lKF3yamLip
LpzIILbRBAbRl6Dgu3zAstoqRaHmKYFBCoieSWh8P/iY/1r2LYNegoTgaDm8q1xf
gRLkrE2WM0dD+aLeEBNFzRRHrCJx+6nqtPU9cLpnqaeUkUshXWVpRwQmCdg9WnZl
vjWVNVMkjvuUIYri7PQJaZKtUj+RFynIlwItelaYQ5sxWmo/br/s6rft4jliEY5G
5XcEhTUM62sIyDIspIpXoYEKhcMyxMW2m3GdyMHsGO9ngC1ma0ZlY1g3x1zrX/+8
QiOGR7ecJeqM6WLr3Aa3rlxtzeqEqk4zmMCd0zakBA1/knYd9VxGCoYTXD/rfKTi
HwJYySHQIcJ3WeXFL2bzEQO7e8aFd7On2vx/N8URtEgWp9b7cCp1m1j+dTHSKc6R
p57cxvfFkqr2rYCQQtEBYqq/OUjy/MAAmpZfHtiELT3x+ZQ4YqknRhYLRyguowut
OJ4Q3ZkDHf0Mifwczxln/04IYWBVTrc6DjPouhVSkYDVZ3rSq7Oy1OblPgv/KCEe
3yEst6SmMJHeLP7NLN17EMBwFIuXz/Rn/K3dHooMsR5PD2scrmjqDWTUQx2eSHBh
+uHUy2pM7VltheujM0wdIXD2mf7oT760MPdKLwg+NN8FGjwkQTF/PvwI+UlKeA4N
Taay6mPHb97xbLLQaRwCBiHZS95OzXpXhG8tN/bmnn86qWXBEqi8Q8333yf5q2+v
03URQzBrDw4geB2jkspatb4FgGLa28rdeXlbocWChiELQ12Exd5S34d6Kb+n6RoP
9ezQCnY1NANGIuaNDbjgA9qwhGcBPhUET3sD8zxWaK2DZD4dJyGQzZHXSjyb3cft
7qqvqGyspECYXadCZp5DDzWJyapTQViyy6eFZpsh6auuSiGGuEOb5XrqRTIOrGp6
pNBMaW2MUD9jCK4qLBmrCk1nuBmmv5FpeHg2Zl1ukA6QdXdFxvusL+vYejx/zrRj
7NodhGaG7NTCLnqKA3vOhfRrbSAdI2ks/OI4jJskXVIKWjhOHWsGofq3MYh4sfo0
dkNsxMvoga5pTuKKTaXZOWiUfiRDyJiJIKTilVJi3NoEzITkbpmYNUxykAiv72/o
7CWbbZSQPWNAcrx1BXCvYlx9jM/hDwUkLo0IK7EoMwjgbov2kYOjScCYs/fyS7iU
baEFH/tKXVVcYUh9FpApuG19TObye9RKF3bsZrTCbgAjlagb0ZDojvEOZJ8I91DD
zh1PSiIipFQhqcvKJZQDUQkARn4yucCrpxcER5RvrJqKA6WItf4lfZQD00ljnjAi
vI1k3O3OvfyJW/00zkelt5TdEfsZXLdFHXrLiAyPSgx1KBTpjj41HoMHvAXC7UKX
Vw2Nqc4luVUEUg0br46cIOekn3OsabqVn9e7jaHj7AUk58D7DahF0EJZOCnUmD/O
oqBGI3Wnhl2sSGgw9t/v47ZeokHjqoSyFxJDn5H+tA+oChM+c7xznYc4omhMsnVY
ZFcG7NrAPo824l5Y7mfhW9Aa5OVIE6csIpyxe8ZYz83Wih+iwa/Tld/uEXDkptoI
szO7Km1JXQ4Yd9JK3M4BpNugRPrXw8y60LkkXu7mbVvBdsfGP84uCpoa7l+htRXf
FGabUTFXzB/38ll3mFpg/i+hG791WLc1N2rzp69Ggn+wUrTBhTSEGwTfP3GBtTvV
1uk6FRUmW1X71/QoShRNyaLnW7AEPbwLx3e4k936UmQlZtpJVTg6Zbur+fCqXDdg
r8hr6S+mCKxjJpmv9yB5uIm1VXZSTYyVlPebGhUodLnMu050L41bqSziHYXYp/xS
bgq+h9nOaeegu0oqR3FWg693AIpTzThODJ9lrXwOicyftP4ObqT9ouUg31sw+FZu
d89sxkhKdKFnYCRQTgmw8EWp90dlLr8cM6bJFTzW/0zQWYrNseCi7JUIh3dn32LR
c7SbUwOGXShmFv39lRBb7C7O25x3NdjD3snGebzbPnLN8MDlmNzQDFuE9sV0GP1Q
5xHh146hPZJPOzAZksj8UZ+J7OQ6b84SnPtXw/muJ8EvgV0dfzqWIkwwvB0xBImu
MpTOTnFzx13IBI3KJWOJh9IlPzA0H7T+fui9eBXEKrfuobmeIs2NB8fp3Wo+0fAC
O6HPRujIuiDqujaw2QK2m36rXYByZVVufyQ6EQvQGpKBUjfBW5xcC77+nnHsW+BY
3Y0Ro83V3pwV3yMq9BW1wtWwSVd6OhK008UHx+GBqGsQ6DsdruIKOFyQihQMoaMl
H0kJPPxJx40Ll4Yeqg/FCPOo+gxZXLP5hAtsPnCTeFUDffC4E/n8zgtDvsupKTXx
iW+z3adu8JLEnXXCN1KGNi7Dj9oTvaDkmxINmHdnanQKOty9f0C/H3lcmFEyxlVN
r73ivHLt5knv+thZ2rs87pUMLHhG46lERlnd5ioPfSbPilyvW9BhS+CsmbKCDgzX
y6qc9yTNzoiEtLsZ1CUJk7BGscTbc3uvyK4pgPZxzKxX0ap9EYXsfD0mcI7nLCXz
9ndGHQKV6YYxs8SGSZ7qTXFKWE4wgdMdM7WVPLO1EjBU3Yu5JrZS7MY7wVvO8OkU
QBAkOJZ+/W93L1ctBOJMc0AQV4wNkFMAg+zlbIljsDPcHgosXL7SAc1NjPhR1wFN
Nz2OIrTcDU7cCJM03xXuWPRkyTuDkcsz1XCsLBezjrhtm42yvKjh5Nx+MgGsFkPN
70LfGzwyNgjKjbTD33MOYlVZ86C8Qx6fZ7U3CcfbJUeY8MmSMaU5jbSBtzm6o6RZ
HxbRUbVuqX00VnHoGBooh0/cRJYZtm/NlC2WQ9dIH9oAFacA22sf7rX96mkoofxJ
GxtN0x48k9R/doBqESf41ZMKVuOggStjahkikutvkRqdu1n8Cqt/cY/psohGAsb4
tTjNHgoXXXNi7D5SQa5i7gjiSp9Qj2W0ezOwOrkXjFJVmnI2aBXDVfeAfgwx2Xp9
bc8Z37ZoIMdkgYEYLAlV446bmHBL2tzKXI9mJB2lHT6+OPBxtvuBUA8jzjZBJnlr
w1u6xNLJ6/NLg8IrrNdnv76F7wABYLn4ieRT0zPiCIBBh5bwH05zIfXAYz22Fua0
s707i6VMreAIDow7LCIeLsrgjnPndMFsOZKLkElPXwQhVaPHBopif3tgWB4VTV97
IooPWXNydsbLNz1Di6/Wx+zWLNY75hVXhUFBsO6EaHJeYVJukAtQVJGKkowDZMc1
rpr3amrWWz8HtR5OJ0P54UrmvAoXkdewL7BXwz4dP1V6abbDunEzQokhQmqtov9e
KWnpdefYE/TUMZVkPQj/b7H9UIphnBFl6F97Tl6+UDYiqh5T1BjuIlkcKOKDRWT8
aWVS3a1v7hx7+U1WNND2534XacEGUkEniq+rv/YhzS6X0EfTpWlPJHBqLAW+1RDV
jHK/y+8CAyeAThQgi/k4jB4dzEDsEP+j+PD0Xtjsg2UIZk3G5j+a+6L3fbmtxLAf
nTZfHMq0kYiV5A0WUSztJBmREbrOzgNDUT+HCtbKd5GCb5Qu5RZ6hweE4mI+nXet
F+yyzR47CIrbNsxoQ240C65xqNTkabNuAga1GwzPFx3xMDCXHCTRPgevORJmXEf1
Jxrv1+iSOz6o9L6CTbDqAUR4/VboWq1dayJ/fD0XUO5Mny44ksyHWqnVbcBha41z
VDtR9KsQ1lJvv+MtNnxdaiaAjdpaAtkAeQmtyn1fbbmkfLlV7Ew9i3FKpmZ2htPe
S/vL2pguY6Rh6SufJ5peVanBubH32al1iEdDDAlY9f5ChUo9lT45MLJZNV0oWIkb
S12s7ivx5q01SkClfIyvONQirLX1rVmVIoxPEstZlztBLAViwcQIzxtGFPJ+41Ka
oN8KUAaVoC1o4lqfstyeMfnCaGi8AdX6tmCyCkPoWBg8zQjEzMs1IrbPXNcQpYvO
73AgBWv0/syRCZsZYTaQwxF61eyQJ57nk5sOeK6qNmp0UGrh0P5O6Fuw6TuserdH
/PT/sk9/bcyXuz6FGs8Id1zDTliATOu9JV0F4649HPma2i5gSb4FvbwY28uBbCaX
VriWRgKf7dvHiyMh+ewoxiuGWU9U5cX7m8x2RUxtfaYfABQQouPdvOZHly5OXQ8P
H7CJxvhSoPxnFpB3A500KuJCBlemkUEdqH6DzuHjUvahfqZtSEhV6rxDN8buFU+l
jSvgrAsSJFNOOmsCfinbXqfOSDAAjUUfH5n0Sr+0SejvEEMcLpH8SFDq3ifY0bL2
CTnrDNSd1IGW8zo0zGBwurEp/ttpEd8q+bbt6WUtlNnWlrO9/QOURoQjAikQxSd7
IF8Mb3n7HJ4DQYjQw48rr16YRrZEqxDrHYsCn8wYgoW1rixrbAbEe31cTob+GVZU
ELT/96Mz3qw/0RFhVc9AgX5bWA6yNCMeHNiQyB4xwi4Af5JS3hmOFX0Ovfn0zeaP
6Xs/S6L47UU0OcPjspbc7xKHGMflhwjjdIj9bHU8t1mZOGJGxc79rzHXBD9fRckh
CeinxS6bVP8LAPnb8hMl/lIcYF0EQrKD0GNcRqKTgcQiPikC/6FgNkxevLL0xSqR
a7iNYxEu3C1P7JsrIRGcLWKI+ufU2fFno0X67nFw6hA7O5wLyHLLL2VYR7zUVFiG
3vDUSMZoD94j4wikfH2+TLslEzhMWojoveKjaiivph5rmWpf2AzNDTj8kQNZZQSw
EDuGQBdpZL9b/GQTcxYsuUKyy64wT/GOIN/sFyx9g8GBu4wwQQdyCifwor0TNCdK
3ATuDKtbUZGL+waURgdziuliOnHCCgMD7OpqoiT5KbWolaw51yp+sGeAtj3wxFpf
xgspuojcF4aCmoyffct2h0Q8jG1O/fwpVrh0SD/MjPOPcV4QThDCgQ4T9i/we0kX
8NdfwNR2VST8GmDxsCI+a9DsrGkTqT7LlIigaZM+jTmuBJJPeSOBiCAECOCAUJ8R
CyC9LyEGR0Nh86yjc77k+PvTIuF7Z1fFWpkIgv5ggQh6FZLPBywJtm1wlMaJevCq
s4wwC/8Zz/tRKiIk5lTVhBVfWLx+dCyfEGhLivF/GndcOfgPwLF/mqwuj2Vf3AZ5
yOxKgMY3mYrq6qAQ051XWpqCUkh/gKJqPwFfuKwnQkYsfJONP4LTAqKKgXJapycD
V9WaNydsNV9+4QGU3N9W3KFUIK3aezrQ0KiJtPAxvQzKqFTnJJKUecEP8xtBdB/B
/kKx2Ekt6sBQ/FVFimB41LYlMeNtX6kHdYkb3EItELi25sBDRgPWcYOwMN3MKxWO
S7ZtpETJ+bTB8fr+r47Ccvl2hQs6WU/TDXmzLG5Qt6rbS0El9uQxEmjRHYf6IwpM
nkx66DtzWI0Loj2Dop7X/texVp32YGLaaOpGhP2TIJ3L5wu9sD5M+5zaLbN0PB/I
9RjDNbJHw0LOFEidfi/A4fGympwmpk713+NCiXJaq2XzVNaYqgi40gnZDxuRA4Tl
mHBzEXjBxIefMJULDnsu//WqVk2PFonkXh6A/3cmDra/ZEx+AoekbZGeidABD+OW
VNGR9u++aix7DUhq5XCoYEI4mBbmvJZSUgupOwYlqJ2pLv5HOhquNk6WtMujqSzh
Ekdcky4FWFZIrIRsmOVU5oBzDjD+rFW1ZHsyNkowaGAM8kSo/wxFPunnoANaymCt
L/V5mdrMpEdk4WLTFxgF26+YIqz7HZ7JtkgSfcoaLsRGc7o3nqlUfvR9OseI6kNm
OqzOY2pRFjQ8KBHkJhI+gqrEKtrsEuAh8gI8y5UIYcT6uom9BDlnI0eDiMC0P1NC
b6bhCKL0wQJBQ0QlkhbSZiMBEWCfurTAc5wHlvEwgBKoOKseQwRzWgMwScy3cx8y
9kJ/uBRJAG5G/XUn2GMEmdza9418YtE9TItn2hrxSU4yIp9ftGX5bljA/gqsRINx
KyPoaI2wEWazP2JDMRePntxXiApAR7+Rj7bjQNwnRR780vYdhYGHUbkAZ1PQXq6g
ZJ6v8+7b3AeJBHaQC5OmAVMfmp776MKEi3Zm1JhcUbzI9ggIAwlj6XMCYEnc5fld
t1z2dkgTD1AaM4ppwfAvmO8dxMv0k47PCpoQAhzc525o5/2Ko7eiJgWsLaVRS8xR
/mlk5adx/TtJbN+GcpU+aO3mt9dHL5EdO8AIQYpNt+ZyATWbuo2T/s/pw7GjkDO+
xJV0k4Kl90WBDaXf/ujOlP9YaqT0kjpzn/WKk9M1Ih0hdkIVffwhhlyAWH5+D7MN
wZQB36Gvtc/PV9WeVB9Xu/6G5yK/4DmqsHrRY7wyGc6Lgl+gORU9shJcS8WgED9y
Is+6egHb3xiG2oYrMa3x7JZsAk1Wx4dEOCpLLI1IK0TLtUXEIp71tOpGsXd2B5Cg
iKZ50wg/foyxWEICvUhzDMRfgC65UW5zOgn3Ao9z3CUb9UrOFLIIcnuv9nrmVkrY
u1d/rVVFWUjhQ50CqdamGnIbj1FcIHy+u94KHxu9y3dV7LoYAQe+47ioIV74Hgde
Esy1mJ0o+awrJldQefr3BCcjKzC2o/IXl+Ip9MhxBPBzpgv7VhOfLVayGjmYuNmv
gdg24X5Mbw8/2wm8yqJHYGrZ7doy3+EUVf35pO3WGD+sZpqUUDqc34c7zhQRAob2
xL+L2OewfxX+mWP0gDrb8WkC06Dw/2v4ZweGC0EvlwvJ5gkNHDxQhuq95mUaWy6L
vl6hM5/wXFcOm6xWwg0Fd5DHppF5b2htEcOBq9vzWDCh/yqI8MTwi9g+hcy+RSSV
NayajqF/aWvBFuwqMXuY0Dsxb0UsyHvalYf+i/AWMakME8HTCtlXf79wCq36n3Ov
VyO+x/HmC0EMkv5ifG7HdPXrQs5T8HZzz9I1UyCP0P+X+hO418WQtahij/nsQqOE
wGBwRi0DGEsTnMeLFSRddEWGAigUFV+0us0rAzVxwz5Lv53zRnEhfXOic3zRrH3L
wvBahNgAiz8UXpN6VoPvxARLqUoNPi8jd2t93ud5I8l3uzVad54hX9rfYhKO6OoU
ssU/M60ouoNGcyBvF7OcYCGrUcv1TQE7gkGCpLLKdqm06Kxo5JI+wMlxwf1HWed4
XV8d2BU/Xgo9r7/FrYRltyo2JWac/oAK0+5R9sdC511bQ7L6evSdS2agFdwkVmrv
45Y+i6qsaCTTFo+dDYc52lYKzfPOrBwmhb8g7GZsSFOluonSbraFiIFf2VUbO9q2
VVhVfRYxncFxMF1NYq4gB8LluR6jZ3e5RmrrybY4iY9UyN1G2wNUVCJbaW416E+t
PXkLEcApWoAhpelQWzJcyGeP9BurmpiMqeJttdrXVl5XvK6xY/AeKxR6ISI0Wm7Y
LfOoWA+VxY93O/wXUVxNUhzinTAw7uL1/TFY9gIm/k1gPEKd6PYTQKsj6sTmytgY
YcPlfhc/CUxl9lVR5jzsrVzrK5xu9QuR+MSzJ1uTKMrGC2na29wcQnjZ/t46Pbtw
AtGZTHx+gOVU80yIJLnpAzYhlUWJlXVJKcapNcZexb2SkV0U17AZf+uf0ArCSamv
5z1yDwStFV1GhadvDF52dXSJCItIEjmKk7EW2bAuAcwDWg0Sqc6+0KczXgEPI1Pb
3LlGvFeLIMdwYmu1Y8Ji5pHRbmFeDZkFBrgNtfK1hOP93V0LBFbTMyr+VUeXbMV6
jcznM1y8NTswuNMgSc0OlLqlUHQ274QwClXrOttGKSIoKnq+CiG0MX1QJV9qfYll
YDoV+M9yGM2lRmZdFbIHJsrztCsxEPDUKnWBwdBt89fpfD/lH70T5GwGS68WLjXt
/qJND8mhBxORUfIMx01TrJ+Kui59TskWjVR36P3/FOsHH/4oaOkpIFjlCcC0nS7U
E+Yn6Gi4nrCfgOo8om0oZjaSu2OmRDDPM00OMX7Xzq6R95JTlejSSrbZvPd+AJWO
lwCHVLNvVM5VoTB9ha8lQkcwD8jt1sK6VBbuiIIScpLzj3J0xdJsj+/1GUIth1NZ
abLlzOLu2z47LOceFnEHyIiIMNVyGTgwVWsCsBUiPYCJ/1TSaDWptgPVp//SzzaY
NmwBIMGyc1C4qhA5hckZu86w8yVoFC87FwYyNn7y/rZ2oOMvgkPg+I0wfPWHpoQ0
hxnzCfLGYad5ec9A+qmnXJwRsGuUJpIBBRaU8CgN+A9Yny1MdvcOni5v/2mY+C23
JRtPnVLmPtUSm77ZRY450zbtLrSXzquA+rgoHKL1mK9g5NbqlkEC77YNJvxA/VMH
UIITxwXPVAH7adwyiMIGg8XY+S1knikhjXSgdNQjJax1l0nIk7YeLjEAidbSotZy
33Kbnr9WcA5tmirAUAvmxLQZxJevvkRd0O8dRpcVNA0kp5J0Y6lebS41aInItya5
cBhLHOvxxlMilocinP/miZGF+kyGpT83AHxfVfg1wqPjDAEgSbAJn7gbA2/nyQPp
WOvt/BKFF3phG+PXosIRzptsCQ1XUVm/vKK9p2IUaleCaYU2a8W4UbaC43DbPkiV
L8FOh4v9bWKUaPdgebM+j23QaEL/W/ee5NjAhms0WE0OD3cDG9wMB+y/i99IDLFW
fsa5XcerNENQrvMcz2iGCObFRL9z3lVdiE966BidewWS+WY/0S9gd6O+Fbc+ZZaS
UqGM0gx/uYN2XqWkDoJ2axyfd84anOBr0yycYTqXhx4jg9ie5RspxW9cq/wIzxHZ
jirGM5QCh1/8adi/pbLQn2FOEa43ZrQiZJg4wJBt1l63KGBIN/HGgsPcCHfFNNoT
FtbFHUp4QpQG04Qkjy82KFQZwznNQC0hudiBLkXZ5LU1/NYKFhuUptvH5uQxmX6X
TR2yC9D5wno53jafIcJkko7rTfEqQTCj2mEKZuv9l/vY9REuxyWX/H0NsHfUCCdH
uuNgPG8Iu+PUxNnn3JxyZO/tSTlZj0lYgSTrSx93b7knyu5E0VlYA3T27+H1dCBJ
rFeqchgNhQ899O77P7bHUy4+xpgZdm9j+VatNHuupJ5BZ6zf8eaG6SDhLsZOjB/V
tU7GqOlcARiZZCDjDnNkSVrAgkMMMT90au/oXTaH2I3zN67U1UehdETm64xzpjej
KqwlPPgGjEk0OIDvuGHaeNezbqv0CDL+xlEo5qNBuqDCD3nhwZVVGB+syur1xwZ7
qq/2nn2ih4TUfEqxR1XxkWDuP5z24u5mLSJf3bHCjkYKNLckCZsNoTTngjWaB2qs
6VvXmNPHQc2MeVIRffxnMZ/y/4bTSiJmKJjaYwNyiIwJZrYSQbWFs+JVTkGDgGP2
XuR9QwcTEIHzA9Cv5yjwZcatZ700qVQDo4yOpA0qP/+wewY2JTNzvACpTmf52rWV
c4udqKywmvNQlwC051RgRJgeZyFER7bVRFFFIYYISLAKmRJYQ9bJYJy2Qj1J+V5C
c9dcjRE81cFRjsWKb5aLHQagi8pR9M7+oYCTY/u4h2oOV6GgrhnIwaDpqjln6F+T
1xB2FsrbTMHA5lMHSA6EGHaNATm6nIEFeOIOaG6NLMcIy4pwb8trPWiqKFyy77Ya
6Iig+Eus3o6J2jFzzww1bRbW1DeKA7H+I6C6kexkENxjoudrfBtCsOUg+8rwHoQW
sBRsTkpsQOb8/OeguVdukejzhs8JYgAo6DQHGaWiMxVBibeEIQgZvrKiMKexetKK
Y3BhwMOU/lrnDxnG3U9Ge0SJUrvutF1pbaoC5gOk/4DwjYKHX+A0ff6bpW7tSRky
tgtdRYsnjRhFE7DP1egdtnoLp+gvJdSvBVbW3E78gE8f5M7avTfDrTaqN2cFvlv3
P6L8jZefRGnzjw4smaBqzFjIoKHGTjsfnVGx9EJyvplG0rnlT2QLuU5ewQmABw6L
XBkKyqpeYrMYuehsJ417WU/U+oSZRGJnSCP37rNUq6UysbwT9il0OwnoReYkYo9+
tpb44LWhZbt4eJ2RldNg2Q74FwX2O4H+A0mwhL9GOn/clzquVb2ORjQIqEJ0BqN9
9J6z0ykg7SBh7TezzORD9KPKKARa4HIu4LPVZ+sqET1tKhRO+tqv8sREQfDRyUT+
xPrOSDdQj9GBtvMUEmH1P2thBV1/nt7TKeJ3OkYQF4aJbI8FLzIk4qTvQKnQ1wwk
7L/mEb1xeZp0TaBHeOqZI2alTFh2MXPP89n+PGTT7ImkGuo1qp9zIdX1VaZEoXa1
PlMA1qnQ+wMr4yl505Uh+p3OFOjhIYf3pwcn0JDQoHETlOACBYmBnAyMKi4TT09S
ycLMtYN3PcYgu6oCNBTs0cm9RYAp8JhJY5Q3TDIPiWfB+/QFJEB8xkxp85WsmSPH
FCwwsEhAtlDRMvKqd83AfpgamA49IgxPUIawbEQugbW5/chXJOuRaYgAtSizfFg3
MUgvJVw69DADJCjmlDwpCI2Q3FKubt23QScEq/S6o3ub8D2USDI9RcvCvg0MWcz8
3a7SqM1XbrQFRftgBsYTNjdGtonfRSLdSrumJdCDyvR0pbC8/m3Bc9CVDjE2lDUV
RbfTWGTiDaFtRtUWODQO1fbG6AOA6J6rSE5nVMoJRE3fGNjPwylGzyKVt9ezPo9V
IdkXeqTY7chiC6wmTcW9YU0qiwtwMnOzIZ7l16IkmZHNLFYSR3KmhyvieVaXDhP8
VTgOrWG6hJMaivl13183Jonha9QwjFqJjToiDTF9r3L/WPK6rsh6Bl06UwAxJa84
wPpdcB/J8ByCOSLaL86TGzcoJziIWVJYWVg+XrDrbSGBAyuSYP9hXvTyMq5vAZAS
GB2vCBlg3/zVj9RR/i8y6i4lmvUYsGKgg8dJJNp26tVqHXfRyovXyaih7r3UI9ra
celKtVUZJj8a4rbVLY4oLaTY17QQQl+nTsJzCMFCPNnrWmTDxVujfc6jinlmOQj1
8tKHQS6M/XOdb0OO21Lr3YTpV+/Qef2Y3ziMQjxmzCd3oMm0/aLfOrL2bzDMq0wY
XIfEL88DM3h6926F70uzRpECJE+6z60Ku/uqlE4WzOy9zYysUgclaWldAgPJ0eBh
PLnkvVQM37u8FjgVHGIPaWdmqcnqZ2PIAw5tcvFDyzpkJmARHvXT4LRHzqOTexnY
+Vd8ZpjzQlRh1nKBWQoPTsfjvCTkr7miXlaLBqKx6UaJI9N9BTWzI7FLuEKKnNZf
FZyQczDyetKW7cEroArjNe/Cjg+EDYAIgrEoyzVpzXR6huDpXjDksMuOUXMwVwJ1
zCp9K5qjG8Uiz47D7veABvdow0YS0X+M9bxGGFKRx/fzKk0iSiu2nborQqbAN34/
ocgH5afFFTykkdjeG4CqwTYBk7USaLBmS8tbLoW8GG/M0duLtmLRr3LKDGLR8u3C
oH3rrKhdzOJr52T8GTqvNR/ycvwhmaZEkspOE8qlwh4Ex0PGWqg8kFePvzcxyVM3
75SCTmvuwChwkrdzFJJ4Et6C18Y7BH71E/2134G2fMPuVqNOCdFC3BkmOV8nKHt9
p1Qa2NeCHZ9V3Bwz9Ls/jU8vIzG1P11ja7j983Y5Ej7kphN5NMUHp3dOIacCBeJX
3zNdMVgEtLX6MtNfbdkebS1NFw41NzkrQZBZqsb+YtcByA/+imkmXFpxFpvj5L4e
0YfM+DnafByhcgu1uq9Gi7dxF34kz+KY6LXC1zRjz0xYKhUS45HfaZjg2q3B1iXy
GE14py6STv580WiLkuhOVtDvrFRud2auDXXG7U1iPNZmS2x+N1OGv4NnOQkNl5Jh
WX0Y5yBbaYWW94FipQmRX040TbIDi/CbYhk4NsYM+MPsbeTjtqFEAViwlkSq6S0F
yeEmHh1du7SsOghp2T/FjHphxUu3b9HjFYeOz9+RMze7GFSjKQbazohcucHEiWWU
kn4DCJ/op7tkdUFdoWbR9rGhH/coUqElza/KQR8g2ZbylomgXg4RNSYTBlVFb7Dh
4fIOTTJWFJfi43AvnZUg60j0uOPrAEKPzk1v2sIwYo8pw/CS+aZLXVRyq4OSwVJa
wVs5zCw91XFTvfH0NG8/g9Tu2VKXsjfLZNT0Zc8zJ0JTRW5dq2ju0hjf36yBl9Dc
oG48ztc7ukjb5n0NM+HZJQWyEpKSo1HVCqCT/lkV1HQayt82Fpgvo+brP4Xf3c4P
915nhyi2LS/ULoiuTYS2vehPks1w9IgW9tNJZ8w1/NmnRTyFzX2VAZ8JhYqtKD6B
YJE/R1RGQZrxg8VVwEIXo2EZQDdVeMbRAAbnltb0uh3483xuz0ylwhZJ3k4eCYPH
GN68HenFIpL+9Jm5C8bLUg+Y4VFJC/4xV4f9VU2juEQMKNKEYXjyi3LKL3/dk4Ax
E2UHE2obAnCUYo+6bBzfByYfsNn29LkxLb46Q+rMQYek3tl+sTHKUClo+a4HcaD0
IFIFGzzGo2BSITsSaYj6ra4O6YiBZQWJ0KgmBkqvvb6yqllt39NxE26lzgKTlzOe
RI6YtDy8c0RSFVK/37Kuzr5XD16cK1UyXr4m5ocaUKO9Nkc86mRlDevuEkfW2Yd/
WPw9SriEJzW6n9zjaKj42ZrQUIXo/IxVFBdidJ19wTl/vY8Pia7p7p3PyPyW1ZLL
2H0lp2LBJudjqiQq4YNGTloGOMUTOWnebpYX0fjLwyPwueSUpY1d5Kl0L7+yZsUd
OSwbScLfh9Vwb5W7izRngnD+lZApVWt2mjrXBOswfv9LAZUUfiCbY28ecwQn4Y/W
Vz4dQWttmylCsO4Nf/MBgs+09H1dcJos8CCc8Cywg0XLzMdSVCZEI2sAd7idk9PZ
3u2AZ5GbqSh7LTGE6jGcwby+FeKuMnadCPVBla8govALsTYB8j/I0/a7zwlU1sHZ
1kndnR5nHmt0pT7I98/2dfTZhsKOBqmci+NQVtPz06YI2L17Td4hS8mXSGHuFgsz
813GX2ezdqpaYP3dqpi1vOYxEPlkSr+PjuMqPfqmkoC93E1bdPzouPUuP4CwWEBT
ZuSG/qWISkVEebFKhEdfgtX0L7HZEg9sQhtbhWxyyuE2reD8eWeS7reRBD73eamN
FguxSfRsap7PgyeLAYjveFDsK/TVQGkJvzAQTRo6owFcCLEfPMe/YSMHE8cKLRI8
ymmvvbS9tL9FiJHEQvDR/+aF1M3dQS/X3L2mPSidIk7qCuVsP+oPti+SaLa7bhp3
XsTm8xBVSf7ER3xGGpZgZ6v72cuHmk4SAwWlMEnBlGJbGBfgOz7/YMsYZ1VmX4BD
sYW1f8eMOy2z8bkETPRGN4lFf/GURwW7FYIOWHZSPfcwxlFbBHm/DLdFA42HRtMX
/7hhAu2bnhKrQVi8eikvtG02kl6f8khsoHsb5KJA1mxKbFcbrLs+/S39oqWX0nem
L3Z/USpPykKMlRfSb5xjXImHtE933Vj22AJ5ZWjNuby5XbACw7tO7Pe+MoRNMeBU
kx8hTyPoCzFiSUnbJCZi4iRu9lo2Mfrl4/4phHMLAteAauDAatMPbrzya9UCTN9o
Iw1A41f8XvJeHaxzQ+WK4ldyLFXUahTG09SreZhn6t2lFVWyQxKSpfYpMd6IrnXA
73byPxcWMPMAUhahMuzjagRW++bCBqq9hW8v51E3l/4He2MxYvevroFnj6JhLInW
+8P8Svx8RtnYK7zDf1xsAc8y9HmizO5cPA8Io6jUQ541bjtOICGeYbZrRN4R8N2n
iMy832534lOhjU6uEt618oLxWdIzEGxLLvLGsWifuDFmlVnqBCfiLWhB5D1vfp4d
+cv14ENjBB3lyDgw+UsNthUSGRGiFEG/jWt9gIRI67XlvLLjwuPhilnnFKolnKnU
/4Q8gaHhMirz7WEDC5L0ZGBVuLNzais9PZX+KhSEyNyKRGsWtmEuBDkW34WixuJf
jYlJlFbUu8uoUq53sIBGz8cdns43rf6isUd3Xy9vgZYMYkvwyTtj0jcBW5Y9VxBN
6PNi8wYadS9sUnNvOkVuagXiMv4IJnBNdFDTCd5IEFk7f06pIKWQ8DmOSxYcCZLO
G65a28l66Qyhlde1ZCro4Ws/l6CDsnXtXQVucT2K6tE1nPhQF7zEc+ngQHRJ32vl
vezOhSbxIfYy5SEn7C4jIihf/+A5cu7cIpe2gxc7zs0XiPT0LyT4psQKM7E7OZMW
MuGMrweVc9Mw2NTi1KekM1kvK/xTYpCeITHlZho1KlpGqc5wsJq17ZpGm/X0XGnN
U7ut/HKU2yKyNS9Ub05rqJDO33OxPgoYTJdBnUPGrLYVZJT1MtQm9JT6hQPXYF+i
z6qV3SDiACRDXe3+7Cx4/fCrUk+tZ5F8y/fVqhDQElcXxc+yPGUpSgt9T8Cv1kFi
ek2SVK2CgehD869oM+wPE3DBbOLbD61NbrRiU0oNEZ+Ruv4QbKgzNVpeTO8BHAy1
fUWSmLOjX4OjjCy9Ew4jjHBLHO1ffEoq1W4MyMzWhaL/cEv5sAlXN6QC52+XzNRZ
gypLzQRZiil+iiJ6e1eaZ896cRggmYF5U1PiUq1p/VEsONvu3zyCx/X1pH8mUIL7
SWQqfRSJxWRRMjggjVcB0vg2QYRP84dxTvPT5LAMtCrhKkix1g5266wXYyAyX6sr
ME2RxEBucgXlhAZw/87or81E61j2Qb30XCtAJw8lu1eAgJ6/HlBMEQ4ciTRwZZp+
q1JRq+DEoePx6euo3RbT2Cm0ldV3dKXf8o2lMXrkModmuap8lQRjcLQCpI+vEf5w
VczwoE7L+ed7kTbo3pJwwkFlM33JNMZNCcynz4dz15NiWH2i6cslCHS+Lb8xshIM
wQJLIF6sjQWi6+lfGgDBDe8Nz6HTocwvuinrRnbgUSy/Eqs540vQDFNUYt+lzs2q
RTv2gMqL3dSu9EiUy8rsh772g6hDvUnRMYTHS3Zgj55FtSdfNuAv32MKxxk/t3lO
T2/HcSZIPHp4epzXvoKflQSlMAX3CHWyEYXXWBRnr7dV8CODhbzXEc1WKz/KWAmp
AthBU5ZDZx2TrOhaJtA5rCEV1rdFkNHyCIaNoxYwmirAYmX4x0C6o5VBOGrdlUE/
oFYe4KLZOFyxdlCF8Ofi9cpV+Onkgrj4P4ezrHz6S5q0byMVgJsU8FPW0lXmjCL+
2SsvqyxSusUpDcqX4tuv0jvZTIdsfh7smFojew8ib1q8+mz8IeXoamQbbIgacK3m
H5l/r8myQSemtudNnmc/0+SRWNDxSAwJrU8Owx0JbxbtO/29qjmuFyU5NsQG5D0u
s+jeS/sUWNbLoqNOi7UkdDwtjEG3iT5Ph6TjDYBNKd2rxN4E397rOvm5Jji85PVh
LTxEEV38hcLo11AfJ5PGxRblVSEnygOKLPN1PpbHMCJ9gdA1V2CJIphOHTeTo4dK
UHvmC6ViCIv4gQxDGTCPOhOKA2mGlzaY6V5npRkBT+LFT0Yjnk9kXQ8gHrXCv9nQ
lORPbNv7a/6pdsyWjl9v44OxMhbNPz91r80+IYSzV4s2MbBkY1M5s7R6XgqXZoJZ
4KPuGKc3OLFCqa04hUggqeNwSF+MPZPT0I/JvKABtnXkW3+zEhG33wkNRoyAlPO8
1l4bxFaKsWUR5DXBFhFYjzHGNGeNSJ4Fq4FYCzwYH9W2EnImMrZjrKpiuLcO8IiR
bjkuQr9kM3Opl6Uux0demzA9D525GM/PqWLYZwbjBfa3hPQg27beW+Bpw6klTNJu
fath2TStp/BEsjJTy+/XQrhrKA438/6qMm+lm8h0+xATomqSvfK3WM63bFIc2CH5
Vt5axtcm3AruurlTnzYiKeFgFuK8cs/kY4PU3mWmmZcvIL02ix1ecwiHbMUZv/TK
WIyzYo+AVFVmE/SZ3PlzwsnUvCCS4UktKnovoJU2zz/qhL8geLDLvpSVknqYtGOM
yVIBOXoSgSRckV3fRFHJvrIhSfK4Z6Z6fPxQCbRA4pW1UPaahbsr9xVE+stna1Nj
k8H3SmAP8GD2WpfkkB0DypOnsDROZgt/9qPVb1eHvJ+dSJ5iWUGbu3WpjLygrVCm
fUPwqdEzTP69398T8S14xR/f0Da1sDDAfuiicwuyHXnT8IRvGDFjk+Xn9JRVpyxW
DPpoi3/5iYWKaWiyv3ZHWfkBruku54vrjkZyuzj4jBIT2GOTayg+KLtTT2kpda0w
OeUqnfKwMp0R9cEedmE4UdAVAvuXOn8h/jo/b6WayApWZLBrnYn9MEcxXIjy4di3
I+6nKM+vo6nTTpXQs6XAwmkWlIHXMnp6d1fWLqhUdWbYy6UXi+oZC5ONKpwCU3HQ
q1E9y4guYyBdRnxQorolzBgjoPkJxFJtCoDOMB6a8G5pf4BU/Whx/6W5sROYINLl
XcF4tQcCRNbtAIYCu7zsjh81BQoPimb1GUhcZSxyXNGiUclRAXGoJJhbSIHHNBIb
r3+GQEAnhAbyoPmL1eFktElGPTFZwfQO4QToYPTNci8N5XLxOuuNIGX1ws7yHbzE
XErFe/3jFYw+sISOa1IWN09Ajul4qOa2boZraXH7On2i14eybF8jpKzuZJXQeMle
OtIYqYQWGAR0OuzD9NFn8zq2g4we5WgofLocu6EdMvamq6SBNB/IEXwm3ekLQiAE
xGAIqxv+SU5BDmbq/WvDBoZgke85rnqC80MgmoXGS73yHa/Y02pjKEdPYMMYvhOZ
uX0DtKvtyb9cwFTni+11oNXO64ka8ALUz5Qa6rBVFM/XekuYzr/kRikQs8XVuOFZ
QKxxsGhcLIz8t6h6v4b1K7UOC0br4Y6spRsCKM8ehz0odPmn95Op7oPnY+kzGMqF
qg+m9JSPcLQO35vpH7q3IYcsJOiyHhWMGKY5Lb4i4ROvtXtDNw926OsELgCVMhNi
G7akzdp/RH4oRPEN/I1J+gNnJGH/5wb7jvGSQVkhVF+MIpf4dVtUGM+/thtvN5f7
wfgWjHbmH83kq0H6Ir0tTScHnGfMLSqiJPe9dG8UJxNreOPrFlWOCW72CARVis9f
ekojzQVkpAUv86w+9hneP5wZS+ApZVCytq9PzF/GzU5hYHNRo1T5jFzfuyZhfKPX
QTmcoxq6d7DzTguBi+JkBs6wxyeXvgYb+Bvx39pyqt3fFQOnVsWibqt9q5s7cIiv
37kKFtDlA1GUIyCtHN9GdlvPDD55TXrSHcaftcbvEEmrdAQXmuXC/agZRIbvBwiJ
p7aPfKlwGLkYhUJuvYCA7EZOgUtK3MY0PadwbMdwP8Y+YFM0shb3c79mLKwA2Kyg
K8nxIayAb8iXAnzrZ5TZQ+Key303rP0XbAVHkgn7JSSSwGKI+pT1mALZX7TKajar
wj6A3y39RTcexhKrSE1ebKLIfwFljuxLz7Efvu2ZMz7uhvkkspzUvd8ssT8NfHDa
aG0+PCXLkKB++Es3OpjycYTcIIbP1QBa0bGNgHzb8fg8oA8MsTG0yCerU1AvG2WZ
XqH5TvvHIHQuE9rrK5svYzneB0x10sKIr7sgBKvVgvTHXebTcb244zcEo5AIIGdm
E/vTOUQWlAlGot6wWTGrzEcqYPi2B40Upq6PEeS4/984OP3KtQVn7oRT9v7IITea
NyVajBal/TXs7vhnDLfYj1EgOuHinukF6KXgaWMI7bmZ8LlIu7s8qzq84VLriHt5
Gvzlv6eMpzW2rBaCgEUSMTBb4pH08pJRBCnRDilCuiQw6wN3ByAaZwGTI5NYrV/H
eCQYTMlA30Ca+sUsBAZbqf7n2XZyFS/KKlLzjnKKo4l8zrdL6zCCiyNYVJ1dCQuo
699l+Wrr0F0hrS5HMey3Qr8ARRUWsjpYnTLKZnMd/9i/07PuOpA932oeqcfE1I5l
y57UazrjBY6acT9i3rBKejxGmK3Q/q14cAqE7WFe5Pc8ICgkQNJnaj2cGxUzReOo
Jnwsj+umE4VTY2zcun9vcb7+T8YSAtjgBloKqxSz3h2pA5AQFA2bcYr4d1jv23LC
jE3f0lAcJ3JjBSWiLGnbXYj8SR9JSOXUrcE/PC4Y+ILx76coNFY2brPeJej/9HyF
oBHSK4HnMAOefU34y8GBmZEgnrOCa4a6uAHpnhcBOLzYOKF23vcCjFaqB2atKVny
sKi8wkNFsvqiR6MaAJghLABIvzgy6VPIocxoChlG1/wrn861XFEX/2F9qHlgMpNt
596vugh1z5GATscqKSGitXRmi1Co4x06lqDLirfsCRl3sdagsP15Hegn6ZF+IIVp
fdx8MEYmdp92MPg9x7Kte78jkZmlYx6jNqcNSUYtz7cppTiSRimal00KJyp+M3MO
fKkpG4Ng00I4jhBvv4TFiEJPuAhow1HwVpJ00FY4WVYyvRKiQiCTZ4M6CkCW7vjG
+TY2IECAXHZtI5AYnb2nkBn0HwTZohbgci+UgjyTJzRurORSHAI64AZQKZf9+0gs
KyE5QrXd8Q+UmiA6L/tGWP09zOXpcLaUfUiPlYjDqnlCru6VSJtsidBcaMOkbPZL
C+zz8B+2c87ssHEG0t2obO41Fz7o6bS9v8gr/Pi/xpmGXKuqYwjVp9EkRsrwMO/V
aT27st7BRdRwawcMZmcgbim2ZYHdRX3uo773zB5z9qP/CQ/POQBwlESdEvmtbetQ
0oB4O5USRUMd2cg+NUmML3/dG0ZMVWCgy8SQlT1EQl3Ir9k6hLbMPLtk7VpC63l8
+YUO+OBBLIps+uo9tz/nSrfy9p2XjJqxRJVyDeLlzdhxOCtFuq57xnfPr7H90kfy
G6s5BRjM26Gz9SaC02ICQhIr2D9GIb7FhoIwuZq1nX5WZzH0/Y7rE7L1jA6hbGlA
VC4uZ88jJFVhzYUOxQjvicF/ng6TcIpI7W3Qh4cjVIodLUh0fiEwDsghpO2VdcLz
gafGN0hSkBXZfxKbw2VuDHgKnr6apNB0xGdAWjPFXylLcgJErTM6F4qlRTSGu7r5
DZx1DtUHq1EgSDbOVtv6h5sKGmU9ZeOFntNjipuTP5/2oMmdh+YBHFUr/d0QiTkq
DzprPqEriGmFqclktABCFdbBzKdxCYmLJZv/nAyCGs7TRHjiMK+rULyi6ADlGlOA
KwQxCPHZK1Sbwwk2KXjh0/dkTa2lLyqdo/tn/h+LRAAYJieAZ484+cavhBr/CPHH
rwxIdB7tdrcgiMdSVdVaX08FylLn7iu9256DPU7NNmxf7IaTmG7+JGBfXQXabLUP
KLE/OZ9QcI0t16YiAot8smGYkXzy2c3gpVtEgXo+hFDrTg4XqAHdzoa0Hw1jBX3d
8Z8Tv9pwWXLnFh51Xaiba1F78GLZ0yUYoSulKHcwj7H7i2AYmo3dqBBnK4bhf4Vs
gTREc7dPMJmN+dxcv8igV1m1guvGkNJ8Hfd/UTb2Ngli8ZIa/hYahtsSqT+Lf4Tc
VxqMtWH7O6959fxzoUVVquBO88yxs/6mzIm8qXBwUwWy/V9Tk0aEzATd0kTRmGFQ
ym6fkDHTS6RHm5QKmnkzsLY8iPx5QQsz377jmQhemshbYjWpb8OHEvcLsZAV47Or
4et2DPuHLxvi4RfKDqSPSMa8rakYKz2wAMGu0iv1WoVTuEXkYTYxi4xUfvdeMpS/
+TC2u6zjosaEDu5gMLbH6kHrvgbt/82fZkmgolsTn8kuS3ShbR14/KFDJh/x3ciz
Av1m0VSnj6oJdHLmN6JfQsk5/q2cLRiTQoM7/t0oTx3uEalDDeQPuIwKvaG/SWrj
FL+glGKRtDHgIcS0vPCnkHiFS3JBRRUqE2E8RN4aL+CK4i8X/KXw2+Lla7N+FjIK
NhXI8odpAJ8Pns4cesr5pZRkYH+UsUInW03e6ylazjx6L8HN02o9lbyKY9AXFYjR
NeHFg43cPoMELGQMARiKPNLtYMrYV5HcUOTFL85ycJ4DQaQ29rg2kiQZVEaMpdCl
8Nk9rkqx+XO31JGGF48/cdw/75+C8JPwV3DkPM8dpG/SYOjCYBf3kY9HceaUoMXR
2+GFQT3teW7u16buyo1dRBlCHp/Mp6wKoSBuDGahJN1L7wDfD2ZMJZwCWyqSoZWd
zPAxa4IBfbC+YFLV8/+Nvi15A/3c/GXhkQofDXoy9uTtru0Keq+0zEMqK/C/5vu1
jhhsD23m9MJUn5BRLblhiH6647Dbtwa5lxA+RFVc7en3PleFi4TgUMbpknh5znv8
OetyEWGfxWuw4aIwdK4fmEACb54On+R8/NL7dDX3sedUfHdPzkUH35+O06L9EO1z
PH6jaIHB3qrpEnkI65ENUmXa7vxYWmJLmhCtnwex5/bUwRabXt2eglQIQ1pM3Ule
uyR/5HPO5CE6k8HR6bC3bxd3BJjycqEi2MqGG+D9PJR+qCq7o1xMbZHfHcWtJifD
n90U6Vah3PX93gqUntmN7DpS4yUQCFipIlawyd2QWnt/PZmczlO2ygaglrn/83q/
CnHi5kUax49A46qjKs6GBP2zR6K/5bd5JI3S/fkUKAlGiniDgRkZM4MbTHTaoONi
jBVL4k62T+cx7Xv0NYGZfVi8zHHWrEF0NUnySpX9ZFJGaG8skhZBaPRY31qvq4PM
WTi4YyHHMfwoRR0d7pbSkHyV6+xV7yOL7+XgZ5d7AUCXRuj7vjcjdNqSJKYq7/a8
d4tDGK+6SbYPhatB2bTuEC9CCp6Y5VbRrlvl54x5dTjctKlO/tzlXtN4ALu4gLH7
e7nrJrluqLW0HfGhsNaPjnua2NXJG4KqOZgEU6Ky2YL5ZbhuELe4RwBHUYu3sfFK
a809g66fd0q0j3q3rNfrD0p1IyCfK69pAzCvtKxCWn+vkYlRvKRgPcyvu5ejXoHp
57JWBfVALm28Xf4nRl0SUfuejanS5Bv4SSlzvv9ZEPq24TApb3YA2ATDpwPzgKIE
gkpYy/oaFU9ZtCeLkcnv8jIEjkS2YOfymZG9djCMtoeJeP2xJMWrWxIcVIIrEv55
z8hExDns9BKWHB0PC3rRq1KGJoNKixMdo+gwyu3uaxGO3qeIt3fb6i5pht9CNTrv
8IATE1lopin1tZBMmy0RafXCFQILh8kiOj62ukcZmM9TnnSEM+R1RhfU+AJbNOI5
Edh91sx1b3gCi0w1pjNmHgN7ABV3HgDOPAB7Qh8OazB9Nu3FUN/1tmmrwkqugo3Y
d0EtzkBsIkSsdhY65ggcvemRYKrej29eAivnOes2ntNTzAQEtlQhxYTYb8KsNFwQ
08V6Ge2fLAXPRFmo7Gr8GgqGafEHa0qXHNz/Ds7BDlqe4c+B4PhqqQAszMXuYT2s
hICsMO/PUaI60PtBf9aPEKRiQ+h2xeQyuVP/Ot9pmSNdtaRfDwO1e3uAXCeoka7l
xU/LeRIo7B3sqZSrUEADTc+s0duqI0IjEo8VtnQKVqgpaQ6VulCV1FryDyqNHMrI
wS7YMJhlOrZBi4yMAgems7H4klN/8dhZeJtD1LxPkzZBjJH+AzT8LNHvxdLSJTTQ
UWxokf247+RJt+y67c5Ix69vDJZCfoie4mfa3UE/qXk6XSXP8rWY3fmgpAAqLMX8
gz5kCkNOlVyxX4vKXfV/duG0c6cIyaEseurssebl/AoIBtMWvEyb8IT4XPcAPBrP
c/q4BFv0NkTc9w9qUgVThmlsayEdCXiMr89Y6gWDg3po1ytWxHrDRCoKNf3L7raV
3Stazx3Hyf2yDjm6HsWEKeZ+GS6iquDHU+XGHLElE28rPX7ctuqdrpHDfqFvF1ck
oCfBc35FP/0ERnyixvIn8uodA8UOvqb1ykPNOh6qwng/rPVxpB5z37RxR4zNku4x
9mv65tf4NVPneupPVwGiqjKnUwU45eTEx7p250Gh0JwlF7r8ZtAk7U+ZZzNvNf9R
+dwAGVByjgvSUPwq1d2U+3WUkRbsfmCjnVy0z4H+s3zjJuDELW0e0BGpmGVD+ZT/
RFzClzszBaz7Ymx3PSxqSzmseix/f6XTFYGiGRlUJx8viP9K/sizSfY3G/kLao3S
l5Jg656aP5FoWkONjmk4/vuyy5T9a6nViajVH623PPSqFPSmULNYZA/78dniGODh
9Qb9QNCL9YviRZi6+Es87FwEAQ65avvMVf6bdbMfNx5ChJ2V87uSkQw78KwYqrY/
NH32AtJmihixBnPZtnIopVcSHgqSu/QROddEY4+iljT8ffMTHfd27ugg/Ki6ODrg
hKlvZlOtuvskF0f5HeesRXagRxxxG++oekYACuR5YyJt/epe3sX92JEMkReTJnpa
mL+JbzFS9Mduo8z0tKZ5GlyMw3S5BjzBBAPrjCFAqHKHCyH4tQXUYoTlDDSzQ9NY
tzxsIAh6IhdrTpBt1B+OO0pWrVa6M51SBwYSRNQr8bXl3iDBzSCNfwQZlVhNw3du
GfNa+RkwVQPGwKzlep/+K2auaVdbmfEaF4NrXUFrNEsE1g40DvTDVZzA5UpGRTrw
HVEIJRg9D/bWEO6jRNKmb5quxbdduuTgurBdw1QmQ8lZi3GDYNpILV4HzTIzQE0u
seFm2+1ZXOWaK267phynYEQzRSWns5WELHB29FSt+/qqj6NxkZcgFyv/3zb6NWYC
dX55kMG7xx9xwMuRVJDhKxW0i6RXMPZB4t2NIROJMb3WN/ummBUoht5GZXrFvWeA
AC4qff8mCPBRAywQghVXYQ7PgLsGZjxeqBe62ByNt4RY5f4VkQq52WUwKxiR7iBu
o7V3XhMIa9RnHmHQYzqtzT1qePbpir05PLY6NCUHrcg34Cigy8JEFmAQ6zBiaVqh
mnM4d4eynFj9a1GGTa32Mkw/wpCnjMYz4Rbjpa+KrGhwLi1CkxccfLh4KzmuFSWw
s2Ti/LqC/6tzIcKE9nbIvqVgZVtljwbXcWqDNQZb1aVKt+t0T2GZHMW6cxkTv+vw
6N0Ol7JRMI9KvAguTVwBM2+0n+PhWaQ+fmApL38LVUTS4M6jfY6uMhS9kLHm86ny
ysmqAARuk/deTGn5FUOhhDHmIrot+xbrtbtTogOrMLSDQLxeKIV9x0b7utI2eJa+
wxtrGgbwGt5PecOqx+IG/qN+h5pg74E3QkJ50EIlyWX+F3pcmVPyeSG+82ZBR/eS
Pi+LZfOBq3EhFPQCH7JnToTSPK8sw3OX4u0Q0dHWEvQ1SRV6J8YIM//n0R942HfK
P6NhbLZuB3owkr0QugMwLJU2cfnjfHeGBTfdZdnoxMSlOYfU2ZEfddW7G8tY1VzV
4IVxpI8KZG5EnQj1p0kZl9lp6yY4/WyeO3gPW3jTqyW89pOk+xqt1YJjoiXd9bGT
3CN3RNuIgK8TxvuKYt1U0Xy9GZJEYu01lBFChK2ccYUbyEAEPF0ptex1GgvLQwnH
vdZbtGJgZSmW9sn4F01EQPdmadeR/1Mz+yVFfp4i3OGmS51G8zf5+LpvKyOvqE6V
eVMT7aR4EPL7ZUyHZBzr3KPXqtjE+jHPAM9M6sY+19lKNzekHVTqE3653H1dRBlk
B7FWGi6Cpx24wM14UH9H4mIzUFsfL8WwIcLa7eYN9gEGzTiakzV48CmswOL68ZYO
+zvsVaMl1xLuo63HqZAGy84Bsd/jmTug999iZcm+UydoEywp/cjHqyMDCfJPDx2C
NknoQKjiDRlfLZnlOYqjxS47cffFEn68+qSe4nrVjRXy1MXUN7dUqnxDDeewXvBH
NBXPcZMM/VDaMNSJ1FNxmNgLLD0MQm0xUQcgL1VEmG0s/P8KUu7XpiH3UX5IKS0k
mxUy8IBv76YFxJuXDriJK2EKpuJYOK6YqtwBW2ONppY9pyFpEy4kvzKpP8eDyHUn
cSXdIFdosZEMNt1OvPaXH+mujzzkVwvQy55pC+mpVU0cKwWs9bJxFKY1LeUh/jLk
2OWXh+q3csHUBowVjwG4g3y0bnbLaJ11VaOoJG4W+DHYRGgQ3fQ9Nv9A2IeTuAVJ
j/IUpVkBQ3+P/riNGcfTZf+jnFvM0KbqTGJD1EwzRpyCiOaTvh+ExmYdBoWE5dmL
7wccEe4Z6REPC+8T3exLits4KMSOkoRXg5MAkC0nsFWHyvQR3q733RIN/ij8P2L9
h0QqaFzeJaN+8CaXYMOgZC6s7Ol8Ygs7e5NTx2RsJcN2204aM9AJV0G9LpaEMHVQ
Y51sLsjH3uUMuDk9oMjNjTXZ60wI9nannmtPtX2vmdPpRbBjYLBN7J6YhyBYm1vz
V94u3yg0k4iKB/qvkcr6u7LsYotn62WOAwvIyeUIJQGzQXDm9eza5q2kydxgoDOp
wxNzbAHBT254+JLZoUO0p/WFsmxWXdVLW8v2dpUhhD11OuQiz7DzE82l/bYbe1l5
G0RFcs/+f3u8Gyyi1GCQ9ZbW2hcf0g2QhuAxoi7fN4NNNV8u1eEK5ThcAWTfnq2q
viqqjCH9nQVqMVm7nbik5QXUsX6ATp2nZCJ8jgAT08R11tC0RPCHaCbf+YkPRMLV
OVvh8QF1NsaD0I4AaoDRQItht4p4JEu4+yqn+9gQ003MGww86WourglgRwiAvLiH
OxPxJ5042g79Z2lFYmBzAPx3Iv/j0a8V4OqxE/vSQQySTun0DZAiVtcVS+gtptki
L3m62GqyLAEkVX31Md23ku0FeXj09ByL/JHKCq4Llpj94H/cPiCfUC9lx+OzSelI
z5nas3oS/9ZOZ8bClkzcmDoYheUxayUw25AvYLANskcXMa3TpAZt1srfVyCHLLth
YxOK/QvUtmhS3LXgDCuK4Ds1v16bWhTTm76LJ5QdYmFQWMfNP7S+kJybcmxFjkV0
jS2zcr5KDEqYw3BN5rpUftOv3hg4cyPdx6ijOb7Ocjv3nChTLAFZLjt4Nkrfrx+K
OuVbsRVdyXGCbkoEjvl0Jol90ZFk8EfDAMF184zlSReDg9f5+yvNK1Vk/YaCwh9m
gJWdn8BkZtsngRu7vywQ6qT+oUEyrezQgR6JygMHqwk/xolRQEkD7UKXOaoAyl8y
9+tC5Z7qzfFKKpYck0ILRvtyiqh9uEPshQLYTLQLpsqTKY7qFWsn7l2VaDnZOAgK
thg4BO7GIi3bnY5sFEymGusDHYIR1vjphCKP0hYuu2PJZsSDNqo8opsL9dJPh+pQ
XWBl65f62uTbmIvoPv4CjmK0aI4oAyN3SM6m2AFDYqY5hCzT/68rHwOHlall++ax
N1QZvTiD2JYjosEgEJ5tLcnKfuGNVhOYr6t323ULezgQYbupKAXD5rk18RL8keJP
TLte6H2vSw+8sF0/Ncr7Bg1fYZnIkq02i8dZw+0vIBPmTsLwxd5tr7LtQxgPG+WU
yhQDkx/eaIhaPY0d5AN1+7Yb6tIGAfte0AvFOOza8B1TWhgdJLWSgLC4FeD5XqR0
bk5Tz+4ybXOrfl6bHzSyhYapetTcwjmsOVSNT7vGb5C4jasQkKXzSWoi8V/ufoeq
uE9247WNcHMWRZ2OBcexRTCw7owqf2OZi5grOkQ8q9YcoCLERZ5Xoz0KfQf9elaA
/TqDyQHlUwjf9pkh00dFgS49JeuVg/3rg8CWMmQ5puI+wS/ibQRuLnGThonoj/V5
WUR06/qdoFaSU01+dXyP6qkVtngqCOgKhAewdBU+2upNXwNsAlY/x8ZLmVrIkY3Y
gRNswDMzxfhA06p8B+ABWCFW30EeH9Uc18OCDBdD1Wdcd5qPCYJicoi9BwssoH6K
oMR3/bq/UYXMiT211UwADMv1HhNbRyf3ZpzOuTO5hnj9STlFJe/kUKWliUSDXPn1
jMRLtrJPAH5Hpl946IdZCfmXeS7KP98fmvdDJ/Tcrc7HO6FQ+KUlK8joVhvPk/8v
NCJiJOuZpyiRUzJYUrd/yvgHoNVgyCCp2vXAi6z2bPIN7hVLqUG9hNucQ2VEb2Du
EfpufFZ5xdbecsKfNKmaA1weAmS+B7xkRyZvF0MakgwSNvdNESqX/A48bseTN88a
v/AvmlQQ2lerD0RdSfXyKG5zj86DVXFT5IxNz06rDv5lyxmCALDumqzHRXhVx2V9
UcPa9L1AUGxyw2Ax4z3qiVo3PY6cxYGZEXDZzfO8axwUyxtPcTwgJhUXLz83Gcuw
FHTpviCaO19NsXOLN+lH0uUEl3mehuYyZlWxUBgGoqethhR7fydwoQe2BAAmTCCE
ubdsQCpQp7vRYbysueAgwBmWbIkHVr6bBB8qpp7qzSCbsUju4YnK4/k4zpvL24KV
EjWDqV/GHvjCj3UTeY+E1Ej273wXgdAra5kfea7p2A3/ZnunjtLn+2xbRwk4onpu
O22IJ/18lAtwycg6Prvv9CyVXsFNQeQBiiykOQB4max555HDdQV5dI0OmDfRXNxO
efIZCW5F8Ekm8l++NjmU8F8rtsHarS0HFANM0QU7yQjpY6/sl+WXyrj9N/Yr/8k6
BC5xQvKxxjoM60vHRpnSLuHb8aDKKRAkvT+T4UDpDlkj7xfuUnl8KgBlJ/n9l34b
dtF93pXgDlHNG5tHefXy8At1X2dP3KwWisdcoSezbgKJJKvLw6cpXk7mzMk+UObN
/wyBSktqdesSbYJtVU2cOzsRE1VCMlsCZ7+KmwUdLTQ19OTmvPqSP+FOGZPI65dO
qJQN2w6rWPdncow/MbxC/JxlpgMG0wfYVqOQYW/NxhM3fOHJdBTnnRtLA0rFc7r1
tLC3SJPh4oykV7bPT3wBYUqL/GYoDaAfgArioDnnMrPJRaOs/I1qKBEl6fQttkiT
67ZyEjBla8qEoWb4J858i9IcTVPok8Yb2PsNWT5Rpe6FiTOlT89696RAkGcBvelK
1YTTxRXjPGqpAK7FeMAEobE7/DFsqx5H2Vvcfrv2o84P9aHxBv8u82vjvUxD1Fgk
4umycEk0uPcu74nOJT59GlE/j53EpZfhcp9Tw0yGNouGHGbd5y1sTPj03gSnhajq
xwesOy65mUsC3PJSY3Keq8gRcaYtptJ/n7H3PtlpWFqpdHZhOg3Q963V8ZWRPcjQ
ix7KeWAvhvyTgE7cgCPuqeT+1lKWCj0ljraRVfQjvoDXnTNEYQQuonFHTztb0IVl
q6TBxYpkMU+dURjH9reBDnrAQ1kSzQYk2V7AjRtWgz+1kF09A978TL3vhtdO05VL
Ta2DNVJKeIcRHj0f6+z+Pw2TnYx/gJ99tHQF6TkjwZoSOaG1M07UY/3quVnxSSBY
tRaJSSjtIzSp1hLaT9HTDeRMPypRKnB3KFMzemc32GIp0NrmjiZGE+YHJ9bnrjjE
diu7YBEsoIup8oeLBIJl1OgA0zCyvDbsw+0fXOTDKjuM/fqPmWgpmb+wLYM7GCAf
lM5Uy6wmxeb5oq3uRlac2LUdM+jS9LCbQzOZstUW3tcLeCIZ1WEVl6toJ6yTWl92
8LAwSaaNHa4AJf5TdaQfknK4SYLQimgkyj9UhqOp9Pc4+j+Ik8c2fK2KdlhVbe9W
d/fFhFp3Q34JIpkrsf1ecHPbv0A2g6Pid9zghTA6jMIqMK4cCMnONzpBa1uXW8ED
0AgHjbMsfUbZC9CM62zTgYFHHM+mxSsC9VIPDvajQJgAwln0yNMY4JZg6X9oDUaV
r97d7CQ2hQeolVJ51WLAAbGbpMC5equmEQ6as5z5KILxivhh+AJNEUQ6hWcVnkhh
56t+kCHo25hC5HdpYsBCeTZnLJiz70x+DCx1D81g/q96IrQgaWhm38gjFaBrXH+j
hYY2ZPXXVTKhXH3gL23w1mk1jlbf1Lhi7NXFwdxtN2a+4+5+BGEXhSyk909ADkrn
NNjRURC335l+0yUeNTWgB3A7dcv694tqqXzWn//kZWeWasIdrqtNcyDoNh6/lehg
Gz5DPea4lp9EI2ljvATbslkJHS20yaZskrWUUR07biZufnZKrx3tul/P1uqvlK+I
sYCHCr9NlDlPy4q1t6Ma3eo+MEsfotOqfF5vkVhvYk2Z6EvS/JgqUNCw2GUolBKS
+dke5o+gCmt97qFoPI0iXtfGFFrL6PexG8+xVeC4ugNwCrGUYF2/CtYVn+/+0XFq
SP7ZjjdQLFr2tLk9xZYJa6FgGab4TKI8d2eyEKVj1w7NIMYg7DBjLidxpmc5Qy1t
6+c7T9G5rCp2dc0qjssGl6evaEO6k1p36qEWGM/S0CLO/aywqXcj1SenIYs4o4lJ
f4+fBZsrNr0nbk4vdgEvs0x4LRm3YRrLnOajclbUqgpRSyv8cH+JoSX9l8qVCYNc
3nswbr2E8LMXdtsLsgNPUUovWs8/Fdd3j2G/5R83gV8wwA/TXHc2Jek8r2TdQtuy
GeVj5Gw61C9icVgB4fiAGJOsQRwkxIsvLQNdz8P7aUHRAZmUJiZ4ClMHaPOabPyB
8a8vKpfAgyFHfDcqczBLLxGN/+EZsiV76A5BDpgZvwSGFDaarJR0OS7L+8m6J+90
Tczxr7MrLFBwL2sgxlTPSPruGtAo4QJXYFTXUPaVZ9UlOs5hFvolKdZ+syTnEuzI
dhvfnrNFuMdXVw+deZWv544MbQZ4sRQuVxV0fCI/bMirf8ie+bjbGFUjC9tctEHC
BcvcUmxMqKlPmmPXHChRe0PsZc4FOxSC1YmbVWyL3F067pHkQ+fogXJZuPeRnumA
NJ5ubBX1YVqnOU4JwpetHQ2lbooxPYJ6n48oHFyerhOIUbpSp/xnV+Nlwt9vTjlA
Ip14pwdtSQCIYxmXM+nN4HAGu1+9AA8CmdwFpfAjROvBsW9IS/wn55NwlMcWff7b
xjtp82V++nOYgvc918ChaqiLNb3q2IibT2C0yzYXLrV9ovFkcm0xv88NviYjIeop
fauMYSL7CwNpL6daLkyKt8ReQRsaOPZkHrwYD7wofIN1BrrLSBLfkq7SCLagTi8B
zsjoar4A4aQNJoeoR15LNr1QTVhBqMnJlgNuHlddV1xyD4kUePXWw8+MJBqqVGCn
b8h9e91YByTxa/45fCVpGmrp8dTuvLPqmjIIg4u83Ji6AtTNw3KQY0nYu35ZzoC2
IO99XRQqQEWdQWmkq8nUel4ufkuIhi545v4JCzcR6fbEhiWXpzY2eIwC6ENEd4Ng
peIdcVnqrOHX8eZCF0leiUZ6ESbfAtHw0uXYmOGA2WaqroztsoBjMkpR5mS1pJGP
N7iV3nef0wNDv+il0u4u8H3xx/gRZltfGv1WRWWZycOQnmuKlPGLK9VN9lCDFZHZ
gUmw+GW/7WeP23DHsmAe7YmPO4JbTMaDhcc3rT1BnHFEShOtdLb08dHFNUDe53ms
DHPr8VUgR4YcutMiFYd+m/duPJi/3IgEcppy4Ui/s0CXxgwCvMZL68tHszc80FYj
w4noTPLyeNW7pgtwlN7lr4qu0zE6kxW0AqdGV+KDIrGQ5bvUI2KT6AA5cAZj0+gB
MbiJ1DXNYYb2+BMu/yIVlfzoZc4zaXEhYVpufpX3ClxRzMIBF7P355ceBixn1CRk
CqnqS6HmnOBcJ2ln5bgtPO/5UYvazXusp1TCF+FICccqScNYWztlZeR1fkLE3Oo2
yBcs0SMbd7eJ+0ucALh46/9F+DvTEB+EUAn58ojlA6Og1HkrZO5hQoSCTJ2hIA1R
vbsLXNZqdVR8DRW5PRupZ5w5Z2L4iCuHeqa46ZFZnHIjzVO7I//VAIo+HLUOfapI
4/NDtzpVxe7RDHwOSy2Zs313PEITVCNqmzkrQ7HW/aD0ZsMxGmpQq6BFN83kbcKJ
jCkCNMDjUbmbzS/GKK0S8kvfukeWp/de7e6Pzd/5423LJCLmv3S/CCibBp00qRVY
fBJx5HO6FH8uxCSHCR/Fg1O+MeHGyZNyZe0JS+cHPt8fev6Y0OSu3rBq5BH75BmU
LQGpbl2+yzWJHEarteg+0zv1RzwyaQtt2XNlfafsalynrzurPWA1I4Jo2oykwZIs
fX+5Hg7tKi9eDhVMb6JruBkcYykj+KDpYt4XZFw9YOGD9cYHVnT8Hdb7K9d9jUkN
wlZ8mNr006CGIP05zleWB8+ENkZHV4i8vNGl/cFj20h/f0M5HZL3Eh2d+f24aFBa
l1mfR62G3KX21cvQaHbrLYFxUD4UwQS2Pfetfr4j3uxhOH0Ko53xFKfWkAEtTinr
155rFd4X4PCZjHiq6RMvqoB3QBDGc0NrO0xyNOPrwAWAgg4vs+R9H4OyrUAlIgGF
S5AIl5hzEaQBz+Scw5hiHDVQHp7YKKtL+4FGYErmypji7X5D7Y+wWT7WorBWUt6v
3YWjLF/3OCCId8CETzRNWtVjciYFX5HMU6pP2qDXpR16I4GQxY28vZBV1penjrga
tp8HqZIGj2izyNe/6V/Bs6K/bGp9XOwKA0wi4srnvkxniAW4AeJThQ7A279WKee3
ttrKLLXF7CLyk3/ncJyZNteF3OpbHk+WHm1oOTHD6HEqKwKz5RH5JO5EnZUWydVB
TOmJLpRlfHMaeV2UDbBF39JKTvn0qqB5DfVxhilylE4Vg2RXVMcdb789JUzAZQpC
Bdo65rQrOgUj5JSQhFCDgOc7jJ5lA7tjnSRPa72udQo/hgSyte1xc0aYwXVbtiTA
HFAyGesceh9envfAogQKKrkiAsVKAHpeezLtpaZHcJ8WM7UjZFoBTZ+HGTwCW/qt
A4aRMo071KcWo2kAdgJ4KmTdeGzWh4u/QoidLh5LVlD2J19XVHTvGvG2tQ2at6t4
iEAcEmKHtrJOTnU7pLPRUjJFX+XmK+YjSlKmZ9t2ZmJYchR3pOA28gYKoYjHK5y8
Hb36ysy7d34J/GN8TyytOl3r4dmlqPq55Rr5U1FQZm2t9BRiw6fxOK5qQFdGvJb8
CvKEgagYZTU05SMjeZ41Znu5DFEmyZ/krn4JVF8L6QjdAFnt8eemXWQqS8HaDuhL
5hmggtqKRYNtj+lvylPqr+qKgHNCf4iULSSeIXAs80CidThmabTn7ElIRGVGioZK
ltl4z4htVo9R/MqzituDClUG+zpnbvP+dK7MGEwT1EIWCyM+L45rr2Ysjm1omJTR
rr2OQKGehuvEveLZh9mkb2YJ5oRqoUC7DVKLt2qIM98Kb6TUtpWGA+VzaovmDdJV
RN9a34QReOXXKL+PyoyFO4zC95vjDNeV20alSrvXDJCl30PnSyTcJbJHBTNWwcob
mSAJ9c3bMJBn2ZErkT5cRWT/gV4CoHb35LbumEKRKignBE+r/YCTbyEGyZr8u9Dj
yfRfaIkZU7COJrLpBES5NAm9uORY/edFVlC3qkSPytTM10kQrJ9clKhExIcsRW8d
MGmzc9l9PrCvJuaXl5P6yVqjzISniHwoWlZRFqSqdoKynKPQOLEAZXJCghNlY3wW
ekRiziwU79Fde8LJW/4JviWJJaweQTbvD+fBS/hHBLIi10/moy/sQhu9WvJ52wel
9wqwLb49Sm1yMCpq59jgPhQu82X7Jtf+OqR6CVtGLGV7axozovFT6u8oTPEd+T+N
k3IYh7H5fAwWjyBjI6atUQw2H2TMNR0RZ8LTzE6hsWRntACm6DFqeobTs52+eXT1
qiQllFv2Z/RQhBAc2rakr3AVFpOvaw0aRrXP7LjfBJqj9Y9463MDUJJa+mrm74is
+RgpigEFJzm7P9gtQ1laFAFpNV6accfsveGD2FzFgqOXtA9OIcuRnpvHSfhe1YnC
xKOwFdOGHihTKlUOzsUAZ32lAqqjvugFn/6jHG2Z2E+IU43Dx4yXC9xvfWmLEapL
C2hTBNAjOinItXsmXjAOMgElRqXxRcAJjoCKEJuh/FXmW7RFBzE+5VCFclu5XsG5
BNDFlM8YBeNNR7lCmXc+o7hxh7al9UB5V0SHB5rPT3ke9NVwcrG/onOJ8whtmICp
+QblIZfECWRJE4PJggoF+GS2cWoSyXA1yUZYOuMa5PC0QfCeRagJSC9aZ6bBHEqI
ynWCp1OOwgQuLi9iwSPvQxa92W2EvBNlQpxmtnNqAhsorMsG7iy4AZ61+YNJeJrj
CnAYsYxz3W+eNTGUVwMqbzlhwpP74ObsOCt6wSRP8y++9Jbj+Pb+pMoBKPeQaoly
Pr3Ut6mHfP74pdZLtIEOnJhg6V5igeqz5qWUEds49IAyYBK8Y0lk8MYORsiR4OOd
IjccrLbOtjr5F1JW3KIdjcX/CssVPBt5Kf46j4ffHqrhUPGdU2hKl0NTDNko3EdV
wEIH0o2Jlh1lZ+mQqUTEadt54cHJ1rXIKxmGKURux+ihEf26qCTJ+2CDiAkbK6aN
yWZP1myqFc5G4M8nZgnh0nYHBfAp2bG67lrhdyXsQuNBiRucEzBkHuzSeoA9CUIr
RBFi3g7On1xO5y5c93NbJAvM7OX6cNaJVwAMonf9Dm5UvsMJ2SvSLC0JKu2IkCAy
R+/Tg1zTMtSeVFnoI0urena57tAptINHS57qe3gVmBqEnVCHwJL29/6MLYdB5XyA
HAiy3HuphKAeCnfKi07lZHI/xzJFWkjxJnEeGvb5eXwiilLSx6hv7ObjNZgM2nfd
D/XFkbafeN+phiZpVo8DdUUtiIPG5skcwytNiOYaWlHMPpxfRMxWHyYjcgfWVoTo
N0TvV7OyO0kNHYD6TH1SKED/DkBYWXZxYUVJBtj5fk7AF4fCxXsI4/hhxEIMvJYG
uuQRFVqWSbV3QETFh5aj8TOLKi493YHkyblyMVWl0OS0JIvdV4wSNvLcpFjhHrQ4
Yu1yD//s5WOdIjuxEKB6d/31CisXI3jEQluSOxgHSpkSxfyjNc75JaZhnJxurGtN
ONPQwXOfKv+fg/hadSKhveON43SzEvtWnFqOFP8LQ+9o/asxuP3KqZS51rOwTDkl
xstY25mjSqO1sSNhu1n5D9XcyaD5fcWl9F9ajGZ54d9CdBek6WanFMAdWZjW9yxj
VnGKYB/eHcezsm2dHVqD6KKBqZn1rDN5SsBbIfzXhnk3XVkihdpbC/PcX10cVsT3
UDzIiYBT0M9s+RHxfdvKW9JSWYClyPvjoX7OAhdge/tDsxRjRlcgDHYNq3HScXlM
hXa1ndCHxo4PQ2r7FzEVdLEJvxqX+MuXNMHMmgIG1cChRz3TCCCIpd6JK1rxPnJU
pmgiz6AIvj6P+AtUr5aUb8Ds81QMpPxFakuOA/90hgChFjda6NY5jEoIiCC7TgDH
3oBAlmK2Ul31PSHjHZNR5AcnFyWxMFxmobSIRLU16UQrk9J3b8jXjx6b/IgZTIEu
huUhTLdgmb1t8hhO5gKunO6ddcIGZC4hupPXoZKmRfAdu30imXcWZpcuncq+/Aeq
kqGPd19rCsEi+U8h/e6kAW0pXeHr+wYRk3hUZdo0/egzQZXkCEzm51gz8EDptdpw
Or3QZyLAY+9FEg3CI0lDtjM6seBdEcEHn6tY87kCl2gHhUlsm5F7d1MTZ88CzTVZ
ArM3lZ5LqopCfe5aejYPNUkOIceUi4E6sMJlqdrrUV3OZgb++KqZG7njLFxkaeH6
q3YUcGBONFER3+sMi/cosGusMfNZ/SFtGsyWyy0vhf+OYSYnYBiiWGXky2GbuuUA
fx2w/X0y0E1NXeOddl3ZFa01bdoNSVzx36qsUf6iLcMgo4qb8WnFHybuq+D4eWuc
6c3LqG0ZU/8bliDvMiQLClR274ikSLy32Vilt+5Ak0I4y51/IZVFuBuRZHdt94Vq
A6w0lcF10n3ZDDpjzRRbJ/coCKmfuo79TW6TsVJjXP8sMUqmbf+TpOR4IEeNezKS
V3QVjWzGArKSgoJVkS2Mnn8DVDJKvTK2xx9gzGu2jNumEykBRgYw7M5jQqLe2twV
m2t2tvNrLFUcucIFQ6RXPJ8zvsQL1ITe44GqDeNasb0eg6gMS+1dqZwHK8tXuLts
fuUufVK0XgqgrvlHT635bUIMwz9ddn/ii7X0nnRC08J8rkS/TQVCOjqq4PMyYKAM
RuxhNJ6KhGEXrUtUg2qWoKpv7RYBzTt/87TEkURaw59gQDCLO6hZq+ZCazZQfYlB
0Xi/j1m61xldj8yvlxl/iW0vQmA4/lQsv9m8koz066bPKUjNFJgzSfmP8pBggpgj
mccXA1lCrShF7LlDGhDwbbSSg22Nzb3AcqBSIHVC5HhTYX4E/hz7nagqxvC/vMXl
9ab3nfMcWQrgGR3XC1Jg6mP825LHqI/QqSEABxj9HYyevDh1p0hhNGH6xEiiYy34
SDKBEpG1r2pINeNFDApyD50fEEZ8bJ8/53GYMsA0BEspLoXW5g/qDtAq2sGB10XQ
ufvzCumcaLe+1lw+EmcwZ3EAx1Pi0WWZqER4e+LPKS0ipYVbT04+qJ15dZKT4SQ1
Y6gVsLsMGVO04IvcEpmHllstF1VAhfIqLy9Doa/+B2bPg+mobQrFoq3cNgeDK24M
YMDO/T6Jmffq2USQ9kViKRRan+a6xb4y30jSjE+/aHTAS6uzkRdcQeYFMCtqUzf7
nUnj4P0DTJgMsMj4DPjezJgFUA+wyCpnvjEa5eG1kXqqQ6hh2L28mfRW7HagVq/+
9/6yFosb8S31HdcXGrCOLwbIRP4yC47/6/ZcywEfz/P8FJ2XJTdIRkSI0hUCMCx8
KuEarLDuwVD0RnRjYuRatlr1wWpBmOdmfq4zN/UNuTQ2txqX7Bjg1sh+qPL/PuO4
u/Wtkg/X+X1zqvldkPyWHr0bMwyil0n2uZqXrwAkSm6Pf2xV6pBK3u35lC9XAMjS
M0ldT2ifBvBTobXzLbxpxx0lnZEdMzS2X88aAe5ndyeiLSXsYVKK3J0sPD+YCdxH
WhgCnq9ncOMXcBP/gwn124pXxTNrKD2Yi6oN/lgZ7hbq8iEA32tRDD0gBc+cVPCA
JmC7rcJjW+Tnzfks2pG4N9UKCVFWZISGG6lBIDrlM0IHbWhmVedzOFV9WgVsAG9f
+NOsf3hGjAbGlLQ+NEqcIuIsP2dj5F/On1kqXWGKh2r2tEp31s9rbwLtEYkEG5Hr
XVi1JJ+xP55gtVcX+WARPazUfdeCSEJZcmRpgIWbjJM3TUZS48hP1gFZpzxzCKkK
0Y9wSvhFCcl9J0RnDrpHvOf2iiUU+nelN1qpd3GjQDVNIs3axVzb3RBvBrlDHZ5g
kmjznvaX0J/bVaXZr1/XsJ1osOffpsoKmHIkzcKh9RpZ7w1nBEzC2HjEkuAKclbb
EUdpbC3UeFEKu0VtQjeolbkIEvdf/OPg/HP+tniEFaicRGdq0TVS2qtv17dN4P8x
1yjQ59HLhUF30WHPSQHHq39B1ynYsDAIPs3nUu2I7LHqerqLy95Fm9Kq07rpad8W
QmGxyO/Uax4kBgOpbGEmS/mhRSC8fTbmdESlDKRuXvKKRvQqiFQKFYaAGgbcqtDS
xg2r1M47g+fqm+xxVxXa8BLgJ3VWMN+mvjUFN7UHMzsYWT5w6sjshb3jpAekUOM3
84LYxVPFzp4eybzdyzsrWamAYwslso6fj6aBUF+rTwJ59C1M8R8g+ihso9r+nCbz
NP1m+13RM8L4Ljznzz6Crv+SI9OSO5Cm0evDztCC+BhiTm0LmeTRyTEOxSm62h3Z
2Ar4soHeBxtWoS4u1YwP9o1lmmp4yBlpCih5Ew6Rz9uzTeKq6oifVgYDMMk5ONxx
y+6yuTJMbl26v2/8e5OE2y0N9HnlBXQEmUGMSLLE/I74ReMlM3/6azfWX0FAbvj+
ZfzLJeO2tk4pbDsvgmHW2ikU8q/YYzzskg1dRmTgsh+cmZpKVvSen829r4EbZ0ev
hR55A6Q36NbJMyxWics21pyR42af0JdQnAe1X2GyJKdX0r7rOoIMpieoiA0Gpooj
NhPcvSlMXhBPLMCOhU9SNM6KD6jvGOUsUXTeD40chcyreXB84tpfw0zT2Jo+rrz4
ApMOFpr/a6r7Yh/qvEysgduyYVJH8JebZO/ILARfVcUjHZ1za1fnJNTdxtPAzDWM
s+/pLE/Zjd+ptXQfTFg9rcGkZKRvVAfXcS8rBVuwDV08PIVnFssS4G0wWdb9fBIe
aodGbPtMdyGLiD7kc8Uj/xqtYfkTX6YtRQJ63lPXWvEQQhAiq1CFV61Sh5359Vm5
BfkTWxmVx0aiLwb2EVIRgjc7MM5NqiztiW5YUZbQ0hJTGAmM9Z9E7/o+8uYRH6L4
LluOF7awXktUWvLnQX4hH6uYtBGZzrBY/TPfpMC5PdPnhh9WqQvspqR1nOZdXqqN
cWMERB/Z2qbVATb4mT6MnL/klFUfsGvkNmTjWKUG0rTN4sQ0exDTDTRFSSHRgIoC
9lOTig6YBCpCGJREzorUX+v+Fik/1/Wu8jvDC9pONg4vReXyAaR5O8Z14a81ebVg
vgl0065uoNtblTPMIGNSHSZuveta/wnZZ6fHiDan8HglHEvDzEPGOhH5t2sR+CiY
dVJLSqQ9MXxT4P/GU5nNC4dqpXBb902qRuVQmykYJVownalBIlEZIKRoHz5RBr+/
fU5wpgRLkVC+e0wdIOGsIjqzsQGYs9Vsowi5YEev6Qp5lEFa32ku3xYj3thHWlkf
x9UCO7Slawuljsj0qUgF0U9yjrx/q+01FrlUFaM9sJqtatWT08XE6H7Z23nsk7Du
CyFk3GrxlTIDcbYdwbfIbJX6KWlsEq+COIq58bP1/HlpCjG0OPQ5LHr1FNwf6/j7
wW7zGDhjSrsGmoXOP0gKo+TKvxCYHkr68anCdn3YtapFi1nfhXvWue3E/7c1cWvS
fTxBZ3dHm14/hOGW+Z3xj7npf9ICZPLHR98iljC3MtsqVfOyMtRDvolxJdnLNTo0
EFQureBtOAVtMhfbHBHpTaJgQZdna7ta/76EoVsgjPjyYYdP9CN7wBavdhVXqFiU
z/NehEt21GP/9anI89hi5Mvc1M5Yy+NBdEl7A33f46OYLDwM6kv05jXHScarvYzg
6IXu+vRBu8e0TkGraKyuCHrMNSMVZGCQZWE5a1O1OwzZMT8y+DMzhQ365qN0+8JS
dpvOIQh9iAfQKXxOpHwIvywobc8t8Crhr64SJp78cEk2xhT658LRRkbG1sS2iuC6
140hEcHkGqPrcAdiBZp0f/pm3FI9+5ae2qaELGaHC+T1jVIb6skppkMJeix2u01S
s6sdLWTrB2yxlG+o6QxDoPuknBkxZ2SATvc+PpmGWbLDP/Vp2jqFczWFpJnLv5th
lYCT2JMdQuRr4ZpZ4RRO0UysRoMZqpVykwP5LALPu0X/s/O9a98S/G1y8oRDP4KU
57zkeRjCadlvzfnHeIuaV8zDX7vKH/IFWkKZww1AwjY9xxd5q0pUqETlgpKMlbek
HAcKx8CWMjRF7eOnj0vT2o24F7mAAY7EF/6xUxbzp1K230pYd31Zfy5MEgW71SXd
pFFj+r9KwXB0TsD4KXop6hbA9K/66hBEscq447G6LlIfYdqHJKpJ36IP4hGJmbyV
pwgjzP86bC4eOFYcMVxii+6wwuGB0p1UG8C3zni73JQKmcLzZzo9o0B8rSSXZePl
Dy7j8nIYGeu6pglPlpeENF8HD6R1xi9WG+WkTZMk3gXOaY2OQTzvpjelqb56YYOX
M+os/wIOTYdsM7oNfcm1QvEkRcPMYZBFXLGAS1bItFvkD2fzyzAiHem32nb1V4kL
KobvSNzW5/4WJd1KBgaQW/6gaJ4sIFoYg5lEu4zW7uxtqE5dVCq3WH57hNICLahS
5VOooHjsMwiPNz36RrGLxIiHfNEWZgia2h/DabZLft7EKuGos2yPlp4dgH1xPBb6
7+2JCruJ5x1BI2BUu6zwjaETXNilgLZY152aXOXGlcD9tX6QLegyJHmuChnd252M
jtU1pv6jzWZB4Hh5Q72HK5KRshoPr9UowGxsU3/3p+DVG4cD04+Kbdj13WkLdylS
Z4ZiPTwidlMVU2+mvXLT2GLs4jLoOBfJHYTe5gIEEtc9cCd/bztzHRVfnC3et8Om
MDWTXa+FW4o1qQjF2BldNZ1GJDVHNX+4J+B28e6zHQmYhb8lT8Q4AXf7kM8vNAoJ
i/qxNiioqSGgQnH+bfOykEmyqVAV7u2VEvBAnTmy0p+b8YOw3pZEuECgqk1toL4b
5EMRvs8yj8IuKKBwrn1R9CftPU3PU54mvmKJOVVMc4CIbrZU/EAUQLd8GxTY9o57
t7A6EibM3skWSOll2TYKBXaH4sfhGJucUKBhjydC1D7zLL0tTmsLfFCNWXeOcZID
5UGQPoAFsjmJfiWSZl9n7O77doddcfzeOgWOfhSBcSYSDQQyMJrHgBJlt/A6q3kw
jzaVLEYHsGmGY+pNYzBKy2xvtDdef04DY6pXEcnNO1ss+bJaW8sqxG9GksYiiVce
N9a4vj2ArZWy0IC1epYowgLvm1XIX/ZWR+8L7/Wvp5dkT0Hq8W40li2suPZkCquy
h7XTgcAL2zv73v2H2M0wA+BDmWbJsW4ucmPQp2YlEFUE9BJ1cSKY8e2UUqmlCcsX
9BiNDagXVFWpDGZAhnjnBiDyiIy7m20k4uPoOnRwuCM0IM+0lYY7HkHmsqIAz0ai
/v5e6irRgc6zwCRrd+G78hxjgydrEtpDm8OCiEUBPkjfB3zzJEsIc72tsnmoEdDx
kl0FtYFrXNJBEpIjtMMCZuqx5VEGpoNC5lw24/0uKrIoEW1g9aUwrYKZQI56ViVf
NbetTpjzD3t8WtmNwYqSj80+ZPzVF8u5wSdAUvJYgI+gBKKxa+OQDhXawKD73Gte
hlJ9mYruKWU/UtS/MbQaoQAyJgOxWYMfhX0TJqmRShLpMgREINKIlUJUQdVsNRd3
V+cwn55U0jdv6Ib/rRE/QE97K+0/XuEKgj/hL7oE+Ujm5FDZ5EmkmLGcENpG7L6U
NvYhMmEYpk+s+VuibPiDsilyr9xhhaId399KBtTP2MEgyAIGlyxGSR1oMWopr0K1
5uBZPfg0+WJohM5Pto18CO0+A9ySt8WaBYYBBjh7+6MWKeFJ3y5XtNntL/Wulcr1
Q0Ade4zZmf73d+s4ES2WRy1L5fCUL3noJyDEj7sfJtmwuEawAadyhXAQEO6G1yyH
zu+sz4CzditTdb14z7IbDsOzrJ8SXThgvVof1Qw48+ZfN+dzlnNRHOWJFstO9CZ8
EVp+McsW/qX2XA6srgAP0acyEF6IM/StavMvkDBfL1O/jtE098GwpCeZK6BQVcUo
yIwI+xBceCUBZ3K3LNqwxmkjvvemqPcV6B8zdiOOQ/NpQic9k8Y4AIZTFg3Dnd+m
u96gr7rOV2tcnrAPO1PUHokNh3hn9d95wz3kkM+31IINLsoDXL7iaD9Mov6TMyZo
OnvW13bWw7VJY8xzloGeOQKgyW6eLj6+BxyayQjbl2ELBNlIwBGxL6Bg5xmnLCRd
xsdv+pZAP0KIOytwr3qYd+yxNdChRGTvONHkRxPO7YruPh2CjIq+znTMKx9uAJJl
pwfI+nGRd6y96eRyQLQelSN8xiN3N6G1GpgKc5PczLl9f2AqMC9Apy3jLiNhjxzp
neggM6P+QYn3A+72IIUU9zKkJ8F0w9JL2J5FRx0PGCCWlrusl7I6DGgISZ2IPWut
QolATRKCfKDaIChwDvllNK6jnJcRhDvR57kApe/k7g0SqHN9TLpHCSXe4vvf2CS4
qmiGcZUYwIpzz16KEKizcZiXhqnnaTr47blrbfxggYhpgkWDp+VUtz1Zwy299aYp
evK8x0ryZ1H/O4PocZa81+rovyDyrBaj8JSKj+c8Y7s6EBIJiWmyUY3s4j7nMQgy
2F9PEZ9FKGydogwBDl91QBRLyWM1KZYFPJaMwEzHmHtqGF3qt9eu3qzm132LNcuk
kypKj57Kzo/I4R/LFippCCUhW5C9AArJpkNGI0SM0muJX0yaBWZrt22WH0og6c9f
IXcAI3RO5KiUXLjUgYQ1+MMnoE5UcSECoBQK7YnVySHPJgr8x4WDIwiRDvfjDSQU
HyG0084uTft+DGW5jTHYthdfv+6XPVEcLUoTTTEW/vM6LjB4eYL9/QXZDkpJF3gU
j3XdqajI6slfLlEtH3bw1LagpmBYkTDYGEtY1MqZLM3BzHVSQTcx7y1OdIFOaZhA
mDc0lNewfud3sO8F1c/TTwiXjndHE+RpqJRyvoNQmDDu2vdHNVaagJ5SrjViWjD3
5dzvxtIsmXWDyBD+vqMlmENkmYDQ7GK6gFGPlLU5MbsSiHNcYeytP20V7m66YG4A
zyOQztPEmUJvmZdK+6o4UN9hQXPWZCI+5GdV7aRXK+3FuCAd51LDb81JeNVfncz5
uqwy8awVFbbHUAwU9r8JuQyZ9B+lZvXx0TJtYqJyqSHYcX984eAOo9fQXURAL6Kv
cFEsdxA4OHzstiHIjlPefWv6PSPv4zr/CiwKswGrbOT3wokkQtzRV3Y+HZ1imrfu
wZbQhwCjCrvS4cR4E2oU+jYF3wF5YgaE1eMTJ1IXSIdyY7kY5qgpZtwWK4OW9EcH
eHmYeTESn/2lGHFMHS2cVOeZEiT3zn+1gDsToaJuEYFvGnhAaNeFUg6lKmquYyDW
kQsBCXfiiCtuwqwtNB+/AwLym57le25n+Q2aklzPa8pm7StxvWBdrRcm6s42qwrN
xqHbBLgOm0jzT2ffaIkY4Ey266Ai+fPIreRkdYS8G00WuQX5Zf3RBUZ+VSodC9+Z
TfA0db/KUw76sh/HIXjZ0SS5XU6msawZOOK1lrWKaWfP1TtlfvmmNlWksScgefSR
xaYKEVhpc0y3/wHFbnQ2GTcaHUX8ghC087si3TcQ7nEETrEI2Vw5ENeO9ofNE/T3
bBA74jmv/fSHGF9KunuQSsDM7ZVukJuBRlAsKhb9Y0XNGSIcEHGv4MUOosLUC0f3
ZdlI+gN0UrFTT3T+1zpNOGnCSOnIYv/KaeQ5TITfOlDH9Ef94ml7XXnN/YTcwrX2
0DA5VFbvDnMmupaaSFETPplx/Tcd/yvAvHQSnAQHJQM+zqPIut1OzvGcATdy8Upd
ClOFTHdlRLCxjYfvMFaCZ5e/3qOJAv80AY5eYn6UKoFmvqqBcKuK0a0gZGJqtpGd
wYiGiIqyzkN7EbAACmDFo971abpEaGMd45QO/ykz9gBFd2XBnGdNAGfIYVahNeBm
PUTalEa0ySAy9wZF451ioK2YU2p+UG3N4B6oKc+aq/tqkrq+Ab+EWfhfxBlDlnL2
8Be+GH00D0wHKk9lmf82DcA63PglSIRrX3NRjTcejxYBVYFB2Ex7UfaPDNdn6Fpv
QSqzNcggkB4Ap5FA+1Gb44KWgostrB2kSVv5DRBJ3i5mBY8goyXnumf0DMMThwDe
g79UH+U2ZU3VdhBwpgy05cVfkGJsobclEdfkTLGkJT+YMthe2P86E+Qpu9ldoCBx
jVUilQ9a/QB8OsrixwyU+vgU06xTXTV0XkhdFneFlFvRmKJvnJNE6koSykWgg7IU
S6xBtCLkDxAKA7423dXJi9BdLH0+Z8yTjKP9krTgAJnmeldpGSI0+i3+/Nz1whgW
S2FlaKfO9Yiy9AeqwJORR+UnWPgwxEBa+nm5P9ceDrhfaSAZZcY2tBj1mYEKy2K4
oMupRjS4KYG/0Zk3PaNJiuRMy7ZooyDvC6cHOFimEyIk/Xw7jfKnmPDnCPbqrhYD
IQfHhBpYGJL11VJ4leHx1xEhieGGHmWTsnRf4LLIZpIIjl9r6fqeXivp7kCBPB93
DP4ap11IHmely6tr0IhTYer+6n1lNUEVuslCBDZy+jSWeqHtmtz+Tukhdw12E5ZH
SizpgSUHlPSY2FtTL4gd8hFyaajK4E8DCECRHq62+jNvYMw+D/e4tyhVex9yFPh8
rBjRJjrepBAeCn8FqNSuqND8nz1PPNx+lpQUGFGIvvusGZwcy5v4rbtIcfShbEdC
ctvgsv8pYB6EYJ9VMlw8aPhaXtsVfSy8ADH9mgVoFh8rjFY/+k00QxygTX6ehN/P
xntBwBTlhmekKRRQFDMIViQWjJpc77yezcfyVng01nncM/hjK0WmGP1gyzz+PDIy
iY74AS2fy4U4tdfZyFYDX5zHWrPocdAHv8gmozxfkcz5vPvabnczEFmJ37Srh5BQ
6sO+H6v5ZIrvLKTx1L17YlFKJ9OSIDkIJRRThqW+xRK5l6glWUTGHffBYsNCJiiC
3tIs4bA5iWPuSlRj8uuKWLSonJsglr2TTgDH16jC0/buZ5gl7Ugylk0aj8EPgOvm
7Cjngh+IH6H86WMKtXatfOIzFEc4moAYEVCw+zE2bwRky1eK2AxAr81IPNOkycAD
uPsxmmj7gbSoEFSSCGulEAFNi7Yfc0XMoa9p9AVj4JZgvgw6EltV49E5rLuoxsS1
49qCTaZM9VyTjVNnSNg3m+EVdrkq0GDX5fj5WVLHEfpCPI51A1s5iBa2DxC1Rnsz
8jtX6y9v4Yaz4s/mvr2j4IljdcZ4EkLkCsu8W2cGcZz1Q208Y/J1+2dHnQnuGnn1
vprV7xwYeASF0UhHswgBzJANmnZ5k2d5org6PuwfWGwYU3EAFfoJAO53fyFYpW9I
Bcjg6qshFt28YYLVbzbrzgOUJSfTyHyMtKm1eCR/WHNi1VaTEcGiiidJMtUD9vgV
GWtKjCSnug9sGc9ixtewe93oN7JeRhwWO0Xxv+9ugQoqUzVe0mlytmy3HFpfYCWN
+SPbAMZhjce2p7mVzYqdGZcGedgL4ZCtn/Mgz1hGeTTgMtqhKo9AJUNJTa2K33FS
0R2NV2IssiHxt74Re8jbuHME1qsdiiwVq+FPNYha+HadWzh4TiqXpOpSNpGGfpe3
3vCWTIDByUhfXy9x1A/m493LI68n5XMnCr5sp/O7fqKLoZatazodcBFqmYwDKrN0
iZwFGDdPZTGVnFPKh9LOruDaHEjQJi2Stq8T410X89zFlNAmLpdxp8VqASCzHFDe
NvFENB/J84a6JFHVmp9WG/MITF/L4fzI2GmwHhgJUloJRCWm6jET2UYFPO9LA3JD
sHQaXtVAhho6aa1r27nxJrCprQW693Hz5F5SFchoBdhKGDNSQHjPbUb5s73O1mXy
QWU/vGxCUT8lCyqC3KpVq60kjJsEwCetnvRXHIU1zz5RVAoM0ixi2jo9FZ/NuSs+
HKLwjJV4oZ9zGzr+JKY5Zr5dEY1eVsQWpr6tkZzQGmaZMjwEJLlgkYQ+FcLAwo1I
+JPWnR/9FkdgtQVrEDCTzRifQsRi7uRUWSBaUN/KgriRVOPApLxC22oeL3ftI2kF
3Vw0VoD4FY/EN8su7QAXrs1JC261rpSEddHq9XYtVMj27Yo8Akev09iypYzQhfM6
BMiVAuWAaZpCgCwSXLgi9e+iWDR3gJqme/HHc2OicIapmRaWAsjuOrMPaNNNEmBU
FzsPmTAhyW1//1ZAesWVf1e4aqSrQcBojmQu0ABEv9jvuxNP6FRBaRAuc4o6YxOP
/cy0/kvnBNEZKK5r2ArYfYkRjC/Tg5G6my60a7DyxCItU5BUCqAixJ5ZLkVLMhfr
+RXvlZnwxRTQXJqUAa3f7+JEJkbfM75VlHP2AjBYeIFfvcv3Zzgyb7m2r2NgAg5E
BPTfxdOpX87sJdE2HnC5MwNafoDRicLtxEv/3talVQVi1ghNkMGRM+LyVKZSuY2d
AJcBnSuB5T7sjebAdNOhA0G76PiNHvbi/11Wmf+5WDhFyJ2biEVtFTQkgkNe2j/v
PwFldF/f0nBXdJtHwd7rUwc8BUnRri23VVRWDVv20EP+4iJqNiJKfLFVTjIWeQ8Z
spTsplDEHIAj5PT8qQgU7Pe9Ke0aY84fE9Q9xnIIpvG2sGo1bGsF09ayBFj6k0kG
KKTbnSYE3uXmxWkYFOSD8OpwBc+yi2y2wG2JeevTS9xE49mmN8Fezrv9K65+EAOf
La9anxFyekkql9ZRclz0d+sXY0+hwrAL8xfgdzxVbRTaMe7mrUCyVX8m2WInhL84
nDizhIPed7OPCADth4L2V4Yldhtq2gsiUkr/+U0D4z9q6oU2jnwVHRTt5kf0qmQw
QmE2ctpAqy++Ws2WK5+AjF2nFNb/+iAdmUd9z/+zwWUB7jOHY4AtC82k8BUGkoJo
QH5YdSW8zHR1e0TxO7tbdx7I7rR+3r/Y2OCgd+BXvZtuELsscWyWT8Tw97d4tvjG
QizImgTiZPxtZOtXEoFoVVe6Ij+anDcRgmruN+JfwvzU1VNbfF5aOlseJfCeszW3
bLnFaQRl9VKkSmwyVTWQyyeOuxxPUqy6ssNv6nCA7TeUII/ntlsM+RvzA4xTpT+U
9FNbpv0AKWKZF4/hV4J/686RWrKPP1+7A1QtlgtPStPRUpKMqm6vsrHujsAUa/bH
O+MqbKDbt1JtWWltXsGp899kPS23Knz8MF3+Ya5Pkc/Zc9/akDHRpRUy+JjZ/UVU
KPHtNIBbwpmUvXr+nM8WlW9ZOMf0Wh2sLLbv9yIfR3YgeefObT04OcffFHUOecbi
7hDTOGaBsybThf0i1mwbhFqNIdkYNcVug0/H1uWDGVxIya4aLyb10ySYUHt+YDmN
ti9qPgGats5CSF+HA9A9cSR/OB2w55/zju6viNiORHdm1jd06pAcmifPmBmX0uEj
+3SXkHDiSVO5mOPXappVr7QS/i4iIc2QSmxMzDsUq4mlzV4gUSOzLqNkVcWyqXx2
PCRVhGYrTsD1uLIMzpWfypUYbYDTmbmBgJJEmSMeuq2jrn6pGvz2n7q+FegT/whR
zQ399zQwKNHF3WkTpDqL4AWP9ixeAGmZ9EUtqeAf3yDy0rLAyic5MIl4ZdTX3RKw
X6/RzX1VFlfnhmIDgsLAV3lJ8A6XqIyF3pD30vFXuMMUSFWbw73mcBHHExVvxpya
ei/pGUqEY7ZWDwWOmHZIGvg4H7SfzjUPKBolRdKGxqAZ18o+uuZt80TtSVSIay+P
PQ9wE5bKcdeuSetdr/Vk4btry8bWldXvVXooERNQd17XGnZnDQw+BxUzlELbAwg7
j8XpdQFcb/TnJxzW3QY86W/qQ1TWT25UK3a3JjcImr29sz29fRpd2MvLO9Rt5NSs
HErJjd9yXW5GW4o0m4pPmXHJfKdwoM8Khu3Hy5oTe9WhZswwRFWP1T5IKULZcuOw
HwCRFpUrho3/tXmu5s7fO0pobHEVmV6DMvlF+QHqSq00zoi8LxHSCz/+YGoi1JX9
ywzwu5GCM1tqXD+CT1j/1mvqySOwtDXtwupXvmEz8YWvtPygXfjsl/JHV6+sGrgA
UPLOPNOye5vhFbVYXFHNvPu5RXZQjmxAdh/cLpeWXRkVqFnWhiz5vGyxS/6LijtJ
N/Ox8zt5D4ZQCSlAG6bFwLcHe7bAnc3/f8Kf0KFbkMJlO/81lg4lTdkzCwb+NwPj
NzpN1oz8UvU+I893uWnZw1XpFmOmS7UxYlRDZhTKTgdphHnfT9905KhM5vaHRcoa
+ah5s1NLG3L95wyMsAVmaxVp8hSN61nDO43m1wTi9wUoASGSo9YZ4Sj3/iyTuuX+
6THhgfCNgfdNtLUFNtBQwoEk0zA+TiehfLUusjuy25pRsUOLtcEdbQk2T/qw9clW
oOE99r3hE+XXlRlV3IhUIwIgFUEVgth4FJ6/zmB1ZNECjn8tKcVW37eyiKlikdAx
RE9Vij0+A0EmVj3r5dLhcdQNrpox82wKFYqEGg2dxTZ5WSqLcSLiqfWepP9Loizh
QpgbMg/mgXZu003Wis8BAxm8veYMl0JSxdf82h9Wh2agjvWG8HYbf1XwRIKzyJB4
FaVnNP0/fogkD8piBkmmP9WFHB0oT9WIYkmVzRTRqzlM9bd8/w557KK5Uc0eCUnp
1r/Amkwjlclz5EjZzqe1EZgByglenz4bgODbY2tGRHSO247P3T4tnbwaQCDNXWl6
0z7OaaH3YhznPWZHIoB/SFAM8C8YswKS1Bp45M6ZFtpHA2tnWFmcV9KGNAHOYEe7
23L8M/5dSjDI6qjspT0hp5irQjbnRjIis30XBPtuYzqlkuLPHq1bTuQj9QsMtau6
pNS2jKoCtIdkdTOjyE+qgeLKHSpU7x6ygZK4sX+fUru0bw4xGNcdrVvzLtJnnmAC
3ZBAKWzzriCvYdGPq2xhOHRzska1vmdCENFxgPf2DQGBiHhOUEjf5GEwBeo3Bj5Q
zYMNblf+qI37oBnG8KxyM65eYfjPT0CW870Cuee0GEfIC5wWhGF0R8+Ima0Y8mEL
NPk416zAullnfO3Qcx/2L6XXkOUl5id3s5cc4/k+KIhvJNqKqqmGxOTC0T4xtbpO
sRVv9f0FBd02OfyYWHeRxuDf1Rkh77fxXVykR4HCTmLHgP7L7XfDohVELztMNjjq
9+jKQv2x2AZMLHFxO5zgaddM8jY6QLDVNhdzhsXEDb97kpqAAlgDfekvMCk56qWb
iopfP1m7iBiIEpT70DJbI4RW9fwk49XYY6a9seYeffR5r4O+2Ni0tw+QuiibMWrf
7SAxBUzEpXF28Elfp+O3bVtAbrUgCDeMCUcCM7A26LfBVrfMpNvhV+zVicsh3P7c
9tESczmzUKntamYO1wBOxjz8aL059PbYK0gaLAYHHjy2sf9rioCKMF4p4RRSdHzw
DpotjhTDex6uPNj6p4qkmzbeaQ3kMxNyEWCl8WpGC3rARXqWMR58mie/qR2SrKaE
JlqXXgI3y4spnVl3zeh3GF6YD4CID4deFoJS/O71N0p6cOUJYlBALbDz18eEoQWO
gu4odIfQPGmQzKw6cLc0YY/DNYCNIh3eAx+mEdXDtnBEEznyFH0+jKScyx9Wa2qU
IH/ERUkFjHs2QLLKXQzKFIYFT1jw6kdKnWRTPHMqmjOwTZvW0vkybf5CP8bw/qAH
tD+s1uUSIGHRL5aU6K+XdZnblqKRRJJ7dcx3vYqH62Tfp+ocvL6Pk8GK0th3CPQx
WgEe7ErOf3diR3eQHKjmngVh8c3qSRtdgfFkgMx3X12uk/kZ0RU0ghH2lTTOlmux
oNNqs/9ot94fjPQXNM+gKXv8vrkieiNNjSFHMGCAwf8n2BEUZDbo7/vErsymi57M
fgA6ruSh6FLAz9h1B8r+bCzckp6eEcfHej041opZbsUUrpDAxkbpygeDdxnao14E
+ArnxJxcE/C7VgeSThSDdi8lAhAPLnpIvD2gM3PU1R165TKoDwv1K8XDJ6R+zKfx
0j9w0KLEz8T7Fd/g5ckaGg46G3G4+bv9Vvqjd7BQiNazlzSd7vTbFQhQE9r55Y6G
vtTnKO4MVIcobQB2RIUcVC91EAXKKIARlsa4Z88rndBtTivoRwuhEr0+7EcjIOpD
OWytAMlyWsle9hsw/P0YKDG1t/fqNTC+doSdvT9AnHBXSYQSXYaZZ/1ZZhY1fXuD
r0RJMjPerjiuFRCnhkTUzOQb9Z0729CQ7gQkNtlxQzXFPFZOB5MbFdiJUB6k97Hm
GLjZOFbdmq3sJmTvwH8U7Nn0v1orLtaAJmtZvO+jsNEyAcpL4cUi/OW+yB8RvEN0
35ImeK87qHDXOqHIjb2m0ADgyn9+Ruv5Et0/Fe1whjv980y8Hgqo2kV9k4iKQJ8l
YxQhlNyIWjjyuncZTpVleDpxEW8IbGA66HrimOzhNJD7yYjtk5VeKDJeLAddLGB3
nON6Maq6FycTwjs8X8BJGjlCNtjqJbdMbHgMpRsXTeoFjY8Stb9ycueqNj6pOf48
9yoQru7Ow4JrKNYSDhVwta+BmCDQXSXAQhhyywut+09bjAf4TtblVf6YIw/QcQLi
KNQSecPQ30lDa7ksnE5pUYZr45r4kYxADVAQDH1XKKJQvbbqFxTkKuv0Rp0erS6D
qLlCcqbkGxdomsC5Lpe2HcN2VMiJZ175lpVojnBLHVl/ymHDnhcB7VJzN3afTqzW
YZa5AJMpbI3IqUyy8LaXdwKGrjqYRPWOBqCQyrkm3CldtNFRpnEpqJ2nBsq/D+ZF
gih8Wv/xrpTIbhsVwhLtMKrPaNvUDIEA1xS2wpMu14hnorPpwKngImCVMgPmTd+i
LIJSC5/hvYleUlLI4aToJTaax8pVDidfQEx0WUlw+fRedHc7UEeDyXM+dm3GU9jx
InhqsE4tnrhAEsIsXr2rLcYzCeNbI23LvbZEu8q5gagRyJKQsGXDoIQX51qNOqRy
ODuYSTQafZ/qhpalMEVIYQd7X0I+AyE9IZJg2iW9ExaJykllyB4iba+E/5Eex8aq
dPvEyRK102GggLS2dS1RSLoHL4uZ059A/mGMG+C3lGVEUCzlLgZq+V/HxDHd89o8
qKi6XltmY3Iq6wpPXQa80jBQRTLbLxIIfgWSJN3yROfES0CWJEAyht/tML9Wqc0U
mL/nyuBb19HIix2SBkH/GdkO6DXt4092NoZ2U7d9P8XgR5NVVwL3W6oZNGeY2yhP
P0j0MIUhXsaEBI1ThR8STJLs0O7YpNKetfpeKFjTsOvj0r8hMYkpAA9PEYQDKuQ+
3277v7/t4pxyR4ijXyNYReIF0X6vClS5VE5OG+TgenTssUmId6Htk2j04Fni4+JK
V+Xz1SzHxTALraZcCs8VgKgJrsg+cABJX2yJBQ4Q7QAhLTKNFM2zUCaXkp3gCmcC
vG8bWARDBJw8WfAXPMe0V2bgeOHTMjlQ7G0vSgsTt9UfMWuSIHrqmEiQ0bvVZIjX
MO2/cU5SHum/pFlcrFfppZ5EmSW62RoVVgK3ehUGqxSNHMDX+J2lI6kPCajSJ5+k
dz7gN/2m5Jm82q4mpc9K7iWQkB0zrKerTXyx0oDWh5VI7bGWIfwZE4fRqzM5brDk
3JygZcRpnPbKPjXxWd32uLcV1jIQaC0zQ0ByDSQ04exF6Fy7Ny+sz+gXvtQbCAGn
lI7R9GmD8lxEDf8mb+A05cnpX/pmg5I7sdEZ6MwHQ+Z8NJ1+InksZTOocsyiPoJc
Wu83fcKkbRa22NpP7j/LVJIy9Y1XG26GWodEtcQiHphJ36PLyI93/HMFED/i8DNK
QOabaIzis1KcoMJFVw85vChlcE1Ecehbg0PJtNgXu6ujDa6HxDVSX5MgHLrnfz0J
dx+WDsCT/UHGEbl11ReahoALNvVcLQYEREwmDwZHjHJ8Ywhglx3nXdl8HrKK1H3B
+JupWXPHTxQugWgZJulBetK5m94AEWzWVV8hV5YEjngyduyFeCZoiGurLB/SzwLJ
B+yOyKphaM5/Gl33qMBE8OgpfsAWhfd/asU66kODTVO1DbqmlfCNOQDY25AXM/2Y
IBYTq5kpiUmdcyXN5NN+7Yhv8EQWLiV+eQy7LIT9BWoQ4Cx3sqLrkWUI9bAIZ6QW
E+CIG/lwhtAIi/RReJ2Op7s0idqN7W74wkF0PqBSd5wfrJ4Q/Yc6AX6NQ//G/XAL
bcMdRc6CSMLbM5RhbLLAeIgXxBBl7aaIWYeQiAWowKYwL/a4eyisGNaA7zjI+EGM
Qj1KZLnqfBKzb5T/awjRzWxGAcjl2Y4caC+TXYeyVkMaNQh1+unTSehrPehcX1r/
TnU9KPFXDVhMGZXVlCtioqtitd5+qj1IDBTur8CZeEfiI5Y6zNZ/aZ9pbNDmqQqZ
iCrBXIWa4JCiJ821br8wF9qLgAuyahq4vsTIj9mL34FOnsjhwS3/CxM9vzrkwDp5
AN4arCYeN2ORK2VcNEtQnX8LpCC+0Z4dHiOkXIRLuyeQo+4eeMUOLqawupTHFqAN
qqJQ8gTjXc+1OjscAoMpUva/ZJN0Fncn3hAXIkH11EhSrAsNGyqPdhxoVzJye7Zn
IyY0X3S6hauNXJOVIfJ3g7ngwhS+YvSSGcrD/IGLbJ9Kzse9zPILdAc+16dNJ2E/
nwheGe+JIVy6YEmSlNE3SXN7lrSBzoXpgU0xum7j/yFtrmH6nBILb0+EVSOahWKy
PYfN93W8GcMv/p2R7/d1XaIlixjQp8sDapkW1TdVt6RCTCOhGvHn3IskNHHAf12G
ieuAF7ZWSHpBk+YALMiTpenwmBlambyBWB8xDbu1VgUrGyFH6P0smIDAhb4WDpuU
o/mwWYSivOREU3Q1FAFpccOOFoUQLVioOYWGq3PbL3zHAS5hWk6pIOofNiFAhjUU
piuVzFXStcplofye0+HWwirgUbw7Boeai6/FXKhjVaCK8/fL4keAtzzjHPeJqe9c
V1QhxNUwR4AGLNyRM6F88mcMDQe//VX/8om8U3Gd5a0wCqdbAJuF3U2ToPfL1teZ
hOWFJ1kRd/y/qw0bfnGOTqUwER893Zg6CfeWF+3I/ICLX5WikJpeRogkhXXOtSnD
vg1xiY+kcf7O7MJd3MzYardPdT0FylbuIZ5Hyj1VwdHFQvO2lY5KLTloerR4mKAX
7pVFWcInxmMlNZ5hJ5W79aH0Z4daSUTK4W0ctfzHRdU88yqoMsXpyDHj0GLprYiO
ovQWH1k0xe+4j6B6T+KzbNkFGnUiKDQuv9bLYsyrCUqy03ixdnGWaD43PqZLel3F
YAkAK5Bei76ffpxbo5+CC/mQPBWUcn9kKNMn5UMg9BUDG8nygPqLf/eDejAoU9Sb
y6lm9WikTIjU3G+SDFQahBIQeUnAMGm2FAWgHP9sXhRXpV5Bb9OBCRNMSCXXQLVw
qoLGLhaiFZc+r9D2XrDVxUvFw0U+ruLhztp/FCeIl9hdgyP7h23B1xC0dio9h+7o
xu98Ya6WrVUSK6q8ZAjUFm00xn6aXEr2VtvXwfFExtK2g95VWULdHz7Z8dETXY8D
DUjvmosp1HufcX69WlyRx74oNFrrjFmoI+ZWBbAhyo1J5QNfkP9lr/FgqvgoSFc3
an2FBHzYtCrjxq30cu5kPCqGdh5SkRXCE1Tosz/31nS5j0WqeTnVM9+z+m5aGiuO
wqzLwAb1AwLz6lSZzK8Cpa2ihHEzj6jlYOuazHoSObzPIzhq7CYo7965SexJ1YgI
dODMPEzF2DlO5WXnQKxaJmv6j05Zd5P+qkaFtKnVipKb4oB2L+osC2NHYQpmSDiu
k5gUBPA0bJWkKEzScufM6G3x9cdiJTr04+Bgk97RSw4S8pzpfVrbNbbnKuSLFvzo
35WpVBgdgsOletuTEbvZWCO+plyGY5itd/Epl/aL7JN5rFJdi4Ezn/02CUwjFDX2
M8d0Hmglz5VXWy5rAasUZCiVUEiFInsfDCsAbH+aHgc+VLYIWyZiv/FrD0/LnEwT
8wMzrulOWCBAhdzeimJgCSiLp+jYkDypIU7u2Jn8OfEF0GI/5/BmXXHSG7VMJt0a
9SbxPkGJKHNpm7s3M3+sQiA9nW8VF2pANnw7weZjhCBIl94nUyaLO4l6fYYJRlx5
ue4nJzOqbWiETXRVYjgIhzHJbDu3hGXVHdnLof/hFcLQT+AWZSwBlHm8rgwRczpW
wEmKNok5vZxBvooRiE6GNfVj63OxF1D8T/0qrk6vaDOTO6J7hkxal79lTe1CbC7U
+BYZrmlgeUNh1A26NvYkq1hk3WOe3oEGzznSNJheTtXcm7zDLbuVji0WvTZK1rIc
6mCqVl3HZDC53K6Zy+4i1OcYW/6tg3sPanfatOhDC67xb6UjSnZruLvcUoGv8gCj
MUJrdJgYysZLfuJ8KFMAjDgKj3FM/o36t6KpHWykvgvW9eG7OfthC2zGpmGr1PBW
Ek6Tq/fq66ZyhUJ+xe4sC+jDlBSc1+XWLCIFYiUsYGrox/zZo8N/85skdnKLVUwe
njsPF/jbfBb7IwIja7FLiQkgt3g6BpZACYKO+5gKZuosphPw7lVF4Fab8mASkZnJ
K9DCxUf73aExjcGFkQJ8HtMPg0KCDiQjo94F9uyqpmNUOiybucZ8iA8NmuN/d9fj
NeeFbyFoYQYKVj6qNBHdT3fagwh87YHIW8SAqaNLn0/UrcSw73pFbCitl4k+Dcts
FFt/TsDKf04STmNjk+L3+qJxli1lYvPDCKdadYhVkErT+ekFsUZh+kKpEbww7Nch
kur3y66bAUtC1dRxKqLVSEs8oSruBVKyQRqeFvio4KLjawhnyaTeiFkhZ1YfpcNk
vcYjf6C7KriDQ0AhK1WrOGESshqHSfD1ilUZWD8Is1lFuDP1hnqTQnVIHPKe9U5+
p09ErMIuMv2w0YwNGcmdU4NKgVezogE7Jzb6ie+liC9p5MkTBtJboa4q3m16jxsp
ZHSnTQcHPYGqP3i/XtwH1WKs65iG+YHtwLYQEzmNxqR/Cm3n0w1mMpUutFYbfkF6
N8YB7PKoFLfNzl/eJk2fuIvwNcjuYZSNF7AsOEPSHBp0DPhGVnaJ0zIve6vcYcZM
l1s970ZyAdsuxYDXD+uNJkFRwVbkw83y1HFNAMp5GoIvAKhppg5pK4omAkiRLDRH
bbLXC14sHxKtOhgIA3HdHwx8/3m4+VzCxiVO69xz6NAV19Flk5xDbgZ2nVaZ/UbN
znxRcQ7HA+l0giUOH4cO3oCNtDFV+47qZN6MWczJG2Rl8Lw/3f5lviAQcJZyM0p+
VS8MzQiZpCYkOZaA2rPGb8+fq5JFx3zPdzrSKoOvkjEMVMNk3UPfBP/Ad1D5tf0e
+G/4zwYSAwqxyJwBef4CKvAKI6T27nen2OczTWu0tVgAWKfbnOdRbREBXtVfXkEF
qrdMT7Ox6s4t6sfuphiOLSixFNFqR6ga6VkYcgy7+g8EWlI2cRV8uEtnkdFPiJTO
PLlibtF3C34esQPl/F95byAu7nvIx/P+u9gxjy8oIP7TCUTZUS6KJ61F14bzYEV3
s3+9Ony2eZO0Jduij0ccYWzQL4QBa3ipXfiTnGePOy8GksReXBoK9iVTJ67RY6Lb
iAsMzPqr5t39xEpQbTzDnVdbOguM/VGV22kG2LYtioMDutITaxan9LPzaBZsPTPK
qNCWD1UMrn2E8ECQ0H7dgg0KVwD/nDVRrz9XBFJtsc8mBX5pMthmBWI0hhPUIKZS
nFw6aM205Lz7Ah6InNv63arT6OQN4unDH7Pz3MFiExomS+oyKjnOMx1V46TQmESu
86JAvb6XjcIQY15zyIFSpMRdDyyLWvzx5IWCow9yBZnxo7Y2bYdE6+4H9HQDaZUs
Wqf+wfCfv0ODxKIStHDxzLRWZKt/8CTipZsaO4POnmYSQJnRhx5hh2JmF++Ad2TM
lggDrZejWYLo0JhkdVcuwg3YJven1B+Mz2sGMG8kOIq8kAHlvEuTG+1rQppcfIlQ
cZTDXXI/cilcH5ZWAFtc89IZ7huDSNv36MDj1WtfVfM572/ns25h7Vflh+ioWfYa
7ZhUCL3MZMHY9qeu99JBXRxzhsGTs7KW0nKNQZkdjjvxblYLefa78VNH7L8qOH34
L4DJn1ZLNgVUhLd8sR3r6n59dak1FihgDigLTPGVfm64ZMXZ7pRVMxzcAnq6pEEb
xe+634VSrTez2xbFQn89w8xGMhnO4pqLyta2BfV/ESnw7hGdMciZJAxSw7+ePdU0
VCprfapSD8rhq5uyzBCOQs5WB32zZR1EPQEyzwe9V3MTvp//qhHtS/tCuO+4OfLh
sVkKRthwNqIg9n/z5BwRqYvu51uRK+A0OzhE5k+RkCBYIvD0xA1iOG7A+LnagfNd
5u/xBazEFVMKzQqmg+0kflbZCCwKq1ObLCmVx3b+KJp8zwOFKMKpnIB3a2ZzGQBF
uUL5fNI/9yraD/4Eg+xe13LyuDZ4wrjOmGvQhtm7EsJ7GjBfws4tNht2dtgWMhQX
cZlGNdPK8Re7zWpuBz9OQvEeArCUe6gHKXq8pkX4dgbdJtTvumC8qPlalZOVHcgl
ED+0+S3HMPFOzTpOy7MXdw8cATRRfUQtQ4OM53ZzJ4jWRfrB1W90h5Xi10jtXFFY
NyVq8/I8v3iSwlG3sV13RHlbyFOWDa5P/U/1gWjQfA6rCbAr5lHGSvq1KiBriLDs
gS2WkdbBOKL5lLnGEGqKPYorS8JV7+W3Xf2DRxsB/z58tMmlUcy4yz/h6McWagKW
28fa16IsCqfMdffEBRNRxh4EBoJWUkDwzntBS66pHvNaAnZ8OwbeUYzyVHqMS+Cz
qwj5gn1ttKGDOqx4s9atM6UC0z9I+lvmWa+5cshR/U9PVov4KYWmRQXYnAlZB0gG
R4horKBkR6pE4a8qb27B6LkrYCM0v/fzuUE4E/6iE+4ZkO/h6VZeIIeDBmoyx1Ry
F+4DEVgLdW2cGOK7l2Bpb6qHgWYHeTBCbd9xSRQA1b1ZHB0SEsh489o7ADMu2auB
CEL12CGJJEN3vrkwP8M6HIDrJ967g8JMnI/XTGFaFH8/+nqlvz+3WP3xqJk9vDGA
rdIJ/R1h+5iPNOilmKdLt1xEGIiqHFvHZ+ilhEzSHf4SbNLRCi3Z0L+w1JUwUTRI
y0V905H+/f5M72S2Hwz+LF83hmYcJLiyx92xSdlD8Y3sHe8wRgLKqBiody4i6gSA
HVql7xT1KrWtptRKvf2P4CXLgcL2aIABHiPHT1kQth/YxQiIDU9T4R0pMekiIVKA
2QDT7S/Ku8HBTkodIgunllmct0r5n/wi/DHtOIFImBEPg+JeAgf7YSAOpmZfac0j
cld5NEseofPRHqzUAVrXxzBPowUhdHfu347dC7Qs3BHnbEacT7GWXkJGtLJGCszK
j1mS+9K+fQFakl5R6Ju9V+IxEOx2L8WgLxR87QHRJAoJ1S47xliHUYycv+m9wP+0
LhPVvv9w51Yxb2ZaZFbrA0RrUWckQRYL57piEryn/wgYq2P8i4qQS8RApJ4DxGml
PrLt1bQ3NapVom0xmiLBLkp5+HgUcKIQVw5YAnASc4Cflzju5+V97zsQz5a0m8hC
5nZ3Vaw1oTfQhU52a5r8VA6y7JXr2Nvhzyhs2yedWd4mlXa6xs1qS/voQadYAmD1
+aZ2LUoHotketPLscYFEYcO1BFqblHmCdm9qanGlXFicN/pvyB+pCzizGcdByLlu
dVhwttYfjm+oyj0hNPrf8sr6xmNRvO8wGoIbqJC1OwFPRZkW3+kSU44oFR8YheZI
MCvQ6DDzqPBOBGPvRCXv5hOXgGsX+UX9P2+Qrd9yNCGoxAhoJjk1Y7TY5BAABzxg
tGs6r86D90wNVQInb3PzahPUpPB5MCM4KLMH/vCwjUcenV2BJl46m1an8fMTX1Ne
c5iLpccglk+YBJGk/zAbfKnVhIlO0GuP5+3Kj/imqj8yTSfRMq5wxkfv85DSwkY0
R8Bowv64tCrVUR/+kPEWI02upXwbg8Bt9Qp/gddrw+l/8D86HPm/bj+opAyAg6re
6wbUr/dvK8WkGil22QVCLUj2vmI0b+H2QDZRUjUUYpYFNFteVjmbxtenDIwRvzao
o4dIqS06VoxdRo8j01b954euTJDjtT/d1VfoerVjYmRkWRMOkyvGNwKO6pY/7/eo
HgR7o+P8L/8xvvtbBAgP+zPFhYNJMTROlolUnZE8DsSUTUyT+ikdrqZSV3xSBJ9q
dCjlTsTNZX134FIuCxigBFeWhSQVy73YdxB0LLALE+NG2tkGW3eiPyOCpraohTZa
poL0VmbbHsZczDPvTFR+mv/1M+zBk3pnwK7s3dlMj8ZExmFp4BZvasfrpknkaqDW
dj5cKPHtAaGdxTRrulkvyC9OV0jRBr1gBlocZtuRIgVY5zZjnySpxuhr21HkJGAf
hzrbAIpJub3n/606zEgYJLkznqCZBLXXbwa18Na/rGemSnekC7nKnpiWlZYoZw6n
lRFNFr0EWomoORSpMjYUZaCfeY/kiCq94B1xfJkkJh/DEB0fPqgWRBjYKH2TLHih
HGuZPgpdUUFP7rhF09x7oDm6G4sA2imKaNPYRb2rsboHjciIvBzMh/X8o8krYcRe
6YamK8Gc5ahELVjsSevBlPTXQzCaAWRiyCq0+797sH1BU7XZ0Y4LN9wl3ZOp2v7P
esjbeGxXKLno14q6wZsI6G+eXLQ4IjifNa1Lmfn75dj//sSEKM5JvVuD5r3M4dRU
b+LBJqRnexgczX6q5NgaL7kwYW8nqKFjUVGdsZai/Z97YD9PU4LHjnHvJg1OsIj3
lli0HwfVy7V7SIl/wi00QYnJyB6duPoTFuWO/mjfroTD/hKAtRgx3CBxsF2HTAV3
I9ZqOpc0gL7SOhc3yihTcoJbbjbzeEz76Mq6/oCSjBEEGH9usY2ZtxcRneGWWcLO
ZaqN8/sPwzHFOb3QLGtmrzagd1VwRHZn3n6q+ZuHbEX2m8PRByN6WC7Fin19rbd4
biCZhasaauSanndlPDv+NzZpeDHJMr0gWwOdZ795O5gB/CpnaIiiB2VUvpZaHLVR
4MpyYKphTwmLB4iUxvQVMfcgUiZriX69aLgd2zalSx/61sNAPGsYsRsjC0QcgxUE
ZZS+sGc1fguAXOaM2Tr8wS2o9o98uUQBZXlfUZKP+K5cHZfxZrpKuo8MVvZVojDU
LRv65+uvB2nLl2rlIzjRzpg6QoCY+OBUXgRtKh85JDAogI+0HWUPsAebiPaAplVk
kyXCjukuEzlewFUeBhzdBHUHn1CVmqd8vgHdojDU/X6OSisseoSQ76L/Dv5BPcQ1
XqwN6rhpIokraJv2DOqgZsqYeo3prFshYzKtkKYdVDtv2OH+UwTib7nhP1y0M9d4
t6QHlzcU5uDvWO6we1Sm6hRQePOMl2MACttJGxgTwCgxS4aWuf7JPn1HPDpSmWj5
DJo/8yrk684QJEXCqZtzgdmdYRbeRLl/cXNDt2hx4gzEQsUTrjWZGlb8dUokJ3iW
1ZzybG7FIg8ryUU4dfRkAKX+XN3LoXSOkKEkiIladIB8kknMdnklNVrQkUfXThOO
4F/aY3bgLewbFs/JJyuEvIukmI9wI42+g/EZO+Mtto0pYPsr/J1HrJTdKnLS6L06
BlJMQ9EqA5c3ORMQye4vi7UYtefLphNcKYtt5AU1mrCWrpqcEi62GEgYQHSEPde1
+4iS/0FBMzROStg5SzSWAzAGpWMADmLm2qPWe17ex9ZpqKN4PUH73nx+w2R1BVwC
9uoo4wk9rBQFCmnllMOLxWQVB/JjN5EBRD2jifcM022vwRltFDqPI3DTO2/UcVMQ
0ItT3NRpuXOslgEf1D9Edb1Y3j7mbFGHDg8zDJ/KFE8INQnDYXbIYlGWMSayH8kP
iGjf5EoTVuv71h+2qdXlfGqTyfYfVqqDDbtdxGSro4OoXBVT6p3A6L/iT9py/ebH
+nU6h9ulmCtxrhRkV1OCEyWUqPCsey+N8OeTxNwQCFmSbl/IXc97UK6TKiWaJgIQ
DB7FGgfjEbuPFB5/lPX7nrcS4eDeNjVy4rnfb7vxD8Fv6eo0UgPatj27Fqb2+kxq
OV3gseKm6TmV//6da7xAjWiF4b3vxsyRbgoi6yQJ4xnex/rNkUGGd5P8Hp5ctJZO
YZlxRZC5o2qJoXd5oEgOelbDTygSSZkq0P7zoC2/YwH9L+61e/qw4UMvWgdtpBTg
zO3N/n1B67MmbSsvlhBN1zSocf9sjafxCm0NcYB4pMlv2UhydoqbtQH8iD5dq7kx
LyfmhRcHx2PoW7gb+apsWmfkZM0uK72YLBXBiPPmgHYpsKBjpfubzuHgLqlUkkWv
tlot62Za53cb8ed8WQhCY1Dd5VpeezAzxZwBhwxnl5zSl3E3PRlFlsfZcxSdN6pR
j4XoaUfnduREQ6rb0aU4pfkfnCx7OG3YK5xL2vE19o5NijKQBmKCmvfynjYUBNOK
QF3vzflc1ETRFrU6rQhHk9CVdf7Q4clDEUtK9X6Fmc6HyQve6svOlkx5r0WT2j7J
ATIDXvNWvNLk2lccD7dQqzWCElLeuRep/cyuO0aXiVDtVcUpJdK3pNQh0oJDErEK
sKmq4BCfKyxUMZsOSP5i9cV776ndRtVw4D1DnX2sxM4Mww9J4H+m7k2CiL9QXr9O
AvolDjXGMqIPXnyJSmOmJb5KLtSVw9VQtyMID3U4JObUTceaBcRLBXnCKHK4rcVH
Bxui2W+MAurF6+SG40yVdIvrpijyi17S9jUWOoHtSyIVo+fOqt7wZXHCxOcpqG3u
EJZLGOkNtq4VLxqVjCb6Nl2EFLgq91/DtGf5MxJaz6n0pbOXpzPKHEcM1eUanlSr
ZJiXVPHYlW0W93FsMPvVbzdu45w3DvA3hAwZsQhibZx+sm6HAMyzREgqJOehTciU
IaJfKcLmQP2ab5xPCMMlaqDZx9moNbpbzkNVlwpJTUHjmYV9dR6JF6ul2FpOu7Fq
mia5sH25b5HyUT6weJTfWK6OrYiCGiGNav1ZOqu0UD/R5iw0MRuYjDIVP+rw853U
bjxTthUQUWaOYGtgBCVzFSXhuZ2Jpg/8OROWvEcDWCrl2tfdN9uXKIimqaFe4DnZ
4cpwRwiHpsj6bdB4QhOerwSUQgRuc0mQc77N9M2e0clqTUTNnv95P+9eTRdqtXoW
j62RTEWmlQZ1Qo9qqAoW4V6wFE5p/gX3vYZaSBNtN9Oxsg5Rb6B2Ob4j+jV96bt8
Epb0ikuOedc93edVGhLZxDfPEY+FcITYsvH4ebvNe6NyecIFVwKoXJfVCqxbpTxS
q94nSe22s4y2o8dad2PMTrjVlwa90JqBlsPDQxo642x1at5+yoGam8F4RMopD735
nQz4/Pq9qEyxzv4h2DI1VTa6/NwJGW7dSlF09jXyJK/90v/LVPLto0B+pTJWPz1I
+InSrQ3OpGSG+1wbgwuusCabn6MTLOSiAtV84S41ddt9cs3UK1vdoYxYRJptgvp0
tM4ZHfiUW8CjKe0wm+sxr3cFLWydf1mRN0SmDS+NQVjjoLmOxWV3NFnnMUxDd8pH
YTqn9s3OUYv6m76liX+AGZQHWWKFxbdX/3Cj+jyY7JdJEev2dzbkEsLEJzzLaKnv
K1GHF3YTtNmiOZB7VWiIMBzjN7EasDWSUuqt23M+N1kW+ISJCtz6ZGEKbUlZmQC8
QT+E5XjxNQGh14ZgrScugMPjUF+JhxhtNFrcsTLmmDO0SGL6S1/7maPikqEzx5hU
No6ImJ3HA3i/WtA6qHevQSEUU4foG1BdHgeEloCooTWRgUJa2yM5uYMCHewb07s3
8gwB100lLsTgasYSqfeXxVDYrBgVpmT+kLcPAIr6m6zLbdteYP1Wpnw/BxeXn8xs
GlgPKXVP/vkR/7WzGZYq49JSc4xJPzOmiViW2iKQqBaCpx7ZToPPKH8fgV+hSZb0
kdsRIqcH8dWAVEkgc3dFgofWefllX4PnBof6H0X6UuIKh7GITqJ+GJyoecYChYeM
hkMv/U0WFAZ3mcEoKzu0xeyxjr0GWjRXxFNdpMOy4tVVC1MfY4efl7m9L9fqzh4V
xgEUQOlfsTKlKuV5AUK2UUXgKDdYbxc4QHD8LaKuqbsgMoMGQHP40B47Mc6rueUz
9NAAJ2LXaYjWdVFNRFn/Ir/FH2HXAS7/uTFS01hX+YkIan9Q3Kem3AujtMIQEhv/
6WWFbsuY4K2QQXH4+NFRBd0/puCgAjY2J+xhfCDa6LFWAZN2ryGbfToEAT9Ig6V3
Pj9ECs0RP7N3Cg1IlaytFCi12Ao3fJOrp8QLPEJJdWIIdYt0ktOHlq8e0b3ApXw3
AY7LMy7B3SsxluW40c5GQwh8PyoestMKDShBsmevq9PWY79i73HLBiulG1zt0nHr
8erdvUuilRFpUtM+3722xNIDNJMZwEcEyINMPL8YO1sgUFFIh2VUS7bc3GE0UysY
r9NvD6P2q2w2n+VBwoqmAd8oL8FqiI+ES0O7CKw9SJ+kzhsNlUiiZbnR2NtlRRzi
WWMMMakGQW+QK/5Ikn4m8IECe7A2M72tegGXob8TEFMJhUErLwOfEdfKAHzI/mmq
agzYgPsyKkaHu6APHh/5QNd+wuuJlwZgaf+Fkq3hhrQ+lXgSvSk1dbaya2PBVo6k
2C9lwPvp0qOyziuE+nbT5kUxgvxpKERISzFmRWDrjND+OYp6Xt6xDaRS7vUlbruy
JezSHo5c3k2URL99QtcOWwfoSsqw1Z6VvsF3ZJS9r0HvL5jhHkp/Y8gdpqN3e/ix
LpeVGB7BfQsCXZllY2Cfmty0yY0a5ABFJmDzMNLe41I6ahmCd40qSk6dX2oABylI
SjYCOgPi/cOYiJvPVQhcbQ+ZEkEeNxMMJQFYJt0mNYGEVxyqiPrFlvzyB/BFjgkd
2cJRfnp7Js1koFx8Rf8OOFQw4tX5fP/kkckpFeb5AaEYx2iHr/OCwkFdKIgS33eY
KNz7SRzfsQFjizTkAb0wG8RjP62r3Aw0o+z2CE7W7uBzvl5kjAaIt3IZCTg15sOe
awvDlx5ZZ79P7sLlpRikLiKI1cxlGyOjbbKhF9DP53Uae44Tl05Ijk4kpZh9cP1L
B62L94ZFXOThBjveqOfzX3QRj+bFpzwGtEzZEay2rRztP01Nn2vDTRQUng+Q/pKq
AZ3qaVZwo7jjGy56IAfFb29aMv7NqRWOhFJzZ6C8P6NJhJgELqxOiRj4bfUJV60m
CZ0hQtslAPrdrL1isR0gMgRNNtRQOKP0RyLGOcRgVxp2vCYstBCIgn1Dy0HRKLU0
HVZYAPacOO/vJKN0MLEe/IziqPzEAOexNCWJ3Pa5EyRhqHkelZKB04wu2c7pwAYl
rRYEOepHQy8vMhUySxdP/dvzJxl5t94RHN18jXPOePWHNuO2LlVeES39C22fehye
TCn8oxND7gLAKg2nmOM1j5pOPBPKFyeYzS7K9hn81D/wM3ARm7reS5IuYFtpScqn
aWZEJ5hlOx6eA/OSiHimtMv2DxTbfjTEk8AjH8pkUX9FDFNpK8Pr5JSX0ift5/rg
rqzMr1PxXm5abIbAsq1PTCbPtEui2yI0X+yyT/RSPt8PIgDr25q7yPo15GpsWNXg
FQEV7nX7vWbkuTXN9sirfDt8OaBCx5TRtf5fwzUXWx39U2y7Pa0jnuHZWB2EAUrx
B1NCnmfSYp4dNOm9j+1P8153Rm5UJilvNxAhXjSE5Hxm7+EjnTXsFtbQl6f51z3Q
YBm89+/XAcewsqnTHJIjcEDmcNAAEjx2M8tyRP7hADKKtYpDQvAnwchMfQv2YTcJ
Hgn/ojzP+l9mDZ2vq0C6MMNQJnamvH5QxvSlSa8xZkqHdXho1R/jlCicr7iLN3R/
5DmQp9RwzuvyynyOMZrOVuyOidixTp9GIH3S8lupPNvQ8BgM0csMgSr8seceDGpt
Z6rOhWcFzN78UTU6Nwq+cZs5OgEzg1hbi4ITSmTjNcgltudOOfjLiHrV3WresTdn
HZCSxkJrsx0qWTLbDUPkt6j2pHeLWO/TqOG1/8J3ZKjBTnBfjJUKTEy2GL5DkIbr
/eRzXS45lKRZyjCjyF9jffBAAVsKRkcWE8Ez3CwLINEYT6mrUYddidkZwPyoxtxY
pCgfd1ygUvwrOJ7B04juryr0zkZ6sAAqTkkVt7cI+9FPygG3Jk58QQihgR0ExPwA
ovcFIjyGYor6vbpFXK1geT5rkcP0BAgpNOg3m9AmItKmouaBI3FgBvMEiFWkKEe9
aTdJ8Bdbe06/4dNg1318WQpb5ij3xYmHQhdW+TVkbOfixtXRfOsU36oO0gq2tREW
v/irrIWH0XL9VjKSCE4iqNCxFD4iDAYn/THcaT/OBQ7II+ulIxxME6AQd0NttpfZ
nuwl9p41lmwYTD6c8cPCVoORv/go9UF6bbiqcUofd5JS4PptmcGqRSv54ptU/Eqs
aWsNjz1Tv2Z+/xNwwkGsRaRTswkTMDzuaebU9ExhW41Pp2B1jQmxpupIUYQy0fW5
f1c6CFYasrVWMyGloU0ndSJ0l4KBYOlbJmHJY5Sgn993VXwgk7f7mWWrkTzWfkhI
bRvjnnLLkYfwprjv+dILOpJ50Ki0+hkCsGbVk3w8RVm0xQjzmm1M6HjalviCGj+i
kVN9aGvwMJNT77DzMYT3iGAgxUPfLoU41kqc6lpp8S3B65F0hPfe7ic7/5/ZgDv9
bz6nwLbBtHM+kTtfBjVz3UTo/pRFsReIZmgLLJSfEnVOOTNw8Ol33sFG6fAfVTdc
PYpxhkJw1Rr9oY9M/h664h7CzT6z4PTXdMl7WMqD3lu4T1sTyFKbNGVp8Faba9lQ
Iq+VjfrgYJB6ToOvUePKv6iCy8wP3Q5QVxAzFDzSkHVShxiyhEX97iTi2hmyAEas
kORe5ZSPsydymbxLmVNLPKOAmajiU4BxrFHu0/2+OerEP7Erw9CA8dDHKeaV9tIx
+szFXCGMDeunChj5gbtLu5FUhNvrmIpglZl2D7UHYN5qxolOWmkerVtgc/Z7EjW9
LOOipZsZD+2CEHX71lQ5KrfNLK++c4/VcjGclEjIjF0R00xuWI3YkHv6j1dHyqYl
yPaJ+/9nKRt3LJYQ4XUbI5lCeOII0bXVjr+Q7eNwrAuFq5ScLSYGBPtFtPcvTuh7
LVlWnqFU4ONR9o8xFTBdiLnYuMq2hJpRo6JJwyg060fJD9jJS9E0vckEi+bes+km
g0m9zGMIsxMckm/ubjBEvAyU76ixCl4j8e45UbrhqLm7+W2t7beMyZIgjp+sajQQ
3MPxp8g7d0h6nVLdv3499c1RsWOAfM1DQMKE5VNFX/9oWh3e7UXwm3Y080cXz8V4
0f5YLnP5TUZbicCtVmbLClSFax2cIkcRVKER5ypcRvdOH+otJuHUkIygXh8hg2mp
tm6Vl3gpbV2Gxyjwhi40c5NEzLH0dDPUYmY2VGbK7AdM7eAE6UTT1fazOAYSc1Up
//c3/SRbl0bvQB659/RWo+/ryBu2R+1/epA8HMhRzNFvf7eZB1Y6nefRdR9nkiU9
KQX7/lbkyGC72ERYWGIJj+Iczrgu3XW/Fd8Z8DC2qrbR1WRO6MYT5Y10AqMeSjus
licu/YcQu/8QmW+CD26rZMdRVCReoQX6dYqblpOUSfp8FTUnJXL+9nlCrCle2vxu
kQj2sHxMPpOrAD01iq3yueSsOHv6PhknO4Gkcaf7ZBJ+htgveR2+HpbDKkzAQ+/H
OXmRmlov3nSxxZxoWrKYeB0kR7RCFvzNVEI0/KtBELWFwDMcDtEb3yW9mdF5l31F
xfhKd9TTTMBT75l6mvwe+E0yZ3Mgh13rBalQsCMVifsvhA05APJXr1o8dF7VITNr
Q4RRUMDRLxMo3lDXjJRPlkG4Z5QMhJpK+WdOz/bgYOTznlegtAYvN9C7K9ZRpdnl
aKekbHSVE3tRxC/DYQRanyRAVAUL5J18IQSzSihCR7N5jBLxjYiqcDz0/+nTw26B
/teehX6BaxHzO7fzzqQyBzz6UOq754ltTqMYoVxF6leK0qwlv3ODjUZZlavZqDm0
sWqXKLMJHOS1KlMunj5jsglqkV3XGHxY54T76leFpt49yEpgAUuBL+VbeUihGSK5
K6dVxO8aHm/oQURRZKMdvEQK9NzzB+DurWDoeEum3YrD027wYqjC/GXGPrEPn4Rd
1fWgKNDbnUBbNRxbV4gnBbOjN0vtr2xWOeWQ/WlC5zvp1x/LLX77RQPa5ywVeh83
DZf4c/c/+u63iw8wJDB8hQBAVdLjK1CN0Vpc8nfjCBSAgLNMHeh0vXT8vBM9uThE
KMHmYzXYU/NZgU38wQDhg/qyuvJ14bXzx2leDG3NPceI+PSsebWgjJR5EcFqddyj
oQdbrhEBw8t+e2e1YbR8AWerV66uMZw9Xshh0Md3GI+sDneZnaMYF/CSv+DUwsHd
7tsNfSxdYIP8O6pzA1NA+v2Y+tPERqY3Fdpiy6B4ZG0I6diXj1EvhTdzzzwiasus
q/YMHXU296Tsf78HcACTQ+bPOsjAYK+nhofJZhPFQA5Nv6ujiDTtJgEzno1GBcxP
IoLtdLDtmmVpsoulIN1TaOQiqWhKVg4i4vKzca0CB8Fw9IqFxGyhLvqsT2DyckYC
GChMuZDmjtnv3PsJF7JtgE2KkZwy7ImE48Ppo2yZI63wkK1IvZVNaDbNKq3W1X6u
SOpxRa44YpBVNO6awh6AZz+Lup4ORUy88B/S4va4nUtFQut5dS+l+ecbkbW4m/Jy
soLpUYLdnGHlhR9nmpAReMIxDDjlVtNcfjZSf5X0DuJua14//OMROf33SyfDlqr3
LttRh7kWz0hiEootXDYQTGhkUXwSbvJyqAP2UQZYzRFiyHNVcXnkAgXifpdSfL3b
x1IezNMh2LNSVikV2slITZj0PrmT7VuPvRHQAGkb6Z1Q9u+HTv1XNbHWdI1UYhbU
PC27m0A/d7SYgQs8hRqiQfnkNQMLX7RZG/BH4jN3SgcW+gdo27biosJeB8tn0u0g
XN3vk9Z8mzyrp1omQs8ssHssDp7ZT86G1hgyyKX3NRQZpJprJFMFXLg7D6n5MJMG
JE8FDRIRwDzYNu8X2b0KKUIsrkPie9QpKjSKH8lm93zmxzIL17L4g7LkjBJBi46Q
GAqOUq0X7msKI4l6Xe0BvA2ZXaxhYf2Yix6xc/8yCpa/BFdp/5dzAUkAQ7n4vkLM
WvrtSBr4DLUEF9FjgJn113vOobVQmbIYzABNphDkNwvZ8BdAWbscO3QHENmmwW7c
We1g2nBbsRFdWSqd2NJQsgE1TCkBX0uCiT0+gmqYAzD9rQkrhuhkFQOascYBTl0A
tvEu+5Rywqt5KdXvxkUBT9lBc5/GMhAEUxYm6IwhDGBI3cwBN97D3GtiNmT2zV/j
23/PwAO/EIt4RwO8+4LJHqoMHgaTtqmXTeoFY0j2998iYxb77dqdkIV4r5T+/MgG
iA4LMhAFRh/gGGDQlHPAd8yKljlNVD49xO4iwMSWz9cKJztuByT3Gociu5QPojcJ
LYnJQds1VE1oW9IBlfCz4iL0Hr/sRlB7DUQrGL0K6eqDUuTCsSkeRJ5oBq5IYvFG
IpzyHP0Dfcu3+kItpOKjtEbHrIomHAFAIXbyHKCGnODHgHy5u/0d4ABYVZsztCwy
Hh/oTnJrYSAjveq1edIoObiaKnFGO5O6lzqomTldUaskVkFQJIB59BmK2mTV7UDR
ZnDL8yrDs4p1AXD8JYVyTeoXBereCY9Ev1J7ec+E0DEDY+E41jeFxguc9LACB15E
M55/HazmkzRR48/EDJRpzaqUH7wAvUlLSEVxNBI/tV1ggK25p+4ARUkdEgjhrxF/
KGge6tIrriY7DrJUExARBAYE10L32x04D4/yNotmXt/1cR8hamH3Ch0vqJJ++4vy
SsquIVrYUACYQTCNkYmVvqFJrUevY6ii+05olTxS0Azf8deIgtJS1XGZSrz5a8sL
x4GBwf699z64Bd2RJLclhBhG9WfOjIE6cvQZ6kCMM7tq2DrT5vRgXWgAkAZY9wa6
C6l6WW4oQe66Z2n7QhVXL3YU2v68AD7lOpvEBMCFWvOP7+LCHM9pLVj9MBywbmpd
qqcEF+F77thxOwZTJKiWEbredXNopDZ2G8U2etCBObUbM0QAmNiW6AUbQwEmkAkf
B/jEL6an9kAj9ToaxNcb4VbQZO2Htn2yw6vY7yvgk1BDdGy7A9vzCJLhUUVzPuk3
r7wIHL6a3g0dFFJj6lp4xMaLP4HbcbD3FaSUbHs/v0P/ig2NXYndoPo7buBkuDYX
0gAvFby7KchJPEe13/M1t59A6K7JpOM8PlVP5EfoMjpp+kOnRsj/wWz9ZsazxlpQ
skHYllieQ8tZ32n+JcFcryMsysBCOjqs6gxEHwNyqDZJtflhoV4378N/l0quBFvB
L8YiCMyrtu02Qzu8FG82Krfh/lgbN8CPYyYdJ6LyiL9n3FTuHq4dWMIKz9pi1Kqn
lIT31v3Yz7PSHFwbDI3Qa5lYZaX4d62JAGbhV1GU2udnu8NVMuxbWzlW/wz8xK8P
QA4M4i5e9CSuN4k8ZVOKuXfTzaJEaLa1nz8cEj1O8DMORXPWbntsqbQ7HgN0YNAk
pscEHXFJRwp1ovFuf/n78K/wEOAgeolVzBCY+66OiKuBDA+iJxWEnvZJf9eyDaxi
qpyj0gPV0ks8cYoQ16d2X9uCpkpyjk0VR3kLATDWgx9RQgufRy79+tvG0t7EGW0w
OuWsarnghIE8c9FAn2JkEFrtvFxJ08ig7Sp2ski5v37a2hzixDVVN5eVtMsHCzx8
GkKYj2ygHJjNvR+8cVPPYwVpfuBecz7MMlWxwEbt4CacXP99Ay7kBSM4tEOrSlE0
ZRIpYHpPTGrTrna4Cd+/leTyyyDzkh/Bfk1qu/WPUiHVPalJas9xsS+b+einTTcE
LVyWnrX17c7oE/2ZfuhtvntvUMlCg21E+mJZTRPWs+j43+B26YR3xwIL0T3EUTrd
bxLsG5C/Om3kHG+e4axbDrJyMgnEITbuELBX3cqS37vV4YRo+falDIApGC1Fiii2
bAlbHQ6eNkYBjhwjnrjAqpCUJmeGzMNIn2uKlhptLNzYhYb9grTnu3BM6gfh0AYp
G/lqeLg1z4nLmfbSArbzOuNilSnWmBcl1GSM2I/N0WnOXZUu+hOODi/hatEtP9h4
qBG9qmn7ajAe6+ytwsFscsXIIkdYqSdab14MtGOU8bHuHDlHrMWb+hOi7a/+lNr/
UtHBM7nB/hYU5JEQgaFzSy0EY8aLtiz2Y1lohgi236HhhQ2qfgVVKTpKp9gbvVUW
+yiBfIVWEAwOi3LdEY4FdcLzjLimMxaeEc1JE4yDgmxbLXs5hVCmhqdVAbIAlPC6
BMDQqSLenl5AyMTGcCpohXWmK9yoB7RU0vZEnVa2d/z/ATkGN8g+4mgOWwDVa4Av
hUx6kEqLTOhsjjGqosrdg9+ZYitrMbzGbQfJzkQJpppAwWSaz7usacVnRyuypkF4
8Op21KMN6ohOODp0+FgVMhjV1KfR9NsjGT+rxvouxOc7QxM3ep6ObGOsUXRBoIi4
TOpIz7igb1ZolCyjJVgP7/YNH07f0VMUoXkzgPADqUZl8oY/kHWRWoIGHpaMhJqv
51lWvmlq5azHj3wTDKcoW1j4dOrnmAugjg2hjEV6Vgdbo/CkDmYdC0AZ0QEAmMbk
JH7Vi15RLZBqWwsFmx+zAoRl58L107w1BXq0ACVOgfTTPYaWN9seX6My8ysWIq6Y
QYjYadZkWrc9wlPYoexJcY9tUJMbMYkqKyeqwpQ1gQp83d9ljAAQ8wRVFu7Zfv/B
6AvIroUIjeV2gXjgRaXke0Su3vTiLRwWScnrcffp67zLKrrz5Bx4gYgpuGfQD6af
UTEU5Pt3315smcfKmt0ZvgZr9dv/26J1eOhUibPbSfW6krzZErg4UVWKImVuR3G0
QItUyaPfUIWuQoD9u/xzLo1M5Xsw5k/BzaVBpo64bi8OxtlYlGx4OaJaL/2LEBPh
IV5HIVwQdaVcGmwkf1lvt5p88J0eNqFhuNdsc9ssbdOI5oNDV7zFKTwjCIolnHiD
EvEkBm5oRzMEJWXFo3DFfXtNOBxj8z6oQI9WcCPK3bhVgG6QZ3zZGQ73NvvtBeBg
X9se21798AsmF+Q2ISbWTW/tTZ5oVscQ0OHFXYqPiRvymyd9MO1lT2tYY3NRqWVR
nMvTQleb9YD5UTWwkMVngV2sA4H9z1sCDH3eUCGGJKbZtR0gpSonzFYJby0bQUQZ
z1PdNmvKu1Th8JPs5ris8YDPzkmFPBdZXB39/4ERkIi7vMfzq8/gVb4KOPjGl8qj
XZBKBAh+sc4KFrpMbBmimQWV7b17n9WlQWtI3zH9mX4NMy1hYb5YMcQ8QVdJQw8j
Rz9QBRTT86DTVLRL57+5oCW9vkHQT0ieEmM37jKETvpTfONNcfCgH8seM4VqWeA2
0pclAp+TmD+XQw6I6J/r7UP2zLjRuGVuj1kw5ZRcPeFlPFoW6O3YCIrudCrnTuZx
74bnDpLsUxzgCu6eslohaZxPJnJk+EA+5GirF1Uf9015ymAI6ZT5ZjuqOTlSX4CJ
NkG6nM3Urx+cKWwQ7T8laAWc+dJEH16Z4BBsZxJW+O4KX/nd0JcdaUEqMG9Nx+eY
uHoQ1b+oPHmB3EZOpOz8VByhH/SPuNuq86Jht1vlRQOazXDanxtstEUPh97+HwXr
mqiliaOrDdomYmfo4YAeEy+Gk2yaV3Rc+ks011dwqgNTv/4O8H/x8mAnuR2FxS1R
NBDiCGg4swwGZ+kObkvlP6u5Nq9APl69wWhSoZHx0EYLJtX90Hnr9cPlRn+j+/LX
ErA16whx7SgOtpDwe6vJzfhlt5unZSOb0TpG++99DSjIxlLCgo+HkQF958QIJFbN
A6FoR1ZXTiIhQzOoW6S2u0Zkn8RuqC+VpbukLfHiNon4q8jDdh5tpgsIhA5aPCT8
D+ixGMhfBFyJGOqaY51wncpKkh/o6j38/OBOr8DWbmgJWlN3YW6ZyUtoiiCxgTE2
7dDSzZl+Rz9q9oCEjOawuatZCgB/fglDIHRiYws/5dxemlkcAPw/6g0x1fmIPzT/
ocsyCe1EvgPWQ1rG6WOpzZLCmtvKjoGYzCzCDDkdTw4r5QXI3yeW4MmrRPxFpW/Y
esWJ9YpzIIOasTstLgmj9ytevfGkBcJ7NMcWX/VBapEiO4Ou343rswu2hU0sYfZi
Czrn6bRZCmfQ+1wtRLCvVFE3ogefDclzYTp4FgGphmsdm31k4TYYfMI0cRsul5l2
EWzCPAg+a2CpmHwJ8qDugKkHg9eBarPBynP42oiXlMGTO1d+ZTi7w8sTuBWRbQhv
0yKstn2lTnCtPMlqNAyvfLE9dzNo3XFjnd3HIFhNXuaihyrQXE2zZtklKDRnaSFs
nuxVkxwMJwKniRPGFnhfJ/GTTqVw8eXW/QJpy3PK82Z3z9KwXIxgHuNU2zyowIE0
jF99desCxqNT/8ZfVcqw3OjQXt69jrkBEalL81XaugMh81nAKM/VAmvVqcSsLpeO
T7tKZ2s75iNY0/6nWkDQnrd2xNnG2d6fhnbg/A5+eK0PVwUNbawfAOKCgJeOgA2i
YtAiEMu6mdHDInv0w6TDXfQ9kcGdxOjsuAVar5LTJh6PZ1nLwU63FB22vD9MMewf
y6iMgwbFvEnASwzvbLtcpTVmdDkXLIzrs+gI7Kw8vgpUQJi1laj+JifCPvm/7g1n
sUl4ZW4cW76bbl75Qy2ofdLgy/t6LbLQijLRjU+GPUg8sCL74TP5xlaJANlM8WUW
vKyhNvXXZzkvBe2cuKDUhgHEQYxn2orODJEgFZeWOR7nvKIs7GnBVLkWXAwnYAdp
C1o/AZYloUltZKIMfD5vBV4hkUFPNZ8ZabaaGXyoG5gFY0+fNG5hiEQVmRrgt/Cr
bl6TNiEbDAC/GHyKavvyqN/2cyIrC3A2vckymmN7zdAGfxNK2pjGdCVHKIkqAMIB
heYstMw2rFidLJ77+kCEgHkZ+xbGJH1zWPK9p5IHOJ9e2QHN9UOUnv15LodGd/7X
62jKmPKf6rwnxD7qsevVevVPPVTYdEhtZ5gy5jn+1SchtFzmv3UgoRrxcune5Lq5
Mp0sVwjYveXCZ8AnCxbL/3SF3TJ2201pGozTdp25HygZyuzT80fugbTNQL8vxPx9
tC0b317OtYG9XocUcVZAg0Y2lx/iirsFWQjCuEOEDCQVS8k8kzPcFSOjb+iRMQJt
tCm7rbGCl41CJtFvoayutWYB+SMW6r+38pgltj3HGmunIdMtMhlsZrNZs89bbzSw
6O6bDl9quZdBhGmh0AS0EcfNHU7IoHcby9WGmzBzwMHV2AplxDQlG+Y/AHEC3FmO
lIIBAqdl/ZFegI3pYhiD0+kyacpXJw+DS1aZnBMJVFX1nFlVPDS1A4UcAD9FepgI
DI1OXGlHTlOBQXpXORvw4bM/nRpemZVcOkIkRUNSMWbGAcRXNDxIpGnsPhw4VEaY
WlfDGDN2WKb0ddaOzWslIfgcnhPIQr9bbEkUMFT4FEUKvsuk0Ge8fuZAwA5zUssh
IHR4Yv6+SMYefRYmANOluRW0kdrreBSTi64I8h+oPlkcd6Nav09FdWnB1ncI2lL8
DIQeGjMpEo8mCAG37K5P7vqVzQVoNEuEnGZ4DSZuLbrUPv8MRXAELbKwY9hhxlh4
atXsVuhNgGCu6mMYTgKdRvnGJu0ZLZZ/hGCi7TuRC115g/H8SghcDVTWy8fAtpRH
fiJtOlLO2zs6Idt0GRf+TbwWCtaQZX7o3y4UZ3RYuxK1DOkM7T4XB83/RW+Yk04D
2M4f+Ev+s0wANQg3gvW53t2OdngZAn8fHUF3/AWp4deWm/kMRpZixJCxkbXY0w6J
jqFEA6PY3Al/f6iEAVVEZeBr5vwp1SRg7blVJBMTAjnZ7Hu3gw4Qp0w+MeLyjSZh
c3zNMMDZCgMu/fz2/M+aLx0q15JCJwrHPPTfGnS6wyhZuU61cVWOPFCfqF/VYAnq
l3OuqvpAJxyCA5Z2qK7NlzsnuE4ocKMtHu0sszjDldQUl8gWJ8LwO9KV4HCvt6f6
vYR0DcBxlaQpd3oF0PiAXfXygdBBbIMEZ46FF/c484e//qcX76q0PUIEDVot9tGq
epVVKwrG4KEt9D2EvxP3XEXSKPCdKLh6BIKELC9gFE20YRYXtW8I1vhltUAt/F8C
18uMzo6Iddgx2+GqBr0TF7iavbcXJDCaXGNkwbfG0fQcdhBJx3ECvJgT7YmBsuhQ
mhZNqbceStZOPj5g3v22G0uXDRDq3GmMlnZyVALDfdDgrJbHCoIvU8BR1vqPTHwh
EHwq9JRnrc/g0cnExLKTHrhVrvnHJs+mp6xF3OCOkoy8xKxlfBFmNgC0DamTeKfV
faBlW/ysazt1RunB/jF8ZBP7EK7yRKsRAoOrGiTYBc9Ojkb6JJqpP9cX6Py7wFl2
9FnsADEc87kzo3pensagQkeYJtnM2uCK4+odPgLnRBiW9D6YDDEf6lIlo8bjJtDT
/ugXKrKwyFx1IiJpHQTG4QudFTS0/OLBqnY/Kgr1yRbAnNoIzwMX7SjgkMOv66l8
ZV2PzTFI0FLwLfBjcHiUjBO3cZwy+i+MDmbhKwIku59dewLVtcGS0kdwpXmG8CP5
k8xOuiJvhevQHvAX2yEV9IidaK4BIl9c+J9ET2KdoJX+Ay1BLR3YlD/+ain2f60O
CvUcuw4Z6Wh9NyXoYebCVWr4sjKUcilAYbT0IB3/W1QUb3Qy3iA9crzxuAVNfA/a
BxH4ywWOdmxp9LPWfZF7mPDC8D1yZS31UIrsal/t57IlDi1j1bluzUTSBWhiAouC
lAyY/yrPOMBFq9XzujrxxEkCEzf+JBCnAmBJFbi11tLX2ARwTYXKrhCmyXiVH7bv
z9nDRLZ612DomwXe6KQg1P50vA9luP+8L1/XEHpQHhfc5K/YX5w1xeWjLSENw99U
XiLcDXa2Uit8ENvPA0HNezLdDKdEdAO174zev1SUW3hsRn0oUYImRNbtDEg/vTtw
ypfw+FH9T93fYlNAMKezGxAHtJZ/gu87nfvtAxqGNP9F/tjOjC+sx4OkMDpt4U07
izEceUUT5tTZ05hpWKjFRvNAHynSjsrJgtbIEil2Ua5mVZYFqr9i6SePqhmCcVjH
ucjXAZvLcdbp9AFJrBF5MWuNzXWS8E9m/9e6wy0z6MA6ODvt4qcrOVUgQwFy7eA2
d09UnuoAnVOHT72cNoVlcUT5vBc4XeZ00HP2E8idM+kTRxZtlEZNZ5GZ26AU0kqy
FIu9wzynGW/Gle/lsWhCxdFq/N71DzOsPfpbCbYivqoJpw/y+VFEjwKN+S8g6a9V
Gy+ekchwFN0oGGhDZwJBv5neFQEb/reWnrXn2AQ3epLAKpu5g5xMmqgOqvaZ44wt
PFW61DHCetpr0jgwj1j/CRRTCHCkx66h0KUMqhFV4E3FdjXn2woP058bTaz44HCO
ndkymzFt5v/0gU4GF1YvF7uJTjCVQbtPwvXbw/pUgwK5U0YY9BT3oNnQJcvdr6h5
YvRVjvYLb061FkHiNskJwjRu/oOsNY3HTCN087cJANAtDPR87nXROJrG1+LMeMCP
qsQcK6tu4y/2/3i9A9oheJXfOzlHVUz9pz+DgoHPLBLa/g7g9ylyTFh1qtgjx/k4
WTdR2hld2S6S7JYP+oq7pJAiZTO2keCepPWammzIgg57M3U+fc5FIyauw46oi9g4
RlXrozjL5p9GumzNgkKwKssG8XInR7hDGH6K1knjj16IlvZ8PEFVly5NmuejuJgT
IMtMMPrebPXqggLPJoLtd99l+B3RFfWwGNCTpK2Oki2g2XsM3inAL1V0Q9s6YwW4
nLdV+m+1KLPYq7CHP7W8mWd5j3/I3Ka7v2iVek9dDLabqFui65vLQGFSkUwqpf3u
d8/+HFGupIp4gUnw5sjVsXkSTz4RP6GrJmVpYdZ2aHeRhsSoo0VZqIfwkMSVYDSx
CPWDQ4NLYeJ8y1rCrTMV0jQZ+gBvumPm1QzhR+XE0zMeHd3MYM5FtKldtpIT1fwh
WKzEsE3dtZvQmasQwrqDBgDUugLG0MDdkmofq4l35BNxjd1nrSFiR2GGJ4X6loAL
QZhyrwPLc0qXU84/kz0ejB2jCNfUhBvsbh/rt6iKBnfa+WP+l9K9kK0ERjxDZDyK
z2wESbYLuoHtELMoF6dLBMh/u8ytbxITFR/ss1bs7nBv/BE2pz1lfJBrfb0sMLaa
AG19A/InrTLt+0e+ceBDRKBt0CswXn0oMu66h3y9nY5f9LUaclHtqNmp7ZaRh7Ty
5Tw+PYCy8rr+jjGw2bW7nKr8u+R2Suq5xOr6JF0gBwl2YFWKvsFHNgWkv6aU4Ij3
vGBcH5gDigX+3bx5Q8GqFMGOqBT0Uvbzu91fn7Vsfiqr2wygNAYWZKBQ5DdQ6lDM
mafmTWniQBUrIwaKf+fvSBZC88ApSvGjvCDysAMFpaSXXVbokf/teegyFatVDtWF
PAe+LupPtVOje5NAwRzPIxg9K/74OD8w69jv6jt/sJYJfjh0YvvqAp0ZUw7txtye
Qlxr6ciiJOPKEqwu9CFDQnfX0ao47EvR4Hlyv05sce9Zlgpmqu1r5Paz7XNZif/I
tS5fAS3WekirupppbofWA7MAOpWNRgAeatg762uoA4NosNSAeb50Sv+UO+XxKEjC
91QcIV2CxqZPr0Ypnh+NjrWhptNREfOuxrLJr4LKGUjE50NcqtN9dMzjEJosGW13
3k9CX7lP2hcg0zTAU3OrWmm+dwj/wfewOdn1COVj9BVTm90LnYjk69G06/cjyHgv
+un/L5RFy+rgD4+5FWN8/ES8z/MCGZ16N4AdP9jIn/mm/usS7RQXSDfQ8heQegFV
TjLdX7kNEF26I2Z4EeqZDQ3nMa92gtkA1O5QTgApvt/eVB6VCVzY2kNgSy82R5U7
f4BuIKso6G8VU9O0R4oueq75ZCa4V5x5E6Tp4rulPLHexaIksPaBZOMsEgUCCak6
QafA4RZKztACX1VXKOlyQj9YJUeY3ytbxialpxMqNlL9WaQ4k0Sl8w8jXDpgHT7h
O9RdNWZb7ZtxCBlUIrM8pxCCr9cDvCqEMmE+6krQsstGkkwEhMKBG1H+c0Nycd+l
ADtXiGaWF+FezF5MxDU7foTFfrZhB59ka3w17/f2QWIFmlJS8Bn+Ce9DEvcetfis
Y1kZo+m9igjesjZkgXjQ6yXFUzsU8VeCXt3hfMo/+m6sH7Ez5EXufolVUyF8jVPP
3yrMV03QBdmTcgdyQO0c47GW5Eugv1pO+dvhUv4pNLrCDGiPVMFU3CG243GW0biR
Mnaz5tK0Att5tBpie6WJX/MGx+KpH8WwOGTwjzXe6x2zFbxjM8NrlvLDa0vPoFTd
+Xuo+HW39Mj+2q0LHHEyaWuhtHKjZCqtahrq7+uf0aZP2ABLhVXq9tRvHkuordfU
BW7ZDUzRHlrLTg0SD1CwtRvHCFWjkFD6jLBMnlgL1G8yhd0gYE1MQ8HEJBKqNxdH
XjUfQvKQWsh2FVK+HDPVoyrh1kJq022XkDowT27q546kxdf1Pj00ZHmAc8HmtfAY
L6OObwA2yDtmuVV3WmP6GM9gTvbt8AehzCo7tqV9jUH56RC82JSfGFFFMrwWTA4l
8ZzsXtA45azlsLBtByYUlJrP/tmKPfX+kFcnIk/4teLnF7ufP+2TrwvAU83GZM1G
8rZ5m5j50WgOy9PQtavY3p4/1C7SHvzRfMhQk4x9qRUfyk9iP9XRIk4ghB44mdg/
P27iVpBsKg/HnSZAhjTLQ8h2iZHCS7Jt4OHkHeZRvOvhkyUqeypcmuVWSbWd+aUK
x9E0b0/8jCDjFTIjDzmPgb82Cayw/GGvyA58NwB9dpX7SFOXpgEWwSMBk1XkZMe8
9TbGRLWDrfEDMalyzKG7C7DTNP9dkomqlJ2Gydi0uUn1sHjyBQSo9vzTSfTchFnW
rTJ0wZfsk6NYKacws2EH/WpLjzdwySVI9nbGMXLEIBD24//u6MaheQxs+KibndWC
h2+HQIRST4MG9mDLhoCWISIvv2s4FAAxyk1fTRsfONZKdTEhj4u0iCUVyjQ/LlNl
poRD+Qgkt2eCE5kC3vWKSsJMxNDf6C3nnJl5t/QWvvnTlwMUWOHDUK4PYKFJVw8w
2DaFFYL0I/EgMCuz/YRBeVLMX3aDV+VYdAVo9NnvgmySfHAlAOAC+S5om0DxQp8m
fJHl4A7I65QGeZ7R7bju2YAQqhVyabrm/jQJQ+FyDJWJgQCxkdBxE2f9Twc79ZWc
NPL6EFLi4TFZsO09EKBPSXsz8c5G/DhNXmtNSTXBVzo/HhyNsLhPB41ccFHOpD+C
o2O4tXD3oN2NlBjpyw4BwAazJkggFn0+INnOQM/ShQzAoB2LAphN4eFX1W8hsSMA
clbhO1GuHMWr1Yflf97PyEQ8q04t5ml1Jz/Bj+nPaUycuyoNL3cB3g1n/jOxvlly
XA7n+Dat/byJDR5+JEOhxW/MRDjAwT1PIcx4adeWB7XKQbk6fIWgeu1iSedqpyuv
meQG/qh62SmMZwHdzKiTkTow4UGT4AYp0r1y2EorjCM8tFO8RgKBICxiGiAiNsE7
+/h84v39ZcTDAb+IFfsBuvfrdEr16q0LEAfMPuReNrxoucQ6mxoZlUK5toIXyfqD
E7tk7BBQrHDxeYCzBjB8HlPRsZYp7eGfOOVdE66F8UXct6tX5YmwZfqu2Xch7UZ0
MjSgLq83TZzpXsOksjecy6QMfvM2HT6VGhN4PrU6V1iG9oMzltEduZVOj+q8pq2D
dQ4+x6f08NlJ+QY1aS2nC3FtQnH5av3H7yG/4lwHZlJILk/lliVsl/36KJ1nqfva
/0B1Kq0pD4AtQU/vT6hV+kQFsN+ZV/WrSbhADFkBSZM12VXhgpL0id2q/CPGFFFZ
ODnTuXc8UMfZHaTkNJMfaf76JUl/kLUEoTrtzfjmTQg3XcaW7MIBmKLXt25B28EF
W3O3ANpO5E7oGoMUzxR44kGTQttCtTPROTeKX1Uui8/+L81iLpl7j4vFcCLNAe8o
hhYRvuaKvzNUoixFq8DOLIBU43uaYyxv/JvoCJY5KoSJM5w1ZeiOdse0YenS8j6L
IuxIHJ+JdGPZZcDC/lFzOk+V9btRsITTr+24QqfMYTtA99oMfT4gKaLvc6ftI4fo
Pdgpgpb/Q+dvdwG/Ad5zy/kaEov8n5vCkHBeLTUkzEe+zaza4alXxBAk/ikIjFiR
qgFej0muDZenfroddLhC6yt5TXOO9MgdbnF1guAucalJzy5oLM67Aw/JpsESDSO8
wyf2nckibAVEyjafbhf3WiTxGUUVhl0FTBLvsQZniaTkS778/AuUfzDeHiQr47MD
uBttqnHmRc9n7i95Vot/173FHtk+yaPVyccVUuztB6wfzHEpx/YwQjipXAYQGIRt
GSFAT7gU6KITyIE1EJAnlzUibVtK7ZrO76hQBRx3tyvAjSEfqx/EdIpO+5nnf9+E
EoYbSiI45B/xQgjKsepiZTAivbCApnwXI4nCI/07KF3zya21oRBUVOhVAYUW4ul0
WHvawP4mq61vPvnSjET2xJsCb/YSrbY9xQ6WEb2aKnXePQzJNYdlMWR9EBrlkJoh
ra4N6JI6TGbLwRTJuzWYagh6G+OsRFDC6Nob4JyMiSNZEho3z0w2VOexog7lKy+S
alSU0hVVNa45Iosz10U7QjZODXDhK75w/V4fuNge3UwABMKL/6tvqaVFrS6BHMJe
mUqP2UwtwXQfm7sQruhZ+Z4K2nqOvgQ3bA5mqVuajWlbL+7RF0S45adc0uhDVORi
TyRJUbJ0js7b9c/beh0ixGwefSUyY894TspKTCy+V/6+zbwUNAgW1HNgmQzvkf0J
e4uJA8S2SCWfpVXx/I6hscBx32KY1VEQVwRNU4uB5en75TFTaq0TWTDiLfFxtFxF
YNNBcKoLItJH24HOWC3fAfPjoPXHyeFwPZa/x/YoYqXN0B16pOsl1tjCT+immGUd
TPwy8J2rnQTFNuhgXbzn9cg+vwRdwbGwX7IYLr4sYwG6MEnITrMvBSpu/k7Hwtv6
kxqIgtoSYiOYa1NGpwnoThCyTxzfMFVCIlhg0kfq1HI2cZvkqPMY/oq6A2/lISRT
FgnGjgSfELvvk9aifTWXcWq0kBxsDjkPSNmOEbl5K1QZfoPwNofCdxOaFulj4zr0
K3GJFcHSmkLuv0kAVCzimR1b1ZoJYhTQCmE40ZI5eYQ7YOx9kHl20m1p9LE2M5vf
CFS0wGW9/WMwpBaWJh76JVqgvu+sT4WlnPCS6zQbTrVYZeV74bpGWxWKqQ6OSn5b
2g2d0MfzDZr0uHKgkFVFuodMhSRvY7li27CN35na417zuf8M8UROLd8pBTIXwXAH
Yh8cGt5NCDxrC0h5K4KzRPohAtmr7fei1WdrOAjm2S53d7UgvpbSIdPrQzMp5Xmp
SyH8PvjVox4VqrcpIxgC4SvcmiKBByIeqTmSNuS6lmnIzH6Rem2sEb+fwinBXu/5
WwCtW3ltMgZfDfXcQgHS/ujPvV4X0cOMB/stiYkceK/iRVL+5kQkQtbeWXWPsqfH
lpgM0ZeJkybCgsLlTdhovSG44//Roi5d3do8+WrtguWXeNbwY8BR9gC3vcUffl5L
Rccjk0pavnnA40Sfy1Kgyol12NtlhTKrbTVX110NlfwwVIElHXpFXF1ruQUan7sP
Ref3uv19Sf2V74ZmBEA4IFdSKhxBNME7iaV45MTfcd5zkokEjC4276qL+pO4aK1E
39tid2+tRJmac+Sjnto4mqd4prQozqOsq+JMGZhMoSQBwUat/Xsj5YGQfjhsBVh1
GhU8DVQ/nmotqrlmwiy71sITrOwH/Et57ltSZXaGNw+Q2c79teyw6J/TbbgrMtEF
5vMBDSjLScGCQ7AkS24fZU+hD32iR/1S9N4hnS1AGMDx1vganycyNOfoalvu0Rhl
0LYoyyeUyF9VnjA4RkbGNgjL+M8s+TGFDryh7CVjXV6lQDMwKcdfTfz+0byMnUye
coU+vOhlPvZIfyFBgjtMYthekwbGrwdrhlPiBkc6F/eJJ3JL8Bxf5D/3nvU2zncZ
HpUipo4+iD74N7H/DvEFQC/pWroMYwo9cgPEdcydGI1AZHHV+cGskUKT8wftgoVE
2tuR7HnlUOiuoe8Pv/mbCUpjF9Yo2HxYpteAMlO1XV+w2y/53YBZJ7dA414B3StY
6UBGRvNGgiorf5waeugB7WEDqjGsFD13aE8SGhDeNKKe87Nex+GZzeR76aLrDUh2
P+wyPsAvEp7sXW7yStgiMdh3Nwa9U1e8KZ493RfwBOumx3+83STiOO7r/5DqgGys
msRErdqefua/Xkzd9WYBGoN5UQRZTh0L2dNZTs2WOWY2P8/EuPe8e5y6Wr5erWPC
Vfffj5YJRqrEOsUTA+SXOpXVFpgo4rTVe+wb7lz8letZjrwMjrYCZ5xmS/YoXZE9
pTPwz1lqVOAhGJDbCVahsAdsBW0yCT/b36wiL8xfBdUfvDlMkrQtuEWFEpKAyYhx
2WfO6Z5VSkr1nP/XaPjKQNftlDO/kEjnWS8SsKp9vIdVeDxghFHXEnWWt+bMNoZ7
qYJ+k5csKMYwNgcff0+7o4/iU9umv5dO/3bqdnXtHtkefOTJeFchodhstVybf+Ya
/JovaHNkllRohOoNEw+UpbBFW7FntAAD6BExju/4uh8l5GTmOq2Zr3+O09oVxkB9
akHapj/x/ze06KWk6pR+KLz74i6SknnWxnfQtHsb+FiOBbAbQlF1O8/IuO911qHW
O4puDHUpPsuzJJIliUr1IfnpD+YYD3+oglNilyn8e/XW2bV0WtjiW69Kk8G5hGmS
nzk8mHokI6pCSGm+AyQJ7sMDdynHknGTFOObzHt7BmCXdj+hIOwk+AaRy98Phrt9
jzblVzezZpmE/XeGvwFq65hZRIy4+50ZNCBWMTV7vqelz2riDJJ7L/tPZxATM3z0
P4xl/dhwz+mBOs63gVd0X/t40HwSw5hMs3UOU1UkcacvcTBJrcgIlOuY1UJxL5zs
Vcj15eaXbVocD89fk68wSDvVR6foIFvdySLs8qrWgB2if1QNAsF9z8pJfQsU3jqG
EVHM9F/vNMfYnnwL1E3+AMzPBJEaLumuBIuYgqNYIW7zE2CN2Mer9Tz7Zj9GBVsC
MFFDggVVoWz6kGcejtrF0CAkv2GAGgz2uubmFMFrKEh10zYjcCQ/U4+WL2ZdQAJP
fTEywKLuQMhDRwIgDUct5dbH+OI6mMkWF2022iqrHy/YN7uLqEROoW2gypZhyv1L
h5FE+1GuF9ipA8xRYjQJOFivfW243uiirwRhBRSLPYWxjK2vK5sugZEzOq7NAaH8
w31VDyIh7E7SuSJAHmiNE/NTrtd9MITr2D2vDEhiUB3qNGou4r+L5IQLiZFJls8r
sMahw+X9oaQmeEEBD/aqPZpzxjr+Cz9tjJFVuRjguavvX+UY8oiUvbxKo6mAXSs5
vZnu9pOJ6Z74V9dY67e6ZCJLsioORkfLhwmn7heQuxxAZYGiHU4TZ2gl/os71b5P
ztVrUpz2rJbCYzVDR3NwM+9GCJSWQgW5/aUysPk3lkiQpbeRg4IKNN/SszuUjR+w
yHf1MlXR+SeF7ydNe8bcXf2ul40yx9hN6ThP+A0eO4blvzIMtzi5YFyWCI+qlMdI
RWCEPTwvRjR5Q0+5O7P5YFfliv/s7Ikb09e/AGD8J1q3wTj4X9YKzhBaKr17eFkq
EUFDUTF6reErmGIA5jB2l4Jju+qf4RgOii/ak8fOgHOyF+8r1YtYsPvooQmOmPlR
pdht5iVp3BLOqoh5ciNxeWx13hPzPQuF6NG2lsg0OxDKNNwDpTd696CcWkzj4OJq
xMtjtFE5CZumwfiJ/1u1CgDo+3BSvzlXnLsZnT9TsVbppyglN6YZ0d0WkH2u+id0
Oop6we8Veug2poXJuT+JdjR+OTsJTs+vOwicu0RTIwBCpl9E9bk8/87iL1jb9DFA
W+DgzmGHtl/GXy8TDnF0FXvVuKX9WvUERVkeFjeEmQT1JG5ECyBdCKCVHC8VBhIe
7/MflLf9Zf2PJSF6S8YXMtDprSXUMl32trQyXJDnHuxtkbZywuO2xsoOli8C4ov3
ufuOpoVipa9KOSnucsQcZp0sNdQFTNIVFNwgHQW2TxJaF5Bmm6yWzLJRczR6Hj1q
YJUwUpO3olkKhjlW806wbP7EoHy1s5w8bsz3vPfpCMB+j/kJxhAh5uA2TyemzmCZ
ZFps5rEVTPge/el0wtebyawHvJvBWIJgwvon76VMkXJVrPo4+iT4/pRtp43rQQ+1
ULX7VcWr5ml1NumneAgioboSp3dNr3Bb1Ob90ie6CcuCGe7HGhu5It1kkU+TuIWJ
Z1D90NAju6AmkVvMWDO6om4O2uzwD4G895aM7ePzMHu5HLV5tS+VpgEgMvsN0xEw
kp0urgrc7AO1xDT3m7XQJX6vOz4hbUtdn21wUkjRLBjMn5EicqxcOb9ToHZp/QB2
XNkV0guxiV6m6nfxEyMUOH5UgrPcxzK+4eOGx5PyjARtGc83gj1rsM7JEUzLT5lI
2EVN8bJArDK1wxIj0lcZpg6v+qONf+tojc1ANc9ZB+cKPiy+vyOcVFn811mX515J
jgC/YOBp4/dxCSo3hjgSTGgsJ4h4UkfCSKdg8fOR+V5WbWy9Zg3O2e0F2hZMR10S
wltsE8ZPM5PFxmloqBOb8uxzXzi7/SCOSVk7tUExTjo1F+ZC4DG5esuScTusy/Lj
vJpnuwLkihHhPtti00loSnJtCxBlRYJ/5WzfIpDOJ+Qx9tEa8z2JkXskd0lpFxue
sDkNsT52DYVBkGgqFfgmp8/1K5fwQbkn83m1oV/Q81OyppP4OGRJGKKmckydehr7
xcjw9FGxcUPMaFV8mLESCbKaYchSPhz9DzU29bQKkFrFF89Z+/Tg6rPBToNbkzx4
6f4cOTxy1h3swuv6gXeXcIICaxv5APA7Dn2xeOu/1XUz6c9SE5Z8/Jksy9sFMXcZ
EzfZUlQz+eSZKxGWqso/F7hzVs9RAU8DPhCu1MldqsJM5Zm3uupN8awYkeX9rPpl
6nmopHQHuMKUe9E1MIA3P89CTKxXMlHYVh69vFqdOJ16lY7V1Ae6GBDl8bArAGC7
J7qOxze+jbzWAEg+CYWJ4gpEQzEc0u21ges61Vf3Cb6wA3vWJ3JwBQo1qLLMpNoT
zGPAmgyPlXB6FsNBfZenxlLWGzlfOOU4sjykWJX4jYW+eVRJ0k9WFIgidQV0R802
nxPCITNXMia39mnt7AhJ+X3EAq9mdNBMT+aqtNjzuaqiyNZNur2YIlEiZyJtNJz0
98HnFIOWc7vuZwe5nugZ3leeDib0w1Yk5Zx0BWWh5O//vGQo7jGBw1M0wTEsSMgo
rKMnXbDgZSginJICjkMjc36xnh7qVFBlHfd/Kx9kaU0tS6BPuT2RaUiffv75+sOF
BhQx1zgkghCKvK8IcapvK9xEfHnoNd9KcsvKtNtct00eRGgAih7uhCkfIGmk/dCJ
KPw2iltLNAUpfmGqUlQrwhBm+MVT1oprPyGDGC4hHgESSVBNEi5djLGhrmFu9TNZ
dDgseeJxdVKnFzkdo0jZ47TI+KFcs6HlUYk0djS9w40gKTZv6lryxscy0hbTTINI
v+iH6qN6CwWugFr7kWfXEb28izMbIwNissmqGds9cYUfJwMU91y1gJNwTdgSephh
5DKgCEy4YYJ9AipPzAZ5Czm55ZTKb73mEI90+NQNqtlLiNIkwhOut/sbD76JPj2u
ajxMpNk2NMhYRBOmdeNcvTHwMHr0Tg487/oJymloT+tEqww7IJC6hizkX5Dpq+d8
0PlAdnoH/ftIb8YE7CpsI7+V2mD+wMp2gkfwEfTSAeoOe/B+33QJZAtSq7tcfjsN
LQ96M/IRCmVLHQJEsTMy884Ax9oo5JCThP9aaJ5xE73vrm64hgCoMbZ2J55RF+Dr
Il9ymrSC4GRcCRTFSOnN72j1nDdgLa8EkDB5s5IPf6g59t7h/cYXMPjA7NuSj98w
gAoW6TbnROWxnwlLL2ArFOE2Q6FVUOeGfL6pGalnd1dCnlwr/Df2Z0/ZsUE8JNrb
mGdBPBj+2dh/Ps0b3tMcQOiT71jzHvs40Vxbnyyc/fUi46u2qfZh9mMbwXQ3Toxb
VlyzYpnNp/UZCeG7B0sXvKziDfb2bXgQ3urDvcbU6WqjBDrGeyiGo+d4+KBGGZdY
KKB0f+gGc6hiDboFbeEE4AtIdxfUIeB1d29yzkvihtsGYZJ+tCTwbFMYyiwcexeQ
J+O3gMSHvr19ee0jDsRm+cQ8rszeYiZEGK1m3elge3gN+GOGm8RUuYblEJ2AbXd6
Oti68HpO+HBEJSVVotQgTAFGly4snD3v1UrKxZDv4IDH3gv7yikFUc4L1VAr0FJt
Vd04WTN/ZsoFd5Uv1e/H/N5UQziA9oCPO9g7zsgfRsKCcrV7xg04lt27tICpAnrN
ie2YsEFBHJssxnK57I8xpxqHL/gRrduAMw1e2sfrPu0wuK03kvvKOue27yWD2tdS
C/Wjc6ggAuQOxz9p+38tsuL+PHNYjpwrS8UjdAiJH6/24w4QPpbn7CZ8+AdA0cud
L2usNl3koh10rfdqm9CC3LBHoEINLIjFEXGMZUNZM1RndFbH5laVmzwD5uVuLXhq
dZgz9/bYxs4Bb+9iYq9QwfbY9C7m0Ryg2sxocINi5HPSrfTXqi4A3dBL5L1b2ZTv
tmmyTKEO5Xmg6hEZMvrK0TYtRUQ9l2Ps6BJzbWc1sQbUCMJvBe1MdsXBvu++pF/g
MXgwaKKarB/Y+H2l/3iqxD8Rnb1Q9/S4BlZUY51RAotEgmDTaFVDV8IS3d0m8GC1
z7JAMyzGvprOLCoZcA95WXj9uOu4xW3avN52JTFZ29NzwHvwnRBsZ53sB4zdxjHm
lWCfmCJDoay+smvO2v+U3LzptwjhaP/naZWGuNwORsc35wpCFGPitHUk4ILmy0hA
oZWsSO2PKaF2MRL6IbzN6/0clLvBMWh4nZaDaTlOpnFHkYIxOgHdVhD787ka7jli
zUOzUnuhz75Bu3X80xMDlPjRa+i4mr/8Dl36q43GoXIPaN41bncNLJEIMvuQCEMY
xHmd2WdkTjNG8f/x1uT4Cg7t+6dc/mVaAaIK/Eeu36bmAwAR100lF+Oc3Qr+5I5j
JpJXtvRfRORH0bCSEguSRxyPGGSYEk18VnMx5p26sxKKL0eY+Z+WKk4SbrIzyK7J
R1aGEghY5Fd2DLvtnTL6eqfCrDS+ytt7Hz/PjK1oPM4pnPJmzpWUlnoATvsgwHQb
vXM5o0Y3/6sNoQU/wIJKemG8BCgye0DP3GZ3lbkPJU3+qp4bVARAwtEjMiiItzYr
h+zhNbeyUqkXw3wyBTjh0rzanLunNJQU8BSC121v7+q29TE0bguOK6Rs7a9gg7gM
n9Qy38gjkXijvj/AftaqrjOH6Mb69khTzG9chMpClwTiFnsEgSfq3UM64hLMKjLO
tJZX9bgleiW3awl6YRadGVItKF2GR4brPc08riYKPu6LxVTXeqc7Ez+yRzBkQ9pl
B5fbkVbH5KsNdJ+rBNhhrP6cGNQuQnTO4ZAyT9URRKUcyhqKZ6yrwx+7XhcCDv+u
0ZdclYu72rosIZIrzebZfSKcQuNQ/f9uqZqrxDbTynxyTiUnbX0zKPL/b/JYAdCO
RCuh8bHfHXspePLidyqOgSOVnxz4ovQ4tDHkYIwAXMTHc6a0wgTXaKadldrjGHXv
LwDSCBlKHsGwQEXaO03L4b5M/X4WCjXg4YmMxeMp1zjvMgz0A8Cn3LIdKFFGYAeT
iRKmF0qVj1hpebtRZ2TwxFa7dT+nqVRD98Xgqoe8M+SCMI77tThXAaFqHASncb/+
BC5bybMKEykRzjVfb2daMorPqlSEBnU3g9XFomwV0LnekkEiF2eyl8NvBGp3ZqZc
mxKUEHu2FIvbbM3C33ifl9ivnnqyTIff8/nkOfsx5tBuwrachnPGl6yhGfsliMFJ
eqvfZZk1f2FuyqD4iOfTgVc3ny3tRPzDKuPksV0kdU1A3LY0wOsEuUoWlqh/JT1B
ROcP5vrxGjJSuKrXA2/CEtGgTfa+r8ZLBf+qjMKwNPu3tze9SxCIl8nkpuFzzmwJ
BBx5HQUHX9KtwTF2/+2/T7RwJmA58vwbGi+rGXalgD3my9vQBt++XBp9hOIvBJz+
+mjq9rNNw7wP6sZ8rpen/hAFRsLseh0cw4avVb6O2BRjn0q5jDfl7BlftgMvIZYO
Jb1w+kqlHE1Z2akq4tc9YsgXbaDgvF2OXG98jqCptw5qKVuAN1Ie4HWZz/L0Mprr
Y8Kl8k+OdS279wonYMFuGKbqZIOgnc7uUh82Dfv8oCRoP5hXfyHe1cmYeHBU+f5J
nxXek1Wgiq7+uRVOfsB+UT5+A4UvfFO+Cdiiit+tlwgjpLfV3PpK5uuP+1oh97AR
88HEK5nSXpfDeyaGIyalAvNqy7r9cIc2OLlTP1H+NjiDjrG4zjvYpBvVsuG4lYhA
8llmO3QBzIyCeqRWT9PJyg0s/0snFa1Ewu2fOcsbJYY9FHWEEHEPSL+Cf08zVDQ8
tXccoZj0Y4r7/RuiEwg3ZhQvkIlFnzYJRf/flAXJgqoQ36SDnkFJ946P5vQiCgP+
OXbjySrbc2ACuh5ZohpEzBgpix/3dXAggF5gbvLICvnKlGkELRrNC220wETuZXAl
oCRmG35HY664DWw5HqAP1oYp3IeTCZJckgPRb2sFyUHPYQPpzVenxvynEeDrMICw
Dc8nO55bT1nOmtlkoSVnZ1yw+3QYNYKkeGuj757H5WDRpjz/9VusfCQtX6qvHYfo
yqfHR+czYjDUcuzTOAT2R4doRtgK9oAxTkZZ9XeV35BzYIj0sGms3r/3BJD4+dgv
aDeRSQo0LNvpxccHOCih8+FT9butEiNfrg2LzlYf7CBgoKoQG3uvgIgcbMZcGSqS
ncyd0XpcHThW0Z1FGnwVhf+rfeMiESA/7CbgfPOym12War7w+KQAYpYA462+WNVG
ISDRAaFBJWwOWpCG6Jl23gLMTNBkV7V7qQa2l+WOsuz0zeKrlzLCIp+anLjLkfJW
cZaWi5N9m4QXYubvgbgSnyvXt+itpF5gxqcL5RwHrwq1LTwNkCPv/ENhMh3hqD3D
eC3y2DJ89vTFsDCfQ2yBNMET1tK+L/6LipGdH970Ck8BwzcX9VdHWQRwJsPvkn7l
SapnKcCkcEgyAq8W34XCoiO5KxIn9tYshdOmbQM8L4qW8QWosnTOx5EXwRAdL3/S
NxV5UYQjSFkZKyf6+w43qhsDoGXg1y4lIhlHGUdx2fR5T2mG41v94OTELrXOTM/e
OiOZheuEdG/miA0giR1lBPXiawOb1nAok1GPQhRrN5B2EbfpkS4gSHoEMkVNtrre
N080gMZ4pHONYqf5flTe5OBSJtcbaY1CP5VCOVZ8E56rJRfn+wGNYAkAtKjtItdO
2rbvV9/qF/SsZrWyumxPPu4FkX2oKCD/VUau1bAtZ2OXwn3tQQG5OYvEuXR+OzjO
pCb3H1NGZGS/WF8pfbMJOXRF2jtzpc9W8+848uo9eGMVDp2v/fKBqc+95YFdC2aa
Yl2RLtsXZTPkXC9IDPTn3iiWLgxu3ID7CmfUopscl8ksPhwio++AWl+gxSx/5oNM
hwa55QX83V5COluXzY+HLBJjt/EelWgWQdMPfiCzWbVJCQaRxbKxeu6/JkwTlDKR
Y1C0JIoFBSkqbpodSSo9X4cY99XIP3SCMEE/cEequ18Crw88h36QwO5ybxn6Xc/2
V5lEp2YcTiEYjCUjmJ9m8ilASbJ6h2yIhmHdZmJfY5GBDqG9/yy0pP7w8dPz36Xm
XwUz4FQNG+rdEAlzyMmbIFYS9qVxD02eLIg67zpcOXuz6ohZQmTWKOEnXpzDx/yl
flDHXht1Qy1E2hjJmtPk9nArM0+Wmh7t9h1TuRaozjlVzLAiNamiUNcrlbQSh43d
3+gjByvXXlr+H/fzPf12ZmvSnOT+3YddUFWL0m+cHLspQa8MOZ1GlTZb9plgPa8Z
5aWX+pmaeK89OxHydL9m7bLTZDryeqrJ0w8tApXjdXEE008BVmUxIb4y8CNYMz1K
lnD8JLppyZs21R0ZPxdfqjsGndIFjSOJPwHhdkiL3CZCoBbc7eR/zuPwjiShJRPD
5Ab5qtpas7VyceGId/MhhnQpzGi/qdyArE68EhPknADp20njxVwxM3bUeyb9MVcq
398d1l4KYgw05Y2y37978S60saFPa/+r9LkIfTW8kPltT7NEj1vKC+w5Bu0pUAEc
xifptJH0yf2OFtd0jkXuJmbFNwOuyLOlFbroYBoSY4FD+a8TSAaelbu9w6dpuH5Y
lgnrRp5rVkaF3fhioEA8kGbtEUONI+wgUPchS4qUlEy+tAUXxnh0x3HlnQzden/i
OLtJa/pJiQqcz/IAFV0hsn0aB9zp+N4HSUHjRq3u0iMfkoQVTCgzfKxAyTRTkhGR
XOK+RBvtf4UrkbGieo7slcDd9tc9PdOetV45/jBPz9W7qcQdqzi3Q91pfcUq2q47
JWqy1HzV8fkh4eJMvc1SWpE/Q7o3nn5S9VkWePsmUFDgcISkutuv3UFGhDwtFXwv
UjtDeOQKL8btDcd9dGnHwnnTswycz6wpmModQ5ik7jbzn6werHL1MMvANI8l+lQv
aU4uUZ4x03K5WuEjlk0CtSH3d9mhsYCVLdHQ6nQVtcdf3mXIIhubulRRhccml/YY
9LEEkChtqy38E4nRRexrGhKjKwvchFsSFPNUwcGRwt5I7I1RaZwkPDWy5bE4F7vz
dR8tO21rnbhE1CYIEqDBtQGgN+zwTmslsdxKb6PVxy0I0iU/TAOSd3uvbOwiCL3Z
0W4zbbfishylvZG5/jDXcu0m8cfMdYKQSD2UYo01dNl4ihIKfShtRUvU6m4CbXZF
HbaJh1HtjrB6UJij0/qsdssqJsR9QV3LPaMid+kf3GSyjzpE87Vu9KTcu8f+UcaF
McmpcA74VksLC0gBSyf4hivYNUsQSiLyP2QzHuMAX9UDQkg7WuLr4O8Rg8/aWDkU
l1anBw/zGG2hCL37Lun6QG1qLvOmMVSVj4RQRkS7oCiMD6W+rjcBS3vzWPFh5K9C
Xt35MOS7Da+uwn4jCpC2Or/zY4TuV330+J6ESwKXfgmrw+0OJP1g/TntVi7gGl6z
ck6wO8M4HAC72whbTqJRbs/UrXfr0K6lwTRqAgBRZ6hYCmWVi0Kk1BqGzGPtbZPW
b6IPBjEdHX9bTd/G/YCa/J/HXvwB9kHrglTNwN6ffsBP7KF246OPu0TFUKOdbizS
wGVJtboQZRJhycw2gXyrDyD3YQmt1Cb/jmkMZpdenm580NtgoTzEmCwwQGO4qruy
CadKUa4euOJv6qJeb2WbcNsSHS6U4QTO0D3z6tyOel8CAefiVXQ5BmLOhuRSsoWI
ZQo8cvVcX5u86gt8faZhqLNIz8j/f1r7Ei5/jncjBJdBbPU0R7djEnNiNdKtUgWz
ZFbnGtGFsn+fCkFZtTYGfo/vxeIrmjDtTTWp2xlJePaojD3ZlLLSkwE+7hotB9Y+
CaYsHj7BOI4olM5BudrSDV2KpjtxWxeVERXEKMPsyLBr8jD+Mw+SH7BG7pGWN9lm
jbwL3fEV7ZhvGrmOUcYaD+dJxHw1BAjm7volM8jC8GSBBSPi4sJOC0+hCLr6Srzh
TFwForoWRjLs2odmf0A692rLAoPIbr6b/80puTVCHLXE0Eu/kcWVbqvMYTsS4SHe
DZAXHM7a33kmIjYaRMzFuMkV1CHctIUAybuAMKjH8Vm3SBYccNlTtbeaOgmRSXN2
9T5tLWCvgLCawkuooMC1QGqB4/VtSDBoOmdvfHdShSgkBxD6eG090unbP9/7VkFq
1/sTFXdQ9/w1/DQvv8Fd2Ay2fRqqOusj/7NeijB60ILpPdICALj+eLMA5UJTh3QL
VQ4QoGNNysjZVkNt1zSSWJdo3odf4UoIjPBmA75pPFGumeppLroaKgGyl52CyaWW
hQrjgh30VFWMk3fDdXN42fjY1LTFucd1eto3CsApm4hQxNIIw3iGzun1MpHaAKjg
UBB/Yw4/m2ZMN/8xQjPST/az7D6/5wMIwyhgxZQZkFf3zBpuj28wfFicsrmGsaM3
+iK1BZ5i+Q0k+dMkLtT8oqKFBoRtlDbj6SdiPdPh7g8qaznUWAAleW9vPwvuwL0z
LF5RqE7JkOODF76KuH412lEZhdAaGY9Dzu/c29hVOLKflKBZ4+xYbYCj4phNfHj6
K1ogrV4A4vBmivoY6oZod1DmJQ5NBhTUoFue2/Rcs1RClZMosWIvsvRyWOBGt+WS
7GmluEwjqTBZ1KqHAZT2b+8XW4MXeZd0eB2UOY/PPAn+7t+3GbGPcBoY0GmKvZm8
/rHwJ6bdvuSoD6b34QI0nQyd5FP8sWqQBX6a8Tg7w8vQ4sOAeKOOcYuREULt8k8Z
A1wFO0a4p1umGrW6RcqS97BQAWoog3H22yKZURVuL83v97F4XSSmfAyQFwVPj48A
zVzLNJbsBm2rAoizd2PyHgSQJjSvPkblYfxsVYeII2vDQMIt4KRj0Kd9cnXBjRBq
KfdlMblQeMZ1OF/lMq2Xet2xrRqtfLGOrt2/HtDo5wQDtmzUuYdS81tHTfJbp8aW
rTSCvbYeqPleb/6SqDMFaWV/3ZlPOnvy0PLKjyyv/Lfxu5p02PD/kHICdyQjKbo/
dLBFrvyPChqG8ePoFjsEztdQQPS9PfLE9H4D0RlCW4EwkeyYoCuW8/AzKDIuzlgU
RU2ub01wr9s2FFmZ3fmfEARhuxcO583IQSZcOOIRooNgehSAwayMOfWx5FgY66r/
k+IM1WMvke0enfC4En74RKFg6lBFMwI20JKbbmVZX5O6CPW7aexJy7hdkGp2XBo+
ZK79NI0P+KZt8LA/hacXvhz+CAeH06wgdfUF8E4KBa7Ur7eXYzcFID9wlgnNuY54
/OqElVc0MVGgcPDdQnXVK1Hc7y25neFo+MEVXpFUckHOyJWlBwnVs1UEgjzzqO+x
q99O+7awIqAIxpYgWfWxJn2cJEdrqZHpHY7zxcZxT9T8XQD2lF7HsWqWvsBJ1N1N
lSs1L/rVzMhXlA3flDzzo4Pe0z9ziO8tMaeks0JkOp8q5MkZtmLQZZet3b/hZ/MT
xP+7yv1zlj3Ho6YJ0pqdofqqCm2kpIVCUIb/4NIo8sC93hU8ilK2Ii1k8Coe15Mo
nO++Hx7lbl+wOZgl96fjBrsetxtPXvrNsgbzdRQSxOcCxCkpa7AD2qTcsrNAtBqC
2c5Ba0YFTWhDvHfHfn2iEo+K5qdeXAMRVPjGbt3zF+PO/PJORvvdQNTIla03uFdD
vqcmqMxV71MB/ZC7/1YdwKUlqK7OgsXyVIv6yevWUaEmYO5Q7jj7eNEzH4rFeyiQ
nffF4OmwsIchb1s3mExuqY6fMQG9ySVtSX71JowMREdUm3qAJDonF/oGAUYaxG8G
OJiFX6dSUpwoxuyIBVt58S8yxggfy+Ok0pgaRuGdxTHg+XOWyLmTf+Yn3rTNKuu9
7Xl3z/6Q69h8t/12HGN7ShyswonwkM51AV8F9sLryM2NGMyiNA0cKlV6zxXOIU+z
GNvKO22L3e2D+quhWkD/96dF4hSTV8mRQtLY/hZ588U1Mbqu7hj37CQZa1NEv2u9
yycb9plihQKcFuVI1y4ARVxudpdFgO72/uXw6cYjw4ykazZo2Oo8H++6nK9grd/G
S2TqiVT5jVBzoklRsG3y/0PLqBcqwoIaa4kqHqsPK2xBhUMRSkNIM8eDjrnvTssL
7yaxvDK+I6hND1uKgNzQIli9NEwBfxYk4wzy5ZGvTKc+1jiEbG4OHtI27KeODcE+
/qH0W83aKGPiAeYb78/zOJ9cex5E8aZihsaPZxc0ML2G9RY/XnI2Z31L/1LfnwNu
Xt58BE9gdjD1RCfdOfGN96eeAJDiI2aoevn9ji0IHtTdefbR63Ko9tYHMCesctOZ
58jiFhKx6ITHeTrBXnpMXD6C1kA6hpbxoiO0Bwr5iM97KjB3AUKyOjsTo3LLR7cB
1/E5wbBpGq7seDBG6QRGCDMPqgXzCRuCb57BtUHhBbnclciHUap2KExW6jsz8L8F
F/zeJ2NItJ5aWtEEyxHhocqngTqvqIynOiKMVx7ydQv9G6nz+TAteA6XDxw+EzVi
5hf2KR00EXXiUuDRtj9FkTEaWolDq6npY7XrTJLY4kHTn/eBxb0cWucIFNmTG7nR
+n6mhju4xN5rWK7EA3RGGb1j5tlcPR5KRbZd6TUjB5CgmEy+DtTERU5ooPSvaiJG
yt7yL/p+VsUNmxAEiviRzSBolfQ7DsANfZTropCaLPkeIwWAAyHsmkShjpgXKNfT
Fh6HCg+eFYxOVeHAuRqV8XdIXyT3eovXeHGhxiNoW749GXs7g2wnnT09NwhoPkwe
kFl7/brU6sPUEIO3gsKn20Zfak+dKl1sYXEEB9/Chw0Wwumi2nX6z5OUn5zqyaW7
qobMXMk+687TQIFeEDz4uF2xkFeDRG9ilPvXwcW2RnE3qn8pz+A8kQUkfx0uuslr
U4tdBUOx/r/wD/kAzNZegBaL915TVCrx08OexfRh17+0NnHcUU47otQeKvBg3CG+
nRf3S5auxnxzf1FF/QVpfjUYyzHc9/Yv8hp6KN4I8Ai77LHkywkJb1XrJrdIwZKe
HvsTdrdmVHdUjz8HK3KUngWntzk7vujGnxfAiF5V6Gt7lQATISa02eDzWwsVhBUn
hP5486Bye9i9x/l5o0aVpP3yNWSikGBzydMFT5tGVLiqjrCK1V8/sqYG2AHVdgDd
nqYT2KzgKOc7mc40sVuFqftXr5jwNFsJk6UreQoB9ZSnBNzfbUyUJnXoOhAqGHPn
L1ZFouq6g+f6h/X+Fa7t2fGrdtH7K6m4Ort/Vqa54GRm1t2OWz0iQ6h5Wd2Zlxs7
wbj+eLCI/kw2/SOl0Vjcum8E0UOUAxlq4kZgaZgcAd6YtTETz683sZMuVl05TtW2
Vo6FM3/2WbbKN9o7UKyvS8twqvYtGue2q0X5GK0IvZfdpzpR14uxbs032pj85F1b
ORg3fWB5hxWF/5rucx57QsF+F86SWY+5ozGWWOEy9qoZP+L/wOwhksnTXY3bEtIb
eqsb5lKPDn6foC/L/ITY03ruMsdBbnyNNwd85iZQ6L0YpJRd0VXfLbHfeUEivev0
oiOqrptv6+6fklhnm8HwrHzlJbVpbsDA/kMHm8FHaMRSHxNfvNqC8o0XYOmbwbNF
ydMH4kq7EgtOuSedaj837DkRuvkK866TmSTv5h7PbcbpZSJvtjWFPOoapXEFIKLr
EPpl0S+FWrfqDFBZlHFBoP09rl86MzoAozA0rd829sIDdfTPtFtg6vgw8xMJD/1s
l96/EU0DKvdR6o3P/SKyUVvUoSixh8lgJ6rGMfNpDtCnqwkl69t7y27T42lCScW/
0wNapcz+pvLMjB9kFr+WQz/2nkFHtKJXYy2kpHY+s1pksk15rnPBf1ZI37nj/rAH
d8oK5kB1MizqwvGEUW5GGRuoOTc2BpGpaJ0vsNEU9einyttqKnM0i9szpTJl3WUa
zSQhNxeeE5nsGfdpAxK0fenecxS2Sd6q63YHWdgI4jYJKC3askhufxvkg3426fLl
LJyMcHKjNjkp2xQchKsm27/RlxVi7bgu/lGlJjVJ+Eta7hP9kOm3K3pducU+3MCb
7sUqB5e0hqBnYCckBbUOCfhO72/5VwATqmRm+KXqZtiMKTomW/NCwf5BpafKjTe8
5er8qWZakKFACH5MK+tAsdTQ80UgYSpxPEQ9yYj1iQsWke1GEJO2hTdoJL5XgrO5
zB7PDcT8aT6as3h5eyNhsg054fuiItrve2buRcFEZh64bC3YMkmQbU9CpuABMwFH
6kNnXGjUIO7wbnyDuMcek4so7pNldQRf54kbe4Z5djGmQnq5Q15DclskuzYkON32
IpTypg7XihwxfnIub9tMVHo7t2OfiEtCa+vBn7zX18x82mArfN2ki+1v0j45amKm
YlJ9x9AwJ6DxRUI0wM3LV72Q4czmCk7UXUoAbdWX7m8r58mDLsbEBLnKjyZnn9vf
/Aj4YorIKV69K/6/JXzqz0aAfdsHj/2xr91bQa/sxJZf5I3A/sHyxAem0ee2wU1e
pq0reGuaWFRxflxkg4i76756FSjVFMNM5IxeQ7EyJnAC603xff62piZUn9ZfoDDo
lnm5LpaqOB8PyBgNm+VmiG7mvQ/If/aC8kK6kwRlhNwj1v0Tqx3PNsjtdnc8VS4k
CYIQw5rBnrkWWnIPndQrcxRohx4eqFz0cL0NAJHjfsE2MKyC26XckaFoO/PCfayH
78L2o4Ivg5z5RnbB7dzoPJZKGV97kaiJE+oPzuNz55okBYuZ8wk4O4d6Sf7uUCAD
w8qSScrtjtLfXRXiTF7rjo/re/y1wCt3ARGl3YM8mLnI28DTN4gIZE2Cp4erbgk0
ydhG5H29l7XMLXThe1kyziBtlvszMCKzcvGP5h8d/WU4WRNbVq/CyMkLePEvGNTW
mv5E+bzU2FZVdwr9S+eqQ2fMbYMdXDMzhChwfMeIyV33ZemlPWF0sacLMWklZc2Y
N+7TqAwgx8h0HjI+I6t7OxflbefXlV+rmCsueKlpg/oLsnyq293WSDvjTjgHdTqn
/IIEMYhms8wglJ3Dwz6oTHQw2oiXgin7fU1NXHm3+cnm+qMiqiusG9WWL1cCsT9U
HLANUdmh55CoIklBGkLBS1ZMh2QwOsnikBRp7RF2wdQtvZcmZkE6xCpWNqPV02Rf
4Ia4W0RCN33/xK+AsnOajJfuGc3SUgNmoIx52/dwcyWoW0OyhgZdmVMl+5IhDbwz
DFmYGlyeRmJ8GNwiNOcZZxBftvuIPp4eEVvTXTQw5srQ7emF7vnRKOQ7qAvXmPco
usZwOKM1ClW8DXN7zSKLDo/DzOf3gxcPZim8RzT6tFGUeW+vW5l1hH4ddcbt7W3w
D2M6LQVy0u91Ai0+74KAKQt9Xi4eh6odaMnLLbk3G4CCw/P/sfqAJTLLhm0WLRFJ
7+qFwzcMLBLH77sMx94Eo2SeOdT9MjwoUUYmNmJ5pMPx1tpK9aAoJhmtHpbfqodg
YMcMlpPZp2lGHEDK9hfvGn9SuRDwgP5hdztwRCY2vfo7d6/LTI6ECtPpqvSDGZfx
GuIin8bGAOVVmTV6TzJwQyyht5LgQfFWmmvqKSstPGr9j1J2fInIIFAeMtk5iMoE
nmC1z9HVqa3ULEqGUe+TM5y4jwx0AQWqIn08UyJ6IyUWIj9gxtAGGSh+hwbdJoAC
Rrj7u8VAUMhUwIvdolEF7TlNwkQNt41ayo5HfvOIuqge9MJk2GLymw8WpZl2fq+N
xH89pcpfqauUHudVC+YhA8FY6vGfcRgijj1qxBfgkPBjrkv90mjkMVTPy7aIUdZL
8igFBZnaLCm+FSSTqMsf1NwAaW5GN/cNKhSN7GLl9cpO1JtG5KFAcLliqDtlZl4l
ZsST8qAxUUyFld+wRNsDOryMpBtyV11SbKuAOKEfN6SmfPsG9abjl4mLUEDblgTP
Yj5fpXn3Sv5f4R2xw5iOylXvPfb/d9/zQA8L+DmgjE8556N4NIX4P/cubUQS26DD
k5EhUu7jAOPdNTpuKPEipbHIZ6UUTjI4ev/78PclCWrNEnTQj9PmikA9fKBPU9Kz
JPTjrxF9O2YsPZdxK3ySNm5wl7o9ynaEC+/7rmgIaed+/UzLzX09jKStXhRoUnt2
d1j2lSaQ1LJa7HvJ8f91LB/6uveHl6UwaDX/y8X/ahO/NWulEOz0HFc8qTvGiTss
Gz/bnQD47bL7OSCT2jLGFflIQcLWoMDJ0uVaCDlp7GdQnCJqJEaE1K7UnCd48+aE
txHuf+ishePOLmn8FkWIKqOzV1hESMt9D6I5rBvwrSWfaCTxoWej63TXFTwzuwSo
kCuV2H9zXJHLTU1lFmHGTal/nUTd5enu20I/lqGgFx4RRhmlcMWpIYcZmjrHwd9o
FLQs0ucL8JtjAc9YGTuPK9g49q7uD4UgjdjCvVkbbMpetss7kkiFOJ4xq3SGxCQp
QlrI4Jvma8D/mH98Yn6SFzgQGrp32+EyEJMsf02PUP/pIkuMI6A+KgCTRQ3UN8MU
NvUbTQ5lCSKzjDyGQpxJ0CzCBrerd0AG/OTJKConE0MPoRgdpXkG7+W01tYtKkB6
kLL6Rh4WjJu4Q5qpgLXBdE8n3oGhqKJox9GS16ES79/mCXpTdgtdR6sVOD09Sq1B
rZrr+P8WPR+dMVXeKDIg1aBygFE31ivB+RcuJGf3n9T5LVxaqOA+9Wzs9V5ZteII
aATJc/+iuC011gXfyUMbjg4kObO4Xx8ZjyGhx+3zK+dka2+vMsdAfLT/uarLjxSN
/luEBuFGTybUvbBO1wBQA+d9FXJB91DVRlGDybHHMpTe28Pp2ZrjEZF0t5WD05bl
hQXu4U7KUjEkme8Tp91sSGgdQyyQvR9wctI80nAdit6KhV1I+kPcSHhfly/kbR60
fiMsTY2QMAWvs2PwxXHR5Esv/v8Fad2jjXTX2czSVO8IXNsiGrSslTKwQe197pkZ
jXYSb+4iCgNlJEFeQkxiBgl++R6hKvtQyFP7Z1eQPG3jObWhvjihznqOwadyad4R
095Vfzu6yuivm20oFtK37xY/SU9B1ocM+Xuryl+pXFDtfJLwZ0RV/jxuhnl3ijTi
/5nt7nb8HvQ7wmc6Aug0i8d1qFsTKd4bwmJ2sWtj7jfVqvsHAPOkn3nmLuEMz/zN
F4vhgf3zBh4GoTjWK2OHs9lRQdNOixIyMu6oNn8WJrk3aYsgOqRiVjAAO/g+CTBT
h/PZSCU5W9XSZTjhaGQqjamr2g/a13SnErFSjHwHaP5v55Y5zs8SeaJ5nMStypSe
wZJZcoSOQ5RG1CmZ57eWCxkMp852nyEjZUZhC7eOMfkYzkNiQCpuGtiO6dNijyGi
z27op8nHtQvRxrOnZ3pyWjpq04TcLTvhZ1EYf34v1Yx1yei8PeO24fU4nQMJBzQ5
HT2ltklsmStCWV0WyCeBQtQpM1Afw+su4RSbT1GAaESqiJ9WiYalimqbxROHQxqp
iBA46BjCi6jbnBOfRbzMaUewIt20g+GQ9W9aHjQutem/6iBM1Xpsg5FvKHg2n8PH
/YYISzHuKSpdNtKY2la/CRcubvFvTh2bDAI6Y7MlaOVQQy6RhdfBiFIz5Y2O7wtj
LHSRCI/bHuFhJ0JQUX3T8s/LjZ+jFOl5+0H6s2/kDeBeIF2uDx64f0N81875zB0y
xTCCNzniq+gOm4XBCoyG9GZMP3nAGvpYB/JxTro5rsYtR+XxuEAWzIFiTdAFU2gk
VSHa6+tZQwWGsCD0mY/AhklW6Zg+2BUzvIZ+ediejW3hABeP9lLoMAH1vmX+h14T
Kie6rDwtxWaNALMLzDlHSODCRQWsegw6cEnE6pW9ubAdkJ4TzRczSW6pF/0eq0JH
0runjzrX62awc7teu0gXiM3Ll83cCLDBeI6VWJBmi8wwH2AKaYf58tklJu/yr4h7
gsN1/PQ6A5F6VsMeXRRxc/SF8j8qN3r6ut+COKjmtDRnaQdhaebC480B+MWwerUh
sSrr6nYJ+/kx04PzVF2SeOeBIscwbq22fsReaWDqCESczZRqLhLq99VzPoGgtYz5
TrZSVgprVj1Jwx3cVksbzLYSukxvGCCwFF6Y+GUyHfhmwMjI49oo3mjVrmk4//ET
3GIiCu+IGRPNqOululhrkd8tfFszldD7489Ulj5PAPtssWV1yfMeIY25HY6stVOa
Lvm10gf4VVn6j3la2mg3rvYJneRkge5D/Ew7+QV+HPmHIvvOsxXVIzRWsPyCeyMg
eXuUwx13hjGf3r+0pDcXVMAGR0Jo2+yPPSrm5jTG54b6MotFtDgi8wBJL7UUjdjF
+O2DD1qGbO08G0spJGosl3ORVhmt+3spiDP5ozqt2f7ecbaT/wXl0/gD1IVcnUMN
ukkAVuTbwZd/ungnqJg1uCiAPydbKNtIti4R3ieuk0EvnceeJwmsI2YGlu21Dx27
hHdskxSO9LGVH8686pcYoKrnkjpBdOqkx2yWdSnBNkyPr/iGmuxIvAuejjHy5AeW
1yE+KQetUy6dJ8EdI5xezLFEi/1q69CRzie86X/H0HDIPhxPPtM6va1e6D6MrX+z
muJx6X+0HZU0nk4Tza9Nh3Ad1XSp/BchEgIsvL+ndUQNYudwhWnVVuzWp4ZY4QK6
e/Fmqtg5UgZ8nTGykFmzgKKicdcIYkgYt9Sjq6KRQPmAuix/aooAQEC4MntArPIe
5InrZfkVqF4s9LWQdkm5JZQU8vP9xohaEMECF69qcKmm8xXyqXptP+7b36mPm6wo
CR5P60LRFM/wDfEDjNq/gMYX84+uMaW1MYna+KhotDNNT20EYY+9H+orwv2p+wdw
CILBSQJ6XdbBre+OMQCyiZbrFoyv/oMH1/E/GCHND+ah0jOPaPU/WoogLptGcCKh
zfZtQ3cf9NzO185sdBhyPrF4XTt6795KfuY6xy7t8STwJrBVgj3gBiNne75Z80zh
CceW9nMIG5LHMioCtFezM8apOqdpjWi1CS7U4qsj+nCRjCJd5/+5F9/qj1ceVAkx
lN78VYG7GfLguKSpcfztvIzADf3VXHD7T5l3lj65XX/bX20/pc1tQgBQuLucv2BI
bAPIGPRvTXbwwJU4wl4xt05XsgqHTks0XkKijoqmAssy8tJczNBe5c0VtffoHZae
AcU3JFFm9oNNM4B+R5N0UHi9149AsQDrqi8DySrT1mVtRdBQNTXpUxryNsHZAwOs
mdvoaF37HNQn0fRYC5AmqRF70ZWHwQAxqi5gZGsuJfq2STNScDJbYVdHdAMK6UXp
YfN7mAAvxHQS+PbIcUUg3R24Bhhck8o//ES9VGg4enZqV5VUCg7HBzu0TkEsIjIx
WxfVT83wxfFIYKu7ej5QBeac4e+W6rS0b4grof1pLFfQS2zrbwxda3LQ3gYvY18g
WonfzGBm4kgLpCuT0OdakSJIzq8CEfE+KpohOn+mA6sPhDnHpJcQt7wURkvVmlhd
DAn24WyeZHW9hAlkpz04IevDRPoNPG8Atr6DItWru8/mLkHfsP+ldhq0jGOd2DX1
gGUw1VYQSO3eyItdMbmV+wywrRCGLALgecx7WgVKF5QEpmGOVPbwb9eiWO5sFBZT
IfrYjyk6O/cMjK+XjUC3wfXFM9g4ByMZsbi3Ht2saxnhzV8PSSe74PatEnnexlzo
jtB/VbpTpbkE8qqA/2usmCKkVxDX/knONrLylak/UNoGLB0PiPU0DkFlraa+p8UM
MZtW9e32z2I2SmxVw5nkVHZpOuLuDScdwfJZQWE27WTAVJSFKBwlLll/0Zcmdd5X
tUkJekGcrGDtLFsjREqejL3LzdSL05WfbpVPU6ydqUSDq1OBIbsukIEj7sU/zL4Y
LBKCfl2qn6zvrpSZjie3ZCBvfAydwlhLnCcHy3UBbRt1auflFNXu1GFMv8/FZe4l
eVFVdp9XI6j1A60oVG7EoB8WwUqkRzJ1HMSyPFxFtWt0RCAaYePN3cutzyi6y8lv
FtaIp5iHy2XWZ2rC5XA2GjG0jwW+nkRmwlpfdWu5wbFRVMMU60+JV3XHJIOYZ67R
l4mO8nL4ZineF8ZBRoMWuXAQXobBH0u2GUd2DRvZ9Oo792li/LdJJETnBnz9MjqV
IQsAWtYsbk2xrkZ/kGfKt33Qzi/Ivx8ZQrx09BICxSkZ1jcA0lvBXc+68+c/sXTA
ktfuHphfsQUnQHsISyQz+mHEytmae9w94uaW/i1MI19/fl0+ETy1nxcUuIygA+PR
SmPC/SYDCuQ1UJQ6EkPLPUCaiCdUq9Tf2uk2u3AHSrhW13qKeuuBDy9QPSgGSw57
fsQ5/ZhjFBj3RGtJWGRvi9MzxKaYnV1neS8DK5D5KevvFcbiTIwHTQ8OgyYi4V2S
Dlef2TPtg6v2mTwEwW/6aJJLEQhFGE3o0Bibs3qhvlIox1lKQd3WVfxcS8WKgC3Z
QEeG0ieYU55aRwRe8CNHggQvYH1e6SBvcurA4Lo6xhHehe/GJ/Y4meSfPFPGjqaW
+MSsJ+roQBOyTug0S7xbe9WMLYI7OQ/7AJzsvEsKtyXVdfU3z3pA710oz9pXfxoP
Pq4Y99n7TO27Q9/22D6AdUsWJPJ7P9PlgEW0vs29ArScJ9MhqEhK7xd3bRQJcKZe
7qs8e+/mdxy3PMFtYz8yo9asJKD+Pk6ZxCPEZjjN6M/EzxvYvCPC5bT+SDJIrWjx
O5nW9PGKTVrNIkUWNaPdog23RRhclReQnULHkjGPar5y+TOEIIapwis9u97PreB3
1G/4VTxXqawTz3nMDp7qK6O4iwcqcIQPJpRqSdCce1VHuh4961aIxWCMET82xjQC
TZN/CG3j4NvJw3iIgHJFb1IZ/mFr4p/k4hvlbHo1dtl37AL29sY57b6nv+AIkrM3
hzINzkGLoCMGLh8bjmSzf7y4osPdLcO2wE91VlMKElr4MBgTIuW/ZAmiSszCSndQ
R1Ac/2kv4QONIDwnO2T65RGvvjFjbicr3YzmvkgaMuZI1m9+dgm9yg5Ze8C56XnO
U6GMEzxAfaHXByiFNgC8Ybo9LyXvXe8r69/nPK1W4ws4O4ZROQYZ1D+n3D1nLw3/
fXK3lENmhiVG8ok5nhMxM54bGWsxWLb2GKablBBO1S97UjALqO40hZibcyk/j678
xV3RL+L11UoIvQT75i25V+9EQ8nTHmSSOGUcuF5+dMcnZRT9owGS2nQ1havNVNMe
8H7GZCjvxJQeQhgN0+amp9J0KCJOws3L0gbOCuYm6rnrcHJM57MDGzco63sx/OVz
Jw2AyY1tiIDdSzlRf477bWCNO4SPVlxwRs6F9RCo9v23dfx2Lsjak8v2qciHbRQc
p94idW0TMSEAByKou0Hdal8fmn/zQeJgSm8ZfEL2sIBxB0UPWOMldpWAdUl1okzF
6a/7h83FV0XY/MrgakFO6pbSRW8Ol7BAfXhQxvpvH2URjTtnFxMskOByVhJdFaRU
QQh0kOYCYaRT9HuV5lEICWtKl2aQaQCA5T3AIM+fFgTXEBCMvDc1iRQsTZUmcCCh
AvLZ3CRvLebEe4ONvoGj3rcE4NaKX7waqp15UMcEPbkHUfLPfBsKstrTxZzxSwcE
ZMJNfDDj61hrgppX6DE4BU7zy2yOQ9aEOGWPm9IZ/D12uZ9px+Jz0ene8z82Mr5/
mcZ+Q3Yb/AZYiogWv4XBd4Ee0LHA7j7zFXPyYS7MA+OvbG/tlL/AvzSSz8HN8iws
pzqCsrmQvc1Oc4axie/309flxSYyKrAE1X5u8S9K/PJPxZZdR4mdwIYGvRKTIfJV
RkwkYTUyY5UnjmxH2PgxS8lErooNpz19C182tCeSsOSNTQiIJCPGWRv7OR3qn2WZ
jb5d0I6sxuOoU30SNLFOZT8xPTqwTEA3j4Bd7imBcUY3mGWDkvkYLMS0vAF8JYoZ
Zr1vKnkHm8Wt0I+G4LnfBg2tGnYDMskpWKhcb2VMC+KzT6eOAofO99G9hLO4JHmb
5yNOV+eQr8wY4cWFRCJnJlCPe/vHPzwKbG2LJ+7+76oqxOwT1YRkFNv9oHQSqrgq
MFaB4/Xjj8WixEaqEq22AF8g3Cnwtc4OhDEC3Hxed7FP0BOgUZkBDsNeUdyizKJD
BNorAKylx9unbbKBHGFTZH4FnH6myfAjlPnG2GmgR6J38D3W4rGAqtwxsUCKrvbp
KyqYuDV8e/xwKsPN/zl0ZASmZ+o35u9GoiHHEIg+6AVftZdkAhUKUjQ9UZZUkdb5
JFTjY6Q3BzBqig+yLYvhQTj7ZnUBAvtwGE3zfes9HVZE6nDBMCqody+Ko71AaVa+
VAwm9ldmgYuZ+14Xn9UvdkGiGW8XuVnHleaChLpSTKWrCQckiXA6QnnTuo6/wwQ6
zLaOVas1+Eb1JUE/1QjM7knTFSn3jizBtC0AwJU70ETwQLAqeQ7fUoGsHUyQfhGx
tx6wIOpAv3tlERaKTDqRBw6hEbIjJoUq9FtpBVOBtFUPuGKGdePnaT9DUyBWR4+K
Sg38tuBYksIDABubSx9JDd/HdebyK0FQmpRMj4qSXwjEgNmV/zq7he5qOkboXfk6
vimLLi6u5xiiZ3uYZvEKK8sDtq7pD/lj2QkZq5TJ91vDwLUqhhBDet2rBOE8bezo
q5xyL5Fbg1kxaVw4ZeJ6FuchUNORMgA/dQ2z7mzifUk4iuOAo87Olp0P1PSdIQzm
NQ6tg+OPELlirQsn9gAhhH3GyJLalfw4fMkCsdKkNRpCdWhV/uet7KchMn7zOK9P
F4WxrOTwNqxrQOdg/174WqddQ1E3HsDJOD3K0/B45qsFmfDWnTRYzijXQ7LFpCy6
7IP8j4xhvX7iQBlFls/X9aFwjLzxgTuACkSCrbzVePvkCyHgTI3LMidmgdvqd3qd
w5v4r2N24eq9rt6Bc3ncwCn1+AQXPcu2N8ZYj6G4G6VdQBFvx1Ets+SZqUYLfGiq
7w5eeUcOZkanICIKrQ8VofhynIqxbqrS4xjGsRp+Cv4Nb89orwD3fmjWjrPSO3pf
KBn6uOITXHuYHwLRQI6GKwSk/ABDFcxaYuJ9itDo8ofmZbyGiYNU9H5r9Rol1/1e
OKGNfeMIrle7CML/jY6JyK396xVdtdqtGi98qvO57/rpGMcYhixQ8CG+UTeBxzU/
6cmg9L51EbuOPG6/8IMoPX+L0Z+jyP93WuAGqe6nLkcOYwrI3Gukjptvvxcyvi8y
+fpLjSgkgmoY8egXccwOKmQZ8ZSdn+95g/J19SnKdLVUzd+UOfWO5buNRHMZ5dRQ
wEui3xVC1WZp6j/IODQrC54ihE5O5uE2s6N77BXz2yT39Y8t+iHJ0OWC/pEr5V+l
smVjyT/KF5bQgfLZ+ZWufnJSUjws1v5MIPc/LKYYo12GNd2fYgo/Jzc96nwrnVOX
Epqfyd94CB2+pLehGDqNC/Q09NvI20urvUiwWaMd9wYjWelmCQJLvN2lsD43hoqj
okUfkQU6t8muVgERCSoa/wj/PnFswztbA0JcXqpdlTlMPhAvDUakQJU4NngieUt8
Kaci2jALMmBApL4lecQkUqHsxTOyXA47VdcsAIQFFCyK7Xnwwp0RmVI8Wgq2Y5VI
s1YjAqAh8nXwURIksi3kBVdVBjwpFqguO8rJeKuf6tiycUXn+bI0Ay1c5hOTjzuC
gjQZCgaHEm1Vrsdj0vS7Jr2M+tfqYcLMrrV2rQD04SyAWVoPykjP2Gre8l/1ppj3
b8fTbW3uhn7LHxZG7RkfpV3Nb+/ow05ybppoJ3oZy7LTSZyfLg1iv0SueJ+8kbWM
cy1M8CMQe1+xVA5HOI+Ua6envD0+sMmYOtnuv648/JRy0VgBaNkl/6v+6osTZ0cU
gkjQ/77s15tkqPAll70DcRuIQY7eKUcr9GEbzFzgbLCuBbR1jAMTE+vUPXef992C
4OKIv2WvEDAjmQpIa0mIISkV6fdOz1NW2a7+RKvG1gz2RGIXjedwKDZiEKuVvGVi
oZSQIaIUifd1tdMUAN0CHgie+U1i7uoQfndxFD1M7+DuF7LnOJ7HUVbZLncwXb9P
G+G33T5Or3yPrQfBGCIchFpd2t3aDU/h9eg0NfHbfV+LyMmdSpwoCuRQjofvEcIa
3hYicFdMeXG7AmlIaC8K6ChehzpFrKyxwT62RAIqVg4xWZzZ0DNZzJlBbRPx6Bxf
p/2SEf5KXEAewZAakvIyb1HYrawjLe0IrSfGFBWBNkaCBFwJ5HhsQGk4QoupW1Th
oVeucEuADGtowOArpADVsFClMo2+rNxjXy4dso5kcNZqbMVuhK784IISYGi3IRnF
ubDG4ztnDvZxDhjIYeBOLhbxBbVGWKHwyiPv+NdpJW6KK0ryppXskz5/ioILP0Ba
V2A+BWHeOiDNssIIST8IEOC15ZrcUonJS0cOJvOlVNYvjmewO86m802rrx1DXorD
u1OiqfiwYJR+BUvNwNc2dleomZdVQX++3HOZWjoLPTt+sjOr9rt6aqm0Blv1xUw3
prSbA1MRIXkF+wvamX2LW/klYj9xrLutbpzbKtAlXLMQh1+/TVmuYivSyVVXkDoc
Mvb9uR4TvYEBSzMCPpK4bxQOxAFII32CrxqDHBdomoY4p5e6oF7WowQq40v6QuAQ
a08/afUZcDZeW+ovIs8JsclKz8gd8mx6gtXAm4fP1cw8USKSN3xGlmXTInikSbea
0QPKsZ67YUQymZ0wQQxC2f/jLOy9DXugpC2zqXvHHqQQ8yU/9PNUsOIiEXR2tTV2
9VUjbJ23WTC+gUFBtdg43MgzaEnjW07u+RmkroTxM/cPFVsEX2PcK80nWkKIEHZ/
lm++65UDZGh4YmmpBaC1c+r+jrNsf0ZD3FOvHpi/2lYp2bJq1d+BJP0eMACebj9D
Y8abfWQYv8Ogb3J6NtAXvDM9G5wdtnOssmrnbWgoVtIETTmD/VQiyOgsFKUrNXE7
JqICoJk4x6TlXM6t3DtLWf7v0hX/v+6rw2oEkaSPhd/Ku6IKyhpYI/ccN4WMC0vY
ONzUFtK9JE/t+GwWE8RAWEz/Y8sIpsaH8Ou+ydNzjA7zm/NNrwONYpbq0WepbntR
KjGeSY8T6y1kmtAebAsCDtckfSSDxg0c09TmH9qq7b5HZ1v7R8qkiiMSGSVvgH69
4tLkBDLK73fJn6k+8wVcJkRb3XjY2BwFQ7LDWqpPLfsnatVfcVILa0V9OLhupf6H
qqUbZTHQN1fuhYQHQwLGBNzTjPPE+DLrOwH75gdR5xzDnL0rly1/w4AVO5AAihZl
29M4HB+xJob3bLR6k0/RrFJZWKpBHntSXvtY3BCICjH86XXSMFTNQ+MtT7n7Nvv6
khYHZ7idtRBbLFSenr2ac7S7+3YOiUfEtyM3Lj9Nld5/AbUwgzbZCGe/maVMVIlh
XCVIib1g5Drrc2cJDIbqsjXOu/QIA1rUXGJxGMJ73rTReJl9s8IN/yDBnjmXgH60
sX75of77UtBfMDwpOHAo0RmRzenHweFnimockfidSr0G8ymYkKEF/53QAfUWean2
8Vo1Uwx4mvw8nAwObKB4BxTaPOzAaOt3QsmdbyMpUwSmDWoUHo2eVV52MmDOV/RG
d16dRSktF7Sa/zR6utDeD2fKwAkHN+URDPZUDjyTzplxJ8WjtIO8FZ5nicSse/ee
ZN0d09ITLv9AtvEkOt/ztVWHl/atPEnX5rhar/SD/5PYrPtzku4h1zfhg/m4kS6q
lsanbOoxyQXNoDNgIgMZjiB0GrbQLtUovNxvS9fHZZoYxmjHt0wDqze36ctnjk55
8l+K9C6hyZNjwpvPSE31T0Wo1Z8TTlODNbLFJDBE9gjXqUE1420sdn/UzoDGY4GA
1u7LwhwVbExBkCSylLEak+qY2YX+zpIpDc709xydgM6Rmet0VgizpnahxyFj+6Um
sejblaEgrX7g+uLqYb/+EEX6Usl9YbJLJyqbmm+xFFZkCHQWzVQA6buD/qvK/yMe
4ukJ48DK7K1obaHkNm1zi3h40n0/Kk/TKbf5YOHgADVmwMQNEiTqvbq4bcU16ynD
kIzudIsYiikDd1mJOW9DewD6dI2UqMJV0TaHIqezApD2GDi4sWDjMY+lJowyeNrS
uPaBwHKbKV35xJncnGJcmYtj2bpvd5w3bBElxoUp3s6wddIDNdWdz4b31xUHTm6R
d9hFhl5580Ib20TcrGvD+pvyqeNicD5Wn6qSqjoyvgzRrE24YVhDxiY6yKaIEjSZ
T/x3za8/T0i0R8JM3+iSBDNgfS0buxWYN0NgO8IyISVLGO1rS5AqKZhFhVjWp2kI
XKrkVgKactKqBz/CaVux5tZK90rlQD2zBPJFBmFUrepbWkbx8uOi7XTq18b+HhQr
CL0LaRVknCSazEHG29YDvJN7E85Z3Li+gdVdj/MF3UK/7JHFoIPMFhmvt6D3yMzR
xgGclo6mMhLIr4I5RvAFG95if94TASEk1/lmgE0/DZ6JKM4jeZRlptkZgmi6c85b
vqZj2JjwJKElrOn/rGXr3A4lXzAbrBd4ww445TqhlqJsdBrA88Ldzuy5xFNafAd8
nH9tSR87I/JchNY16Moh1nyg7ihBXMTyOVWhDVKtmdBHQTLAOcQ3Cn97+ghjFq94
F2rjdrUVkKVVXnqEIEiDGNYv0Xl867LkfNvJkfpMEDh657iXacLgElXR0G3yLvJm
rTJCuwWq67PcHGpgJPUGV2I+1LfeyOvgMCthjBAB9Bjatj5rgoZ7V4nVex98nYRy
LuYMVQGQ1ZNa1cJyvPZ6ddDwzdZseNbwcccmsTjGN/vvRY9ezYWfpEeANugEzKuR
4qtlAs0OpS4mtajaSfqKDO6Qwi48NTqVi7ryG5a4OI3JjgAf6V2VHy97S5OYIrrQ
DrjSSkGygCKznXyMwtaC0w8OqYSUUGrYLXLS+Bjm0u/XRRQu0o9PxcoBt7JV9v0H
3FeTVYavJteNzzT7UK7npuGOywxNbkiVGCHUMEwdojCp32TGEmDcL5/PMatvl+Hb
3YMPPQD2yVhH1FGtYM2HMq6r3esWBXCx8ezP/SCnyFVQdGQQdJvhC6LAkbxyNag7
2Z8JzkuShsJsj9sgtTHr06Er8QQYr2zgLGwZVAoGPrbzy8n3NQv4Es1L3AxnAAy/
jGlRAXAu/pC5rK85VvIP9xoA1kazPoYbOuxaDGeU7gxxuSLWHE92DKdyXGv+cHys
hWlnqB5b1uthZRAuaP65X+zcVmFcfr2kK+aaECzp68UXxDqq1cpADPW80gBGf5nC
j1RZJ6Vni1A1aPf3Xcur1/VyxBzCmIGkovkfsDwRZ/tu9+klqKNVSj/NamXTz+8Q
SVtWgrFQ1NG4wyIulFU/8ikud2PxyNOEhYcHx9gxTmFCWCyUrfVQxJfmfiJjGr7T
N8JScJQ0upeS1e052AMZf7hr8o+jqCjq5x/5+/JAR+p2Q9xlXJqfh8dNz8AjUSZf
2i494W0yjK9jJWM6sQBkG4Zmfn7DYfksQliWX6RoGfEHpp++BEUijuJ51OC50HOE
YPbC1m1JIXUSUGOiWUlernJP74Tpym8WGXqxdSn4qLMF3U4QtfES/0YtnmmuLdv/
oc0zHSbPukCce1o7ma+08rC4OAyL4j2kvmSajwDgIzaQAeKduVBLZ8ubOPAg8EJG
ouuMY+XQUG7INvIOdAMI34+tc2HrVu8RFDQihYqEwqqrQbxqCvWoGG20s/vLsn0O
8IFwPZ22Uut73aZaW3C2ayIa2wNjOFqHabGvr46NzgdGotNFGwz7VENk3ey9z/SF
QzT6Db/51AzFCnBDGlymLNsi4NadstX0N9YWhT33vGh32Uh46EiSMQ2w9MtgJFct
Whcku0Mgv7XtrbhkOgs/jyk7dMVLZ8PavjpqPX/XGPQRB9voBqIgh+1oBYhV3K4s
ozOx+Q1IwQWPbbuqvfIee305VOWflgGBrEiqXtvvS/I+3k5aCO48iJrP8oONFJ/3
oifMuViqGiVTR4KcmIeLjmeDEya5aN/KmuZ+jWoGD1JlwbLHW158Dyqzlp1UIiS7
aSdFnRTDaZEmrlNYPN6BpgJM2UnAv1WPvfewW0NN9dwecB2IJ379+0l7jDpPc1hD
B58jwY1Ona3BGmZNm9cfGSFnGNv/H+eMEW46wXdf0Ne9PE9Wa3l0V9JfPfjowje5
y2jMmmMt+My74MbJ8eBHbukjgnM3kvrFFxjZuXB3b8q4XHV/NOpuRSBc5bE7HOt0
tqWJsrr+coJ3cffLuwgT6104pC6Wna9qLIDJGnUWXGRV3szwm5ld1LzTZpBjEBSs
Ly+n50uxRPLb46+wGHwztoSwe4AaOT+U0LjQ7xyOIGawzFz8uCPa8T9J/yKSU3MQ
5ApEXXgXNoGcKZAUSSSfGTrkPhK8s4eF8leIpnfku8TwxtOowFggMZb/5CTauvaV
mQATK0ccl4tUMa/vYZdWBrJDUZS5KuOgPasZMctbT11QegAscaLBGMOEuPrOujs8
ZXiBwwRSRClFqRCKCXYSGF7oxO9y3QF3k/aScYnE7L+dgGLlROwyKtCTI/xM23w5
2Lfy8gnO3JgBGeok5QFFaLxW1Hup0sWQKZc6q3WgSeMQpw05Efv+h3JXrLp65zlD
SeuTlBbQKCOg41bucKOQW4XJQHdWCbbz2oROZ40geINYsxorjT+uv0jRr8PeZXvf
Wne/3njx3/ZjEW1XR9Nv7yeWttl+FL7ln3gaDBfjUNmaE/Afmn+Egu8BIALi5EZc
Ns68E6smFUgDKrwSGzw1Dt+K6y25f84Y6K7NvS4A2ysICRDQbGcKKj6RY7JPpTEv
Lj/u0fA/TDl+OyhlESDjVE2Z+Gs7H9BybON4PXSmSXWOiQUs8BrtsGhq7d1RRMYN
6bU/QtVejU1q/OwjIEwh+zhR8zbGJwJsvBA6tH7Le45RfuHdhc6HUGHDxY7F8ILA
+TL91FgsE3dXhq4fcROIknBClAtPQbo8ABDAc9Tl+1KXxnfilCs8VPaT6fHgbFRh
+40moq/Du4Q9jH+PZ9X6Ad9V3yXqtYcHJ3UVYa0T13tCifok4Yi3DyDI7uHKL18K
PqOiAThyLj3dO083pDbWNBpNMEhSxGd8yXX+FMMtLos2pI/rc88ptaNQ2z40XB+H
qoBZt1OhfxxM6elMr88wLTNcfE/Psy6IINZSTK9+Dckqqi+OO1it8nSCOaVSxKuw
+E0xJFOeskod2caa9Hv9K6ULXl8xuHxNBl6DSvNtkfq/tdeL+Oiix8SV/47Vtydk
TXA2skPU+FsazqS99w3DZcqkfxj368oh/7GiJlQUWo9xjq/c8IwGYmftw4P4LrsC
d+gQfsiXmzEXXEJE0x00/X0dVCWoglIBGvtS1do0Qx1mVoyhV2Q7SrcsU+arS4Jw
2aYDJ4xHaczlMaX4N72NVDVwGBRt2HmRu/W4WGAqyDo0Okydi5niTse+RSB8k54z
op5IdyVfd/uRbze9epKkZDI8gTWkZNebkQVoeSuXgmnzVd0Aq1uJjFzYXiOikDGV
QyxamJfinrCL7qyjHlqOtmGiA6Qt2ie+J0xn5GRLD8entgUoIqK2Fm5acHE+QCqu
BwxF8eHMTSwEtPMjOSyHSaZAyyiz3yD+X88iFD3txKF7Phc/70399epP2YSlCpKw
R0VOJi2eN50Vz+QLa5nIlBY+t9t2bwo50a/ZAL16EnMh5uD1tDmA3bH4B+aDrJ2o
VQTEgQGucz7/K6qeMSbJIgRhEGCkajzLM3goLarkNb6EsYLwHZUXCzkjCU2Hzs00
mJdaBO+ANe/T4AZzYs1ADfYp7+2DGTEghmK5RDF6jyby8mPt6DvCDgpwXz7AYt9a
JE9QR65yTXO6GLRTQ0Kn6TuNF+6fZ3ixNxMMHIVdVHByZnbbFb6/H7Ep42cXejW1
VcAj8//lchgDnHVqUjzJ4leG/sj4YEuAyjgArFyYZslD6Udg8bGKHeR05nJzWutx
Y0GQizfImgH6TDleRBVtPVC9zHkGaFVvqCraC+Clos4Q3ZHsvPnJEO4bqNR/0n6W
m/cBLY5t6YHo0/EhyS+vjFm94ahKEhgCdwKmeMCasaYb7ChhtqULQxsX8Kto5P7V
7PmJFWRaow1xDIaYIgz7LceVY3XTC+4YVmrH2jsBYoHqSUdkt3RM48hepX5NyxC1
GOwfwtXhudbF+ZXyZm35bSM4zv2uKD5YgbIXreNRFRuNhw2SlGWMdpX4tNuBwso/
giviGj0B1cO/p1qIg8NsSoVSsrOfC44rnrCC4bqWFAKoe984WzTysp4wUXzvxST5
nyu5jQutWHc+PDiKFZAcvXZptzlhsv3vifiidtwWU+X5+J4E+CWhrgqX22a2FzG6
PILJ8IGmtQGWufhZk8AgbO4ZTcnXxqff+wQWK1oQM+sHNxsTuZZjy2xTeJFOIFk1
zY5m2AF8o7EGeF6EKxYxrUtDioQPjmSgAa6cM8RepWMaYZyw0vN5GlCGKZISVwXh
yaKUYOoTghETt9ssu7hY/TT4oa4AkajATFUJum4Vl1ehfi+Yf266V674K+Um4Prl
cCYNa+U+gsTKk/A2eHhdPZ4QQdcItn8+2AaUefouCdKxLfWM6+8WZ39CYb4cLYnN
FUFqOBvGKjoFPlYFzuZhw+AvJsOKbTjH7eH3ho2uEe4bQtAqRg+eAWRv3IFbKgCe
MHtYcR5RIsG9A8NWYNuYnOA/w36MrLP5u+Ilrz3yM4+jo1kN497SjQVZmHPERbX4
i/y8shWgZuYga2iQhjLCB8FKKymvEs2DDhWKdHYxumC3TBi/MqBLgICJ89ZageDf
v1QoNCmzn9kYhH250YrMN0wO0wQeQSfJefViHsXgfC482qXHUxXRxbhQtX8AL786
XYdtjpH/cy8Zq2KnM6d2x7/cUn4njTDtya93FXNCx0R6znxCUORERcW6scPM0kvG
1NkTAyUiiVzrAkyjKZbSgJFnLMq4IZXMiz82oaI37rZGt8M5DNx+0zc+2jD03rv3
/xzXn7lKaOelZsXYp19sRo2y7Eu3L86nW30El7cCQ2VuV4l8ZdB5SLcOoP2vmomg
QyPrEBvmcuYQkSexSIQkfaSM+HAB9ZxoF3VtW6OOGzHOFw4x7RwpKze0cj1LeufV
2gaCqJ2xxJtifv5/yrNdie/04KqEncHl4leBpBZkWU88zXpTtRF70LDkUgKxotE/
5GBzM0W/T0ByWNcAkrJindff7pN5Idd3sTGChyLRVs/ooD7rtvhJpwZvdp9w09v7
lpTFa6/J/bfN7C8PTTK6uLDmPUOij724sLONPfOoI6gG2kCq8o0aFO+ow5tQKsxn
42VerzgnQScm2qjT/GpeFVQhtHCu6LOCGSXPw2sW3G9LITbpwB2USIyYt9YZOIAC
7lvNjUXDb0oMwh8eFCgXzTV+gSbo9qeLwUhkTPIy2M74CfeTESw11J0pf7DjQRm4
MywSqPhOXbvVXlItxr3HdivKlt4mPzGV+Na04oIMfXNb1bt2ZMN1RwH2FrJrBJYa
0OzobZ8qjCiWQWO/obb8ZoS6SwUYkjD7xxoJ1+lgXU5iz2F1/FDcvwhNEPpoSCG0
rAt+gpNoVvLv4qe+KHebc4WuspVGbunCXzpsvXC6MttYeI9G/S4ZGTL+xOnsfsp0
IZqT9MBi3p3R9vTAkSbM5dZtcpTJXRMp79ZPXxBrl3eRcx203KwomQUE06YsbZ6r
vlZqFw+w2Wo1jsuEQtWOWiXUs92XbBURz9pyMu2CixvkJHBLVzNKgJe6ui02nx/Q
BbMV+2J5vVloms65bEIBnAfZVPzbnp9tJKxt6FnRhfu5FG6IpiSLjtC0LbyRwZl1
sfVxwsNUF/VghKJCAzXypOYdSdX66w9mP+ZcfV8jvd6p2BTrMEPN6v/pwVerjCzf
ywfN1R9VqwhrGmVhMOejSXEGtcBrfASpmsdgHErH2mwXZk5oeqjK2suAU9vymbSw
3dtPFrcSHrp0XkcUySNBE3krNCbyyoKV/r5oVZuubkH6rxhVb8m5UK2WgqqwVeGS
8h/Rcr4Nner+kSkjHdY/QT1aPOel1WYzBCqCpN+yYLNtdFm5WiOcce4+a/mog8Ef
vBYPjdAg+Ptq/HokNSzUCu5RJibHPl1QRuLvTqofr1Lkjp+72sKiwFtsNaE8FmAq
pHw1uyoJZ/aAnvppjM8uYxhMnzmoaoaIsBSpgsDpghx6KBk+EQGFxUH4TmukNd9x
E13hcfIbyCwNjplBS1Xn590NCcx/XILU4fGTVCSLwN1HSnH/b5rBBmb0zP4cCEaE
3rpzk+dMwd6L8qwopxhaDiBYv3dqPOFFCrDgB8ymPeCFX2ooCkAunFPTME0fCj3w
bCnlUgGJ4GaJX/x87JSDY5K8IO9wbRFW7DxJpM2PpIP6DPGjOxQlmENuFPe2hkhl
HYOauVK+wyzsDjwH6e5hVBOli9AHJjDjy3ebVyO/biIkfMf4PREgltwZJnApQ3dx
gxf8j833Lzt6F3+zQfsPvZG5P/+4IRM512KHjMME9dUaUc+mh8CqIlckhrcs4WKF
GqS0L7UonWiTtQnp29s4OAnPIv4HIoe4Xs0sZ5dWmmJlwJdzOEYZVwAmtEN5NHyy
smPFqG9siM6svNmiCHuRSIEv/wBLjliS7PPUwZTrfDLIh0bJEgXVLSkY4+DsWFur
K6fdOt6BuuN/Vq/c/4CvKYWJLh/CQg9qpIwC6MOavIJB5Ex+SC1QaSfnHtc/ppau
jmCr9QkvOkAMk4SsO657DN2wWoMqqfjPSLu+GLar91QP5JFxVZ9vHqJPZlfmlogQ
sH5ZGQAbJiGouLKHPGXMiTX57zHnJLBUt/g3mKwbbo4kR6Qu/GHXagkG9TTP53uF
QbVHoJH63Q4G1yz2Mjh0y90Ve25iniYXFAFw7528+GRFocD7V5VoAVVzlm+RtMQc
+Fq2zUeC3q3j1nL+qXO5iGWO6ds57wCWYflaU4UB+MIqerX+jayZSe9jk5Qvuctc
YApRREFtr7yiGHjllxmXqcfhxgxbArV7ol6uW4KVvjGF5g9TyRu6oc7f8dQBoXAy
urnbMwL1Os8rcyaLqzi09BL/2AvRQt+CFV06cIAkBXgwSc76ubCgmOhJHgbS8zL4
AI+kTuCvcR/gtO0/bjRMQoib75DJitF7OQSNxNmEiI0j+fBDp/Yiz6zms325LvA7
uZIraP1x0/qhie36z1CUtKLLEU5gcO1/kQ3hdsF0U1yAoPacD8lcMxqqsIHjaSUm
NC/bvsNg9WJC3ZAGsOf53WvLf4+yWvUHFUq8Ubd9ZruXrHfUJYKUPc6AnVlAIjH9
JV4dVWZHLbm4u+NTVZEH7c5s1pTdwu/jxn234RI83GW8vbxHzrEW9sgI3bpcHwvP
obrDQNqM4WnG8b4trXJF6MkJukLiyu+wOC2kPlQqXuaMtM8TzA+1MSBGlCStWid2
HFYf0kqrbT3dGkEF8Tij7MDuN92cG9lEOPMLIE1FFpCUtzjG7DSKW4hvFMlT5snD
yHKSu8mOJCaqOVBX+uWJJanvxDIbsBZc6pGInKOZL2mDsgwvkysabE7OKC9iY9uq
pCfIuR4V6fIoqtDx7mZy2ZZth55Eh8XaPzwzk+HJ5XfWOkIuNVTI+n+djHyQo5CZ
YSpKAZCZH6g2KAhyt2zSb42JEFgw1ODZHNXQNwlzT9KR82grDGMvMizrzMxHvYhN
7BJUi9/arLDHft9tImCt4/uyBMgUjha3Un2H1QGrbeDQf8r7UEOLd8FZsXqfxbBr
MZh/PsYSDp0hbEsnX47yLzL9wT+uv2B8mXQQrcyTdfEVVJzsW/TjnVO1OIxlGO4+
s8pTJ2AdtyIRlo8GDlZM0voiNlFfPTeGUnZ97Ylp9QQqVpwR6Gdb8I0LMcHb3u0z
CoFxOQcaKTpPIMJ98KhVGzJiKX5+zLyA2JeYevUcfRCsYgoa/V7x8V4CR7+cmYqb
IssDKvQ9K+gWDuYaDoqgSvDklpGqiE4NecDQyW+SdaVSEf1e5Kf7bf6w4Bm5Kw8H
6KIOkFvfvXVclGr5FgoI17e0J8zA8eOv9ur8oNfjHM4NCV6iuYqQtW+zsUcavbeB
ZReySMyHauySfP9Fd+E1wSb527ttt/SU8bHNNOr/cNnWCVCeTvP1DuGVUjtcBHmD
Or1Q2ee/OnU7scxpAYw2oTDOd9XlD+GrB/Qcg4ED6KIVjNonpkNhrP3WrqUb0Fww
MbNXwYLdwBBtXS7WGqLOQz8aJ363/YXxrwJl79kiexTC5UxIR3kZNt1n2YF6nHFa
6K6JRmEZYw/Zj2ZmqVdHMS7sLjvdIQwZTjfWaQaxQ8+OA7gJ7x9qUE/K7u9s0rzU
3lnKjw0yXITcWqOL4P+NLcKESsr+Rf0dxgZffzYHwcVwR/nyVjPeGrycRqItseEg
kERPrYOuj5NV3A1m7RfeFSJ/gGV+mgihvFJEZUJVZsYpvjsNpGPCaLUEilZUyuGR
8t0jTCOocDk1q8PrAtYVAEFtSnq88hNnQJ8hnWC1ttj+YzoCgoBkBY+AHyFsT37A
xBKVB7LnsbtzVUaVb1YkPsrUcfU5W36lU/JUsGRTKP9+zRJ18ldQFVwDaOkIHg7c
AapuNx6G4XuYvTjfmlZHrSvgZ/ZsrRwQYV/zgpBD4uyeIfAH3WOFe9JiNI/Lz7Zl
LcXK/UUQjCXSTKWDyQj6IaEbCM79yYDff6a9jhYjX8CGkrofx2m4VOkFcjMA5BHe
DuvvgtX/4IzlxUewq9NyW0uIu9aGz4HO0dc70UGblZOutQleJhd84jo3ywB8zeWp
P5R3PGtpHNCCIozlI4txWQcAmgpEbPTLJxXFyeIeeJhSfrxW1p6PXJ4zTjDERodN
vNUvdziBLwnnGGzCwVQ7qwnflmaHslB0czykiJ1xsm6YpSkXofMK6w5os4gsqkdO
tawGzh0Ftzqyanf9dIv7V+TkKGxeWKByOh4dQC9RRjYlMjRIvyjd8MPqwr/4YVbY
yKWDUwmJTG/b3S6FHpgo7oadEGxh04uubNfIaJU1PMeiEVdpRhV+HlUDLIcjMFGr
H0Pn+fWmG/wulgizX4N+sOI+JNTmoW2dpoTMxIcqZ9VbCQA/OMuRiEdrWunssmS2
Y7BmgAOpxtobrL3/zBiFTjkjg5GQb6GwS6pb3j4fb68TYPtDJRpLKcjZjBCKejdB
rF3NCM179GF8B2DzcMu3gOO9Bi1DTYzdSNpUdX8esW1y6odtss0oQdZGnT1TUbiE
8+zPoovrbA24cbE5Ux6XECr2NjbimxZrDdTIwmUtmkn44oDrjEDsooGMkCh3RD+d
JjXU39pRLyCSVUoXNlONwSRZCe4YjF8YeD2RoRb2FxLvU3F4Qr5vGktjhGPyYMNd
9JBtSwRE24IwSo12etEuIX4v0j4vvBQxVsO37+kL7lYQ1FThcUf9J86tFfSaAlGY
y53B2Z2/JMvKJkVPtPC2k/dE/tpvXTqN0GCjsZJ72Prp7LHXHBpj3jiymfSM5cax
Bj1Zihyp2r4bYRabyVeTZf5uN6AtcJWwvZV7oeDXCTrvu/htTupfydPT/vJhMkW5
bCg2uNSiWymwsRdIz7kvshx91KIOYUPS/cMr7zERy/b9OW3YT+fcyXkVEl+yoC7B
3RI4zwGm2nN/+JBrErUgFWI/7Us0H2F83GfR+2I9dpptZQx+Xt5oITHGiz2dokpM
NhjN/9c1INu43Oun/d1ucuzQlnmrWepMCe066LyCcfvEU29pLFGYJR3uTJzjjl/j
DZCn3Quw974Hn4ZgEozIcxftmD+fBYdwoxR4S/jTvu3RG9GHBLmgDNThAKhARNCl
Q8Na1DWFm3bE7a8snhQ+ygm0UbtDiclEBKozVyu1WWktxzQS2k/VQqKzFPSApkc5
VSN+oHu/MnYtW9dB5uy1Fus61DC/xSHSdim1UPhzLhn5FHuWrkbRmiLfMfP+H2yO
oBbHdc9WM/qyrsxRdhR1cVElZqwnNIhgPHxEE3psXL5HDiUIMES6RArp4xAzrUOH
A3IozoWDuBKKOqXX4yCAOkYjq3gmYWi7vMSuPtvNq0JH9EFfCpCQUdyByVgqPVuM
jaPVOILpUq57TUAa8b22RJergNIOp3t4sToCMk5a+SEL1I+PzPzgvuFel71n9Ss0
a7URx5fS5C1i4lcdTP0GoYIALl+8BTYOm/Iz4udddNv5HuEW+bZSZ+ySFfPFzEaO
bYNt9L3l/wYjKMkWkEpvaDAvO+cEMJI+FQXtcj31g7FS24QyUFgVOds0hKjLrYDq
+wZw1hd00Jy4kgKj9sPFga9LudvEZeqPUX+UUvaHL/qAsZunGvqJcApFNBuul/b9
tbI4T12ggR+Afy8uDFn0uFKJ1NSaIfjSEtHbtYxStWPEZb3bIdog09H2i5mKU6Ke
DT0fMbjCniLnpeyWoQd90s7wg5PjZ6nd9GUT7MQ94/fs8fWw0sNVtppkgvCzF27M
Sw0cY4ZvFTxiT9DggGKohvsD4y30HNxj9hOhnNIZj8mP8OWKDcGFuXcDvXIAUfGf
1/CUB3GF3BfGkq+3+vPuYE5P4bJ+4MBcekUQSokWIDjj4Pjdj1/d+SoEWEo1GEgp
nm7KWllYD3SCReLqJ7fF2omdwJj6kHoesSnyWZ7G5MQp7t/RVAyLz61mDU3+13Sg
vaiMAW607wniHg7o50ea2/yJTB8T3RqRUjVr8ulBYs3QMdVTRiX6e2+beP97qpMI
t42dditmYGCW5tKqMcXgJic1RUA2fok0+louOQu9SlUkoXlCaC7U6DFrF6nUYw1t
u44kZ25SSoRpLwCJ7x/AJhgC9Q52SnuGt0G48ZRXAuRH8P3+hY231G1H1Fxu6UY1
LrkoDXGXtuk0OvmJGfxEAYH/fpjAILJsYlHI/4COq7Hm8rJlCNkz7TfSi6+KNtoK
wkeG7DK92u7ND13nsmaStqlh8WCOoyZSq6a1QbXVVcaNdoLZMqdjULdWWCPWdaxQ
CGV1130iwHYwkT5nmezTZyx3uFYJXzgnX2KQhG2kcu1Y/Ux27UfnbukVm2fH4Ikw
5tAo5taMov4ZgKqxj75u7AYam6MFiccJc6pbVhBQZ6JHnGLVL876b9WES6KPuRJ9
G1Jx340Rj2NvSnZTsUpPwwcPu6QdgVRKNQZrbpMyFtBcTto8NxNAViwsa+eM/qfp
h83rXmhzafuVmibDJ9yTUUbefuWqm6Ly3cASZshvJx23E7+35bSNxsmaY540l8U4
+SEAhLVD9xI+lwsKuXlFiREKLYcPO9BKY/fB8fLFU6rU7D6uEh7WrTS89KqeeuMv
1c/GhCgV4MFitNVX08IFYBKJlM/NMByDgpB0yVlT7HpFybL83LdyLrbBPKse2AaQ
15iYr346HetdiihMy5uFUIQERwBnmcgQwqwejEasqlfCh1qxt8aLdvq0KvWjzP1i
kz10QaOZuBTd0hlwxC1cYc9qLvxktM2gOMpdD4lVpdUy6tFMBACowPn2xpu/12YN
iIYXZ6B5mTZC4LHiA4b3WiVt0V38f+uNTY33S8WgVuhuU6ew9Fbv8bgYe2f/tni9
IQXGKkTRoZ7sNv2jtmaK798NE0RJEIWVH0bpkHyw490y06hxhOEFyfT+RVJMeh2R
16DkixHGYh2EDO4XWzLPGBOiJrCwV5NWf8xQUDVfyB8xaAx60IJLYHwL6sja741G
/WP3CFwtJCMdyNryyHQWNM7rye3juZCOgNg5icf1/3l8v+mXDWLfJehcOzz4agiH
1jgNzSku11QuvBjIPm6ElhcyNEca6M0UUi0BvcwTUSPgcm5uastRgzug0g754Jf6
ehgxRdXfaj78Hqe7WG7q0yVRGy7a0gtRoP0PhAk/AKa9uaM6bPjlxcFaZNhKpKeZ
ozG8rGkbwazE7on9MGq2o7xsbvAypsRSIH+4k4albWZHCsdVl3wIhcBvmLmh+/9a
LUR/xZD+PuUINhH2V8TYdCD3lJE/7qZNAqrbFtOzJAi9l3Uf3CgnVleIgkd8jiQ5
/6vbSDjeGCEJRsSzhndNhiJ9hYZPUyPKTMc5m9Ouo88ePc0RFDQgplpJ2sxAD/SF
0BtF8CsZ7hfwMvhzSgrWRl8+ySI5yyT6bxyCi5ZdkL8WluXUH1lrnmMjxNE8rDR6
FbsV243cSaV081EjVsOe5c8VOG0Wdt92Mg1Snj2mh6o5DHdoWOhubDjd2EbnRcHj
6egtiH+aQA9u2NMmcaF20oyDFu9ywZ9fmLwjRd2Bnzd9s/sNDyg27uD+J8jUB+8J
90lbiZFaTKq5vkh2/FucR1CW/ZGa9bEFXjucABBIy15VHA5k2fAabdD2vR7Tr7no
oyBYZru2JnR+8ETV2JlbZxZWpuwDGjB8HA9GykwzBejwkY+mHcWyA0Xg9SXsrXUv
J54adnJCo4aDEYyf652sMACR6y23LKthruwt6SMcylWkcRVMenNjp1M34Qg3b6Pi
2bDKxWqFX2cdJ7SUizhdMmE1f7ZYOnIO21AL64FsA9DA57p6dFTYeUmgPV+d8N2l
nhrY4F9g/krLxQAvUB/I9xEdofliCLxvv8zrleXS7tzmMmxt7Caz3k612dFLfe7D
YUQipnZpHlDU2GMWVHnl0GN9Me9YgUIiO3lzpYK0ZdDnnLZTNVgAteHkeTj4VAmU
jZEjyOELyt7QlzDQMNf2UVh/09NngbuFAQSKyFWPm9refscwnG4EHlv+rsIN7qMO
uMCX0m/Xi2iyRyr32OiwxZCw/WAk+7jIcXWtEuPL7D3MPgbs22N8H4L3R6snfWMa
JDgF07ymZq3OBxvmZRBljqSAGDbMgPFTo+4a5y8FKRE6iENs4uD5sKZgQtAqvDR7
lXcOOQRCNGJMuQXKK5aTC7mZCfLvJC1N0Xb2s4dxNlDviYzTli+nca0Bf08VxUsd
hknKwJWUUL+nDm5brW/e1GGSybVvh9eJj20YqIVeI3688Jy4yRYWkW9a4GkdB8Gh
LjnMrICkikI0gbhqaVnZ0OuyKzbDW0PLQGlxlYp8q3elyuEmYr0o5H1XMV6JmUc8
z/T+ecKPexm1DMtSy7/6xtcFbXvD+vPQgTmtc3MWunUDQCFMq/5H3Lg5hse5fjCk
xanQw3BagPOmbTGjTET0k08S9uTgF8u+Ngdup17fj6P+3FMW17rzhXou2CMOsCo5
8ub6RIHWeqT/p33yojQTpWaaga4O8HMW+viWFpke7FqUHeKXPDRUakKnXYYq8Uix
iYZ8Da0v1lBQrzDbalZZXsaWaFLsJRjRW+Thq2W1u1zj09IvCY1DIomnxJVEBgtN
/W9SkmCiBrsqWJddVdqJNV4vlWVQOy/G60MeB3GAVhLupmaoxi6/EbPcPK+Gm9pQ
V1E5i6TKlSALgNKqoz+++2HjcALPapd13E/HdHcYtrAQXWJ7sFQd+rkqjIQftE/j
g2vzQ1IkKjqioFrDyjndOXMyxLZi+QlX8KKyzlRUDPPntrIyzw1aR6LZWri+1t6g
guXA3R+eu/u8WaDpZBgaKQGa7/NOVJKwT43UE7KzKV6gWhnKolukKo6rJZO3g81D
mQ6lYLmq1rorzhcBmV9DEEgP2iMn77ixO8XbM4VvnD866tVyP/QyXY/R2F/DR1an
6fGMNL7/d657lyVSW8rUDRJ3XDj/ccxuaLT6CbGfFfZIYjIkHItLO2KkMCM8ykA8
SMtIts/fbPY1oTFaPBFXpa2kQbEb39cI3enFJ8Zfry8aV0LbSG+21fRTas1fBENE
/c2BU/NIQZn1GGtez2Pkc05JNbNoRjrZibTAeqltX84ybj/7UbKi15wEFOdE7k8r
3cozbl/W6ixu/f8BQ1R2357Cf6CWA0ctNmzt3NDYEXB6roSwIKcyXJNiCx9dpPko
stMh5vQ2PIdHGFjiifzmOxgtgS7Ie1xhIjLulYWpfOPt6iSHRd4wiYtkiExhry9P
irN1hw31x8wyGeS0ktHyUsqYvfbqLVmg4y9t/BRcye/Radsk2ErKIvthBk9R9Kpf
Snh70/imotQVaZHks/o+dshbzDyxBIGiXvs8WnjAb+uU7wwJvM+QVy5ajOBArjlZ
Q49t3Z+1ujSHIs81yyrot+VVqq3RPL9uE5rO8GQ4AIVnylLg2zGdWQGDKMkB/9E1
Ow3LFYhLGUWh5/JQZ1u9ud8z0HW39Nhd7FClAgntKDcRxLR9/qHMf5n46Cl1J8nA
PBaGQiB2Myx1v7V0TAFS2Pn+u5EVJn9VF/YvW9L2cUvR5srfJW1WMTWVWrEI+9RS
WtETZGp2ysUMbuW1MQjMoXyH4z8RfZZc/1PAy2FoM1pwgjBMf/SDk5psy0lEN7tI
bkCeDBze2bQednS1Ud65m4HEpdIDxhQ9Dv2k20oRyk1+rkCy5hF3QesDC7wloBfv
iMpTqVS+2Dobow0R8JDz0R/XUZMMvt9Feyk5mmcu+zuGHBgK0jI9uYTZ5jt/IPYt
BEscRfoMPBKPZLYT2hPcpNYaZ1houlHFvGLVNKtElkJKWAK05CjObojet/xp39It
SON/WqqJdYve5JCq089wGH1WQY2sVseSA9tUBr6YZ3B1OftPmOXEwjA2Dr8F3tLU
fxMV0IUHMHlugK+2FfuQTWjnR/noRGJsz62+9Du5znNMOtJGvZB7YpEC4+NSLoX/
2wqVOA48/Da1syTTJZhb1gXd5AcklQcPNYE9hASdnmSaWA4SrRiaQV6hGjQcEEAH
dddPx7NkYBeAByb8X3rTCLrmuwAA7ZcaeNgh90EB+SnGlFxiza6vOPhSmqfrEY5G
yl/d9EmJ9LwZGIYBsj9atQUnwiFryNKpJ62khY6PeANGDgKmAd7JY4baFugJMOUP
mdzc8nDj4iU2kAPg85Zh5/univQ8SSArJXSlHTWL9PymzFcxZwjW0vAA8uS+eP4f
NY47kP08mqB6qSQj6CDc0mgNsFBH8ftJtcmoynl+MEfzzp8fQe5iI5UQu2ZS/cR+
ClRAfVJvD5YB8YjbgtwTo4fLZngHUUmREt90tS6kGZug2PTwiM/Zg1COp78i2XVO
ARvfbJzfV+eh8KsNp8KnHeEWavyaqpwfhrdyIn6a1JWwVbb4tOXBZx0jldN2a+4l
beJrmGVd48IEVrF2Fr8jpWOR/0dSC+Zj9MzLOX1GpejSrFxd50wjsOcvJowGBosA
LeB3GdD+c3xvPnrZ4LhwVBQg4OPy+05/7JVHBjmNRJ3dRiWsC1Qi4X7WjGmppENk
v3Pi25Q5Rga3e5e1LsmcC0ls/EW5WvEmJmyF2kBfeV2CJn+e+TjwVinUc1znaveX
DO6ndf9RgzZoySsZQFsksil59bJVREdb0lqBWSP7e4I40s0S2LE6U+0a5MTBZKCj
Fao90IrdN+CmKcahZw2/JPSimZyufczaYsLJ6fir93i1fccOFwsqJynHtgO+CuKR
7gQbg0y6XLLH5BJ+e+bsJ/3AXbzzgkUajQvfobFQjsIeYSzw2d9i+DPPLfGd+QRV
uN+OP2qzYaKxpRu7AfqgJj8GUqzo+ZdYhebpsm6FIPqGwnfXBKj3g70GMDa/HcgX
XLP+xlLzDL/chJa20QUmWSUfqDTS7+OX7UKwm0coceddu4p01w3ki0/rtrmX+bef
lxbCpahax/8Mr1XmU8QRQ3F2zJ2ndNtieiERLbb4kGXiWOMaenUipBh35ZM0VURf
yMbmOoZYNX+mZN/Jc0ivJ9gD2RcEI48RUcF6ZisHEsZd5xRy37UiPgr+zdXrzt+z
lQG8f18ajpGBORxXv0pv4mCDQtEWYolrce/QylihemN3IjYGDnlxA996GUoqF9//
274j2vm2VOBtFh8zIriZCBpuCQBuxc6nFhU42gNDLd+JYIzt0rzspt1pwvbSsYe0
Fi0drXbQohaexr8IKMP80xn1GrIPUeIemo/mpwPni1bTtkVPoJWCI7ZCr2ey4kce
5o/eLpgr5vCZqrQr0jYpzFQiBz/zsKfvPAECbUgwIc1gwt1B32Zbc0DeTZm9df6j
JKa/5QQcdyttijhQL+m9j3zNlLNmJUhF/PG1FUQxrZ49weGnLddWGlziFSZmYzXV
LKE+h3xOtmN7M8RZ20IyDURHTXimCCPVWklchd9znCG9sOU89W08GDXQxUR8JXZ8
zHoBTOFzjYMbKXK8mP07kmh/K6HL6PwGymjna31+TSgEhD4R3IiU46x9UtRulNrV
k/eLvqCD464oyKRK0UPGg0Xxqga8PMq5Yva1OZxEBr8ANK1d8dRnqTK8UXie2mvB
JwDzkEIE02cvmJ7MqyUiuxzo8fB2i7IE+iQiFmGlW9WhFyQXgVXd0Y+pmCs7Nup4
g0tt/p9vmF0XsiW3ZcRZIaRyJvvcsKeHd0pSql5KB1pdvDl6j4i3a5TnVTjkYtHv
wntBlXruIvz03lsfqidoraQ0CYmKSfhk9YeUNchhZ3duEjqZlvwOdAM8csmTF77e
El2fw/uwtAl9uJH6nKcj3rw5uUwOx8RlLNeheckQWiaBj6Gt6prFY+teceD23Pdj
Z6hYNdMLnwy44DlXM8JUsBa4YKpPcqlCDI+KFgF00kVk9C7sImuVG/xTN3bO2Eqi
bcSCxLrw535qs7paZliUyENt6JE5VCpDR1T2gjKcbavdoFDwJZVBajwqydmq2BiX
L5XdaRi4xn4sXg4VQH/U5k+cxX2ErcIAZ3ACmahoG1/CEEzz7jZvqUwwN0tsLx49
XEy9mT1w5ekoTue+RUxjU8pTsjMPvAYArUVOIyIxmQT+jRNS/RbMhIEzVLglu83n
iH2vbbE9mG0kGv9PV4C2Ar0gzmlWq+CobXxeqMF621Ig2+aXHnPW/tpxGmkJg9M2
DuiJq8qynLdVehAFUEz9gC89xmGM/jbF670xsgbEjTqEvGoDcMl5UrHxkrBvcPe/
+swrvf5JAx/3guQWj5tzXB8VzRCfcIpSTptKDD77Opid3aTBrPgO3lZFulEB05WQ
F1f+qvEBQKlk+HO5sBEZIx4WrjXSxtIDwmgrF3dwsTt6mqcBdzuC50flj/WhCjGq
5G+Gh/5w1wUMp929bJ4KDwnW7JPojyk0FQG81V1d5MvdqHVzMnNPEjSRu94y97/j
zJ9hRuzpuhBxLywFSqXdNXK3fbzgrOgaUQ6amqgietHn6Q/oCpUXQyEn5tBNAT5F
Q02jwBL2Nq9RQKwNyUqcDHb63s6W8wf735Tgl1byko6CUA36zvEMVC6bLTbjmKuu
ArF0dSfJyN1c9NLx+T87Xp/Iyvl61wsfw+WwDe4SzylxJaJFRjfi/VWHUykicVOW
Hrolb5MccMA6HHpkxEiMOy7pAYkcRV7+gRpMceHLZ1kkGdsJfA9AxCseNvzf2Uxr
588jPUcdIqdxGxMbHkJXdAxzEdRpSEbHLIU+JE0QD0iNym/R04cTvzczdlfZRwKb
GeBsbw1plm1j5hCLVm1YijawUobANZIWcRJZfUsc6/2t0SiZsYK+aOlt5e7n0o4a
pVR+RtN6B6JX+OP4p04X437oZOrrG4UTNVg/Y5s1bqxjjvrP7oLIL/+Bdsq16EwT
USIFQZnwZPX7VKRE5Ja+acAfeY9SSfqtlQbAVATjjrWl/s0BBH26JCdGsSMT/jcO
dIYizPPGBEdZ6Oed3e3vnmrt/AX4FVcSkyPgbHilcARdBvqy/pMvTPM17Pgv9vN6
FT2d6gjtWgdF1KJ3bZwk9qU7j3hz3k8M0vjzbdtGvgkNH8VQEY17wL5rA/OckRL/
MPLNZEFaTx3Th4HXKYTSgO274GLBnB3OrQtAe/OVqbnsPgUn60Px3KQUcJU1816l
ApZ2VNLZsWQ58hW6mBDnv4CsCyj2U3temGb6rJU/+8E6HcBw3tzkfz3a01ysaDi7
ZQTkmUOUb+nMfkZ+SEwErnpxuSyeLY8tW95ozERpzTvNZr+6JrLWZakHB8JG8v1q
sjV1jbJlBetBB5P0ZZ+Fwhj/qmYlwA+FTqWuDLoTjjd5eVRr/2vuupBNK0Qhfld5
uazU72wexayRPSJIjTmx88uTeWaujXv5uMEyXwACg5Qz+fOu/rzHq5YY5Eu2IyAD
t5ujQfe901nQkJ3XhZIDstkv31EB9jYlYWLjL75p4j7L4rGVr8gZLhcn3uwUDZvz
y1gTqTT/5O8SeRdERpXnyvsUxbu68v2bM6Xu28gbpTTRwVGBroJOyS5k6lu1KTW7
wHb944Nvr+sCiTmYzoQtTwya6PUZMMbhxnSzWH9BpZluoUNXV3m3Z8a28NW4jvbW
QZRvgaAJoI2cpkzEKW3CUbJry3arV7G+Fi3TY5wmP3xyT2t/jGhP1k0UA4RSBnNU
L+VpFV47lRoUhhOS3IHu8JNpk795YhFXUZQiMu4UDP6QOuJ0puiBVehV2gGjlgQT
wJIOS7/CDwK47AuUmHKv2AZOTjcDOGuQqDJMoJ/rUjixYNug/kpxDYfylRJ446nn
6opd+3+lemuc19MUy0TUBLATVtiy67ebkV2HU6duKwx98bX2LfzoyUSdnJef1MQb
W/mJxGDzu91NFibLATt3/uKux4hdwthBGvaaVU7yPyvOqfYjEoBWVdrbvJ37yxBn
TkZWhDeeYNCMCxAajQzAvf6s2HVfts8J+Z/JrN/1AKu4HXH0LS8UbbGYph8B/8FW
FoDP+HI2Feq10xggn54PHVwYyNd3htBjRKIdkkxrW8pgrtOQhDlYSkMYr+FZHHO5
2QV5Q/oaQyCifTPUbXFgHbV2wWjW0bFZNkqdXQ5BXIaeuX+wJgAyA5wPC+gCL3f/
Rp2bNvoK1THMbVRNBT9fszJR7suGOn4zPdqVpnsjDvOSO4KZzV5/jNscsCU1vlZI
qm6VHrCFQh34Xt30P9ExZkQjT/ghKOu/lVCXp50b3578G+mD1JSQ/aBIq9Ld1e8a
csTdS4ZgbS+cepMUcjWEK/Cryh93ZtYihv0wUFNSM14SNmP1EsBaVhwBLdd7Ltvu
Wq2D1TVbkUPTfLRxB/DjMUsSNwKn9YCT6EgWFiGayGyvg7XdMe3W3RC68DeyFB2N
5mCeGrRor6Oan8tGOy8dgVS2GDLLKmZ5gDxIhddub5J0xvx7ZxnwQ4paDQ5XsGVk
RGSoDLOcuWyCgJkhnTrpLZJjlrm4c9mhu7FN9h4LAi/MvRg57nxA5DONCFTFyRRL
BekJgeaLdYBpOtCQ+vMLDoug15F6jSrCk9qxOivd7VepR0WeErvqz2q92F9dDRNE
iKRRzLDFNwESQlWJGhFEYF3Z6jxpNZ9gfFLCSdUV3uZhR4rX49JYisX8RJ9zni5/
EULAhrxDRaHBj/U8lPRUGjQKNZe4/AiTa9E1xYagFkXE5R3k9OodpaisxSFn/Ewh
YJYxmniT2d5Ztxz2m2guRWrZF0TbkaQhOZZSrpFja8k6/rOH4g/+IjSqBd/ebPKg
mRsHQKJk/hgmLQ8wzEp+cW+as68BWcD7NzXoxDJImd6W+wKYsuMMbVDNOFiFV6o6
OG9AvDzJSGPJhK+GuMBrVaZK1bamr+nuVoYWvA6q4CIbsCnVHUNq6/qSzPVilcY8
rRqDYGzGPVWOd98W2SGGHglnPALEogRUJe9HfHyr5bPnIB+cDw2Bi1qFz0HLj9xu
pnlKm3BPd6/VcMu/4niZtJuP9h/VSdUO1D1g1ExNUoCAHWMpSMgfbfishEASmdkc
1TxuyHbmdaPyJq6vLZvXzH4fm7WtDcqflQ0eNSXaIXAWIhRCPrZMMjpVQk428h58
MWdnAFhIFjDApAb4axryxy4v+ZpBDJvZeXKxQy4jEOO76Qhg1D4kS1abFRDgwPkR
k/L7mG7l4KFFyQzVtgMinATj5iTJam2sPgiAR8A0hTnT6PA4OdAeJK6z8hAM3yOf
JUG7SN27nsezDeXH5EU3Ro3UzdTW9ip3/OrGpOS4xXbyX32m6jzEX7utKQFKYw0C
AFftEJD2vB8ADUPhIXAb/CFm5XUEM8SPyLODtIa3zybsu3wb0dQY9oVw4qHDrxjs
YttxgtO+uFGp0mvLemEVhbBOhYf4A9oSEOjgWFAz6tIN/R0pbPUzP2zcvgDO5yMM
MLpd6H+eVWjx546vQkqZLY4mVFjm2mODe/4ZES2oQuiY/H31/ijk4b3REN2jIrG0
QSPXypmbct8JVNEqkD0zakc2MlihBcDqfD4HvPv8Ar2tyq66kM1Ou26mqJdV/Wrl
z/jkk9DAg2YXQmq1s+FjLG0Jt5OSXa+jfn+/rzQ3rXUiRnF+QygKjVxqtry8lCYZ
Rfz/aqLtlpeh06Vus91UIglWjoxg6/VR8SCIk8ANoybW1MYBxPpYGGxwuQeWPNtJ
W1dB/x6eINqVG2Xt1EdgWBKlmGN3jsJA1OhtsCpX15OFREA3a+sAuPn3L8wsc+04
45CXgoQnTTGurFiw2N60nAxv++4A0CXK5uIN1qnqpSf2iF6IC3nH8NBrj5HUPeQH
OnrBZ91+upcuL5xG5aT2e/RIZIruZ+7hJf9fR4VmXndFW2yqrxNszdnrIFzBvyB0
8z1vbWgs4pT/uerpbiKsI//QQcMygxEz41mhuksboCqTX6OznzvqoNOCOuED3CR8
jPm45Gx0c3fFjp3v4xfRuszTqF9MQLEqkNpBCvc/9VSlAPtTKp+Y6dtE/TBOX4ho
vZjNA6jbgFcs4IfZFoR99RObHoveWUnEQ3o6MUT+S6+MavI/Whz9WvCWAYIGdsOB
dU76f4CtdE3uJD8HcAtHXeLFztchsJG5IjcAu919Dw6UPHvqXF+J7/nLpky77rMU
s+RjRW0NV2gc81a8s45uC4M4BJwvSJKlhsFKiW+XRiDoojSPUGY3gDn9OYAohJKM
EOB724iKoTqKRITTT7AabeySeeb4UjusQ37tFCaOgO9YiJeBVLUngsyWsClFmbjF
Fe/qT3hgw2nLn4y3D0Ym7KNEKI4qsoRs3Oa7SWuzq3IEwRpCLYi0hwgUDs9ePewk
mLGMXC9wLJOyJSbI0RawfM5Fqt9l52HicpuSnOYfYQz+HpeIGlRK3kMdMGWN7PhO
bkial97DxexMNRfXfyGJu6YhrfiVdIJFNdGzuBtYxR/jfUU03dUn2wIkcRAXLKEQ
YXgXS9Tb23scyOlyq/FViJAT19GJhOIBNxiWIoa9YsjXDmcVISkDMa1ifObAgC3Y
Ini7hoeOz0Atg1/9VNjzzyRcu0vsMD3fkk64xLoOaMb9JWYcP5L7DGgjdXB9cK5U
zzTfhJxdXacHJjW5qv8ULYWb1d7JIB2FInWSR7isCDyOapJ78xojms6FP1CBGnPK
wLy2Oi06o5sl944YFCIPnIjp/G94iYFzmjAgq1k0ynV/ka6wKMfjb4k1nYvRohbe
PWqRWliatd93kkgIGF8IoDGp1hiaLs1bAKX69tlq76FC1ijOONCNG8nNWbORQdiq
p9qANc6PnjVXTlwigPZoFxiDnnHLuhWC0FK3EZoqMCSj3y0pKgEDtRBNcZBKJP4h
DRfEc3pZOLEQ37UggBXh92/Gv8zvrkTMMMm1xFKFFklsOjceNNdH0A30dps2Ju7G
wFSrrj2C7P/3qS2yjTYyYxCFuwok6SWbcuIJCmZMhed4ADXjZQX+FFwFugXayftQ
WxhgY5ESFPVlcRKUIuveo/eDNRLEOYJ2AAXkY8Rxh8WEw4RiEJt/CRkuDxTHM4jc
BIH5Z3tA2x8j8fyXKEkbmQc8X/AT3kPQz7YgCbTTqsj3CGkP9g/ojUlk9GA7v8Jr
zXrhDwtAk2LhHAEtsKQ1y68SjCYInZnKXk3uSdquVav72XgoVh3H/SD9AcxIJdS3
0izGadTsDocF9m0hEYyiE21aa0udG4j40f3XgP/tdT76QYIGb6sW7q490fRE/pAD
QxZZRhQd8QHkNVJag9soeNSpDOTMoYsKsAG0K8ttsQpmI9DpCRGwDSXShnP15qIj
8tRVbEEJjLQO+1b2usRm/UrBScVJ93pDvC5Ul1ox9VIsuODrN45HQ/cOrLDl89zb
YxkJvweoV3qL1O/v0JJL58gXpO7lP8EJT6I+BmozCH+lFL31SFKwnJlDxG+URUZa
NsYukrBpnG2gUqTRbvJyDa+EOhlO0eeOOkLqS9fa+zV/8bo3A3ui/GAGFMzv/v3a
9gsr/h36Wu93wICDVtQfqAB/yJAObHsNdicmQ80s1VTvlhRUHa1DLQSRGmnzf+XN
zqkN+h8rPMPT5jvovBJpFMfSJZajbjKzOjNMbm658li6mwYq4U8OkHLgD2CFrzyk
riJMCA7+RJLK081DO1h64mEEknfRYuO5MeSwecw7jvEAUX/oTEUjRJN3KXzafr6m
RK7RYBEkv9sRd/I2cIm4MbrfoSldeJGfaOgqbnh9seREXF/aJUT5uQs81ZJdhJeG
0KS35bUtGvFdWaNPpTomSdyMJvvYnZC2yHDeIgO/xMgbcN9vomyA4/XqWSw0qmFC
ssigD9R6mydEXzYu2lOWmj4xBCogF+BusDPO/YL3K6KPAcYKN8MTPFuMeNLWg1g4
lVZZywUxtvKRy5Kf2kT/3wKKOlpVXIZ/pe0i3XFXBhWs8GicY1LSJQn7+FNjH/fu
5AOZELkiBPvq27BKNftNoYwKM3XkMUUQv1EmLng3Wk7T5iUG76bq7xuAppVu/vnR
Q7ZrcqW7EnISYW1O7Bso8525Mt1GgW9BntTuLBa1wWTs88lqxhkjUjYJ0ISkdLu7
TE5QP06QdsZwkf0xWXjcnEX2XiKLalCiFb+mwVO5x57KognhIDgDDwj3/epXyMT6
3Nu2f6RgYjyVWqPbPqgaqrB2GH/4YDCdp/umr7mXh/pyBZYvdtypGwN91ramMZrd
3fsXtv2SsF+A6OCQbW4PgI1nkx/DPRTxrG64nabws9bkpolFOhyVU7Ml1Qt80VZC
WBrN8BY7USlZzcD4oyQmreeotMAbG1v+GqNy7PKi4m0ubVk90cAWRhBNoJeg+hxV
jlZ6UOTcC9d63vWAIOWEHuA9nD5HMlkCvCAyeY+AOKCYQQzuXFrERVNmb7S3vQr4
gn60u+Qo0zXSrZy1xPRz3QStd+TifZBvwMVA0gvFPwGNVxWxFBwF/lP0TRxY9G4f
kkMWm43Q1RWfZHRh67R/urZwhfEgxnEbRRzSWn39/3ARiHytAaFowoo8STy/pLx7
jRoxIP1VZjoUjvw7o7oexQ2MGJLC1yMmdLBBiFpBuedlxM67Ioc+L78Rzyfao0It
ly5fCTJAWSmEUVIpCSL7kIi3lxLJ583ffvl8ZXVdNx6z/PotjHd0ktMWtFoNxqqj
AyrjkLfXTrbAXxqg1wuv8fZzQeVM1qRf8Gw230QFs3Ik9TmZUJ91zMaGrhHeUHk1
m8GctM4rJg+tPGLjJgdcDvumNZA4q0l36y3G3ufBYiWIIRraUo9zyIvu7fViKqX4
VJp+RsBQJekTsoUx+zzpsWsT8/mHb80QDLPnhHggILNCRAu/9YokQZlR9pGq75Aq
aHxkn+zkYFy3nuNT8d8ZR3GZioNTtYsIMRNNaWFEtlc+XSxeQRK9k8h1cG+lfrqQ
9O1YHNXd14XK046DyXlI8w6w4Q/q5/I7G7Aq+znQgQQO7s4WY2Yie3gokWEm8mB0
IVVJ7wGa9LY7wvPHZiWNgWLGE5wNN7tuV3+RH7vIjQrVkHHgF3UjsVphpRaEm9Sf
Yu+jKsz6Tdzo80h5kB1SaB3b7UtTwG1nphiPG8Dq7w1lkIQMlDlNHhNu0HxWUSqH
p3iHXrrW/B7+/xziIsNi/d4SNyXu7D5v55/byRkXdURYRa0sgYBWDCUrmGpIEFk0
c/msJXM08d8MzFwNDW/inPbbKFxrtH/1faSLhgIYuJThC9dlPq+ee8EWda4L0prU
+TC1ygLUj218W7fgLMCIMFJo1zdAgdFYwvXR9Vu1YUCUcLERn44D+sRywssI93PW
t7TJ5Nd2tNP8XzfEZkYyrbA+Zhp428lzT8+STEzy5mEbqHlkLOgus+lu59AzkVgi
AuIUZP6P9Hq6vct1Ik4BGDlb+kF4s78vb1hkvx49fRN+NrFdOHmdSqTg0QT0F4Ad
r94xrwS2rc4jfHRwEBgWBtXzouRnVmY1FCeHePN0j8qsoFgvRseKeABeRvpdVSll
iGy+Ofxw34Ncs1C6309ThR9MIWtVfdU4adL94ldupBkZKHX2jeiAclTcBCFzPzHN
Jnp1Mz/tjIpgnVpL7WoOO72Xhpd9LjyVzSsShR68CrYg00AzmTmr3Z4pBd2OHvuR
2fvWlCUj+rOmORdZzsb7GhR4gQJjY5i00JZc1U8dLPGefvQvxxGxbXSDkhjFOjWW
spHDqz0BeN4KuUGYhOqFATPSKKwgMvGhp/q6mJP+WnGDN4sSa0Xk83PpQRfdLyDf
3EM41xcvfGnALU7wHx3HcZ/bUWyH5NnOQy3mY6uN97basVt/KN2++ZRHaxyH8FGd
ozOCECBC7eCP4qtFOWKvTX+h2n7p6QA4xcTSCEW4ftvp/MtS6wm4HC9cKx8MZ4Os
APo9KjmHM+YBHmxbWFOtoGPZBpAEc0UPZgM3GZkCkSPVg9q8I3ObeC+A1jmHk7H3
88FbmyVD6mSSlmoGWvV+wcZrsdEaZwXOvnaQ7iT7aqPDYTR5d6xkWV0tlbfH/E2b
SwUf5HnprYEStLNCi/PLCM4hx1DXcApH4JBzK5iiO9SdcXjeMENCWvwx2d76Wuua
vRAcpH5OWFAYh7j8xlrBGADVWl0mryFS1Cw9Zym8DQqvodria8qR4sXd+Mv5BaXG
1RFTBBW7Jt4Mjf9oKdpUrcHmT6Vt/sfFVNb14QFeT/8+eR+Bez9l1a9b8uyS2Zj/
J5N87svLDA6aVYlRdW/OENViC4HT65IOl5ZLuYsTuI8HUMyV1485xjudTNNoL7Em
3jh9WOGgPPN9ryG71eAhRzSkMDJHqeSjNH6fkH20ERqNXnYt3dXAdisSfTJpf6fC
QcbQa7g+2XnGw2Sn8ZoB286bPnrwRm7fcdqclF8IhBsjMxGIFlQzgAx/LC0NMFIQ
k/YI5QhR9ahhNWecAdRIm8HMYMd+ZqKrQRtmd/2YffDMFe1dSGL3fnYbdOoJPDiD
/d0Z6cnFjcGd5ZtGkE3T044+Bxj0gkCgnkPWvB7HldhfnTjr5pjTeiAL6+TTFkbI
QhCA98mdc3BgYsGzeDL6Gsrcn1ItZ0gw8TZ/FEk5uhvzz5A3yv9ngxK+9gwCvvo9
QulaexEU5h9h1ikMLIhhIfDp0jWF0xHwtc0aFekFK4dT/F4Ag6dt6kR/m/A3PYBG
f5duuENxtHWo5rxOVgxvaXNcs/ESw3mUVZQ3qKwqdKToldSTrGQumjxR26W0mS+d
+FQx9cToBC8hFU6VmWPNgK1q/EqeYdrDJ9td4lULo9TFQg4V6B34dY7YkL0SopHi
KWEsqYZ7a4AdAnmWyrhw0pxcWfQn+IolRlJ1TNGZllidKmY9hCxxCJ/L+Bf5FKt7
7O3XJhbhdqvbFX0c33X3dE2HSgpfeWcE4/Mn6C092Rx/y4tJUkqZyg8+s09S4MGX
memPQV0ppNpIo5R6u2+H+YGzqXb/KViC40EZoiq23duZGxpFnt2gnpCHVbgRSes9
dM8ECBQOshGMfePYhQAWLoaKgOERQqPYk2MBokR/F7t43VPkJLEiVgRJXKVVuykD
F0V2/169ombu+h9IimoJ7pvLrLwMYNKCmB5P6xIiALQxfap6dNh1HlDztk0x5R9C
Pb7lTLT2qmOmmJaF6JSX3yg5ktNOOkutV6ptkoINSNLuxkG58wM43+Toss7/aNnG
Ljm835FdCA8fsRk3nwXVPqoY8GdJTfXucqyhA+a6u/NLzPp7QmmXRX6rFD+M4Aio
6bIwpUigRIvwr7jmmqwqZnnzl4Qv186xGyXjI3INY2rQ7j/67ogGyRWVcPEzNuw/
vQOuvIukCrCgIZLKPSXSTBZ/aUMdz4PiB6UKx7TFAlNS20EUqR5D3co0un/sxu/E
buhAz0T6Yy5VUVSuG4ayplGHc4q2xyIS1o1BjhTGPN0xZjNxBccuPBEGvKiNk12X
gK/f/8XYPVGRSBQG8Sfc7FL6DWfvxe4kQPUtIZN1aHLIajmCbAmjUkYIQ5r9CNWV
tgmiBVvw3gyiMgEodex29W9TH/IWitEdvBaQNm8QbTGaqh1uftHMERE8Qjp1oI4y
BWr2aLRKCk92b3UMbCu7mzHhn004MR8XLKCgAoTD4ecao6jpoYSlAPGoEHVN7dJs
pUltEhTUOzwoz9CPDAEb+8ss1IGpqE2lOcodHIQRDYMMzG8K1HKU7rRueK3dmLYm
1CyA9+un5f0jU0b2e1/eAGUl06y8ZzWLbMml7L7rjybCG4QKelh81MRBEFVZs7Tq
twjXiMGIQbIuRFJmcRZUMeE1xewFx72V4WrRfHxtHc5vr1a7K/r6l+QsqL+mP4/d
mcRx180t31u58JHKt7/Rc0U0/gD+8s9UKk/Uc4wzok/Y8nYmjqQrZ+vImGcLzz5a
iuNoTC/QJZFvpCX6D6BEMkazfo71c1v0uKJQJi/wt3R/SzY9Hp87ttiFpW7HclMA
gBARXmr0FwfB0NkEnWv4jpI+qf8wEb+3mMReRkS4DhKhO0uz9Er2X12dCer+e2cl
fzqKG2eoUowgYBXYJvVXo4avZDHdAetE0KsIdTskEv+aSeqT+VqEGbM5MQvT0wbi
y6i8aZ+/yI5ORuUGnvvvJ6OR+OzXetsNiyLLs/uzl+Pue3wRtkBNop+M6vdD32TM
UEZCzjvU+37QViO0hybU00nOwUS3Dbs00f2bw29ztMRQg4UY9yfeaT4jIYECrcpA
qt22Q9JwrZEB+oxRsyf3Bhs2UvLgubvUjbnrfzWoGiNlLdIQYXAKQSEAnwlYjBC/
Rj9IYUANijowZ3v3Cgj3w1lJ4NAHJdthW8kOlQEnNi73g7BnsEE+4usqbEax1cAo
fM6lGo/duDd8JE8MLB//MQSs727VVnkAljCTchmsbrFsAiPQ7o+U8c9OEUMC25oL
jIsoK+AV6WiY8RwG1uTgK0JFhA4yT3yTihyhqh2i+EI7XjDyQW0+4YR6yFgxCiF5
8QIcrlHDvmxJH8M/3f5D5hL9P6TB0YJCX3uc/sUAop/lLKydQPCZ0kX7UUGx1DHm
RmRaOHcDIG8Fz5Lk9D3mjpPIsGnkEqgAnxKOmwEP5ZihR5PX+f4dIkbhFQxwIcJ2
KUmOQl1P06VTbeT0z6w6T0mKVICyd5VXmMBwe+5maauQnxJALXGueB9VLp4eTXmU
aqcimmjN5dQ2RxTGpIcNQ1+mo5wOxKzJioflvJRoNMYaI1We54E8Dnj4fdYXnvxZ
3pDX52ar/fqU7MMXzJtJnldFx0bEB1kD2SM61or165GgiH5L9AUq9bmy2wfb9wxX
c/sw3VT2064TWWYIBBzBjerw8lRdGYfP5o6RC4yL7/JZbtGGtyMN9wqIoLGb733b
N5oTeWcF4H1TFe62Lcl3pkVx2ZwV5TlyrIk50FBNGB7QGuyxezjc4J6SVZnU8TQn
/JYIduz/h1n/g7lMd6OmcsRs1U5wVz1EJs72VuybGv6jNhaH/M3+jnpViOZNg/1I
2Uee3HiF8HZZrQdhG83Wn5mzLZAvAuVQA/oCkchGhlCt3ukiJMDQ60rm2HmySaOI
9s3r3Wm5fFOtlPml/iNxJGrrvp2cM9MtGwWwcHsVFg2lfwllH13v6mSvoEfCOHes
See0THlBsr0VvOwjSurunAPofINOhor1fJ+gX+HGSLuwCKja1gRswAZEWXTfrMY2
ofbZ4xEmCx2qq8GgFHfCuE/we8xww0hJN8sy9RAxghtpj0ib2o3MfrMclAbwxuKC
FnVa/NEpUh4QUzJ3642KP1gQFXrEoEIeCOcVSPzguHsMfAt8dq7O9Xz2uty1fZRI
/2UAvJk4lxEmBXtp8bQEr56imJ2BN6WrOMzCVXul5R8j7Yb8lBiTC6SeOrTAIeby
vtxug6BaCJhWlvF2NwEF1LHydr4Zl5C3n+rdeOdR/gmRcWVNkcdnOGNqHGlaAwjW
fmDsw+AQr/lUltZ33RQtCey3zHYDhfPo8CkFrG07TKWL8Ht6FzIpRB8yIfZU+uCD
tra/aVmQSQrNQbWc6/H7ahcJViEsa1pDQyLTR8W4PH3JwMT7clLvP83ji6Os7is9
Ka0LifuVibmqtWij5orQko0vP5+3WKr82iJSrQBYRLHRpnxThf8d1RfTe+guc++M
rgdND0372uh4JBCrA5ElJw24cSGY6vd1smMMnACsz2gzms3Zsw/A5YJP3qnKgW78
UnNal6jCm7Wz6UR3xBUsKOolYPTecp1Dul+uFIOrao+PBV+Vg0kOJAHcaMXt0Wxh
RfltA1fOkHya0pI0Na1r3LDIk+lP//83B0iH3s8O19YDtXfSNGx34lfA9h60gFTn
1/1Iu3CUV+Gde0ejwVi7sNE7ynQkzHrlteEaA+zW1GSJROzJm1UIiwXwgb8YGn27
KgroDwPMphWi72udyCqyAXdf96oWTWPx/+FHfvyZ0ZepeIpwyUcu2EGEKbVzkutR
m2hegHlAHYkkLMVu5xXv3mjfnahR+K9LruK9/TeK6TurhNP+IM3Tt21bYMWm9wZO
QNh8sys/gFBpYJSPAlOC3+zp0xf/OLRJlPamUd+768ORm0sUxtv6eCavHxSZEeFE
Iij7mmJj97AZ8G442a9Bwxico9nrOoY1+4wFou1ChWai/pNHmyWOZqrSbsLQdQi0
CjziFMX5rQ7N1ZVd+8hvDxhY1XoHfjy0tlrvn66Kf/iEFShpZ+L5LnIOxut4Iak9
v4EJrxGIilfy6RKdEwdy1htClZ0cW/JDRrVXATcmQhjEacGV67gMpTxGKlRjjgyw
7QFFLUV6cj3zCNGgjHrKehMt05rfl+LC+1gMKrjeOXPBHaJ3NEmeDwaNPISw43x+
XyUOSzddRDd79F9PoeF5xpXABtvU66kB6Oiq3kBJA/TC6uwfo6nFQDHAhCvnoxdi
e2W1HzDDuQG3K80QU15p6PnbABzlpzuWidQO0kM8sWiZetaUjKbVcrpTRc2wdxSj
2RF1NNyP+YEYQKE+axhxFps6geJsCRubu5MMYIkEaykXy87xXADNTShdZ8RkMCrk
cJmMYZBkXzSRiwEWJ+jVA12A8abDhPr49/1PhZxaBTYQWJuqNdvemZAK3FXDD4mM
OfcgFMDngl8CBDL0HiigHtLOp87EC9zAIV+1sgH7jd9+bDCfQNL4cNxieZjUcmB5
Gz3JSJJ3PB5IL3MZ08n6XRq8Y7dfKbd0s2CgdP1ZxqUZY7orLOUqa+3QyMjB4yrl
ttaIDKfpUh2bPTgsuPKpOkUKpdvuTAfg4DR5ikQipILzeVMIIlIVNpprgo1cr+Vs
h5UV4Ej5brRiRt3hz5HQUqBT/+mSSWoEqXBTmarbenvUej0hhJ6S3UkBCybrbYQz
K5abXakex+yI3WXcp5MdhJEBrinz1K7iBoRUhWoORkCQ+p9HmW1Wra9308rcfh8P
ZyY3o6X4vrgKGeILzKBNnB2n8USYTvB+azj8+/AhINp+fB2be2sgOs2r6+RbwmRg
+vaDh6aYGnuNLEG6AS0LHSWufSph0YcAuoCbsCUgw/Md5/qdcnhskkSoEFk7U3oX
e9cnqrVCmx91j8zjUzborCSJV8ight+mgRZLRvFSEJDuYDoA/haoPAd60bBnPMtl
gcUZXW4RuuJx54IRmhHGc1FQ/zsg3uB1wV6PwqKTDxh0p3Ldjroq5wSy9OBFCiqz
HJyI/x21ZsMylfVlQ6m4k/6xEznnl1ChdAJtqXvGzrNqR9zLu5TZH6l9RGYBJDtz
1R3pGpBCxy70nvbTYaX8Y4MzQ7kRGT5SOCczw8Splse6wGpRJIORS+tnBS41Kgck
mSwtKAbJJHcOECBBvTKMOydd/WYMwRJBP+Y3X4E9E8Xl74V/tyOmi6qkaE3HSMGc
92oUuIxqeq5caHBdFQNJ25nav89Z0FprXRbDgI5o+X92J/rAWeR2fdoX5QsX4Mz4
R6eIkltBUmazqmXtHMBGxcZfEXSLJxIGHaYoQ40/T172JNunxRLdinz2IBGu7iby
0U14P6nJhcmZ0nC/H9mW8hzyLwqHEs03FbOwFKiuglrSu/4/GIH1bkun4U4QEfw9
W8CziU8UGc/3nFAhg54qplFXW3Gz3DOn39GWIdQWgY6moRCaqAoixmpjzOG0jc3x
+4gtdzT0u4lrwac04KReKaNbJ0BrDpYLKrXHGgDtTS04U2h4QMK4HQRw5TWyQIEo
CXgBSu9b8flyHNKBcCaN84lb7Px+y8RSHlDAYp2DFhKxg7G1L1STgMcBwgRHBs/s
pb4tl2mZQO4punLKpb0uWJdfVX0+vOHLqUBh1MQff5WBTqyjTW5cZkIhTX9CvxMx
99Y99cAwAdYvb3FLHkGRM8+SUktjc3c2r9QSGjHbVb9ChHfVtLSTiiunVEMP0wGk
1S0Mi7i5KOjSa5edmvJshNK0h2LzjLzYpHduBCTjDIE+/eHzuTX57euxhUyoxd+F
1nF1tPK4tcAQoHmwg+RQL8X3xUfd/tf8+BD8kLmDnBCYXgg9PR4sTPRyPY3/ETZT
RlcZGKfom96Sfw3RC3ig3gnzBVXO0eeI7U/GH2WFTLpGANSt6RBIBeY+d9PmfF0m
+qMCoZoo5kB/dLVfU0/+Dhl0nC2YcP9GoYhbDX6jWOPlog4ZNpJVam1ay7D7vPrS
DygVNwY0wM48pWoFIFnVOzMQkZRXv1Grvova0DDIC8+GY2tj18ZgryV8eB6TYi3n
ilBfflNmK3A+qIkpb94GhLE/rMu2lZPMyJGwURi7EsdqTk2UTPuW0/Y5e3C+57Xi
z3fGxG7zyS2SA8zWP1SCv5BnTmXOy+a8CCUhKFRidWQ6kqoqtibxhxy2hnQM9esL
KewgaAaVMVLTZtbTyGn/FeQ2cA+DhM/CTmH+oJfDZ73dwsrPB5yxWDr7HeH79sgF
dtEHqzlCcTg8jGoJtxdQXNYBJSj9Bi9rUhG5Nq1zzArOZwW1DKXrxwLUoDVk3uSS
e3wPeuSFRlNolYu5ORrJ5tv67im28kxN9w4mpaVj52dCU86UbdHTLFSy0oqAMDPo
6C8Mk8Q4jrt7mp4r1tWHD0jY2UH68JbtQU9XJLdIX83sKSad9v53135aaQwMpJPZ
odtOTzHWHiDMIdpbLeCuae20cL/k603d9bVX0VuL7/PTyvqaOnr0qgTEqICNRcss
FycVJyBpFXpwDI5a+ATRpaQKIrNOsV8AYM8u9pHmG03uVOF9SLVg7itmvLiYBdNz
e164PNSBbdycajqLGlrBDQ3PjHqcY7/6IxCcAb6Cx0SgRWcTdgcz+HNRNRz2mEF6
71DYyoETAO4lPtg32LtxNyvHwmsZZZJi8BmHaEDyZZXgxRlAet9CnqUXiK80swPV
YlkvcAXzQ3uali8l/2vlYpeMHt65mM9YboRLpkdlXnJgw0CfgFEu2O2tkmXpyNmF
l2FJESngGmpQDx2T2JzT+poxnOnuv1CryoqNPvcL9VHrQEHhXScn+ito1a4WEMQ+
6PbIHH9Ns8kq44QHDhGQfdQsdKXh3rxofjcfFBKruMZU96kgeCYAF6QmDHgJQlc5
RPhtUn4Surj3q0HhCF8Koipt3H/oylwuhKG9TuGVaCzLpDPOtQIBDuEDHgps7kWL
gXovmloLn/9Fb9e3xM5v79/m3vWiQWW7JyllXBha1RTsziacT2aXGaRFR4KH319G
xXCm5qFnq4Ew3mMnk0+4QkoQbS/73ywGP0B7iOoixBqyoFKTHAxbdGU9tVToIrm5
mw5IOkHKZGYYazCfoeu1gE10fpQnBtRGT11NMtnVztoYlPTw/O44K5rikhHkUOZ7
HKN+pVyW8jmjKsxxW78uLBa3B/u4BwWOhg/+Y9i40pexd1T2n6Gi7EVF59iT8v9i
icJ63R85tEe5F8u8+gQdagIxaidlQjnudRbPUZbXmpSevEZybbfaety1xNVCsraw
RgBmdWb6HCYJxa4Zzz7PMkL5cPsqW92Eqe9H8NFlzfBJ00NUv6BJsXIf3DmG4DG9
vxWlGUoLqOSfo8/j1+xESaMo4SEci4O0cOgZqXQdlEDpdM+b2hAxOckDhgVJ/Eyy
FigawSm8hwtvmm0kLoZxDVTBxK57fH1e+Gszi0A7hmBqcM4rsgogEHYuC6Yd4Shl
hiyt0q/8ud7EXEvvAF+lkvD5iDcUg1ispGkodLABPjmnarUzl3tSY/hySai/vrE2
0pYBBfcB4GAK6J05iQ2P3yn+zTUmEi77+msYJgZz613Cyyu3JF+Gv2vMqgyx+9a9
imK97QtlO1FAO5+mwGiGQwZzyEFnqsLhkZrNQsoqEwCWI2cBCzzQeAK88GhgIYL2
TdJI0CVyw3DeRO3kReG6t6Pzad4gjEcyLwi+6bLaF4wSHf4lpAKpt/JvgDvqvb7C
Cq/dUs6w3jE4sXc2xvYIpQR/CHDn1A+2574eGytAQ5QklCWVg9dwnQD8BU2l2qKq
XPr/84If3jNSWmCxKagi6Fkwzw6vNR/qvRTugSjoiElALN8KneWhVBg+N/J6Bx/K
yk/YQje/5BFEuTLg1+7hvSZC6QQ+X8kbyxJKO8DAMfLcdLCAdDhVD8x9uLD51Q1/
XIoijd8baVfghdnF6wSXJVWYDqck9GRvgN7I7Hz7fsG5zWcHgMc5ZUNdhnwobWjh
SfMmhisIqaNZ1YJibnOVtmaV3KDL34IQJv15PCD19eWX5MLJqI5emxQsTtsSngiv
W6dC1aUMgnm+FufTjvJnwRKIkk8aFnE1kKxgRUHaU1uXWCBAY/zd2VfSKctSaVzc
0VlZhx554zG8Zr2RFjgnuEzmDZDEPtl5+NW92Bdz1kTUWi5baTFxN1A5bcLquui5
vhpbq+Bdb2ONPfqhQFg0LaFFdRA9vo8KCZlnhTa8qjHvXCB0F6oat9zH8XIZVIAF
fGKdxT1g0szd4NpGmTtM0aU4lRlrT6eFTRQ8N6xG9J+1z36fCoAVfQC6+NdTEc9x
9G2ShvFCxnNj4GNko1s2Hotbed4AeD6MwPUX45OuoY+ZTQbECPeKoAFX4MsptQ/f
e9Qwo1t3IeoGHfNgRW6aaUj6Xll4Y4GAQtdYTy/fz1SwicxWylJsFp4s4JBkTCrq
pyzrcfFvEWMQwrewEGthUOUkjrdo/CsjucAd+eV7hVOs7GbgmTMKFzofRnbo+kL1
kldOIopfc23zOGhBR4F6y2tK9GrsQPwvN8+T7of/wpA7HHxrLWV673GCWr8kRMBR
HXk2aQT8rCN8q3XRqn62JOft6HseBiuf2ltsa8jpkqspkWM/8mXqaEBbCKY/+zzy
wJkMtkklQlZ4kDy6zyRfOVEVgOUhf6CVCkgwNg1CMhopB/UR+K0wh7V/SlRzlghH
IapXCp8qKdC6MlWghHVwOUCWMmYrkgPYLqaHeQHs75D2zhDsWmPUTJLf81ApKKE2
4SSRkGW0ZuqHTa4pOVESDYYUweYk+ZwrIm0aPcfHOFPQQeKEtFdNXQ/RtvoSGqr2
D+kM+9cU1KboOQIQptpqSIpQhllmgn8lOqD2roINdX8m/e67dmBmeq+YDrU38/qc
USzwblRoXdt102sAzZuAGI5g8KCelqR8fwTXexQln78gideZq009pdDt0ESrrvgy
mOw915xljNe0X2Yp3TYQNF8v5n8T+Z0RFizCaKdXIKV7OdtgX/X1A2y5ZUi0Z8hj
d9/ZzqE+ZEpLxfx5Ntgk02j5ZElLKiXBYDCW4wGbHejLGUhdqF6if/wGFkYIQiWK
G3RHcEbNr/Z2plC0oRTguuARER8r96UVotA37xRrvkxSntWwOBlIYkTi5/F5mKfb
Wlkn9bfQ0ogqqCQPCLThnK9IFnnzWYISa6u0ApFxQBEeHGhx5HWw7QNhIqGzzxJi
3rPZr5W4o8TwH3HoXrGkqZnqy9++q2LJdKVmofIAl/NiBmRiD4Edxn9XEeFYvZBU
zB+lrZ/98CA9HjhWRSEdALJa4f5YJ/dm0lwAuT/tREp8KTXRKTWpg7m2llCnky8/
fW6J+YX0RJc7xlxg2NbTB1YI6LH/lSV3c0t6tMr6VpdRuw1eqDUoLfudqTxDeWKp
cvONQSkjGrsUQh6YywdJBhXP4UwBmNx6mI2tsHd0D1o14VFlAFfd3MFrOGGWS3qz
HdGZ2J62R1iapsm3rFZ3zNUVzmYhoHPlhxAEd2ENuHfx3bc4Iri82zMz3t+8U4r8
RRI7b8hqQq9hs86sNa0Qp+60f+4YaZx3N42fhJefSuPXym41oLJLx1D4p4MHta8t
xTxvHyn2Pbrlo/jCL4lvplmLl45d5n1H5FUV2KJKGrl6z6qPqFgnjQeRjGYgZ78J
cIJ274Z+egoZIDV1oYdaJoqwYk+31vuFiN1w1xmv7n7RZM1SFu63aM3Eytak9meE
6cK6EMIfef0YC2FE8FOY8K7YqWIAp4i5ZnlHbwGwaZ121CO7zopMIoy3KjSwWVuB
mUAN1Y3rbL/PxpEAUJkwubosx8QGWDuwA9n9Uck8Vjy/hWfJUTVfb5fnQdSHTeQx
koZjUoFxEoT6pDNtPCohcE8z8G61fkuUYy0NA8RfnT8lIoQWJdALwxbEI8pQGHRX
qB/IGrv1lPptmPFCJeEJCzCdfqCaaSXHSHl/CzzTvxmNkpIjwWkx/8AIkaSBvOXB
c8EqN7vuXH85vpNnjQbGNTVaIGCpVkIiYbUzEdfQ28/xrS8TVb1hNiovdeY55ccB
R/hyMM/QBJXW+o2hzZuc5ZlewSKJjfXpe6xAmYoX/6mdS8w/XjxxAagaOrbGteYE
Tg2b0vGxmndIcpjNO/qb33xiuFLd8LpOPuH22VeAnRS/DUFAwfydUFyZxXMdb03N
2MKdN+FJnp/1YRYeZniWYa1URhZWmjODFMqBPxtZAs3nl+rqXXKD19Lt16F5crAn
kmnTf3WyJtuTkvR8TebfK7cl4fCvKO3/vvdqqAbZaBrApgB1awOPgB9bFglqdg7t
ohps/XrhzM+zyWm1N6m24wF8rb22+NzdH2CevoEoPDOBizvo0WdlTrr+v57T0P6e
1eu/iG0JJgtzJT/UG96mrWHNCbNQaZqtbEWrEkzhNhBHBbYyp+Dypu5E8bksXutK
MFBkAoGHeySPFp8dLXS7hpQKeGeUp99jhbvVZYDMV4lDlvNYamV4g6RzpLA2OSvN
K2WCGbUO0wtIcI9Av8zWnYTpXeJd/KLxrRgmcCNnV5w5a7dOwdbEE5j16Yhsmw1D
hs2u7AwEz76z05YXAEQ9jwxt+X4vrOb7CEb+6z0gex8fuWgLXNcngFAYhFKApoYt
C0pzOxY1sgbuMry+ABfopnWYf/fQzzQ3S6s5OZ9sTQDx6fF80b3ktK6nAwL+ORQa
QHDiVRkosJ6vPTMYlKF4jdt+9KpcQGCnfEHGOVYDB4y/u/+2ORXklaBSXmtQeAm4
Yz+JtbFcKDT+Y/LHKE2b0IcM0MPgXPIozHq4hQTOXLvzUhJRNfwL1oSsOMU71r5/
RDhuR+4GaT6KAI01UCx295MoHCMWP+SsNBeNW8kaqMfgZ2F5MMGD+3gl1UBos39v
tChZqyCGhyKWFoTnMqxgmtssDzg3GbKh42LVaZGAqph//gGNOI+H9uwVrS/LmDNV
i0ZatyR7R1w9VhfSAkzRbROQUG9Oj3u7I+vRxZpCp17QB4Pl3lmWL9+TehTbEzQ+
20l+prf7UloYSFv+ojGouLOMd8S5JyrIESi0kngXJ2V6GFSnm7cdFZS6Hn+Klx5s
DA+wYo4fnMdyM9xGY4bAkaft6a4fYOIFkL9c5hrJrmYpAm2SG28kavwnUbijkouk
xTv0DonHkhLTpSgSzE3QA3Vx0tzAnFxo1p6Cqx7kzdHvyc2KOglsY5uFawH5u6Hr
dNAmfn1eEx4+Aom2+2mr12kUNqLL5ED0Jn26SOYL603t+dBfL99I6KhouwoSnX6d
58jCsyuhqmlA2pm7e/6uj2hlOoZfjKgBY2asMVzJGnw0Hx9GT4yhXOzC+hTEZzId
CIYmGLOXuk0aXvHcHpKF/jwTt6A+BchLBd7RXwxg/ftkhR6V0sAwoGJk1DmvOQLT
owzbFMsP4NRxtSdEwnIkS7mhrs8DKxLg7E4rLQRQJs15bzX89O+sFizRRA00MxLV
cKef4+Iew2/KhDbsIW3AN0AX4htuD9PT6BHYRWvkQn4dtF7I4mUxIdAPHSKF9KVA
YlUxtKNhEgPq/wTYQOFrKq2BFXEDVdQZ8H1p80D236YV5EH6otpSP0dZFIM/E3aM
MFxRQGVf9vPO492t3Z5rMF9GdXtjq67SSyiT3dtXHFPrQCxg6SLJ3rq6ACCMamrw
VFtx7naO9lumrSXLZJnjS/IcjXdtw/qjdXfCDFKe6Jk5A+0sUF8FSyRASu9TNlE0
nmFDkheBhFxpe+awfKNAdgTFn5iL+pBTbpoG1Wz1hvg3vfltx8Ms+HWPUkuZrHBK
RZ/dXLcHem+nU00+FtLXfMfgfw2jwp4DNEtFreJjGGoIbFo4CdqU9G2+qaKZYUfi
KBCE2NSo3WSuxYHwechigKI8FdTB701bbxb/82WBhq0Ph8LMZLq8adovC/v7oDEQ
jRwMM5S5DvyDgHFt8N5tEuMgjIh0vyWNDV+LUfT64SOJItVbKlj9dC2CmICkFhqr
79g7WcMFbzFFCiKDlGIDb1r4wWLWzMkzS5axH2iqLkqcx8jJSqqge1pOJuku7d46
OzE/cP3VjP9G1IqBrhplVOD634nCJ7X5xwzDl0WL6xCflKYlLXbk6/0cssW3UNZB
w0Dg0fkFVecuwkqeMcbGqNX4dAvs6UDc3BJS1ISnOCUUgbBmZBgzMh/GRy7fJhME
qd9FfelTsKlDyxcd+RSzo6d44GqbvkQHuyQBbewAeisj67Le3SBXK+HYURhsUhFy
X2NDvjZkbGTFY2nCX9MeDzi2Gm8r9Jr6t08DECwF7a6anGZg7EyG4siT0p0iLhM9
1BC4vbj5O9BMp4wyxZyjhL5G8fvAMm+UcpKT1nIal0kObkQRiO0sY54D9curRK9m
3/JEdxQrCaUgQgEHHpiI3iYjg2VZKeSzEMpzVl9zRr0BvxaQFG1QJyCRPCOk6enq
fueVidA4jB3UIzsbXHPIzPoSRJoXMET1PVlYUesSmtPvI1lQBzrVibPiZtqNUVaM
0q9F5igDYzO3ts6GvbvKhuQPFYA1ERH0qhlef8uo5E550N3o4yDMGdFi3Dda4Vnx
AXEEwF4wk8ABdjWVK0zGlowNDah1vTWWGsrIC665lBpREcA3qXtrwX8r/WV0fzry
FsvVkSIkX7A9e2gno9onAYGPirsXvsrNIqcIl0f7ptE+nki0WcTH9c6UZtA6xifv
u7xdua0YBEygDWXcBWGyD3aYneFXTbH+QbjYNR75cLEp2uZY2Qm9JToTYCzYEX/8
KJ9QmA9TLBBDPJY5KhlvNWqPpYtxGcfczXwkuSCwodJoq2NF7kbV7E39bIrXLWBe
jMgZt90wDlmXI2beKjRKfBBB+bEKR8fD3mwIf7hNIjOe40CJTjmMSrGeLNDJSPbO
0iiLrSGUz/oeOlqTuwuKFE+8g4i3dmtAq7O3q9vWoVIxQZsFfPLi1MIoFnntJM9F
s6vBBOCJgXhPWzKP2Eayd5/1TLzCKVE81ZnpRSyja3pxAM6lUvBYtLv2PCQk0HQ+
/l+UwBS7F77p1Mtyu7AOROAtz4UfdgvTuH6QwpXLH15hHCr5MolUtXJi4Oj8s8qN
YxkshSUzArA77241FXsXfg7WVniRp35E2z1YXZjub3GMHp8rry/f4Ys8ARkBhHdj
H53p5D2XdpK+x4k4R86bfc5lsrCn+c1au+lMEGuuc3et1q6KbsyhMAH2CTxSqkxr
TXmsuFNFR3za0BYmhP/UoiOPlDFGLMFxgsWTLQcemqcV7T4S7wtwtUv0h1yEDWIM
fcfcRRVJkMGoZ2qNhy67cq9ZRo+RVfV4TIs+zeZnVm67wg0IZ3beBBAPx1JNlZPQ
FVLDaLSnR3AWyQFu/h/qYjkTf1YOAXsMQ4Z2ZoL4JPCJ/h5YI2In4vrKlUrTkLgA
xd1QTueeaH+APA+J6fvmpyY5e/20Fecz/l6YVddCfbl9hHuwZ1r7Z0h7L+Eur6EN
99zxV9lW+xohWraG+La9/xk9gTT7hyexRNxN+EFrwWsK7jXEA4+hga1gqiYJixht
di9VedE04gA91UCTwDKP+RwXEBMQEJBh7NQAQRa4eO5u0Q9bh9r9Bsc1VO6zmWsL
RH2ndBz1PH+imKrBzl4Uwnojffh6BO7w7DBMVO4mvaVG7nCroxDQFz8whBn3yZ1Q
oboaja4Bw3rjHJQvJj9bPoloOx5rC0iPzTViMWl6dWsCF9gon3zfv83a3Si7LgU8
V94SUaAdTmcAeJ3GusaR85Yur4gMfvMnX/tLHtjvxtXoGFib6kGVXzNyyITj2qhw
hJVIO9xMEl2SdgQKHUXdPB69rVhz1n3d1hFuKqGbMRRSRoQoZuwhirmMD64udOoV
eHxsw6SHtlh1SOEIxEJOmEi8WeXXfOjz2MRvhG3Ysi7jY9QCpPXXN3b2bUSaK6CS
ST4sMwd9EllDKb1ouYx1WK7LdC0HtZnybUJZ/eRyIYkOsta6xAt5TN9yO4xCICDy
2F/rSDC9D+hfRi7c58O4rG3UWdJwktbx3qa9jVKutXqOhpctsUJamjgKEHgzg8E7
Zj4IfpLnonCZ1z5D2gGU3O55BWzws/vAF1cbPGuFtv0gXBgXpxYiBdoRYhDmy2ii
m5QeLJWisfqQNRKjJTAiBLAXK15lQ2IFmrTCUT2HRzUVE0W2m7grNauVwiE36yaq
V9+ipFM6QqLw/43g6hvo5+Lg2Fp5Jic0iXOsFA7cj0kHdU3W6eT+jC0S3hTSWDVV
a9+CFlYOQ0jJHptYBgu5WxFBC25EMKlgPXL/lLgGarGv2srHo4PG7Q7i3/WeIxQQ
YYppEasTlRitjsTL9CmIQCbsvTq9E31We4t89ukaF+g4NRp72hzwpJfEFEI4OAlN
WJgZxlRUm0cID10MGTdcgSQ5YExKCG8vCfpzHfyGSY8vHfo11R/hwh139saFWG80
1BU/J3Czxz0QKyAZ1Ni+Et8/oB4hOjEdy0ngVYdOs9JMpHEctvGbUpX3xQzsThWs
L61rOOf+spk6q+t2EvHVLR/MrG9aMASxLLT7jOw2YbNW8YhYNapj4tJgI7KVy7NH
DHA9JC8BTJEezq1PVBPCO45XWGtW3SYrWnyFLU+zZkDsEhehnfUGB/wK2LqXUPW7
DCi3DJz7tPQmJ7LfqbOt9misVzEO5+0o9cexLilNMYQ7lCEo5NDUWBxdmqE+Mkov
VjDdAd9YwTnl0E1/3yBB4RylvK4SHvzfOEoTUdZcgdo+kGWMyQDkK1LrTq1mgc0Y
ux7NrjWvPZRb21xT6uML9sDeIlby8qOJiFIfHPG6ZRlE+czqzeHcRO3/EjhYlyrH
GvXO07gd4hDEGuQ6HA0jO21vNvoSSUbPYyvLD11tnWRTLoymAKnxxGXAYCxrSlWm
IEnoCVAv6AWKuwzerJk1Pt5oLWy3N1IInnEJW7WqgQIRnAsB+Tm1okdgQOlwPz8S
zPMilarmuOxkDRDFMW9k81/k+YX4AFRjUW90dfjOY7vuw9IL2ultsmtmjkeKyoZQ
Z5UqKGW3h7uShWmvcl2in+OiZWE21p7cHk9OjbFhY0pkG2EN5Rpn95j0xihEOn0h
/i48IinST8z3N7K6HSlsIt3yc108M+EbRJqKVHkT13xK5pBtmPpee/J9+nQekBOJ
wVm0yNbKNlusbke07WTHdjds6fW4XTQoZaulsnMsOZWWIFgxifkyorGe+QFh2erT
0LAHwf74mbeiZ3zYIQbavlefrkyd2u3TUU4Fqb0ixb+RdhXdZjHncyPpci8oAT3S
O6LSuYd42dqdgXx+SUlYteFqUYDpeVIh6icPfscQGf0/QsuBof9ZVrf0MLOUfNlX
8cA72b2rioXwoojUrWb/vfUvwFj7wvNqSHE3MZuuTQM5ZgGV6sQdCCKUsRNKMwH1
P0GGN9oF4LqtPu3xRTBV5W3yPvUv4TnXW+Pn6LAAaJcV4ndbkk16/lb5EaGF/40v
hThcgg0ZbYzV+bqvWVA0PaJRck0g2o3HvMiZ9C+ND/rHUJCG2R1DzGfwFEdDBa/2
FcEc35LCO7m/Q1KLFbd2c/kL28IT+kIxAVvRos0shBA/XNP6cFYYxfOVSp98tJKW
v/SAptM4vb847boSwg45qUmX+UEqNHDXlVS5S27R6De6PS0bJPfGjf0rL3xFGR88
Lstn0BszShyk76zzF0BfewXmUUvqsmeseJtLNARq5DM3RLXzueAO4nzVPIZKMJ16
Mkfn8hE07uOZBun2PB6cTMcolWDojvU4e+TCZzcBkkTKhnXavnGKukk8Bz+0eLUh
hQMofT2F858uLeVEzGyu1btEjSPh/vn7T6NIpg9zX0cuhrheIHtVqKiU81xTMMas
u9BmuMeKwoapRUuG4NS/LPCydvb8k8/b/sZIHQs4ngP3Hk/3Lxb94DnFuWAVAovN
tBpxna/RC0ovqvmxEsgG1qKFaK92sWksD7eQcD7oK6gGShcmG4xIqFDZ0ce6CcVb
zAHlHGYs8c8zoVqpOdLfS0j8XDyMKdaTSA/x4Z9GRXV8UizbEQmuHYfGCcZykUxg
9Q6lQpE9qK9C6x44LMEuU8JJ34+RhQhhAzAH4QCaY/euSqrSn4GVhpQHOVW0ABqI
egBumEzmxV2f9b56Uu7Xo+6w7iDBwDylvOI5vUvDA9sKAI2Ch+1skxnhE9HX0UUH
9fCnSoD4HjivVV/3J7Gdl4dLvRH71EOhC27Xvpng0YxrClkjBgK7gdYenD8tvy++
E1cpM3L7gshwS3UAuJ1Xk1khjcXJEN34pxkVHnag0FBJvboolu8TgQrbwyPLvvEA
zDFvWklK29neuxeFyZIi1Z45il3sZJGDVDPrdmNV17+ma4ztKjW7K9dFlghfl8ye
Sph+PoaWOwnl61cdImYW2rjiDJNdGrPdf3i/fKLG96f7zPfmJQPZm7sCAcF4sbLV
mU0C/dddfCQvIZ00TrVwp6Mz3GarWk5d3rhpErcdV25kt9GXu4UsFAaWAH+L0h43
zog3uFFCkDz07qZhXVxrXjae8UAzHBg5N8d0mHaIVKawpBea1447o088WuXSLoF3
bdVeeTnpwXIFs4v9HFayD9RRfTpVgyBYR8schHbhaZYr5/5dgJJgae0DzI2nVcOg
0sCOj/dzLbn3QtL0ctuIGEXEVAlbTuU1spCQjgRXWVkbaZQahVewmkruk/LIzK3z
ooU7MOSdaZFESMsQtF+8KxI0C+lzZBZ7BuZyyS0qmTp4OXAsE0ALldEKRAhddzKs
2lFzd5a8K9mC9v8in70jVaHeRKlHxGl8GB+nFZhdOkCMd6vvSpQUaoXWxRa5tvs4
ZYtc5oNduBbgYZNsCrAd5cetakkLLUj48ftDK39q6K5KZ2JkDyiut8sWK4R4e6t1
N7WBCkZOo4Debf7kRkGmFguJzPJDYvnjkE1oRo76T6noy0koecrRz/jJyfKK8bSF
hRBLyxV2Z+xXDCaLQ5Oor87KMzVhk2xHgh3rJmSUYLTEYCHXEB1b0hyzOB/0Bbt2
IKIpGbil3zdX/GjWQuVm0AlszzFnYY7ZA4qIQaIO6pZbZvQfV0OG1SaAtCU8JnSO
AgdSaADRBkmRFbnGNuQuO16fVjac/wbSTN5g7aaL0uMYRhA7E1ps8tutisnzn0Ng
Hu0Vd4lAfMRpYoQh9yatP47T6mcB51BzmJ8bR0q0d1VDDGipb+0YW+PzhpWbNsPg
AzwT/Yn8Ws1Wf1nh9b2T10AV4+ffxgHyijsEOumet5tHqwxzfNEXG3odUH8/kYke
a0dyiiVi/ekeJa9Dv9BRDoewCgOcvbdaPkG7+8L6L0y/0aUyH+6LZgbr4rx3gbvb
EMEos4L8CdUnK3TFRQkKDmm3nvAYdDlPeTrtXacVRHAKos9/fV7kQC7mXUG3063k
rX6g/XB3ZFnBpUpwk8llgTetVhmlOXKeROidQe+IhTs6HzsweHjjP58QxbrijDMF
YMqpWsQOPFS8j+y2eb3erDSW7aA9csof6qygC8jAW72nWFkdgkplyX71gVG8UuQO
Wmg/XWEjLrTPf1xVh5i7fybXpxbBraD4WXZqcfN9i6mecroZtHMRjNOVuTxrB2MB
GLe/GocRSpzkX4djqYsT5S2Yg4atvZYF824SGO/jYzTieQt5qnRD/WxkHSdmZWxB
hraeqdcP3FNTdBCzo85tDwWcQQhXQZ5ejM1n6hJGOtPpWQgFuCTIpESRuEsMlSbE
6e3e+xMlsugc1cvT7eACA1jg8XMI3IWhWnLFCq3YeW9HtPvx4LEslKalQGpAQrhv
0DEJe5gf4Uy4HRld4jZe4+3tCv9Og4HbeT/Cj7zovbF8dOMJEivs0yFyzkarChdh
CxfG8Ip6FCYLrmpffMpLB5/uTUJWPHIjGihggwxRhz7nkUryaTqJB0JTWVyvIRNT
C+rodbYNVCIJmjR9RXB/i5MFsaGFCoM8CGsrbsZsNkgFz9Cx3rFY7K+LpP/vWoBp
xSCXy7jnIwYn3hLxKMWA0G+bxfXGt7xwJMMmRNWipGdFM336JCoMcFypjfezEOqs
VeGm5TDajr4BXwi0IUQZg3ROaKiBJNMQ7VFHbmmupFLbedxSxoEoAcBqr6fJoZvo
qoOxjMDs/Z+C7wyz9XYJgJl65SQx5ZLc5nUHIgcj4Al/5yBhl6SvUWVtFVsZ4hb3
9pabGwt2uamzCNaBwkUL8Hv/AEMueOBDIQIlZPKcTMwMJzc2K4xtuxxfurn1cn3N
ZUzg/zhH54i+8/yPLxxkS0UBr/3mrlTOCPvviu3tuqg6ktig+wBlEP0pK9Oz2Mi4
zqWU0nxPas97T6vNydDL7mqsENnCoVNSmsZpjvVGcKmIHbyvKEtX90QhdqCmUKic
PGo80IiNHUXjNqWnUU7KOT0ulbMEfq3KBALpsykH1EMr5yyI+mEYDIUXJQCW2OvI
g39ZHoT77FJYFZXk221i+YWOngw9dHMkm+G8+aIF7AIA0hDyQxxzncwLr0vp8aVb
WEUj14IYhIF+ukqTSmCQe/ciXqjRu543FOPNN0waUSEKs0OEtsBNOeaNYhJ8pNV/
taPZcHojlPvdwX9hI/7TA61s6RCx+py+DZ2gTC5RDfxWXAnm2TOqQcGLJdm2bpB+
wwd6ryJN73ZPPrU1BD3fkonvW3CIEA/TPhQ2OJwte3iXAuGvfIpqwR8pfXpqz9AE
cOx2usaOnkT5O0XUp/dfcwTJmmM35ZiTuK/RdREL54dCO4TOt52l6mAKk167RFsN
DvEQ1UKGnbzGmHgPX1wjyPe5zKIb4VMiOd3kOoBQHPNCxoiV9+kiIzPtX7D6kxnM
wftmMKWveOJ7mZG2ypqd2DKAzAbm0LwAcWpKo4QEZzYsVUS5dNGe7l6grcueggL3
kbGw865qpJvaJTqX7bmOKjg1UpBfWnScm8y9Hrb3AONVyFdZP0P6TFaXwzpP9C5S
4bDha8iAlMKF0BIgIwyAff5tsILmuSA0AN2VebeMywYNQ6n/vxiAUf2si0uZNTrM
JRloKNbZJ542IcmXlP4n54onezBJkihsD3BhuNwEQx9N8MMqQ4RbTG8AP0R4d9Pl
ppsRgzzcHyV3TgTTWdCaTeiZxHTPrF3MErnKWKyJoFxuXYNsNlVemU7lhTOh8RqA
XX/niQHin/w6rAIu4aJBNOCuvKKdeTejHB/0ReQZcBAoHU1/Vta/GMWa9SOnS2SL
THsbt0hHD8Cl/ohCQueZ7GOp3VJJgqMsKtBLE0h0JPR7pz8HKeYApkTBP827kV7g
2OvncL4La2U1wLPjlXr15j7yfWAKqkr7P6RQvBQe9hD1YP5ZLtDPWz+dRmEyesl/
wx1CYZTCsDy5MgXtQqRW4gx7uj9EtB8MaxMwMrd8R0LpWA1sROv9FbmbYi1EGTtX
CU2Ths++jIME10iVUlZdxs49m38THVSMmaUd4a5sjiPQozTYkS8lVRRchsPH9fBz
+yBBKbTbvEhKboD+5L++YorlEDAPVpztDb6Yr5QSB8ItHgY9MnbabCMSjCIcjoCh
jX8LHkDq6Yv5YaS+uGd2XeqJ8FRQadkXWA7ZwBT7e27ob1HU0lfDzuz7vU9rFP9/
/+JqgWApknv2qwkoaTUEzqEHDKMp9HgZmye3TDtfj2EjUOIvZWTTjxYH7pQzMw9N
xVlUyF9KeiB+OP8wAf1lOIW0bl0zSvyH3v55CuUterigA2LPLizzCtVRlXk5p6nk
yNdD1Nb6yelUtdU3Oq2q78gtsx5P4M7xKn0AWsPANjQ/WY16nsSsJRsjnyzn88Y9
pFmZD88gLc77ybn2MSyA6aeCoCxvpYh1IJUBDkRjNltZ3c+1IZJq4E97kqdwqq9q
p6/59gs0J2YfS4zLTG4NUOE67SgTJhaLZLjQ83EIRi7b07aihWcJ4ts+XSKnGduG
aDLTIjzN9egNnD1k/8SNXsi8shbZQeyoTmpOc3BDpKZsduzy77H+BuHZDMro1Hmw
mZZa2lN+Ge7lhS8HpiCOBk053Vzk8NjCV6Twuwgnkfk7311qIMSc1ptTXQYMbFQi
0kWAiDNKRKoohZa5cayD4wO2qxMsMysimKiCisZUpEIsxRe7d8x4XFx556H9x7m/
Y/uGszCzmVQnNVOiDnoD1spyUgeYYu5tApRwdZmbV3mCGtM2TzHW3thJCl1hXsHo
slbI+NABdd9dOCQ4zIZGJhfGAcSDJhAjKFxccVtUsgLThS8DWfqrjJIyRSWfBI27
E+5yM1bQHfOVmOAsgsASQOGWyIH6CqKqOE9Ybch9Y3TLDDyKHAfeOBGposM6kTGp
X4ZDdCBqoGaODwGvEK52ZbYcQv4X6uBrjv+aofLbV+ity+m0P40JB+ZTJ2/gP2Gs
ikfFRLAobu6d7kb5xl8uvolHDqz6M7wIuAldfysYcxXVCurJV0Zs1eVykjyThEGk
qLTZZ349hDTHKYVwETi1eHD8bpEquhLIUB+ja1zZxmKpFno27w6ZMHRBJ63Ya+9e
uXdXfDIT10MBxh6O0y/rJS662TLagmvcrxKMza8U85Uw44+f9jARlvI2eDmHJwIR
zBUbLk1a8oEf6pNrcNAIaZPT1hbBYYrwUK5RnDJQOdSgwDrUDbZIZxCh6U6hYReq
aMQH2GVuYr7mRSb2BjvHf4j4TSD7oKYOVC/c5kRHX8QX9q5/EpAvu+w+L2P8o5Iq
dN8ljdsBq9TZEtos0B6WDUPZ2IEFNLS/BMhUog+bG8R5wScUj7zMl47KfK8O1QB+
NLojQMH9YJAWP5FpxfTg+x+gw6nwcJh6lwne7sYGa/iS4FNHQ+QtKTvInrdXuI5P
nxorGOYH65/krwRGKe21jRQanuZL5Qr6AYVbv07xfup/FYiRPDYwzWagIfUIMnpl
8ejuUA08Lf+v8KzRS+4m62JCxkSlz36QxncDFV4IoPbQLyk4oud459PpIc6PffJq
V2tWm9wcrWIoEhT6jwbqLYghiVV/jdtkWG+eHW2V4tYRbBdn14SlHfQcx04lpHcD
jA+jd6XS7Z57Mj0cKha6zUvHp3c+PCfcmkg574+0iL5/DF3AkdxMHAoayoUQHidx
souGBw8/f1Lbcfq4wgpAGeE1PyTvCk9A6jDnpKa4/+lGxrudqMKTVuEa3TzVG2nk
xAJYXBcVvhomNr+X3r1t6QP8y/SmCuk7305yPXI0NWvxVbQEFn68qoFKi7FenwHS
1vGditATqCWeTYYjNhrWmvHrlAWaCz4O+iew5dkDNPb3dO2rR5FClEb2yCdhUvLu
/e2OWlY2nqP1zWYzXukYGnLjbk3Qis+vju40cvOKFBjiYZqZPL9ls+e8maSCY3JE
i4t36MFWGP0E9secjBcZDLJmUGw1g76EnPGNEIDGCjfCR5KQrUJQqpCWqTpGt3tW
RTS4YP+2gutKTiVYogslMiGaPw3P2pNdhGZvHQ967/LVtxHcVqf1IgL7JvavDBSV
gw1DbTL/235mz/wnaS9lp2GNdoBE+C5R7zFE7lJtrVJ22/zN/PSrFw5r8r0ltD2V
8Qx6eP/pt6InGgx+DIqrjGouysub4+QtbUZ0jmVvvOcfmMfCRTtEoKfdBIOEuTni
ngz8pOpmS7HKUgYq2yUuy3+VZGs3Z/ZLtWTZaBBYVNLNRDsKjIzvVK5rcYPsUWPO
HRONQnOw+PZGvYu+NHTGWX2LCc1qa39y4RUkZfFdBBZ1nIamGIeg4X1IaL/ASd6B
1T4rDpixju462dcoceJCP33qTy1kThU4YIyzGknJd6VgRqy7VWzycyndNbsTr2gr
hP9xRXByOwyeahLr9LakkF+hqA2yNjXvm+AGUgDkjxPEan1UL48XeDojg2Qwd3wA
sDK1gwfgPBVDqByxuWvR/LoTbdpInmj0hUZLr8pTum9rVXhSpKYOuuxVxstJ6ld7
Ve3pXZJ1JHbuA8H9qZ6zexJlovC5m/NBbUseI/mRInSS/aX0aH7upEjsjXiYm+t+
VPf7tJroa0nI0AQtdxM0BL3HNeY29+gVloGMDOmP6In1olLg0XWDzqv4jNM7U7KK
fYd0t4/uwaH+N+EOQTm/Pl5uaK/9Y+Dn9W2D29H7/YWf3yyoLAXC8lAHDBGxDZH1
Y4qI9F+qJuT4W09igLLVM3zeCSRZU070F6NBBbjTnpFEkcEn0dMMuouRr6pdVcSd
6IV+v1Ggt+9qtszSpMK5vI1DRRNJ6JkGqQz9khSdJR1+GZjGN1Nh2n04fyyBDaZX
X5jwsjLhY2YLqvIn7u/ygkrFc8jUAlIg/12n/CrpYbh2/d3VvlDgAiwC+Fmd7/TA
wnHqX0tDgBKqfEjN/hDF4Jg5jlGvIlbsHo1g0tytwD5IQxgIqXFKlreYm06XWvsL
/NdwTzVuNy7XzNZ752RzxJFlxBBglDpxksrLikcI2NldoST+2wZcmu1RExBJ4idg
17N/FcSmsyOo6Wg8+VsP1FpEy9cjDaKaAHBO0eWbvbvjohAx4IY66JqOgLliKKn6
vmivSt2u+mpmGvf8XW4QnJd8mBy/s6jzE2gbJ17aPjNwwHg219pvQsHhIsWFUGeG
ko8TzHAnrQ2ArlBk777ytVvaKfw4g4Sc3put1YEu6dT3O9eF1XRnhmcnYNWc9+Qj
/SX9sVqIwYUmH2+2fXf4hst+P9Lqqcf6+kfW3W51r5C32FnaBD2EMy2TvPau2CBB
SUFlYlxrMoJEZbQ4JnfMVkCh0MJgUHYJkG9QKNdBkdoOI9q3roYeQOvFn4zwtIP/
NB4YiqNwzdYcnL64jKm6ZfBxaFp0PVVdqg6C+0fMWnsKmy8oachjS3jKcJXWhHv+
vBJPTlSuL4nzUJ84hLPL/hPnA9rsxYEM3ARbSDb5X+Ko+8vptMIUPHRbKkEdwDem
z/taNX4Wsc4RVto37c8Rl9Ns5NkfCi+izvqT4HyZcHEhmBMYUwAJyW82+opbApQb
oIbnKNUtQoMRIiKKWqN4dOP1nGQtY2dXLRHfqpbxtjFNTAaBdUl8bcLrnzByuf+F
UWNCSgNIAJdpwUQlRKuH1Jn6yDEKnro9m4TkHOc2eBe+GqnEIx82LoDL+bgajU+2
1VVPGTo2GU7ihPqj4Du3iBJ390/LpPs3JhWtrxxV5OtRQc30v2jZQ9bvaPtUnUqq
DoGkxzjimZW9OrK2sL7c+brsM7TNFF0Ad4YTs0SzJeHAGCCMTPN4hFD3cqCwvwkT
8d8/hdG1lEjoFCffQ32OPQCypCQqRIciX0lJbEExk/onNdvVI+Gb27nO6rD2NEvp
U+WJLRneHDDBSAwhdEYXDrvo8OmgfRGv4l3BV+96A3KsxjI8mP8G6jVZFWgqjhMH
2HGVXLdXqz8X6O/dJr5fhGP+I6XMRCvjeGvzXV5UMw2c+dTfmUy0qSet0FgwnZf6
SGQ4XAhLXvhYuW7lK/tS73WvzWliKROYdGDvb1dNmyRKXH/XOELsVZ2wYXU1R2RS
VoPD0eyqjxErnQw3VRH7swsA139DKXZmZIu5erH5fPWrtL/0UIcCw7thGzyumtab
F64l1SYNyGS1VtEh0fvOK5XMFoO2thmExsco2yLT8x+snPllw8GqpoWige5hAb0I
x6s/dJv7oJyhVUCxO/j0LJ+SthX3p8+2NCo7pm4su9XUt5FUcKBRObS/Q2JYtEJ8
FHK84yG1O7FkeNe1gcC7c2P5s1iaRGN2b3rOJZzvNUjPKDra/4IZcekDl2Q4bOW9
THqia2MbJJjvS562ZLaE3/RRv1Vkjy3fRZJcKL2p9IaYowj6Bb9Ls2Dw/gcYJj1Q
icLm+gpLGqV6ZJNIXJZzBU+RUydvaeHCDnxtlGpnwX3qBHjpk46uyX/D0aw/tprg
JFilOVAOnKfFYkaom6EFwWFnqJEMojB04LEXEkwrgrDIR3O0KALxNzK7uwxy3nfx
ho9bAhiRrhUcwdKSZoupsDjbmDrkz8BRSTBeaxNkKuVd7U94QbIkbrvZWypwOsLQ
1Dvvn8NTfXp6qj8AsbTmpDVQ+HxYJVPP7/rUvUUXhFMv5OWpSkfOakAIJKEuqbU+
oWvGGy+HMDpf3scJ5vzBa7Vf9/0bfhIJJv5lCcX/Oc1BtkMiQ/NIyt6OEl3mNtG4
8+GW7PhKr4FPWAigVYCdMIvXXCNSAJzoz62Mrktu7rIx5oNTpakavkIr2jskjELk
FGtYOf5vUNcnr4Nx9nzrX4PCrPQq+jjduT/UmVoVGTj0SsplJLDzAmbpRBdcSoKh
GsJJ3yVFgiKBJBQrL54mOr2u6U/1puAJrW9YYErfIpwO6VFUJPviyFX7JZXKAxUZ
RN5Ea0c34YN8ePpKFjvlnPZBSqeTqrWruCIDMPwQpjD8qTZd6x8mNs+ds4/blj4K
UbBqPzkG9DVTm/36gEyCQyrHTKN0e9b+ohWkqpVyLn646Utnlw4jhOCCLWhu5yTn
L/62X9oMG9BrJl3+gjCCayiWa+q033yA3EjVCzCkbM71ymIcTtOV+ZDkp9FW1qBs
yc85St3b3GvjmXh2Qt9AnkXF19NnVq0Cp5MB6StZcmwckmsddUcv81na8wsFMzjN
Vn1PkbJAUcH+sU/vTD8eUen32exTX8L3UumJP1SlOWUndRSSXf59xmsQmGt2ge6T
df8E1EKLz2OFkmWANtWIqHOAHqwtnI0ex1Mh/DF9JI2zxvoNVToyUxT1h8e1mvLr
3SOJyNIHaE5bAL3v8+HzeLwI1h5R+0G0YY24zU33FGWX4Dylrn2NsZaDJvSAkjW/
fZq6U6XdkPX5tRiyjj/C2bUnW2dasjiS0Cot4Elqo9pb1/zQ/mZ+2WmeTmJfmvYe
ojtG/9LMhCKxU+SJqgUUdsLoxOYt5OS/F0KFc6KYg+1e2XNS1OEqyPJZ5f3tGAzo
aYykgLiJciyP87n8ZeOSMx07n0DBuQAtcZ2AQqpsrzHWdAzqn7m846GTVZzTBV4q
aOESB7N8GFMAMW31klfXGWzMiyzj/zQlvvGcN1nokrzq0lj6YksrYotNvjjotLN6
Gi+/QGMJ6gMBYMUnceIGHh9ViidmxcBqeT5wFG2XTEmM4shLdu50YvyjbAp8NLCf
4YV1WYRw/LHMAqhFwe6hBNn1GoK3kBHgoKE1fXRAMusyORzXgYtItVO/HCiLD1dI
NWuzsu5MTfvSwQ6rU2WShAsOjJTlstz4oP/AHUTg8iBcnX0X47UfUSzuJgdkG5o/
+4SiOXhCU9sVqkIfE01u8fKo6k8t5ghUqGrbWY1ig750TtYihgU3q9Nlt04VFwQB
OsPBMHNiJmnzkYU3bdGFOLtyGAuP9NA+P821WqD855T85jzvjLlKJCGJDsWBpRyH
8eabvrdhEAMNt2Or2GwQrZkAK38vTYtk1Csw/Bx6A/sVvtQDmZLppdemMFhfyyEE
MIHzGBFl49qrP5axd1/NwEXzXhKan0dVHwrCXdQfeHGSVgeyIt6ATbhwz+bHk/ek
ELvaHZQmkIt6mQ28XzxlokKdIxaSUD+5PQAa/7GkkEqb3GYbVmfp5vYzouOxdRBw
UxfmKCteoE4SdqjMuxIkOGuhsSSrrrJEfehsolc+eMmdy6+mchVhOhjUDfZHDd6E
h1g5SknS4STrT2s0IOOjUJzN920hSdBwZgGAUnJsMtcZep15INhyBnGdbx2+VuQ9
pQl89ZXtlvqnvbPXYbO9aioen/VYg52zio4MKvKBl0+312+X0rWdf1dqH5YfYfi7
zKX+cKpCFQmz26wIWHIIYO0K7zbpB7+inUr9T3UzyBiW2ZG+5JCdFk1egpZ1uCsu
wHA9nS0bDRppuG121lyFWBLKT7eosNu3iOb03epcu5oEFiqGuK6iCppVxilTWpaS
VtCr6EMawLdhwWk3rizGXknYvnvU0p8YBEwPoqJm5vqsInpBz1Syr8elgO+nzXZe
1A+JDajimfAApmJCUUnVvufM6S3x0ynBDdqLuaRMobN7Y22P1yMH9opmTfuCsjPE
cmtXFa6q2dFdS0C64HwucFdhxLvoa/3rq4ldmjQjGUPQyabvhzmDnoMNUGrlxDWU
t91RFv/9I/OXfLssP21IZg3IvDQ1oY4ugiwcMKOSmc0KNoPyQHmMob4GVsaJ85Dr
HdhUDMX5KqDPuTAcdcuoDFLgFQqA+T61fAVPIH2IDxGtHYlABchIgwKHySW3K0li
iCku6/nB81I5vYVuk4vaOB2HTXSAlX7acewWPf3u17Cr9WIj9QR6HdUufC+5ypfE
T08VOH7REb5/WEV3dUsXm7g5voAyXsLzEYwLftg8BhU+jtlDZYt3l48MvIjOzlVQ
SOyQvEFQcxwinjcgA17yxR46J3Pfcm14xRUZ2jzSIoHnubN4gps9qRySsbZNlqeG
OLtlzPUEdlGtm60fK6lDaFK9ig5fzzJXRVRSa0Ler6jnwiqiFmAnpqGNh1VPvc1K
gI3ILG61cmpEEI2hgAKhSVJ0oVYQns0utunACNIzxNFL5hHCf2HHLsQoLTkuyO2Q
x48xmG0JEEE4ojpQ6dkzEYGVyBHEKrXs/HXI4uBtEENb5wxF7GoUKjW4aHnPE0LJ
j0XuYaRHy93h5Kd85F2G+Q3BCIFnPTtJhsR51e1Mr/FRwp9XRn0PedBOBXd0AW97
aYUH+rhc+tWDPKrn09l2D0f1ZGh/DS7hPmP6t6evlvP69kY4frIeUVgW1YstAC9U
wGEM09NNVfTZQmhcf3OC0WGQSM0GtDy2mpxK3MXc/Lm3sBO7ZZmouvv5SnjuYlW2
g+m2RzmDtA1A+NO+6ANpBW+RFPBSv8+xa+Zb2ob0seg7CH1bvscamYkn1giAESMc
BlQNu5IsjPR/KI9974qcNx8qUiOrd/59PyM0tMq07BpZ4+efSOlbu7c8sL0UPiz2
ZXVa93iXrWFd5tiZaDRcThkwbjywOTf00BIPvdR0s60XHSwfRSRNBrdIlIqzUa94
3u+QivYZITbJjrg3k6Qw8W8q9jB5xefMYM6YkW8sVapM033n69rw53a5qXGdnIbL
c4zrNv9RupddDRVhmQ4V+AkPIs9U4W8hzxbsGaLIQ1s43eE2m4LlUqTUFj6jGDAv
QJv0uivX3Q/yJZPB2L1hVnlYqpHvcxLZtRzJKz4GEDMPgOUYjEBlEAltl/VeYDPi
MemXysr0uSnjE/d9r6MYMxv2DVOMCxR/aIBsaw0y9Z9umnLatFBa3K88lfTcea9u
6m33K91fYVte399DZT/Brq+Tsv0Gcr+0uzOqzORGihk1Eb4CfahJvL97+fVSRiAg
sKx5OR03RKG/wuOORbaYoAawprwcWXmwq9flpEn7tz9RqM7KEzTezhVwWyAkovD7
HXC6YcWh6AiODfgiuW+XiDjV4/XEVS9wfQWdurlTjre3dP/fd3Gdymq/S1yk2QB4
zr0aAUJ6mDYZAI4AJnGe7SeSA9GYlT3B8pBcxTbiMCTkjOccHR6LkFpJT57Q0mhO
dV/VAzLaLyVlpp8lBkgGaciUtkFhkigbPCOQb7jUx1cLLUZb+HGaCu8Yf0u/gxVb
PSx05CbWTk0wJPCyW/dcaJNH+RlAEvM3ku8YQ9gRtq97poSxuTQpddUzb7EbkUIt
OLVY6kgwBGJHC6swJ/yjPBM4Oc5zvpogjaf6G69x+O5edPgfKP7rEsNhAUEEpHvU
XryF/xKAMsCIYNRqBFIeg5sVQRfrFKVXXj9i1GeByPNuQFN+1YdrjYJP2ZxOHGDs
ivILjipsoqfAK0GbGKqnOtjMzKhaEqQEqP8Nsx0GuQcre/EEIqh05eJY1GtwHCCF
ueqgfQnaQDwnbd5jRpkSZ16eOFI3LDfauaRaQeo17yflvl02Q+n0bE4vsCJj8c6a
rb/jMM3L8EgJDs0OXqU9+zxwCR8/iQM+1SQm28chlpmKwzFsx1enawGj48nOkT3Z
/udU3umxCDs0TBDhPOPfvAmr6pwwvnuPl3wyOKmaD/LnzyCRO25wg8gKJY9rpgVv
JXfsdHIgWCpo3eiN+BVa7XjJPhx82q0zCKN8ZrXJ0TXU/rum0Q7tsYTotArNXxy1
xTHyWFrLlL0TqKswdtsP94DLOv0WJ5fqyMY8LHjPbvFe7sbYWQskEY/wg6VMpy7O
Hqeo4NYOavDzTa0D1HH8GiJEb3wS1G7snhiT+mAdwaaIAfy5/9rFXFbvdtQFLvcg
Df2l1Zds9IH8/wTluLHrkHILz8vRvjbvC0bMX9ksgBmjkwux5L35AfvdOYf+xku9
TcUe8ORFgrLFEis6uvCxo/UVe4CswoGArECkOEwTljLKExjv6085d3adatzq+8KY
Bz6BfQ46ZWjJXMaTCYvCj0Gspe4WdmVBNEmyXQKwME33MwHhFLodUpbhbStu0KzQ
iB1PGThIeKwxIPMbSkyL8oX03D1eER2ME6aONWDqdJoOxkUz3dqa54RiRpA2caJY
LDXiAvrCwtFU9cVspPjTeCPCcQrkMhd8c/Gunf/AQyva+2fNo6MIh/Sb6X8HCJPg
hEdX6/dRXGLZhmuVwbD5pEJ/WurFa1ZqDVTqjSafTbstYC8I4z8kzmbo4rsSMPjp
MfuZ2Pft0vcll5XuDL3NT+sHUOARax4xzHxIUGhV66euzHI9BRz6NMR16wdx1fIl
6EXekxep+cS2tk7X2FIO8Vl54Kly7Wcm+xIE2i2IFwzXMzMHtiFFal/8XBDVu0BX
lhGtUnjsPCAEBpr7KlfcmJz+Fi6tOO0isdnM4md5ATh4lClyn+agyKkpD3c6rat4
MqUPVLavmzwpxoPahXt7N4n4QmrYH54oNaSGTrypILVAlTpma2AA39ykBnRFMMvQ
sv0/aCIYmB5SO4EIebjgXg1y72l0VVHg0KQs8xIr3EnZo93kU2vRWooqV/V/e17J
HoklJg8nCYZCIt4rJJBKfAKNXvV85FHitA1JsfM6JWZYUjFmJP/uDGsAoTij9g6w
umrSmYXQgrF+oin5Q+PwdED0vNdClHRgoQ88BMdTmnPZc+znAZ7i/JGbwNYWSa60
UqvRYrZch6QbfxtBevh1IwQFI5R79HcuCBNExdTT2eKd3eLcI5bqe7q6K3+vXSmi
FOBWNZtZYTQouotQ6pLUcNVoB8tG4iivUKREmZgypLZXcEUfN93oCPLgBJCaC0Uj
ZRM4rhRBBaoOUUDC9UfZsAF9FfZS5GK7Ry91JyduM2xUTj/aEd5JvcIGu3QC9lEz
sML1F3aVJVYFvwg+nbn22YUvZoFgoRno07VVgxC0uWvpZB+/b9Pbj516UK7NUT1K
59D3jyHG2pzKJC7Czle+Or8XL1Uh3RS+p+B3FiaWEi6gM+NtioDM/kgOejDh05Lx
N4bNZCVfAelwv4x8ZdQcPcr/y8IlWfziTdRF2zWJ+wVCsVYLGkUOMYLElxZU8nyY
Qf5EczRdWTUm0n7xJQVtnX41JaN7P/iJxr9az77cVlNxNvCrT97HmftYdxN214ul
R/WPUkfUGhv8dAfXA+Bjp8jYQgaK+gjnj+shzOwKpt41RwKQUDD79Iw0KvbYZy/n
zTL0moCDbq6z7rYeL6p3fhMd/YhZsNOeLRk0rXmACY1GA6Myp1TWkA9obQLxE/kg
lijq8MDt8JyG5q3/G2X6dj4nrJDBqoBk4KJKSpEapW3oY145szlTXUEK/Q2H4psp
BGzku9HvymYySbdc7QWb89ol05Cmfbi6uKhZhaKm2H+fBrLqjqRVqjzBevWtFsEk
08DwHuAQC0BV8ekdMe8VxEDHsi5cOJ474WNZF40rS1EKa/m3NRXiDqP64s68JIoJ
TWj8G+W3D6ijJ4gfV7Iaj5OAHgNPSQDXL0BVgZXmOW2zSZyT2sTXyKy2Nq6NFKEK
ALu/jZ8yDciKDl5FvS1IBO58lFyXF9vFRnmqL80fdBS2hGk1OtPBPQFkHKijMayf
ueyHQl00NwqLEzq3PVODuPWf5VT6nfChTHkvMWqO2x+ZYzg2+Gudn7RTW3Ti2G/G
qXOSD3gd0uizGa+/8kYCr87lXr6mI/vaJ/YbDURvSarIxSEH/geWYXIbU7+GpEVv
csaeCQEJvnYmxWIKutM/aMeHjtOzuONwYewuovmeJYUqvDEhL1bzw7z+oKtn9Rnv
v+/161YZ1ELzihuzGbVgFtssGe73OniNPE29J/T4USi88yAhQe9Y9qK5p6SLyY4i
m+Zm2oW6U+p/Q2F3x8Ftxko+eAWl3y7ew2QYYq98nf/oVhcwpLPbMj5gc6eoR1nY
XsJVRccI5JU5xBfcQlDNy4cgqoqRLWbl/DyOX3enKTkaZkh9fL1SA8BobLNq48W5
IwKlYPhe9C62LkRj0OcRI49O9TihN1LXHNx1D7UwxfDcEqVUL5y4zWsKYjzJX1rj
kYy4B3LBOxSzt9+C1wW+iNDVCrhoCTNxfrXJtsxpAa7EJJ9eejZHoIQzMFwYKjq3
nIxSzUwtJkcvTWb2UPMEfgYwjmYwGdmX/vpWL9ekJslelYwgbm4dMchKAUkZ4pa9
v/KHdL5jQEcWnOP5mwLkuw87lvFJFnORaRnHOHMbeB66oBjfxE/rogPcVxIV36LS
iLG0AXZy0pU2r2Hx+yCh8GUfZMyez0oySBt5CqFkUB2gb2VzidY8jA3or9UtSvAL
nD9GSdZq6RYr55pR6uMDaMWsbfeUbF93EG3qbAf2NUjBIRH6WA4EnQMfBJbSF8RL
X6IcMHtM73SiynxLk8YgldqgXl43esh5gmQttEUNzptJoNRTDaBalNk84Vnky1Xg
PavAbjNrYdiGI0NLJbMl9xxIjMz4m9T70S/fwXYFMzmq8EYbCFdpk1Xt9jw5gb2V
2x3YJxKmT7VYiu7L1rHT870jX83ihUixrpwPzkFrJcYOrKg1G23GTRNIbMT048Jl
0ywwMrRSNbKzQBocSgsI/mOiTg7kwDPL5zSUE+fwOh/o2J4qGJrEQpegoh5SSnxN
HqKvxBzYHyYkqbQjqK8QgwRuW2zhpEwGiJSDfGurlEDCvNDVbE5zkbQd55rQUEfp
1ZN9MmgbUkeD//VgXfQ+KgZMVBAaH69LBhzov79Kohhl2XeFUHH9LgZV2BNsR7jQ
BqxxSerQSq4akUtSy03qgDN5bJpqVgP/ifYdb0v5TIxnArMeWH9EvCUkXJRx1vSd
vdzfcQ/y+8uam5Z8XBAQS+N5aAtErz3SV5kKXzpi5TdExM8SYbMNsEqvXu9sglXM
SeCRxjAaaitMDGF7S+7YPwtinliFPgyLnPN+9pP4WwkO3IkMvpPBZuXbpAYlGm+w
FJbPyVRncugaeDIrTeZlvIH3Ddvx60TUWsh17xOpRW70HJwpSI08JCgjPnjMMwU3
JbaoRCpnWyyvibArKjdJfOSkEd4bShSqTifVSMkdjeJMcqaT47mng+fKWZbvuown
iTMXixxV7ECpH2qtHbQ0NvpMAGTCllGtynIkVPCOmTCEznb5kDpyQpMsZiJxsMAA
y+lvclIGYZ4stPRTjix5bot2czARxtPN/YIZ91pqVmosigXD27nIsKHMncUrhbnF
YLNyLGwfadwV/NqueeiOst7T+BxfcksRcLZZMqwG27eE5amksEgXTjnQiJJtm/oQ
ffEIYjqIpF+5SRwFIpk06g7u/LPn5l0F7LHFef/t+p1Qkx+IoX+Mgscq0bBBFFsE
tFF9wbvKtJZ4/1knLalVNWVbuJcieBs3K4E4wt0/ibflZhkjNKCnKB7V7nBDUE1J
uTLedYDcXGuo81zxAl1TmPCoa0l6dqSkbzf4rVyolKYoDFf4m/CBeCnaVWsJm3bk
kmantX7SwHrZ5xfZWoji7In5BzPm7N6V2+KaAUuZ5R+A6pATeKD+3XEJPjsl9i/r
QYecioL9aMxuv8hislFt+XFXdGCrgGnR3bLGT447tMf1vHY607yLHwocim205EoM
mGvANFNKFPELXkj7QSe0fLB3UiA/zMQ620aiT3oRgO+BsCKaFELTVGoqd7VdZfJ/
sknD3GDsojFoSBt84N7Y6UC874GwbDgx/qh7lgUpih5OSZw3VzGW33ybiLCnWYdS
Q97Ypg5vBsbP7VqwgMLwm9l5nBRJ3lx7LkBK23dciIDkYY6sn0KHFlPIPy5aX0Yb
f7NZYa5MD9dhIX0Ka3e64EivFKtw72EDTWrwu7zdOrDyNepifxdjsMmofKaT7QTX
Duq7jHkmw3kbJ5e3cOtsXd6viqbvWFh9gKkcb9GSkmrk9+cfqtn72QFFb63O0Abj
MH61JgntZqgy9LR/YAjXnIvJQUGmEQUnA/cGHjy9Bne7DS9gamxwLgJKEL2lVfo6
EWRJsQmjP3Ot/Hy6BIbgK79anT0b05WoFIZQtoA+liRjVV/znayT+f5F0jJFTkDr
uS/UEwiMf/zeeA5lNE7AW6YvxMAHeuyNMYrZ+eSnOUXJ2gkYNqMwGFJ1GTJDEgGL
ByXXiJ6wLlNkBwdQz5sUGjbZ2nBIHMfFeRUd6m4b9PztoDun4ths0NZA2TpoPHUX
sozP2GnQUsfNQ1SMlh/85yAueGJOiPYolRGw7sWgC1qN6u1qFVua7aYn7VXEhFef
y/+Bx+ufEG69yeqE/NrqM7KdnowIi+yT1Mmf9CdCGhIHKnN1AEQAs0sa7H0Ozvtv
zFf0hoWsMORh7W2MqXVDGUPft39JWuaDxXXsRP4dS71ejKJcenWoLMNSw823809c
GWjbHlhw8NfQbTLhuJ6rfn9xrd87umaMQM7gf6hK4AraCK1ivKfQ1zj5S6fFtkab
jdCqIUpogk5/PBBnALaAPgsB6V05MPNE1oQvE+ZhmSFjObTZKQBOUBCJoE1QjDp2
cWeiR+uZBH9DSnN183Is+QYUraR7LrPPTTTNr7uqibVYD/silfNCWbziXslDzd+j
l4QCyACTJe5kVtjGU1urLhBD3pxqoSex9sXJ7TG6w4CtBffPONeiNoO0kPmc1ccz
V9RqCYRy7hJJqcgAapr4qkny/+rNy+X6Z+O/jB4sq/OMk3TBG/3Yx+3ZuaadK+Zc
HRU9+Unu1UQXK2wyMAuNKwvnJgjSFHuymU3EL1gRBUeBqP5w+Qfn+DMISInmqizl
TC+wfZ0XaZa8JkUIbKWCLN586vPOdUONa0tDMtwexYUSBoAqXadXq3sRlfw6c+8V
2ALIhjBMSN/OrYEzC1ltoGIDZv8ychpS5QEEwPtJARdYymmYeHdjNUKzmnzkm0dG
100IeXPvqlQgyD9Qr0ec7tyPE1VIwP+YhWrc31jyzkSPz5BJMoUHC9D7k0t8KDfn
o70SmBJpy5NDa4DVa5O9CtymBdt3GfSiyPMEK2sOKlho0M9h11+XALIRRv24zTGw
AHShJpryR9NyR6CRLVhEVN1wxQXXhyFH5yviGptv1sj9o9NZoPMkQ+CNjEyafEgN
Sa3RRr8ntmeu4v+0LHv4vhbWjOKz3qd9YdRTyeoiC67C4V4Wk3L79IVtF68H5nPo
1LHPCTl/DDzNQRTev43yIYqIX752OwoaACE1BZdMOStIjEwqzwpCsRr2PwbIJ92I
U5cNL7genOsDxjJKXuhULSgGJhDf+xdFR/aDBq+JzmFn4KNROtNYyDS2vPILH3z1
zCjc+8V8Q7BDoGbARJCfhbJ52rXdE7wzhGFLwfmw0SHqWzWyrSO1bbMpfqsmjAEz
h/5QE76sg/eGxOtfadgZ+bxgLr4Bylsuoiv0HsxBlrsO34wYUwYG+KfHzNZtaXBf
hbqA+kF7yVy3qMK/e7JoduQ4oDb7SqIT5JBHGznJihsf3T1f6hXaJ704CAlqkdnr
xzsq2gBiS/KZkZG3scwNsHgGdCaX9HhXO2RJx3l9Pezd8Ch/pk+YDOvH+YySRyNq
pT3r71M6hMP68MShDv6/kPUO5k7Zi3GrUAh5pNr9QUFgjyTvP+DUXAHvc0oK0eS/
cTYoAIfSIInKnOzMlpSZNSvtW81P6zsNc9na8s2Mmf7O1b/4IbfPCuQBQZzd/deM
muG82IpjTyj4ah/+MyxsP1eVhr+38S6nK2y+o+aG8mqZ6Nl2+JJ/L1EhlTfWdq1S
iTf3yeGOF3KVgP/lYvLtpItU5JovVnhVDgHJqy2ev1CWFZzYn/59dsLS3cx6elgc
UG+sDkXPREyOULUHwEY44r7JvFnTSX+F7kX+33fGpbrPH2yOUYAQ4iA/KBGjNA3W
ok6S5D3EYHhOLV/MkShles5QL1CeipGgGgn8csH1MtIi3fKTf7rIfgh4jh3QgPWY
V+j/pfCfcd1NLKRulfwHmKbRZ/Hbeom4suo1EUHird55JaOATqaY1Q58GrUVP0bN
mMRv87VRGRjMLy7HsEjp5YETWwU9ho32psWogkXZnugsKCsSMIt5N1MgIDRl9y+x
FnxmRbASBzaP+L0GC/4O8rDOJ3MVy0nQzaSpUO1JWOkn7INhO3s8cm/9BZdKeYgt
nQ8n0dYLzBl3srOYrYQm94wicLLn/fw23lkilU3Q2btw/yO1qi9h+cE3ulTb4KbH
QE8+FJQnWHarjfpFjOQuReqXIhQaTl1ZbLTCcYFoVBCZoKpbpHNrDIItNUlJuJ1Q
TjoPLY4CdNbJh54tCDDzqBnlQnwAR1DIgKz3Oin3wz2QITYpCeniHzEjBdqtpmg5
8I4J/z4qfa95Bmvk4S1qhrSfVOKmwUnVpUcaVi6YF+Dpj7n3l1M0lFFMp11gKf1P
/Ti8GA943C9SWrIODeGuHa7gIADFrsTMqicpwWeUU8s2jMz6kOX8osBkXc8kFulo
4JmBB3l/+gsM9TmOqSiSv8djK8QgPSWKLLD8jnfqbY3yawQTQzhlzGRS2serjXnG
rl5yhgdyLbtXVRuKLM3he44zw85XqRIqlXSOQ39zorP/t84bm7T2j3N6L9HaZ5js
OKuYZ8iXH4oEKeBVrxjzXYY11+TuRtq/a5DpFM0PAlgNd8xuZUu0OgIAEZZ0d5ci
V0mhmDr44SA/vYeuNMl3KPE9vmfBzmIZpOgFKb/4/Gi3i0WtDJYigqvEtRuupGFt
oy+2AK35UdE7vTOVOcziTXwSXh3WE/UWbnBb/TMsgGrG6Q70aYAqUT0hZf9alYxM
Ipv5YidkORiyEqf8+2PcYAzghiprb8YuhvzuyGyE7XbX3nOQ1fRNBjHR+fUbW9/s
BUADXXNCJhIvVXF8+UC+DqxuFJzCoH1BSrzSU65jWUGKg0gmQnNWT0hBZrAADYHD
egVUMDg/6kCROGy95CXq5/CxF2J+imieNvjubszcJBI67Q7zGYXnNOpKT3DZAsOX
gRj/PQJLvJZydPQ+V9VaxnWbyVmHy+htL2vI3IYHMWGTwWVX/+Ph1L+vUa2Zo99G
zmikykA53hVQ9LgNFaB9be2wFoae3XRKvprHjWODz2AXloFAvtWd8ZcnHqPWkQNX
CVL06rY4QcQA13LNg0w7coo0GI5faRTEF2ZqgiFGMhzt3zjRa7yVceWYnqFRNW+J
QVja2opH+cc0U9jaQynN9yHrrAz8uYSdkxDJuuiSRwY3KFlIQ27DyuUEPHSw0qVS
F0IgiuA2zZqi0kM9o33/77xRQnVJf64vkB3QFuUKWkGZ2iuo7LfQAmcD0qatOa10
Iox8WXZjQgc+heM/K0kia9pAW5Ft4j+z9WfOEWOCxQimPI5+A4sity4hrsBK/Nyz
UkcmYTsm/Uzdv+far567LCEeRJKgLyvIxD5FGIksL41grOm/ksENSujB8k09lKNW
V2VfxAmcFtphxTc+ONcNq4e6+SRajxfgfWL6/ZpZ4P/ym6XMUzuUi2o3WmAeXZaT
EKQBUXjxTMS7uZeC1XxaYPzayx68woY8WYZzU7YqNi0NmQKDmDeu7f0rhuQI1LmC
rPcYfLtWiZSbG3VBz8+dIOH5WfAQg8K1p47wZSfmcsYdsCQVYwzg5STZt9JvI9Ac
f+T3vuof4abGF+a7bGuLzbbn7TRy78dadd1uQxCq/Y23uHeASsLYJA5rlIZ86Ciy
hOYi+vw/aOUcY5ncMPwB2ueSbx/ZsJa8MpWfImOzEdf4LZa9TTLNJO4dnUHZLDnG
ZjTnYQhnv1puwjg1nBdbUoauid2GD9mDtjMP/P5JXtcYVdC9GikTlwtP+l1k3Act
vnFizhAHt5z7u8oqFq/WE5Vadf9JrgViCUcmqs6CoBE8R5whEkjU9/y99C6cINXf
HaFtEvFsmvbZzgcnNJ+gVvITDt4fM8lvb0GOSISKQj/JChezhVz0q1MJsGgFSdaO
INFSDwkmiDgjPqEry3FHHC3C6N9ipJDcJd+WYCKQtQW9rqRIqMF7AWPLOAjN/vg1
CO1djPyH4mizmK+I//h++d4CHOc5iPLTkiE+RSSbb/1laBOwavjt6MxmMJmDEjqq
rxDVpV19J9t8VK8LBvgyAsUV+p2XguUaRUbE6P8+P4unv7MvHsiwo9uP/10YGnUn
5/+l33jKbwKxoJMTJkl3XyTOFLyuyEKRRYdf6SnHLfJFHA98cECh5VfgADwdoKMO
pDQiSaupSEHxf4lWXGD6+W/EGFCHUXneTSB/qnntBgri2xyVKZNeIm9OTVXXr9OC
GiUGfdLs+59u4SlP6rBCCax5TyyHzAWicjrdBxglywp2YmQ0juPnKgwypuS0goRz
mvj9JYhT0LKpHNunQK22OhOT4SZt6qun8Xjwve0N5HcucMnKntStDTTC5rNoJoAb
H01OER6ib7Cfn/i9HEy/nXhQ01Z114125iButeFNMF+OF7XEAowjwKwUfFuT+aVR
7Ff2fcbD0sT/IiheRcvaCaIv5RjJZp3+/AOdrVzH6hCIV2cZ+USKjoLFb/4EYFFp
M5IhmYaKQGzFcKckt3h2rJmM0p+5b61/xyVeMIMwbFGF0gCvBhdmQvU0IQ/sLqtX
oeb03qpCMrPw7FjkN45wUnlsW3VArNl4klZLRp8FogKcxgkWTRyDruVnuHJfp2y+
j8tm/nwY+/UU1bBssnrQK4UiNVpZlOuowGJULxs38ZOFocuOBOVP4NQCa/tUqFgw
3/ju30bIxn2WYT0RMB4Vho4N5LA4gYQZnDsbSnwQZevISDUR1flTBdu+v0we5ul/
P/VmpvlClxVrQeX1EEFzoKEcFcJ1Pw085t4E7MbyfzeiLS+i9QORegmHJkseDJEy
bHzzmqxpJmObCyugAPAEvu3D5Np2AnJyU3qCo6EeVqsjbzaQOTrZ9ysZ1Ng1ovqR
rXq2Mhnrl5vdm947z4NMzcyydRyXCEmQjsKn2SG/Bpxs/F6IUqWDo8CmDDs4JnRU
t5u9Q0hQkVormf1Z7ewq2OefMe5fxOazjtM6cnTGGVovkRrub9Q6JPYhILwa41Ss
OiSPjP7Gy6woy+sriVHw6lBM3zONerh6CEvOrBGb3snUBPlY1mh86Lrur2AT9bLE
2lBYnwCOVgbPHw/OJnV2bwPobmsA9rdTiQXekg3xFp2CNugCjjkgDDvyskf5HsNs
HJQUsPXPh0ckdrj/9+JSFPGHyurMEICgDne833lK8EGmAGBopluyb+jMDdHVunYR
CYtdmu4zxV/FMMaLDrUorB/PN2wVMxjzRBPEZw1tT3evBglAQb4SoDxNSvF68drQ
QeML+LVShWbieNW6M9NI+MRz9nU9PSNy+C25Yry8/I68wP7WlEN8hzv9F/Ss0VMh
kb/hS+Hrnjp26l4kHY+3kOaN3aesyUPcwiRY/wHAJRPE0wd3z3tA2SrtXHbW2BTp
tp9sdUKB2zHIecHXnC66nqyFK23hQakE8q162yhtC0WD37A091X7oIW81hD/KDhA
vUgOIqTGVDq03d8luMRCEovUtkIsJwevK6YY4QgWzKvpIBsNhP2Dt5OOzC00kJcs
Y0OELax0xuhba0QknApuL5W/viQyb2uCg4H5SEaFLDDz+64+8HGX6RShU40/aNiF
8Np/ItlU38xEUrtDnPQzzQ1luj1iTCzHldLqNTuO/eQ1H4cxK2q9G+Fu6vqQV379
+SUA1s7oRZWJAeEoQCjHhyBeVMLw2tZS6n0BHwuLrlTIttm6BgNkwMCLwxmVIEHD
qdaASeTYqultnQZk2o8obNa2rhyAJL5Li2ddOTqw/NXUaPnLkCF5ihQfVs+OXgTQ
6cRtqZZRvpIkUKO3QtzWYMz2BEUb1M1fyDHhGI5i+aFXFqf97nqA+6opzNElws5P
8Dn+CW7uA2VgK/JkkQTtxJ8/uh0HB/RNEu9KeVq7Sy5jMeBx74ZzmrDo8GwCIWQb
cI0TmrsxkJtQ3NAiGHUpHNklbSyUAVxmk4WEYlYZUOlJC0BOXLJQ/6tZMAB107l6
SP+sKd3Bi8PkujRfocYjc5NV/bbgkQiSfbb5bnc0FVH83Tcs7KnNkaiEZ3reJ1/H
wUM2IeUnqIwLcIsKYcnovgrar+QhKaiDau0BVcw9lChSVjVOwTEq2NTSrY8Ic0hf
/g0b98G0GAtgv/RHJ9rGF8tEzTEAM08JsizkVvcvgtW+pfB/kJbs9voXFAqXNnrD
sG6xF4NkTYub2qBPqfKGDWooe+BQlH+CZ3A/PjYHYBNL7oS91wNoRJCWf5H9XA+1
feqY9hzx57UcTlmtMT9XqnqZZ27UW4AGAu0tPFonZP1usf1mvPWfxUGbNona4CRh
AZ7xJa+xXAK3eCpCrlx3mGERPobDRlTlEEpLrep7dQxL9JxQULOmBu4PLDEFkFc1
DbwOUdGquUVRmOGCBloY8SiKG5rwUqGCiczj7bEEUySuDVtMbyDO5rLOWk4YwVP0
MJ4Na+8pXVnvY5g74NWSmff/TGco3IKYFH7MbMEFtxm90UnBNE6ELq1/RRU99yEW
7I820Ad5NZzlvrVjv7/QWvLx30LbvGepxwBtcWAWjy033hkxMCN1auNhqRhnT+so
Q9fpob2pY+m7HOiTl1u2XiF4qgctqRjEbMqsDz/ejWCXGtxnXtiGpRZpFS1bmnbr
X4+2f2qBRig6RTv9f0x1AHA3R8okacu1C0EgModr6GwWu+1G1w3kJnov2Unownbj
aQN4S6hyjz27DpX+Q4nwUNXd8V3RTs9wWqBDxA+F9us8rGOJm177oWKKcQK74rgg
/NfK5yCg4jZ9p9GVdYj0piNndcYk2MGLBB8iOU5uam8NEpq2d6TadFWeptr8kVnv
kKIs8uoiAlGYAlbyNRGjQhSCu2qwfdKaixTIqmXeQRzFbKa9G9ItA36/u61FK8yT
2xxtyHw4h78BmRads4xijlLTf/+/ejGF2xRalp3tjg6wPF7YbQHK9R/Lr6bDIpTA
CXUb0Vkbv5RL2Hyz3QoodzdRUh/JUZnMVF1ag6QSwNcY66tGF2gYxYludRpluTBy
f8M0pfldfArW4JbDBxRnPgdVRiXOKnfkdv0Ex1po3ng/TIN4p2xbV7NlmGt/L1yo
stjlGDTiOH6q7dL3yYIYO1aSOgbrApdAecKEm/JBXoaA1OLAE+VUWV9t0OHsJ3ON
N1Bob2c5UgdxbK/3ZhNug1tXlKP/OpJdImCd5lkhwx85Ewy5axvzQmX8WP+M3dw1
V7PyUMZgFjkEr9TiMGKK4JsFqNchxgh4tSz6VvY7hSaqaWHMDqFOqsVQ5VFBri9k
K+5nn7TcD085lTmydXAvTB97VX2yzGzNGisQfuBOn66gX8eQY08QYc65sPAkQDSA
1bjR0vS37wjzw+qhOH51HD0s9TUo9HVxVEpopFnAMn/9BodLYAZBsSNxDbEINLHa
k2xvGfqtTzsjz2ghHR61hWUfBRtfVE7bIfIQCu7Ysd51FUzosHFuxDLQof2rAxo/
RO4ejFGl/fjaH7jJqjI8G9lnC4/uKE6R+1Ymxl2aziqpUf0BOCN9KTYRn+sr8Hu/
gZ8TQJXt+hmJJ0+iFlKwTSyiiWweBZSRBWFXcLoMimAEiXNiUKaXyEz7EVyFaVLc
83jNi+XtBJCJMClY8/ouPFRrpqQIFkSejHHuakZ1xfMGv3B1usgqUsWCZzoET0Ig
8FidnpY6hGZtU4TOlo5jHEP2zMhuxarZFDmZFoJfg1eO1m2R3belrMwM+29hnE+t
2CNq8ho9VJomdwKbyx0ZA+OL3WFSjWTnVPjX6SUuh3Tj71n82NrDzlMq76/t2/Nq
Yfi5RJyyLKJlqvNiZo/W5uTJ+tfHYYZZCgmDxcFh/mKNlJ3fKrIeAyb3b0/AhLCJ
xPT/UzNq/zoRhU/NxqKyvryCS9hO2bnPunWk/V85NTEf9j3hIoCgQ5Kx6G1ETVM7
frxG7k7hWEBrARj+18Mcx1jyMJscG7UYiw7nyFVU6aiw0BGZofW6B8RkNdHDneAT
dPexdC6A4LBRmV1srzZ31vZ7Tn/ATf0LUBI9ONiELFsAu+nSmkKDYa3fcfYhpyia
Q3on9XrUSo49ziTNdGfcVacFgiw1CBqVUIC7ze8rcvkCIKVEHpgt32vfDRseZ94W
460GLCdlu8CuZWQ0QH2eC9VItxEO4q71x3A2C+dYTNKHpA0oEnRo6geit+4Nk8th
eh1AVoc969XLdp9+a5lQsS8yfyimvaNrMCttvfGfCBljRfZOvFychJItqp3O35oP
L1rD5KMiU3ngl7peJeWs6nEWEA4WYb2bDNlNBEKrBiKgSq1gDl3lXFnasjlKKWEU
fcNZ9kigLCLSjmRuDsByiQt+ze1QWojfaNKuTk3iNP4SUe+FdFMOPOgdZ/Xxopjf
hijHqvPU+FRPEf0sntaos+SOThDjyAn73NlRnlgt6KKfyEjwGMWv4LCfPreWSQvV
1GgtRSdLAAhcDM1sKk6k0OVwKAixsICa+XMEi69TOe8/rI1IBk0Cr+6TiqJT8RJY
upz9Xbc//uss1Hg7ZjfPM1JtKVFWaWYjivL1OmeUefgIaWbnhIU7t2IqknXh5iHU
47WrconEgQX2lwO4/CVQ60ZnEZx3KmklRLQvejpAcIyYI15ZRNwjcwWVZXRDulA0
JVfayFeCaoE7oarcRfE5jKHdnn3klW6IX6jhrMUk8ydsqeMAOBKACzMFZEnSCZCP
dRwB1iNILN/5mc+HTNfrLNdJGqGYVKeXNxNoDaXkNTZC9Ie86iUlQMXeSZVLLHfa
6oWG6RJhBAksQlc9EGdmxDYgW9f9IwFyvusnIsbpsVz60l6iBwxRq6eV0/uBQCYM
0zO3fBAdQeDQk4gSaXUlBVGYuodI/WmVVV0QGcmpLBqld/fuQMqqmT+u5oXnWUGn
WHXrAmrdcCKXw/OLQmd5aLSvXzHTgst8bMKOV+dVfWsQMyfl9/GfNk++jm1NRe1X
xA9PwYcSWlCAdes6X3P8zdWtDRU+LBhvKkusQmIyQLPFKhNkI499ERXU4i/VvM2F
z87Y2il9Tuc1sSJ5SCpezaXe7Ytd9ANEzzJrwd+X8M1fbTQhSBlQ8nPH9uRua7f/
VE2TWYWN42xCZ6YjU9mIj0/93uT5tm2Up3J+aQ9Vy0ER0cfiqP0flbh63gAGPLr6
T2WWNvSy6zifHa0coRuhRsvfhrvIPAc8cOd/4IBzi2MM1KfDV0dXWYkiGz+m4y1u
coHFaIXD2eTl7ytiMAxV8jnY0EFx5PG0Oz/rFdf2+ExSNKU5LnDgQk45LsEL7+mv
vD6LqcuBYSIB3+rzRHfSQ+7vEoIuyAH22dufFo88YhrxsjzyY5MqOzRO67YNAhry
Cq6hPqhcc9Ci8RP7Hl+bPK7WebwjB365JMCXTQ4bkWMprFr7bw0+8JZwNWD4JXkt
uKGFYUqxd7Ngx0BG8tbvpIQmbY9vkB72qtGb6RZfVGmuosZXyORrX5P2bNEe+Hm3
k8Ss0O6M0iPlRqBNTyNbFEC1HLnq/dAqfQaEgPv4++K7fwTyN0BFR6OhZWPQ2+g8
x2xmbng+Iz+MoiKq7HyjuqlGuHL+P1wNo0jRTYZNWvL0qbVfjR0Qn3yIhh6eLhUH
s+N4Fq0kPLxrextq63lTB+yXJp6lrykbxSfmmVfdHQcedzei36UF8TZEww4GDCdb
LVt0NDCqN5mzBkNzsCuAnwQFR6oV/1bwTpFu5aPydCMfCfVxaaonmDGg9aNys5r0
zWXoS7V7RU4ZtnPvmG/n9XbdmMaG6YlqaarX1ODmRtEkLTYfIpuaUOj8mksdqmDI
Vd0532YkzYORqPue7aASWNNlzOPaOrMtCTsrHT3b3CT2VAIzoWpxvMEGa2N6eZE7
zpKE66NzQ+BhIORsnxf8holUKnY8YToiUt0Pz92wVk1+7bTeehhLEXosgVaWv7+8
TklRCb6t4l/4MmR+/Fq6XrtcNQUMykdcFWR4mZQLqmE8fgZFL/rvswGuu2eyoN1A
SpNpsLOBSWctQvIULns1PjjIabSycsDY1AfvgUjIPzQ/lzC3IzPLW+Gde/iGlf6X
WAZVGceaeDhcX0K30AYRa8ZfyddoXF25y1AHkE1EF3G7TOei8PUkZ6sMQnO3j8hW
zxwn2g5kpuMPhWc3/SZUyXMfGHTKEoYa4kcpL1P0YFFZ6C/fXGazgQypX5dYWdie
FgBLosSK5uufbmlxbJldHmOCsrNUzEAws3mPppRT7hCBRPJRerJf/2rVOp4wnQlf
YbVl0gHQWen0sljz4Zzqixg4fXbfRs0OtLxq5pMqkqhgcyMV3G191YRXh4DiKHbU
8D1FvLcP3bsM5JLTcEDtync0QYtBRmYXGOuIqxPSZEuHlHSjVwaX3SpSDo9Tu1Vp
vd1UXYcRV1mpSlnCYGdofa0cO6bh0NzbvT2cPp3I3vhWhf8R1Bum03WB9v8bILS+
QuBREcqTquOURpMkRa3158cxc2u71BB8f+eef9PxVaVzdmMzKnzZOznPAqvJtIYS
Z0pO1knNBBCuUc0Mv9WdCCch/iXlCTgFzXagAtmrxcnXXf7wU0xtvGxtBBzmK/f4
LdzvPSrioRPEOgacDJBv1Je9zCF9A3QxO6ZcJk2lK3CKqlXQM8cKh6eydQUkc/w1
i6cEntgiWQXoI1Myy9QMQiRQ0z1kKijv46K8leuA43cpC9fQzwgS5sfHpA8G3AtV
d5lKgi39DkPmE9zVKata7QMeCHxnC7aQ9GzNybh+f/wKp4Mdku+/OUsn8BKgLOYO
nj8JSwd6Zt2/tfGXrTR7U+MNgdkd9J/+RdS/Pp1LHLaB6tSDwg2gdjQIW3NDwYk8
UmwWMJ2oY/UQ4hNIzzyqtEJ9CfqCi2fUAvf1Xi7a8zAIwHqpejZq2ejChGyfDJxo
haP6elJk1JzIKQFqKtXOlQ0ivBXge6Crl971jJPSlszNe+aw3rlcAp3rnqHZSYvA
R91dRDCKVux2PZdaORiJrO9CEcy8X3Hy+e6yM2KAE0QN2aJ3ePSaWU6MIjgwejov
z2ulXg9TaXwS2z1SxOXQtP3uZPxvAUAq19x0PW2qW8dUp4avVNF903gH7UnfrI1x
zVpXLtDMnHm+rq7c2bcQw4xvoH2iYSrW+rHeiAJdoLYCkpxNPZL+7QgKGH0Zd2L1
3kH31WpSoXm6zH22GLEZueKbROQ0dD9eD9oWpZkqwKNVBEjDBFbhSGJqmeMo9Q/I
tZP0iB0UHfbFHf/6xlO610XLvgZPigDgonuwWBhaAFjj8d1XBeIRzhdqQr+OaA3Y
H1Vy419Lz61GxtqRjDP9VfTdJpWbTzKuxwHFDUa7HbFUueFu+jmL8uTCNmGELp5g
yP+0yOUglob+jARxef0kkfeOv+HAvzMOuhI5QkrfPRiAIYS2x2AiM3notiS5fCMC
PXeP+8GazNNC56Vyf99AKqBxDkZlWPkgoswR+WqZuIvG/0DlmXjMr1vS/XdnSg44
b7OzeWkizZHpA6o6sTgHNPnfGCCk+c3Fj3cQZOIGQoi6G6NcciXdzt75MU4EW87h
pMHiVTVueKvX86OD+9RD0KTuqJiVZWAfCI0mKPy7K5Mj0BzJ0BFqKIxheTl2Zm0y
tiEJcZGbWbb8aqfS0Nwad3/ENxDmmtQ3iUm4PbTPJFxqaaJ1/GujpZQBXUVul7Mf
E7W7Cv526LR5xO4DJYHe0X2wp8SW21ZjZ/TYY3VZxgn41SQI0ia63+/OsOXFbC6z
XtxHJrc99nLJrnWlN8dLNSLbf3iD5UE7i4Amw1DbprK6x2oUua/hj43/Dk/UGA8t
AaCm+l5HoU4wUruAqyG76cJ1GwJEXGNtFo0Nb8ViTuTcNCJCrVF9MYVIsqC/4CTB
GKaVrfb3R7YevHWdGyHKN8yT0nF6LF4KhzbbzLSQf+qKZadNVT2WT1BKQSJ7Opfj
td+P+N8+jWtenHWJCJ5lBBsk/EEX2F7nZNWuZZ0ZAw+5hGdckHXJqb8CAeH42ys9
0eiUyXUsvQtMmMXq4AXZMvFcwv2sC+OhQFUmtRrHL4Thk3cMqr9ub5buHAOZtyLO
Rf2zPNTD6amcUq6lv6g3xsIVHlU8B+/0NBgxYfS26w3KFBKzuamKzeaRnG+Ms5UT
/kZoM5tLXDjFoNz89oV2GgxEl+8zbvJZ02wETEPZVAcBc5gq2f2xt2ffyV6Qm5X2
VnJKUBGwnqp/gsRGaL6jCZ4Yd2Ln97jZ52nIvAfvEvFd0VSR9oq/WdMwGPSZMAxB
qU6QxxEjo3REnaq2HBDkWWb1zTM7PS59MCPZHIFPtNJMlV16+tsh6q79rSpKV9X9
IdYz3g/WUqClbaW4XjSW46OKEQlGjzTgg7yCzwAPkefzNvZPy6vcTCwIIVO4kuCc
EClriw9OTEgd4oDJPQdEn5GEfu/Ar5jXAvTMRzuJRkLvBjCxIfS4gzLU9Yj88sYm
Pf3zIWkor0MdMivgTzFEio64p9Ys8ibiGvvbMEFDppxKTsrACnDmEQ/Vo+YPevCM
A95NugPeGJcbQ7/kWZF9i33qqAoHdYWBKG+/TeaBbmjGuaMWmrZpLbPDuP94xuPc
uROA+im5q6bi26+746j8k9rw8+meaiJaSsSwQmq0RupqzgYqAKgJrrhXqPM+lZqd
0+1HmYdeU/2Uqal639COD59i4KGUfoUzDvk/FcTVibWUWmfMmKR/4N0Msd9wPkdS
w2uDavM3n2UVC5jwEQc7ChWPfj7dvwSmi3X08RiK1ACCooZ41lsoAe/C2eE6eWf/
YO3GfCpJ3JXuv+QfnYbjV4s0ybCY0i2hvKe0GF0YTcB5xO6BM+Bb+RsIyqyeVhzA
aattmTFngSvSz8F2o0yvVsC1X8v2kF83H5R7UqY19Wk/gUbrDkMSQ9sY4n/9iPJW
t/OAsTrnKjTcvIGqiQ7Vxn5wxanuVQTrwzoj2GuParXjLeF4ysmnLEV1Z2bK2OZU
eEPC3OoD+joNL1BxcCMzA9Nu/7A1vBkoGYDVnlzxzv3V2wLRhiC8XRzh3GR6pskS
5g2PEnAt2STDDVRXRpoedPOraUmUv8WDCgzk/3vyKP+iC84M4G3V8mmxrv4UdqoU
w1Gm8OBYDzhyxwbsXM18nT6CsLwvKmqD3xHlJu+XRHiD1Q4OUeGWukgpVkypW1vr
wKmHLdZUo84t1Fbmb5THbxpP7oVJaz5w36ZvUBlGzyeANEoxt82Hjh/slpRSQsnx
pXg7qWVqgCTHnFx9MG3ne4RzpL7NlIr78uEmdqAYoaDtnt1GqaouH4H4/gUDOc+I
x/aQaJQYTTPsOWTtFz0ZS1/JUL8HNzuT8JngqWMbVzSzVNnhAF6wORFvMb7AVapN
Zsmv1uNAHkQzParo+sGrJSIllHd36A4NdR0OoM+tJqyLfKkmREZZ+VdsClkgWQvp
1FjyLRYsARdsEP3kQrRROnczZ1QYSQt6cgpFm7BASq96Agi84H3chMoP1U++bizg
u5S8WE7cugqOLIhoz4A3y14lWEgbjawkAz5ZBj9Mqur1GhNy9LBGXCO4QyqdN52r
zhpHv0tHNm5XwNx+wcr2ZLxRX8l9z/KFi4q4fmsJk3F0iOHOUDDrU2r0BWKN0JJG
KV69HKjJ0zamHwa+MWDiu1/XX33hDrHbr2lemKrYOAt4iNqheiYQrfxtCgHZXkZQ
Z43w7HeeHw23GRPQe9wg5pGNq2eN1bNuzylehIdDh4C+qETBXberO9JvfEM/INSf
Qwv87c2y/fZJUmfYBlHa9wzC51HT0/uGav1Km9/TpCw29ODkUPylrHYHzuURFJDP
85rKMDkpLTkneLUZqdMYnaE4DZn2OFuhL7f9WMyY9k3XCt8w3NtWB/lsr8lour5Y
3PzqQmX8FT2F/d3N4Y1o5+zDWnFG6cS3l2IQwFIEt7g7df2jeY8UuJaiDjYCTVEQ
EwWb+Ov2hjU8vH3mnVqPz3IknoSf9I+9BJIvYY7DJ/xlWcKoTcC3F+QMiCvE8Ys7
5dAn/vSzGKhjmR6JLZzpUzdYOIuDlpTPuQrVxw5gbOCzswtKhcY4wt9dLli7K+zB
ywBJCRQy7la2zIlU1wnOZs1Af/USK3OrlCwVaQfhSj4wZ05gFqYQXGJ+6m87fmFZ
Q4qSRvv2zfs2OQpL5c94So22zYufL/e0AcojISTqQk3mvaOyWaY93rf3IaaSzRHE
A1POO1U26DppP/uACRMz3KxJKF7kJKjjL7r4Niohoq7hoO2tQQ4d3nUuDS8f1ZYU
o8ISQ4c8KB/13a0xiLeB3sdWr+P0fnatvTjfOCqbLk+FuggcsEN8uQQCSJP+YNP8
p8GilkY4QK/Qfv4rEkS2RVkRZg0EUcdZRirRjpI8nuE2mDEBhxVofCVaspdhqMXs
ICvBwwxrdbg7HvyCEvmT6XFyoletHS5OR9Ye7spUFPym4I3jBObYBPWr+T14OYtl
Q+osyjrif/kdcjJ2x7O9k+FQVCyxANkzJlhg2tER/uaL9rZ1bLxw+KRIOWkKNA+T
YTcv9LcDRIJSx7k6585hOX52OfiD3Qk/cgeINf0q9+KsjgOvLc8ibZTc20Vs5Qz0
pEoHCRthUgZmoT7M5b7W2xyMcOJTOB8NrfP1NQ7PtBTCmtIVIQ8Ax+iOdkPU0BAF
MqNOqQDdELv7gwwHszPaVOgoh0KA3CkuunzjoEr37sANsLB6Z4LHdpXjcHJEVT7v
Kjfv+KHvYFlsRGnUdpWKYDkEuMEj+xHrtTzagtx7ycnasudci1rl/SBhjduF+L+7
ywgeE67hFGrSBE7QF+XYjAC5e/iz0e+EdDYOYM9/qZf7wN10n3cVSO1gbyRSoVBR
78fe3eKLt2WPRPP20lxzUbUc5FGMkD0RqxUewk+NsYR9vqz1mq1kL8No3PIrZJob
fiza4nNhXKGynLGSG2L0FF/awW8NEpCv7GmBirvxFxwhau5+ZOK7EU+qoLKhkJkn
lQk9dWQRyLKgKAO2qxfL83ErsDPtVt6p4QW64OhLqKCFUSb1Jcidd1qAI1ccqVp4
2mpViA47qlFn86J83qZJqLiKqALnUv7efsXgImY0+oR5U2O/lKDCN/XrXgffcVVC
2S4v8+qqDEEOE8yZTvuZtRKDxKnEMWw5BC3/SVDieAKtrhDd1yg0tjy26Stxpldw
Bk+2ES2hX5PiEIxt7DSQt9qWyQUWXZNFMCSyQS8Xbg9EpwFMdL8v50TABJxDxD1v
iIVQE2LD680j4LLA5nhd5EbqZaQOznBOe0FDjXTtwf+zeGpk28cJlwuzcxmJ2soQ
lgPXIOpGJuRqObIauwsXg3i9+L06Vjz9HLnnxMfDK4KFyoZOfIillXexMkeeRzTG
8Mh4rsJzHh1tVe9YX2kXzRYRpw7dwED4op/6QXF1xTTHL7AZWZH/oRH1+jOTNZQy
FiG6vUEYdlsqXLk8GumlpGaweDagSN3bl4BjuaNdAplizs6Yy34wipoBPcKeR9AZ
EWyvBsPZVeXw/QOyF/Txxo6eTzVbhkZgLnFoi15rGUgqtmG0/XGp3Ha704OHzJxe
k1IddgaYiQpV62mkeozdnJbcY6DxFPUy9fZuiiUdSEGU8PYx1Vj3wgsJw7DVGF2o
/dSAiRuxHU1mWlBOZMfqI1F8q0dzsEaVVwjt8OxbbIS/ZmhBigdSF+9nuKx7owYJ
2LG3BF2GauMvQVTh8NyMfSqKRygb7kGvM7Iq9m7GPwmbJrNxhn5KVCotY/PJ/9Rt
v4SzxV6GO0rErFh/+d97WJYuqQAbIj37q2l/jbewnKGAl4WCcZJ/ncEXaa7dEq7l
ZaRyFDIpJdxEpudqIR0JkHLESEYo7RmVjjUeswuwa6fFu58j3GM7JjCQSqMSTCnM
ldjUUe9qGb6lVoTvgk+yzABmRi1Nv6xxDjg9uJnBoAE2i0HP+wDqhmQ8c/NFE/g2
1DRHHC4qDPWFRsVbGDW5P29mrHDy6NyFKNk2QhTqu6C5PbiKXzu6PwmyyXwyTMUj
rd0VKl5pS1S+VHkkHVVfUdDjSgini5ArEDyDcEsUZ0zcLTaysOKr+ZTtPjBxy4Og
NgRI590rRIWAd/Ly1wOXdfpH6qN0VzoqOTK8eaiJK2vBHnDuc8fvZAjI4f4WnSL2
C0/Z/+dYCg9NVqstxLSJ/DYhppMM/gaZP7ptGa0IuSDingTkcp7XHGGHu8ASmoQG
SLzOoK3gEcN+6dfgsf6C5ycTLeX4Z40BZx0BrmY5EwwuCi8NkJS8jTmLhE/11jAw
JQmUousJ7kqkPgbmjum/qr3YsxtnUf+FKh6EndUWQ1FLEZVS3mNgUmYVR8Nh9Nqu
McBzsjxlY20BvWY2o7K6YnSQl5/R8bKw+t6hLtbcOTfxikMO3XMNXhiYPkqIcZve
FdIXR55ng05EmBqDP2S376VrE8j5WtDyekYYGR9WoZoo168B+sv1m0h3r5vigkjc
SVBOdIFdLTX0VKWArbtQKo4yex5gwE3GC3w4Uv/RHyBInhlfJWV6QFHUXcDfpewi
B7d1oOdSd/tGDflqL1J5HnjGTAjCjM7VNluKbKQm7mOCoCXPA8wYwRT5embm6/CI
1E9SU52VdGJoTeV0h93D5VFEgnoBZW4uI5kgpoOBVUreSxVwjT+I8XHQAWfN7Zj6
6+4C+l2i0Jk8F5ANJPUfKdzm57tzkp3BE3m0QjJitLl0RMg92HAsVhisx9YDtsmc
1i0p5wUefiXCEbzSR7uP9ahz8Ot0PhY3Yh+ong0+UFDUe2OojA9smmMbzrv25qG3
67OGf3Yb7AWr192kXiHQXkEUo/oAy47EHD1mxilg0P1hgWUUynSE/i0yYX/Oxyx2
pTaAMDfaT7jIqDnHRmpDdwKsVm5wx18At+tjQkoJ/rr5Qnou+PhAK0JmrNa1okci
Lx/8KIabpiZiw3xc/B9QgmV9h7acJ4jAuVIabTiGN4qL/JTIGujNaTXM1fk1NB/N
aZJPjf7aZlVad1/wVlsyH0vuPjC/ibBjzsKfVWwDRxUvqwS6M7rRtlspFWdOUW2k
JraZ6SAmv+FuJsDLMDRrV1SJHBy+RK1rey46NQGqOBjnhahO91k1CfciMxyKK2OW
ELYX6F6V9OEn7AQZSo49UPQ5Zrxo71BBOxpfwLwfvppPOjQdKVUwuYpYzIdOdmHP
851atSzz2Uy3MYmQ9n2XraVrvNY1h1VpKRBH9CaL7JMkJ7uWx0V4Bly4+Z8H16Tk
loToZH25KRwK8P5TalZQRaJhfuthRbUHazZGzc8LXkB0SKLS4PkRpIrA+rmmEpCh
ZcoYWlC0hRD7s1glvWWDl1I7Va1p62K1O/hiWQRrVpsHxkkTKLEKe2tmCol3e4p/
Aelyidje5gt8II3chKF30pch1KFzRMCyKVtznqlc6aC0vltAuxFCNGyhV+RfcGIw
UfGLTC8UWdMi3TsjjFFknp5vHmV2pw6650yGN4wU+M0izxe6LHnfPgUAH353lrUQ
4qrJ85JGu7BfbAoSqTeCF1XW/Y0JnUv/c7GqcqNyHFZi1tZzqKJkGxz93ykcD3FO
5WEKrVAvta5hbTZi3ayzei9Wg4HFWKWl/jDNPOHCuN+DVuRcrqFjNEGbhAKBbc+C
Br6Zltz9GOXtT1CjfEbbJYWXvGd1rtHj82iTCIPXt/Qiimo+zxVwsXZnX42Zs3/v
edeiclG13UfifnkG1ybOm4uv1o81jkLWD/O5ypVGugE/0wbmD4U+L0P43g8vnHMA
BHQ6DRkfLylCR0+fa1J3WYznm4jER8Vmye907l0ZyCOYmHLGyzYxZiGXxG+VLzQP
qjqQSMp7dOrS3vQ/BfekDRxIBDedRim11V7cvEJZ/GHIcPy7qqlZ4odYuZSPgPdI
9cHASelQnqjMVN1ewP3meerFyriBs/vLl7QH8xZsTYCZqCRLgOAWAo6G/6ESTt6B
0V7QmlP8YZniB4216hcGY8PW4My3PMA03OarMrpMNBDwKoToZZsLwr3RoG0+p0j4
2NyLrMd7u9xeRnA+LIt303HNhJHAMgumQOXNJO1LjXMIYzqDbDY6Gtat214Xug/T
Sl0N2LT7s4qXkOnYwF5sEcqTkTMbhG6QQL+c1BmnNScSZ4NfD2idkrGc7IuVyHLh
yTMFFm4Dk9u4fN0Lhl2YB0bOawUbId/ZbUFpIl50iU/9RH7YTr/nBg7VpzPLo8Gx
6A6jEza/tWOn5EAMme5eUg7h06D8XxWhWBKyHzyalAhpxSNNVLKKxIHAJydYaCvw
kSEExTCZTbNSUYldzxKEBGXR14VuoTiwCSOvpLOrbEzZ5UsOORCoqWjKsl+SZQWH
joLo+xVy9mcFBa0JgnZknRWz218Nrt4P0J4YrZd5fd5H4BDvj1zoQScjdkEsY+6w
yIW1p/GUVT/k+EVJe2FUfBxBYiiieqrllN3xQmD+ZHd467vx9+IasXs8sWKbSRVg
6q3q2ewHIH2lsOxJD7OnGODo115tH9LZU5LZ3IiDJu04lT915nqvSSC1N6g0KM4W
Pv4P+v4nYmrYSr8gNy6WICpqQL9+mHHlZxs4oX+E6jgO1mzU8kFKrcI8vgD3UY36
VLILrzK5J6Awg3uGjcpBjhm4HjfZlaWmmbFdzoHQYpi0kVzBl57VdoUxsKekdNlA
jj1+QsWMnoXWutweEot1/eiFIj3SUfk9FDpLuROJ6Qf/ch8G/N79QhsEps+0mEea
J4+lHYjPiOu9RWD+EzGu937zCp5cZTp/Eefj6DVtgyE6KaoJ0zhoemg/ewbk2MM0
T5ayF7wsXZCrjEeWdTnbuIcCncEfLIfLgRL1yhjwz4zov/L6KgrdAXtaghajcBBG
Oxl3/YjzCmHIsFzWGgOqWC3ciR3mzjmXYC+8tkpuwy6sH0daPA/YFnXd0QXTwiJo
85f6tFfSw8gucLMWOT/l7JRecfHY4LdI30z9AymGXkNMI9dYFPiAmVdfk2ZQb29U
P2CMxo9ZUm/ph8FpiYgsVRBgsXnmmC1+01OC5+CZ1+zEXxTZZ1wm63pxwUB4GS0o
nkVQBCXIbR8qjeBP+s8xL2eklfUXfwhPlVISzeCy4/IkJM/PmETkj4QIbd0tUx5d
TtIJaaXkXYgovFX4+4bQfBrrAxXWIaBzhfaS8ZcWq8WnOksdWvT4eVTPB7OSAbp2
c0X7TKpDYJJW6iaeqm4efbnoutbG+jGQTUIDLQ13v9/+O2StZKCZ17u3RMv/WvPO
cuEvNH9VnHobusbplU1/cuLlg75gCuAspl6thTqJSDGZL4CUEax+2Kc7yvImjz/3
sMvo1nLnabzpoZfH3nsTiXvAg5zJFGGqOAkY/Y/rFhwZ+DaoMhYwzlzeAMz6gV9x
/C/qB/0d1vAy1qNn9+8U6YSoJ/QMDBbDi9UG8BTKbbWMSPPtMOZ1/U2mgbJ8uG1Y
nEV5co+2j1hgEbqu0KpPWPzkNUiU4xdk7ApqIdkUTUsf+bDrUbL8yvuVUThhzbBj
KjZ/1b1W+83xXcUcHrI3vkgjJX8Gn8tTIlKcpjtBdBC/hqo9jq0GEh4TPNzyli/3
9wtLgl+n8UAHPJOAidOM1KnzaYTFsjaqlCTZSQT2GP3mUa2qw3jenJhLEjIizHnl
WR0RLJLLAS0Pf2hqHPo+pA5frfTz6AKAjBRa0HSGoFCkZ39LNQqSMmC8xMVtqwcN
TfOiMzs80Z5lRXxb3K+s9YtZCb8DHNjWSdrvdrjNjuE/3MGF7/S8y4Y77ujb24Rt
GjGLR4OKhryu8OdsqLwF/WdYls08/cTOZVMe4Hy1NflrlIPbonfxWhT8NaIA58AO
awZuB91lmenfvzRPCZtg40CUsTdpLoHcIPz+S11/Ru3mjXWeVnY/QwNDMDvcM4n5
iD79GQSzoxm27KjvH9784zHYAK/54ofLdYoAfr8EIpAYcuTxaeI6DkVvvIxmDizX
bWO94aeCasWVhkV1rxAz2jPySvKvFTSucrjDeysIeDSRrRbOAECM9iNPRlnBDbbl
han6vbR5loAzgNvcaJq391wv4vifyk0UVyr5diTTNk6ELjPFefcdNVZfq2+tHHQS
viQqjW8emsXnjT6VJYTVZSK2vHIHOi5r57xU3zpnBNTlR8ojp33HnGGIlLpIHQGj
D4fwChyUiRcnosSiENJR5SF36mHJdljGOeziUY4gTJRXt9AojUb1QuYGNNK7ov4A
NbqynaVIxnbPMf5H2LaAjoMJU4eNT0qJBss8E+WPuw9Sf5UInH3Xau08k6WWLl2s
hQxnD4VcLI7D8l1ki4cFyPENQH14YtAUiW/oLlfhgRwlxDYo2q0ZRUh9hw1TvNRa
8TyTKgCqMZZSWKXt2OMkLnfvO8ZRfG8QdwYhMVQgeRoJq26HnXhoFPbjqhnPgsvQ
MI/7HgEH72REldCALp0w2sJbN9lTnBboIanu+13dWAoUp1xvVGwFfVDkTpWSjipt
4p8IhEJm7fL/eYr5kelzyr04UU7hQ6Oz3mLDl2Yq5zt/TVQa47nTxO8Fl3VDeUI6
rxeqw8efCH8eJgr1W4+gQDMN2MBWZtcmB+H6z68OShdXIBNhQDqOll/oyQby0UTf
YKb1FGAVWgIWlz54m117i2e1fGo5M6gVV5BCuN7vOr1S7YZWLmUsdnK4WvF0JNrP
idCzTom9YCtLSqsMF1t2eWpe6BNp4q05QOr/5w5N3ZTqGXvSk3g+GJu7JVJTfsSs
xvNJ7YeQCej6wWNr3/WlDBD/mPSqewGEUR9gDyI+Sk1VjXbKSdN4BKdunTYJ5UVS
VU9E1TsdazpfrWPC4DHuDOmEkQ72M1i1eB4OBVt34pW8mb0t+s5AHn+9rMOSV/ZR
A3mFvaQt1WlIf3ODCtDbeX5Hm8Qm5gVpFFCcRpR5XQQX8w/Gt+lRYVeP5jfU+0FV
iNG2mbDIbx+hSlgkSQDznRuNOUojSbZJBOZhD2h7gXYQI2yr+yWXowp6ZsSQpPJ1
GJ9YqpGL1XknJzABCVJkPf/LqihRWVbblbaTuAI2bhWwl4Mq8/WrytcjdBzwQsQj
sJIkToIhJbV/A8V7NqTERCNRPLrklNxfS6tWtt2Yzlxx6mQDgqSGL9Xi7h/bsA8s
1e7ehFhHHqT4q6CbraHnDL653nNWAacoDzxlIhf+oD2EMJBnHcKCAuSkJAt/uXUB
HbOgEJVXTNs9mKByD5ZVq2O7CgLSc8sh2auaHOWp0UQ+k4Q7qL9Ub27KA0GjUn9e
KdfDdghxF1SEEiejuowh4g1vlvF1Ht2MdgdSDg7vzTJzzxvuefOFJ+9jsq36mk/L
n6/GKpBQILFT8dbhWaT3HLktIvRCg4QrTb+H9IkY6KI2OymMfzI2ESMAheIpyaa7
bhLgkVEkzgZ43btZFeBqLpORGH4YJt/y4/YmL48EGTRuADzNqe3E2hYGf9p7P3Ed
ympozdUShXnjHVmOGB5f0so6m7mdKilTYXfsmQBRMQ1zeL5d4kjW8eNct5Q6B/tf
F6a/F4L9XCE2oZYq2guz6UqkRxyWNuDdGC8bw3zcGJra0UNT3Zv0jxHvDGUyuQO3
2j3BJA5oZvqBcRKipT36hFeNNYQ2soqv1M1+R7QhBe/4267f4EKtSecrszW3DSMw
ytv1U1jEf069W5v60gfdKsKxvqgCDUhlD7VuKEZzPy10Z+eyf0xVOvPCcXMa0x0U
5EdqIpG5u5So721e3IQA4+MW4vQLXaZUL78dLv2RwVsrhJJwf9jws5zYl+P6VPjH
KtK0UX6Zp6Xv9uglvQQNpCQXQ5YVPX0k9HuSLUmtZoIcMQIsdZMAlOp0j5ZJrafs
mA+G61vcQFmEyM5XpV4MqkBAQyWudeXC09pbmWbXK59+v9Vy9ksBBKYCiotuvJI7
ycgZtRpZBCCql4e3i9YL6cfMgBF3coUe5nyhx21FZ1bmVVkFBJ5oGSLx/1kmdwbQ
mAwkysEt3/WOiIx2WVhF/8eXdzOmVetfHCE+umoTLudfWWSlaNLOBYIL4HCclyAe
ynpGMAfc5JhzTbi80fDIxZ9awhSyZ/J9mq0vHnTNUaSGJOHyJDSQMYbFJaegp7mB
kZPlEGfXNYXum8L1W314nIVLzj7I6cPTtyWoMRkFaOKXSn0IeBY546CDOqi71I9N
sXBHsDvs3S2tWlmjoAh0ayeG8SWkf4X6D0jEIU469QalWEbDD/RzmGU9WlVTU3jr
p6ZhMbuorRX6FfTPGM1PQSYt53KW/c7u+7orDU0w83Kgf7BZyNFVzqKjgpJbsynY
1Qsw+84rMUwvGXkSrEPF0oHFjO8egse118IpiBWmJ99uzGEArAQMjKjdZ+RgraI8
qFW6SwLOI9mmvOeV/DBsCFFL6xbIeZ5KjNkGoTx1mqws9kb7ljgkhYToCr2pWu5e
VTI0QYWXI41531TWYdustWao0/Msa687p7fxmjLNtSUc1eo5608MulEDSmq6qzJg
BoS4OwSNgKRqFKk37oQbbHGvhe7/1ynT4acCiiIfPwqDwPYDFa9Dnm4sA4rsxkh7
B0l6eNdLCxxphoG2qMaDcvKsbVN70ra6txXzFmDbTMx6SPVDVTbG/icbYUn8C2h3
PkGOysvHR3dPYc52eE6EsbTZetMJrFHz+vehWLq42jltFIllE4DBZ7YTf/GAzik8
lnzo8p3OWK5lsQbgvrZQG9XFwd61OjM0npJFZfdP9GpfEOvNqigeZUdgXk9uf+8s
EdwFroHlD0I3iAUD2r+HpmyvfUp/QMwbuUcj97mODqMO3vR2a6kJw/KrkRv2zRk/
bw1bzpbF2mamp6Z5937i52pZWCSGWhgx8Q9ZiINc2t1hZVXcncHC1gXSxk6jN7ef
HxtM5mojV5bYw4N6pAbgCF7WMjz9IcLQJsMQ+HI4TxxcVQvckapt1oR3Q5qTP8zk
Wrob7kAb45FbGhEUhPxxUtDz0KArBVRhht5amTHEwrxu2o6kg30AnrvxySoZlftO
HcD92Deg57MwTNZhLNKpvdYyHeKEFr50N2A1Y8ItCxgU7v6tPy2ckoTPe4UCidXC
pYRnLg9tL+4xq5TKmdQ/CSkdB7AZwOHEu9/it11Vba4n390JzQgUavE6l0CUQ9Q7
v9+YeO3TSZIvOHaJvXwx9B0JHXqXUfyXfU735jtCEOz+WR6okeXsXBUlX6zGqdjZ
fi3VegY4JK4XVf4ZjYqmd5I5Z5KJ+TbMgNMBLFzYtw6YVDA1MhOgkYJh+bZSsKfJ
b1gWXUtLp0wBmU2rX+8nnxV+BFHA2i42ltSj0mv6WwAtn7VtLPi1qt8RGTrgpwxf
1akUm6MiWiwxeqT2OkxJ8gIr3hvQ7IftMNuBX3HgdWNOGNkIjRD/hZTGZ3MS57TD
4p8ZQauHCFfFahZLlP3JYq8qpNhbIIMnbXeLYBYyKvbny3LDBvYspByg+GvUYUCx
rMF/xxiedOd7YcR0NiQhTXGgjdtmB31YXSScytY599GoKT9KJU+a3PQGHDxoGBtw
5DowB0StbN47F7h46NXw22AYu2xWcuCGIBXhKf5jd10qRnfLwSCV7o0s++nt4KNb
cIcWqw3/eTFRMAHlEMpcFrr9Du5p82qLzCVGLgQk5Y/161VkFfxXE+1rJoQ6d//y
mOwP/oMThijU4m81FCIlhexlRxP+JdRgiSKXvs6KyYPJkI3syFh8UyqR59lfXP34
Us5WNcUwFjY7DieQKToXcgONudW8pQw2/kb9UG7A/2RQqbkLv6h2Zk+cJvm+K/94
UjyX23l9aYdibvC+l+o5xn0/BvamgKCWUet0V5zUWNhaoZ2D4foewjzd23dkyjZF
CLoJyDBEkCmO7C+11Ik0Xn2gFynAHnMP8NH+MQ2BrioFdyqGkEoRPc1yidKPD19B
97tzS41cv1NIwvrnKwxVXKalkPfJercpPlpjgLaQ8jOYc8wFoOwMaPB+wVatTEJ5
HjMSvnErwoEM9/8VGHC5HweMQFvW2wSXt7V9vC2iPaAfK+3cbBxLGyl3P29ehNWI
lZe5xIOrwO2ONt7naHH6wXacTofS9rkxpKuSyEIIRx+cgDQAJdvij6PZry2V4G/9
KeVDYlnULr6bZCD5Nof4bowNoCrSIAfT3KT7+wQf9v98RDETSVgj+6c7dQXzl+HS
1uE7AeqW0l3GtRUgaFiA6Dq1OBshFoW/Lxv/xunM5h1pL0tTDtjS5YCIq7fR/dI6
xNBR2a6T9/kqU1jieuBWy/u6fhHodySzcsisAAt3+1Bgp2WyjCygY5ZIN+QuAMdW
UY/SKywHUlvKVQZ0AYFzcNdKqu/CF1SKp4jUlO/couPJlDCLQBiQkBvGfuQZvxim
vb11nEgJkiunUwWUzN40VFpIf/YvrrgZV7RCXwhfgtmRkCef+MMhjNEIycGUtcaX
JehHmld8w1W5/vMbuSGeXztO/CNtD0q/mXOpDowrPtfEw2RvC8T7V/YtlNVfM8Vu
MvzZeq/Q6sw9qhKPbTkoz5JO9Yy/03xtngvOJhpFeUc8Z3ISDrnwl1XPWSMkjDg3
FpTx/W3q7pZd7FP3/qSYTzgtrVzW4y4Lug1H/rjmn3YiG4yBblzi/T0adjxGBUvV
vKDtjzLa2Uz3LdOo7T1m2wsi9VYAxbZQdRMCKqn2ly6PU9AKZSuBQOc6C9JIUIvX
FCNWV6HBNgt7BZzgcElqOjm4rUsCRi7J/J29eMiR7Cf4RnQIRfjRzRRGGQZeKG8P
2TfZxmnkY6yRfMJC12b0ujrJxuAYfftxxjcVu/k6uxsuVoJZ5olshQvGopetY90Z
70y45K/ZW3+LxjD622oe+vwpd8B8/nLGG5M+r1anjly7+earBHdBP6AgpeDN13Jk
SGZfk9jb1Eb/LQ/GPNlndG9ymiZrV+3QOztEm3ufFWvWfQ802fXzgJHygQ21DYwg
UlDIYt8gYx5FldHOUEiGrpK2PwQCStlyws4CN2fh9i94JNll2cYMo7D3SCriLb7W
Adspz48ayErWtkN+Aei1r9lnypN+QgQCDpByG8vCylhM6g4tfchPmdjKNVvo4HnD
PLtH+g9R+JJAut3Q3PEfNRSW9npZQBq3C2lyahZVfkH4ALffpKh/QSYbRgFs54TO
8mCtbBWcZOfAzneiSutCQkhUAM4ETyJLcH1RFAJ/rlwPL7spWfKw7Qq1uiN+hOQ1
kjjVR+C1wF6quYTZTvLj6L5srI7+SENFA4p2hHJ+werGu8IQ0jK/V3HOCnr0wxkt
6h3TWcRZ3J+yqhZzOuT0cEUFWZHH8SqlIUJpi1hLeXPz/Te8Zay3V5GRo1L8MkCC
BFbVEju9sYjSquXIg7SgdrdI8kRmxPsJ9VyvUNadOSE+Aaj0EsUCKkzzWJjNyeH0
O74cIXk6sNVIV04Lzy/n36J1dgq5PJJ5sgyj1kBBgf6aQ+ebjS9J40vojOZ0y449
aWUz8eBy7rgOAofFcstACczE60vKsRXWcDk8RuNC024iB4NFBduX9mtJ8QCavc/Y
fDk7tI6o9c/cbw6aSjmDvrhNs/XlfxwmwYEPcTcpBzxr3UyL3yEG0H3uFRkn+QjA
hLwnpyngNI04sudgoph6TkYiPBaKWQNOK0YNTe+62icdTaie3uJ9A6X/du20pHC6
c9tJlpoQNJsOfZyz/wH/TWDJ9A9rxu8BWQx3jUKkquoa3K4d84z9qHKRY2RKJG9a
hU1dufxmVxAhcy6xhqI1/cP9do4E3FzD+z7RCXFPuVWrRT+TkVhPcw2TWa4ilz2/
u9Ius4fwbpnFKh+5heehqJhpu70S0AxLBC1Vgumxs6Vq44WBpGpHLBH+YhmFSreh
JZr9UEKui81f7WABfcaDBmRaCyPKKeCm+RiwukI5Jgog+InMtVjYox+J8xGvH1AQ
gUyszVtF1EtNR50qC4WfdPtrlGnwYUbG8OGhfEu4OPcr1qWUXsEiyOZtblv2MxHj
jWLNIto45PrW2Q0lrqfit9B/j5sVkRsjBGv5hbz+vvybZpQ7oPlLJ2cUtrQvNfON
GTL9Q4WFrRsIPfWQo0+8V6MFmUGqG6GimRTavWw4ProEF41PJ7tIN06etrlg25LE
2NgVHbezM2a3DzzBq9XP0OICptkwn8N/cfQ+gTNeTbPcDwXo3AdqnPaUUTWKdXEQ
PoLh+6HbK/7y8i+SeRcwyVYj+y1raCNojjsUkd3DzWI78MbYGHN/rZfYucW6W+aY
XvhR/CSOY5PujHyiVK6rehkiu6/9LLz5+ilbLn0dji3pRNBoOIf+t8eHXaD6i/iR
xx06Ew0wVP53kZ+/d85fT+Nl5Co2DlV+LzmVtLNGdbRRse+RkDCenMK9Lyg5hDJM
hMyeNOI0NoLnbzRIPK/deUwIikhYjvpmiQ5uCbM6zIw5xryO3WNCJhCPzxlpHu4+
oPRqzhP1UIzWmojxZuVW5pe9iF4VTr5/V275eUD4wmq4//c33ucbVWqFHp1yokXG
1rGpcpgMl6h+nklIdzuF45CxuW8FesQuXJp0MuIWFNxiNPz/nRDipGGVS5W6uYn9
n/9Hgm4fPXHd/FBGEXt0kr6XK1WhKeuQeNaFX3MleTZ6QPa4xCi4ORBDaB0xl64T
8Un+ZQq3JiaVrrMKl3Gen8ArltCUGV22z3otmC8lII8wfeoK0VUDqbQlj4SUo1FG
K0qUOU8VkrUwRoKrXU30x2zfUFeNFy8i3KZtboycY1n266NJ50ELe96s++vlBEGS
xLnvmBLDeKy+nuKX3zAvSKdHZIRSHzlImNqW7+7uChtcnJRQ4D/HicQ0PibOhBn4
AwNg485am6sJ/JbxkVovdX+l5735rVUj1xidG5Kc0yWFV6s3igBDayDj+Pr9Zesa
fAlozZiVTXNTbsR+KDT20xo+h8GEBaKcs9viSXi8iiBSw70e38YgJFnko9/Akwy4
BfUbP8Vy/UNh9XA7GcHT+7XMiF3y0tk0p17xyqaREbIEavNqVHQgXufXChR1xchP
qmmpen7S3v3klxiGCjXF4LM3dzEYH9ootRidu/j7DX9xoHKCGcDw/LfwJ2sXHC52
q/iSOQGF/4meiAtHW+FsoXCmvU9+sadKejp5jXzlX3SJCb0TCXAZi2Bz6pU2piBh
US+B7Gz9PMgfnscKIpvQU13ruJcnNi57nNXACtnkmMjTrD/xcWpsfXPZW2ckX5FK
ajTm7YihEJjDuQHarlzYhqwwmnWlBzn+xGUv0FhbfVtc/K7bU+vaXELvQkT/sKlG
iEqIBltFVmHPjeiuBs++szfUL//yROOpoFFYI54aOg1H7f6TQr/jS50b/i1WVA0l
W2AoLu1/TmsXNLYPaBghYWVSBwfabnvFjkAcDZa1pw6pSaUWhv3lepYpi5NkZCJA
0aJ8LOAWomRvbtTj9lCVwsx0wS87s+cHqnnKDuWOXl32dC5Qi8KBy112taHkdCF5
eeWj8OTCa6yWkL5UK6cdRMSk2CTlTb3cL90FTvfcn8vN/iLCrU9MXpSHGI+DZ8Fg
pRjtXNQAt5VF9S8zHmK3xPc871qySIGPKyCjesOq2tICPxb127FKAvxDORn7WdOc
F3e+pLT7D1cT7lLeMEvUlY95NOBYaPh9sf3dJmUiq7rRLOd9lquGrv9uhaVmGNCu
CYUCl2XvLIjavbjPaXzArPcZf3CkgCXJxMR49JL2NOc5B8q0Lo4db70lKg7yrC0h
MEGxf6boxozzPlcjK0rM+1c81fkWbO3Qe3If7OypoywO6PLg8rcBgv94zlkAW8fM
iFw5/PHgvpOA0iRB36ITwdz6IvlfUTNHhr1W+fvMtubnxB9FwvzRPHIop0DLozBR
TzrYFYc9h+rAez4EiPsmnx6OkyNEKC6jpgWH9kGN8AaL4EjicW+npoqyHiE0Q1lY
vWNxFfgCLoMaJj8k5gEMK7boJNyoIfrTfe8P6Ww/OQckWgMhxb2G+aW/egJWpj5w
1pjKyT9th3gXrgtaEcsLxsizH7/rmbRa4XOTdrK36nI9R68bjY2ust7VooXKuJGP
yavbyOg8s68QOO/7TT1OM1oGfgJl/XOO8lmdmlPQvslYbz99ASD0lI7ChN7hDL38
SQELBAFWs3owrU7tSsxSJ7mbRvy0Uu4Eddk8wtS6RQcQrrzShq6H2qsZPVa63XcL
t+pJzagl8ZwDZRfPjv2XCYKAl8ri3tcvlHrBRHODZMOcej4Q33Xu6xNo5vpYlIBw
GmGZ2I3eEW8e2zbZhavduPshdjPwdN7kzXmzfMElT7qPriTf6tLXjDxj1BpMJwiX
cchDQnUVkDLGLBmOAlhrAoIBxUKP/OalQz8+J9Y5cggn6ftemxKmmmpqtxpiiL2g
Ak1yXTvpjFehPDdp8k8L3qzCDsvnjjhHyiKMzPMH3mfkiiBRoeSShHg6el3pBMPL
R8O/E+HMEmh453P7uI2ih+xuNToH6wRWN8OgyvGHWWhtJRdbKZ9HR/IanJfIQUF2
peZPYE9MNEmDPmHLXJV5lRXmC4/kAKwoAE7jbKIu6P3gaqudRwSTy0xZ1ozF0S1t
aTqsrZq/z+88N6Do0DQm9MH1FOTIuH1K0xzmQZkUluGvpPmtHAnmm+IE3d13VAaf
96GH4O8JOeLj30DZJu37SdjA1N3A2fR0x1BYMMuMimIV5kndcpHby/8SX8nPRFYO
zVmm37guPT7fudc14AudKTq/1ACYHSUvRsDio/IWfSaMRY9RwLjLYtfsuuerqW2O
eEXBrNt/IDhL30ZK0zz3AoFzUFSrooNRLxHwtCO/9MBFNwv64H609TC40Llugp/B
gnRP9VwmZA+Rh5dnu+Kn6c0wC2BhCDW1e2Nh3bTNc6gVTKML+JUFfvQK3BOrIvwm
6J4pI7xRSNDrpKi9cvbxPQdbYsXqbR0RPLGjxBezCduWR3tg23EpM2nyIGGU6vJT
ibrrq+1rZ2rm7GUDjN0yJO5fNcd2ZcIXMcuGb+BjcPmtjSKeCIgl5JGr7S3lV/G6
QiJzWc77pzds/UljVXqERiNV6C8aTEGQPcXUXGt9Cox0eUmQas9+dfrz7b8HYWTd
av5EEeIa+INE1qGdq1VsOFB4hyvdel/y3wNgtCs18KXsrhNBhltrumQdyl/sp768
IsImdkfqRs8Ld2oGstNgkFxRDSSrkJAyUHyWD8DIQn95FFWV8PeGvUd1LjgoJJ3L
OFJ3FBH8IdXYlGDJPP8TGVhg/HQ9XDK8+nx+uPe6IyANd2sYVmisVvlbfI6E/GXP
0dbZeTr0OC4sSQ1WhkOSe6tZcIzaLDQsgR5f32GZunw74jdDyxpC5iVWPYt3QyiX
5vzKwKf8BFHjo+eHQ08v9Y2q2Fs0//JyVM3DJnSnS11ve1dB30GiGckk5hYk6+gK
Z5vmpLYMVKVixlt15LL6jRDumsg2/8+j27fv0BIqUoPKVakY/DlpfHtQoy4PBx74
2fuTxUusiK8ZRB0gDm91feu6wgIweFy9V/Z0ID5voKWKHMgn2Rk1R4oCuUKkumlt
hb6fkBKIViEKSwJvwS8nYHXKktz+60WYv5ZP12zTD2onAzXokgDPy+pPTSeU5Wcx
U1gqHXbX9lnwjF8S0SAhX/KxpAaFjkW2wpGbHH9LJVsbTpR5vBVg4BdK3Em+Dawy
Z5+uxmqKTAyFUm2VgAjNzVn8K1tIS+GORwq6ZSgIaNkupKmukOtnysgyWdFajYrd
3IK8gQrQwod5Q/XVkEMtg4Mr7lEj9YZUQxRETAxJYskoKx8ysXuoedy2nOTcWVv4
BKnLYo7L8nntFizc7n1NKStgAN8NCh8wI7YHpfsL1YED8Ps0zbOY6iMM8R6MsNiC
VHbMDWWIuXGfbVorIrvSVruhR4Ks23YNbTtkgvwd9YJ2Qk1IjUnDLYss0kNg8b9i
2n6zyJzN3J80iGWG9/bFllY4GZaKYULLhblsl4WNnP7jsXc3mD6x3AVmJFOirkdl
aNmRGJifh9IAsiyOblfC5viXLBAd7JmRzuNdx5VypKBV2U2rh9JcIpRfYxOcJc6g
3Tl4V0mvQDs6ynF9QbA1NRm6m7RL/3v0HjAzD1fSO/rzrVdtfW+2FgNGWb1DgFVS
DGStc9jUwSDUCV+xhWEYcEeFu/drlYRPju4aF+SraRN+MZ8tJht8YghAtADb7HdH
wANMvEVaVaETKTK+eN/NC7qy8N0i/K+phgDovKnABkO0x707uSz/ywveD2C+hVCc
ZVujzSsBVySS2MoLFjkPpHwoyWYPcmlwNK8w97FcIisxTaRxMkr5pcjb27eXAXdu
JuKBNXpV/vJ8OVTdxCSib3sIeHwDNHMJFhPccWh2LEq9LEeHW3b+IEB0pNxnFsli
Y6COPeX8iswF6UKk5HCZxcgYLxXunAnA0X1EHk4ttXCe5S/P95r4EXgHhnRkmR5x
VDPaaiC+SXv8SDm43zUjSb3rW7K5fxmeVkmvDUSoR6xdTu7vTvF+WT6me1RrECWv
TrkPNs/rinS6W1SzaZiHx7jRiWGq6FUyNx+n39Lmb3H1kOTnzNx61DMzr+39B+RZ
9NS84fwO1Fwu8N7QOn9r0qOOEmcGStP0iDekfx1IarP0yIgfT9I1tUHKLkvvy0ef
UHrX7Qf5kh8yLAmcYW9qyhISufDKwa06mm0LdUZtmsicX9D1UAQxbKfI57Sgx/fI
DLCEl6o9quL1LG0gf3hiU8UIFq4h+h4s+LTZaGD/yZeIlJx6nSmBCM0B/i6gh6kC
sdFbWQ3IXapf9zXPUB480y6CPdq7nwzer27bsXM/aGuYCUHvi+FJchWvnEYEgWZZ
GrBHZoYuUZooerHjPRrDKhHN4MFnQ7aWSh/vQ3yuQOwUyMQ23I4BVDZ6SFsobSN+
gP3RyCWGe3cxEaOFjAlX6T1LfygGKjBg/0RSswlbV5YzpRQYbF4FRvSH2pzr8jzh
59gCw28p+mdWPF/o4APNwv1fmuMggBzTrJsAJO8Dp0Kz+md0ktL4ethyd3gjCZsN
3k/E+AGq2oeWYeZ50nWpHR1H5O1TmlCvRpJRnwZR7z/8Q1dAhqPvVq/m6BNNHRPB
7MeHXbZMoizMac9kqsAtfzIhyIYKegSvqjwGGLipsjeHos6PdgRkPqKLmH8Yp18K
nyj0dxUYdfi4LRo9QGZ5HDPd8iDFrpG/Ysa0oPMM2QJzmzYi4Lax5ytssm9XusgA
kD0aKP2kYu+BgT/PDwQNXtTSrYjcBT6WBJPCyOIQMO2u/Dh4zv+4FgIlNwIMuf+W
JI7+5TBLZi063wdJlQYaTkHL8rA2y4OX965ezDmFsH4ZdJb6ZCsLPuPJeeTQfI83
H3XOhILqSq1rwELJ5yIHQfN7l0lsBJK83OZdr163Z8eUXb//+IRzXkw+3MvNWki+
K58TYeYXPy1IUm4/QAK1cgmRuwuJ3Vf6aU5saevdj1uB0AiNd1ZcDLYIbQDxZjvN
DKwAuf2WY2oLzaUGt47jcSFQJlpgA6n1GQG8NhwA7xFCcot3VXOHlk45+titCWAo
xFpGJO8CJdsTbc5bjh0926ql1I17KOegm3MoAYebv+qpY0K45+/PZ2h8qOJtQNKs
ZZfpjlFg+0cqxbanCJguE8YOYNBjTyZIxi80Kfrk4wKxCZhw4117+fybbcHM2Lci
4a74DS+33ZGQ3R8ojT1Y6L5+lf4vt4jB9+lXze+HMrCo8arQ7GVYT4V0blauQowX
2wN9cqpeF9LuFZjPd5TsO24IlZfOkIz0RwsiXXvjCArDuA2V+GyMlmj0a9ZJT/KB
Q4dNoc1RX7VWSviBxvfNXMb0sKO56n55A8bs+yH5nAsBlHTSnt/kLlDOuHpvxb2p
fuYv+fC3M9iJmCACaMU01HA10AQ0MTEka+zNmsA3JIVgTRIcWa9h0FLd2NHT1QxH
O17187Tmspz5hJAfh5OOeHWfGbYlyg/Lz7Q/8y0gZ6WyZykJAwgPD5v9IvYYLVV3
AXWxv7xq/gvyRjsuXcNFyYGWcXDa2NdJYlZqvKLa3/KzTTEJZGZiuYTqSZN9052B
XKOyPtbw54Zl55o3bS0veRgkqYsFp6aBxcnJhp/c358yoWXK1MZCo6BlmYk2Zx8f
A4+YmLX++jadBeJ0VZZel6HWBcNAE1lgXU2gYcVtFtrMEDDWG7YUqj3z5NnuRaQf
fLMTWflhr5LRjqjoMueHYQ0T8uiW2dPUsT0QuNmfIEebII5+s60thC9o+8G2+hSt
plD7mAdpjONy6xXi9QqxA6QtdT6KT99xuh9mW7FB2Vp1J5UpqBw7WloVbEAE5Zld
TWmF8Zs5jLV9R1ukb8qt7NE/oyVxe76tOuOCw0OyXUycUvHSbzkgck3U2q2v08M3
ZLw9CaPeX64ZZjEdXiul8fnEY0FoVhWtLSFAiStd7Uh46rcaAta588vITnH8hjtF
Zts+Cp/RnPMpxD/pEGx5m0CTHeUyK87QImyFVYxGoobW/tRqfptegovhtLNMBm4t
JePgvBSbuEZr5P7EaBeiktJrNNY2DE6LVhN9Cy4J1KUpboeDg4V8wDrEy8eCjn6u
t1qs6PK90OMglaMF/+k9kHUgelwyBTUe0aIpB/ypklAs5yAnRFvhe7UJViXcl0m/
RsRT/8aD3cjUORCPmp0gD7RoUIPzdoh0hkzEP/Vi6lcxLsS91BbMm2EVln/YgROK
J/jQVUWHVwaLCJ4mGLu9zcOUtw6jvXU9ujZ90XV5cL6gmpvZUo//+8W1F6Upvz0N
BFb+kN29OL22LKXwSdnTDakj9S0Utf2RYd33jj8XGq8PqquiHWkZUFNeVQUum+yk
c4fM2UHLO+2TABuws7FlLzYV0UqXUWhPkd1wer6q22iTXgtgiqS12J6rkkxErbeH
ByzjZDLGEmAqwhRuHmiRvdGkmLk/lA/hdXG7VlIiTT3Z9DUmmt5MPq4LIPTDMdCQ
aXbRpzrb0fYgBabDz3zEFRuVbHoOpOf9yw1iZLurny09mdMlYnN0zD/J+BV4vuHJ
RrL78mYwWf0UBKey/moNKf9ROSG9JxnuV8bfe0nPkQrbZBXmiV8izl1fWbXjQmr5
ZM5QVPmIOStq9Ogrs9dedJlVNeBqxXjrjbx0S9b4vXYN5U5FSjpdHu7XrnGas9fh
1NBpL4xVoIPBG+sWzuYk4kTlP27AseHQg/g5RSK2/pz7QJBH+ohxW5gJAOqWfLaY
hp6F9bZ3AAfw7u/Fv7XlGM5S50fKtC7VVZMQCDDCzD2r9fMQZI50CtlOIujbhSDQ
T/BVzj7M7+OhY0irKdCFjuUtFuHEcAo2zh0OX1dMMz6yxpyEJ+Icg0Hi74tv4QD4
OqDU+FPoTvDeo22bJaXxy+qm53Iyh/v1NA1/tiX9KrcKkbRutW2/S0y3/JmYg22I
NfsIKC9LFGyFTXRe8hPWjI/ORVMjlp+ZKYYSHpz2gNsmR0NPdWLO/gLm8/ago0dt
t73HDxP1sEb3ZORp8G3msn9rVgC4ezBHQOy9OfsPyyKFrUKQeh9nsENXChnC+uJK
sYpY6UGcB8g5NXlvdXY92i0M8cDl2nm6Ifw8ntimS/REHExIXH6CVfxPMHgVNlNd
z6539X8SSiKj83Ip1HmfJX9GWlDL8eKS8OKySsR7QDzDRzv2fKUd7MSrG9X6TnQp
sHn98YJ1LelPRTT3MnRZsGZP8/Mj9eIhUZETzoHHp29zoryIAW18/8Xnw3Xpizou
zPA9MRcovHqqCWO9slrDZcNl5RLeZYaS+KKxMZRl6ieyGvbMkoV/wpMON5j/pdLI
N/4hBG02Z+F3mwjuc/Rg9TY0x2DrlR2FqGShNphXBTHEw3Vrk2zp6Vqzt2dTbzCc
UylBDj6SyfG9WiPRrdfeBf+P/wn1HZMaKVTbvtXByvNrCz6L82/8tX2wnk2xy+la
yfsg6wJcNgcmQVjkzzIRjoquZun2zSG02Y2jBxqFteG3lL+rmV0n9rGH+1bQJ2Gq
Ilsp/QfWK9OTaguOkM5q/jKQAhDLIMdLOPucW4G2XOrZe9F0wACcVQtvE5Hmp4um
kgzdi2q4zbN8DVUaLmM11TyliJ2zFVBy4teJRl21B+Tq5CMZauo9eeO3X/+32OyK
NSYgnqrT1eR4RMW27cSnjS366eWwRyjSY3JfLqreVyc9Bmt/h5DGQdl8aAAD4Ed3
tWz/eS1cAhzWh32XQoh2L1OWQSQAOZO96XUfmmhzx+nvSMa6flTca1+ShGiYVXAg
1D2usZnhrtGvqwQyG6BcEixm6c1cr9gYrJVs/ioqOWOdufiBJ0EFXO9QxpJ5lDEE
426HDMEbT98EBT0ZGcpzNanpxsxCwD7OBQvoxofgixSKyu4wrYOaGZqjxigYa2Mf
bLH0Y/sSHKYBY5g0Ldi1Z8EMCzCgM9mFPJ5qLNw9SbLJzDi4knU7dXiy7UyL90ve
S8X8CIC9D5jbjEz6tkgGjdDxp50zAho2rPpjAEptf5L4HP7BvY4bPPHj8mRmy05+
kmiT4Kc+4Rg1oqgoN4Up9JFSx2NU6G69jY55TMkbTb0vVUnsNeRdzR72HD87yREo
rtZVz4wUvHeBb/PZxZwKN1oiUlh7UBC4bnLd0w6FJh676W98WHWFo6JLQsgJvHNU
6D6G+peGuZowaZ6wQbi1IYX00DxOWTLkNRVJ6b5LoPPAhjdh0CdiSoHSSGXKolnI
Lp/ix4IaMytyAqykLfJv+n79iSgPAFFoYQii8uT0D/f6Z7EEm1ez/5OmfWOh9mSJ
xzUiFYAuqNdh8qvtskEZqPzVeU6tYLpsbWL2bWh/QosED72XxLc+wNbT/X2Fosgl
m16E+NOBazfNuk3HtAaKtdQ/bbq1LqK3CrU/+gm+FUCe2T0WnUksDQC9i6u6UDWe
M3/5mprWKJyud+JMIOXMFQMJRQXjNUhJEYInFUMUw71SI7qHqVHjCmlJ1tiJV7Dk
XouDKCRlzU2u3GhSQdACYQwhCSfYDSjzUe/Y5SG8Qh9fg1h8GXupkeHPKFJ0NF4Q
b5G8UROkhH9N8eLiyDPGgrWdpv0wKEu07V35GF91lyXi+JkFUYUkdo21FFbSee7b
h6Y1wcCPE/W7fKXKNWmF0SYZ+KcqonZl5NZXhtNDRbS2fqtpL2i40pdLlOROniGd
heEJrAaUj14eRSfTOfjl1YYM3cVopUEWhevPexO14TS1XDSAViJ7GCiGAzojo2wy
3cHYPT1aLmge+4+3Darb2ei91ZcSXJjAdDvXuYEi9V8R1zRY1ATBz46odk4SjWQ7
tVcuzZl8R+hecWCTR7sf45o/ylG3zSjkPvV+HSVwGnnx4iiDMncDmbBvgL0lIe6z
V3/gnrlILJQ04Mne791+EEhWYYxhkM3WgrQup1Rhf7fik7nOeQHkAYwIKK9KlHqR
vocp0Br1COvPbCw267EeszmjUO3OIYhIv+ghi6e7NKIKHSBbpaIOOQyW/5Op3egf
g3sh44fFfbU8oY7xX04tmfI7kn/tIRlfPutP5j4bJkKjNjsFdMgAFlwhHUn2GXGN
GSsXjGIGzikU1hu2UF8qI9PRXBS3C6oqJTFiKtleUR5ZftErm8dzDLMaVMW5A/jh
3mVUd55sopSEY9PET6j9KYKPQczqww0Ik7Y1jIVn/Yw9w5HRT9W2xHfR/UcMm6mv
oC/6nr0p37htLcayaRAHz+kWO4ejFB0Vb5rNedH80QFDnRrBEkhkgnFRne9U3W6t
Yc30/+J/cIOjPUsQ2hNZwXtbK8ra9PPgZVqt+1JOYyCs2TLB32JfjjyLCJsQniLi
Ltwl1/O2sqJJezeJxOjZE07IIUeZn/YoS/DLh/2w5c/SpiL3p7xQ3fDIDgQKl6rN
5ZyRdQHglfvscMSiaecnECi7QuL3H38QhPMeS8MIoUGS4bjHuwMlmBhPND2acbOV
GHMAGe8JfTQRtVKJ10yorunq3geGbxDHx2kbQbNggAYFtCE9liTuVAGegZ9UK1iZ
LNaRx4nI4N+mufPrkGCF+lMsMjCgsTWqWtxjwUggO94AR9YtYfaohlFgMjSCZFJG
nkczmdp9x8UWfRsSoXZyQUcS0QWhKzIjHdVLU1lhO277aexGeEf+eOXbAS1U+Nw4
yhgbpet3j7RE7n6i+suGjX6GdryPiGtmU7tJ/jiBqFM1aKTDy8bp4ANhFF9o3c40
BrN0Uc1JdrV1yZuh4/+2UM6KkfrVzWpAxrG4BJkiT+L3jKSIjtO5OoXB8DMcWbC8
O7wGbm4aWQ8AVAemRTMHZSpKfZMuV2NZR2nXk5O/VByCCvktAL+tT8C+doSMmP4J
DaFxsoEm2+WhVzDErQa6UhlSp0gSNVCn39t/J+422gbHGcDzKejpt9w48mJNp68C
eDi6plNJm532h2eSuI/1Tmb8lwojGztz/wCZmGXrhqnDX44i3biNpecIwS13thGi
mY/RG+yTPQkU2Pudblz9UvKDH5TnAPuCbxoceAC9Y6+QjkB4HOZvpFF67yUEK/ng
Z/CH5Ca0LcFDolK27xLB8hcgD2wrF2V1BXtkP1Iq4nYyrYgpA6s3ESLDJrVnNxNV
ahawffuNg5q3n5mpBVU2dGRBNvRXI2ZyEvTeT5KDvEJJXk/9BMSr+ordd8Jcg0Zb
EzDmr9r/G0lEkOKbLC7DRZ+AFAFhixainQ25WXEpdKfB9fwdo0CVE6UfUNkF32RC
GAZG2fMnu2CJPCTAANqxTF482n/vGPdUCXvX7UPpQlNfEk40sOtC4NP7tS71a0UP
MZ4QbZkhIsLgo6iBqzR28XzUotZa5OBoPFiEGKksW+FCsTqHVBkfMjMzxx7aAuBe
mz7n1ZQ9XuVc9+KtXo60MnUKkmrS0SnOQIQ6bg17k8mLShCYuXWR1uu5RBBEx8vP
4lfBSb5+0bvMpz+WmVeewMmcy3IOOCMui1RLk0TLB92CbCTKzA16hRXUwQLcrVfD
YwJX406EorRfwsZDoFRq54zOFn2Oa++E4N9XC7X3cf1pmiFHWr4ZinEtcmBTRaia
NaNP8kR0qHhXxnFFhRL0gPSk0Vk6uMd0HPEnSbVr27wKV4bFPpzkANlXwa+k51nx
Ivm7+/laOJKM8K/7HPEGJdgk0l8GegUS1wPdIZ1kO/10dgKdYZHBr7ghBBZxzrCg
LDCVi1ELozM6zuMjj1u1+3o5I150Iu+lqngBB6PtNkUmWf5PJ9+RjYtA3jjdIkV8
frzzDgCeDBPWXX+xkKZtDjNB1eYDr1p070OWCE2O98Jey7Kubp61ggwXQwqEWcQr
2wkNknRlfQzNO/Cg+1oB1Lcn62F0sgzUn6pzGUiyBgxH9yrii+hhVzgVGfpfBIDC
sch/z6dqYhLVCCU4aBTFZAXxpbGwBjAwK+qCZqiF5NPoWKdtqS3JxMWR0gYmjdHI
5T/nUQiH/h1dBfQ7BM1gtSBURwYfpym6q4LMEg1n6Ul3uJBnuXMAgZi580FJyqX9
kQjJNsWChoxtCHl1FeWeYh+09YesGWrPvdNGZfLWAd92zODl5Tvi2pVzwXPpBYNf
jHauAFdCgTQJepmGJnLZvSeOSZnT9UwWifEip+Ph2uE7O7nWdZ8Nn4/vlAW6QEsH
0xSgLGqyxWMopDOBuuCZzs7+W9SC+g2a6UXMEQ6X+1lQ6b8C+7ndbrg5X1MMmgh2
OKWhy90u3JG6VQVX4CWy/SogMMOmaBoypI+VkYfnjraKT3CWYaaAw1Z2vJ5jtpNt
66w8wLNce7ZhAZGQ3H5CA0pJlhpcq+FSAe660+HAaQXs54uPrmry0O/8i4ZncN/+
VHrVE33GSAOfrHjkGzJtmJo04hImAAVHBKK2/BotR2VkKYj2L/mjARAbwty5aV2t
H6Jg8G2XEYB8S5ZsmB6E8INu8vWZu29/PUch836tccsVfJA4o5lQe3sB4Tgh9/m0
Bq/05HI7xaa5fJUFe3BodH1Sb7qVpSYFA2lTH09nOCph3z+EfweBStlNDxjNDOXK
ntUiAUXJETNa3xAhExfXIg8YcWcf4mBNtwgNBCaFQtinvg7ZjKAifi2A5oVqVkDp
eKjJFl/RrElXMxf2Eaptyj7sAe9GoT7+E/fiuizZYW5JyEsHR5VYJuJ9Msiq43xY
gavNmbnxxB0ukxndc07VoyS6DwVkwAN6QW/gPVGoA88sSP5qcAsJkshLeWT1K2oy
StdBVeeAgOHXmn8JJI5eeX6WsVgBB7XyBGAtlH8XQ7BfmHBbe5UfUgxIUVLFmGA5
aWnfHhPUwEkZQ9RcMeDlM3pX89pVI3TN+O3HcRc9PFNl4E9Sgp1T6HXP8VbRd/Rx
NlPGKUunozZSRPXZ3/GD1+B0tEtCbMQCJaDdEQA/Q9OWI58W83/soVvT5DHS7BDR
kPpp9D8eN2uenTeEbWwVhJIVt9anlWs81X0Nc1J/40VJ7okCNmm/kE4bCg+27h1k
qLMruOGIhfXWUGMQVMfUdvuTMrNa5Y6I92xL1OUGJ0uv8ZJvzf/8LoRBx3cgmbhI
768dZTF18gkp06+6WCX4f0mWRrOqtcrM/bOg7KnP5NCJSarAwzLBF2Iqbc573xxZ
Y3LIgh5Ioz2IMJuohKawTZk4OVLacrKwqZwUXxBjtOYH3fjrohwujjQ7InAgTNeM
Nq3CqaJvNALuNsdGlct6JFSvC5shb2wnQV68MooSOVznIeJtUg9KqYoKHFRT1e2k
zM4PJZmkAhSIZuprf1pqiAb8mKFhWVYG+DWkOW/zmdaXSrjEOlZ0HbKk0YrRY2W/
6ywyCYjMSRVXR+tyA1xZFqmgh6QXFE6LEP85C6zoEAm0yyW6GNGHrEgaYQGD+T9N
UTfNU9UiqTp9/mF17h88PoqvNBcxTToscxLrGy7c+MHyPz+v6qH9imYt/MERTDws
B0ScXFjTcQ/7igIRBNZJ6RCoW24rlInLujHbDaOM65B2k4YM+3mPirLvnlbqmh9N
d79pBm9eqkrkwo+Zq2DvFfM5PXxOcQm9oQAqLGxQWa3u6Jl70FMd4WcJsI8kpEnO
RtRF9MgHJpFRaQ+zxX04Gi0G+LlpqULzGKzxV2oLEVDMvCI0iCrVmb2DqHy4LBPp
d5nbnDrZQW3zWf1aYjdIsFTdbVwAnkqdlUaZ1NMA5V3EpZncZko77HpEL1dBdjgE
Xely8qfkd//JTFo46NFSp/2TqrCsZlsqljLsQWq0Ebs+rMGoO2z/xU9LAkLYf+L3
+6mahtHQf7S51jhzPyZKk6davlHihKm1rVEzpB/yVIr2XVyngiFnMXM2EmhrcW+U
fi67qoLkHYtj1DrJ+VRJDXzFQx2HLbVesg3nwu1BszxodMt7JdOCF+lDn1/EMiEd
9Wz7rCUDDNOtjyhR2Q+ivezrU43kqtXnwxowyAk2lzxo/3R8hJE1x3EcrCkfz6+H
fv/vb+mf4oaIiw451cOErycBsJgQr549fTTthRsEmGAVb75YitRpIKEVyBKMwUXu
teG6dV+A0GDijaPBQ68/A2nsTW9QUNTckbi/8BDlc5G01JyfkwNefuLeuDf6+MLy
kg1YNbNQqjxpP0Q1jBs/n7FggxLgRSXoCdNVm3Ar0rev1UaskCEl47/ZGztCRtcO
mhABL9AiLMFyWl0WaAclAPDBzKqpUC7Uj63EM/VeBf5psDAA2c/A69474JKqsdfo
nGJlqyBvPa797X5rU/9ccdX+7O1fYlhi8GI+ZyQqNpayC9JXbyU1wEfEk2ivKwSB
yLwPxXk9szWGRfV5kC3GPf1p7fKiov0CXqeZ6KcUtF1jR8jaYsMfyIoj0Dbds/ro
0RZrcdYPnDFGMwfDqXHCIFYJkY4SCPyh9Ns8tb6WrPzJIoX75dlJPE3y9P8BqUJN
GpnhsVKBqPEfwZAT1s77AmUm/cMg5Gcptc11pIhaIMt90InuXvdZo66Ye6Dyd/Xa
OV3v9/Zojnp+Hu7gs2QNdfRJ6fmOROaa4Qfzx9uZcAksXGXqswXR5P7YVQkG/sgQ
iMUWeW/kKwjDg3D8/9OugJWFqxxiDZA/kD5WRxOnzHxNUPQdfFD2RwIYMoQH4cMF
YHmlORLY336k6CYlvBgi/QTBsBttOtRc+LAWJS3FQuCbFmUzSXNQpy8h82Mj+If1
tmzA/dYMZ3CxDGD8SSmTFhw7VX4CXGmW9UxDuSgAmWTete//kcG4iZpyKphd9VYy
AY82+znn6S4k2BFwDTdKncBemKWrtEssAELZ1+H2gFB8NDYryY9WUqzamBIAZsIB
7gMJFdODIbpDLis1arKg6bVppq6F0jtEKMzLQK0olRYValNLYUigHg7styD3sec+
QnjHcUfF7wMy7IkaZiFXRVCz0UWgYfG9L3rNFRRCOL9Ch3z68JWBHf+YLJ2pAUdE
7eOB38MNQgtl4bBqwI3uc7891V6yZKbaZGLrNiT85KmELEO5frWTPN0KnHh8lWMH
LlgyF3U4MQn+DQ8C1gj8sg50IR8aypYqcV7M27Oy3l4E8qty/wHhls3yP3ENYVkv
mxD45xT3Lx+vqq44UkLbnwJ8QS2nvC8khGq0HD9bsXeCYScaOZ+A4rDYd71Yf5y7
7Wo0Rtd4yGQ6ueYVMkiyAgjQZ9c2jvLT5ozhnZxePsfe+8wD5UMX3BQwuhz1opgB
XYcab5/pWJUutCJWMsxGkOHgUj48gZPTvcpm3ekI9Z/kKJL8mL14SjkI4RE5KuR7
IxZukIuEsM2xBVnAezoJmIJAiOJ/QDZ4hjU2sdb2UE/jTQM67srjkHxcdd1tyktI
w0aR4lYM24w1T+kE9mygowIxCi/LgrGlI8qEzJft1Z32dzwGTtARNMDJCApYWIjK
mAg9bvd519GCUcgEmynKlNC95gRGchpSKN5lZA9G95sZJKyGuRmIzEKkJjjsgA9P
DCL8vtx12WxoU6l0YH9cGciYpQwAGjW91AuulLQ5iC5/YhWA8Zo9u3PEH0IdzHGr
1yocBEgnEMxw6KCsa+fTgaiEqNGIaVnl+kN712hOsmsM7iQOPvbQRKzPRlqi8HGd
RDxqScdjD+heW9KN/0VNVGMraNao8bOF8rjMnn1SJbR4zTjLgK36uNrqU8akDKZg
6x4OBJasFaUofv//SlHW143da9yfcgYatZDVeP5jUoeBXQN4tRfbFAsx6IGNbkoy
OE9dVS+ZVQWdoP+VWCuTq2Thf2/E4WBYvJnZbNrFsdpNjgrv2Y3NIVRqp7xS2j+0
Rylruu9P67mtCgjaitBmM2AkBUBw/Qph8rWL+Y14A1rCpGTwjAfjDvXPdirWLLrF
joug4jVH4sx1ZVlp12IrNcn37NxAl17tqKG3OKZg/LwINXT03PydBXbYFnO4ocRe
8jJftqaueSrURvEMom3Z82x7s2m6aO5XcWNN0DGB+oPEkkcFJXrG7VC8Zl4Cem1k
byn/wDpbh616hJtQWys52D8yx5TvKHQpdSa6sjT5Ju0ZAcmTBER9phkb03hBC60w
H5Xpc1NXAEbFLAt5H2JYZMEF+DTteZBQA06QGjBQO97wVOsGfmIsBEv9T/MQqWgh
nNNip76wzTLpV2o6rAC9vfF04BejABEQi3UQRqwQ6PNw84YOQE2nY11iDb9+yhEe
sa/w4An8NCouTKeMSx37fysISxdJFaS1MrMGMa9EMOI5oYX/0hcHa7dh64lol2kt
qbzH5ZKK1YwhKq9rvYipIv3/hakXEnHVQxmd4dRoBE5r/ales5ceCSRXHJ2DZWdq
C4wP17ClIgcQUoWTUJwYQJEC8ALqsm7eDzazHWuhoZV55AdHTjC7k0N9t5b95ofV
KBL98uCHlEpjFgymDkCzhJd6hwvLLTOQL/M2kem30NhX3lyCFTfywbdBGV9jyfeK
1tjx6TpqNHiST2eqqizqf7NiKND7QhfIyUdcIu/LPx2q3d72aXHoY8gJbCMCRK9l
9Dq90SQgAKxJSP9n5mnMOU6Pd7WiCtZ19E0DGDqlg5KpD14ORmCmTpGoBf3pm9e5
LdNe7WyIi01pARpfbaTMsGlZ/po9SnGydcHMAA5S0mlFa4admG0qeMR0UsMNm0CU
xlJElQw4wDNmuE4Ct8WjJ6XyeY/12WlhJNu3KRTbfjxi7+6pLKEXBkZooLqKxVK/
BGJneGYFUj/PsiuWdkJtoPM4LmBmQsPfBOy3GAwGPfXYzSd/+sisVGquSz58E6/3
5JLDWos71cZz2pgCG5JuPak+8HHVAbMrq/OSGsxNeeDu2HoTFxy8FXIll4ukZrUK
8LttDG8KrqhyKeMMZVm3c2buJxUgmpqA1TX0oUTr0qQ4cP4Sl/tpPKZgblko7yXl
Fr0xVAp/T5VE8ivp23D7VJ2s8jpqNHPS6ZD5J0f91oQPyY0CLz4zdnEbpMxVJXQs
2B+qEd9Ls03CaOJsTdIZYPdNu/h9N4fUs/FM8X4s2PYgf8klu1IgNTZXjsVkwEKy
pR2XrGLEBWUTHVhzjjCuZ8yQt3yqExTT+vxcsvMll/jG0XiqNxeAgZ37mX7hTPlV
37caKkUrG5XKfnle+Hhz2/5Jz0zP8fukZF9GBmPwOsEh73IReN4JXv6uROMBOR05
GPLDSe3k+YhGU60p5oNyLgR4N+d4nhwBw1fGbZX1bdl2u1kLf/de/393bDJ/tz43
VtspAEHIxLalkpRaymnmxRyl3Pz3Gbbyaq86iysA7URY2Kxg4fDIjp+lBu/TGlYg
tQHWjbhmyQWiUdw9fTM9Oby5ih7Rjua+OD+7ZsSMBZq2Ec+XtpNCuQtXObD2BdjF
1rBAYoZASaJ3HoISr2H7yQVKqp2a57LgrTVBCyWnKTh4s2nCD/yJh1QlPW7eHGOq
U48WY30byz/NvYKuvsXyJAnz9dqF7igLbUEJqNEkK6yJ8LwMTXcjAO8PCr2lgoQ8
OMF8ysDup4Nu94PlpkUgeainVujfLcqFR22UfStAZ02CROA6nq5W6gz/Oee5SUc7
YJaldnncC10Ipci4hoFoPy90mboDwd0zwKgKYX8/Hm7VR8kmGhuRWelEnpTZStFZ
nL5XlJdiVFejDEtYzf+lqfDlPBNlWDqmOSIPKFP2PafhP9v+3XE/kbZ0fkGwszm+
gouxdXZZVipNn0UIqXmsUPLpFEt0NiFb/wB3ZOmF6n03u3CQ5I3pXkVUC3LhHV0H
/K9hMxxo+byWXwrMHFuVvITKll1/BGcfYKqZ1uJ7rpZLUmowDU4pJpo7EbROt1Vw
lXhXRysqm9Ul1tcNJFQoIrpEqRcu/45B+wBWJBSs8r9RTtOt4lOsCOUCGiJoiBzE
vjlW34k+pamZOQWlVlbnX/qRjHnUysbEkYvINOiFqyxt+Twd3Y97fh/xEclTQ0lQ
c0jy75xo2AYOFt6MCaGEncDpAd2UeHvYEOWUubUUpLRvEoYCaIo/MtzMLSCw7M+z
N+83itTBVRBiiitrn7W5NoOwO2wr5L0cUsi0bw5TKBvpLaRv4cMVHTiXdsKdvtG6
v6yz/6cv1qaKfil/UjJdL/aXlVsa4K09FdUwypiNIG+tm7Xk5noeGE4xbCrcHBRj
a1t6injBxMU8t06OSNW7ehkEPrd6km6QewpgdIH4Z29AcBLsln5v7g6325XEQ9TB
mmyg2Vp4P4jb6ZRXQ5Xy2niqFn92agDimL9ct5263+ezfvxJM4n4680zAH/UCDE2
bDoqYLQqioCGelmDWGMymXALuj8EM1syGrThxano6CIXFtX2nXorO4mynMAY81tJ
aZHpFMk0XGVkUfWEpnr6ePw7jLGLBb8qd5I1RaOLAi8kT9C9tHNls0e+9JTA39yH
UC4I4k1KI5TNU3UFI4tLR3J3XkPrsB1ao7ZzAzeIrjOkobj88XfrZOHj3nUsvn8c
A+YtV27sveCOEjZutQ9ZjTwpP5wAbrITZjhSACSiytBnJ3JaV1Qnm6uGW2PxkJIb
lgZj+kL+0vikVwoNke9JthVSxzLzT0A7jB05+Mx5mVm2FF0j1tszreoJmv6MbMb9
cjb5hR4gLLuJU2Ha/S3xelvB8PHzirF1GmChEFoPSUH/r8EJ+qPEIg4hnP9buCYi
uktnmUhKc9z7/Z0i3WkSxsVhCF8RnP2V6ZLiLz2VqmezVsz0IZCXjGyH3j7xLeSc
RKZh5ySMJ3V4+uDoUDrD+Z3oFEFMtacDQuqH2acPAl8zKoHQ7IM8rmpk5Lwo4rhb
e1ELvNDKIPHCV+JD6DE0AOIG57n9LcpUdRxfzT8Y+c158w2/HxCHe0VFCvsp/eS/
2pMnzByjOWftpZpHmualnjcQOUuoWpqEfZKNgWwM7Sv/5ok59UfPEE3GB/CztU7P
Ma6hmlVczDe6w+2hyZ6IKADaxQVxratCAuZqWJW1QK+IKAIhdvuTKmQjBaQq9TS5
DYwWnKlz3hLGW3rCXRjlrCOCbcHZpxYOr8qLgSaoMEhG++K0rN1rdr/uOSGqWcp/
3wn9EypV737QRZTrEFAs+R6f/epPiYtHsugNg+Ds9aj6PpWLxciVS1b9VyVty6TE
KbJjK7FBntc4vzKBMnOyPZg5OfJ4IL+fThWXt9SLZy+6/VQoaFzJzZSBiLfcmwLq
+EFSTnUQlPSWymeBMIQvJvjq1ijSn5le/5TzBZpf5B2SbrN1bfRGRsLIObhR/xDw
EoiZgEsWbWBzkK4+egF1xAxR3P61qZBZOzgkRtxdtFaYjNKEFkap6f2WltkhzBH6
3sw/0LEcpq1/XkJ/IQDGjR0XOTphqsXCj4ksklEBwlToYZIQZt9ZpCJcaWoBqM0H
Vr3NmGf5mIeWWTV2yr51K93Ry5hQWvXtmiXoaHxPI4Bs1u1wtRbvNSjI9ji48aP8
VWBhveCKRdPyjCpRiIrmMjxX07kJm/XUT2kEF/SHUBE4yVz+q2aPyCP+lT0jMzr7
MCIWUNJL7/dW1TV4jLvFuTG2UaQEuOuI4/apHmfcxrSvd+YUQ4wm/WEZ2UGY/HRe
jTdS9snqrQllD4Go5/LvqcnmEJRjvdMPT/hyyDd5BIMmKjSiGsR7KVu9PlvlWPwy
zuvviFySy36haSGU1V2+4yfrUmbFTUw88Xi0Hxl9PrPldbQbs5M4EmBTjt/PQBU4
jRb8uqDd8p42TR7ZmzWdtQ6t/ycmnxNKB2HH1EVpNIV29PIBMLxbYnGl85Iiuopj
+1VbgUNUrv1E1Ybr7BViv//UmrsyPIou07ZoqRt6uKE41s/E3p7Dw1rwTLQgsvJL
ro8SyncMfeQfvn/jL8u/8kxxhPV4tSq44k4nfexXglUcaLk+BFHp2KqmtLi5QrFC
jLioaZw20LZlvaca3XCLWOnLdyAdddUnPccZK2ZLlumGIcgyGERBMi68ZmlfCWIb
FYoUSJsy/5rYdJBEZTuG9xGEFJNETSIahyUcCaN6E06YvtisYPCLkmBUhvOIte3M
BP6pDxGUj1Wmdo6bXa6BIIo895266pqxmrkw1v2EhrEPWKHHizLU5qROtJwioLEm
ryyab5cFIpcNDlgmV/WL6mL9ucU+BqFBXiJpQvENve1mUkcv/ciRyVd9Et17Xug/
sA2ElQ0tjljsUoawVcxTIBHwjnNMKvEavl8rf1EVSgMs3w+R8wvN5h3i86UErlkt
fKYQj9hDVWvywAND9NkYC+aFMWKn4dGNnF5T5pCwhgM3g0CLoV1Ae446UBMaM6vk
vKBOJx60W4a5B3sROEtcaJJQ3s65Ajd9TupN2Z7/VOtBt84fpfGSXCl1QJDVjyF4
8x42Lcf1z8VC0m5NSoE68f2LUZFOxgIeCapim+GrVedcHdCBAJ/RultIsOLDnfVp
PScKFZN3lvFvZEAhJFuLf7UWQG13xZadi+tS2UFXoe7NeluXeolqcxhfaDnQsG2/
Yg2bba/6RtxSlTCsBYdQREnornz80POvkps6rshMYsbkxxygiUQFPycYTcwCQ5J0
PtVZb8RJwq8MHIYqZUOfJw1RQOgr4SOCPIQJFIzu9f5Su/J72ntwG+ud4B/Uqxsp
V1Zv37+5pfrPbbtV+CYYEjR1DaLF7FoGtwyVOexOdN7RYiZ9QG6v4bm92ceafFiT
VqmMg8or5ABmLdF0v+P2Ad/vVl8OWSGdbmopPJTDAlYAV2WZbGchjX0oJgbbAWMU
mhGgQuw3UY22Oqr3+cWX9ogmOIRyABTSks2TsB5hQefh24kTgWHinMebmlD3xfAO
V7qBV3HMSTfHTXiXZP28zJXJrKPfrK2qg5pfljh51asXY4yj3lxk1TEHNMMiqasw
/aNrJgSJp13+53Fs3nSGhziWsX3xyWIaTFxc4R2hkHIXFkQBcYjtGwz67mS4C/kB
jL1CEL21K8sUF9u28X1URAp3nZp7PfGX+YdpRf9nF4/j0q2oPdNYxcxilAfBjthh
55nWlh0cG6sBUcMDruJFAPmiYvN5Ng0x8GxYyzQ5Y3D97siAPGCSAibUqr+N0gSU
G+Tpm1M4pffOGnbkniw5aiJQTzY2vKGoVjF6scYIh0Nm0qXOGb+5dIYyvmgTwLLR
Eei5ynW29/o21ZBPfazyCDExfQo8CH7/jfquiDb+qo/ULRVCmt5zdFkl1Ysb/arP
OVRj9z6O9Kc5X1xhui2PTG1zwJDL54P/BNULp/0+//tKD+kWbqoeyWzJm6fq6gzS
arGp2IFFbu/X4OlBhh03wKqKBaEp6IQYQUk22QEPMrOretH9mpo4dDBgv/RzbRqz
zhW+CitcPBJy9fRVldYHgegaWMcQX6uMF28TS7szHGWeE58fzSuG7JjUpCX7S/5X
BNWwFFRPTqzLYEI5BfpwkraBj383DV4jvUnNPaKYw7nXZJO0szxfFngsNtaGiif+
oUUuJ+6BPijrCNgymp17rFqyAZ5yslp2aYnIg5hJix+tvuVK0bVAkNsJrhqBjnvw
BguccUwY78mSO/YYFa5XTRWJoJYB+r1xiNe4NT7TuCFQhsdufURPhqcAJnDG3PHE
CJWuUee96I3+35+Cv1YaJdYkmrHDiQySgMh86KUdBA0IWvWq+Rwlo6i785ZsqPQP
WB0agZ3s3ahLDyexnstunv0REXPNOLCszzzpRf2LNDRAcKZM6Dm2BjZralcNhrEd
g375Kn9S7HVCb8qr89qZNBa7B6Wq8v3T0b1kYchjVwx562MdFwlOV+hCFfTef6QU
8p3ucQeMjMHNe2JgUrUhaaFiZ90iw3f0gLdRbZXVownUeItNX7FvWBSli4RIGDTZ
epDi4F8//LCdNNytA4mMok8xIpoiW82osLKXKtKi9/N2fUHv2gHaL9tm2qF9nWr8
lh19Tf4Q/z7sfjrrCII0pv8IByn+3FC+0A+EUJSYdy1D7VajKPAQDoAHHaGg8edv
bXg7JX0KGzUCU9JVzpL7zsnAlY1dVkpuJXMLZ+RtKejnnfMdSCZwpNUsgxNTq6x8
HB9SlyieduoZ6A9OW/THwhBNMQaKWo4zY28NsDtudHy/w9ZQIO7M7FPDrA5dUVUY
PYAsHS2wNCDBHCBEKTQdXCduqcy2Q0NdsdHlBcOpF5ujlBnFuEhwLStRqp5FGli+
B0ymY6tTuij3GemvnIOL1lWHDF38DDpFfh/vUty7wzvgDz3uqNVgxLmwuRV6ursb
Et63R9b/ZXkSH6cvw+DOtEqFFTSvUuKjaLbH4oAB4R8/VyLsGdsAupa+l5jhFm44
qXzbFWAR6u1ZQQyYlckltfY7YxmbrJ5E0UvDHcY7owAu07u+hN1lt/IlTj7HV4xn
AI10sqqTaQmJCaQ+0xV71m7oivtBaX+Hve9xw1kYE7tiJKU8aQQmmAn/SkdQRJAF
bqkhlz8P6WZzhwl/fW+c46ZdDCYY/O58P19LZa24InCkh9aCMptLXTiEFgpdMV48
YChno+QXM0JHIXTnv3bM88FLUqKHIo4639lo96+ecyfUNm1CWdC/E/0BPlypmsT3
/zHmXf3OPWb2FRT+FpjBY6cMq4xR350DABkdp2R9NrmCCg2vlVeLUshG6luO90HQ
i2mYx1zO7QsHC4kpXDkTDIz1NjxAFIrtFzwxGA1Q2uQbtfColjXR8/hngiJSrePy
UfG8dSSEDV1Df+FZiSWzPHZeAEboCW3YIb/hB8doiV855zuhWBCqSYQkubqibAft
XCy/SsK+2ySPWupUlOpnSte78EEZKiuSvxQOkBOBHkLVAe72bGQgmd0CkEYhsdRK
IlmVxF0ymjhHzipeK6i6a6B8boEFGksNMrSkPwdbMBezJEvoKG2Iefr6MJjZevh/
GqWhEcUXKOr8GaMOu9VAr2lc0lvETKzt0tVPDFo7G0V7FPT5gBRcdCtgYkEX8Yfr
OyjHBN/n+dAkSBYfifRXG70Kao6HPQHMkFHhxRdtpAKh0FH/nOU+r4MdW1j0YK3D
Im9FXEfzCUhc7k95opDWeA92yiLM4GJQIPbVlouq4csuK/T+97t/uIoItgAc80Q3
v5sg22Y1t2xu7XvoF6N1qtqS3aXlsoVa0JBms3h67hSs0OKLZXDviqrMmZ/tU9U8
Fngf1fOKW3A8Y36OFUiZ34/9xiJRHPi+hKkrBiD/3evpX5JHZXPXiqzHBvY7fGgF
7ZZZ5mMWK/4sp2n1a7wWZlmT+9rhwGiOA/f3xPWFbtpqfYWrYVFORZQKiLv4DV/7
wwwyDFDiyCogJZwYcGBOneSlUR2rQly7KMim2KNMbvd3UfK/GLxfTCgY7r2Pd115
CFc90jdwZe2V9L9O4vart6klNwsIJy9m4OKr/ivBqfMinsJ2yR0z2nk8SFB/+Blx
w6tksi7Kd+M890o7ivWmMYwrMplXOdx4joms7QJLJC4QSR6eL4GAlaGHg9gz0OA+
33Tb7HZaplOShVXKKS6H73LdrZXDpeyctKPmxK2eRKo6Xn7mh4VkFMWrJutv6pMI
uuJzv8ijDk9qEyIfwq8t7D8vJ/OHXNxMRtm0fPgNNMf/we50BArnk0cEnAIeWnH4
XypGMW8YVb9WMOQbtsqN5KUToWw4frUl9nkL7LFGicXuBRQ2SiTy8IEPP1aqEom1
v6l3cpdrJ8eVZh7IyS1bb2VpdBhc8MRYOXgd47UmncDSMSkcb2rDv9O4lAn0N+iJ
caoxSt0diz3npfSB61A7nEYRaB7moHxP8yB3WGtFOCE2iPGrsqN/RbfJsVKqGyYZ
RLxRiwZWMNxU9Xkn7Xn0/3x27XfTEbaOtKnX3k3xqeTmXsW6TUP+A3HWqV0PJjYV
OIsoZ8Bh9nq2kDkx2pifmObYzjWrxAvrzsj3NUrK41XTxW0oN6ulV7+N/cMafqcX
kcmYSh9rHHxuKlz32auBTuYYEhR87slHZF5LCMTQ027ym3Iz1ofvknJ8uAKX3W2S
WjMntVeQHdpx6wrnZRHLGnfo7D5VoZbHCL9EpllC0V7aePY15n6UYFKKi4fM/4rm
CSkUqNo36+2tlJcgmfl69xnawDA+gu4pSgCMBZQwN2Y26O2xaAd6zKrbFipvm270
13Xh9ux9C3vCt24h8/AfYwF81pTZjqFxAeOg4xDr72BvlHex+rMKKsYVb3oPLJH/
IuUZwWsB6S44ZGD/NfD6e+HKSzIp6KID0VRtRVCl/+upJuSSKhZ4w/ND77Kw/VS/
yFN1VbF/K+M5YlVFlXCe/hclni0uONcWbWr8tKIO/x30c9TXYKoygNomqDC0YxuH
I8vLITtPC5PFDL3oY2tfDS/w/j1kZZtzXsml+QTRw1QQOVzakoLVPAYyJVuHJLm+
G/J8wotzoh7ZOG6o0uX2pKgYbq8Quzt1EPJEgQ3Jp0AnqT8RYGfiYYWVqClquVlm
K45zqhdfz9Y+U6GMwZZzIo2kyqC4AcUg8UvutEoKa8L0aOr7uwRXAzVXJSAu2l5f
q4HFPsLVDYa8kpPnFkhSybV9Mqaae6mywl/eKsHtgy5vmQ0sP2+T65mVCjDMCoXC
ZMkxOSLhvlUEyVHUxNjoSiML33QxmBYXN9ld8WxuL35u9Qv0wfv2OKu+12c0sHNb
qy7H3NW2+/Dcw3NjYzHc/XAiTVUJfPefVrS0G+jAKb2wXGTdTKN2euKpVt5EO18A
oWaI/xf2WvGpL1yahvC/vWDe7mmtVLrJ7W/B3jpIz3SqBwVXeOG0xLWYyvZGYYG7
0Gj876j04q2uum9m9Fj4waQ1Izq7WYvbzjz9RKuQXA7aZzVWRLC8qW4Qu6gP9B5u
MQS96nX8oCe/wTTkLm18xv+lk5sFl9yyHqc1i9MLie/U6+c6rBXvFZWqZIKGoHjD
063BOlmllEKT7gVIwV0L6ABJ+qXM6Z/yURR4Bv+LjWphSmgXPmQUygiu8S2AJJ+u
BTGtJbtXUZxHpa84odtmwqHzGII9icgDiX5rz7xddznBD6zviVi6LXbEfOYctwM5
AmYqd2PNVxWvjsu6Qp4ah55GLLW5BhfLcz2ivBiDBmekodvpDSB9Vtb4yYSmo369
G2MDG015O4Cj1pZHfyEVXdlIQsd1TWJxjSCv2AOV6SKEayKZRMaeKRCbs6eRXQHw
KpWo/wdvDUlXjeNDXQBY7ALCU3ZKuJPzLwQUjV0w+Fb+b/k5DPJUMzUynD01O/vR
g4akTBPYGzDM5UueWIVfp/WhPduwU2bzLpvisL4FwYnOgMXlkVAv2uOVeK7JgeEB
cmZ+YCKBZVdU6EUAb1Fu3INcH/SrajdUqtbioSwqCCihn8NBG1GhK7Yv5Br6SK9A
WtC+X0j/balzuFAWgaMZ5voFF8n+/LzKgFbaVQGI/wODCM7fRkFZ9YPU46G3FWwv
UjcJIPq5Map/5XVIR4kQmaWp1xI+uwu7MgFXPO226+0jKRhmUMpGMwvcrI6Sp1rM
/PFjEId8xN205eSAL4k4FKnpdQxZaeGeCkq22BRcg5BlvFftY+l9SrfE71divZYe
gzmW+6lK6UpNAE2szdR3i+CewLO/TJ9RaIbHBcNmw/24RLEv7ZTDcfLPhLomU2oP
bSdr/Lj4wpZ8+f1Ag9KgA3Ya0i13NwnPSnSghKbBEbPtPsV9iDSeNxPrny4MkB7C
PR5FYXltnDPV7m4CH2aITEpL9QxG7yrxrX8GV96QCoMrZhLTgLrIy+TZ5UVmr8t2
nF8+gT8Cn00rkygksBrbRqRZHYuRS4z8Vjcf/z9s63mFVYecpiDx626XIcegGO6s
j5LCa3hbqvCXEW4Y5X/yvPDhpWs/9v3afR5KfzBL0Pd3rG/p6oPPe8F2s/X9g51E
RsXDYno7GjXs8Z7bb+fxBcIc5a63H55CcFPjiHRqWZCk/TnO8vUqydPI6bw4fyrU
UvlPbpQ0uuZ/3hvUkM06b1Jl31eX5ZSuw2DW8eAh6ZhHbM1t03s2Lk0LFEqLsu88
tz8vtKFjxcvRdnkUwGDlZncvRK+4ajBrjUy3DvXRz4UWygmIEBIMpRaWdEYMj1Fh
onG6Ums9Pi7IZdZTq4oMLIVqd+9/oBm77NqtlRqyL4NQlreiIJiK/DdacDPuSB4r
ePodnnnbTtbb1QHPZincQb1Grh6c1mEQyJ74LgL+Ncw7TYgomvclZ45PYqFX3QyN
APfaR7Cw0e9ZFflUhwScdJ/2prALMK9gxNkxS8TB1LJb5OIEQqDIz+cEbHk6s1Ag
TVJ7sXGPPjnqjiohi86utx5mtZzGRIMaTnG/XiF4znP22mhWO6GvPKozXznyFni4
H88TyjnOFylSAAcjIeccIK5E3sUKMLZTPaU6qXZBH0k2kVTUW6mPmHpQXmbHhioI
xD4NRexnU8NYshk94vOPZZM2eHALyfreSTZbTWFXuCoETtfojXQSqulovXP5NFO/
DDwJjkjs58bPCMdMXrQEPX2sl06Si5lbUngbPpsGFMJMxO1/D82G3vFIUHPmiq6K
025EwWygOt6v7JRONQBJdjWlSJ2FRUR9JKq9I0xOohWs9N25U21iLy5n0yBDDHDd
EmXEt+DDGOzhPaoQttfsPQTE+Gswt6y/1rh3TBipRca819brJl45SFGs3a4O/mU7
5TtN2VWfN32fg+CDDdSPzRA5n/Y0zQ0H2qr8augluHJk8rfJXZlJMwq/qj/D6G/I
HfiyAIDl0qvvAwXeNbDF4iUrqPKSyYag71ROaai7l3awRMkyRv0B0FkKJ+FNXvqa
I1Kn6qVgESvb/kRzKjbDtBzjy9PAhIXZrIyGBelyAoFsGniT7bFwNeavvERoTJRl
DcfDnFYz1TlN4XCuwLDNrTppRDm8nkjmIOVCIZ4AjkH8X8+w/C7GUsjbrPfSgsPj
7b9brdkpTpCwqU9qOW4uF8WSo3HU9va5uODNIBiTl70qLKgKHAtUOd2dn9mVzkww
ZSp665u22OglNdqRphK29MnmMEPng40i29lQ5zKKEhA2rMBvHCPJYFPRivOTaLWR
/IdOCzFGbIL4EoczFoRL4w3Oxz9DltL4gxZh0XOU0hbsu9Ryu/HVMy11L9oiC51o
j3gg59BgxUfui8CrH0rneV3va4YPkNgrP9N7UOHtpPmBDASZ2aV3LdyQph4ZsHzy
vYRJIjJlWlj9LwjZ5EWJagkblf5dX7nV8Rf/yMLjo9/w7agipLREqQ7rroGHG4EO
6CbRW8ZONT+fG6Z0y9hV9QIYkKDdjX9cTztid7jcwJEmCtUDuvsD1D6Hg6spc7TM
vG3YjXpWo8KGMYi8czFXX0zerTXlu+Asj7ddN+cBdVzVRLk37sLDa+PLF/95LYyU
zLUjFPbXlOvNm8HgqZX3EEN1VORnD9Bh0WgL7IVRUhuAjFvTinia725nYVM4OlNl
S+0eA4axMSeQMFNK0ynZ3ofCBAEsPSce2Jr43JbiagM9TNnkJzOvPiummf1z3jNt
+WKDcJ6rQLrdZzK+qJLXbBzqC6V/JhePpEAtA998MW4dz5X16bpI82C9MXVJLlW4
3UabWTfmN0GmAp+xB37wqw96AQKS7EVBu4Nt4bBCUXwBVwcTOsBZ1l+U9fht8sKJ
q04k8CrQt9nG3si2AD3J+Qo28AZj4MKqC8QpIL7Fp6H1VFdnN2Qp3EiauqniHhSM
sc5Ww305XPDlDoboKYMe16nokiQoYdnvwnJph+6hVXfE3KHle48p2CPbypE6qIQ2
JqyFWyINdEcYNRW+X5JbABQJxee2klH50oilWiwSJkmG5GZpLh5p4V5PNq1+UgPR
44gmR89i/49aNV+WwuRaavNFzsIg7JD1Jn3ZqcWb8PkWhphnH5uwcnaDGdVfaic0
lRB4QGRkaTFWl9Fgp7JvF3WQKsEj0nZZWCokQTmxxt91xstsCWacn0fKw8bjUhPX
WpGKH/THC2VFz7Pr/PlaGK1YWyGCIM5RyA7yIQUdTn3Slqu+mhfeJ3b31GDVd+j+
s9Z0Y95LZkl9a6yMxN08ZLJE9vVnd0LjEoXMA05d+5v8ePotYMHV4MWBq93S4EhY
r1h/Th8rEe+5LWgg9GTNXF46i2tzC9Mu1ok4PoY/TmwmMwbyUGX8jUJ+NKM/ic9a
y6FeuYAzuUDMw+USP9qo6o3psqW0lt7ofpfdyLcCFyJlBSVRghrGz4vzXyekTEVb
Z5paQliobyawvO5v6k+7ORniIbCLfMuDKuJS9sQbl/xMviKOHzDc2VIclk/8NT2c
KlvQUe7RylhA5t1A8KJll8vriiW4WGJIDoE//bzdO/tpDH4S1hZryk9byi4xwWiP
f6c0/ohx9UDsibmu/MmsIeZNzjOSUtIIo3N3m1CdC6GGNseT4NJMTspRPiLaG1iA
KiaTh6zjf+fGNe51TvLvpQk9IjPlWln5SMklmT6eQaC4kVoh/63AmF8LLpcICO7O
uY4V1RiYh7lPT2wm5L+X+ZwIdS9xjHentzmgl4WM0HKOfzv/FJh4W3EaXfs5D3UI
9DBWEm35goFZwe4AU7EGEMqkd3GgsfB/Bzfxe3pMpRXpNXJmG+pP+gvfJkVrvJvB
zrm2YQJHWux8ElxWDGJ5s6LBItgv4722cvwEOs7czs3voJM9Fq/crv8nJvzfx6Vp
gvWoYMXiWg5A4N/qDYggkGNkx6r4Iirp3jpc6fEJdMxl5Nk3a6Qx+DE57DGPPfp9
7aVZ53tU/k7DNfdRa0Xfcd5eI6BiAL1EOHcMA9G5i8XNs3zVWlUJlyFYczFxkOUJ
pctYJ1st+m2NdUtIeCkswpwutwOMetdZtXa5co3cSxFOEpLL0K/ZQZtgvkWammlQ
dIPPT+ULNVvFrLnqspJptSRYRCdqvcMR6bOyDp1QHEo+SN5oS3uZ6o6XEueP6spG
/pcMfI3H6Zi/YjVjNjqo+Bgz2Yxr0MTta2UqxHp03BD6elzoOrzCoS/YG4dgHNxF
P+cGzg6rRsPezzzpWpOWq1TswMNVH6NBEexgn9yfiGbFA4FNQZBU058F9Sz0HCHK
TO4GiIbVWD24cGNH4IxLieoSSzZtq7eSZdNFMLm+3oW++yok5p/MqsCTHWWqBF5j
ltlwq9SAkaupCUUP3BoBBHNndDBAvl/ZqtrjSKe+4U0OazaopAjaCl2oSMj2KJaQ
fHbTA530ZvNjKeO6gUdjs2sXGY7uAeSAQzxaTps1JQE4IQxhv6Tc4p/F3NqTOLGC
oaONL8J1veiciT85iTwchv8LXzQYA8iUm0ayRthjpSt1+H7UbXWU2mSVw/NNoz/4
wQkeCTAURQ8sFNeQ4JOkOHEyzi+koRxHgYKlkdiZFYwt76vttEDQJFNc0fZO/NmC
2axkNl3QemZ5l0W6T3gfTHa9WomR3szjjJXn7moPprIzLOgcjKQHVELHwvAZgPfL
X2175RUj7QKr9/zYocQTZUHduyBmKNwcuHHM3Futj0pKz0Z4sSyxN8sFim1O0/Az
4dZIogSDmfQKIlBTMwTkF6hYmQsAgZl7S1L5788/20sLdTrw6ER08TIVx5/eOgNd
1Z0hstccFHF33suYiuo8ecdJGmchHZfhWrCGqrxm90HicDuvO/zl3CmJIF8Sy3jz
Rg/CVVkqJcoCzjDQ/fG2vOaY/G4Tpm5VlFCicRdWGuWYrQZvUCm/M3w7WGeKKDDk
p2XIg4avALrK38Gz+Lrew71zf7dDtg8GpCZiGYU+gkv2gdne+JnmqD6sGwP+up5o
2byjY1c8qmfsLis7FfSrzDaUxhozbvJNEzZs5nKBZWrM3DGf3uZhashzr/Hcb8dl
NaCN2NI+PW6Wx3GuyDYBwU75wZWN+vMKhlKMMJM5JEdp+IvpBFJFMqcz/AzYqA3p
moWrJAX5KTaCkrC4/F28JvdvlsUKvSzbRPEqFynCDiCKX2V8nS7iJvltdmmquhJJ
HPfTNDciLiao3r0jg6xNCbJy9FJF4C+7N+LcD0oM/CcGdFpxVnUN1mf6ur/kHJ8B
jcCxHLKTWTT6ZusIPDKx2xdTVq/myV39LabgPJUJA1cUjts/yYEnK6vnQh1lNZEw
IXBlnBLrPfShWPmn+3Iak+GFlnDYpLQTQc1aycpWvlPI517kQi4XNwCWA0zTWKE4
mbMUgLb1sruprfg+vJ3Gu4Yx9H2rl7I3ox5esJL8r9dkunFCgsWg8iHt3FfzWZzP
V6khpkkPYwBYO9QOFlMbp7ihNajSFIcIY0dIRsNfWlbtSBhG34agDh6eDP0mUsZf
c7R+eQqGPEkfr16qbN1+pf+l+8BoBs84fiKMoZSrKzqgZDAKuqZQIcM4lxMyLBfa
mRuhDfqX9xcldEs9Qc93mKeGYiA17ey4UgKmiHwkYkO0cQ2jVwtnkSVJOv0HuT5c
qb3cbSCdDYOZ5LW01rxo1OXTw3gSi04YJjdCF5CgQ4ezdjYlC0Hi2cEP1oRjdNCv
ij2wZ2QA6vgAD36P5UX22djlaVyXKAvmGddkvBCUA7GXULZptapqNNSiR3WBJLry
VWWWvHSc0yZpuqV2s8KA+pS+jYzFbyRNrLAeuPsebdhFUZUW8IJSjs5FpSK1SLtr
SI13sfHUBY1B5kB2UbCghD0Ep1vjsksqEC8iAZ9SuOTdPn0UbgaCi4qbFNXgnmeA
/OnaQuX+82iAxgS70pmBtSCjk5zkz7H0CrXLrFN1RR++Q2P91XMqSaOZX6ml1gef
M/KKfSYulmAYMEXcVbGWM+AOGg0xTslq0a6xfR6gB8b3UGuiLcR8lMDE/68CYuSI
wgpE4sc0b92yzHnvoXH7koj2nj9pQ12G/HMbnab1ksjC2xl8pCDYSfja7aiIbU+P
l5C12IlCJwrMQ7ndLz2PsgZi3OMnDJozl2ro87REsQcrny1NJQMGjYjWG0xlSdbT
EIwijrjzMDJECGf0oL8TSqSGzf3pGg11OstPizYY1ZR4T6R5/DDuAz1DoQChc2UP
NETGEevTz199IzNRCxEPIE28tPPhWaBsq6n4E4/LzHd8vGvTsreuvEhDfDpPsFEQ
JChkdrOdW+W9JYxNhPDDCvkMhZ/MYYhp0fR5jNj+UzLjNFGTSr2kgv8Od46NMG6p
eVsDkVMeJqOYkMQnUk19sNP3wSTA9eCZjOqL9AiAQA+SL1YtRVyNNj7jYSrwptpq
z6U4PUOJ7zjqW0GZ/Spk7ok9ywqSrI306lpiY0rS1kL8SrG31Pnlt/HnJzx426RO
p7EddoC4be1MwObQ2FaNorwQwo7yTEkugNOLxr3fGp4hLfVd2xWIPeys0eac8PJI
Y2YClO5JZf2NFdfC5Z+pwaQe/laUDEPYziF9o77icqsM9x1bl16QE67ejwRypYTP
UpcQ2mYtnarjmbhoj9hKm+dXIy0eR+oAEMPnTqaUj6f0i1+C3dfBj5UEKC5wnD37
V5kgBQZWne1lvP6rx21W48NWJ/rlqdKYIc0rl02A60sggOtnxkZG0a+PCqicrwAc
oyFsjUy1nDBPUqjiKX2+ZhL2SLAVkGCZj9/+0MfTsprqzatm1Obv2HlwRdCogskA
92MRbe7AgpHLFVJPYreKRs5UHPD2H18ZgVhExKIHd6V4YcgzwXmvvUMsZg9klfFW
RTmYszRSAdAWS6xYtO5aoi8nO4KrASrBf1NYIBpQ38OqQUmTLFiH7B82jQzXVF97
kut+Q0WdT79czGS18mgxWyTa5X5dCfmXZiQ18UR4voHSRVJ+7NLPlS1zOJOXZrE2
OeoUnb8QimDnEC0sPYBVOGkbRJYgtCQGewF9lVijwkkhXxbLPreP9liWc7vaPnPj
zV6LG759RyZL7dGimFeDX014Au4zhxox8q6vyWkD1y0FSieBUJGugjoja9jJLBOo
I83HSVcDQmGRiWNm69lsU9vATZ2M9CWkT9x09BnTsvNqs+eTeBvS68GjNHHqocRJ
/6Yt0R2vivFU0AlGC5QkWDMCww6H+jXfywpW1f4+cF3D3fBoQveBMVP0lTPpT213
0mhvrzeApTPf3Yqyv/L6+FVE1M8/Qdy50Uo+spQrYrXSAWKUJL3YfMTODX40N90L
ffa+67e45Url5WwLR5te4+XDvD0in4cpnJXjQG/61Uq3o0ipJrCd32L5fZc/MekX
Xqw8MDC9Z2vLoZU0jKtGwkQVcYns9dmKXM3eEEqwGM5IuUVlpUOSUrUp/1i4XC8Q
L+Vp5uEhEQhD7sd8Ek3dxzwPdZOu35RJLC7Oj/8+F9zROoNrlvDUSCFUhBQ7VC++
IlQ9JubJVDk5ddvkXnQo3DcpJhZ6htjDJkKU1jpRh+6COuRmxVz0Xun2YgPgLo2u
AUxxZ//x2HRRJ5x+fBAFSr1bZt5oydH8q7IoivS7GYauqJ22LKajQrPCioDS5r35
YoC2jGBdVYdj85TrnY18rKI1RLGSsDGlBikCY9c/ptC5oTJj55J49+C/HnsXVlhH
Gxa+SoK5wr/7+GWQ8sfbrzShNMEKw0RrbQFoxHdwy0DoetbBOGU2SdSfYZyJmqYz
QJaHR29dNUvAUD4ROg2vIb5YPjM9RaBsD3+GkF0+2GVoqy+fEuILac2jfZ6B8uQ6
tGfnuVzHd7j4LZCMeqWy8UFpW/PWkkALnKJz7TwSLtXV7v/flWnUjAaNgQfumohg
41rRFvNiU7N9GoGHC658cvGK3WCUjO1A16lKytUPGcFX6fw7WCYyOFTdc0M1DD3L
O6NjPf6nW/Ay7tmbVVFpbiT4P07BJkaAQXtI8WTUSZ4k2uBzNRy8awjebmrqSsmE
dnuBH3HIn8vfV10wkwzyWLsp/ZD8k3fANIjkfSRF7KzUjzrWRhH0kf4E9NjMGAV5
lQ2rUZN5LGSQwI1PwDfslVFct6M7nkJAcJ3scRJo2fEb1ia8pPv0nri0xLTlYs5l
exYPTcFIw5+Y+yvxSRxsjfVG+Ngsran8S3LpSXgPD0A89wb3JXGyd8y6qIm/u5q6
zlbyAnQHsPkGIQY0yB2fUMLrUQLbJugauhL1Ir+7xwIs398DxMaRwJyt7ioHgUQO
Lo8N418u0cIJsTreQ122yvqFoYAsoCE2aVzaoRinFU+/uhHyYD8tGn7/WrrTPtrn
KQQg2AifbOmalUpehb4S5w0qL6iTGa/aYBNyZsqnMAwgjUdV87cGVOeC1CKcD49X
e5mp2zcfW3rmDzQYL0jG6C+AcDoPBigPbWCXU5Rw6Lw21Ex8xf4txYd8QLnFvqUO
Muednq4qyN/NCL0w/+bMk6/Cu4x3n5hXYvbUKZ82+4fir25kQAWgP/96ZAtMLBxy
WgMyYrpsc+B7HxGuXWLZuh5i7wFPQ+Rl8H75UZzfNgvW3ncDi7JkeY8aJcQqQqqE
KVPDWGjj57f3vus5uJzyLpv2UG7xYTyxvLkdJxgiIC5wk26faHEPU/6EGi51ebXy
fKu5JTPIcE/uFqSbV2/5UY3JsVfEF1+iR2ejUY6iXCGLTBAwURBMAlhndu32+NGY
UrTf3Djxzc3DQ2dRPBcNNuL0n/ptix3EUIMSn7PwGBRV8Hwq3JcAzevnk3tNuJ4o
st8V/sHJSMTPcjUGNUKJSTfxA/acL8vB8BQODtMJgomybDPiE7vi+G8WjQ7f3z78
Yw2astRR6dRdFHJfb6YrIYo2SzJVNzV0tLR+icwH0OtVhz0qsL0QnSCT4m7k6d0e
QxQj5TLZ/qJWxInxJjVuyXoYw0c0s+RymoAL6x6JWr3L3fEQdN843lvIB6mGjXgH
ZtkLpFwolTtBmzeoqupCX2PMgA6zfo4S8KfF5FvW7tgb/JXjoRm12FJfBqC9MAMf
eJ0McGLdfc/EJTM0aJLnbsk3AVnDPLie30Iw/GcRTfP+V4zF4q29lyRyAYPqBjZ+
dPxXelGCepT6WLSKvog7JEiVxGPKMUqY6in9Eb0WkuTVBS39IaHwXnS+8aJe1Lv8
c8i0azc55r8Uh9BFSliYoAQXCzGwnmmM8fxJWOiu1yKvAae218hxeQTfFHG+y0MK
wPuuUTJR4eht+iE3ksLOcQQwK/gSSPsEF5L1uIYa9P54Itik9ZEC2iAuGhjJXS5b
R2jKdRgtv5UwX+tiJS9tx/nKaaBkXiQa4qcbflNlXE11y33DTLPtdb0ZxA5BeBhj
XZNf1Etp7hMYyAZIvlJ146MhFE/OFiIMX6ZG4G9thE8vJx0nmtD+fEvj93icU3zb
fsqp8MkzoyX5w2BgsAAzQozegSOhsRAj6ZzVoCfsPF5YJblQzVJUMxHCpDdmOMnk
WwY8dAnCmF6qHsz3ckenfdgJTpP1P05hYfFP3SMkL/5XLr35XZxKgtmwyq+RRLvK
HHQ+d3/V67VkPymCsiE/Apgcg7kWvyFXlaFUZ1jGDvnln45GwCg037OZn9M72DEb
LdNnItIgYXT0F+7M5tzzIuKbr74hPE+sgMcqI66TVyqbks5GSr2nq6gGk2EwWxZT
FYfEJJKPPHouJdJVQamYUOMqODxdlLVDyi6hBEwoeVMlYbpkqu7nSYU81XJchaKK
ymZudYeAj9GR3fMPXbsuSsw0C4EfN8Qrjciw/9MKJbpKygjYYkNk2DYi8MTNsVCW
wIKoIzO32rldegrNDwQiexteW0+eQNia8Daor4TuPdLUMk7Gk3zWuyX279UFxHAj
t0vxIPlL0C7gijInhQePXLaoXC9zTyJYiLjGoIDu+bnufau1+FMAFRcP8swUGVpB
Muzy14cbg4A2S90p+lomUfjFKZC5DsPRinIP1wU/qWFjVMY9MhD0I44GKq8l149a
Iavqohd7627+LC23zcAs2DbiKi73I1H6Oq69kXtHI70386js42UOK3H5h330L0/a
ssji0/r+tA8xHmopKZqJlyPMZ2oXExzYUNW46NmKeTxIyXIlfs+giuYwez+ePJm8
oH+RgqsUEGqBLTPwiB0UE888IlwymMemOxISzOS/iKhveNqd1bVG75QNcvKIbyHb
OLoFocx3T/FuD3FWP251ZxO8KFGGaabU8EjfZdGeF43VPETsV29dzoZeXsxuE6Y0
1ojtr7uFs6XFUmpkxgannd1/+F2RNMD9so3VhRQ1EM1Cp6MEYiMswoktcTjjmOKP
RBOYhbGEuMl/BncCIONxibnfZ3s0bLp3w/rDmpmnp50ILEwDgGA4RUlQnM4XySJ8
YDjIq9rGZVHvVNvli2bZI3XEcUjr+saK7tzHPKQrlGBcXHLKw3Nkj74jWZ68g1qZ
cfFRQqGqfAOpKIjIEBVmtZpWC59/cLt2n8amqqx7dWTMO0I3et8ZQcgHEvDZuUu7
8FyT+V8bxpRYa9f9gz7ePF3RIKKbKX7X3KkYYRBEhfPJTKizsD9K11t1eVKGAfbd
qJr1M+Rn3+mlfK+A41pzJ7znWagzIocZVQEt8dAULAHfpOu42TrLXbTk+WQcKrss
lNh34LYCWsDUyiZitl2FssGLCZpZA3vElLNPELb89ZH1uqT9E2tgHlJwr565qtOr
oKZtu3SoihKTItowHwWsnWbOS01ZgTHkWalxGGyCe6T2KqJGl9al7BSvqIgzLK8H
QVtmZcbff6rI/bDi6uINRHho3GbuDR1SytcUUUD1qOIkpAeA9vq4W2qNN/zfzRdi
/2pJdpzUviwGBD8m+MFtWzOg0GOhxcH6BGItdbiWqeZrHQ13/9qEPfhZDDxEvwPv
VP7PX2RNtESrnzWHZgDZQZ9//WK/Ll/VEqPXA1BPczAMBFvi5gH6SBz1k0kKj211
jp0MPt+aessM6Lj2KDT/k9gtj3VSYysV8PMPC/OuMzFEC8nFav/ItWbWx7Kf63WK
wxY6MV6tfgk4hL0P9M6v/gMY9prPVpTHOAlIq4i2Pii5NAuoQSTsmgPBFsnzjSzV
27FOG+rvVsFi0e6JtIfBbWmtksizGm80dhM0WYTHrFB36pY4qQ7xJo/h5Lad36gK
yUvxLY4xJEnqir0Wifk0uCe4Gzq2NfYT4vH+4/JDUDRg/D3L/DErBqXPXfFR8bjy
PslUr4tC/ZVzNXU0pMqRX1wsD1qF01q6WrVrhAmNfEmJVPMTPAY8m3sTePjYOo+q
D8Hg7IhxdDG9PMJnIg26Sw/wDmeHdWXmJG9pNrhslceX93HNq3B5//rPKwL6GbfY
P04hfx6S+gfMPHAYbYjv798lFK43LBrNaGKnAg5cLjoBazvhg9ntgkrgh9W575tP
sOaThYe6K2Gp1mBopoH7uJMceIhehg+92KPUyoaJ2UidcKFXsIRnbT/Kt+S0eXXL
eFvlZKowhxd7Y9o08urGNl2xQVObFXjhYlkiVor7yVxnMS1g5lGb7poQSidrvhWv
pRvnV7ypTn6KEskRs6ZxMubqk851nle8E9xh8fD1+/i8hEZSCehgQa5FWXUGQT4D
S3N24cMd+gdRazVv0KvVDiOwqoqojyrwPRG05wNRp1Jubp+CbdONwb9KL9vLHB6K
86xbLCkPFzy50tCiz2obJ28siZbxVUNd0/wNud4saori5c4kP2w5h88yvwjHsKqr
Nox9mbIratnuZ98QsKsDTYpjeqCGypsiJ0Yes2AGsaOb7BE8uKM6IPbG/24aYkw0
IAhBxjRF19REp2FjfydftfTzRWQ/Wq+e3Mp2DiJFoHm5R1ccapBqBdX9ai9/+hgj
gyqxpJYAw+yQILN0oDGhRDXXYStdGE4OZculCUyyC6uc+9AWibHB0xRQLWQR2oG3
h3eNMWPIfUPJgzhRiPyNSsnBOYmVftic3p9jCfwhxKrV22I9Qc3X7sVHeD8S2ZUG
lKuNrPrDHCVVO6biKg6XcjX3xgJT65h4CGoP5RBCkFLT2fLoKW/4MAYkA8n5Yh8l
AbsDX/XnB/xPMkp98nC/sKv1JhJeXszf38KtIvhrp5ZEjeekZl3d9PMlsoWXKpPL
SgHvP8YXPJjP1plFM+tcGGRToSMqPIFwtLwAN9D6eEZ4XxFK9h+mkYeryZqsJxf8
sXxRT2rdY4i6XIYnv8iEpKs0mU3Yctchum3t03sHkSeYpbu4cLNeqPBk8G0IrtK4
1s53/jjxAAojfxmx5ij/Djl01FoLjqoHK3Ut1kQsyJ3nztHJf0oQVMamBwWNrS08
0u5vEsfcb633iR1YU9ahRHOl2EI+CDfhKXGADxCOLufKNaTw951BGssfgqI8r5C/
XbhujeHlCKTj3itgdHEmjO27cXwf5Sl0NZojCcFQvRmFVz0DPU9p4Y66fCMS4KAe
AyVIDMWG6Eu2R5bLQsuyOZHbZhHXuZxxMUsHnHT8ZyY/VbUfDsQLwRzUP3x31sHV
LCQDRbWRP+BxgHM2uCSvsMIfMegz3xmWGm24SXXIqhoLOVV6qqXxrrkz8fC+3NoA
iFAdwVeIQkAp2O6VFVvD1bZm41kKFNKinUWqthyTJshsGvb2ZB/eO3hxVaAnMl4Z
0a3gwFN+K1BM541C4GHYj4s9NY4iMBZUmJJ0z9f43z9lsZ+WSNT+GYPkS8Cb5qKl
v28zavJv1HZaOyT8CESJB0C+vzR3W7ry+u5/aoyrTtc3W+/Q/hytxZYYfihFQTO0
nwOr2YxFTKEQHA6wpSG++f11vo/aJcB1+UFUlMjVi79+5YGyKU0N2lPEmvoygcNy
MsMikoSMdcWWGWkbVGqPldJV+I2bfqlkB9X7sTfJhYAfjxOo/nhI7quoKjbAbS/i
mTI3Xf/+z7TlVZel68gCk9iLPup9jdq0gk9jtDJi/1W1CiaHGUeK40KzhiAM/Lk5
p6q2CgNoOkMmcuDJ1Akad/S+80l/oBbLLSSHO9oE4Y3kZR9+khR4/7lWJfnSC4Qa
/vGY4akdwgkzUUgDxhj5WJK8xau8Y+DtG85NABOrhDvu94PqKQWYtMRKrP89hOrr
WpqDv2i8+2dBORrj/esmGuFwEsRwAYurz9K1rhZErIEyJZXIm7JW47IoIZkW2mL5
6jZU/m0wpn5KmPUN2AmCkeLlz9bpN7R2DbuYoHcLLJ5bgWUSJqIC/9HUOiD03ys8
xpyhfN0tFCiL4uWUGdf5TXPgahfJhAr4s8EExkAC7QZsXBIF1BhWkcRXmmODLKgd
E1hLbSnnOsNvMm6ZjoSXG6/m+zARJGWG26R1XmcDghVFi2Wn2pIM1St83XbEi99O
QI8vJXW5OFJmXTpvDe1bs4q9IvS++1Q8YF97O70w6jaT/83TsUTTepZKzQWmNXxk
o4KoBaJxALQZ5m58lNg3IABl6aHketMhqN4pKfN1amRZvoFDgZNzKsxT8wZE4uUu
nIs9+bHbpiN151epAFKnT8HX/IOzK6FXPKn3xGHq2LusPo29b0BWw+bEODJ/yMQ2
XxEjae3QRJxfcNUZlFjQ4dK8hEgmFYQj3GHzUHlDz1z16WkuzDa127dfoCgKi6y4
XtqjvYb3I3wOB0OgC+0u4yKh/eKI9A7ZXN0SR2zkwZ6TbSBkD2UgLmrLtNrMhbZV
RImdF30jielBAzcZOOHEvP4kvbiMBCJdMxomtaInEildm+IqTYe2MmNFpM3sY5Rk
E+i8e/TmJCgK3V/7BtPDy1zT3VKX2tD2i5qct2y0HyIYdVgZMDnwos/5zsUp5Jqh
HASi4Q8akUPqoAs76TpJdFp184YnaIDy1AS4bkXb0K2lwKkxVkV+J1pHuZST6X/H
gu9O3trm9Ve9xt14UKJuN6YNrO67ROzh0mfqNW+zWbCNTm1T6NKMQpaQvx002FTk
edJj67sZLuZ76d4SBgppyNpYwm3FuWKktH7jLisLI7H/gJJGDZQNfeQurGprw/jt
d2BakmKrn7QZgDMV9sEBNsjlmRlJ6LaVU0oihu/0Qy37/RYbQMzdv3FetTg12MgD
mZzZ8oCJYFLmh3g2gscy9Bbj+eMkXPqQf6bJ6+rCDrvPVhebf86psIvg354g0zBl
RbYwBIlwXqBPw/NBpxAeiyz5yiuxASMqLRMgwPfUt2E2uNJYGn/YIoeYxALPFsfn
pkANoFY8ouxXRxJJ7KcV4DwPQ7D9YA6egeRI0lGYhtbJgLFxNoE9Wc2Tgzzim9IT
/zBpD0oIPUvYb5CrzB36reobm/QEJVP834tpJPenTYuE93cJJ2QvCeuepNKTBPZH
gw7txiuPtVDKAqsn2C22aW4ksXFD+/IVT/CWG6nw5sozehhxIZ6jT/CBWeqEz00P
l9CzRdGSwP5oreBCl19Qz8UrWIJgeAXeXIuqQlFNukyZ2W0/34m+k1dwC+Q9BnrJ
BaRBGxoVzoU05AIlgxwaclIgV6bJdt4PHRXQp7RorDIfOBJAizbniYwH0RnasjiN
Z+5RGb7X1Bks4zgqUD33+BmksfO9TPOwmpCs1fh32E5ShQSxi/J9P24Uw/n4X9dX
217aoc90ctxUaKWbsuT16NoVOHjQQuA4cRPv5qNv74vvhQiEOZlLMGnMitG3dHuH
V1cJYMLyzMs9GFgj4enXxT32yDDkXCa9ngzM8SOfoWhgAipXJ1QNVYE80ouq2/L8
r6ld700rFaBzx6d4idHE18P6xvkDLOfgulN7BrcyLAWkFEQLTAd4xw+gUlxwjpv4
jID8rwfgE6a1XGL4U+gWExxdXAGpQocCZpBsrfbZQvSlKGCMdeBDfymp0pLk+uTK
aDDADmZ7Y8LCZyeTWeXefDJsHec9Wyw7nTX7MnAHYtQAHm1fTt2r4Wr+tJvygCIu
4gwXiNmaJ0oC3ewZu6aGUREP/LdiSC14nYlP/FLLbHfDxAj2PZPOMMxqnmDCMkPX
kj9F10z2NGQKTlCjKN3RLdS1ZRxSIHBE6HUX1CNQs++Cbrl23plpiCF1R3JLGmYO
nj9XRWZ+VfJgl8Uf3mVtMQ9AjlLtxw98pSdrMRpQkCF02l8qvXW55FDSPyVlBn+T
6gZaRAwTKkK7yQra0MRLpyd4DEE/nQGN6jAIZ+QJcwiOx0rVqmkO0XtYbPQmTDbR
08wrl9BULJc0dWYsIno7XOAOkrdDT7JmZ+nXpANrWJh025G3y5awUHN+4LTCxHXc
VIde0vRHrvHMB8DZnvhBlLNV61OpQC4Yx1z7vBAlPorko3nB2SHSv50OyE9jbe3P
Ad2ZZWwshIDy/s9gJ+VTuwvVIV5hBTbx0yH3p78eiNMyIiiZeOy5VRq9wi56+v8Q
ghThvFGCKVzbPHeJJyVtX8W4JvNrR5plQ1nmm3gCCOptw1zybxF7V+3qUfaYB+Yj
81IdVt4guNtRbbekAJqLhi6xZX7k/+MdQ/vvnr83w0QMxOhXb2nM8SqEIBng395u
Qyf31GqzDOK2uWONAsIWK2WHGRZ4NRQYN9A2OgSBqLbItu35QA0krumICaoJaTYD
0qm+zaGfd1Koabd9mKlKJKK1AZdWpI9IsPtb2il7pJYDs+EvG71/Qb9oUX8+1ORF
1L3/rEcwbCTrz7AeaVBiuuv/lsVZofihiyogrt+gmlsFq5b9pq3AdvmmhcmyP6Xw
RTzZv4xtRAAqGiVDKlfbkJHDLjPzXIiOovC7pK5gJ6ayRr43hYn+rU8Vuc9oIrFP
fP29NoYeBqIPlVD8OvOQXJogmpBFf8nIy/uCiek/qQTWomT7rWBqjyglmS1AWdIT
W0IZft5Lssr13TDHmU0qU4PXuOSf9kL2XJsFlXljMd3BtzUxUqv7A1rkf4zFBKuq
QBaBcAt/giEDm38RxqxqRHoZKo1PVAjR9JnOWjwR5qPBTd8dOKV0wUkVdR/zssXe
tSza5tH1RzDdafg2+OAjlp6p2a272AsSvdohTkYRO0W+q6pZOJKNihFAmSCrYmwX
XM5tcNp7Ltn9NXmQfWbmVFsxElxQ3Rh9vZWFpW2skQ6O9kBPmTFJKo44RNRdKrOc
IY6i96cn17RZmFjPBDsRM+FZDDrmXb/a1oA0uYHXFwD7EtlvGJBG41DPxVAReiZF
Xmw870fUlYeOxW6gslVOyNkZoDIq01bsZov7KhDTCz9hNP5BUSsLYBRLEzkdR8SE
zAm8QxzvIrJYowPUsdg2wl7aW/UAj5X+r10rTD4/hFBqo6YwPJ9VKXLflkrBbYGf
Rhn9+WhFSVBtfT93uqC1ImjhTqEK7DGoCiBg7DW8XvUlxGn+W13T9cIEkTjqkUXo
ItQSGtDXgka90aixHKBtQqnmFGbzoDgBvxakT6+ZocorFudKzL6ANxV7Z7kY8OFy
nCz3Zoek4+JJyv6LPAK/GDawKl1nuTaUDPf97WKMF4xTcCsk/wmnO7l67RGARwPf
tOc6eSWeWrFc0kRvWvbOmYGBhH7BslIh18UXN07YHeumE4ZZi8a8yculZbuyYmjc
3efIlzbArvRprvyhA3+U2Q8+WN8h4TbUukNazI8IWkKBk44imsdAOxHscOmSeAGS
jzbLyKjtg8UcV/dvaERcDy0rdsW+BwgMhrg2OpHc8mSD3NdYeYJwej4iq0/R17DK
xgHxeB8hO6ZuQuruX/OhCmND5+D6EHDeThQDiNkJdkhErIyhC9V/rbI0EOF5ZuLb
UUhotdwePf9CuFmlrJW5Z9GZ5b8pWaMGc+u9NhzLyjVpljTJhWp/sOL23Eup3kji
BRvR3pAmriCF7IGsFBp7KF4eTTrZmU3qvBz+k/sJ0kgWT6knW8cguHXjYduD+0vb
Q81lM5mfknB+XHUy32weOHoeEcqBROV9oDVQRkgxW5iiMWhRGuPZ+HfslR5/nVFz
9aMRcz/7ndVLQSLdO+Sx4XWdp7cOmEPmsd/eEevYqxz7VYKoRnj54qTgsoxV7BBl
awKrxHX0kpC6+zd4VoceHt3XnY1YD8UEVktQOiwfKp2193z8R4av2kjCoFohRBy0
MqORmLDR3XJYoFxxU/MI9OBiYz5cgGZwDsXug5d3TeUMxiuWn9+n0h7QSdVPiWcX
FGmtJ4nQNfCPoz0toVfVD6GoqGBKmIPEhWia4YSU9jqP3OvSIH+J2J+Nf3R8DvTj
ZMZ9PhUKi27wBOvVDdEkSxLiYiew8OMCW5mE7Rw0U+lwiXOaX8+GbcCxtGiHqIAQ
xgExGFTHt8IDUKZzdOVj78CeQAWDDG3/gWFGcJgbJ6kHueeF74Zou7Rq7eGPye7E
cXagRzVfg/WLF5aA694WcRsW5ijvPG/+qHazJXCgilB2c9Bvlh8jWSucI5xi9Iaj
hSYmC6u7DwOXvcBwQckfsos3q4oeSqvqBj17XQQ1Vx2+Skaxip1qo0SOSRI2FLvl
vMRAwHOoDRCOYdFeqOLKLv6mC4C6xzQotk4U45YjHXEKxGC2jf67xZJ3uyEGOZTO
CVG6JqFF+M+MK1RF191kgrOOtl/7U9dAP7hZHg5Nx+syP5OKxomSNprf+lfIlRnC
ciSVSbjFJFbt5S4ZM9+55KZTMzgggz41cbfKiD0WrxghKDEm5eYwsEuruKvktYJp
LTRfm17Hw37cwPb3Sk523vD+EWGUPkZtt07wGnV5LQu4kKNOoVnR/AwZ3vdVArJg
toRNSWAmH1RyampVb5AlMwvvJy4uD40YJ9JNR45HWfRYIfiM1/mRFaSONUUrP7M1
AD1NVZzqt4RlqkILRBYlIv+R5jrBPQTHhi988oOqdu4p5aF0+o7hv6nZ6xOJabP8
ANxWAOJot63fBvRBrbYQ55WDlm4rhZesdsbz+bMVx349hP3Gxxk7anlCQmqfvlFc
Jccbz4FEH46XvkNDTS1aWU1SoJmNEaFs6lN31zBeWZMQo/dqyq4Yi1XtCsCFfMZU
fOUR+iJWLwzq5LIisE3A5e2nUhK7BQdowj7iRnz1RdVZ/eQnlX0pFYwo8P9lBemr
JEMGCpcEOEHPLn9LcLeUg98Fg5/m3em6KIVVR5Unp0IPahsSTn61TvwjHLVAnTWY
2kmvLWaszQMvm0Qvm+68zB5wEHyx0/GDbmB7gI92JQvCs5f/0AzrdFZs0+CvjV6V
4iSOXpw29PrCXEHoN9o2pz/XhdbhJqXrXqgZ0bRni/MMAfOgAyA0Tm275gT9bRiq
XA8xpCOEo7oj84bTxrMk7z2WCyw2UY8Lx7Iu1t62F8ul8IY+YSFrwRODf1gp8kLS
pyBf0wU8Z7DGL2Qok74JNQUD65u6yISfY9uMEyrVmo8V5jwodvY3XIkOYNn3t+h+
wQRdIhMQgnMeODSgEvRs3doGUbhkUqaqWNS4tCGbfdHLn55PyRCZ5aoUfsvmAK9r
yxmFWEBDTVFCnJXXRAgPwy+a1U0/xjGK6U3jrF9pkLopilDs4O6dnJ1QW7HVmkGN
/55qG93rlMLFZJCmZkVIt4B1m9YLvQLV+4pmG66toW13FfENtRLcJuDLYap7vAkx
Mqc+Y0mfyfklV2eWqIJloSAGmTX95kLyhtnZ35QJ0eJj0X4jF//dpwCvKWPijBww
T2//PNpyQgFe9z4tMSPFZrWtKIamTcZH8G5q8LRMHvu+7p/Jx2iiyvKZIaTxIvB9
R8Tgs8R/JhHWBV/SG7kLGQxomWhKkdTEsC4FiBXltRjdFo5vZD5POiE0Ps/HgHP6
3ZyypBErAa3NGI+BXqqfAMiCHEBRAOWi+OT6q/2BvdtOK5EUA6zdq+VmeAnzZnsc
eURkthF7ZwbxRNSoUsf9bo0fwqrHXCjVsIq32J1ByLh4WZIwGtCh6CYzA6fTzwY3
i2pDVskDI0hRaHt5ybNpBbRkPWuorvET/VroJIoZkBkKXWlyLlowsoFREpI9wJXP
MvQzjp6JEWjomfVA+V2eTZqPP8/Fbgpak/p1p1u4FfCEUSY91pLZfqimlRWsf4VX
Y8MxdaGm/zI88RBZ7ciU1em76wBc0qWT3Lo4N+zC6k9N+sUNYZTSUDpI3WjthGWj
kC681I8vWfEcdnC0syi3ZwuFtymtaYS81qkZPKiaGr/VWly+R5Ujomhh4INqKnQY
G0Aa/pxNFZEbUMKYsgaiaa6XhB3AFzcmse8o7LnskWGaDi9dhqtZAvaTf2Pr4ASr
ZCSHaXmuwXQTH/hhz8LSFUCzplRq5sGIrgBu/9Ci8j3SSXxpnnaMMxgy8myBIIsI
2heSSxTp74wM0k6sopSGzWVp1ncTGvpXjeRseDd3N3EAVIxig0Yt/kRO0sB8LO+f
g8YCtvDMwangShmcNUfVVjWm1UTsCxmiEoo9+eLe70E3tDmzqKfR8ZlF54CXQ1Nm
KLA0Q471DqHNd8G6E07lh9Pc0ae1ArHD7SxkLNa+B7X4uidj4eTs8rDMxUdrMEY4
ukMk70/A3jzgUWGBTubdHd815EijyggOkRBXrhP4MmfiW5bPzF7EABRym4CIVo3Z
ZKUMjoqoG908tjt/aC37UJbd0d4A5ra/t6DIlIZd265h6df84+G2osyq51RmBtBB
qKfyeq8pjB9xxuNbOqAAmHflqDr3SeInDoT+05vKNb6FjWG286rAqN82/lAOew60
4j+qXiTYK764BKEgqJMeoLOexeb9ZtkAOtORsKsp8RsUEvWDQvShECu+yjszkSWf
fvL/XYrb+fmpMVswhFY1Z7KOVlDSkBs5S0tZOaDYxvLd8x55WFdCA3SWbfGNnNhk
rKbyCdJkkdM3nFywJxTYevnQNF+CaHil1Pie3+uL/4n5VpwLdVgOFp6uLFu/F7e6
Lut8FnAyK+3nyFSmZ+o4bmfJKtt2o5wb3bumlpvZiKey7tt6VNnYhdDUzTJJrOIt
O0osyldfyEEdQUGt7iBMQAG4QQ8taNDed+7UhARwLbEFlPeS+kkWIyrCzBILBz9i
Sj2FOuHRzJZp4xhDymjDQjs/DlfBE4MzAvG3fAFU6iM0pIPdnaLRmxnsxXYpWsr5
sR/559s3FbLrjrz+G04GWlZcNSA75EN7mxATFmo5v1X+aW9kYTiLhjRXINPguae3
y0jdJakl48pi9ISodJ0gQEKwKEOd5+QGPVDgqtVbkeTnkYHUWhKFOBLQruhr52K8
sFkKT8uAjcyVjZiZWzIC1ceNy3fBAg60bHW3g9diljygrW0aA6ZRFcpxxvcAGEhT
27R3/k0/emk2lHZiAOIvydXWUrRS2wHVj0yP6zLSMtlAIsYGkMi4D32WMoxLmKQX
SIZ8n+lKka30ChzVgKuwNZBM21DBiTWcGf1Fr5Qb+UoNK8N05qtnsfqYtoSIB7Zn
urzEaQL2Akwxo6fdQ8i0ab6916//RLqVDWm2wGDFrkuBOAJLooZMAN4ReFyGHSEN
Q0cr19UM/KftQBBikT1tSxbmdP/4f3N/a5TPjTfzW7JCjen3UU74Sc60Om+LuVls
EWSBZx9yaany26WBsDE06hzbFFg9OGWqsoo88pzt312cf8EFR+v5VbyM0Lc2wu8Z
CRknYNGyf4x0zdbfHjmDMcMFA92IF+A7gKU56Ln0U491lMRQ4jkz25q8IxBv8IbE
t8jmqC14/xFXpVB7AtVVwWpqkgUA+OHa+PuvdJjxhtfO4iIEMkLLOCSjrwHstHHC
1lMMBTvzuDiXM55y0/LvVRmQd2yg8/9orTyVFy89u0mAyHT4xfnrJiznUrlKmfRf
jjHY+g8vqJNfjG7y2rADgjO749zWpCQIbFB40nMoXAYcBrA3QCWCbmo1C3B8sYyr
qmj9oHgMQV33/TbbNN1raqDRbIjzPpu5IYc4Jxpg5iW5X+jAlT4DgRCdCUldQlGK
MHoNbVm8LlMDMlIFrdTPqSh+nRG/T97Ng5aaiZeV1W8Qs3v1PexIVHqBLPen0xoE
ZH1OjO8t7JPBBEy8Uz/VXlJv3WaIDhvzsQEdx6IDtuyXdESVARzaXfYk+UQ3ZHbM
dUFQixO48XfOqWA9wLLlJVNsPyYd6BDFNIMxz+/tknBun2sGjtC+5A6Pm7S5/7Wy
XxYJvvT2qEOoe7r0l7GpR7uJ1cbvKcsg/elpIEo1RFNpjQm0AhxeCmQJzsagHCj+
8Qo/WLJPIJfSdFp+WKxgeIebr+VLk3IHoykTPW7wrRHOKYZ+ihP27XhUSHDOGVco
qMiMcL6HPzgzd5/2hA6Nbk005ZiB2V0iZiPRr4vPpQwkX44MEfj5SPSKl/sIr0U7
3R1RpoaA9nuweNC3a0AK0VTb+NczI91+Guzg94KtE0UYkXxSvMVJvXUxSPw8BZvT
nuksYU2CEl+CF2bq5ZmpktVTqoU56W1QAQFIDGnCyevJ5FTIa2fZ1v+kekCsjGNz
b56QZmClHrggov66p6xVCA4qijd8BFNbHOPlxObkwtTgxxsLrCO++cEYbqItIYfl
km+F0OgJgtbjRUZqcl40id9tfF2f5WtHGcgY3zoVvtZEzZ/WukeiySeTrBBav5cy
nQ855fbWFQIH+CJfvA7BVGa3P5/rKWsny/Igige6yAdnJFp+DP+kWSPVJRrS0dzn
oRIheNe4SeUJbbobOnCynBJhywb2LO1j1WH1FzPxHo07uUT+vkrAFXJSNs+Lb2LB
hnS92Y2wcnHq+fl1bIDC2185LhV+LOp7kxLb1tm1l0lyn2HQCfwmZmeQYCUSX3Nm
zorUGlSA/XP332vweMWEDuqjttJdvGiBtZ9gVFFG92EZVbhmQQS9lBtubaI5IcLY
4XtHYj4pBNuP0g4QFHGbXOK70q6ZWuwiTX2qIbC5vkBxLuqXN367AeAmbmEtOj4D
wDMVffRUlnfy2EZNYSCV52uZFE0Gp84N8fE1y56wRFIMn7k+URHtkASnYg32bE2Y
yo8P8b7KuwvGlvoY0kHNRgqRDR+gr87jxbGLcZhgHhnERien4PkoBwK+KRRCP8il
J0VrzTtRW/o+EFl6ex4yxLaDWOhWcdkurmacrdJLnjyrE9pUSnH/Pmi4IJX7vrpH
C7c6ByBv1hsu5wNho2in321cncRE+cpnNfso3vvZng5TOOFkCF0TA8ljQHrhdXjo
m2T/Mls5fMzEqNX4kAvXTENBMqws9872yjkKBMy6ld+v7chI4Uy2/FCd/uqAFR0I
RQGWbcxd36JRk8s31vF4XPqWn7+kEsdA9mVvj8u68Wv4u0zg4uCqW3QQ8Fo6w182
5jBU23PbdmfVbr7XcRKKVrHGaoW7vDih2QbG+50KnDslnfGGO8P6ZrGpdcVCcpLa
+q2T5h+GU5NxkEUFLhXF9jJxajzaXr9IwAs9zearbFCtBEz8WibI9bNKiGZ0u0Fj
ZDKhsLjJcj+o6tA4jvEoDvgNlCKSWSQAcbhh/oaylw6rwNgW0/WQNg97TUwZ3Ord
J42ZS3dr62dCmrMEUPCFzxm231YHaMIV2fXVehlDZ65RP97iVgS9HOF4MJeqXyGB
S64DVVyiX6W/mdhkPQS1mM9TWIOiGXBOqj0h+hvk9Q/Ve/3ZfouBL988psf4770K
zC0Mntf7kVRndLT0+wq2oOA0uQTW8haANgWSlZ8Gk7uQhJylyoU4uJ2lOMgFcVr5
D6xv+9fMF5JaLP5qrP9AlmcYRhosu+EmDwYdfUhd8lwkuuy9JbJotMKRt7mbClck
fB9AIu1WCC8acjkAaj4tSdKqn+P/pYBgH0/9WbRzaqOo07lWZ0GfbiavyYjwpd0D
GPSWECk8IMuFxYZ6Rn364YEEUbzeEFQxvqcLMElqCLsmbotNlj+xkDyVoUYsL5V6
i9tVrQiy0GKZRMKjjfIBRTRFvNRULWZPb35rah/YB3YQ8dt89SLaqwZ6zVymV2fc
SHrQrlt58qy5c+EtA6VRcOjBfb0HFu8PUZWn3pDUJbvSYRtauiWW0rwEaWJmddBN
1FyxiTaSxsLxEuHWc92GFmCi7cUxQxO6kMvaw7nHHTsgZ0DmzB/p+Pja+RyaHKrO
9d93LrwMKmGmh8qyw24t1xHzk/jZUlJXxcWbB1Qk3SueDic3q5jbRC1zyylXieZC
+2itx2IB3ZC3y6BG54Z2SsIA0yQXkJIa6sYbMEsg7iNY2LraxYSkXDy5tbBCBb2b
Gl8yiuLb2EOu9PA4Yq1eCG5wqR7P2hE8qK9BDEO649T60aTNRiDG8dKRUg4QBhg3
PDYI8/u7QTd6UynPUY3G+fwWzP0s2fySEsYG+BqQpS1PukZrIydT+CBGVGT6ntyt
6DnkBMhzVU1RNf/+xrSPwyRbQScLjY/yV+B0Dsw/L82NhPW45J75cBjdxwm+wEvv
0/T8fNGCD4LLdsG4medk9hThrjc9i9E0N15CfTvHHr33PcjPqrF7ILf5qgI1orFL
0u8XsdpmlsF8O8XWlg9iTadOf7iPWzIQxyDfRFtIgOyo2cFzg5Wo4o1jNI+xUDJr
0h5FXgWdpWakjmCYZWhvycfMfi3sQWWk9WCJbuKIOTHPgtfjx49V64wVt5Wypox2
nCzm1qKkY0TA0A0mbs93tiKml6gLTOIvL2nK6gx3q4+gYlEWDmawVBhPCoV2bV7u
fd4TGV+PmoakB1qV0cvVpqwEsFA6ZdWUyUXCr0BD30ZBox1KbmtErc0IXbE8XMsp
177/kpQDjlvYqvmYqvJIIwP+X3nW8pS2R0/OWQdyuZc1uQO3P3f8zqN5Na9S3oR0
KMil5xVS4z2llwPANw8MXNN5D2BagJVae4mzDpvgxe1FAX2iHTTGkt1gG23dnlvU
FFPOroQaF+CUhnCY2zmKe/Q6nNpLY2ZTdxl8eAFS9LJ+kArzzKZHW1rcAc2qN6nw
FbF3DyOn0xuD+izIUFVEaz9PbXa4b1wvzEtbzs5EO1RTDBJ0krr+juVChQV4RWvx
P1aCWbSc+TRcOsfAIKvscsIYU38hocnoHyXEtfjeb8gEoVrdUIbKkQW6MMRKT7wr
RxvTBGRxwCk09Gv2pE++VWoFYhPIcv5tQjmrO0BPF3u89kjd5BYA6tLPGIML5pBo
GhMYPCr5aE/A+BJPOFVwurInKdXLy2hlMnEqHAmDl2LPeHJv7DV4iBiMqQB6VSD8
tio6Qo9XCZUTunbSzXlSxtgn1yYYrHicl8YYNwzTS3L6hvKhcZOXwArZdqbSoWbG
3MoTqlNJskcmSUZjEqyfcHkfzzFdL5Y3Dk5pDmIw+SjSnE+CcPAuDCWkxOhNme65
EJRUK+GY4y9T2Ghksnu1NteGCrIDVnh5VIjkPvjTlP3vLAYHz9WRlDfupP13eQ0d
lex8Pkm9ZO5AqpiCoWE6x0yhqCQtXRBk6ElKdyas8e/AzbaA63W9ZCBgsuNEA/BE
yJGSWD2LB1163rLUBN4YWBpYvugVfdIDJ+5P+Xs/3C5orWbeOmjRmT0uddVHTSex
9SCl+wFjPcLy3hsaUXDSE79sLRqGtgHUGQSps7pVfXtXMCjD8Ov69RoM4w8oFMC4
x7XNBUC8Mn+C5u9aJCkAsXP4ELwds1XhYeCA4ODZaxZxt4SeLdNiUQ63VDn7kVcF
xFJdZQjvhk2JQ0jFnJO+xCw3xazxndzQAy/nxhp60r/qERiJQEQPBIUIT5PBzmfS
No+Ayl4JP1kulwDz3JDQWU+shzFNacvqPXSiaNC5djk/P96HbW3nAivhuOrtcFc+
QLpU6PGkpab4XWlZqHNXbVxtv6mc/uh/XrNUAyjLNCu9z8g/EjG9iCgkAPheUf9P
2+X6YbfIPMDMwLPEpBRo+vho+aKQJNytSzQfk9ppgmtIG55m50sqJRHWxPXJ9Svb
WTbF6ncwEDElJ2tfAEiLkKcgNQ8BAjokLJTKhgD75Mq9Eg4dEAH59Fh0hiqqRV53
CE7OiYwjxza6RaSsQM+Y3tEDnjyA0F10NDkK3pmVUvP7qewW5JeKKI7LObJ2fnsO
pFycQyvs8pAOrttRh8mnLL48Esjdu+EHxvNmE4DjbBlmPZJYJuAlhYupmp0Owgzj
WNd0nNhonaTN16KGBiMWEHungo6I4LPqB1N9SwhChmjt3EXOofq+1yWCmC1s2NPF
DHwpHqrTNsWRsiOldvKYb/NmD8nyCxzNSkQpxWQMN5Ufl/PSen/5ZgvcSVZnkyYm
3ODoE6m5tjKGK/eTLuvHZnpz5gTV5fmnS8pipQP468GBkSAqaGB1aQs2SzhUfewX
UYugb0dYs0PG4VoQUp1MyJ5sHCeIwTlvvqemsNzw/IP4PT0p2JFtnm6/1m1nSGg2
JN3co+ktvTbkJ+CiYE9y8KUc7oebijup6IRqTl/NfooNH80WCXn0VbvtvS86yPeV
39cSB0GxDNDD5gp6KC46D0wTUg+g7VrPwP/eJ9tvGn2W02+u5SwZ73kMR6EFAevF
HkyVz32nuD5I4Bp/koDVSIyVgDV9l5qUQIuSD46mo1HvGGyfGgw7e1g4zKq/54cx
yG8yeBdlh05dyQWFHRsfwfvclJkWsO3jkq+jt602IIIj4wXgbduf+k2od5k9d+Sf
74TD9Cyo8eo4EJg3V1cXr/sUhokVUbzolUYIUSKaMatUriJ4T3ihyxsCz7MEYtT+
Z7gCooyYC399zzpj8RzdGVLlncn/JKfwdUTvE7GWjicCYjZ9kdeOPfjB4hvQLvLk
gZOQUY1jYYCWXkoisa6ltpts4tiaJ5H4SzQQpVYWUXRmW0Zjnq5EQ5wS4YFehfUL
INdmeDKPZGq5sPbUGipBV7KLEqMP7JsLXXQLUiAt0FGCQFWfz42xePt6P2rRVaTE
XXjfwayKBb57CjSbYtFyE1OauBjotOX1a0FA7kOxPqEAWvxazhZ+w9nDoe0WFPnz
41Fn48aGfjZyQJ0EZ02wf9LSqhgCEmeKC4kQ1WtzNo/364aDxosK56sAUN4JH0ar
awAP+g+Gpruq0o9xtdRgysecXpntAaAEFLRLp6W2G6WCw3VnKfiaCAPFF0GMGKjE
tToOAMEn6fEqB8Oy2kc1hiY/ZX7KaHRkCNwOW2+b9Eii9/svhsiuFECTGseuNvPt
JlOBiOrUgtCif2xrYdzAXXYr17V9D8YK9N7Ea2Nhtburei8PzMPV/CIZQiLvlJzX
u0XJ6sK/HIv8Y9ZTOIJLQVy3fNatmWfzqkFhXdE3UxehnIvGZ8GJakkU2VY3KZkz
Z5EI8l1qAV8aG+pnEhZDwZkkI3YP/7P+gawfMfF+AAq0KSNmewr4QHMy77JOWAam
KTrACOmrg3592MWwJ2QCJe6VcDNiJJoRWAwsLCJCojja8Ryv+vbiLbH60dl9gvpc
lbfyVBI+C5TtoRJtClOp29SAoN792JJfWg7aOZ3lSg3JnO6jfzc810hlTRcPgWQp
U69vi4O/gfZdaHcr9JP0LAexsgB2oQuZEgSg6zlQew+a8F1o2KNQ1dBmvAwLGfnR
5cgK5eN1T5XrqeXtx8ZUEIvBbLU6oJVEi5QU5yd071SEHANIiUE1BeY6mRPu/QR8
S+73q3r5Ilo3wBQH8HPWu1Hou/RKYyNwV8uINvacQqGEBelBN9JOKUpr1fLPCXNy
p9zGeLWuUX8De7yofzB3uYCHkTFcicQzFWy6/QBIzWHM+kygY5YQ4ZKTlwu9fwaN
7IXMNMEOoMh49j4GRDqlbNtl3JyZWFIquEgfA98dGrrbqrrqCKPxr/HoHQC5/Z1i
DqfR0gnJukrGGJR9YGFyKRR7xGspJUH2diQZ9ebMne1Opn9GOnfByHxIl06nZinV
GkfP1AQYqkY+hHkV544q/62LC3DTTOzXLDGizsa9JHqOLADuSAFEvpO0LqnZHxkD
P+OEKS1owiBDaYeQ9A5JIHChkkfO6hCeuKa9B14ywG89hpvMydRpgTWA4j6RD0RY
CsNal7nq0ueF+ZDMnlcRR/dSYKxsh2LQYa/T/ZUMl+zKVmAJ9rEj5x0gZFNtNsE4
qLojdOriYW66tuD9RdHRtho+TwwA9fe5pymH5r80t2PUfiMATKkRgKxqnH5zfYlP
p0p0KZzcXoO+7gXpQQhj0PiegOjKk1hGuqOfITgN9hBvbJmR5ZMko6ENuU506Obg
jG/tH7Ex1ZAwuiwSUsDswxu5bTIcmXJ+Euxt93cOWG7fv3KVz7CHw83a+UpJ866b
8J5QFW5fDXlj/XFUkmBsJJX2CNN4HCtxcpqK26WPbPleBhDamvwfFiC4yh6nPPEd
bVWoAaNgeT0BaY8uP9Jy5pJk5SxiKp87D2c4t29sLAuONAPawjsfYMTjXPry0QJW
XBzECEuDF+7XkXrCGHBSZO88zEZwrgwN3koELavJAv/dI1p0yQX+gqVBx7uGxWmy
t7z/pAPSen27FydL1MUmHmr/RkVftw22IwWjMzCcZjTwj7+gRPu/ksxnh6Qo550J
JC18kuzxkz087B40mifhbjrDdBPbPxjRHrtT+ikJUiKwslDsv93TnwCrnpx9AIpa
yur1wtEA0CLCGYASfImg+nQXrYX1g/9zc+qgJGEngRnNLlxnSTEIjtML9Ai4E9so
cMgb55k09MXWGlXzp01vfMmJE8m5EMTdNbsEj8Ws/HiR/E6CgiomeDbHzsLxKjjo
/C8gQtftWBJdD5yDh0S/EMPZyS7QG9qAY5tEHgL5LvGtZ0xsLNtYLgeVF9036kzJ
W8ojuGbMtOJwSburxHzARKTj05/qm2RtZWzPWMApgu4i1yBd2jgP3hxfZ23dohsx
GnwexuHCPj37gWAdIpJNEbJ1gRIi7bsltoRxFCB91Wtqm0Y4ZKE4MV9u4pcON5ss
HUoqwovEzRU6YFMulOuwEvye2ttBKqOfNTQDHxzCjOpPwq0OwPTSOY0iSKdXIvEi
0ZFtjQse/DCAZCWYomWIXgN4MMcBugnvIVtMcYSdqGQKnSBy7wVYocax0JnED3gq
IXMMdQWw0uXDU4Vt7204kWz7zZ9Fc9G0K/hR15aLXvJdhvMb2sIv/v4vEyx8Rs3L
GUv1QJLwQT/BToRtWx5p+ZhJ0HdpTkVnxvUNhYnq7FJodrWN8jTEhfEYu4vLSMPJ
FHWHjg1RbO2qcLL/eOcIzbPsCoHIYcblASzqse1dojJrWVC3vv1jYnotGw/PkfZW
8rxb3RE15WgTqxjXdhA/vzMXCGGc+kQ8S5r3lfeAiq1yIsX+qgN00PLvRHNFLl9n
8Ep2/+tdPBciEYfRyM9gkIuQHemffA8t+r4YjhXKZG7kfsvYsPGRtQOd4z0+u9u4
XD8jUHZtu+Sy94dGFDwkyr2F3PfagQfshm1gVssn2mdfFZ36X1YnfkzUmzpw/NMp
AmJhCd2OzCr/JL8EIBFX6krV6J0RJsslg+w6YT2IWQGvRxZ3ASIRBhIjOXOayNwF
7XGqmRTDmroMFbZcqIyogLhRTGjUN8eT8r/KEwkTpn4pWaY7gPvizwaF3eh/lC4/
SfHBTiZGxT3q2B3I4oL5WAgRIOl1TwXzUq+Nc2HT/QzNkFJ5t6ZeFOrQn828iWVe
wxUBgvMiQyonOp/GSV4Rd2kZzf22sAtFRXm56ojp4ugQptwa3A/5Ymui/Zzp1Fcc
BovTQFtTT2qyTMVgflur0ERNYYK1kG4icSwHKKAd3QTOS+Dd/nIovyI7kK8++tdx
4IdrUuvTJPQd4Q9+cTVjjVPbsgzi8ipMCnUsqeP+HPOT+9xzKiK09LvBfuX3ceH6
J6y6Yg8IP1CCD/vrEhKCJ2vyu8BiLc004vQZsEhVzOZZaJbmxkH5JNv+vIIPT1VX
REYDYjij1fGXl7xsXsaShA0PhW1hS8puToWX2gj1uJu8lSSyKBwEyG6xBhvLJo24
nbwowFCq3L3kafbJYbcQVnZBg/mkWytxjgRMCj3OyCnPoLW/jTJBwfHaEMc5hWuo
KIcRrj4EVmQLrRg4Ud9jUUElORugENLj319nHk5zDnUm+GI57GHslvjWj+SwZBHg
CI1ygH2gusxK48IzObt/Liv50VIHWyqpy5MF36ILoEuuEfm6bTWpNfdX+3JqMyAg
BX4PkMIxfq1AHzDoiJWhxD0vs8UXGn9Z6en+1SwkLW2rFsRyUfA9cogSRIyRBt1G
i5/u2b1PO5aiAGBfQhRjA+6ll9oP3p4yGCUZx239bH8RSS+arc/mCxg2F0B3miSS
iBq63flXghJlRuHbY1H6y/KkJzCuLgu8mkjgpVPtEbSjO8zkaPhfIbIov9sC/mEF
RW/qZjJR+e2r19VRA73I0sFlKNtKbn0ivw4RWOHoAjKLvuvDX8xq4IpZUwCrHu03
vBFDlXbIntsdo/D+hh/ErevpxO8/soUrGPOZV/NntrxC9hgO51b5lW59AB9lDSdJ
C++h/BhLU8JQj2UZ3zPsOPAKTN2prWDefsuFkDlbWWzJYF86oDwAHPa0yebbqmVH
JExNV4IFWpXng0Y7ZuS1dDEw126C7NEKD+biE8dk32+gG38wT+1Psem/7SLdAKcC
PZ77IG8wzCzBBgXuHnxya96YdT1i9U5pVw98mDvD2Nkme94RHhWdLWoGfU9t/A49
GHMapTSR+harSeI8vO6TKBDWWjnUOkhqNP+bgBAU6XYfRFQjGU6Y5lj58/WN3nNo
hm9RWgk3GHl6UXr3Kt41UdJpxWFTJLAJfRVcnZf7/wBNC5IfyXL1jIB6KSwPKGGx
hbx4uX6X5LXAJuzBey37Y3mmlSPNCiaNynHYJY9VtzPWR99jXOjlLzbh7UjvnQH8
F+CoqnDjeaPIDX4O3RO6ZdYUEZyzl//hIkTu9R8zlKDblmaLH9zmFWPaxvXa/Txj
Y9Cji4um0qSqdNkHg0NH6+CHC6HsBC1oTzo2SAGaOu16doppHXnrzic6g7i2PjL7
htgGRFJ3I/sJwjRFa9wXZaPdcf/fmZLnbyrIGO5+loBNesApLHe2a8QFoX5E3sH6
rZ2dWHSahxMimMKWFzLIBW15Eyvh5gaA91MmkLbst2kEMVZd5tEZ+Z4VNLWnTkQ2
xjrQ7pQE9BuigDr+BufPp82JpKP8dTh+hwFhFS126YQwnlXuP+OtfV3B5I8RnEGK
nDae9yrSy5oYUi6Sn7pPXbcb3+DBqEBJZEwp9GqLjmopvSX5FYIVcxepS4ecsjfi
akCU5bTAPJ4k0EnMIY28tqW5Rw3ChbQlxc939GZym1NwGMsWwuj25bTgcCvE88lN
nYehXHxjnhpdDrqnDhzHpiN2Xsl9I4z9XY+xamo0ZxDM2bZb1YbZv9wXHWsVStiZ
G8VZUI4IKHuCbRHD6rRp2v4CbE8ATu/sQFM5dKdtwXHsJv+YcvSSyWMg6vJLUGlz
IIHZTMQbnqp0R4K12AylQdE7CPz8IbYIpJMvltyT8VgRmg+hJSj0ESA/S34gbqd8
B9WyiI2GmmtKBZ7Fy4nALBDyLM/uZu5jlqtFNvTKhaEzFljFzJwosNEo3GxO1jPC
d3lP0qbItNk0PdYwlNN1vIgTDQ8ELBZt+Hbr0ScLT58KNq7LvW4Qe7aKhDl0p/2X
xjwg4jFw3X9o4HIlsy6UkBbmU5tGNHpcKsn5ZsgSrp9ZR2Y4LvMwhUdhoo4+h3jU
XleFKdRWCFR0ZG0KYztMsVFuAOntpdEX9CBoxwsdT4N6TfICz+rGrTTrERtG3/ot
IRleT9x4ZU+zhSCMhR4Tb6R65XKMIUlheOiKZEStPjMNFiK/9SMajTWMHgLX7uuz
h0eaAkeaTvU6eGUMIylrD+w/q/Xp/f6PKJaOVeJEB4Hbja8uO/fsykMmBbeWHyPb
oFBDknlPsq8QMornXkLeBQDQMPgR8IJ8G2P8SjemD/iSKGLL8yoLzPbqrEKhJa09
w8XWzn94EPtcNVl5PYl0njrV3211zNZRcCCEitRChdUycz2sNS4ZwzaVIZjIBbXv
BeWi1iL5Mu2jJoyDw5sD+YMntcEI70lVO6caIREvZyfPTV58web+vyAE1M30/47p
2Tjd9qaYvIE3TI2xE4JtUYU1/HxMYBhZIJB8ixXw5RRNNn/svIPVObbADiAhkx2E
mxQGyb+MqQQXWb7WsQ7sXTkfiDEBgn0xW2oOF/m6evmI277EqBStx03Y5CbU62i5
J97VJbQKmbPlLARMZgFQmZaic860ffDe7vdm2HGFlcLGQ483YkiFbIocjGgiqzg6
E4pGjPLnZR9/HrUlTTTnIjyN+7CQ+9s5Tb52e/lJz812F0i4jf9XjInrlbIrkxRK
4gXgeJU7Q6oHyd8qTw7wFy9gBA1Y/lAPe1pN2g4WqAIpiBf8h1XHUAgYWfHpzN/f
oKygnbnIVoV5Pu842fmbJQu2IxUV8D6UhJbb+APFWqwLkbljBiEAMHYKGUTETErq
RbDOvgrAZc0OUyWeJJOhtJaA7RGthiCuTlVfsuZDzebIEZZ6J+YrD9k1z6oRmSvt
/vqcppOBU3ZUqp3qlJuL6pjgIWHVdO+89Ob10DB45ut+ta4lF9fP6fld0FD8RL7n
fBl0ksXJlrSQ8QCyCAdrJKGMTQD+y0fkT5w5C3pVLbYHGNLCuOvdqUklH32MROEU
3C8yPEox9563VKbXX6KIoslh18kqICSLULv/+5+UuYyM7am6zHqJ1YR8cI7uQ2r8
qOAGnnRz8GZ7n1bX74R2wnLVGqDADihtX1i4YQmanhDE8uAPYG2GreGjP3k26AIz
7sO6vwv9OIDrTOV7WaDgSX9XTsszPQnEUnuHLKWwGmA2C1kGUI1D16RpZ6/275KC
TJBhWu2yesxwfM74DK8uZMaKOy8Ogga1DfrjQh7tSOzv+mOI6nIYapoeZ0TL4kPV
qtUJl9cNkryYKByGVlKp54RtMUif+NelLaV2/2FghiuVfUkQWT+lHNaGCYPabIf4
vuGJy6TyyoQon/4NZeUdTnTryCHzeZmN0MRKfQVF4x+Akf2/QfxLyik9bEIF2glX
QXi8MlodpfnIqJdPfHRx6Ek+vUvMCM1NuWdXOzdBlclDlsVbcg+Fq2PaD8QdGxxz
WSI7kUxxazlRcbBOSjf5ckrDb+gLirlmrgXn3r2iBT2NKL/D8PLMJ3S4KXBuie3V
5MbHB12Oc0Ny88YMcUY+wep2MEiEWsTGmo7X3QQesaeErd6JtMH2tQmdnwV10poR
lQOiKNuczIq6Q+3ELk824cNe1nGXguhfzYiuXH504UzT7CiQsxarar7mklQraDqL
l2jdRPgNI92RJtxlEApsv5hkOBylbkqOfGhy2hI/6IRvaWn2IYWD95WokMgKWIP5
0cvj3ai2qj+PRJLpzVBVRbVqukAVaHNPdlqkUkWhVAVqsyMyAJI4Q48yl892Nfkg
94e0jS6jraIT6JPlbnCYLr9mnldUet/atuqf2o/LKXrwVFd1cmkrgFerR/oFyPCy
zxwHWUiTZAqExTGkgmtmA6NOOB79y4/flcenTWTphfKPLzZUs5h9Q1pyo0LIUgFj
3iYD3MHnN9BgA6czibiBj61H0WULTnf2kEVXd/0nrqDz6HG/MLuArxHk3km/kn/e
TAlkeNbRhU97EB2CDKvq5x4s2+BL6d1jQNI2oyd1/J6nA92/CUAH3XMVHLFJVPxk
c2gFOD+zPGqWXfMN654O3kgvUp6V99RPL+NRDiJrrSassuI2BxcLIuJVmSJYrDc/
mcZbIDpB7PspYz3tQPSYyK2RVFCX7DZwPgW2T5OTFPhVjw90o+Dc3T6a1HqglfBZ
K/3vxF6jofkHO73Qj0AXN8mr6hds+BRxl8Qh5IH6gWetuHaq+zzrCTDRJG4+BGbn
jbKvoFd8b82ErugMqOf6ivy6mz1zIGe+BfHtjLVRtkdEKumS0vzquqZjxxfio3w8
2K1KG8DHE3M+7lnS1jNMjnYQZpKm5Vd98iFf83YlGrvMvrfZbGOLbAQ38NuNusOb
hJtfVgIU9hwu4VlFSRa4Yi0S+znU2Y2QHA/mrW+5svj2gGgx1lekS4OBDUg4/rku
1BRnORQsD8CBRY8JRM6f0x1RHMHt0u+O1OaFHH3jHcxW69+a21GPqaRiCtTqXepQ
ZHHk5nb/M75RXIII5/7/ki79vctW01m3BZ8kS71+q4I/o2f+Co0OgTcN8KfFEQnh
0aZCLLilS+Gq8YymEex64r9g5nBVxSwoLkse9ZKyfRzuSkYy2Rr6BbPrkf+tjqBz
b/G7RN6IcJxAvmqj0UJTxdzADlVMMIgntFCLVTq/MJ5UFulhWdCHFC3wA/gpAwOP
5yH6tR/QIe74vtiuGdmjl7uV2jC+Jepf2+mXUf1iaC0vSTho0NWDaUxUDDtuKok1
Rj6FgirI2fxobCUH6P1JfKPYDbfYSZhY68lsFURwPBQS5cFWe5bYqyvbVM5WUvOq
bz/uq81ZHgZHp03jBYRcL9qytgU3gXMn3sT//IIU7EXrPTp+oghm0No03syfJl9U
cDi8Zb8SUtQMQGa5+rkTv32MHMt3hVra+5zgOPyhBWFTJbFPieVTZtrb65Nq9nVj
Lg6XwtBrwtvQuqGr6ZRnH27O4bk6S2vX28ZznGv+FHfhoHr++yHzuCj/1OBE7nD7
JFoE2dFAwEa/V9jyA4HLrGkzl0RGkzev0g38vd9i06rQ2JxK7GkGMkkcQ3Y/ow52
kudkGzQiXCt+7dOSixXhnJe8G7F+KK6S3XM8AnUVDhjg3ThXSx/qbTaXeTR3MQh4
pC71lB3qafeHhx1deRWJt8Mq1UGdaAmoLV4t67Bz2gmwDYU7vQ276EoNcRFAiWlH
+nEPXGqTzz+TybrlsTiIF+dHnQ2UcPycXFLC0fQBmsjXptonLuhHCsxLcxMqvl+B
8Ti4YCc2muFZBLsBYAaDLo9J9DtST0HxgDv1gH2+TwkdYZ0KLhO73fTYcR+hzJvQ
YAjXrtW9FId+sF3O8ucUNPLSRjjkKCpnQ+3zElRUlB2U/6iDeIl2EHPwhoSf2k6W
j+8Gv5SaKL5C8Yod9GOf7ZpF6sENgFbnU6FRLRTPs7fjFBeGxplhhb2hF4y3lR7u
yWtGQfKymEKnKQ4lLCXWL5z81tjqU1nP9CCN3PwyYqnIosXXPw1bxvxPB2ycsAJO
COmjZucvC+fnH+y6/GowmP+1Q/L+0fcYPfH2n5wYt9seFNEINe6Qe11mZ0O3MTNz
+nTnuJvSeaf+gNYi51DhL3EO5o3Urvb85jKtAx/lL2fTgUbSBxLeNm9xBrpohkmF
gW2q44xt8y8lM7l5Jhsa9NuzOwR1uAgZO9o3R2TYbJDeV62xDQPTfBTrXALgy1FL
SiW64kfg+oGjKV5b9uUrs2laHJy8fdYL6s11DpRmE3PiDbI6qyuxvgjgQvW3dXDB
f2QpXWXekSL5SwLe2gJo/K8zH5mZyaWcXtK5dODI3TBNuMhepFM/WfbSkyI3hxrr
CoOgvAimxMjq1Eu/ca+zL47NuaYmPWp8EUs2XybdGDA8d21J2uGyMKQKl2USdELX
mhF4vw4PWNtSW3dvVwhWZvlTq3CLM9vfF2ay9pO3vPU3J0t04ZtUclqjFsaqrDYR
ob5FDzPEN93Kk4ZNsc+Q3Iqt/ucPMm523KHjD3vXuYTTN5SPPdKy/QSicFUbqV3g
d2ReZ/oFcQ/QxfPodUUECczw1J8q/BICd84KNq6Llzn4+4JicATBvbAFP6pxBOO5
cxshPu35v5lDPS22XsLPyctfrt8d5hz0ENaQ2DzE4B1w0zZs8watfGdExqLHEZPI
0zbAB1ZXQWYNAyL3QQ+d/itXfzdn3HvKBfpKU9yltlOoLT91vtktJkUioARd5xnk
/8esUMod3xwp7Mqq03ujEQF6oz8H2O2GuhnJT1PvQT3i4YKdXG8hlXM4Qi+xzCc3
YDFa+0I29m4NV4tMAGO3VO+wI9gs+PMTF+bPediYvmVvEv4GTPQ4T7D2lbov2L6e
1PYh81ugKDJEBE8qIXNnIJYhZEXzuyMG8MEyKF9VBcHGQo53MKO5khVtluRaKyO8
M+HdVinOOOdNjq3mHB/gzZo2MTUwX7FUdGWdDcp9gvIXAXkh+MdQ0PU8G4XumOtP
Kul80oI8K42fRbSMLnAmy5AoeaSqsHDuI3RWOKgRitfKsyKvK9kk/aL26QyBHlt1
Qq4I1IVdF0lyoV5sRenS2xNf6hhFd+DG/RJuwFD5PTQZm679OUnzw3+WKWpztsyH
lCzGFi2c2iud/f9EFYePfUckHCcy2hsovH4+Y3vIQH4B1xcP3mhJyMOGKZZ+LgG8
Oun6zsWV9saK/qk2rzYDIJX4pibJfjLDkw9ZVL1EZjXog/8Du31IWshmrSAyE+1W
2T4LlGg1lGVqXBUdjEH54r09tQ66K1/OC6oBR7OpSjnCwaGWuINLUwSqeXYkhhO7
LrjhttcNMy6uD31t154qYx18trX4K/dAgIA9Kro06PkvKWvbv/x/UX7HwXx+DKw3
oK33wOUaQBDxvHfQ+oFcS7jLqFja1OWVFRVu6FZoDNkL0KmdaiHQ8Pp6nvaV9AYt
3TEToEz2dyhKAHlHS7Lc5YG9VHbhiWi0VLtBycvefAhvsmw5Qg6g3NZJ/8zuMwzB
trSrmpcb+8GBGdu8BMjEbubnLrp5C/x/j7Rp4UH3FRqy2INmDo+91oNffaLnNpfw
C/ixu7TwPK6RSjmwo6RxNrxalba62FY2AzUmDkMC2y+ydcrLti1SoTs8kKqqZw2d
P4jBH0h9h86/DVcJD1UIt7y7KwuKufiDDl9/neT0AORAZYj5/L/WFkC1YUBqbIRO
7Wo4ybla1v0nCRodW26h+pyl8JiVGdkd2s7hrOC5rSqsCBw7nkqKM8iv4TvRJpnN
I6gQUZktrg+K9GUsq0CpgFlFQF/MBGgKYK0hwDLWHvvTObNB4gQoGbdXK9O947vo
1d2tOlZb8FOtM8MugoHaeoh6Em5u+DyPojxT9wqZE7W/GsWfLQvyIzrXv61c7zUB
cx9qBVXIKBQMfEpdtdOyGFCXLJDdCa6rERhYuUidCp4ljXJptUhwXnX6N1CORJq/
skIBQ7HeFBJvV/PRYjJ9lHAzExkUQbyP7z/O7Al6FlooORXazKRvqO4C4Tpl0FyT
FYi7ZIEvNRqFOxu8hl+iggvQfx25eFM01oDOW21CUzwaPv9rVag+C3NSY7tzCAnn
/iLXxMQQqWHrZEyeX+aME1mhs6pryusrh0Sh3zBpbcswXkPvBg94CmySMC3rMtL4
NxpY4YEGSVyayxUMkZFOf60jLxxhrTJqJLhU+83Eb+K1IrWpHrUv9BTIj/fWmSAu
ybBSZhMMSnWaK8JSsZ4z93j2rkjAFoBafPTPfwkG1KJjUCUzJVBB5d5ydUNXB+1k
xWAZiFAdb3S/otuqertblI0Xoh2IvMnT+5gcQIWewsJY/UZQphKFnGa5nHV6XBvL
4nI19r927E1XW+fFmZW+JztdYZRcCCNbcONpSxJsQHm2+bmUOHdH8ZbXwE6Tb56i
HQShJa+K39LWg9iX0xmg2Ju6T3k5EtH5O/PA70lJg0GZB7e3NdNZ02GhmpLV8Rfn
H6PTGfxez1VA1qxDRW7hUJljvlBrAp5KAZB93L51GF/Buq1baEZd5+rDuvYvLoWj
aHl9unXVmD6VMk0uZ4+vm1RKWi2KX++p5ydrJ+ANBprpFHCbckAztgTAgxB1pOpb
kLLaLdEQ0MUdimYXZdlCVdF5farjuyWOp0x6dcXMA47aeCe56lZSvpkbIAxRt7IY
d2uZZTJ9GZKfBwqm1f9Cuyo3Uk08hcnh89FLaKOidhhhopei+zp/79gmUonKULlQ
ualQx4QEKfZtPC6/tnIDIMy6PL1FgP4xbA0dq2YT8CKtH53wV3j5bFwmSiWKSBWx
dukxPbBXTGObynp6p4d2TkFRwRwoFObByiVJUnr3kK3Q1Nb1KdMTJSus7xzYPlbg
WVTCnCNY0Cyhp+W79Et4qSMKMAtBGei1pbsVE9ASikm2A/BYc72sJfyz4uGL2/EF
MKcDiaAniPucoZRB9tfY9sWaLsWuwe/tdOR2ZoiRsyFxU0ocoPhME2gbia0aJ2tE
jfLwVgsloMRyU99ZByxgwByt4P49aofgD4+NwJkvyPrblewO/A+9v4atgfp0YGs3
SJrOxaHn/MaVcPXw5bSIcPZa/QR+rLT1lnwqE9OlCfgvb9BUr3ubr4ygKbauggbi
2Lfe3NvhaCZdtnzCBaEZP2PY+DZLmclQ6jf6iC9cnfCzFj8oyMePtsm34z+QvE+g
GimyDnnFQAKe9lXyxvMdIDWT0lR49Ai49gRnTxy8sXEZ/b/LI7l2TddWMhRkckEW
ZsE7i6IFBVJweIFmPs01C3aQj2xOt67DozPbBBU+5oy4G6N+HvsDSNCVKioqQRcM
nT3ib4iZsNnSyFwgwru+5RFFVP1j6Lax8MnZac6S6bj3Q5OvTNiqqCMY/1cqeCvd
HQj5rXst7QjLKPvdWJxlr8p/b76BzadrKtDdWU+9qNJayDkMpq0T3boslru37mtQ
77ok6eSYb8RN05UvGjY3n9pmAxRMg4UaxEayra2XFJYcOt5lYysTL+wrgfhQBHFG
QIVN7NqKoDMNJVplL++hBbqKlnDyJHX/gijSUQJnGTQcMasCN9EZUZ+KGNvD67Kp
eMHlBamUDbG+2grUO/oKqXB99SBtH6jf2hhAj6FHcSmaTjBb3qUyOpH/LFPDLdGP
J+GkBRFCjeei/6NDq33jU9N9J/pLtYkWNpHEjqnaR0kX9icTOJDlbvAGYCK/YAjD
ShW7uLfDkRq8b2MAdjiQAW+dReStX3JTm5iiHJgShSpEU1KYbfFoKjDvq+K30fSO
6WBa9ss+av/GD4GjnzYXQ94UuDm2ApcA4yLjpEbQf6XYcG6a4jSNWyqx3Ids4vtw
9l4fJ+8HBJRGf4g2oWCUw4lux7eaBChnb/WcUgzXRJDhag838S/IVK9Aen6NG7xC
jEz62ee+Mtn6BeYJlph5fXAAwEcuzK1FY+15jhiBMc3y+2xHrS1+qSolZLT8efof
I7XxZt+VpXasWnWAwGJxDCEUSyynqzJLrpBPlfZ+1jnRLs2ObBvUwODVQTiPxNRc
pQYeb5ZsYcL3SGYr7kVRk96W634Mal2naQBWl8Bv9Ak2HT5p9/fS3VdABKXA61oL
tfWZoeYY9ylsUUoGVU1eQ0O2k+yIYtfCyeJvyc2W3V3EfIHhex5OoQo5SNG9wCcA
IN0G0FrnludEjHDcgpsHmkrwYEGS2HHBhQU3kxUR01Jz5dYvuToofCMSRqPJ6Dgs
K9C9rdZY6CLBUlPGoGj6qgGrDM0lysxOmWXl2JmImV9sS9oiy/5rXEktCIdR85c+
qihjgW63CGvdIJOFJvQs8Jmu1BaHJKSr9YZbm1AOpPrfESZuTPjLhdGkODeMYpUR
yFNqDIRh1DoOb12YkJhtGP6XxOJdUL79T30JgtB3oiWgXHJPl/JmzzqJmhUGqsHt
r+5xFWllwQeitUVanI580XVeY2lC9ZVXTvSkE+DTUhQTqDr/D9emHHgoaoxTknWm
0yQBP/ms0j/ia3A52KlCMIbLzyNW0vlNgVBWt2hURfJttFDphZIAXaJYgZE3FMs2
SvBDJHM64pvU5p5oMBgvG06HVX49fUUx9+mghEP+CPasRnzcmUNR4mu6AxtjWg6j
TZye34Tr7k1VPqqXXRIRJWls+AI89eG9SGNygtwEBtsicpLdvPz7gsvclpl8l8r7
BEupxwzRmnAudnqcoQFXyPYj9IS8zm88PSGwYwQ+3sXFkyNhlI8t+M8gqQKg2RQG
ZYhCa8v4L6zx31ih/2/ZPuz7XH9VRqiCmmCXj89uI7QuJQA4SgfONY9rWTVc22p/
LmiA7elofW9f7ce9TfObluM8sA/XIl/fD9FL+kgAnnZK01Xf3qN7CnsUvFvWaVX3
ut0f2t7z3YoBGfX2ccR92N8Hy9nH/+/hGGvttb8Rc9lmRRKMBMiJN2A6HBAG8hHI
tKQFkZJaKgPdhQezty7g+eW4o77VeTAc1SdXNQKQjZv6GOFTYRbBeD22pPQApUqJ
uecSTgH1n61288eb1fUQujQTs2pfHv6EVoZ7MRBpMX+l46SBD241Fka6K4MYAcDo
5qCiH3DQ3OSrrsSRzeDbaAl89wYQthyKqDAa9JyyzC8JMuczju3oO2orhLXAAIiM
/u07aaN3fcpWuKdL60nOPhjO07bM0g82O6iAl/sEpjsXL1H+sntTx5Ow+4oPGi9x
h6HZZcYyj4n5ElYZMZNM3/1X3u5p0Ooxr2iIgaEUCKw4YcM6wnsoBBFhrXmf5oti
ZZMzWdunfGOs97pZvAGd5r9BuHbJtHHw8F3uE60RrIU9Opfa/+VLcGm723Ty9D3K
U6HLVQCbdhHlIJ/VppzzV+s6uVPkJX9rs9pEhEBOl7xcVZ9OggjhJ/VUdfvlZrA9
h2MhfOKd3XTifytELY79HgeqVFBETxJ57QGA3kxqrSAbMJ0zAiGFguppCXr2kBSj
onQ7uieL20DL7WG7Osgn32VktE49BdZUHmuKQaz5d8OC4mPB4kP/60G6PnQlozev
/HefbnHu00yTsRXNRXiyvdiqiMYKH7GqK294x70NqPEMROzVi1ibYVqeHRd5pp7W
B3oN7owROxJ4Cqr0Gl25CJKlQHZzO5nWkm3H8KuqqdPeO//4ljHG9dr3OHo1uoot
qx4e9nYO1e5tVJH2bN+s/P+1kTwa1zXpbzlhJy5Jo58FY0oR83eCyzh3OeG5+acu
Hr1zH2Ffcd2kogYM/xQ8YocvtOg9Tw1+4ytcAZYkx3FVmkcHwKcoDl00dWmsgiel
JDKIlyZ8225oGxuSOaIVSvdZrpFaX2ifsrLXsmQ+2Vv3IrC9iHOsF8Xb6QJJDuQk
bQ3KUivtgXTIouxy3BnXUScewE6uRfPa3XklVt5Lwsp75gJEN92zM6soI0n7lRds
U4BhrAtK2civaEXO/CnNTq2KvQnf388skcaV31oQdF3PkiPGbuN5JhsXN6OO7WNi
eFHw+MiKnSLmqY7upEQNuh2SsahbilOavIXnHyw/dCC/O2h7rGwMFlSN8f7ud9Er
sGLYc9jDLnrN75gP6SSEpUhQKtpypog2dyyBDwwstzzpZQ3ReNs+sU/eAUIgNTvj
mBPa8gugDrCUQy37tR00k7RyjV2EHUVR7xH7PA80lNXgs959XGk7uBWuMcsCTQjv
M4pkWCg9bEbOGbBK/haQ4xP/3+jAVJbTRB4ReevHD7Et1MSfhGvEzuVIcJaM53yh
AKTs4Q7aNn9dUS7wgHyWBBTr68OKgsJSvTomXX/ReQpAqt1rAuxmXJYF8yCkFMpN
Er27XtJatsrSOh3SJnzUF2ICp4ZT+k+WI/9wAUr9ZhHiBmoJi5hjQcQI7JOlKGhG
BskoiVb4lsudG6dFl+xZ3AwEJKkGkMJu8cp/7mMjXgO1yt3D8BO5svjFHWZIYsH3
Z+ZKoJJhRyD0EPuIpgAKU9vdBSRTmPcKdIYu8uQHcxSrBGY7iunSMkH03NRx2Yqw
4wvN2CG+kEkG3JlyI9KIEdL2fie6yrNqxaLPD+gAI9YKKV0krgUO1djS40SWsnKV
d8ot1yMvimIOyaBPiXAvizZ1wxSyVxGXR/kBFgA7A2eEyLIJeu6MLf1LKZRbYOh6
7ms2JevV3XrHXZbWS2nRxcl8G5q6zksvqCqiWFnImxDvd5RbRzRClemOsVQ/yLMi
4mQci3HlGnBp4AMGY4eIzc4/HMxtLb9aTBVFTsL4CfVUvRWGSdCOLQ8t5gJeUpEw
AreU9FvL9AnU+mmR7CNyVauCPVCouX7W9U3b3gze2if0JNcadw0ky0epRHFyuSaQ
GpW+Jg55hHqo1L4sbsAf1/bt86CUa9U7sZwo4ML8cCpybNnt79Xr/LOhIs3ZFrHy
t5zJMzTD03EgOfFDHO7wM4GawpNaCmTMVH45T+Q/weVcJWc2zUSELyCZIyf36VNy
aFTNVv/Etv6bc6WyER98Z1L/zjqAoLz1EQEKIE/FtbfPQqJRiAo+OItcnKdMx/lY
y5KxADWbqxMAqhinZOoSZ4Ic0YDy3DEbTQ1F7XOvljtl7N0+wAk+S3/r0bUc1NAy
vbpe+j0dV2oSe5GBYPZcax8L5AQEjEp/njstuLJXLUJK+lthRVxWY83LjPSSsrMH
4e+EwnWJR4LAz26Ju9kEPeUXOi51i/pvA0Jel+xNg0pKc8eTS0ggVcTSK9qvXjwe
5SdsuA+SRXtb1SUU4ntQxhn2xETchCOds3aDPRaOpUJTOdXzQJ3fiMKRki1mtiMM
dbvXdypF852jCU2uQCwSn9EUg6qQouHxlbcF1kw3S4kcqQVJz5qFHTvBf0GkXQkO
Z4YvwB/vwPv5133S95DFoHRvtgRiwaonf8/46RUGmoXJK6ZoHh4sY9wjhiXOPBZf
UDQir62aJOULGCo5dRKiS2sLYXoF1N+QKCnI4/BP2MsNcGJk8K8HNBYAih/iH6ac
hcAlJOZAHFy9Xe2HThwsWYlNuXZJPL/QTWVfBim8CcVWEhtfLXa+sXePNjHAEgCP
SoV2yUA2jomhc7k8utfr1uqfixvaE1lnZ6SqDFhve/IvXIFGAscBJrwNDPHMd/zb
DjbGytA/fRnqrRamY8b3+miqvE7DrIHjpYOpmU9JbRAcjHcAqRPtgaeAwGiV4RNd
6EnwiwnZIVoY0X7TKxmhEZJrp910lvjy1atkd+R/SVD4xJn6+iJTtqSTjNON2io7
RSWcduPSmA2ATBPSWmrMRLnvCusDdZtkAs0hDdT9B8n7RORWgk1PFNU8XKy4aOh2
ohyNJ/LDvzeVZUJkoHx9XM6gvlNGDLsL74SZ0QYlfJNOU6r1qjdsTyHh9bQ2jBll
arcWz/uO/pFQ6Psd0yrc5TQvx7Y9TKyVXBYzlo3Kk3rsml70Tr1u/Xu9J2SyaBuJ
ONT+QHXHR4iNeV4GgrbkFwb7/Lj1a5pcffOs7KHnRr3x7kpay0hwDie1ouRRfEH/
X4nsxy8zYJBnZD+HKDUbSZfEfbdMLowJYc7Nbm49JGsmz53hv+8WEcQ4jxE+/nM/
lXtSmRmdwbSkg6qUDTLRYYMqmpMy3QkqEi+F7ilOQatFuX58fABlFQwPFh65G3Ej
jAWemDkGkKogc+E5X+chC8IobM2FFr8KQCIh+XCsmSYL1mOSkq6RZnBk0Gt5LDS9
YZwBu2c7K5AvNOacyvM3Iy24ZAxNmsOn+hxRdV5va2TwTexLCobQHdBwx/bp6rum
duQLa2NR1iNGZv+ZLRyvdIvgbvrGZy25q/thNqW4LIQ0km7oQthLmcQQU4opcEsk
Xy94IhLMIZisx0A1nv44CzxXpG5PIA+qF0kAdWn6LImKJYwPAQ3c2xwO5tUAzHZV
ZU1Y80Z9jZkZHoBA0kGTRuTWsFf8J2KRSb/ZCbTmh14aB+3Q6kLEYpJ7NHUeXkAO
6qeZa+fNuqukJHf53+FW6FH8AS4bcsBeGmz59xh926TgLx21FfN4kTho9Xub0ey9
kunui99kfSbHPfXAiiSawAXf4ct7EYQSrCmiEGzWb1VYLwJM+pa7RUHKp+783PP6
759cIKfF5+DR6rjp4QsbJUZWrAtci+Td9cbgdEIdQ9N5HPsOX9U/X5Gst1R4sz9r
x/HyH5+uw7SngbiaEGA7Twv09ynABFKFn4veKjS07+wTJAujGnzBDFqrz2ZEavRb
OC/5fWS+xKmRYEgzXt70QHxca7Pu5xq32fhjqhH0zPdMOq1gLSVTUZOKjoasrBrR
Ow2rEBn6rA9L4RCIuk+c4M5XDvrELPnrCM0rMhDNiGP3DhdA3KSoxWbO15L9PVrY
VKjfL9JTsfnfZHHstpszKfHdLtLE7krh9BqLs9C6zcvhGW8r9BhuMKXgXJ/oto4V
bN8C+H5olT/3YlEPTJLB3lvXXCYWI+wNVMoGwUQ1C+BUA6dtU5Q5IxOg9z+7hFFE
tRbf+HLxANkoJRrA8jDxO/ggv9Kj1K+WFDTT0lKgEiYU5NQjBe2NBV/6JVuxaoyt
GU4v+4IVMXJknz2iuL88zJcb7oc4JHG71MYrLeKkMNOi03iuolYwx48FOvMH1SX8
jENaIp4suqCRNHb1HVQxbshU5O9ol3S5iIhgb78L4ECp0aTjy9RxY4tE3qW22fTq
z/Iiye0ZUPQ5YwaySXiEu3OEKFfN2IJnxqkO7Pavq++WfCJnBjFLh9WXdMHYVlEx
g216o4Bw1ZX20TSKrw7MmhMK6k3I66895xd8LE7RSofaByfE5AYNYGSSp8wf5RQ9
Iu2SbBbDP2ngJjXhQGUrGK0n/HYSIBI6Wg2acC9QP7cXlheDs45XRh6regM+yAo7
BgNeAuBNUZFHw97KEqCGbgnlYJajK+IGC2XeMzBCCyPj5eSIM04ppXbRIsZM9VRD
FB6ATVXY7kSchjbckxC165AgZchgPirJzJ7a51AmTZsO+rTBMtt4dDx8vTrlCIdN
wZ8FUfGg1X8yyFg4YYkTVHYx5RGmCarLwv7JvSLMpXm71U+xHQMM4sn9ET5iG4/Z
hCLmO05C4jyKCs9CHIeno216ccP7m0wkDQdKh8gIUv+Io3vfj3aIiyzTuVB58aLm
oYEvDeH/2GjxU+ahKcgHxj1mfkQH6XErv2f+y6ebFizjy1nto5G0KeZ6eSCsMLA6
/vIkDaHAslai/p2Cmx/znkeQ4LIgQerntdYFuCqVH06JTtPdKa28PklAabeyjVWA
+/qfitYdFMyBUdPh7Pm7WapkavrGMZy+WE2CvbisME7L2XMxr2CQWn67jHrJC3Y+
TNA8f5BFqi9eGCqNVwT9IZCfN4M+j3+s+/8ARVTelkC+j/QP8lrDn2uRUZOFIJXE
b/QFUtCWUVirKM3k1CBfGWcAaxiGbWMXKr6JFRxXkm5DpbUoBGpPbmHlZaGtvRuT
nau8U0YYjDR+J37wGTvd37cvvU4Y/1O2uA1ecK9SRnbzKx7+F8nVNIL/A9A/2eCQ
ZIPjNpQ964NU/0G/5zhcySRldN+EGE79TxV3TbMPEmjNdblYkRkaYX5+pdl1CC/L
sPhakJqdHM4cK5jp13+NEFpQrbjQ+WjXhXrqyqH8jZ07h+h57HTbND25rrKU5bRV
X+h2AatTEDw5a0t2Ql5p3HhyCIvQnm+FPgXL7on5lcLTyTR/RCpJ3QqeU9/NVbKe
1FlnXTeioweCrrWU9jELOaqy38cNzsK9li6+jbfh6C2z9SdbJ137/dphT6fXOaEm
UO5DK1whSvCy/+DjKCuekJ0WZJAtQPCV/QID7KOpbimUezZu6r+kyg5OL84QlD+E
yZsjdGtRLQ9le1QA9aDzkhjQXcyxmA/7liXzJQKxWfsQ1gU5+FfzI9gLyDy51Kka
vgGyakU3gURu8ilyYG9uW51Acg/FWpnBT/c6q3e2PrZnU3F5Snjsf/nNnWE7yyaa
EPd/IqQxy4e0BBQE3QDgVElLaNTWSA3bsTE+pKDSdC3JiLIxtXAjiuVuSx66HjNv
8Kpa8L88EajF8ccoGU1nmSOTpIEMf8jQPAWslSdG36v9Awrl0hkCZE47LQ0mNAef
AtcXnjyubqoOeDFUysL3JbI0N+J8stTJlndtDYIKBdr9cq1yVtUq3Rtu1tD/9hJC
yGtyxycx+gl95Jz6pCvVFIRnwPelluGv/xvBQvgHNse7tQElE8rbEEmo//52HuvQ
RTiYwz9QqTiHcTRc6Iqu1P9yoT0aZqMtCqDlJ+2Ny5ISYYgtAHs7LRvJfvDpSJjP
mo01A1XCo/2yW1eszVMQNHpeukJ1uIXK8+ZLf85EcSlXCyh14hLrvMXv1S958NDb
FHawuBtW28RBge/e6Hs4kxjGx0oU0pId30YuTudO2SFVgcq7Av/2fxOJUi+JmO0A
dSSMfOT7+pYVAX60eC55Qs0jPw9T2bL+73LscmTjAFO306/eVOJAA0PZEIrc+WNa
fKmpIXdUXsZ40wgAgeO7KIoQ0OLDe9u2VW7w9WFdCCF1n+ZGsMM9A15SMvpjMR/S
zeNutSQNMj5tw6oOhUjbNlBy31OagC7hI0CGZby1qG3I3swvUbhEI3FrxzkOwkgk
NoopEaiTctdnIo8XR4yAcXPGTha+KZbCasL2jkPkcVNY6VoZn1WDj01FYa2bHL/v
rmIc5RtVNgU13Q9ReQViIPQIH5CUMUO44cFvM3PYFlCDmF4+2E8vNAkchG/uWfJp
6daPwiB995yXVGw9383YDwul0Q1gnhObcGAfJMeAGUH/fu1NLqtmnz0wvBxqQk2N
Aa1N9pnOIX5fAl7vXW/PlR8LIRcIe9ahvPakOS+zoXITgCAw5hokWoXhq29CAAUZ
8bwMN+lgQZ1DVWmIkhojlYuVLNV6Xu1YYq/Nbn4vpgg23bCH0wmlfW9jsxw3pfft
Yy5Q8ndRncOWgWYoGC/04zavTpzmC8Ry74TnIw4Rx92C8+THmCO8F5UV4kn6tjS5
qk6cUFnR2KqrEG5ao7wVdSrMNKaTqqse1b0Sw7I1/E42okSwB2Y8Sipwvpwq1gec
ea6APDGf4Y7lQT+jgAmwcfdlFQZJAS33l6rKyXcBA9KvvcBWYnRdEB0YkACypKbc
PbOXy/JC2nTbM29k56TDVLb83DfajAvLUN+muLipxYjq8FORQiaVRpNl6nDQWp9P
zSfzTNgEax5VYo96ELnnvEYu03UxwfAPoMmVGw9d3JUvEHYv4K8+orw93rvKYQwI
HP11wLkTKsVUz0xAYYMbwIdx3tNpG9HfYbWgB13I4Tv+jo1fnJjjcg4HPlEyCsw0
q9xxzLoNeQg8VxEyvY4EVp7CkJrpfyPymr5XxaLuElLxBJbrTMOPxTVb3Bv39U4u
lfruqkHRfqGDJfzafgB/uEEPYHoHWobIh++qvbc/9fIEcsiAWTRjQwwMdTY1aQLw
TkWgkpWfym6lT0qNrU32OOZ64/1HE6/YZ+m1LRDwi/ypkwBVF+gAvOuscivE8uOt
q+FvHioULCcTXFrMASJ+MAUl5s4TCHjGFN59FqX60Uw4JKqiAz1goVM1eKWXf/iM
IWNk7vOC88TWLmtuGpH1VhdUz0U2qrsQqCp7IyUaOzSLCfQM6TEHOl94PDz3l1jE
fjSmw0DpxHp7xxKyDg9Nfp6ZsVv3DIMzADd/9SigAMAbJ35Xr1b7lZWugaFGHcUS
b/04lwBunoZJm8prz8MkyMtW+5ekigEiTeGtBc85acA7l/l7XcHTqi5tbkAOshWT
O7No4OQWekZGogrwmx/cDjm7S/AA417Y69LwQx+yj8lPLlmktaxHPYlnNNBxV33P
YDUaZrcyD0JA4zK+zgLm+R88FMaeOqzk+U9LLoWuJeL5HEtWW2rqk0yQhqewmq4w
1Y9r02QWInSPm7JS5PZXxbHqJ23Dg7Evp0TJ0+1ZwSLc/TjWRNZgPmfysxd537H1
c6lkc1RVQhl1O+Rw+Czxdicuv4krbFPx9FtwH5gKI3LtVI6RNIyP+vipO98Clstt
q9hrl8ylwsImcEiLA95CKrlh1prAatljr6FAZ4FNTR3bExeLHRljrCBh1NZYuwOg
Zvc+mTeMfXSCUMO3zuK+qFGZWWfUuswOZFQHaaDlkmjGK77FD28Vn9p/kun4aGpk
z0mrUs9Ic5csn6wtasPPnBOpe2JNLuA7ia4BNV0YCrXJAdu0pixR+eOaw0sPyYHD
ct+W1/82+fIA4lAc0bKj6IbC/VSAyWTkihWC3Dr/+znyCjNfzTpAZ8IJsF3j2ZgX
iaFcrPBNLJ00+ySyGtXYTQNXYz6aVftCi4t9ZvrdMJ8A6vvFFom1Wwy608uJ3zyR
Uptl9KTjJyLkDGaa0e45TXJgLuPtCcCdDD9ybkbbmQi8EDmZhyy/d7riqXD8ls/a
SnAI5Zb++CiN4PC8hxvpyc1U1RNTxOn7199IytmeAWWrW23e6EmvqXQbuVRgsaUw
dqEp2AJ9M7fm08nXBsGoxPpNKL4hw/wnTMSNolZs29KqDF6Xs782rYNugW3MJYA/
xyMn7dgpVaFdNwMKbmSDl49LdTH+i5jMiE0MPGUyGzEhdUya/G74qJfmKXWKUbXB
SHX6HEP5qF0Np7iT3muO1G+Sw7a5si04qRmYe35tTlbpf8MV7CkavBmiyzVpgLz1
iZGuClmta6mwFmYOAgMG5wbj6nVBWUwQBJdKC5Ksp9V8EDhwOUo3XTfNk7oZRtzD
0ZYgWzKfVdq7OO4p6LmQC1WNiZRehghOY8XlniSoTfsCfCNCwDbDC60egO6uazuF
7OeHxI/vkqORnioBT9wcKK1mZhfSz/GCMNTUJBYG6pZDAK6cdwz6VQN2+48Ve3d5
5DkKf6HTCEnMPAadIaPjPGnebftnkICJedEO/wutV4rw2lxIpXT3lciZ0T/jIovs
+Uke0PgWGVWc+G0ykF4UpQrkBB4IQ6llDiG7drdspm9mzUg/qVLQUGgaIEDfJlh0
6kBCoiZbCHnebr8HBNFIm61woUM5lXMuaZ+XnOX/yYoeVL8NhZsJjxiSxTzFSvRs
aiB8pbMCZv/WPqGSEp1jpkCGJQGXwLlijyQRD+FU0eGAKAxR85nAO+eZNxL8BR41
m6uNI2B7LOVjEQROsnTwtvZFHtgqDkV0/08abR7rSFYd6UDhQphflSefhkOyMD1S
GXeXfw749nLlhfy0ZCvD68XCUUlbvorxi5zTVEGA6YQwv1RfrEtONj+ebcWqqjM7
W0mU0Ucumr+6tj6fpCs7C37IkWIV8+bXYh4eX0UTJ+QiUcT5v9CQ/IHkAw3Z0Wh/
WiWfe8jDklIx8IQE6p+KEI/hW44D0PjQlXwHzs29JVUh9Ru9e59fg0SvKsFRWAc/
Fv9ghN0rcAAstP9bO7FoVN2QSv+3yenPtnfdx+c44+jJIY92Z7VhZRuf4CQPR1+j
RZ7SKn3PjWzSocMA5sRJsI8XaN9i1QvmowfSYlnP1pPX7jVPmdN4BfSib1XMCi1J
J6faWmnzk7o6Ic827oRfzBkyrWVH1ooWL92FN3+VwCk/ZN9rZi7UJFCP+3T43BGt
FZqrcRdI6R3bGcjdf2wyl4dbRvkhNgy/J7EBCjOrZ5O+oLXF+KwQZ0sqL8Fnu4OK
BCxV/H3ahIYdoL+eiRt74oZ8iQ/+kjUVztb754i/lC4GhVZvSurqN58d3gSGNyJg
wD7dSYf3VdLTHLoSQcOgfNE0OdJCEzCRLFOhZXv7yxQIswz8tX4cPPS65vPeXmOO
e1xFjN2PaKQYUwOiLp/guaYJog68m/z+QVOaVDB/U/58lYdMQH+d+mwBkfr8aDOo
Jyx1tiiD/k50q82iti8qw2ZVwMaczMtGkz41X/kPmTrYSkrvLZOfUOTblVQFgbZe
oSpUhNoQ9NTUdWJvzmdkulYZOnKeEsIoZQOpPhrmAp28/1L1kUhO81xCMR3PVkpm
gYIRllUyN8N8Y0Ah2kD3exIDFpFMSDOy/jgoucyid1mxP5ikwKLGRO2En5mqQhVS
OvCcWTuWRXlQfs8aXbcoxZdtoIjZTBRzVY3Jkkr5o1/+dOL6MfsznpPmxmtEqjvb
AmjLoXHIrKUkeC/oEwA1iPGwWMvcsDG1HRtvhF6dMuWOxySNfsqPW/jSwIP15HeX
sjaCdSPBjQbXJbqX5ic8rI8CHZSzT1z27W1QAjGYxKT83Ch9E8X65/wke7iMuMpO
uO7HOvOglBP6D7WJDbHCu7oVCFqoY4OPA0+jPNLHmG1W3JEUOS94zMNn4e5+BZw5
XHKYMtai/gI114bi3g2pjyZ4+d1V+SEoOHrNDKbAYOcasIY0XbuVZl+Uv6MGGl9H
e8wzLnlZuDxj8vZAS5L3SVdJc8lou6NgPgaqM6rgx1Lmq/OpuIQsYd3ScvfIOckK
dpF3bjWip2WT/0lcVsx++WEqTsDI7ThL+dOfiyWIhJei5ElCLDL3YrOYgatANrNr
bVpugnzd5Hngsn8COL83M7nCm2ReBYTnIKvobjIDo5uutcOoHIXjTHWtYahXKb5F
FD/FPiU1xxGVKxmh4GADfy6dNTDFHSEbALGfcyvrgF1NKvQBESTunwBBUHVrIgQ/
bhGk9eeHMxCTtL8ckoZGhwmCL67s0w79NrLTe6Gsy7sI9SwA3K/wnnnxZ2FKQrLR
0zuXfgSZABfzZKaaojQ+SBB1/4568GwoT7b2u9vWWotwCtrAt44zSZIlTxLxTvyL
IL7bRghixlIzWCIdDbBIMzPrsTMjaWSxxOZ0IoHBt2em9NT7ag/0NFXwW0qM/W+b
ryYElCPrt5JCNL+zka28Z0ep42kbgmEcwRTv5mfkCGpLlYoFYVkwkhn6xbfH/Ffv
I4YTCOp0wPweq90YOL3cO2wruFhTrDGAfJ2rMsrbcJvMMFi2diL3p1TNm6fZw3mD
T5ZwBgnNOxD5yVO4m5Ymo2e2QDZVZAKQ8cr9O+fb2tEPmBXPaz0K3DscTxp0JgBA
Q1h1C585mPfNpfmkROSzzt3wpzCl6yamli0rPXzdAqTaWagvfA7zd9k7sP25U7oC
NIXdifFrVbt3F33v13gkpuDIzRlAsJdRo+BEXtNcunsa75G6eeS3VMPFrEWcf52+
+r0nMPK3rYx41D7dWzphRc/bujoVVBqCStGdpgqQyvAJxW807k825zuGeMVkPoQr
nkx2sXLgRTIfLTM6WwIDicNKRo6tZ8z4kTzeQOkZNO2KDAGyaFtD/Rcj2tUwR+hG
hdDqTVxDgB9l0haPPgTpLuWhYEJoMDKkJw1ZVnfPCAxy01gr1XQLscpczPFd/3zu
De+N8njv6ZISICH2k7OQZOeFiJwNalC9CXhYjN4VlaK1KDa+BI9lGN6QFE4FYyYR
+lexP0r3mMoIgNkFbDpPzo9x11QGUCuvqs3M3HoAnu3x5zq1C+kPAe/a04FZbauP
4FwhC0y6lZ7SLdI9+q1dn2RpfuOm5Dn7Co4k8lX3HjHASdJs5XTpriUE5T2TghIb
AzUyKXG4g2MSkXGfqC2v384wAHSIE61WR8dmP/zS5NYZVdvlkhIYOgV0W2jXeR2h
/ndirH8JH+IQrQSWDCZ6oTiy6UEJvsjReEEmKH8VmYyTqc8yf76hXJ0v/bMVghZ5
WIdsRtASn28NYRIOvllmAKLu3QpgmW9LQHIFkuGXT5alNRJyUbeHKF9r0jlgDFDl
mI7F/SzolGGK30unDtqDo4KAk/PSt7y7aXuI/guLIrT8hCd3v1Rv452OFAJTxLaO
VVVHPL0yBrAKq5xEswICWspEctbXBqzgFuwbBzMpNBMhguLzADtX9RpLpDRKF1aR
o/zxItsWdanSYssFNomzw4WrJfCZUcyc7iK3m9F4WfrR2ZpDe58y/ByhmkA+6d+y
mYQwlC9aVIiCyqFWynjsRKhLYWadF4ItihO/qlh1z9WQUSFFvxaFk19kO1wxryDx
JBwrosR5YXE3e+XWK0hzzkKOUYb07bWuczuNMft+1vXdo/MDa3dLALEP/IxDlIo8
G+sovi39vz5wBwwEddZyD3oIsDdUdVue/zoCkGhTeI4DvGDkdz8excg3VaS0sBLF
VyULHVKZqHJ+9gOn1HfBYPouvOU7Uc97QVGwBks7sc9pDmfOnUlqzgj2ngre8z5J
8ngJCYb8/rY4uwcl1RRmbgyirGKzboti4koBV9ArUNuALSXvbLAQTWugpKxugXN2
i0zayE72S+wyXfPOAjx1gfMtC7kvL9UfORNLs8xZ1qcfhcPB2ADATRHvQDwQ4cwE
nCROvS2LwpyRohJKlk5dbvkBmPeuF10NFLXdzppb80ShTf3zNzMKO7p6N83o7Rps
9V62D3btIb6/v2JlDU8AIW6+ooaXQ+rtWr7LBibqVRj3/tM/7ZXqmI9jI62wuJQM
0fk3JeQy4Bfmj3Lm+DoscLz7hLhwrfTc9HCo3HTWauH69pMoU6ciMvXBj5KABXd8
kIfEeFei2cTw8dUEytn/1cltoRM/L/dKmrcy93tYfekvYlBSp8OZJRD6Hfi9DodO
hA6xrqSiE3ntsTo8V9hR+xeqxPlULLFakUDJeTppH83PSkBDXS02cXujU0iBiXCQ
DvaOr0WuVS2vK1CnqqE1RW7+STbPWGewM1UwlmmwCb4FiR6+zXZWOHBTfdVx/JB4
FEQshTccdgfL9K6/KPrrq74QkSTxwQlCKtUeout9Iud8jaXDVVKGkSHLsNniBFuA
J+L91IXTIS+2MFNeBlEpoIXBxNvZmWcEOm8be/HLvzZECOB1Kr4KnbGAiW+Yv4qK
FszH9875oXsLntpo+hdATwvTjRVDcHARDqPnNbLfIgz20ENBY0T5MvgufiJa8rFG
575ZEqhU3mpYdZT6uFztqbjpt3fULF7eyToqUi+5UQss/LHD3wHEFfkn7I6MoP0q
LUe8X+hrkooAcDN2OQd57bd66AlhxEvEqU/ZUdBEZ4mawsIGh3DfHSUIVCgmStKO
zBGYwW1EqtYSdbglM15CqogegdFRFLA6s9w7dWXcp21Ffjroe+vlSLN6WeStfBEt
NhF9ORCUJc3HVwHjAWtuc3iTjOggJulq+T+PFibc4wnjaxMSocTfq55yVFwO1f+R
4Tb/o7DQmLpUN4c54wPJdGyxI/5KukbCiQ2u3jILcZD790+3/y6PmXIe1V1qTmWa
SQpT0VrZ4I1hCo/SWt3uBaC0H/ma3vgFBcGSjsYD1Fda+FqLyra45/SpdmiYN2rf
vdHfGAqsXDNVzXxOLtdX+GbC/v/wsjFNBO4In/k6yYoVX3yRwIimuaJr4Kldiz9b
dRtJZ6/gPFkXkWA4CqdhkVjnbQC5ICZd/AedZf9Ugpl2wvlrhm7fZJHX4UQ1rdcc
IFRVQn3fsv/7+VwFYXWxd/gryvNx+lmN6s1nTxBofzbpa1ASezOl0ICNX2wrrRmi
vS3RfKhl1PE3mOKMnJndgFSfiZiq31ir3+8dJdk33o3fx4SZHHICl9WTsTW2+DDc
do13089PGYdZ6+fb7f4j161s520HKLON13fJ4S7csQcpTn3TT+vw4yNWxugN0ZQr
mSOJjBa/w5vTKRKezxjmb+EwALtz32BZY+rx5Zs/Y9/IiPVVNrbTA488wlRDGqE/
XIAQHJkKcrfRZCtQgU4VbLaiuGV4LtjIFN7N5pgFEFs6YIP6BLKtRUl7OK6BeGlC
obvHTVkqz5F3tdp3APdToOGY2jGs12yk5qbq5swMWN+3LygNSfl+mv1ncmpcBv/f
2RzuBmxudMBg0tipLkDYH+4ol7v8HJqJe8l4uBeurpt+RHfec/WKYm+FWWJjnk1Q
ffwZhWRABDs4y0r7vXZBL+AeGnOeA+LQ/W96ozP8wNmHzoa9KIzuyUNDjeFv1Htt
bfbkHkd4xuJIhwcMhZKbzaieH//mTh+He8eifc7ME0Ov2Idbp1VsVJ2AoWdUM6dU
gF6iE8UCqsqu6BnnuMr/1IIS86TMr0WsLmHnbkTtiKYXClZZ8YEU5gHCeNuou5xS
K0ECkRbhxC44Q5U5Hka/OGN9270bBWNZJkW9oA1eqajwFWcMBibAsNZIJBnGhfAg
xV3AX2Ncm5N8JShKEzZr0nz0wfNCgVAuyvwGHnW1MjBHC37+gtLvkcJRqLDlLxde
sxStvU+rIvaqBiNZqWbI7GF1FniY6JhMz8s31vAJ+G2YL1rignFmPt/smlynu66w
IKthSSsbC0H6k1pqU2NzV8f3hHAHIDWkh+0WhimVQOCtwfQxjW1NIR4A8OiI48L1
KxU5Y/2kBVltHCA0x5cIkQctEajo7J+Xx8VJI4dt6RAUbj7twFVMCedZZfaNoLfV
ah5lHWlKbvJUH3MmWgaoSwh1JEALM7eyeEiHI1V0lwP/IP1ca8HmCfgxZqpm7KMg
cE7VJ/eU9H4uOJQu/BpubQBaKtxgly3E25SIIF+xHglIhKvUneScYR90BcxgyWKB
EM1LpWWYhmYvP0/UZy2XOBUjQiXxHVKkHhty3HI5W+Wf2cBGyqD7AwVSpmHPRaFK
UsqKu9HAv341JCElrAec35mkabdvz0Ld/v34nPMhAm0tut4Z9dR8bhjFaVPNMUsX
VK4uJsRDudQJTBUdiUNuHgp5ifLVULaeAtams3tP+qj2S/68Oe+ArlINJj4g+jFc
lFn3VkbRp413MPe9MW0o7oTY5wdaBoaTBsDRwymq30i5cFxjciXr5WkK2kqhHFd0
VS24r3muiHlVo5pUKWMvzoFEDMQq7Cq/7At3T4KIQNCzlcWVyyktnQOT/yK4uNRn
UwpPxiqPbNzfNBbR6eadHAaNrp+PKmHK5FMs62g1TkVUG75dHYRRb0H5PR/qgUMl
cFFMQlrGQxZqmFmXoApPLN2kyzZ0AHyxWSoNp1r0owxSyQ6iZJ/qlAz0FaEsLviF
hXQQqvjkRInPqb0basr4UKEaYG668IEBy6HkLmb22wjeomlrjW3v3aTiUQZQ2niy
v09Aa2l7eTwqFNiLABiw2sfk5mBSyNSgfP8CFK2/BT6djPd3YSk71wbMluXV7xws
AmMvFEqB8kQvLAevL8XvhiyTv+8BSNHHj4EqzoNmxf5e9Gd+eufXFKd4XvwhQEMu
Fr+Id/hSowExgnbItSBKDWmnDXK2y2sT+fcm+BmzJBJNK6jBifscjyB4HQodlTvU
aPKR4u/qO65M12nYpNII2VTQ5cspHjzSNq8imQIa8Fzd9Vc5U+5jaKb9NL7giQ8n
jMl8yKCAYja/pf6V5IEKFYfXBsv/Ju3wnqjmbfeOvY9sgopmU+/+VhAwpBHC67nB
zT8uTxh/AYDjTAwTs3f2n1hUgw4VLQip1bYPOw8ACvpyhGCTLHFAOAdHZUAYo8w7
EJCuPa37LMrx82aj8b0rgOa3RBXDO3NXynqewEnYcIRjQHRKjVjNGmljpFXZYuNF
kwa4wTtlyDzRY6QBM8KUbKcc3ZpL9OiVJb56Kwc3udUPV6cOi4LkP3IrW3np72h5
qgm3mQjQFKxKRYmFNmanchH7YOBI3qVukOpBaQ03g5ElkFNyi8w0F+GHHNsh7UWx
UVODhqF+leDqqWQHzUWDHISYgy45jxg+c+Ex3LnE4X2UznBdDaOwxDu48jO7Q34T
4Je43SxVvLQ40tk5J+4ivSRGCTVY/kbuaIIDiBfc/PNCwBQObUs7BDEEIdNAgElx
U0qWqoLBxCqsQCPrI30FERDSqYJnZ9v4Ei5Lq0GFXY7XcMtrMwz4S9sF0G1hWtra
/HJcvxiAEhDMXXLJgHA7DChwPek+vz5KodUVBV+yYs/SM6T5QvSf01aO4kEXfqCC
PkzgLyIWJLmyaBH9beXvRQqzqBlK8MDHZy4/Mkp1m8EqWQE3N/7MhZB+0ZNTpDXx
dgAKmQoQFN8/lZmjfZ8G1oH3n8V3ppUpm94efzzdNAzoDR/o07wnfz2hhSHejjqU
61jVTx42lHCmYzTr6s1u9IG+uG84rSoIE1OPaHoUnFyu/jfWAawUjXSZ6wSH7P6H
5R7SGqYWS9cQdRb6P5sRd5aTIYSgr+N+2iZiZ5nMjXsV3J5z1Pxh8hfv7lD7SmvD
YDwSch+1mtimGc6vFMERIr3Lrc03IUXz6bEKi72PwPtNVUOM/4m2bn/OJ5kuRKoj
HBYtjwrBWgiOra8zHHKLq05sttn6WiNR4ZGr8rXlGdR250T3TygyW4j65ub/4Lxw
cAkmVEOl0XZqVACDSmGAXEAaXy0di7QMAOia/531gIIvVSKC26CxjefmrFbO9nAR
frLae+vqicWLC0+to3hSWV6KKPDA780KeBBDuYhFp0sGtVXVDgY0sTrqCyD8buRZ
3mQMW6YqiublkKTnYMIKMpKIYqxnSyfz5Vl2ZkT6kAAgH+NJp1mpMd6YjLvDEgZt
RqauPkm+tR0G4lo09pwlqNHZkvcfTNviPgKgB+NyBlVjxfN8zul6BEOPVz5d2xYW
eYaTK/SHoqkMAJPuhXnNy00j6rF7M7/bMLbSMuSGIr95LtItYBIlVM5CIxO8ev8J
r7Th1jD9dmeL/mwxZ7hzKYNcRzk7pz54a7CPNYuZjaBjpkUYqeIoaloC5vlT25wD
SRJXikFNYnuG3T/T1zSj+YBZznDFa0NK/sUCvBf8IcsYvcJv4mJO/tsw9LvWjIeI
E8DSx2M0LMNkqCo6GQ1n2sCamey6z1Af3LF5lRUagSNGMJ3U6rInQbsNIr063+UD
a5TNzFjoMBCNYg87h6B88ObcVxVqrc5STFoHCsosxNIiLBcC8IPjAe15rrnO3yCd
3CoxZkcjDgUfCdGdYLx5xw9AEnaBuDtyVlwoOh4GHR5O0XxBYLNug3vZuY9B+lkY
OA3FE+Sbfzwm2FcD1uuCfRLBofU+iZ9elkisdR/EhFQX99Sw045ilxHGRB2VefsK
fPAgqN7NjlyQu50+rkGvGzViLfepqQ2CdpqhFnzwbAW1yVdNDXhEuK6KvIKR+qCm
wMHzSuamGN4i951NUgdt80ST4TtCEeFzo7CVzTJTZOssrGwf7LTVH1ZFF2hbYUHd
pewMqm8itNUXjxc6Hl9Uom2GhyVOTq/NeeQjuLtKW32qwOLgTDducqH7IDoXUhGr
JgNZU3VnJCxiaCCwTxQFSAm/WZzzDmpMyq5grciiYDkDAqiwhTvYp2yo/hkbEYYq
GCnAmF9H6ig6gGREkjC78i/URin2TIgQtDQd00iH3olVHqcqGu74A0pwkWl1RXDo
tX1sSaaboVQIJW+YvW4IgLhIRXcDG6Z9p60UhlqMyG1Q+aV5TNdBPPnK3WvPv25H
8kh+U+crFmdNDcrDUiwOdYtDl2GmVN026QANEKx1DdCv+JLg3D7ovy3fUsKE9eph
9kI0ktjKzEjGhqgUwgnD9lnlgiJvf51yaPDWC+b3BcCSlnx2Sua+6/Y/MlxukEyw
nZbJetcKSsISPINFMJn8F49B0oU7q61TIDn80dJ2iBQa1JGhHBFiSA4dy5cx27F8
KSBUG1n5lND63fLlj7MwIF48n0cHdvv2Xy0b3+KAyrE8xCtDsD3u727M2H0pfGV2
eoXLotI4plU0Pha9eztZc1hGAxQ/htej+4rs/ZaWNf1110R87Ls9iVLdwQ26OMyu
K6r5GB2b15HwlH89S6BOsn7rqFXq8JDmt3j1WBfLluKTy9nlacuUvkpaWH4wj9qN
PcZFZnuqx+QWD9uTlFXJJNJIV064FM6KmQdwOdmSQoL/Jo9qEfr5FERlDXTBXQqe
gZXQwlhSHG58HQzmEE8TeHk6nUwb31VvKalLzktdvu+HimQ0bWyjrcP/7Y1+xRMn
jSqP4AnZ69HjPMFgx3lZLqnlBR0zimCZyuKIyj6xe/YrAagK8rX439RP+5/foxh9
Kh/UoYS9rIvWW25t44UdcaHdSPdLVX8YVgSXMGbEzz8Sxzhv9ln9c3DSgekmJt9D
dqyET1Xct6fs0B5yM3XSSAlLErQq193OFMAL/pUIccka3PY0gW7HNOS/l+PWUOHo
iMYSNZfpnFzicHpjPBGB8RSRXqIPx0qhOOGfLcB5TorXJIj4B5k6r22BalwSPxIq
Loj3imsqqOFjgiXzi+TvFYbTRnCLFpWyyMobROg8UH/WUY6F2zfW2nA9bbWCgKYK
QTGg49ZtvEGr5ehsyyP7jII29pFaUZV0F7HAoiTOtCibHLy3pGyo8egvYqGD/qae
HmaW2n8JYb/UjeeHO1+rROfvyLl2+OP6tyHLGMa2iU0SC2iu7EAxKzPd44g20hsn
VumixwBDX7gr3wH2eiono09FCS20jlEuc0xnQxf1mxe95JpgBtWVjQuBg32Z00C8
Ls7+qynsN1BSqhLUQC92Q06+PTLWmn3TtD05xPc1VoiRllTrSGpbmWH6iZrF3Wj6
ANdFrZ2PCw1QwBdvEeuSkvSfKP7laz4weZ9YuCJQEVoszcGUo6rejfo2g5hFb7DF
KtWkuOyL2bb8+r73ncVRmFhAuS6DoxsHy6/fVv2jBw1Ocr6/jADZMyktY89blxgT
1Rx1dZe4aELLA3FxV1dmhFExoqT8b9rGrAf5qORV3aijEn/L+/rlU6TgBLclLnVg
gYuPPZ5SN0GrgOxMbD8i2PRNte1cIibwX58fS/oC3NRNbw/sGR6oDUihJ/EriQm9
sGAIWPjoAiKRdW8jQqbgbwrUrbaNp5voiXwx/Nx6fzCzqcrqACYS5UWqFHJUHpQV
zjn96QhZWR0tePlNvdFCl4dO5dsy6NlhkcKCmpVCj9OSNiHwA34Galc5i89rZOM0
WfXk9dX1o3SseSLhMVs4exThXLU4K2gUoYs15jWOvrOX7QzZ7ORtsCB13wGXViXk
iP8S7LCs8VcijEubxjK1IsstYZ0lXJwRChnH0xjFBNKvFiIYqRu3COK2wzyYGrjk
teXTSaWzLWFgbuSMEkbFIZ3Q+ZlYbbAiTK+KX0LGVVraZGsRtPecCWvbz3j2Kq3l
KQ2qcKQbudWHvvea+Rb/YdF8oanFi9DCmqhME02ID30sZkUEncnLLEOn7M2OlUtT
WMaGEucCjBHwPh+ZaGujC8gdq2iIy/VDAjehJmvpHXwZ3gEkKznsx0kjZgpAiYyp
xwaXz8AFZLkR/KXD4ILPLkG+0sjHjfxGMevlroGt5bQ+BS1oNBcyTj5DzC9SU4+r
R9mT/B4AA9u0UuDI7TfYc10vHxtIMGhz1CFJqHPndCmdgAeitive8cT03jz7+L98
HL8seUAVAuf33UW9mWDD9h9LW8hWDdDM0U0vSUFE9XwOD60a5BuU9wwq7YIg6+7o
Au3UsbSM897IYQi2cTdaJ7ad1hOiGZHubOe6n4Um9XvRpDL216ee567DqbrPHWiT
V+1P3t6lb5+1nfsDDp8fHSJEVAovTtF+P/XpNZvgyiw70SOo0v0m5SeMyQ71JHbv
5Ti0+xQu1zSc/9fg3CG8IexiUWfCnK9t9u/pWVRz6YPvDGqNEhIC4+A9a5VnzocS
VGrrZm0NChhcpFWBam1kaSFSaZYiqK00TyVGVoWAkuM2ovbPx9w3Jh/iNOPilRgm
YA33QIJOxYzVLYheT4BKAmwDJckCCNobkX3D8w62WmXqOKoJ5LvcLZ20I5YpUXzb
cekt4+y0tqwaxjbZ8gSfRQl+SkyOiPs/OrvLYbfQhlpZO8TzOQHPdYBXxWoMyG9Z
J6YARDYwkLHZsVkWObLRaxAfgDAgBUxl2/N2ptqTEMmQZmqRqKD1W79yz/aivxg5
vdY16A6Blvdeypje5IDx4C8Z+AVg/Lu63NW1nnvQp5KvgTAL45UxG/dkMZx6uUFr
WvpD/o6lwt7Tqqn54DOmWx1scWlDu9EmaacXM5Flk+Vd5lpwTPrJ5ExqtBhlYgL5
TxT/qrRB1CyAihuW63N8VYWAjUTVzJpT/1TGWVvhQIp2n7ClmKWQGOKMyed34108
SuXnc9nFareP9U7WV9MkHLP3FTonNBQlop0CcStU3Gshx1JYBUTnyVvoZaUqi6+7
EMlZZksAq38uc9yt2Mv5WkU3GlUF/vbewzCd+XCS83f3/k/qcxNDgYy6aSX4N4/P
28CoDaf0UL5z3zXNzoXujlaB1jZgFvmLxLCVZ3bEaons5JOVyALt8RLHbalR1R1d
2yRRzH/P8QoUMHlVvF8No9uwOMneWEWXXXYkiC+mPzP03IiTv5zrW+I9GxwgtE14
WLzfacgEcbuMw/fH2k/OC/75KasyxmzZX8mMhXgMgSXhWPLwuETNbUfLL4THvSts
nrpC0xXJYjioU9Riye1ruEGu6IqrDjNMQHC8KPe6zjZMS7K90i+Ebmjejv50FP1e
UGJL2YsdPsrZ8+MhaoMxJMD9yzIQ0RcyE0+wQreriw9F8NNSLp4ic58QPIb8G5wz
ZIWioZcWj2vBaUK0/K77141NnyvYAa7tYwEP6lDkWrEwoP7iEOhaAIMJPHeBb8my
x46IgIE4/dzBlgbpcQYw1OWXpzoA9kDd2EZ1NpkW9ikIMVkKb8CyHXGnRtyi46gB
m7HiUVgh1K+hCJo4TR2C6PyLnz25XtQIJO5lWWomr3j4vMFuyDYVe06g6jJNQtXd
6U0up+cSLjpqfB3EzyQ7lZI3ClMjTue/oqlvcMRToETv/CYS9IOGbr6GChUGL9Uk
yn4wb5a92U+RjWbf7anR5DGqJGlGIzDyBN4r/Ocg2RCWncD1Lc0XpYPM2wv68yRr
2YvNWl3sU8hxZxo7XwJGWSKxz5RZLGiUAw2MjVhdJeXjRELd9XL2nPEw50iDf0vL
6vwiO63cns0Dl2nkx5jIl745MhhReu/JTH7TBOWWMcw0SfKUaGw+St/eJLV9H2eB
AdzXFmgvDC70k1w0CjDECoJuzVOD4FzgOpk90ge1V1dB8Z5DltftEu9LrE43Hw7s
vwBls2DoY3PgorrsICiFYw19N0ACq8KkQfGEvKPDhruULd7E2GRl9gUK2CX9jNit
u66oGWJELn3PD9MQNYarh05qDKY2jblUKQjTTjdBZUAbPNiYM303P4hcdIUves8/
bj+mk5nTrwnBBbYavuZ6+HEg/9bQyWWFuzqtYHpuKgvTXr9onVLxvmIc0pzk28IL
AlkOWvwL2T8bU5a9xGJD/ACLMw6mrmBS5VGxP2AnW3maz1atiNRMcQ7cezfIky7D
mQ7R9IUZaPNY9U/97vGH5oziTo16c492dK0oaePoDVP0LouhncgK7T471F5DDB0k
+YD7Z7Mnezy0qomynOA7NDbIOZIafBckUAG8kjKdjPlKtYxRnTDUh3/GTJeQ1FvD
ANDnqiHcjAGWWkdbpvG9TmK7LYDDCclDoWdGdPNx6X3UnfY6xYeHYutHOUNC6EF8
9pTm54/mV+HnirViqpgPgfP9Qp2IHb/KZ9hMARFQZudQzSfRghHZhF4fdd2VKtff
Dkpj6pQGFORzeH85ONc0R9yCFIZqwIbfFI+MMGoi85WjDwZ3kfJhItqbXF41iJSw
ytWZiqYjaSG67iPC0oY7fxZvjbzqXk2cIDZDCWE84KSFtO8jg6uMrxb2gYiY88wm
Wwad8EW8/GbY0UoLv2WY5X0m5qUxHClKNJG013f6nMG+OAdIF0/bnqHv7WPuSu8t
3kkJH+6pmv+YqiF9pnXRap3ntsymH9QdXvL5crAGmeZ8PFNke1osM9NwBSHAhUvi
BGc0ZwLSnHlqICNYma/RolRzYyurnuJXokS9wNcKxRUwttGnslD64FNQwXzMg67e
FCG4fmIp4W/k/OYQVewNHbHvEnKG8STjJX0YGhqEqc4TxIFB/2ubTDGnmlpYwFic
zxfLgJgs6B1YrdKfSF78UD6GJ0vXS65Cnb3iOnXXpnIQg8OfMcPhmIPIsi3GYrI/
qTf3uHdRn4iChiLy0EkLcQpePVLIsm/c5m/yiWi/Tcj344SEkHa+Np5n0cbfH+1w
IC+F8kDGkK1+1V7WdX61jVohru2FlZ8lLmR9qSjIiW2B4UT/p4yW16cOZGfKdN6D
+yzILQ7gRQ2YizUMQA54a7kZGEPjMXAd0nOmFrWimx6AWVHcZm3IS6rFUNvGVOQh
uXepLE+JKPCt2a7uIYVk6vF4mVvNSGX9ysVB4thhWmq8SGSVUuirxKGT/bXUo4ZR
kk0tWwfjfWDgdaHYzHZcQtSkbC1l887vXb69oJsxpRdIzvP+fZgOmwrECN8gOBjn
4HdBxWVmq9MsccUmazNv98h3lvbstglWA6nLyL2E5Z6S9C2qkRQvdqxpItusNjIA
cFNIE/EmJddtIEdGpl8b55m0igr4p9KxWoQlwvLlHf5P0OPAxjbK26tzmw/Y8bsd
q/Ul2VvLwCilycBI84BEai5S1lFnTiKiiyWMqPbaUl0Qk6Bmv03hzcnplNwc6MaP
EVlqADzfytGERdOpADC26WxU9ofYAEWs5TmebI2MYZcWa6yXs4lnqCYr+waZLgxZ
lmE9F96VGhIZ+ul5nIKmfckUVJ112Kddpi8T3CTLRvXECYpgvxCZHQiDl+CZA3wU
qYcup9r8f6WSveUabxw5d61F3w+INFH8TVJBtrsrWhZE/b7GJHypn/WQtj+C+9NY
+I1AneQ0kzLecK0aGM7SM7rrWQ4Z1rqxepwu8nsDUvOaa9lO5p0J1xMOh5uD2aND
3gTRrSoQYzif5wwO4TAY9927lPCaXgMgaHpx70eFjrs9vVYaLGNQnwBPMdTSnklK
PSFXt1E26Suh4Br9Y/abHb5xRQC3rg2hjMNKdChbTk5m/e+lP6r6GAO7AOmiRjTc
fRxjHpF4t/aGW1vU7vC4cGEyPIHZaYBG+Cc8D7LZ3dmrEMkHsmi/yf0BKCTMh7oR
pwYWh53VV7pb2IctbUDlL3HQaIUmKxDpjopeLx0I2KO+iGxwb42L77TJfnVBswoH
MLo9xMu5Kmpmb8GpnDI88qCVOG42X2WxhibREvrY1lB+GPX7La2WF37C8PTU1yyE
1GrUvXCV/+VA5nigrDbfV5kNFsBAgWk6NtY2LOvNbUSiaWbm5H5Nzz6Y7F85kbQv
HV8kyqIwVmbh/86XK+fgvf6xnWNF0zFjKEjMOcOSQksWPwP1PqBAa3F+KwcmKdGi
EMKDmpFQMTeTufQTEZKAwECD8IOJWGOLstSgZbJ9Zd1iKcs1OJsqJy2R9G+/7gbM
tG0fjCdsIhgTIjh7m5Q72WBsAMbnSrtOtYG4MoHF/Qxsg47Z0IOCx9y+OoXxOxoW
BjDuIXgk4zfpJIQCieLKL/dPZj5lVAMnpfnUzLtcAA3NG8FQCrPhYf6MjOy1LMRv
smv19JczLJp7s6TVj3pp4cUHBuob73zLHtQHhP0ZYDK/afBurj1ocZ8ekg7G5rPN
hTo/coPROIiUatfnVPwGUuanIQCdsvAOenMHsZYkigMuauixt08N4ZNnoU9oCTH4
3/ZMojNZgCemymogkp3hRo78nvTp0/3lFgbXu/0fGLJF56jC8zrHHVMikHwh9qUw
VhikWBxqV75Rc55V7hLvPcQl1LfuTi73LJVfU4IA+fxjVinqabl9EZrx4DXUrxIh
BRpguP/M+G1hfBtAqcu4JhNPHw9D0VctnJmskS0ulOUsLZ0wABsa19uroTYCz5j9
CQ+U+sxO7fjR/ZNT2G3CEwwvRq21Okg1SzlOCOe/NXktSjlYL3593gV8KaumtEeV
8HTUIIcGNBhBYmqRuqqci4RZYjCs2U8tFkuv5h6zCfss3dKqnn/XxZiEhJPcjMEO
4xOoaFKNswbeNPaZV+MML9a3iJylf9QFIuUtPT6PfNV5HATvOqmkDHjfTykbwoJ4
v9Zj8hyX6Tbdy/ZRQhC1ijbDiyRAnmhBEp9BlvV570mnpcCyuYDmfQWhZ91DXstP
yocElYgISDV5hst9l4w58NTjqtN5F9IrQSskKmPOSuHyz+jWiBflCMUqa3RxtNIn
qjat2MyLZYVYjTNITAvAhiS9T5DPyvdGtLyVOF/gUdoQ/gDmga59lqwb8yIvDFNT
6+2p8Qd03wMLZMmMZdvo8OdmSCoT+yNGVKamfS1yaD+rPTaSHof80gj4tqBqja2h
udJ0DXCTEJlxcF1MlvCjr0YMnOwuH7J4JEpjhoRyFb4jlSJkugK8jf1Nlx1c1I73
KH3/4oiQTmgFMgyfOHsXtrUuDnem1/GRh0zN6Zn5qHtZt7ZZkalNsu99ksjknCir
OiWRx0XYPXn0Z+seU0mp9/a3bA3/KMa1+uLB3Xxe/7da5SuGVOqk5gTQ9HTgyb6/
DEMqWchaHTNVrjWvmvu5JAxsr0NaTEEXyS2J+eAnQe1164G0oKqN9vTYh05PVQLP
Q8Sw5dR2x0GS72k7+qRj9QsB8lxEGK8r2CbdO1HQ64Fau4pGzTt7m+Baa0dHRL1R
J6jdGD0phwOKIaisITbbOYEhfT8rEFCIZsaoHC5P7EKmvR+23nY5LepbGhqR+FpN
ZwAM9zB5rkCPi1DJA/O0RkQ1L+VyjBiY3k2u6m28w8YuBoAw11S301YC7ym76aKP
PHbMYc1Wxcw/2TAxs1Ri5Vz+RV01HBF5WNsMeArwaSmgYnIR2MWrZfWvQaLqtv1i
pKFcQtO8UTDaPhde1JQbWow+Zvf4Ff7skOMeaZ0N4ClioBbIdnvBNzD1qZXDFQp3
/eqzJX4s6p6xnHu4d+0aIo1b9Mb+JIIYkNdgkTAIEM+m5snJVwqBDV1yQBgo2o4e
czKzqOnnA2DNvasulGZKZ3HUbiIYv3OYuUq6HhD+LmY4Oa6X063YVvKUUpjGEY09
t5B1aPlY2n6JuZFTFliKeFhYERxR5kJKy16fxIX1iMNH9uAvzDep6qERvZ8wkQqd
ly/fKknOAjZfC6hLGMlT3IkkcFPSTkfAtb4fVaMc1nyT1kPNVpY5c1JhnGkPTxuQ
CQCQnKpSTjHq46aL85r3fONRLM2f1wqSESovelprofUhZ4iPS0nDqbu+mODDXf1v
3ztPBSn9N1GQI522OZjttloSatBgEDuVjPWXna8+Dd04WkIsXu+PJ/0bL46Kz76Q
j+jsYAgHkmOvZP50WvIyJPxOJTwmC1NaT+TQZYdyN09HvfQcgX/eYEI9mEziFsDm
aIkLUHYzqZjhqoHMdtChXz5/WO9tr4XyU450LJshig2g0JFEeO2oSv1C9EjS/OoF
vHTpdBQCZMdcLVtsWoMbjAXatYl5GLzPlC0KETBo0+vZSvHirWBgpbaRiDZgdYv1
gFbPv9hwqogrB2gCFsin5bF622zymGIsjAsZAr0nTvIHAp3p2rU+XM9MOnW62MIY
mW7fmGHwv1MDq4IAM65QWSZDAJ+8UyjlM46zMLPq9iuL0Tm3ZAIf2tqPflw2wreD
f5t5COiUJcaqPBg5nqvrp19xbWVftead2wWQCyf85mCpAjveU1C5g9tTRAFmta0x
FP85laiVqnLnfc4oq3yQtJDSaYlA8SNpoDrgIEW48mdHRSd2gRHxSDVha5tsg9py
WPr64u0GQxe3b95GBeVUniePTgm7VhZCM92HQMgncN0NLzxGuDveoMe/Xwx5XFcG
0JQEbepwdgzOJcqSUD7QvZWGtIJ2Aix440+KBtaMC3nfGqXsV7trIK8CpOVvtjQN
Wgn/iZ1bC2/Hd11/ERB0OUGAgGCVwdnkCuaMw1vGTXjAp8qzIYNrTFWJQo4dmiZP
+2BVXK2pmkNqrwUXLC0EHikb0Ju49du40GZU7KidR0TcZoH3reUAVUPctGR1+MH2
yl7AK3Ff2cuVmdSqOnFd5XOI6/R/IUOFU9GWM3F5aFDnx9GDqi0qyoBq6xT5TBmP
wRLv90zM8XG25k/nsfbgrl8IbmkwnzFiq61lkJNCKG4gkSUND+Bop7A7LQHRaC8E
1hYvXSQnJsxuiU40dtVDLXYU90yVOGTPwmaMpUONc4AQntTj/DWnvQ6tIX0xh7eS
ZsRTCclzNKpQu0DPrLZmrtTAUzNLyulZQlESGxSy7gEQ42cL4GaqipWh6oiFJ8dU
dyPrSboYqLLgEOcA1YqXQUULl7fwV219ij707a/7Rg12QYD8RUzKM7cPOTwZLIdE
Awoz75gwVtER6h8vhKbj3nXzGzRSZGf/x1LaCV7lZL+f5XS6LHKWCjew9ETRBRPJ
U3Pq7s+2Z6ZnE5FMtkFscek7QSeHGHIWgWBj79i3noFYDrsi43F/9YpsFMcpSzQO
A5J7t9puzl9DIEgSuLgJHV0ZptOhObYyXO5lCKBPQkDF4TI9MIwjnNCN39sGsSy5
+h1jE0hbGXNYt34sW2ylCFU20Ey2S0F8q4kBd/X7vlt5QLspyMlwDYf1N3+7I9Sv
QvCsupjtEyQsZGhYReOPlYyxI63E/SkVi8BVZt+uXKlUv1IWgc+Us7X8bYMzdwaV
3GOqeUhvt7nbnUEihuX8iJs5MVAcdAOkN6F7DW0bJfHdG3CdsYDyuaYgowZnBJdt
SRCVijwtYkfA4Z1VK1L9stiD9ViqJ4gNnVSl5109IuC/YOmtyj1vNd47gMW1mucU
6dNDvbV0WhSvrn60WdRwdfJQa6JHpme4HlW1Fxx2ynh7RwuGtNjlNLXGy3ji8YGq
HV3CRKa6K/kKE2UwbHhrX8GzD+3SP1MnFzD5dW7Nmrdf8dxpoA8wG1PY52hdTRZ6
W10wBmDlRw74hgjmBq+rQV/hGX1oRBPe+g9jHqIoFENUup5xj7H/gnKawZt+hvO+
dlyPeAB18PcAfK5LywfHs2RzWspNICnvuIeIWVeW0Ku+PwlCtix2R3vWst6UjJmn
HRCShSllblFNWpwO+7qhw+7WA8Q8iMNWty4Zr2fYyOjuhOP4O13m4+STcMel82yA
YgvosQiUBjKrZNavzHXOO8UbCAdcovhyduk1U3JwgiMgGWnjpUd4Inx68RtxZTsY
bEjySk3wuam8YkNzZxmDHQrQH3Ll3m2p9eorV0PBkMfV6pSSjXofOnezY0/7jjb/
Xj2O0GIqzja09fJALF0qZQHLlHviMz2M6M1WIlY8ef6oKLj6aVi5Anas26Mfoerx
lYA+ico3peO24D7t07w3KTSvtOXoXpUbjPRvkZG9BraULDjBIOKb0V2wS++UZJ+r
rw2hf5aZuAjipgU0Nk1y2kTTRSMT6wbIPWf8bwLrFZoO6zCNBQHdwScNhxkpxMXr
9ATodAZLwo+yosYNFKTD7GFjLdir0m2GRkFhxKJroxmQhLqSLfk4CbqumglOv3++
/qXE8OhVfeCTGHU121SBXHvbi7d5E7AqXaj2feetbruxhZUX1SCXYdVPJ9vA1Chz
5EVz3t18Dj1O+S6UBkMYchIy5o2ps2vZeG/SBbqjCkVTKiANi3ymmo9zyeWdABdM
a8GBc//NgFLdJKdEbpxZfpZVY446jEy0Ok/T0KksqdgWDN6qpJWpg+a25zLKuWzA
yK6vDg5hHkBXF1sfteCCC36U5fQyEHTIuStOYUgx0W/Nza6RRwBrhghdoyI5O9HH
TlfN3Hib9/pwpeWlAQYZ/H7AooW1MZArqIRLjSU1AqgC3ng89ynVCANoIpfAPOlK
Aox3Eb+CliU6Wdx9OIH6XP0V0IHYp1hmD4TpBpoiPYGNjJ/0U/d4/4v9zL65Qqfj
bFjmJyAtf3J3KtL4NRE9R0SIiL0fyZKO47v6Ya5UQpBFXNOs75myGpHRn3XEl5lj
LWRLBvVzmkElf1oR7idoK0IPq9X+6z/B4JWJxZetZV8Z9+faQruNznntxuySpvov
7LMhXsivkopN30aqNJp2pT1lJJCjHAi9/GrkQ28rM4uP9o1A7DDOzhLuATWE4/x/
ObpqEMG6a38OinMP/R8JhB0EZmrq9md4mXid4nMFipa3O5dusrDqva1QgnZUVEcG
8cKu4UKdZImE8KVFB/AercnpBUOY/PFBAJlwcujebKCNexJ6PbawkU+YsXX4ypY9
yydYZFn4iY01sOi/jBjInB2uIeZ+CRQboXSdV/oIO4eXbWJvnIeq/nOlZh2eRlb4
isfU5amE9bruQNRMQcpLbzfNoE0ZcFQZlcVsfhqv7XklI6MMXGfx6QNxgZFPDjLB
WSznkSiach4PJhlcBIbfzDG8/7/mG5G4yU61gD/bw9NzN6d+4S0Yn4b5yFc2mJ4/
kAjXdDCfVR6torawnveSk0hqdyRDTZ3WZxbqQ85GoGf+xPdfngOGlP3MN3gfW0eh
AZT3IAqEH+scZS40H/9gU5SD/RECnUdOEjQU6Uxl1sPr/jeS43CeoB3/Ruj7HHJ+
ggorgFslh8Cw6f2lA1K0lUxqWw3CcETZeYX9+WvqiZ/E03HgOHwut4SOGVB3Qo0q
3JO99iON84j7ze5nD/We44QsG/V3spm3eAjIRBIbHhueKS/OZYrYWMrkqmHqLGlc
fmeQJfobIvGSRGKASM+dGstBjPu733nM3r9e40PM1pvCN0ftqKNfdisQuZlqoDH/
hTb2mAYfhfYY0WW93C/z/wTI/n6EYbRUM7a5mbXV4uuiCqOJ8LECzEYbCjdMqUGM
e5bipOAjCf/gFWwzIXdTvDDi3xs6xYI/I/qqXrvTXdOIaJy4cF3blRZOeZvdG/sW
YJ8UVyT2UahGo+MIPPttU20tXdDu8Gvv7Vczns8nEcUqXX+vWg/e9W+lcgg5bxCA
8y/VouPA4Tu5pTKFpb93XSpMaKQZFc3wrtonJneYKTaFAw0BWW8+RY9pqcGpOpkW
mibdK7aWhyYa77J6s0eQMOH7yujbjKN+sJpyKowi9FcWVxk5HFpS2626pFOS0Bx/
uLsGPg1owELeXTsYJTr8zfUFfBm6KJePnzmlK+uCChN98Ew6rVyYTDJ+l6P28A6b
TTduANn6ipxbI6mzbv8mM27tZR9tChBlApuxfhkfgqEUjyzg/DFikloH3zLn29wi
xV9IquvBz5D6mP5rR6Ovj5p9/bMst3YjNkcDLHWex69AzSHlq40E6CLySt29KtGg
UfbWpHp9bpkaZGkdoLJJ/Su0CXxZ7gnKi2d7BJR4FZJfpMGisnkD/S1qFlBeQYQA
b4JElqw9TCygflB9+q+5cyufpJiPVKrZu54xrzatG0gn2opid1UH5Om2/+9/BVCt
g03qAROvY/O2VViHNMmuqy9LHCImSEYPvuyAY03Zx3vkfkcVkIfaSP0/RkltwDZU
4iyYdfHduscixuNY71nKCZGpd1B98P5MSR6X2vaYsaybHEcdm792LaNxPWtWuUhS
sezp52ovebyvDPxphWXr5oUz8+rZF+lv/NVccgEk7Ro2afVXrRSXa32caA2vuTBb
mRqV26iOI0m3m5/jnbyhjtk63SnoeFX3DtH/JQDnrqNKcQkO7I/d3nIqw/R5Z8dS
ybYOOPAOC0hOecfsrvKothSwGEEtywIqcuXuEL9rkV57+ukUzUEEVvvgCxdSO+dF
QHdNelVtd8W3XYPOW5clXqN5JvehJ2j2iYcjVEV/I3DZaFITA5qqNyhNKSTHjvxj
oK0W6hlcvoJjSBtGdHbrOWKWUASQNDwZqUiiUguIuACzdqx1ftRUT9BFqhkJ+MEj
s4AHMOJLc8UnNl+MlHC2RipX4CIVKNBkDUiU3bSYAaqhwlq1O8plbaMbROjY+DOx
ETlo4t1sHIt/i7GaArhOz/EFUOFc6PnRLFUetCoImZb7ac5p6xoKa0QrtvEtg7BC
oeBqO1vrfPdYKeqSBlkc4QRh9XjaFEtI/sj6v3ENcs2V+K0zQT8PBX8QUfQN8hs3
q2Vx9s7StFRkcqxLBAF5pMK1Ft4SXVKw7vTRqU2pwyvOfsxWxUT8j3t0bPTP5Gv7
iFYQkkCbIyA7JJ+HFXBboF+sm1bgVTYTUotx4eoaly3jXxDKgVYz6m/7tWWTE6g+
doDfbgH4G5ZsOhcwAheSBBb5clEefquL/tr1aq3eSe0V8+1qPYh5KeSwbMKmY1Qw
pUiGxXOE18xYtaTU4aYTeB7Hy8wtuepQnw/D+1vrYTtYr7aFEF/3/axJG646sN64
ZW6Jkq4fkPpndN3gqoYcgXwoOgZwV/BIfPKq74j2TSNDLh2hNjixJUZFMpuG+LU6
0xXpe+1G6FBGfjhjinYGdI/Korhz3TZXD1dkhAQRg1oXArAO8TekBH40NFxRdN93
AAAeifQK1yxrpKAJrjRJQAQdkBx1yjKpyIK3CNB2BinKOdcVRwgOz1k7uEO36aIw
PBQqn2VBKjVXuHQ51LAEnnVBBs02dsZnHOgRWf7VMaJ5Zq0soTGcmvfwFjchj+AF
XFaBZ/T9h8R75X/wdnqs01Vm6rJAYQ8uqcmBUhkGQpM1R4lb7m/CCIfEHMsRj8Cv
+nXVemomRpnHmuorTE95DX4Gfm987962fz7J/ILQAjoSnRkdi8IcBteqzTbptrs5
zjbdy6tssX/G/pgMffdcsluIlAR/pc2b5jZEVsn3HCNgUGf/F2OpnHOe8Dsy619A
Ms3XIn014u4HMVN9HSHFX8Y6j8gLIbXRo9X6s4DaICF96yD4MjPJ7Yn+Thwn/Kmf
swFUrfz+N1bFW4NnIuGofj7PVI9jlpvCLEsZlzebuz+4nB5w81XjZ65iicQcYUQQ
fh0EXHqIAnFzNKkomfmgoNC4cjuLuMl3qBNdw+X9nWzHcPL2K3j8GyTt08ip9na+
gMcjhhwVCdG6AmG7qMCnGlOT/miJ2Ki4uEjVdZ6/0rOxVqO/Fhu/NLk1TBC6Ncr3
3k3CQlOt08HjHnzd003qaesjHIrtkpK41ekD+zQhvTXoxpgJ+mVwIbQw5IrIRmAP
FU63S5AoUUNx9vVHKDpWhn063HAWRkvjSqnpAbrk2Z15IF5YBQtQ42nUtKuOw6/u
04OF48uUqN2Et6R9bnanaAOUMViOgmlrUfazMEmgnvbmZCQ9dLCPjVmXy6gZqm6C
tVjatBQTrjMwUyMCFy8LnXdRqrSGptoCzAVoKyfaxVTqBH6gwbqWXXDg+C/fDSi6
+NEdQAuWenOtyiorPA6w7up7xo74iTxghoaZzyXdEF8UgQp2Dg5pNWo9JeplLao9
Mj+Ze5YyaJtjUMrA17ZEJj5NeY8rPf5khir8UfQOUUEusg3MTymr18lrHynjw8V4
S60NdTBzRk15E5VA7/hKfR0a4GNNli0T5g0UwIgZzEAZeNWdeAN1ILfcccGoZ8zO
ZLOVgNqlAgXGOiXI+Fow6NiM4a8FqYFREp0T7xf+LtXLHdCszGdUeq6KmpbeIVKa
AJMJyzPlhYf6qSlM06RIbtECLKqGuFfMToxqliMFkN3QMpJTy0NZNyb65L5g3R39
7EWHfEFPFKHi1CoF7Dz0M8QFV+keGN7dLA7b+K2CcXFQFX6M1Wzf6zN0T0kHT0QJ
XqsF7ZeSCjKyB0o9NIRDL8fz32ILoFHE1BmZl1eZ3kf/+K35wa0obvpfQGpDmxx9
R4q6Nc2sESjE/jzfdZsbhil3o8B/i8Wj13A9pK6pU3Xq7dyYLfVGxFGg7Bu2iWYz
K8O3DWdGh4neXsIzIt5SpJMne4v0R+OXgob0I8xuSwGz5yx9k5MXrk1Vi4rFi7Lm
/iqa8FLCnoNslnqQ3XnLUQY4/b8SjF0oqw9vZI2cEuwsAKHqmw6s+2Nr9rYrq+6p
iNkNXRASWLHyJmfc+VrUjCUfSYL8asvzeWZzWUN/zttE2lhb6kVhg2JA6cKdWly1
hwmeAsbfhoNH87T4VsTy8OMOjP+GEbPnweppzQU+/n3tUHJ73+hJVy9CrFxK7K9+
CnomXqaJuutHa9E46QqN5iqaOlflqosx4o9ozObZjp0v9ikHKzyNLlwtYod3ene1
ySLexvMr2H6whEEcZREnyEiXVstqSXAGBZSWncB5lZku1cwVZC1k0eA4kc8bbTPy
T/E3T8JsH6nKv1U72I1USe9lfeOX5rkABXL4ZOVnwpnBgTi3amBmVqOAEU/dgLe5
ymk0f/fkNUXEjcVZHNdjrb/8FLGYkpxCyxscf6V/ke4aGtdYxhIq7E/fIIJvA79U
ZCXaDBfn02Vx8HLbWQgMTu4/gcXby/xhSc5DNNRqOBGCD1NYMhQfIjkgZsTp0UBq
JDUai9YHxniOslb7gzYZ3tS4kzq6FnSDgip9dlGTdBxoAGqirs7qgc7OnxbaaA0f
ivLeY80jBcgigDl0KZXZp2Vpoq/eDmpudfjy+rtQQqfgVng1Bk/CyyQBomQW2Peg
DwVXpfb840okv9uTE0LuIMvKP98J4jWn/1xwWCGtCgI3JZThCrsJSzSIyilic3o7
HtanY1oj6fysl40GqTfZMKxPthUB2NWc3ZCvVhLJnGV88sgWAC+6P0eU8F4i2K1N
t0FbTDhVpgCfaQxKccah2JbpnKDLFAdjaWqKQUZbl5vf1EBhPS/kubplnMr7CZeM
1hUM2MwS1uvI5h9PAIqcwRkcb9gzUsUgLI9Z2g/J9ZwJoyy0ZjbSgtcqwhr4JiYc
Eg7/oD3SOHJu0Rsa+KsaicCHIjAcnhaN+p7LwRfLl6Ht12sTBiMB944aFDrohUR7
c8VaY8XU0ZXweXJoiwCJitvln2A+LATBZmpLJYojePjUXpL9zFbFJ+6JVC450eBy
0fUf5wFtw7b5kKNeqo23b5cJPR8nK1gS4tiaSoLuTYHcrPuLqtO0iFN5hKm4mjtH
QDExPIFUEOXjba3H7l9A7sjU4CjKtelp7nEHdmcU6MB1lUx8g2bDRGRU6D41PK2e
b/GboAe5cjKXCdNQIlH0cp/kjmRtwb0zWl1ZMlPxJfjWpK8itvaltCrd6QpRN6Al
h/8FNYk1O6xpQ+1n/ybsjxIpB0QQE4N2zQuqaaiHhxB4SH5cuHMJIays95ngJtB1
xBmn6garqYQqszkJavVww6onoJwFLq3sspo6F3kFPGjKL/tKgkksUs1ISCRhCuou
cepE+x2mhN1pfImulCK2IVUU6zyyOqnDnTgiqDZUzfaD8MwYefCz623cINcBbTsD
mfHT+2IjJwobcrmxiLRYwMXsaFStn+naEUWCQbDOWa4TPMD1qeieOzoz3IsdzuwI
o0DsK+MYXQkWO5tmlibcuYpdrtYIhtXOF791ovgT1h/JVrVadNGG+Qt0GevkZFeg
rmambN0hcDtaHv4Vkv1SegX7CR20zQKIDs28Mi5PXCwM1GmqjBBsqjgTyZBVgffZ
jSI0nVYpWSzoLvi/+rR5RQEmM0MEdjuMgWVzCl5I+X6jZEBb8kcRUDT1CY7k/XUL
tW6EUYjDYpqR6cB/iQ+18XbXWWZUh2nojLFlHt1y6cyxYNR9s8Uw4NpM9kjiXB82
agaJd1cQO9PYh8hFF/qWjIMlnjnr2HDBHkTxnSItrJTGkduyCh0lzBziGOjifWn+
gKFrY3z2N98bq2SWV6Ny+xRb5kFfwLE+dVFKIFWNtVFMxaZmeqtcfsF2MjLruEH7
rz5f/JUW9brDfUPGvT0UQeAjO+XxPzn8P3tIsmBkRQQRnCxhyxZgWAhwdkMKyLr9
CV6TvOxyO47Bh9N+EJGW9Vfszxr9RfSJD2ZFHgmmxRCYmpGZOaMROoy7vtXUHwyc
6aFHNtgbTCpxtjy2BjErScI7eoinuJH68TDzBeZMp8dZSgEP7WLZD8Vv+inuwim3
VUJKQb5PQygdJsG05mKs5T49gjMRPghnmX2O0CqbOxs7XfUIt/r0Xt5cYctAxrUw
dZODRu8SeL4Crv2Rv7Vcp2xP6kY5B1VXWqeNaOPZnfFFmOlxyqE+7QRmjCaeEXk8
kTYUvkI5OIDM/U9VAHUh24PNwrehlJWao/JesAp9a/RqIESQPmDrgoTR8RrgRC6v
nvpI/CVvUQlIRgFLnVUkNZcmx4v/hNbu1uX/KQO32liYQz6AIKfVbNh8TDr28QRx
3d1mGo9JovkpX4ZCquRPSWv69NtDt6RJ7cPRNHrO3Yrrw6Z9TYPOfH3J8q5Sxqgh
mAOhTTQ1hWCKrxubkjKB82uTV/zR+XLHk9eZQwHdvvHo0uFJA+YSDB9Qd7hn9Ma4
EHEYEy6Me64STSCnxlA7g3CaR/CmMUIEU3g4pw+ruWOE8UUJ3wQNUPO7I2pYbq0o
wayRY4AT+wSEGAv3llCrgHquG63tjMnYCQSV2cLeFGzgl0/VukQbRsGfwEIHclBs
j0hxcstPvGQVdftaFRgXHoYVQKRV+EifdENFnyWLQxct/Q5Gnrmtj8HfqevHzEME
9Xb2Hof1gltG0gRVbExDPqN8rKubY5HzLlOC8T8GobZdQx7oWKGoYE/IJI9ut6/k
72gGCeIQQv1DNNGUPp7L7r2miUYLpBS2cmeXlvQfx3mFPCgU7adLapOMTW9aDTec
vVljSrZrcddkaDNE/LxDnfPfUlpEDVdJa9ckL7ZGAOOupQjN8eJjS4iMPAoCLITf
Vi7X1TWsFm+UYHEpIREIOriqT2CkMMshy4nNq2FToGJMJpMsw7x5QrscInHD+j0b
gwxRCl6FJOF2gBtYSqFVHbeHbKM0f5F8on4WrxgY9owvtI8d0yEKBpUWTy9J/KrB
f5qkqro/Q9hS/5HfWYgo3nmuhGqxxvGR7O24k/sF5HdrFViwEYEAHmf+JuibYHiS
uTpl6e70cm/FtlSphOSkJ5z7hnce9rG8MrsMvJA0Ev4qudVeH0DgfzEQNUA3yd8X
WUYZ0PNYR8EhmO3nSUUd7XCUJ2hnxuesCXAJAa/xUygTOJUrXexhAkaU26+bUiQW
yzjwrfAj2hsR4tMM04t8AEX11X9mK9xgwP7DNsnpm1Eu/oTQrQ3DoI9nEAALjLdl
0hj8A93Ft6FdwOerpSWA3T97X+1DNdVt0a897NF/q1zEg72kpz4/bZworWnDWYKE
756A9o8o5BODVWVV+oBKxPLl911KoqzSlk8YfEJAOJ0YaGswT5nVT3Xec//UUaUT
yMkaU5tpv+c3/pf6o1TYN6aSYeEnnjLz7i/hpz5Igfdf1Xp81jI2bDZ2bJlrmurk
s8jBZqERVX+0SbgdDw7WNmeNtAPNxUydnwxtSt6JiMy9wSUuW09KA8TYB4+219e1
V2H1jNEt2/mTNvlCgXp6NhFRRunEZ0CAmB2k2EACe1AynfTlb6XsXsobUWrxBUy+
O7iU2WrRqfQSTcTTtKjd6xgjywsB8pdP+O1nfzhTlNR6X2JEb3aCN0LW9EoLNF0G
GBa6BW8t+7rQM6WA302sn7OByyIa7C0VZcp6nalVQB0Bq3dE8fO8g1hqKqNlVe+J
C3yZBGwm9891wZnUfRtl0Ii1x/nzs1HmZ+wNEK355PHCy44iRL7RvJCA+oLHmw0o
1rB2zY6OisxhBW6XwnRB8mI8cZC/N37drqp3Ix4HD24ixqwIIDh8NH9iAZPrSTs7
sJpV2Nsn37SPa091s+0ihUtyoMsB/BycbxsVe/+hfOElr3Y9pa4WQACTf+K1g9gt
e/WColQWZtcEvaEViwh1rt3Av65sTnc/udn4tNHfwFjbUuECwTZ3eZwPwtBsBhdN
2HAk+wWUNIMGvZ3X4pPoPAtvfWEALs5Chm7TAYqDW/RA6FLiATRUKSEE5BL6lGSO
FUH+MXTuIH3EfquMIMbyWXnQGBOtTDv4Kt5Mhs8iNRpyg57eNppc7+m2AZTL7klV
+v84yPb1GP7T0Tj/Qs1AzYAaIu0Ip6UxE8sAXOMVA8CGuVMkMA3rcDq3c9Vwi+5i
J6UnhoK7+pEvnzYAIHRnSqecgY+cs+PrjXHUYKyoFfMkSZ3m5uKdflle3CUHgg6b
3CW1a3BGA4OGEXE7zeV8Bu2bzATLVdq4eGjWB29YjaF0F66pwWVx4ySxfiYTr87A
+EFPOCD44kFCvr++ByB8mKkccKFHb/AzY62tGy/Q9fyAuUZgIv+meW74GoDubu1z
VeWWTISc4kL85TlKLS10QULgvF7P6A0Y8tRLXezOIUlp6RqiUk4f8dAfIom1ucZD
t8IALjrSk+LsIKCcSoV6z/yZtDsa9h5hE9ll80KN94mVZOUh1jMhcqDODK7cX4xk
5rY5FEmMZkxDXwFPjuUTY598tIJUSkYNJORncsFOxwLFIgcwUXmyeLLT0jtrmCGM
D6b1xBntAHXiBqA75f1qdYjOpP0VlViQnEL3A3NstpoE4BMSGeXCRn0WPSZNbyjs
JhZM6Mgfy1LUnn2IIRWdF71HgZhvYFTi+XTpfKhfT6pctbwxm3Vjs7sBWUR1Ecrx
qMoMkXjxM+pbfkMrMIOa7bLFaBYqx1/64SE1MYMhPmKwWKeRBmw4qq2OSQBomvV5
DWfjOSRc63vNVYagHWcLRlr7JZOhqTPnPQYCq3xoMWGFVthWPL8WKD6dtKyrALBh
2xqufvxbi+rugjcayhvH735W8HVBYiyciETvtPRobrpI6FZEQn0jPxmbin3gGPzx
G5owCJ090QDJZ638MFJepyGsd6BnTs8lmBKPqND4miZHpgMsXYwcRo2RcL4SUwi8
/F1CrffcmA7F6FL2iRdc5v060hYW92qrmtVvpSlnHPiKBt0jZp0OoNDWSOy3ZJR0
4+pFN49naeUoXNvA/2lkerXnBNMGzRX/s8ul5ROMQUCj434+E/Ohoi9ngl2p38Wg
02yZZceIWNf9o1lXw908aJ4bRqj0SS9+kViyXdTl1+E+dJ47PAGVD+jBdMqUYjNC
USPqHitHU6cqHAKInjc6Na8emLKJ/RJ4f+Gi0Gl2d4dhnOq3UJRH7H1rl2xy4HMf
XtLTkQLSExagxfLbD+W5mIsceOd0ISnYeDP97L6yDFeqlPn6owGmQ4ks62MepcJR
aqSvzJkSYPEhNbw3nbNnYqf/qWgpXGPK6MXIgRBQ8WSF6DjlAdZqWJ3MXaCbevPU
emraVAIjpSXVVTKWydttldAZizEpp6llIpfb8kcjjdejWUfmtcrB8ZgeXYrUP4/R
oVEnMtWt+wDE1brgVixcpq0PjAQR5r19qtexq1VBJTuTyTwg1YBq2u+/egT9dMNH
nZyirGd2HFvn1lRBUqD+pR0Ou0FoZ+lRNhKc1vpG65meaQEEF1wWQ/C8ZFxJ0RmD
7V1unSKFcRkrB5u2miXGHtGz6mkl4d0WGxQKiEwZebELZzYzjXX5pW9WFQow353e
pBxT5EGUD31atQJlCK4OYQ7Mssjlsvrwxkwiyo/bwfBduuGNpkfNWcaHHsGzwPGZ
AEwrQaTHSilbkD3p9uaSZeQyaxLSbvk5AzJEh0Mt6n6uPYyuiozas64OL5l96Mud
SyDXH/XDtW4nVrfNLtXCGL5hX05z2GsfC8y+SzBZFNFakItKOzawlSswKYAvWpLj
9gE57H9zd8ZwJpPs0gCm3WxvB0O+1GnLJYXKQFPTYP90TfSZbuu95RviJuRO6dLI
6jp6b9hx03cNaDJ/uaEWQxsIsZdg54ZeJRLUmsret0MA+VrYIHRStI5axADE2rTm
BCGM7U/BjKcx5VZsMbG2bT6CHsj0t7N2cwqSMI7iT9Ftihvi/Yz083hK26y1s/w6
d0JeGdbic+V3DObhbOnqqQvT+GSsE+4mQBKFJMvIzTjYSNVJoYEdvigGtykD+Gnb
w/3Y43nEQj+1ZCVDYrC1Bi7aJa8tsVf0GV2erb+88Fb9qcn4joq9LNhOuIWuiKdg
M3IpIt7TarZP2iRkKsMpmO8PhJUbnyudFp3BaUW16as7ap+AnUUuPbVhgurJ+5Fq
H+3ZOpkLYeInJBaL6FVUyG90mWk1kjCJMd6oJMLwN9wCWH14VN1ThVu3ngu6tW0V
hNyPnSifQozCg1hGk+NmeA7PUVzxJgm877TYg284+GGnnIn6ehv8N+h49dNMNeBi
8FDTiWQqWjBSPcqbYRqp1GUu333l69MdVciSD/HU8sInY40ryepgzXM4pyWj2U4/
h82+wGlwa7hNfHfYcSDKcPtRSBlhvSzjP2n5roRbWWPtyesL7l9ldemkd8km2rw7
nsuiEjNMiZ5FFU7Y+D8emnwCAnm3gl7jgporCs+L3v1tTwDpivHqH938rWRJ4f/o
sba2E4JnB7VGrs96JXtvZbEmJZcsncWYySUvee0DZoBobmwNzAEf4jYUlakDnbw9
QnoSAUH5oCd9EEgOLUu5ho2gMshXYONLSQZI6SsZfLLFs0lJhriADbb28vdIpBrc
id5TgBW4acgqKxY42tMMOtGMbpMWzSHz2MaCIaMNCBKl+/b6r9VCmyOKf2J7Q4nL
5BBR/3jgQ8uXrWGH1PN3Udc+9uq8edybSsaGViusbxShHXkTDoU279T05EsiVU5Z
de04laOnEtSg5iN90lp1B1k62giujZsPet1TMY8jSj7zRmMct0GsZM+ZbH+GE0po
YIzAz92MucgP61FcmXyfZBa0gPMbm+2oOlHqwwdEvnqMVw8Lg2gzlhEXud4JAj0E
wHVMoEDEaBuX3dQg1RHhoiwDLHcDTwVhvUtx7v6dWo3OLwmBnEJ1Lu0vVyoPfqNf
GdE1NJR/9UBO+p4TSjxC+186Nzrn0bdmF5/OfcdED7+Kym31qLS2W0Q++MOYp+VN
JlEms+ZGD90nKYtfqaAATvG3WsahkMYDfXQsDzDVVaCapgDVJITABKxK4/KO7Z37
8nXvBIDXqs5hpJDMb4Vierj2eTe26ugOKGmWGycCeA9YEph7e5ruJm88HaH0koyf
J1Vf20tSOniylaJ7JjKDsHobPUz6vpN3CCMp7Qbgh/9ot4Ap7owDrh+KGNXrTjqN
TVhTUVOVwAbf2PIZsHR4SJUemMc3VRzt+7QGVnpbFpBuBUgrEkRFf0va+5j/ruMM
gGpDxH78xUsrARrgJWolgjrH5XVzcB0umEmfyfmjGtT5cGBCJ3+ys4pApoqa2egr
1YemNi2XEyXJjFS+KeMamSDZF4GrDvhaPKHxBRiuJYi8fqEUG7PMYOXikmvk8cX1
wXcZ65dCAAX+/cuczKwutmpb8jccx477vzbiUzBCfti/fxOTrU2xZ1HZxldSsL/k
QxUoC+TSio1GGGSwUK7YDw+8j6FH11MdTtNU9If8pSIoFVD8BzRZEXidCSIsKer2
y1bgekZLWRaEtT3FRwciXzskAfEuAS3sivQxRzJPmmh+ZBg7qFtq0h2kqwoTMAOZ
2Jpl44eqhsYqvCpUrtxwSdR16gpyYRuIyRwr3uyXYCojWnn2COuv+LShYVSiXzSK
K3kKO0orGoIBGd8Y+SQ81VjYoubeLzAUWhzvEKFJRS2aGjPxQ1JAEclu2l/cUuRq
R0mMYB+uP5X/B5tvMa4pGKE4Ey5sK2zbHZB+dkh9fTziMqnKvI2dKeitXbv9OoxJ
+lGS1J8RDjggrpxM3DepomOI49+o+wGMmVz7JrSploqmjpl+VJGjTpiTKbDg5qWw
dXzPOUJ/zd+kSVKbF3QDUnMCKJ1bJrTJqaIsoNrrpPTvP318Ht95Zs3YSgNgMWoC
l+avd4b0vy0sLEC8BYZcabdDDAVbTgvXNAhACN6L0/dl+KdlgDFjlhJIrCMUb6Vr
OCJvn7l8ymGE/Sap25EopPdp+d5xIml2hFRHw3/mSA0AuOwuoNzlVRfBvp+cuwbL
rTjzQCW1KhN2Gqk69Lg5biW8ndzYrH78KSJCLO/prP6F3S6GjmMeyrpk8FsloCTd
YoTuvn3qEPoNz76e2AoTKYaY/KgLwpsJ6RcB2rrojqb7hvBNsMBdLal4vZHx80MR
ykdawMAwaStlwQyksHuYEBnLR5+BZ00vYEOETjN2BQO9L/F0k4p9r5B5EJ3OJZjx
403kHMU5lWl4+KCSg0rNgtsxxa6EJwa4z3hjSZNfH8G/OXDsYhq1XjMuXR7Vu5it
ZO1KYmTteQHs4ALHGq0/1U6q+QrDUrr2z2fpnpivu6RdV0FW7L7nQBrM4fXSrjWx
bJ4kmTHo3YjlMrGwxSy/Z4N5Wz6wxvwP98TlFA/TNKuxmOeL0bf3P6MNEHx13Vkw
HOp+/d1X0HFWVUXaKewKS9OAu/7OVggwmLxV5/vFNjT1Z9NcfK2i8B/sEz6oeRU2
S9Rk7cjgBemCb7FlgA9gbZewrdG1sMAmrI9tk6kwahS12736Vd1DQWbty5y0BGz+
j6vV1kxIBgYjTi+AjHO5QbL7CMefwNxqPumMRJOuyzBlrn71W07IlCswVbHFb3P+
SnZ8YnNLddQEE46lCcrteWwTrFroyJeAmYtOt2pr/gNH0QxpCMHh14WaF5QiANGl
/OUekKU/A49QDEDIsW+gZy8e8+vIYFyz2zmb28Pl5OgGwZWynVgXooa1yKELUXHs
POk+zBav7HP7F+k9/Uh38VlkqHwz1BP6qsukhmxHce+yL5NSAJnHLeSWcbifl1Kq
TPjJiIz4k/cpMSb3prNDdygpxXfDJLzgcll2eRoGgZdc/xyBlNKMINcJUNURKUcc
LeOWS+n0H2AsnePU1L5cri5LUmdAli8RW+RXowHkrCNSQoNKyJIdSaGL3c1h2fT9
VbojoVLVyPmHwmuI1coK1b5kkTyohuyDovJoAfOLDOmgnUnx72DdW56MADHjJkkZ
7jQJjY1pIBUaZbtpsmPITaoNXD6/0yl6vpNHBmNcmEx9qbkdeJT9G/lsOZ6iJH5O
tfMMv/MATLDCbLMpiLSOnjxrLDl1kmLj02Q9Y20P3qLnk+jRjigSwSGiQhlIi7Wl
x+c3w5Y9lqHsgMISE5E7kY9mm8nizMxLN8QdoL1ppS5cUFWp7hkYrZc9me9VlSYm
GwKrmqtAzrUjYNlLaUTX/vPHiAODzck8ctJkCuWpW7wcMx9hd3oxwze0+HerluLn
8+f/sqf289cre6Sz6FRFc5HnOPu21wT+sszxslirYoc95Gxblr5gFt1QoH1bI31N
C+QV4MGLxue5sEXTeTHTlMjiKfVeFTUtHHSPSsyyjq+t6SLFJEhDCgK72g562OPt
M+FM4EZX8hPqxFuxU0XB5wwT0YP2tiKW2P33xLu2iCYEKpfh6uqJdCHjpxeGpeFP
v1MpTDMNG6zE4LFQ+acJVW1BRbH4v/VFA/OxD56OLls5baQRE8XtMys1M2BkZECZ
/uKpUu73ITQnmucVAlv1+ntLN/c/hTgFAUP/dBONnnbBIM8EvHotjKoAyMVKmXCN
C/6yGuwF73NO9NRv//UgQIDs50oGLPI0NFAqfuGjHBN1hZjfLaEMlVMoGhOLyQq5
PlV9zFFpbX3rywwBgjjkMoCmfOJ+4mUDQyvRUWV0nncg3VAaAmhrihD4iqv9CCGt
y/jyT/lOcOzoONrlLsXAMxlM2r9DIp6NdnKSIldzQdDNa6PpAvn7ZCmvsUpvTH2u
hH8POkEkj6uzbnNxRoNRSWPMlEFfElMP57VUBWz+LQ63o+UBOYnye3ewAQ+798yS
PZzyVTAKtPJ/0X1sd1StpUckD/A8oK7Jv2wH2NaKDWrxPT7CrHf1dFJrtn2jlXB1
Ms5qJZjsftWzPosqBEibNcgaag7JVJ1cnQR786BKEN8ZqTXQiImWE8t/RsFDOeM0
Zk4enENj8Rkp8EdQxCTHxtKmFhcjAoED2hxHWERrBGvof8yX+BZtRd3XxoIGyBg4
T0aeVXz2qbUUBZoadMrdPno2cYLNsRbTnKGixAFHbzahzVhjKjHwGDsQDewqZK6o
Vgii4UzZ45av9Wjbqc8+HZXY7mOmmSvm1ulyhzfYT4eflRIGU7w5z4uYspTqgoLu
3tL7zOD5DhMUjp9XQewMapeDtHxCJS8sQdKsXwkbPbQiHH6y7rMQbNks1Bd3qzaT
nOe3WpUDdScTHYwYG697cPAKEypfT2ZyKOzcpVfTVBM4Lzv65gaqK5G2CFKF3/vb
ODGkFpDhEHzC5fHTwoT/jaCCxGbwihrhlg5h+IWtLUw2yzYq3Scp9jRpOt/pmeXC
JVeZs79k0hXYC6QoKVioTLkZ9TIjHneL+mdk8mkeWk9IVvzlppsTqC/BBFNLx4r4
cRuc/5IJek5hEestFKysgiN+IqAg5L/r7ShB881Jykiy8rAMq6rQds4P8zmTZbIs
yXx5WaihF0FsT5+iLXiDZ55p3H4NC15SQuZf+K2BIWuE41UeDflQRvuMJXpx0SIU
x7HzAG23XyMPIkFpo6Gfp77kwAFkenbjnaRFpdQ04rJlkCNUqBVVoIR4teGvXvRo
Oi6/ahRoYRhhhyp3a81DoT03Jp6f3FaT7CRVr3KJPybXfrKhO3Zw0k+Y0SAbSdrH
83GB9LF3arjrOeEuZpzbSLEpf5msnQsehegQ4/wKPIT09ZTgJJOuDItlnVMl+MiW
RVVzrbSWeBc6vpTY6lLr4rJdGeQ9UvyalT6sIw5WiSoDM0+oX15fs1BqK6fqeHuI
CgN8CpSAe3XRzUPss4vOvUtwKdK5zpBcxUE7oDymweEV/n7rVjlYM43C15r9a+Yw
w+Lahyna2Sds5rSzUStCPTy646hu7Src4P1TPeI2+pKdAjxOngAKf0yKQZZVMEjh
0oFNSVuWA0tQpLWi4DXJck7st2I3QPloY8uwcsv+4BJ95l5/TNJNI2sYIt7DRMm1
aIlKLcwTt+Y+mphR6EjOcp8e909FBu8CHl9p8S4B2gaPItNlwHrJEznKZZgG5OTY
5SMFTaImT1HOoX+qORxexvip7M1dj6lXEThIGyTPvD25lfPJF9ooMk4APGJJJAhe
MZ0JBYQ7jM+Ii39hxfFzFAQtBVueoe7CgXci9zHpSybOuFpMri3LUjLwsYfFdYTN
4afl4PAvH9N0ngh6tx5vFCyhHmHOBIgLztUOJbAItqDbDXdkhVrBwlDssz1MnhXi
r4nu0PX/iibK3wAer7Lfuyhnvt+3lvGii9cmbXWhHzg0hOCJ3VKEmMSxvQ9+Mizi
L0DWpYebPRw2fF2LXyAX9lHxbnuKSg4auV9+Ygf1IwLKJS3IfHY6NKZSra4WbOJ8
Csy3NDmUDmX+MckXKvqF5Zj6N191xqNGd0euqR/G67l/egWrFhaofJ8tRl7uwtCP
MI4wiRVEKxacG8GcDq3uV99a+0RmXWssys6RZEdrHaqBFPzdwCPN5j4PTNXChqZe
9OxoSXwltKn+pfwTX8Gh6Hf+LRSK0BXw4tJbK/lMb7PPwXLBZ2oGht5YrWTWre+N
g6yyJ9FR8Tiwch/N2w8l5LQgcl1stovXZbKr38kq5MXZiv1AyWFbGB6mw53j8rgF
CiVSwPFs4/PMjOySh0L8UJTZtYpo6eARp134wC4EG/tTYXM663nsAywHSaQshhMY
nxIIzGgHZLSQ0CwM1p+bzexJ2H2SlJqNpz1G9dKephYXp4DDTtnM6YTAveOshCcO
dZFjapVgziv7sN98ch+zlNLjNiohHHB4AHvfX8yDvEbFXN5CBDwucpd3bbez1rzH
0SAbkYqD5VQzijzCxpsVraWyCkT9OUWUW1wTPRdoLeKnDfXNXYMg0MAcZ8rbJsjn
CxReu73Y9MDVHwAlm7RnYO1HGCR0nvC+YklBBWuedTmTXlat6piEPVwU8Z61IGfD
J3IoyVrV7uemAt/8xa+xVAGPLFDKh+68Cn37o7NxA/UwBIj/Jk9eHCoCXsnOBCPo
L3pnsBE86PeVSkQf+k3+R1fJCXAJstArn2P9RlEAKW6ZwcmAQoFMMjIzULILmCif
YF6/w2Q64SBqObVMoCjFVQK6ggDmxvyYiRg0EDma5ceyjDRwBvdP0U8cmU4FY4JA
zLI6OyzkeF9Dyf3qZb41zWISwCONN4XCwX1D0X62J21YDloFdBHLNDu167DNGNw4
dNdHmP27zmQr44m4SmfgWuXewSa2SFNK1qmXGALvPtKd72xZ/XAtHOsSWj5TZIZ+
Kz6bR9Z+lM1k4rRBJt1hicxr+Hx4oBrdXKzKOv1sP7zfLVz2BIgiPhd2Jllk8AY/
VJ0ix/e3GtECMhEYG24UujqsBe1WvRBAcsbiC1VDHMqzf/kMvByVhvNwicVpj54k
2JAR3N+BLgMaQivUYhaNLOWkXtGY8LdEkwZW6YcnxpE23WJK95NRzOsYjQPgC4SW
wGNOVCmjtaTHHhCFkLFX+eNa2cbTjM/oCjSvuFXu2rDmmtzBX1iG724HfcKeKlqs
PiaGMFLWaj7L5ejgBQ35nDiDOiw+hXolpVcguG78sqlPyVoNtMFIw75DfOKdDMaH
fY0LGhL5flRwnfgBiUAyfE8JSwvjXZ/BrhCZhUZ67eOmEMcpkUu9HaGQxOZiphP7
YB6useMGjEzefoz2TIihremarpCXLazZHME2/83p67H0W6fNb5awVqKLuzHYDLWy
SKRUDIauUOwq+dSsLJlWHU16RCE4hD/ytW/CVaMEDiTIzC+Z3SAOlhcNtpNEeEuD
nyGmOg+MSWrYnK9Z8I8FrM0JZkyDwARytwGu5dy3BRhyzDMm1rgGq/OCbaGRRJE9
rh8NAmFK8Nsst/uw5tWPW9w5IIe2ai9tWgxweC1jYescvC61FH9PDiYfJjLavg15
5Kk2fZEmnj9rp5eXoLvXcvz32UY6F7DBIoHevTugQedd1rhDMyCOYSF/2/PeJf6m
xsnSZiHLuZjo0e6gRIZ6r2QDswkYAg5bbS6+Fg2+Kn7ejBxHIvVpHc2tqk3wX2pp
IOxcsRJRIHXLiUyXzyQOa1V0KNp38nrhRxKlzGl3jGvDGwJxL34+AxYdzEvop12d
emQCLvqrBsRHArLch3R/BdZdnS7IICYons37fwyr6hKe5KbJ+Ns5UpcDcLTyQczV
pHM2JDNw2+RneaeniWRnwAoJCm0oObKhn6Ctj1PFtrgQNG/SMlN6L2IwpMQ0UWSK
jVUQ4dTdbcoknVO7sSTODTuHkTbv68/oUHmNJ55oWLdmFIvcTsEtdqYoopD9wF9l
Aa46k50FcVcZwFNjcwY+/f9s0mommfmv+pSwoMdbahi4j3XrtEdu4lk2jG4YWb1P
ga3qA3BgsIYkUQDpZniUrWtFj4dDNJTjKG/eZ4c031o32zzP+UNHOBQHPuOFKMTQ
DNYcI9O4mRPfxJjhjHFriHfpir6AOBNCjL/6ZRAfVHldQKJTMh4YAI+4Z1sj9P70
UjHnX7N1Z+7FIuktYMivxUQ+LXJf89PspHIEkTgN5yFKfSgoZkz+TbmmYLhHVToz
tEUd8F4skfJdx+WEEik+NKC+sYvCjEC9ny2g0BGMEaA8zU/WjGRUgchtGJTyNZYu
44T6Thgdj3H/Za3gVzsSrxk7IxNIjpp5Q1fPk2h3++Y5ZwVoCk+LxXbT/g1TGKbu
coPWyMO3qDkH2HDqRTxpKi9Vyf7spoIAwxMRnXzc9Rf8UYQSeWz6v/5pHt21MjmQ
6yMQq8WfqK7io3pJ/FLxPBLRkcCqLXiHMRI16BaR9YzYjZ2IGEX/DTrta8nayIJS
xGTiutRNrADJbX6JXN0YjbHfLPozPFCvbi2HEI4+nVmPzyf6mN0DUd5eq6T+vOUy
q6giK3WOp3czw0rZAk8gX5K/6FEaTOajwQbDXGVT+zQz/5f4P0RmWXCDXDsh8Tgp
yNhUn7kCx9GhzgHPXCkSu9o1w9sDTdlAKeKOSHB0p3Btj+omq3fQDb05FeqGGZVc
KEIfFsUC3WID483vFQAU/Dn4MpmmWMy7I/msncGVkMEowLifml9/UD2bCkpyGh09
wYzWrfecg65DGFVw6zn/H3rCahd3HGkOkBpHUq6JBuo91wrwi8MgRE53PSMmpMA0
7dV6h3Y6h2GonX103EsrKQg1u2KR2qEkZFixKfqLwbwf3r+PfcoScOuU+0XqqNGL
zMhZSebGNtYipB95v0mPZ0njCLu/0NPyBkGfra3phO6cV4S67Qde3JdsNlDd6vZv
kHSL60av3XksWuvTa+wyr2zZ95UA8lF0HRCiY4jZ34wVBSLV7dCmC7gvRX8zSUfE
GSJ7VC/F4a8F07WMLfaKqdKSlxnEKH96+HQ0JsLx0eXCiPaXspbNuZdjzOoOnlwC
2lH6qb0ZxZ3GjOp80bkH7uAG7hVpHqEzALJ4axl6cy3k73fOZFdRIRgw+OCHHPlj
0hLihQSHIPxl+U1fsgJ03y2tryF6Bg/yiPZuAlSpmChAP6mgJHiQBspp0SvjcYxC
1RLPK+j6XWntyTHi2C3urycELy2Q9kq1XneNuSz14gnn1vmZq9ELWEbCud4165TG
mY6I6V9O9hBar1jdvGx4R5PPG0qpax8Pp4qjedIsMWt+IjHsrr1tq1rurYtVOxW2
gpt3tqI2TgdkSGhDMBYQETfPz8YGZvaR1YomAh57gCllZO0czRLeuDZmI5k3dVKG
qM6U11UrEwZDOxtcr1Myi+KSTGXmtOKloKSXz8IF6WB1lcafbf3EHRY0JUfhH5Mu
zpDdv+vL133M+xg5FivwisFoGFUIs6sXThIQ95N91LO44Kk0ryaim3aOw+dhQ3Lv
6yw3Um749qBlvdfZ1LuA9Ifq6EK+8dayEXJStL8DMJ51QlNQmPHvhAC7alErQAwc
2PB0GR3+dujOnl4avFx0E0Dpd+YsvTguLBwRcMWND+pMJ7BrHsxitZcHCuncirDR
n52UJCOSg9//3o/mi9pPo53DIhNYP6qp7S1ijtP7o+Haml+N54THNad+cfjsjXGp
tVljuub4ghAwfMqTq8LA1PxLzL6FUGGDNAEaZi/2mWWLOKrdMTtC5JPevAIXP2el
QnsGKo42p237NyN/ox4EdNqqlbgjXDIOKOZQhHTWGrCnpHWLhw1c0AFCaIS9hpg+
38kxF86MLVF8B/w86xzVQbmN48IDmY59sVHG0SOPoeu1vi66aTni0TCvZP0nESL5
h/C7aRZ+3mPb/ST8Ff+yAPQKvWBX4a39RvmG/Pkt4RN27EH3VPy4tS4XUlcbldic
i4oCYJvrHWG1NXpapiTWw3UM3P13i1QdRKhfKGx9JheyrSRYtyd47Qpy9dFJQojH
Av4lFXC9KG4zj+Zyd+cUKga3H5ZAEaBdTZgNqic2mgmpFRCLKUB6E06W/fHDSgfp
zjAMemCEncjjAZbjWgCdLZPmGk4uk9pFnTlR9OfYOSrXQViz3YYwJtvsE1QSzlG/
aMUX3mQl5pSy1+XoHD4XZBablp8mT11BdiKgiRh21TV8JGOLQVnwTUGnJXFGNqoS
auQOWf9GWWXYkjW8oT7ZGLdFm+qQjmXRK2Gj/wSlBRrUpYo3TlIuZmXT2O6Uq5sH
Cb4DtvxIm7czZu2VQuj29H2DnVGazrOH7s2QGIIqzsdWDWPQUATQnYvt6wP1HhWi
aQKNUGNiSZUg7spR2z9A+RbkMPd1th41H6DyqE5YhXFCW8etVwiRA6P0Gj12chp+
OohhtCcnU977dpCAieZL7nPVIcKbaRlrsr68JT37PI8h+tVo1gzNPOXg1AiPXfxX
MrTFGO0Gvewfe2aOfPbFePacdFqWdE6A3IECYLeg/Dgw7E02s5No+w4OhkSf0vXA
t5N/kM2EeH45b9BC/BlxUK+yVrzocP2Ocr7/Ko8UTtzDxt40f+inzVzI+jx1+In/
W6moyy0UrUC6RpVFHmO33o37qZrgb5yLd09777swjm68BygNu3ekreioCZXids0M
7RSJzKzW6tdNCC+ZL1dlTPR/ZnHAxBBCP7A72qVZAeyYCxpId0rCiD0eNc59jfg6
2BFL82cP7WEzZR6tpZkI7CoJfjwD3IC9Z8UC6m+eE543tcTVC9umQVWYViz5D9g1
MoNT585eHbvcixJMHvz0HG5LcjuZ3Q8Dv2y7iT/Tf9PakFvrxW1v+G6BID6gWACe
Ziv6B2BSaL4jwo7183s+msZnZfD5Q2ouXrNUV+vUwE3a/dqXcHbmZZ8ql6gErwzz
1s0rcgcO3MQGzdApkghj4/0q1S1bR6Ui66qi4IYz6h7140sISx1K+7otNYtIWLNi
sPjvke8O2Nqlu4PTdcUlOHIKAJ/3oNLmCvXTFE+N6SQf/vbIHwxugx8hEMtsISn6
qkZXqOYqt5lRjUo/qFwP4M6CLvc/31dlre0q3cSTzgo5oudqkYhyKHCz4FstvpLh
g92E6QIcQV2aK2TsC99ZwFcVearSVEb9V8sBx6Ew4ihQqsu7IoUKOjNDEl9Ic3Pd
NvD26z88AGk0B/Ii5l7AuQu6YzR43Ot4GX42LkwBDmPpJdDF+H2ouqlQliwaimnk
YTrs5EpE//+iVZkRcniMwxV91BMULz4NxedKQfFo1JG6FipmU8NlPq3moTW9hzWG
V9V5sDq//DUABoGUEZFGY3B2OQC4A9jPLEnpOmOMdujXDh6uGjaR/gaPhdCI/zZN
zdzrRGxyoe9KP8Hy/LphxYtB9bD/bsdWXOfMxIRURH/mYVxYC/IZ//W0N/IkBVSd
0qNP2eWk8VlvS605Ny2NX5UdamedhSIu4I+ByVlA7/PWEMXrGeFU2ZwEYAWpykWM
aTki7hvQTqKMmyf227QzOpRiDBKasST00OaxpgQGb9yz2vp6T+iGDDXVZ50pXoUN
6BEk58bMo+gMzjou7vfHeFLKsdgHf9G58A6uPphBmdZ+qSigtkej3BHQtAehXe0c
CSCsqQaVpNmwAGA+Nz6OOvQ8nvSu9IYoYB7Z8oBDnW821lZnMyM7j2Wx4jvChKlp
qptzDV8BjofuUHOoLeGGtDRAPu5JURhPXpfMeR6NTG0V9xEZB2i7VHZg5Dds5LK0
rLvzkZrRZtwKcROOtAbjzSvKv+KzTaIv1Fizl3/tcxIMBYLn0YOy5wv5KzVQNWEa
4lRyyth1pWfHMCBvKo8NkKjW7/ArxiJ5cOE8hcD75/2RviAqftTBoOt9YvAKBb7B
l/v/DlTbUfhQWL73eUooHfDsvbvMz1uVzWFY89WKoEHKfevAAdzJdsjH7owaE/1B
fbB/lMqygN/KKO4u7J5F94aYovObJJ8l3gybWe00TpAoi5C9dXXrvJIKL6OC5bOt
uHCYC07QTmCy7BhvcdWj+jsztYKiFK7zHb9z65otqvx6hHyj3Zh8G9YgPw6g+vq9
tTnFkomza0A+n9Z/NV6uOFkzBIbpeQHkDvH+//1048PST2oGa047Pz/WHhDf45NB
RdlxsuFCcBHMlZp0uFFnczISdBgRgJbQDe/5JASEUV8e8FDRE2uhmpAF+SeaR5et
GjTbSUfex4N/3azjuZsJ9uOjQowZGNK4IwccDUdixbbYxk/U8judbC4h64F4cI2I
Y4TDljR31ZG2XxWEnVHiwI4Yis740nQ0FEIItrLBZ6/x9EFPOTVBVk0zSYRvgOAw
m259NVfclVnHs14+02nWciGHVsT1Jmwa4dJqw6mr2qk+ntYCNQ3TRgYDDo0ifv9Q
GW76qw4Ar9cbKF7L0+zxgi9Fme4HRs70tZ0jR8SkDXoCw+UZ8bJ5Mgfgn7nj41hc
56BKaQjj4OCM4GCfB1sLGviUCsRvUsSoB0UvyEmMcWD1VaerO+BWT0QxS0qy+lSF
L7ZhxSiLEhF2zpfWCaKbJecLmxSMhUEWpiDdZegVBBCbICgkptZkFAYqF9oE+w9O
i0hBGvsNsg4qHJh1vPTbH9RagGelojEbBzHrxSyHdyYB5Qs1qd5pi0n755InBQ4f
jLoO7c9EAHNi7qzTKCe7C+pprf9efpiVGKhUuN4oy4Lk1aRzGQhIVLA7p1+F1CGK
JM4qdL8gwhY7ycSaaViAeyyYdfzgctr3ZfdDA1o8e/SXMjAg8XxJZsYLyfvBfhWY
prahKZjtGxXkrzQjrTcF5ocySmHrWSfRxz1YfROmF5lcK7R427ZTAD6nIoeX+fUZ
hAbi0sxkD/LJFZlvCtj8ghU+UfV5VDh0ljqyd0HkzzEeX9C96epVW7BFwUoE3axj
K8iElwSryTg5982FIVg3VK8Bq3CJ1f11/hIoLohmH5kOSVm0940l90MiLZbGkTmb
wAPM1auhusG/VNdIZkT4CRz7wVv1kli/nlTJrR7GYKu2ojHx70DZc29/3KR24RZN
k25EnU+cfXIXZpMoLewf8IWwyWz6O9OaOWOQEUiq4+IieNwJNfqiL38UKGuW0NOt
4SR4eqCrAp1feANnpGCCHYwED0BolQ7EgJkYjjn6AQdJwbjY25IMfKI7NIYLE8Ok
6c8Gh7htaAsyNNx9qoUK5PHujX95SjCDk+mYcSa7N+XEeQ7hrhDu4usEWec4da4T
Vk/fF3LAvqynIvtAWdmREhr8Udcuv7N7tKPnyrrgV5tibmafQrn80+P5R5z/tsZ8
TFeLk6DtP5iOJKE+q8HBXRMBrZqLnp+HJzHlICuFQlT80/naw1GO+D+jD/7oi3uY
Z9y8up1tcpYCjQm8kJmnQqud2ySbV1AOkbfFrOSHnz+EhuXXbdQITora2OqAEZ2s
pEaA9s0Uxe6zItNbkJblkh/GAT48eowS9CXOvv4PK9uxCz70l4Nw2lv/2z63wGxz
hWTpHtId5E+PY+EBzTZQxTQUpEIaH0sxGEPx2Eo+WbRgfsdmrdET/EHkyBs1QD6e
3KZ3a/QzNVPOVfhXyj2yiBOEj9Mu2b3uACwyz4DNO399eBKIXFxG3Mz5o+wX3PsZ
+CueR3TZfzosvt96Mhi+peXkEYMkEND4TtgwP9jlpHQ4s0AgxZAlZQpAmeMyTTAI
oXWXapm3xX/KYy7ND1tgmXDAFZMkemppbDEgJuSrvpDaZmyTCNB9SoqeVynlLEmh
BsDWGUrz38vuDK/zQiY6rhYsIR/DGLU8CR1t4UO9NrkmlMlrXuxzVTiv4YNegF0j
5ESEZTejwD7wax6SW4lA2wuJfUgZHI88tFMUG0Muko2EM080+5PHI7mbfuVQa/D5
GIxThfVIhpjA42VdAXNLByKzGp9SjjIsPmYWxB/gwgvPfDZXo0ekbH+4zRbfr6iN
WNnZ1kHvFXFaFr4yyeqrOkJJqo2byNAnEs5IW7pWXuAVxOBu2znQQIQ+lkKibE+e
g188m1zEcJmCwAlXsFDPwtenAGP5cog2xhwAEpjGAkCOvD2k8EIXvvMxhbG3P1Rx
SCjA21GvrcXlkxgFTu3IivwJnr/vjtGs1bCq6AYPyZlfvRJUCeZaBoMrUiHujdzt
sBBPoGutzbsLnKUVEbDToUQSPppvzy2+mKG/D5tknykAbrDBQMMurvWnS5BV/GTN
UMb5cD+ltCZ4lmvXYGu6DRHtWr4bfoxNONm4/mpMnHOhZ/zA8DQlW4MwuFNiiFB9
IojSjlEFn0DEuRlDoQ+rhdBu+uE7tIzw4DknVli/oYg1NT5nMI1Mz2Vl08n09C+f
9e38xng/Diee8CQ3m7Ht3v/M9Pc2qW4VvwTyJwF8RUD3aQon+SSPOjTcT+zW+DDh
0XbICXjevqssXaI09x3t/NL0dxGjaULxOUi+xH/IYAhrrrmUHGY0axbXYndF9nqO
nZOMBOcTMiCmiZXDfDScDSFX+k7YvqfBiAVf3vwC8rfiDIiVP9sHD3oKPsBBGSqR
kGBmcDGTeKbn1grSru50nUjbSMP2FU167qZEmJTk7GbcXlCifvBUf62o3Z6fwtmK
QyVOY1CuamMqDjl2jDakOwazaFHj7x9t+zsaXwff3Rv/zPQp0bXcSa9ta2bqj0Xj
NHMz48+octu6KINdo0c00mBCU//2BKN4tYVQ4T7vWkKb6hiv4Z/1vUqTmwHOTopi
dxNwUnm5D+sfhWRtIywiQAyt9Ksvh95xbVC3d1TppdGm3m7uQBbSgfNLSJkIaqPe
hx3H2rkDuDOuvf95HmC5WPwtLkR/cuROb3Q2I/9f2OHt7sjdcU+XsLPGqsE4uNai
qQ6/advijRtdwdJWqQGpwuXCNzdAXhMxOCFS31oGdE+VNt8136VnhqbQiE0tLgBA
Vm75XI4M7JgvIhmzW3mxyDROUdQFLo64YMkS0aziypK30T0maeh+mk5vVQgja9l1
DqE9HU5Wox8LgjzjqcAO96Lo4ifnBEh5Ot0a1lVOZRja2/XA8qfO9HwumXdmYCjx
AYHkzwG77kStKprLOb0jOQFoiuc8S5knMiQSRFRJdCdAVmAWNXNlsEKCgJzcfUo2
2ZAtYiFIAk9M5uSltsJWSLFvQg+/hupPr9kfSGqBj1zfwNBZBu8erpUK0mzfZcQ8
rc90gaXDXY2NeFHU4heCMGtlNSRskNIkQMkDykDkrrz7lY8J39k/3OKjgTR81j1q
xr28wnRGfZ79MfCkKgC9WVlGBS+Huw6O13KWsTc0XcYr8jiyjOoznPAKvYanMKK7
cb0CiFLf2xH9pR28ihk+2PEXDbyLdoFHwark7MdCfuvat/xDqx01BWQSx7q05yS4
MG8p2qJqB3Wv/7IkDsKA7bfSixV2Rte+qjonIemKxaZbgUzwGgDB5LLpHvWm8JkG
9UIBul/UpmLtvA85BGnFyYPCqxFcenI5r+z0kX7C6QdeASItZTvZKI+KAAQX923Y
vs2TRB4y9wrIq4vRTeE2UCGw7UUTKGNIHxt7mSNXlBqeZnC7/h7nkZEDdvc07mZs
g8bFR9RyOIaplqrvEXtooM+HtItakwSSTc79d4WG6wcHY54XcZysujdX7ItP8Ewd
AV25put1U2F+Otq5LDWm82NHeWP9MCoJx6WraJFxHzw8TdtlO0mgy8nct2Q9Sbo1
kvMRDYzlYyYBG3YNu4YzdPHByLnOATmOgCMGacL1RowyBxKBkcoXj5+DzzMJMGSH
5mqDEDEW4Afb/hUO/EQOMPvv2tcAqBHLbZzUB5HS3cKm+8bKwFN5iyPtci3Jk0f3
PxvQnt5Uxf9DC30pWjBxfAY4rsadZ7nv2MUYhaSQYvd3ccHXzivveWB/Qu9RBt4Y
/aVXbCedo/kY21ooyP8VPNrdsBXvm9hjWNSY6e7y1y3IqGL7u/DgcA5tV/Dg1cDu
t6yANTb6nIbVTFMTBfQj+cBtEx3CACn4U1MM6LNo7uOrGrF8IeSj3U1lfMZhMHtI
8NnX3w4wZux0Ww8S1bC38bTJMCsCn4bfUA/yCMbkp0+D9Vo0e5xdLEcScQK2+Qoy
ob48IAin2z/8VYH1dfyUkA2E6N/wfM1n8GzWSYatGVxCzHNHg6b+1tdlrRM3Nadf
1WE0fktdCRoRcbRHJ1xO8wo7ictsMfBPXZG9eGbgKPSTJV7wc6kT6IX3opO6/TZM
rDi4a+7kHynUPr5tqP0BM+tJutggvfYHwFeCahrX1ZKs/oYEd6JcxpKy6hT6ER+y
jaB1mS79uISuVDVFnWoy04DH8u1J2sPtXGVTWA924W+BAGXO14/d1nEjikPCPyJO
VoItRgN92eXE5EDBEuJEaZr3gVPO9ulitefkxRTirA4PMQ2BH6Ld9Adxk2z9KFyb
1KD5TH++0axRtQE8+pxikmIzVUperY+gGAYFj1IFqkBPJK4ILRqOH4uWvPykstHy
Q9tno1+6dvkhGbKTqTD8XOAcZ861k7BXN/imSsO/i8vk/HhvKvDhB/iNMDL9cJKW
AYl7bZ69/OhljW6y1JExWPOhED0OeduH4NUAX+xAKEwQbi5qJ5fWesofEC+MQj8X
A05OgulXAlKqryosXdlC/fvotZJAvCjLuCPQTVTymofxsn+8MbWSxht1ufLmIDj3
xpCgp9TvxM0eXiaWPvNl14LrBSUlu3UhJr+KoY+w/8pOVtV13+Gx8LaBRqtSxUbT
R5veonoiQLJrzAF4ny8C4n1owncxUmhzyIZsGpJxvm2Yqi7w4Kla/U1YAZMR6dJr
i0fdDWz3D2k9sFqFo77QIh4AgeQlAyT8wgABe1hVF327m5IFjA96WSi1V5P1V0zP
fUWgf1RNLO4c6MUc0NNkX1kuInWCmkVvvCGvx32lM4GmF0g/paZgHMqPFCKOEj0p
/v11wZt6tEMo79/l3UOOnpTLrBfCDn9IWM4za9Wx9Heb16U0zvuCVBcmA3WHYmRy
b8M4cN7dNnLCXgtfj5sW0CRj5cdV5tDTLbhqCMFYiJA7cJT50g05uSFBrOq5rVwL
NptptrThpONdLVWZ2Pa1i7Glc0Jq248omI4uB5YtIZIRc/qHTe/2BZKdNT/Z6sAb
0G9bnbXcYDPvJ9Ty7Ew6XwSj92dLKXB20vZD+bta/DEv2N/NSjdZ5UcSlnqnHx3z
7bxPcMUSP2idtAHcLMRZ/Lz47Rm7QdVhbDGBHAuev/+E+z5aQobL11SjBW+K3j4k
j0Ok2s/nFRUIKqUCxFmZYPOE7GwC6+Z4OxLy1Ep9R4ZGDAzerC51Ky1qWrsxDzTc
8wNRAMwfYcxDV1i+/GrxdmMEQtxfIyUxdQWsOEel8ZQL9W5m9WMWIKG87WY3Lzb0
YVYTUs4TDCRZN2mucm5B+eXFPqxnllbp40l61uabLbDqMUYEyicnhtMSnSiw0J0S
D9hydTvN7vM4xLnBGdD5q0Cn/WXan8TahubM7EpKAqYkRcZZc40u2f7Ud8Rk8ydX
Uca6jBmy6IKV459biujv2dHgP/bbdxzGzofz+g2zr4UU/F5+YdcGqxu8J45eIlHo
MWYRdPb3+tHKvDoqqzSPDCgNnwqH9gu1yj2xKOimskBUdgpV2lh0nAtIIMOlGwol
3sZ28P6tE4eNc48Ysl1ftxBGGMb6ZZgrGR7pVgVGlkqP9IpNCD7DB/6cNmd7ep8f
Rq5Mso+rTszRroq2f+MEpVdt7vQNmqtX1bi6rPoNFO43c8x69o9i0RkWEACEnB0t
CEZyEUIPjy2b0ALL2Ne761aWCBt0kzBYUuwReb1xcpAux4WvzrxuYFYksv7egBmQ
oqhTLk7+2/i5rjx94kS1O5MNI0ZAHRhBCCK2tYseIL9BZL/v5YHVv+xD1T66V1j4
dDkZs5WsJrApAeN8gFECY9hvYLLihHSQMOg5hjpt34NEqDt3y7IYnfUP8Vt3InSp
yF7VXCcHaVKoH20vH2cW6FJNfMuGYYByg4PfEHMGJo30vh/n+Dmvu14YQaixWedj
x2ennj682uVoaK0rtD497/RZqJKrBzUOUexgaY475qPyNTlEnPKSoAiF8cPybyo2
aP5LMVRgI9vyDIKek7IR9U8CZLHrgJ4I5It+8LzgvwKbT0pkVDnrBhbjBI9s3OG/
VsC+TSthPM1Bp9SOxB720zEoefEF9GUfznorCCANGNI8/UvMy9vNTsShMk8Ruqql
oLn6z++q9a+J3FLkXQEi6n8kCTy6I516MrbOTVJzzKQQqN57bmbT+qurR37SkOdd
lCeGm3USFkhON3SIryD7spvN7YG0aXstjVnFdTRQoUq7gV+DSJC4QahP1h3sr1mF
/0elTBo9fUqXSUZNnstEsheKz9kXvq7/Up+rGdlYfwaWPznJJ57pf45U6GpI6zfr
QAlELfJsK709BneCl/VNjKQzPmQ977c/XB55JPgCC78S9DDtiS0lXxzDa1aX5GMG
vdZXDSWkrxKM88LHDevzHghoW1xoChvfPWPpN3QGONJ0YQMZ6IMCe27I6yyo0jOT
O3dnHCxnQZEeB71Q4fE+gDU7ncX53fpwICBJtBIFy0KZa8jPme7Q9ZXF2Jer/mnn
By+tH8OLJVHMpoKJvxUl/IZ9cp2R4Rj0MSmHeLwTq7riVBjUMDYeiLqqa6QNeXwj
lkhXyaHyApM6ReREOU8XgsNrf5/SY6N8ZiGHuGiCIECOKsmIP5YwHa0h2JM6lahk
VHcKmjpC4VtzZd8yWSk+bFIzuFimmM6N1TUpmv+dQ67gCSqnw0YmfBvEQf64t2o3
XEM8UTaLUUll3959DSqBWT6ki7tu5/0M+u0WdHvhjEw/5ZEP35b1D1QTrxi/X1JP
a+YIbMy5wk1fAefsjwpV5edu9ikczMPv8+k0pchrEtijIzdQnhd/QVBBs2ZcZsDZ
RpXo3v82Je3kDbLRjmPjmoT316XLXly9XZyh3HsGiShcPRj6l70X5n4SWOEjwh4N
p9jGHZIiaiHxc0ST2rWgCzr3ZwkGFJsMNRa5/IecYUhQWY50q0MVPnVUQQUO9vaY
4qXy4xiRLZkMQe6BJ4dCwibfj2nS+u27W+njjLsufkTrTj7XGPRAVFShd4fzxQfs
ovZCldv35h8nsGeaPaRyKBCcDNiQ16V3x0ywcwrQGlaDP2b71luQOVor71NgIzbK
eRasKaeTQzx3RtF1/im82kTstvBxnC7qS/pnuayzQ8+rpwleXH6zqiD25tNIHLHy
lhnPeBpDTWRv40yaDqF9+OPgXARByxQ+DEAsZkXiUEPqgQtNL8BOFhyungURKjZw
f1SWZbBuX3QTcyBKABDuBJuUjuMEhHKLBVs46oncHE+FNurp4su+1RXkEkEAJ//B
X6zooQiy0lK88zJ/o30eBW7dQp5QNmQ9ZPYgrdGXf+vkDHOP+H++zrfeTbCNFe+r
rmsekdGvKA33l3hXrghLJ4FA66zMIKMrMhoXMHcbxKw/6KghenEtrNeYkLtvjPOL
tNOYvvvGrHVTv7YljGmwvryr1YZ44UwrkG3FFrNDtKH+uBLgkDJPbHJw0GdHK1w5
EEa3h6Rc1TDThB0/r9+EVNEEFp8CNbQPg28bpp3+WYEZJNhSXdt3OOyAasWu/CvN
a5agSuvx1jyFIBYRNXDCGIFal0fAI/Fh1AwUniOUXDKeoFwxdKe7hEKTG/sHtSPM
VHvOmsY3lzwAqUMWigrujL3B5r6VwhqDS969flxmYoJ94RGxPnI9YI+F8cYirvi+
DhXyLb2KiQLOpOUHkBUgGCWBCpXDf7/3+hc3+VYJAhtmOz5CLOR80CLnfPAugFF6
g5FB9kzYwMIIRux+U42xM0sY1mtaAmiN4mInAaqIK+77J1rrRA2+slLSkcVEcFuX
LaDE3I5yPGbBoe/UnuhTLVhGBtPlcf0QIUpLFKOJ8hqtmtFLLcS3iqhZhysybuAJ
Px7mvRJtLxnhLF6XIjdPOcW/ksC1mNVa7pEFSmofGK4bOhkhhdMBYbEtHMzaDHGN
aneniGRcdu2wD6r45Q0h4Y1gUrO1mS0vbILDmzo3MxDbF0z5IH2VFRGjT8t4Kszf
wXOZaEqr6X6Uxi0W/Dz98EGKdTCU0sowmRRGtdARppJpvy1VhRXDssRWdYTuGwTl
gwYI3XF6m2Gkg+v8wP2zb2mUFWOLZzrk1i6ZtMAFc0zgYBlvBkUkAiYk6GuJK9Hj
SWYDKnny9ycxX+9vkvipuk7KXw/QOQzJVnEVYYx9eJNAUEUIkuSrZycqmFxCyVqD
+RcHteBIVEN6ZJbaFew06K4ZxkwfSBPjVYsjYJ2fbGXWHrMy0Tmm+NEYNB//uA1L
qeup9shqEGNX/SxvrhfM/UueBlcgVJ4pOIvWL8GfI3ABeETJ3uSmk8pm4R/x7m8v
uPWRYiLS8kQ2SePg93PdkDUpJN2sX0Jy1dFD1wNV+nCsroWjq+m8XKwT8rhXF2nJ
LxjnGnrB6V/GblPtlWKUwdrtljoQrNYMqcwI6yoRrP2h0urm5xJq55cqJAgP9efq
o6MqiyfcRXHzs+nTEdRqDM6FFWCiZ3sGjYJLIuL9AMMpQ8MLkGfFWNpsEH28IuZn
OqbNljTND8cxuBsrKgiK3ROCCmkRkG1W8ppPGf2cplTnp62de9nkW9ZnjVYJ0E+K
86yUWL698AaQIu0Xz/Sy562Kztbfdw4lXwf4WlzUbugWjbVwKFHYjAbeCxoESZME
5MrT1nfPa/FpkART0mV55Los9QsRopilwh3fr3B9gpazRQzRGSfMbGaALgcrK39e
uo3OOUTOY3oVMf+ypj+y8JP3zHthAiCemQ240OQjtbuCflipD38sTPT0/FXOxD0Z
dhdkvZh5uY/hCHpwJTj6r2ehMskocn6yRpTu67Zb7Sq+zi8gf2qne2iLgX6OQj/G
9CN0b3Cj9KHuFyAg1I9eIvbHXIXxD+vCMMipVmdyGVhf5F5qep6XJ99OjIMw2SPr
FTVlqdo1B2krcApznwyunqkpK6kHOq3mzPJbplYF1gpeTfmAvC/D4Ds86PUP8+NW
P+8n0USBU+fZGGj57rPX/2qeM5u/pyF1hXo2T/XuynNm5wL8SITsezyMpoUjFmNN
FRCrxG8r5EHXEgN726fLQlhpnfllfs0NDDyAyPjHyAsZ/oaOBYYdmVb2P543CYKJ
Ar2PiMUppX/UBT6L2dUsl9pcHxlHbenLjswGk1MkShFbsce7EjuJgTjG1t/ThsRb
Hk8nglXel6T4uGmNdpRvWfcfPJxCb/RnFEau9vR8owwdCL/62Bn0b7CikOfE83k2
ZuBAyPfzpP6B3E85pl1qDq3KM+SIigK8Lt0SxvR5mWiSXpsMhawNk5D9FbaWZZQV
UMmG68qELfXTxGcIJcqrKYR0JHRo+p4u7mrLy21rGdp3cRNQHco30KRtDZSYuAqw
9B1muuM13yKkql31DrWebaY10hR1exOcFxi8JCkrRUUEn/5aiD6ULpzgszKSPNBI
niCeAV2rZCdxrdBkfWcxJXg43E305F04Noi9n6APL1ikXqMOmMfc41fqf0joVNdf
ZKbL3CPDrT6TbSfxD++DAUqCELt25rpueWgzxGqWKuAtphKJTpy19i0GtBlc4RrU
EN5JfhGCqzEG/Eju/h+SYCH3a6+TEbsqqUbzsX1DQKiZUFAZL7jrI3lqlmEcZOMc
1ZS/N31U9VAHF5ckGk0mP3bmDNAqiZgRqOKttGuXzuZAYGwHyBFQCMvQ0vXQhqpA
1nwGt8wUf6Ma5lhHUASv341KDiVpJltR/hP6mPjv06vSF4WpnCgtCjLd4cxBLoRT
AC78SqNT8MDos4mR+rBgHkASkEjzYszIXbzCNvURsRgCXjm6Vmx6tW9BHTB7qqjl
d+lB27pmYbcvS7GrsFGts8KR6YS3927ssppixGbYeLfQ33awonWEv5aMiyYCeuAD
tF+qEHz9mv87laWlrJQsBVynor7HKokCYpuF/9ncVJunvr16INAzI+ZlaD1qX5/V
M8ZokYTLocBezDXlMYgMoK/GP68uv5oxOm06QxR+Y34rrovnr7mluccwhB0Y6kib
Tmw28NhXQNzx+9eBhaeeJ4hARTnmx7/OVqNsNhGqUjHgt2vbpOWilgQjBzj1wsT6
cPhywAZgRk1eD/Y2dKKTDDHpcCXNbmw4zeW/WfqoaU0KmPjuSXig7a4NMBrkH3cK
jqe6paJRH+wgPIwx0aKJMfnUc0IqNQKOVYcqJ647y16F7iGqwvukD1DSpeHL2n+c
p7pK2xvpPUgbHKkv7m2P9u5FB8FBQ5gB5aj2rFjTIrtOT7LHeZGunkgjEOE5crt/
X6zho/dmN3Z+SJc92sUr8+kadoqYsJY8tenWgpFiO8JA+V4NvDkmBbtZg+TrHXFU
T90slCutg5FNiwLX8ESIa6XjYsR7mU8bzPQzMHJjNc5dr4NzG6A5wadD7IE8xZOl
9/EhPgusCkdjCK+Rh16bgl+JGEqtMs0Mx4X1Kp1ITgDcd4pdjNvTxQ5RTzddX1u1
Z2QHiwMTJu9bmRXnFSM/HoEMsAKgIiNI0k51FxGaRHSFh09oa+VL9AAPPDzn/Cdt
OLtjZdajSDJuYxAlfHcyhLNXJIl+iTlf3Cv53/t5WABzTig78T4XM1MHb+e8sJs2
NSdYpB+Vt18yJ6GmpV8k48ZXAAhDOiCAq3tf+2BcdZODOD208oW3g15KHtLefMJb
AIjjzSq3XeHsS125fd6mf7f24VHA8TFYaXU95m1JtSuwERLqAxY1mXdPFw/2OFXb
jXE15lxDRd2iR5O20dPYi9zJuGipbrUc5GAIC5I1XnuxVOkHcMWrb8CW68ulE1T1
0LNBEm9zJ8ZcGQLvnMdQ/0edZpTxhNc6SPvtz/3Tsi+TQI5hnV9JeexV44ZDaIub
vNTrzb7BNDKWXhsjrjwtXxSBi7PUsyEviHfql+ngZ4fVpg7yYwdYQojGRJndBYZF
ZolefewW5/OxwSsZyrxFvBqYhHYXqHvqkWVFGHw3aSUXO7/y3pc4UtQj+e6gENk0
F+ix5sTKh+sWFMOJ6FPt9JnuTUGvcMJ7GCxzdzFVrR2+mnFs8tpDBJggU469ZTBc
NaaZv4epG0oONfrk3Xl6WE+gZNztrUe2rFOowKOP7iWjdBwkbEgseCPp+FbVPJiT
ib8bZ+3z1c9du8LKt4KfkHY+MfhTftvXl0nJZ3/RcBeyXFJK22REGKsir5E9Z8GV
o5HmFJ/kBaVIn2lPGvk2p//G0Kh4SDkc86PzWfrnbfmOO+q3ONZyzvKURpHNC91O
sG4qe2Fyiz3O2LNTZ4KWUVZAwZIPAuI6yF48GoRwA1mMKrtejOQfxo8zLY1xOAAg
fzP2w0jJMtkVJajhzUuzB3Z+VEBAc+7BJlGDrvYSQP/z6TshpVDmA5YcIdHuUnHg
rf2sDpQQUQgoEAe4qAQAx1+JK/ubOLjCinQPaLyiqKz+J5HIEpr6SILqmX5Grcws
cpep730Y7gCt4PDUSLhkVxYjQ0BPIY6QApKhELn4xoAXapQxMrbB+qYN9+XyIU42
jRMma4nQIfDvIrMHLMPWLn9KriO2+iqb1FyfAnqvVBJTtElgp1Uozdqhql3g3hLP
2R00QJP04KWQ2a9gQLooES+seTbOJAnwUlT1EPZAG1oK60RUYgOluMRU6Ev79qps
zFmuCjlZFkrrRf5ajNM3HX6TeMEWsBGwE1bEmeqTEb6Ftzi+JdyBGXcUwL3Z7+7f
qK6oaMmOmtP+EwXg2/yiAM3Egz1xrFNr5phe93LKhHVcXbLlwdlVryiMGpD/97OY
fbqSyl78vrGODmoOSJ8pJEN4bfLFZvdlYE/D9UI4TMiRlxhMaGspkFaJbBnqE5Yc
83BwaFbokvS203EXNczL6gL4cA9d3vnZkNHmi68owMODHoaTeWoALZ+1r2o5j4ga
34IZyRC+K+4mE6sB+f+qSXOPaX4ywlBbFY5rn3vnoKXpz2/3TljMfGOJkC5/R8o7
WVWztviOTg6Kt8V3FbKnIo5yE3YmuwlAL5hpiG5hlc725Qnrr0Z/zhpCXm44/5wb
6sO1z4HfDcu2gh/udjvUDN2NENk5y9ny8mjz1qXWWaYxJNJwOfl7w1Sta2Pidx4g
WAxJbKu+Qs+yxoz604r8dIb/P1ggcGuuYqQ8rofB7iDj1BW/0URF/IJbJck7oueZ
T0KP6mCkt9Z9dffFj3zXCFl7G+QZUCAxjdrboV3ph6jfbJimQYvT+IUdY3yHflm4
FltAA9XMR/+d/x1DXiwRcCQ2zl+6WkkrYfHWOcGzH+45N/KazJP56y3KaxJruTzt
3GPIhGtVEUN11iXsRXaOEexz8lHGQc3CO+miqKbonkUE9VNUaD3P3Kjxk5q3CS3l
IF1ZaRcPUxvfcByrV38NAcRRyIurpqT07BFMz+jjRZNPVdaXCgdRA8ff/ovLi8jS
PRUkvMhQiCOk1vKLjnKdTsiZM8VXJd3dIVfjgjnomtrOn5poPAeaE24coGNEPWMz
lTXLpUPztE34eiMaf6c/Z0n3ijlGfEpasGnN/8/k8QULcXriKCmBT3ZpGPKeOmh1
4xHXZMDPq9eGvFrWaSB0UasDyMW0wv8+1tyElVTt4FTaWh+L/CGpVwfMwLhyFqXQ
PFlga6lD9rOOc/ukXi7dA4MQGeri1/Sm1rneBPRiee2EgjNr7G3XwTUwmGz5WPW0
rGd3CDWg8+ntyjLyoU+pjgO+ysA4HBpL5P/sj7ICaqZe7QFiSRkbJiRyS8bzxevt
Mk9b1AJLetW6gQAS29cOlUlHFmSlOt2cWL1+tGo69CeG/8slUVjAUUwIq78OpCwL
fSH9lkuudEIWhTM6RlNT5W9jKSC6ywgoKBFB0ZJVWJP3DNLJHNdfGULtjt/YtMWA
SwCqJ0hxQXE/jg3LkF6T2JZ2RzrqT/aLbvUwvrNRo0mbdxF5VbAZUxVaYky2sp2s
TePhOGvsAf/RQ7dVrzR+a2HozilCXF1yoHb+hCA1J4FZC8FJSeqIEb0bC7CggC8b
wZlpYARpmdQIAhQ8ss5jnvVkESZdMDB6C1PgaUbhGHLAlxlsZiPZg6cMezV8MAMC
swYCAXyGzG9tuN7tCDBI0BrwGiKeCE1tBCnVcroW7oQyGQRJhBBdIMkVHJ29cYeH
D6wsV+Utcd2Wszl/1jZjH/PYNhbGotJG1G0lxoqaJPIeqqSs43OtC3Ag4JOlszA2
kU6eVsl2TSaZA2J7QE6AerHpQWY8Gn2/OjKy/0hY/Eh/k8xO5yuUtiG1/uGShFF6
yKY2DCaiH7M1OIdko40aNkBQlNhFpLswnxvY+nJNDT5x3WGTNHsRGWKdUO0hssuj
AnPEnY/qgeZHOiQ8VwCoA+EU0pN15qerixOThigUsAb6gVnw7liHlK6kbigYedpT
Ym2XH9bnVifCEMbsB9UsPK4ok3xwTbWWdiSHHwbVjoi8pmr4RQKkXm6orjjroq+3
SgvjL2//wsaftfrZ/nsq8py8M9r/iUgK7nPfy1HGcnLMcH1T7U8FUEyIVuM4cXUy
DSH9lxhYI3ZtBatyBMbc8Dtm2qEm+/g5CHjSLsbcfFCwmu9td2uAYzrhDPTJHCWX
3osdSF5RltukaYsR2J5vpoJilbXXGl2XVnvlyVM46ldNhIjMcJ5OlYt3fQu2G33R
fdV0nMBPATkmb+QNMCXZ+PXu244RoeXsL9q9FnZRvmy/H5N6LWnVsJIZqbKJlmaX
WzsifXC06JvDfTq5BIoXjPeTPFlnNLJLsCk4B20X+NtsMBN77jU+C/AElVAVF6+0
FUkoRHE/3aTJu7vl32xxxASQL83TG6El/MnUBq4cNpaO9DrNda5/V0o6EEjZsE/T
AsKcX7isonmqho9y+9RVGt6MgCNrGeQPzcd2EGaGRxQ78F+R1gAkZ/qZFWGFsNCX
zliVncO1qxegJmRXowlB1YiY/I1LkLbDFGH7v/DfvomBL9eHA0JoumEWqGTqDviZ
EYQ/RjVO5f/I1yy1QZFNInpPyC2XcjGWldayPmel9uCzS865bsEZ36J5OuUZRMps
ZArzWRkqBe7gUMs4nOoxoXSCQvKJmUu6CvQJfGXQwMLGRrLWONHKRZjpqKr8E3cw
/zyrrll7YKqL60oDkAZ2/IS3rgOmZJZKjqDl7ACY8Lm2MtAHjv8taospwl6CB/CV
9dd+cVF5sYaW/QcxMoUEyws0wXnptQCjuNz2X6Ys/77IeRpa+maDObpz9dNGPUIg
gajB7cWUcZKDZpJRIpI2duyfy+s3eT0Chcq3yRxVBncUWvsvt6Ee411y3DQJ2z8p
cnEoGBCJ8akMwwng7iHvxoWTO3qUg3MJwmqX4lhXt85tSq97yKAPz6dw2Y71ftfC
GjG55ubbL8x/Phvdc1q4UpIC0/DJb/Ut6M4TQaIododv2G++pLPunvQxLeUyc8j0
e944NmdKm/rjvkGf+SwlPWD5kQQXOMWPdMriK9niqPnaT/aRUtPZVlJQC1rRdrNC
fvpt3p86D/vzgCQY5147wlISzxIF+SCYPRq0bSWYUwxeEqJI00qC1npJZnXZiESR
XbnliWnDOOfXy4eLqZVzQtTJ7t+SLYi49gpFmS46VmwxV2QD4vaSCpmJWEZwkzVO
PTcFi+ZnWcpZs9ZkkS3rI2s+cJRAbsgHakaUUgBsLC15dicznZMnZGRZ6EALSEzy
06Sxzrmtfux3WHQD7uHFHrWQ0Y7fycBtOVeei7wIFrIQ05ggK625fG6T7/VLqePw
LffzztpExI1E3hf9bGCSdHIMq0RAYy42MAeggEJ+zWGc9bf+yiJRBb24V4y1lKIZ
UTw2aEnKfR+IgCf5KC5GgVlnRxbRbwHAZooHA1Wk4le0rMkoCmoTC+OirlacnB90
MxobchQ4ZbHIs7tflPNAIAUCHfpt/KO2UawuWOAcEu4xgpEXJESF64W6v/McRcxf
+SoFPkWSpbIJEVsqf6ZKftTLz40tIE7vkDTezH06q8Pn2xQVBFW8uWMfOiwey5z7
CfIAuLzFTL7ol9++soesUfS6wwVeLoDh4gjJXs6kxN17eVDbTBO6hL3KfXgYRmTX
qQuOhhhvAoZthMrYA87cx560Pju4H2Pj8TdM5I1C2cvsY2iMPrlg6kQyrEP5w/S6
tXdU3J8MaYrNLDPgvCJ0sB/BMJNqHlGL5Hh4ee/I5WW0DuIi1A/lbbuSqAg68F3N
wAB/e52cRd/7OI/IxWvk8HeKZ0tVldfTWw3QwT5+qSljt/5YorWzaBM5jq8K9SBR
92FBczUQ02LOXfBzpfOeMyQXUzWQGTxZpLZGAjPQjX/LJhOwq41fOOTsLJlW217V
+BWN0ocy9IJTfglUlEX/PrFMJ5FeYWUXlmOT53oMpHMEoLnBB0HoG7+mGXKl2xiB
aHOpE45xKhmnMa0uuFAZRxTtWZGqumcIfpdUIlEatvDzGLZjdV2tXQ1vj9FaJX2O
eGGSKccKRbDYNPHd7/duCeyXplgQpXMzCHuP0j6pBaewi5OYLxDya6foUxFJlRcA
uFQie4WKZL0CxNEPvpdHctaFkOxEAvfAH1F9ZJ4EnITJkgQ4lgXKMc5tl3HM8Wnb
T70SHDFAITXiXZibKQZX3iliENy5rDsyEkb+ApJAww1z6jq8oJpuN7+YqmweZCMJ
YJurLGey+NqirmwTkpmyDenIreZlj+kTEPFW2adfIbJlorgMURPQhqCUxtpF/OC/
gmlxtVAY2w7aVYjBbgG9FZQgAB+A80X6/oAnfVyNOgWCht/yNtTXiM/97+R+wrOe
pbzq+D6HK5e6MyfHXrIb58OFbSeRctWcg6Glck+KxbteGIqf6BQvHt9Pp2/kQ2pt
jZUHBGgB2BcmbWVhleTsYVOImlxENbe0fvqXO1L0Gfgz/IV2cryKePexy+nWSBDZ
OxV6wp8w/kmj3IijDChh62PwRTfPfFO3BoI46npmryugO0uG/Hvl+XZkUBo4gdhG
5WUH/ibdRIbRywoOkDAdVszsnjhBtwKmJsOtHRX6oXDKZAxQzv22cNapqrSj25JT
IhoO15TLVdGRxyc4m/s3Cc8lSbhEU18QJZrMd6nZVOg588A2UdoavCFTx7GdZXra
4MWVBC8No24EMgPnCBYW498z6sfHauS9NkJNwKNtWildmOYUIBnxlBoUUnLgwomu
6lE58TQI1AtbEmNvemQ1aW4NiT2mHjDa4shFQCA4DCk715KzNx2MnghD3+UGO5Hw
QABkj1gglGmEZF5NddfycJ+fU6Gwr33K2of5Fh/HidyfRhzjG4Sk3BN7203fG2/T
uCIqHiThmOg+S92xDzarfdiVzAVtuz4RViV6YAfYagHj4r3nbtLtesev/k4m5EdG
86kk04ShfofAXowLhOAbODuSCAkQC1z3ur+d8bQ8y08765EUrW7PyuGKqOqbnUmY
1RNvSBN4X8OAHPJvfxOvYwfL2FInBCWnvl5AfBDaRT80jkewx9NNir9Ec7E7KClP
b8acYp7YgY32BVM0Bgk0sMZzgu/nrexOalm5kSfpO4iy60Y52cxFkLP7nUs9gOP2
Dzm1xQUoLE7n3pcXHZbDx1irhJbNafQTuK8MQPw6jDI9IIMr0oOF57I1p7P6zRWe
AO0Ur6xzk3v1tCxdc62LeufK/DikNtMm5og19nCQJZFvVkY4wSZeDfcBBWvmmnM9
wNXGtwl/seacVF1N9CfLEicsAy3grixvcE2aYCVJi3SEpNR2IAPnJxOPow5nDbZk
TTpyTcNiVv+6HDm+IeMK1qPHBFkby3f9K27YEJ0cElGPJw4vgfOgApX2mEJfPNtN
uNTPMDsWEsXHG0s4yHZ7nbpJe4VYvHqlTpAeC7+BI6G2k5V3f+8VvhORCe8FsS1+
X7GPLdfm6vOk7K7GKU6QcHYzevpQhFCYwhwLrwa3G2GqQOSAL43GGSZLgMT0OFGn
qekGiMrLGygVWnnH/oEWbyNP/ATzZezo7tFcQ7XLC3BTV/00otjQXIMe+bqdBwbH
pF9j/2B7bnRxBVriaeg1D2VjEQfjQTb3/s5nk2OJ0o9XW90vvi9L9IQrUutdM8YP
jrqUIe4J9LTR7OMatbKy1jZA57+INfc6eyqlY2zm5xOMKmqv3tDz/EYZ+HXZzL2C
y8JLwtm2KKTuD9f1h4hawdsG5VS5a3wKE5cS5TV4cUz6V9VDLY8h5rEJo0qXh7U9
Ms2JhBue16K9BqrPU4JAQz88xprOgJnCmviyU2J56ebIQWYFDt5YUJQhfB5A01Da
8aev0ee+LdvJ+uzGZgz4K0YKHJzTw6nNYWOdrn7perIt6Ztg5sEp5qxa4qViVa2P
LLapAwPQ41QlfkQ5jy7aqdkxNGfZ5HJqr64MUIe24bXKD4R5Q4S/+35j7K1i7dis
+T1Kf2sd9OmsTKBV4VQKboli/EljBJyXckWrqZQYOOVOTd98CGoM+FC7eqbVIjUk
Y3OuZZuvoxPHz3ezKcH2+jHfmCDRMadUzpsZK7ohKTRJaQPwIKEAmkjsz+vFzoo+
herUdc3UbxNG4WWjWh6YZ5BotJiJ0tYZ++OdcIBPs5Awm8bjSBZVVaLd2CmPfeW5
5nCbTv0YgZktraOW9snVe9mFSWOlAXXK+c/hynCG2Kc7VMSZtvm6Q8qVfOuCbiOF
rIp36wV0HCzHkyZpBYOx41tWDeiPaQLOdfcnlfdUWrAnpI+o5ruiMN+vymgkb8fl
dy1qrn0tlg1rzo3f2DF1BbfWt1aq37PQcqKaznlXnhGZe39lFAK4FIlFkURLe/9U
o9VPYgL9CgGkxn1bt2DfvY4UC6szPMTmyR5dRcteet8Jro0kJxCMTwY82l0yjL6o
CViJ7BZR3toKnpIfP4KX3/0Ql/5et91stPse/1ewMxFB5mGyTCOzb/fSDfA9uh03
XEaoL9QlcVIqZ4aUhv0ulX11dDOok2M4WEKnRi/btcPoRo7hO+b+TcV+D9TvzXad
MSxGBwEifcy7TBXNY4w/DZoYv1SGY7h1TS3YXJqYxzvJaro3g8qkT6uY+nKyi6pR
kpfQ0ATiAEXnSDDgss692n5aDStyNfv8uR+8B/nrjrBAUYsIzKTvgmWXWRltACzL
VbuVx7mu31xQjVbFOWmh0g3T8+1ODWisbhe1GHznxjHcSjkg7dlHztyPvhApUCyF
wHus6FyJ/TR2nutOf3Pxw3WO3VrutakNkfyXX7Vyvcriuu2cz8jw1bi/rE+KjaSO
gz3FfhmI2eRUyqzuw4iwGrmPVtoMnd4/MrYtmo/NmII4cQzxtuSIfsU7GeguCfyN
MT8eu1llqXax6+dpY7UP2XEX8nBfApcRduas1MuEuFWJdNQVLXgKL/2qCdtq4ka0
ICO9hZIP04qSQIZCS8QDlx7kJ9iK9tlvk+BT1TzLPazWNk2h3ql7scYHbPCAMQYX
+RJlgbUPer5itBtIa/knis/UWaIz+uAmUBuzYjXiM37QtOENgTVjDdiqmMa97QoY
04NMSYPFpkIcvM08IR4HwFSMH8AnwUqMp/tu7jiwT5sm9nbLJN0rvvk+51QtdZF5
Fsf/0Cm3f4asCTz4W7XUQKbQmaSVunGFPQXvmvX4S/YEeLSpeTwdrExQEc7eh8tC
5C6OSQfBF6Oe+MsEIdf760i/9QAzUekGeTLYgJzgUfUsZJNhhO5GmarY3ivPIVX+
S36ElrLbipBZRqLqYucXKd2ujq9FBo1nvwYEo6bBWlG8P/DhDgOMcGNBBbTJKq7B
svKp9rmOCZwGXr6IuC3JcGZdj5mQ/mQLHWm3p1cePVBF6PFOMDL2Gbfg24jcyxCD
gwnQHoHD5KWjcnwAd5+5Y/eiLAg0VLZzyqNGWvncrz7/n7yAXyY4S6x3v5cr97Zc
/FYLRagm9+uODb0NNkHYYS8/XLtkN7joSnJNdFuf55l6XN02VyQQydI0FXNNAw9k
o7r63T/0jo3PIdSN0oTTfXPi5fhwCtpGwdlt8dqfHXwxYmrGQUqpgK4IJ0Zgfyws
+ze5U4c5xlLdY+8u1ZFachy/Ddw2qhO1Hd7hHdzlfML2ZADlPDJdrtUzLkYfH42A
AdrkebHewxN5iduJnU+Ae4P9PMmi13yCvcn7kA6CUkW69hqeopkIgvlx777xZS36
p3iyZ4L7OwlA7/qH+rZ2H4rcMqVSZ1l76WVxwvb2kxeEqfJHIl5Q9O0UqV026BPx
WJJ4omc2lBfFc829W5DILpFTbEpQU2XS1jhhaJsA3arboQIAePt2pGZh5SGvtdWt
b2dGv0QWZyz0XYGt7T6LDudDaby+e19PDKtNQSm5YPekEr5NIw6wwCPwLAGhkVoB
4UixE6SIZnR7XxnCTyhk2sN4WJKn2YAMUgHS4QIrf3zDjMhYdm68Vmm0TT79Aod+
ryHu+ySb+0UJhc04VVHdyBdXxIYkvabQCnXro7+1DuIlzLXrS8SsYsAry+cLTHi2
ZdJsQV8wDs0Fcm7iiKS7k2R1+xPxc+Q3nYb4+m0omBP3S9PQb2xY5RzErBGeryXX
EzOXyYCSrN5zOIkUt+fJ3NX6EQnQo2Hr/9GDVNt/pOew4ToF9q90JYQgjWFu/XNF
mrl7R0kEK7AMBDc02vKYisQfA1RTI17F5+aXR8v6WvxfYjd4a+OkVwBIRQnDPt4M
5Yj81fdYRTHhJz33wUMJlxsbuNOi6QvAjTvXC/Z0HUfhC+rRq2YoNpkm1q/vr6vq
FJKMLnx3bEJIncr1gclvHEozPZdoUeEujFNONniv/w2ztet0MD/4ziOx74po7Pjw
0XfW1HruD2ov4WF5CPa1m0S+0Q/Tylpx0W9OA1ULIdgPbmkhkWaqk5g4mpEYCcI7
w0aj8t5vWwomzPts16bRiOldGHdl0v6Q3SIic7rW6BqaYunYunQ+NwCQL1XGi2AY
8NuRAuMqURGTSUTfl4t+kscZs7AZPTkT790Dba2V435UknwTOnLTCdLO8psDAz22
7EET7CsYE8QNHAILEbtvIV59fCY9zCs2OLnIBWxc1FAX0h4OVzO54c0RDgXFswfN
zZkREYRIveMEHy69LiamnVOr34i5qeMZBiIcLiodPdB2BcK0c25WUqeBgeVbKaPo
YwXuR2SpU+Q8yTkQB23JvBpH2jw/s4ce4nM+GdPzC92AyrTv2tiajaYLnyPx3VcY
GtRG4B+XhkmM+ns1zOKikXncQOD4UVB1kZPJ3aArrjqJZLvFalbjQmCczDdObaGy
zjQdytbk2D/0Wtj9lG6FJWrs9noEvG4Bj0EaotThm85+27At8wGd25tbnu6Q1Yhe
EXTZHxgVbRMIHMKzV+JgJEAUVR4ZDWlb3FRuIGcfyT4vGElgw99g19J1HdV7QfCa
tAMNUs6vjL0xHhNszASi8JrApu/SLt4LRte5IPqH9K4OX8Sd5yHYYV18EvpaipM2
PfwRC8g5ZKKFvbuzxJX0BmyINWpgxl5lNjixVr4YzEvTsKTzoG6Q41D4hIhQy1Wu
tEZU2aU4v8tY7mO6RedVDkHtRtBYzZotMH0hvSPw79jN4S/JExBkASNR1H06f1BA
/X8CD/RWG5QOiuBSZr9ZikFW2IEZs+HgP+hb5YRj47Bqa4/y/c3/x1zcgQvvBnJ6
jho/iJJIz63dB9rFe86nMUOeWtfmAOWxPAwzfgElb1rIBc0nqOqBCS78MMP6x1R2
Z6rbTvnE5jtwOG1unXADBC+3fpdKXQ2ITRtJej0ZjQw7vi4usOWTSF4GVieZ3ikf
7RMtqfRyF0v4qc3zAjCFM4EYXRtg6B3uOWWyqoTYz8/b9HrG5W9kaBeOdu6uzZnq
Mc0Q3NBUU9lz4r8kxK2r31Kt03Cb7HkFh71KuXxg4GJMCxJaIvui5A9EP2sc1gMF
GljFIXy4j4exc3kJyxvby+EmnnuU5Reaa5OnBkPSemElBkdKrHi89OKiPsrAxL2j
xxbbjw6dIcTzSYnSNfkvGbVlnIzcTzMG90WoUF0RwODKZ5ygSqn3Pms7+IgpN/Ed
Vm1s6GJHx5OUxJPY/Qe/+c4i6S74Kb8wBOtOd1qevU7bOWsY0NjEJG/MCd8kRy9V
C3Al2Z/dsw0IUKUhmyW30HVVcEoLuCcRIRrznrH/CIHK6nhbpJ+Lw4pmn+F+H5L4
8BaG+zG8xvK5Cjq0Z+9aKlpeHmnDrw7exVnhLReSWZdYnSgW0XFIggi7ee9sX3PK
R3/NNkN930yGXNGYQbN4x45t+UUUi441fxvBBOGn0jVjXyZKKGaICCc64MgTZh2N
apbj6dLPtIMx6F9zSrpyo+ebILenYY22n5zaEgkEigqWR/aHZPPwtnGk2qOJEkC7
EeNF8cErlxmj6cK7A2IqpWG+8PYkU9+eubvUihwIgywNA5TEhqnUcZq8Es6XfteC
O5zYrcGY30uc5HK74x+kOSDifEPZ8gL7OU4aDmYoXxH84/wOIVYQIKyoSD2OofzC
LCAQXSVm1xEPtoicMTW2UTzwn4FoZvKWitcSuUfM9qbHSp06sPtSO+kTObNuhUAk
Z46yBbhiTMjALvgTrwSThR0ZO5n0688Tds89QT+JOYAUPbaXRYrws9B+jD5oXJn4
96zfncAkNq/hj2OEjIqOe4k+j7uVaNQM8tbmhZE7R6vPQIAR6X5/OuhGusNX/VVA
yUusC82wMtCp0Ar14pEJIU6mLB6JTdErRgRrP0Pj2mYc9PLd0dUu7y5MnpdjusxZ
e6g4ec89GkQvqWfKPAW+dqAluy2D82Lyd+Gju1pmFdpk80yfWzocDgivcFlreL41
u7u+jLU+5CVTYzTblC6xhG7H8wfAUPlvTBZOyPlZPnIRu8Wr0lWEsjoM4lTkVgSQ
aqZfq5DtGiIY6qRWq+w3jpuiolutCLa2YjzysDGkWXzrbQ/ZE8RAfsYVPtIJHbem
jIdTzuJbRR/60z7lxWd9tz89HlA9CLfBrEtqOPUHVQfh/AlGkb0WIljCil9ntPbQ
HmJsLPtbfmT6DNYBWc9d3ePEpahdTq0e5Es0pu8quBufdR8aPRKd6LGpPE0Xg/6R
G4xqfIzuXmZ7NXfXEIorbvhucH6OZfWSc9Cg36dZ+/THWetEciF0bC9qov8PKgHN
4A9W6u4M0Xn7zMXDj01r5vGzW158n/efA+UAHWx9GgkcuqRfJ5mF8o7yXcH7PfLl
ngUHxzwIhTbZ08Zr8ahsNwFXOSYvv9tNfiVon9JreMOdUdhgk5MZeNJqlpWJYGIf
4mwpWmNPLF3yFFpaDAwRdVunyfEOUbraF3etlDs6nLVPlnLD/egf2BGTlCKnDcYT
B7odE6KBUg1snGrKA30J9G2k46W28adtRSNhf0wck6zGuRgxsiTFU1XdzUb3Ot4I
UtnAunykYHstmJ/imDr7n3aLaiUC95DM4ni2vTh5DZ601AzrKIDJ67NFkt8xfckx
6QJb1RPkYLX1sXrKMS7oOX0LC6wJw0ONwB83MKq++zKh767FjlNlxhR4pCQyHmj5
Oy+UlpsQbVxuJ+QSiK9wvf8kp08A5YYNAvrvRGdCiWPWF8Z/usY63oUkiocp1YRn
JutIl/X8sL+4GfuDs84rIJX9C2oEUAMQPw26MFO7aalH2uiIHWKkZ43sDnfbI4CU
73EQglsbm6a2mG6aWZKHc79Js4D/nE+8atBc37UiJDtQunKAa3oXlFDHdno7O5v/
WX6CTlnpkKjLwe9XAroKM5PgPkE1z9Tk4aIBY2Uf1sfIU7XeEFf1IaJgcvJeCXtx
I+3LZ5I14jHG5V7YobuXU3tLdhMuPH/jAJESTZAU5vwyMyF22mbhDJJC8ICCkdf/
SgL1qidkHC+/8XRy4C5HQGraZgpqv+GjO7NJiJH4mxhZSAfRx2O5s36QeJhe7mCP
tRIgRWMmFm8cvFBEffmLqtSs3uTPIeQu7Ys1dbHpqSWZ1eEyqVL7PBFtOA2gAIzG
6mN3pg4eAVKZiG+jMMdfLGKP6BmTZ/b+wxVSEuj+CtlXpew9kENIPOPXWV4U5YKh
/2RilWVJ9nmsiBWBuzS5zZA7Jw8XVBWnc103KZlO7UXq33jOJbsYtLPR45D5dCGg
wq+B06YsTSAViD6FaGpZ5saMrGlyEClto/oOKvH4B0LNGB3asMtJ5SpbAFDZhf08
S1iTb+qlK5WPaCoSm4SNa6Rjc8qjNG5fSDE45EOi84eDp++Cg04k4RjNc467bp0D
1Y6n4M/q1KmcV2AzHTylvBakqYr6DTtJ4lk19rnlUUB5T620JppOE7kbF14pp2eQ
nr69Sp98Y0zr14lG6US6FAYk65WYXhYZwbX5Tgght2uggIBxNVXKcVCtSnml1eok
/Lt+1QuTR5ZQyukosWX2A9irhfNwliK8g9FKy3xP920OeIFD6TkOgSr3AS+U+pVZ
Z+UZ31O349neT7kSHvClxqS1f2ificgGOPQzGst+KlbRptac+n8541wIl+h6kTri
EJrBQMoDWGUTTixlc+j/3qYvCMDdnNBN5+xtbLBh82x0cuH9J47SpN95KXEi3PBd
cudPbJGjCU2ByN2rQqtR0jeDXzE4+2LKQZkJpMpTeBkbJE3/+vJYnmk2qEfoS8VV
p51mgqpKzxPsw9Fl7LPA2vKjAdillFKSEYGzqGw5WiDQ0y+Ywo5K8scJGrydrYZw
tLmDTXMzhkzWwS6Xzv2ObtsN2cfggXrfobiWRnJEvDTL8FRVpy+RFFPdq1Pmx+JX
Aq+8N0xNDgPzQjIpdyqlwB5Gw0fZm3G0eoMtsIErUgRBvX+Vy7OBUauqBL8PswLL
HZUEFzo19CufFif5Pcgb0BSJkziYbSCcJRB+h/Dvfy6G4e+jVsDEGUUuRXRMaTd1
mVFbEwYevdVZHVxmysWWhN++PoPmRZZyLjqBVCsbvQ3edHGjJ0A6V8RGWw44ZWNk
xwe7X56Zviw5zIm7XBOKXA2//OWxpooVxYXcKGv2jyWviREIcXKH8AWDACEUtHFh
POjSxJueBqsawKbossRWV2OYQpqSMplhdB3ERzi3fKeI5g7M43p/VeoCDJRRSnzA
B+ZUN2U8N7DXC9fpMYllVntKcR7+XsIE8WJ4xDevzxn6py0m/XB9G5GN2afkXOdc
fZUVg2O3KORvumkHTvidDuw+b1DJM0qoM2frgObZARXalhmILXPogPM+otJ6PUjF
6V5jibjtGoMguoIB+Xe/FxxXu4JEMOR4OgAQT7H6BdUhI4qxI0b1GKPXB4KyqXBC
9cUOtKXmoDzatKHHJZ8BpXGxZ1fGblaQ9WqE/mFv1c2WabZGWjV9gAKCsljZ5im+
c41XLT+z/nFZZRKpWls2tDHTUF+dsatVa5F8Pz8hbemXdPVX40CyIVS/N0gYUc8A
7c9f9cQp+TL0ZbXnaBcQAEV+vE/h3yKTWz6bheVHFh4dy0bLEP92cm2g5MeKZj11
xMWwAsmwsXM3+yPKfeCV2u2GExsPPqS/X1heOQNsq9PARMyTjselNYxXE8uy8rrY
U6C4qglyG4PX2SszPEv6MD9v/ARN9iiBVJRI635+Dx/Kjgdhrk+ArbhFhA8Xc0MH
JdbxFsuVtMkleMLRi/2PLoyTr2yX3NAPvvJwK+s7yu/boOy3+b/v5tTnClwqUw1z
AhH+XKDzvrH4EJlAri8hN45EO8SQWd5yIKAi4ygK0Rzy3yfXWT1AaXnjSn3xHYE4
xRFazPQslWeyZ9NeJg9wpmDsF9Pk2am22B7o7Cp5LQmHn3CUbwCfkJv9rG5CGYOJ
ZDRspvBcyVFKnZXy+30JwGP3zhEdJseZihvWIA5uE/1jXIl0j4rNKEmyG46TZhsu
vYn7EtSq15xfLCblK2OiKn3gD7LCXxCkusgavYmw5lmSvH+seE2F4ES472hkk97w
RWX5BwI118wljQWLN9olueU+k1P4lziFbeZO1Uxc3V5VgS4rPXTojGIdnLppO46h
nYBis4B1T/BjGIZ/OANaqZ6DEOFpwRSh+H3gyzMxSt0hL7NlJZA1cRN2M2IF2x2S
YGd1ncKfDrcE7SSNlNbgthcjVA3CPsCp8rskWCWBwVOiaS0/8qCXps6X0wOceHEC
KzQ+32nDppr7GQ5b0rWU+y44TJro7qKdkJy3s8a5jkKBw24DKhDs8pWtCOBvbUnj
7b8OHHy0KQEE3gzeoDAiOZ0RFgyMVf2VJL5TacODiw1KQ3O7Uk5AWA5BDWMjRDs0
f3lSKqZZx5g1DHLxw3XnzDw+i8MdgGMl8gNZEIYz+5TzzsHm9rco+n4RQ46C5k73
KRo1NzhlMJmBKoB8GcCjXfFKMt7SMPOxQo7alP6jEkxlYIsmfko8GigVsl2UXLCb
T5BkBag+lweD3KZq4tvADeboVDIdEGBtn08Nu0guZyPsXKvLOzMrPMYS9akTDWD8
hFnTBO90h7kLLA+udY2MWtFX9oEuhezBYx/CKxljLjYSEzC6rp/Lj6D79xmgj9fp
s6xKaJjvZyMbcDYqEsLtnyod87ex2NdbAjarTY0MThhBlMk7zGj0n4yISYcOKg3D
804mNwZrEqWkkVThEnsT19oZ2XcQNrRV4WO7RI63R4OLhmaUK04TWXwBq3Cxzs/Q
C7JY5+dbF4H9R0ufYL0xr0qMeDdxddyVZ/3gl9Xrb38jwKSNUtm8h6Zj2k8PPaRq
6nksMjoDmROgwRMdM6cnmaUFEFw4sHSB/iv+FQA8oO81IDJtHnBNjIkcEdFQj9y9
3m9ybBEgJNUPrs+t5GsYTOMDWOb/SXd26ERmHPAsqMNw1WVj0sQXpFfnfLIou2Ls
bqjorBzEDBEfA6tCGwjVQcmibUew/CX5IRSg4SN5IQz9gK6VQbHMxqvjsRXLM1sF
iEC8DnTQNCU5+PeF0DnWSx1ykE6WuD0meDQ32inj2Rra2xS8F9EvXEPOqvoO1r3g
YXDb+lSrv2TwgFGjLETWoXZGJ87KAmGeSCRktO2z50MUYtFIjM+uKO4x1MRVNFEY
OEqjodcql8OAB/g9DPBzM6esrwlf8EylQE1+RvuLtRfFlFgWkdS3Ia01CwsFlusy
4x9veoJSFAjNYcKiGQ6UWhAPnCSEqRN1nUFrJiKBJeQDazUQuwjWvrugGRgs69F3
0aEzC8LnToHBGJMftA4Xhv2s7+KY6lyjJi5uKv6fgdN17XMc6MMpl2KqVN3NAump
A3Yl4+AbdiFRneWkJA7c78ATxw/Ew21GYq5b7y2QOZKnquf/cSGGu97mEJAELLKi
/tVCCp1rWI6tII0CgIKbONct6WCu4n302kq1lMlQwrTo5bko6oLxua3J4fBbLwcx
6/gTtaGmgrpynZV9qTsQPOaBCUKdHevCupAZd9PrBOJlWgwi6r7PAbhc56mZdrge
VUGGD6FwQXxBCLWI5HFLnbTMXlbbbEjxCdhkhjmFb7of5DmpRvGg7ePXJTGkxK1V
gkx6jPQYHlovMZK9J2AnjiHFoBIkjTLDnWuW82JYSAsjuXAveoLSDTEmnay92kdz
uB3kcRbRDxnLj5s3JxI/NY4/xXuliedUoQDKAPEkDNIVEYkmJZ2usQ2ATqJpYsd8
XLMg2L3ieLZfUEIjpAO+KrUZ27pzbJ8F2FFz91KXzG+tl1h2MzX9qt0I45anPgFk
utunRbkiMCszZahWXmUrgkrqM6devOTiSFln0tY1c2lbwM3pY6W1FITuss6YxA4v
zEaF0wzdabYY6Yz7L7iQHndiGJcGdi3nqpfZ4eMRqGz2jDZCsVquqLeOYl+EEZzv
ExOtKh1oozCDd7Rw5CphZ7kzvHLt2KKb3wFVBcx5bI0ZIcwOSJhUSd+rDWNJrAOe
3bbMB9nYzbEMC5icNfg6skdA7zIeB5MldgyfJLxmv2/rkOA/t7Hki6PeturNAjer
S0O7mhGrGIiY3yQX96szabclwwKnXXfdXaqA1JYLci9YbowjJiPV04zffsX54kt/
HKjrkEqssuU+hxgk6dDaOgEpCP3ZnnkVGpeDVwwNczxiosaXIol8/lRhyTGJDUff
QSghzwqRCAs1Rd3KhOXk3z7Z7ORuAB3sIchFug0u7n9YtGcX1XwTuxUjGEm+wl57
K/jknnhaOPH1kF39ZQe6ywDM0urexWFH2q9qM2z/4xiWfxodJfiysn9H7igzL7Vy
SFKdO3OCvxkdhpFECWl8KQJ3nohKdd/YQkLA3Jwr1NRyyXlq5IerxM2lTXGRGOYR
hutQ+J5B7MkOH4xyKv223TdvgN+9k2NEqiV9ySf+cYCMSzLBgsmLqcJ0nHuMZS0t
IAYTCswb9azpT5YO7+577uIADbdl0g32zel+X2MAJMr05sMUMZmVxX014rohlNkv
gdIVtsazAISDTQfa39U4RLTmymXJBkTapr7sBes4LYFr207iQTZ1If9Bynrj5GVY
9OtJSW8Chr//vYMC7zsvKbOkFloH9MPEJHLn1om+h0ElnzWwW0RzZG1hiH8frtwe
hJb1N64udBqsWhEpu7NXaF4m9AWNGBIJWsUz2Dt/dZDEIo8j1dnmxT6GogTw2rjY
qPUXbX4Ce7LNJCAQDtTIQBb15J1BpDU8EQYRR+X+Ku5Tc01MI7nKZQTQszRo3bFX
P5uqFycS2tk8T/XsZ79ZnvfYmHQHC/zlJxO23GOUDmDBW//qo8wWTgmlyN7QIZ/u
tMhyP66Es3aR8/NEp4prSFnsngngeep7F6SwAUIIHrbq0tnFq1KkWxxVEGxnTzh3
Ve/HFzeXvDMlLA6Z23q3ZmnoZkaReCANWHN65cj/KhaxJpK8J6Dj/h1vp2YeX6jI
2rbycsmDQhQAD7POPuBrmIau1I43onc0/rm12SiacENE8Aj5LOEZiYTSW9EEI83R
N4xPqSeq/eS/MuSmlRxTBfC1zuLu/h0I8DfKm8Ilog7bgUBPvUyZ87YvWX8OChR9
4pX3aP7vExDLcdH/JazwtbbZzFhEXAqLdxB04jftHxW8i7fHNyCcoIpY9JSYPSWu
RMC+VsRJRprKcjx5nVmHoSv9TFfUBh68MLAPOvPDbMCEEvgXTK132T3RKw3k8nJu
4o05LIqCvIImF0UX0gXQ0NtZteZV7OuH4uWzi47hJMjDvxQs8Meb5XiXHedFul10
2Z8ZkxVZSs+NsAAygOnP7YURXBl+UMbBhdGQmCry1LFKc8dxiqxkWQ4DnOt48XDk
SmKJJwGEGZPYJaA32V6ZRtXCadNFp+7ad/zQlX+DmUEDooTXHqMd7OcXQl5Oj2dM
TNx+J8Lp5LdF1l3tfAQ9ZezuLVVcQXOKDxuHVoyq9e/Xif9aGjmMN+HZ/Iw4xVn0
PcYIepNR+mkC2D598pbM8LHCB6BAo8QEpzC7ZnmKbG0/nX/VbwYECa+VEhitPAhj
GmVp9itz8wMbeIcZaT6wXtM9Hs7RWgwIytB6qoBSrFXrE41AAi69lZ7w2uwXa7u+
at0mfrOaKH0L+lE6JNk5bvuGFDhHf7zAC2a3nMxXjcEQ/yXiYeNryU3kBzcf1IBX
rQ7ZL+rMjo3L1QzAc8/GlHfKspCdJXgZ0i1fPL9DhGtHqgm9cq0ybjV9iNAohAzL
RdsxOmQk92sTpKZ5gqO0VFtPC31ElV4xlK/NtQ99GBB3bQkPWBHVvRJuSK2Jzl1N
9bLIv3P/IHb7qDIkg/YPuH//116BaWtrOoevrhasOOBPIy3zzBVNtezac1WHNEU6
HaGOGGMpaLJsfGi5fo8wq2eb55QOgsP7cRV390ehhwN4E5YEsfZQDv6NFuJebJQW
DWOtUaNkCJ0Ou2xkcjujmEkaopX3c5Zz9jlCfK/I+lTM5vgQJtg0fMWfJeg9LXNb
PJeuxgmxa//ezgB2X3h3EHLcFwrUXb3bZ/AkJau48MIqZ45RybylPfpQMUh0nE13
gnNNorXX+Ian5DJuPDPukjN0Cbx48zgoM3QH7QbG8JUVIEInRy+owvqTqo6+UfqD
y9WNn4Dxp94Xo+Q+o2iknOOG5jnGkU7aZUhUiUchFwRVtQHsdxrColkCuiXhiNzv
eGUsqlQM1hhRn7tm5FpA2A573lRYuYkMaAEv0F6fZ5n9PACpJm+MaOuRw29XIhPO
R1kkqx7W3i5vbCO1Tv9WlfJQ4N1XKEdzMnlAR5hkF+GN2+oCFWbArIS8isq5PxIt
7dBFkHJigYwBLBcn1CUjYM1fmJfXXEt+dnia0sH2jrl/R7UlmkQLmGBU1ppbpW0n
XRUXqaVmFAdwI73YGJxx+S6UBNW1RwPRZ6tvf5WMkFSoMlUOnZ1ub2CbbSKWQXpc
EXKrSOjayn1nnVMXto9cYHGNfEgHntjf/CRjMf8lK809SfZFlaD82WhM8bDxfJ8N
d1gZxL278tLfTkGNFSZHhwWK8DHUUmPS69LJ9j2R8mmNeoo0h/ctEK1rWix5AZoS
DHg7n9YIQ/QPYhzCupW0HgbRthfbk88SbW4tqAPB56xp9uSBPoKpQPCqgv9mvm7k
RfvE9KWsDM/LJUSbrRi4UOPSsBH2bQ+30U20KWMnWAwQmSvEY2M4z6kwWRb+UceL
IgS2dE8ycv7zMPMe1ArwAlJYDws2PPWCT8HSFMZvYUXkR/mrnyHlS8jBl6quu5su
FSHjIZSHMtf6KWhUoN9l5q6XFrjvALQtOYmQw6ZtcWNzj7QPNJRn/bI+TqZ68ALp
lXub3qnlBaiySJYHohvWxtAx/mx6zx0I/ahxiw2/8IOxn8/bZkFpNDoF/Qtmc0/l
E0EZEf/jjuFoH/X48z6cRzdxU+kPohFhkyP2Q/+DngtqhKGFvdpQ91WzmfI2C4ZN
qZuXZOVO5dyw+cnbmG7Nx71Rafcloupo1+gkDg3G9J0xBY8qFGBhMdqrO4KfXhGI
9tH3X+Uhv+exBh+Y5LcA0GA9kp51XUJRwnXprqDuT3AIjsUFNcMUGBeiJw51nQAS
y10F5QckDyI8YhkgQC0QfhfhnmWyYyaR8MpUl5I2wSMb1JGblnFl+DfYeQpNmHRL
TcnROnZxGh+zQWILAA26wQHdNT5z1avPQrWUcl0i90M6uzx5V8T7hUv1zpt5zcja
9IoZJHv2n2qzxxf/Q+rnc7oe0TdDS+7w3ATsoyxywiIwAsGtbBbd6RDl+W7AqfQz
3Ov/EsQI5aa7M9+/4oNWIRCpP0/9eYfZ2GJeZd5yc7TVZhjyLOc+0ApOjfWXDWtv
9s6kBjjOUIxmww4zZTUB6+rxLG+5QYvs4xEXnwfUSlHCKW49p31ubugKK0nX8YQb
O79a5w6sFpRcceN2U6PJMTFnxiPqR2pjCdiO0aKuZL5Qmqo1K4BBnXD4XlJXFvr5
8QWd2E1vJztW8gan8PIZS4ps6rhmbl+CceXnYK9FkXEW5SJ125RhUg2bQlNO7jSK
frs29+f4jmD/wdn76LTkNcR6p/D/Hk02cCp2Vvu0CrmB0xZUovmKz9sItJNtjpOW
JROjHCI4HbSzZWrdXSwQUlX8leZMZTgPGh8cFvZ5orwCdYgKmyy9UGKrQ2xHhpci
JVPux+8b8KklAofiYaqj6zlSCFoXhqLm6xYoJJS80TgRSoQYPeod0wR1+BNHgbHX
l5j3ojbEtdTwzqo6j0WBK7B46wLbyC7qYo5QpQmTbnX1dKrnT5FyJSEMeduOcshB
xG36zvk6viS2nQCc9D7hRaWKucOTFjRWs5v4UJEoI6SqR76Q1mX23JWlbZtokos+
y/6IdrfY9l2vBvr4zGM8hqn301hlhUxYXmP3Abh9JZVNg8xpAIu6F+QvLHKYSTR8
7h/TNdKXLVX4BBLIxXO+EMUHaIllsWZAK5cs+qtWKWgs4AA0ISZ79Ybs0wbLW+wl
tjduQcZkwNntmEkfP3BMcON5QE9g+CMUZ2HTDqNaq48ALt9vML3LwVBjrrdIru0c
h2KfEgxMRXYKFlXIRaNu2lp4rNPzzDIYamAySb5xE+9/A5nEdAgpDmWhF8RgYYoD
dVXhn7Z1PFnFvRyKKZRAaJyn7/cAi8UFfe+Xl1BGn7DsoCJRfIQCBo+n+6vhs/4N
NuNkeKKoFJVc/LUMiKVumtv2ms9/Nnplrhj+dnp+dKarSjMw8KB7jxxjk2iOD4CG
dTBR6qEsM1RjDW5jPpMdA7XfQ5PSSJDPAjoNEEX9VIHm4pb6liZaSgPclNvf/CVz
7UQqlqK9ALLWTQwueOdufFSl4Kqjh+IRbahkfSR0ZsBRKtgLjuh+Z3nw9Qa63h0Y
s4HXYsY50PIsqAmcdg6GuuIgEvF2J/Y2hGtVRAxubQxqKl4pPJ2mWk5+8ZEjxvGq
NA3GxmgQaGnsugECRZuP82B47qt+nVAYsPm5AbEhLkie80xLKpSClBG1le6HWw5N
0+4nQgC4bexpMnw7uN4M+E9ozHMaMmZVFiNnWsNTsNdNBqCqI29qx8ef7ZjqOHtj
l10uezKkjSImRFJLlYlNgMcaPSc8ruLeDLMaZoo0kv9dnx554Js41bo3sI8Ragpf
TM+ylVs5LCdUzvJSEDnH7Q6oZjxWT/1HfSfk3Mr2y3yyoY4Vie4VRduPh/fIwm1u
SY0gGTQQv+jUSX2MYDb9qiJZ7Y9k57nD0rz2c8kTK9XlYT9jLPFNkTJ725/nP76G
ZUmafEe/2bAmNp7viOTTphaEvhVbR1ZG9ZFrxWrHn5dH1pfCObADxCLH8M0wsYHQ
0r4qgpqlxgtPwGduE3POO/JQXzfYHV8oGbYhkcSMeVJmibPHCwKitT3Ar/V7aOzQ
Et510NrcavUvSombaRBHyJrASsCEbObmJrOVohQm0w6i23CKPXNOLCm2oZZetEfA
PPHU8syYvyPHElFVfPYulsSPwPVvi/EHtLwh9kGITBrhugCwnUm0TgxS2sEag8U8
wuaIwIAXeVDWz51RV/4IwGTPWHdUbfe4l2JTl9NH8XfYJ9XRLtnLVntipmKXw/4Q
Gnw9XuU+v+tO3Fy88vNOBOm3CzKqHAaiQrEMIMV7Uv1QPbAwYLfJJ2o/eQ5z5TfU
Ol4TzVFpH80UjAWGzvdW6yvGm99FaNB7aPX41+GwUHnZ+Dze6jtm6is59S7alEnI
+Fmo0mvoD5wTkilBw3TVhP8OnjKPb+Qjz/L28NVElfYzBXXW+rLEdxgIIlqM98FL
GuaVWRU3yOiUMSQmdsGiFFkc28Iln3UUKuyWEmhimrxrTnTj94pQefftPSnwDGlM
Wu158OumQjoR2w0/uCYJa9E26nNlPjMSKlQHsplnJH8Dx6tRml1hAlLtVfiKZBHI
xBXaSrAS4nROhXNjWxniH4Pef/a//MAQq5787OcLAQBw1dI0c4gkmKsU7gH0k2+N
4vEWkIexdGYESXUDGBCDLmfWvVfEZ7o/assnduTDeIw5mNpKeSyg8dSN2rHKlthX
BVmrH6pP0n8OTCs45oQgriF9oynnJm6RHwCg2LQcynab4wrXnaKWJOouPh5KaqaK
ZHS5fjn8Se7pCtvwwMKW69s21Ff29D0Wqi9cXleagb0rU/VOGbofPSrD80Ao2loC
Iy2AUYchDrqeF3QEEVP6AEOPT+na+0uqRaD5o+maDps2fHbzdIIUYDHpTTLBHVWL
0FoAuyjrnGRrmTzIfHMiEQRZWh6eDvqRqelLj2Vd/sIQYNz+Lih5DsGecXTqRgj9
Ik957Y4wFtEXMxOLPpbyaRUSdL7fBC5Khc4M7ijvUFfZHNpOgnwAUvfOUY1qMg77
pTKEu/hPTnnGKVMbXRfdcPB8uNdug56akrqVCM33X3hrIH335Ct5anwaglkFNVpU
hOXu6CHu2LCXh/mjvFEG7N63cJ8JhSkuEut5Wcb5FloCMhqM9sfoaDSWEqTu/E/1
MJVGNyCFIllCvUIwkD/O2pnF24seX7NurQNVJjufYzwgF5aPI0NJLp+/+vuiJfuz
zry4lDhRTnEthcYq4BRleAvQ6yk1vKbQ89MxGvfYE36eMWhhdX9HalmNZj9WCzr7
ASe5xhe7rm1d4M4klzuHFwqTJwcIRAnHXFu/FQ2W4OUOpxGxzBz/Gwo2EkD6JZgX
rUByg35HP7xbgpevehOGNr9yoBwNKLqd8/oHi/VwC1N0tfvUk0B1Fv8NnHXO3xcf
zBYci5Eg+iskOdXwebX9DkizNF6cTCK0mvKZdNWozrMSe9+U6FVXd4zQTlCST9GL
mA8w20ez/67/qwIB6hY0Cbk+gFiyqUna7AtVGzIusGBszpaiJZBxMMTy2i4kyYBO
Z1pNZyX5QWzyz5PnEKQnUSawvNOH9bIh9YEp3tAswKKTXdPS4fDAYluHqP2m2tFg
PgcSgX0u1V/2QYSNcd7zODlKNiYbxc7kGNDe8yok18v3YnRvf498C6LWMafI6NOc
QpDCgfGi+KNA2XRDiVWs3MGRc1gXroyz/hO9XMuns6kqyXO2hl8e5wmy4SrcGt6D
6ni/a7gRS/NBASITxbQo3ZRc63LG3iQMYIUDv/uq9aaHctDSlrBDtMGCF+MJyUg/
5+JXitMmDOK5EVVR0L6WQGrcXXY5PVjOlTT38NnBF+r5Zk3faEAhoHUrNsGVrgIt
m9p8jZ77KWWZVuYiXWPWJIKcHfkrFjt8MajLEUV77Dhx9h1uGEGJ2PjLeTKz88/l
ynd28IRWtj4Jy3evLJCaI57TYkWizd6RWopQwmcSHqB3SEhqnPQ4EvZakw4+A8hU
itwqr+zQ0yfa0B/ex65tcJbnwKwgoeYpv2+PMV4TE8nGeY1uoQFu8xcVkmbsxj1q
0WB5/XP3oL/9/yY0ZdliFxbCgdT9nOt6Y8fffsc/HtNcUgYdjUtUT9pXTSahcuLk
Bpd/Z6vVzlBlrXkQXRAjrCKHByILLvsUjA1jpZp+G3omV3hnpNFNAe8S6kOJtfFv
Wnl1DWpTTYmBaMFYRLQZwvuWGrKJ51eDSU+PE1msZ8djIBvH7zaBYtyi3rE2AWS5
yMCTBMyV4WAs0/zWWFF4NIQRbyveGm8A1WOlILAxYpgOz1fd6I4dYcSm+nZlSt6e
u7ggq0FzWD7TPSHCQPZRYFq4YuL0NnHX50ke6tdeKFm85Nv7SSf+2feLE0jNsoLD
tpXNjHP8t96CcSidb5MLYH73F2fMOfX/npJy1voU5BFSzPqSRSVcmiXRnBMA/005
nUbl2/f73fr79cKcxRsy42Q8CBa2aXTUaqcrsor7RaqdLZPwS94XZ9G5Ms9Rw4/Q
kMRIRTiuk2MPVHUTZe5vF39w5CTAEwWBQcrz6m+ol+YEF8J3gXiwyoSQb/RKmwR4
meQIoCuyEFeqb9ZsEDmNSTUUw2JWWQDibwFJYLoCfQs4kdonRa/hs1VMaxSBLPmJ
+hL3SducuCF8c1/kK70WultAtok1T7/t+wTKXYqENnIY71IzUNuRa3Et46nPyHCr
bbXYXKV+gfJS6LtW0qkutkVoVRawdWIvK3v5V3T7VDJY6b+9quytHXMLOYAH9Grt
wXeNR/6C7rDKVJK8SKI79dZQ1Mfz7GUrZAPipwvsrMzAsAhyISvpdg/u8ypXDl3u
f+EEn0J7mdge153PQNI++EKJM0vB6tHP1CZJTToFZF0aw68H7kyVQvwjLDwcf43I
fRN+GIdcDHOcQK23zE9bz3sDxX1ZPU31Z/oFgXjM5QpqVX1dvWpIQ13j3vBKPQ/9
3Pj0/MRDzvHo+0ZdyrDAreM/5vJE71oyfp7HlrPln/0pRgGY9r8XJlE4ZWqy8jlW
oGWqlj7xrxfDx4qdND6NsQPcvDXjAAZajlxuP4PkJM6+ZwQlHreuj0ojRXlzEASR
1Ufv0uFUhUPmLQouEDEelnYFeRq/8F+BceWmufz2mRF6PcO0jmtpxwO+9NcjifUI
ikqf5BhXC7vAurilnUGhR0rkwbKTQ1BNfC4q08/fW9rwe/KyXCVn7A0EGGbp2sbu
G8ZiRuLXt7hYXSk1DD75gbKBKSI1E+DJ3JPfv+3jRYSHiHV8lZUOAJU6+zRp7akI
hTP6yU2/qJ2rdNC1uxTc2PjYzeflCMcVjDignJdpYxEVHeY6mSHimFplth75d2Xy
axpfTdVumdyO3/A+RiAp3N7nTLbfMSYyyMEab0rXCKsC4bMTl8ZjXgHu/+HWVtsI
fSXgwSylgwXDNrrTYblLhhap/RuVqKYwrw6aJ0WBkpYjhScnDm4HkqVHD6U6pezW
pu9M7MIuS+uXAoKmPPPgyI+D7fv/tgXf8omcefV68tqaevy4BTVtA3fVcmbMzO5c
h3LtHta+LLGU2xA0/mu45wNE5NIeAaXMvVvbvcNeLtgWBIU5OA5/Z7Cdsl712qWv
M1Gb3leFuZNmpW+BJ8t43vZq3lx3HFZK4hYGye91xbp/uRH3huS6ylHZyK45rRVA
zF4JMClriWN6+fty8u98NPsAVb9CC31fH7iT7mP8qc8XMTidLXscK8p5wx3sr/S7
TJ6MT7aTehpEokVQ1vb++eNf30Hl/+PVd+hsibh+Os9arKm+2+c3ivRAVqrAwgYX
B8zKYlErrqb4Bap/ZanxOIr4kx9g/z3hatfHj6bPx1/sA1BMQbLOugsl7j0qhqoh
kA3MWfUF/BaN8XUOyCya/XaxszJDifquwJFEB/VlgmCQ7Y+lk3jreYQ6Jmy5Hmrm
mHXWmsRpqggocBQW0rs8u4F+mlQkVqjZ9tmYTmZ4IMdfORolrcLKBDLRHmWRO80V
OLSgp+WlEDfxAK6mZ7cQmQ8YwcLTEvL4ZSOPxyLhezXWgi/I1rzpAfPDKzomcZzk
L0rudvxLw1Cs3ZdLCLWyczKp2deCdgiUaDsjD+ZaykXcR9cg80VwLV2kmt3zU6WL
tfwV1Zy61WH7O9ux/aqSHe7XveUsbOMsrmTP84jQYqae1yMV2GWdMbP0h63MFvZ5
WZ1cQYSKW3LS7Ot1cU1/+PYADW27870aqPQswmIC1g1TbHsTArFEg5NMNubiWHaz
Qus5NZ0ZrdPUgFY80xE3lC+EOuSVhoVjJjyEZLdlxESCQdWz91yD0JTKFgQVDw20
I+TurRnjrXi7csHQ14SNYJLfxmwJ4V7pYFofYHaCGSFwhxnY6D4OjMZlUOV9v2bC
B1VgOZNCPauIkIW1lEZEL7WvwOOrSTaDbhOhwg/tWQ096g6EnvaiYgfiGq7y41Qm
9WCWKsf9mfNQiZXFAo1MTZqghTMlqCcBGfkcILkXVhRm+jqdgWr8ShYHivBkQWep
TT+zpw61CCIWEuNH6qzGcjxlrd4bQ9NpGSKLiOQxaF9j1Og/wpS0g5T3tmNmckMx
fVRB03f4/wIL9D14U8TOc0ubnuxEUUKSe9ekEbImgoQRKwp062J1PpByntqv5Qjs
lNsXhAVVzVjhLg+L8ezazLwXoM4oIQd9GATTyX9qIvUvx193OEmpe8rIjyANO1h0
iNVzUdz2PtLMVBlJPR+K6z233SAmPxfPT7VX8FDjcF1CYnNAZn9RDG/vV507iliW
TWuQkrSAPh43gGUxiUcddbQHWP+X2O7BA0eXKFb4r444p0WV58gr9iHvPu/GESaC
oue8xnBVxQtvgAjCskkLmjFk5DD+VgsiDMbtN67bQrxEE6oBgNARf3UH2hLSFChD
oFO3i4ArujdayCjOw9GoKolapz9HdzaaeAljtwtWVrCyY6DJzmt0us6prtbbOouw
JhWnon02ykYyYyFxtGaQG2fqLP4IY2SUZY7jkCt48ZkusHLRYrwtZGK8NLkh/HHp
w2HRdyzZHmXptYe/GCnfSdc/ZHQP6Q7NKO32MqJQTRLBPiL6MKW6XHPrKBRPd5Wk
IcLK2Jcw65DoNHDs/yd2B8AZcKk23xCqwB/qt834w5bqH0ptolxQQj+juLseUusK
+zXgfXwvlyq9YQ0cUwbDtLOZieGHhj5/W1qXYzF1T6SLDtpybNxLPQOoyfiOA/bB
euuT0jLdOsxA2UYhzbMQcOC1sQbHhYFZix0yOQF+aET8e4cJVdI4il1eAS0mGCAC
3Q68VXp/JObfeso9IHp+wo8Psuv3hqK8p1FgDY+GhyS7wYat17AixdRGHhyBojgI
32M/MkVQmhHnKO3kF7/fSat0cmtxvWASk4nqiAdSieOJculLhjfJyyI7UeQvkFsp
oLOHSgzkVd8wtGs8E1Nc3kaG7sIhTiQv1oW6zMocw7sWn3WHeyjFO+1YorIRn2aU
63PfGKIJ/BnFF4QLDC5lfZrw5B1TMu3+nyL2k5Xdrfk14w4kE0E4tpf2dLAcaZ6W
skFrgkZFoMKLBUDXRB36oZl+wbxuFe8lJL/RzTLmPhcEQTYP0AKLQESF/BnFXhcl
xL8D40/hExSuRzKrMdR10MmlZzpSeCrhgcDdLi1qYV2hXvzzSv40Y4oeijpz3ND+
Mi2HAPqYMiiJQrHAtBl1O7Qu4voYMeZT3PUBo0VscXe2ZHPYB2Nv9fOWRR4+qSlv
cnTWWqmRuVZQjXgo+uSWvWJf5IgUBE81ezMiAKJ/7P1UsKDIV+5Oh/zizMXNEKD8
QED9tZbQLuBmvheHSIVJOb93kTYgQOZGFhll6KM6oU0LYRUmMlzEw/IG3cxWmRV9
YI6lV3AjKtdpZff+gHcQZgOO6diHi+i/UpTYJDFFAy052aQf6w7sBFfoM5jG75RJ
+KCfq4l9YJIxpx/df9cyveDcfkGC0Qbo1FZvcJjOqXT/qvS5n0nWXi8HsPTX1XZ6
ap7NDHSsUK76pAVvdMw3MvX/arzD/l/nZinMsd8OZEWjCzeDLlad4UPp2m0hhPO7
qn1oNZdswENQInnsdObXrS5Hl6N/B8IdKB4V515RwCAEcoiQILM6Cf1cMIlCrgge
7gARi/CbID59fmoTddU0CSkN6i4aht2dMocIpJL4BdlJbs9H+5ByVj++2eP7c6rH
bOmME17PkuhvF+PJsYc7WdJ/xFKtkodh5r3JZ7UB/Q0Laptaf367BeXowFFeNrnE
6eZ/ZXknKdeLlaK4wDlphvwFZfVj371u6wflJaVfKBgECleB93Fd9wojaCkcyYKA
KuRWwzPu+TKCvX06UUIdVaPl2bejK+11a1nFLKstV6BHAbt9MnpFXo7WTvrfwbjf
HpTQxf1hVkwkdrqzt9nkAXLjtcU3rFPiaKSr+HqzthaxHkZmuq0t513XSS9LT7yL
7mvv6bxiDIWzsYprfl7i+F+SjWVwi5OZuWBRZqrNGqM5FsPYc2Tr6bQFO7Tbsw95
yteIETYZKGqqChzDRb+tgosJ/0wFdlgwZw+2jceUWdAAC4bsSSq5yQRvbIqNkARy
smJGf59BMVAYAKs2bjHq5mZR+fakDqgElmpUWSWaGGRRQPOre5XUdXwhcT5KEior
a/6k9wMb/xsCvmqZCPujVaIBazrpIDrb822S6HrJ8AFNySRxbcv3B/QzDx9gKZln
QBRX72YLeEZI7dzx5HK5QuJWzFF0/hIDqkbtQYwTSZAN/Laza1qBbLMyI1J5fcdP
aBGfS76L8Y9VAgySByyNeF6JlGKPgazRtO6uYReiwe0k32R4cDrT1TIicFZEqgLQ
lHOPEr6BZora7H9/7/MhqulhdGt0la/JaLGr3G/2xtfPZlx7qcdFleEMxk4h+6hU
ISptq0DDt21J4H3y+gjmq7m/njIzQ8VOs6tojrW6j8mQ9JulePaxseEk8qaJKABx
JiFqySx40Zm/s/tt7Lj1hNNYUCLAdPu4J4yIOVXq/3IcVUFqJEUswNziXqFOo0ge
W6krihPliPQgylhul2FsmpURZ/odEFH3btmtvXfLPA9GwfpjJZaIqe3Pg69zFBJE
3IF5ijA7FSSMYgfC3EGQTnItjh3F+s1cHEsATiJ2P2yUDKhqysBoOosL4R1llA5u
gHPu7M1VrO1/SuwKcjqxO+zsIvGqeGjJq3SVcWNp3wzdhqT9IMxGR6Tkq3n1duOx
RtPY6Y9xr4Bzu57KBmPNjjK6AhZYbOCrMNNRCQHr/pf4N1xhav932HV6TJRU36fc
a0hZW8JHF6AFHFLSYI+8L4252tasVN/vTBCOLOWVGcrJ5TJxxx6aeQFIz91+w7Ii
7tZehvBLk+AEJjjddmSaQ6hLrr/zlNKMQJUD3tvRWSJ8FtpzHysOb0uH6pTUQW6X
HOysfbSC2WdEa39Nvu7w0SP33pA25yGA28h3LA3N0MP3LmYx+PE1ogrSrnN0wSAM
QuQwPZQZT7FeXUowU5keWx39+lCPEXWGSYNI8w/i/siGM+tYl/5yFLUrbIpP3szi
hwdVQEjq4Mg49VmFRbGwQAki0rJuFpQYl8gcVY8bvpQEfoRCKrkr16wEfVmZo0Zt
CCT/AXa9pVi0cAQu14VJfKXnVKI8aWBQ4kh5dyD4KoQxTU58Frp3DyzCtmqnLtQJ
C2+IfkbUNSlssvldD/DRhKJXQhPdyYcTLqqhWjeTRjgHWFfnLipLrj6WSYJal5B/
1+IvJaq4XYC+Z43snvUMuNeDPz4qw3/x2yINfgvEo9YZ1qQ8ddFPvqVdBeY9znWc
3mKV6U8wccvbGdy6ioHpoQzMuvIE/LC/Nn0WrV26O4G5+WMdEvkNvCU9OpTTOuy4
pb8BK29PIaVhwRcXvSxH99fGyrh6lIHf9naybfGdPXmk77fpsUPR3eq7/mUe49IW
UUEaDLn3/9UXb0ZltDrKVzgVI3DFTQFwehqhiqSVy4JIffXJ5uY9VQ2J57mvVKYv
MCDc8pEAxC/sislC3f+FK+Wm3GvA9UpYuBx/S1QNEirasjec8DjNmTr+O4sZNy5r
+hawhaIqzzOfV9bJyjjtR9XqiAZoOE4NUQXDsOyDuiqg3/qtvYA5m3Tk4JCKdu0c
4eW09bdCZffhIIHrogqvNugh2qzJILW1YybMA8Ol2+ziNti5P+qO/e1f9VzgqH79
s8lpiEC48oFZr6D693io8+MpHl5oPUYCtUKrbiuyBHtw0irFhrz2VOp1tetDdBCU
aBS2qYfVr0/z9jNj1NQsbgXJ0EsbEs0DCbK7LZzET+/5gvNK7M/82gJ9gMIQes3Y
AvNOeRHUOAP9A9nl8Pk22iBfFWCTMpKYQLq789ExzVIJ1HOgkLJ5FnpjDPSyUhnR
OXiX2gt1pl31eGJvNJ930FIrpO4MJ+Ihnds/4waER0kE8YqOfVhHAxC5bh+DThq+
9s4ZLc3T5WcsAGlFRA9GMQ/nM55m/6GuM9r/PWFvfGgsAIrDzSAvrNzVLKwi+pew
Xp4c40TkuD/yVXYRp63P01RXxik38gSfaFd/lmGgOodox6QhqxjgP2SMceGhs+NP
tayXuh3kwQeucUywxp/OeKQWhUO3xkbMHe+9xOw6RkrKbDGepCnj29tXR/3Yq2Sv
ykXCvExzLspQrpN/m1Bi4V1ffQ78XxhrLnh3ubEkGdAX15niKh1UkVIKbDSXovvv
Rcf3TnRIKPUBVKovVy4+mryJWwsIAaRtTqD9mhi6qfV/0voFtXz/dC3yMtChkjsm
yUWz2PpGpnN8JtomzuWLCcyGVTZKj16gZUmdH0rifO2lLmQlT5GfCD1D7se1QsbU
4BX6lhcus3DwHzSBSeXChyuT6fhSAEUiBUUfEzBEe1dB6xfeBwbbKdH1jroW+r1i
O4ttxwojUdQNJnbtEC10gWBQHCHzCbCz4FfoEjN116Rxr7F43TwwFlDd3I2PBlb0
AEaHubKG7YDAwoiXVG8sBp5kaIxbH4whRq7mLStl8oJqqibJzjWyyUkxd38SD4XY
rJI73Kb1DtTlmRVUcwATQMNLED2MzAzoCWGFKnD7L7R7rk9p2idIRNdEr27EqQ/h
LANaB3uHSaVlFJhwCD0wZ969kxRF1vQmLsO541WLXbU2uXwS4vAI8nIke1GoaN9d
locaSOEEC4j/jEUhqVnEnuOmt/iuk+t9wTHAJLGMYGcO9P9aoaCOsauAqkFpyGHt
baTRHpcWTaxyx1u8FWhp5gK3YoKu8tm3tcDLxRKpAcKljhhL7Nto7g0ckUftpg5R
FyHArPBYjz2WaEvRBxAOhQbnwfjVS5g4rxeYBDSgizH3fClYUVgIaKExDaGkag40
dAcjObZHkMBRqX3s2hOsIchyBgIcHJ5xe/jM5vZmfzK3f0YKtj6ifbsR+o3LvXDS
7wQwLjaQtLlmsUgWDwWLX8+fLzp2+tMxm0Fe34/sSg9y74aN0YpJNjnKJSxVUvCm
gg/DPopZ/VQY8klYHtKDTeIpQybadP5gUKEl7slFhkonQwEwkR+Os+IN4t6g1W/T
dU4gUNp0N2Nqa7jn1Y84oaRzcgPVgHOyyIMqcGuTB2HgOwls5k91AihlGHuxzlI1
q8iwhoI3UgYLqrageLm++c46EANXnEI04i0lDwIHqwtTyab+tWCiHKHVaDuZM46b
hXBuKnOGOwjGt/dTfWqtoGf1ByT/yk+h68wUlleqIFE8gB2H6Qvl/SQVdBQUF4RF
XWVLsUTZpy41jBEnPR97SibKM+OtwPhPBKvxBHN0ruFbNsPKru9DzrmdmMzwoRNf
KAhLDI4TFSlja/mLf/mYn7pujWDxzA1D7DNPMq9ccLTrAFhMSlX+L1J1OS9HtuPK
DPw7hj1MISxtLRYZSGHROBQuyHjcQ3Z2/faFV+Q0qIMOShMv6DxYO88rpT7uJHOl
1ezSePwclUveGma/rwKzFQvYI/82PLbgEjQG7FwZoIwJwOUn2prTvoqgFBFvNxzL
oxgT8HtqJ2vJMB9aOELPdkNkV0G0WvYPABaykXJZFqjklTw2O3mwYuTxvOZDm6HS
0Xzw4oUDaWo1fRvhyMOi+yWQjOejPhzjnHSfBb8ccpxx0k/LbYVZCnYfJhwulzb6
Tg7mWsZVToUV4hK5UeW+oredmPEHMhLBz9+nOOSln1hfZbRLNoAeLzpsgC+EirDk
gAJUuepyYrhYfGqcIPtkW6TI68Y6s6QScrnOhuLNgipOleJ7TP7P1PgdzQOS9bpj
Hg4yBoOVuepdeeOkDnguOtyGh0IVJJZSoYD5KE/qNtFQOBAMU0yOP0/GgITMdSDh
SUUJOTlHBcEs5Vd8yuuaxHep9vgi/7fsWdzrCAig1GkF4w5qmN4dzse24Ebus7wf
WWZpr1qwKIjYJRm5DAkzNcCtjndXhV4JFg/21tn7xk6b/xUaTGA2uNsPwQ37AV4/
xMPtsSsNeLpOgxQmtceTGzuO8wzRQwDd4fP8Bc/W5zaCflN+U4bUE0yVvn2hycD5
5jAbzz2KqHPcv85R9BTF7yVQVEbaF7t0UL78IrP7gDF8+fm82IVo93ubnkL3bPmo
9i/u+ellCyjDJJ9Rl0wzt/xGHbdlR71QGjIGLm3HPmNbVDVWMLAq75q2EVytM+5l
7MG21QIiEsSxy20usNpRG8cAukOTFe7h8cy4TccERH9SiF6Ib4mVswQKHLMHd+WX
nBzktW/ulFhA7ZmMKdLhbRjpRoRU7MJhVvneFph/ojzK8QfbzQs9yvy7v/JwwWFb
PgiH8zPW3EsJsZ30PWNxkeYf6UpWp9WQB+5VBrGhScm+Kn3631Ve5tzPHYCaL9QB
NgDcq1CHoVsdU3H5WdH7ONt3NB97r88n6NFao9pFaBi7LyJla+ZXh0VVzzQJbisH
NMeo07uu1B1CGchCtnGcajyGoxsktu5dVWZckYtnv16I5kawVgj/ZzQHnHl+IQMq
zC9HPiqubzx3vo0wIoggkxPLO7SU0r0g/D1fadrewphGUpjlh4Y+OWqVAhpNlFtS
BcE/eWSPY7oPTjqYD4ujAon21jsGN3tIh8Q0S+7z/UNu8VYTZNsEJrgoiV7KgXwT
C5o/LSe+c/7B11sE+EGUKosbHFJ/zzeHUaOU9Jqn/S0Yt1axdYdo8apd3CoS/hBp
TcfjXX6DQd9xFF4Witffb4l3NTOzLJF7iop0t0ROyE8UePAWtsTEZgnKFVRtJ6xk
sKMGEYVlEWQ14lKy7POix8gRNrL4QCQkuLNo1SGRmdz3gyTypt2nfCkMED9d0c/b
/GDBzBRHsEzuTrCdcqD7s5PlUf28H6cSSSc/Zg7m49r6ihmHqmy40y7s4n5fD1G5
kW9+x03Dwr/S+Ei1WRvCrD3u+h2xb4bd60IXoZzFGxy1gX9vzgLYgsoNR0eZzc8K
8V+P5IOvunF3idY5eBc26zVC4NjrC9am5lpmDdT9+gIPki6rGE1l1t49/PRu7ncg
TBE+eQbYnuIN24keHfp75efUzBHkGQF8VLLNkGZchNm8RwGYIcP/Q3EhAEZGW87q
nBl2pRWQvNoO6pRNHHS8ydmOnBXbonpUoKLM125wfwXHBii2aBqy0v3bVSrBE76u
TEIq7S46yZByhqk4R3jj83jgIgWjRVVQJTMNJV/Nqov/tg0yPfeQLcHGQboUrb+T
5cpTLr3hF6SCSdb9yI7FTTrE4E7Qn2OyPhSLk+s7G5npYXafY8R6lMSZ/ql19oQL
F+1NM9km1fd4zbGR45o5cmnjUj4Ragaw+mrgsvJ9MZwep3oSu2wcqOzTE58J/yX9
wBtOjJct62Sq83ApXOYYNbBZAyOby1k5diBw/0ugWQ+Ogif5Qr3FCDTwThvOm8U1
h2IIZrmlNurCyNmBwfd/zv5T+6Vpaki/5uB5WCnQoNw59HlsolnU/eWHWlYPNROe
4+q+zCWJd1NtesElpF5rHf2uxwVGBjpEDJ2aYQULJh7P4yJMgpk8ps2dmvoBOTRr
QJcqWiz0ZSAx3coirs3F0Aqo3vx+LIwpPQnhoFWnd5qWrT/zE94OhhQSuBS6/HLl
rROAirvcUseplhI49K13fBUBe23Ir2G1bOFFaeQyYLrYy7g2ejxfbHTt+o8kpCdk
Xc1TJelZ44I5hygCPMiuAEWzqQ5G/np19J/LQcGRS9niQ+BWAIEbgejs6IYpO3Kh
h5ZSj2graie0ZHReEQAqR5YCFcx3XAPrID9cw05lx9UZXjCdzcD/yi3mNrqlnrc2
+JB74D4cVLzvGaVvi799afN/p08caiH0nmTrxW4ijdOKo7TpHWluBNlbWwNK5dpq
/yhgwsKTknIbmpZudIXwZOdRZod2Brbyi7aXYeMTxRb8b1fkfCuVk+ksKOiQZHYz
DNm+BmYpFFbB8U2e0jyTthQQTZk8pLuL86Oj5kPlspH0dBdrByNHfYx1LQQKhVEA
Q/0Zd4JWvhXmPvdYBoxfMqYEV/TYxxONGMmmjEi0DRKjgzSqwNRIv4veC3cAEANu
DwSxE0TX0XVrSQLAviIFc6TKLdom1iIyiIkKq4TtC2y/rgov4ufaxrLY1kfjbotI
ASZDch26e0GsHOHU8RKd8qcFUwFKe3yi8BGTzdKbajrJxP8hhvNfFrPUDTfz6RxW
ln1EO6aoRMKfKenbcDdm9iT2/Y/47NU4NvN2/LMu/8OdEXUXSt4OI4P8FTdJ16S4
w5ZBopPvrZknCADQ4Lpun/ldA+HKMy7aLEeDdaY89x2ZT6A48U7ewSuryPnpESp6
4m1JKKzf3cR1EQ9f7+YhwE+u5OSQn+8l/xgFDDSQ7udk6lpaTstY9Ku8iVt/ZeLG
u00Gk5wQplQPMZeEmsY7UQerwGcc/0kmyUMnXSK2c4LP3idzEeDV/XnT9mUusYI6
XMLa+M0Jt3vTwavSFDaQ89PbBy3JyanG2yRyaGE4Sa+aIDsBpaBKlnupC9hmIGjw
c4IAzq0ahBMxUVPF42pSwuM+4NmjMDSeW/NxpPeC/5k93Be6fcZ6P47mPym5X34F
o9ecq7FH98OeHV7PS0rVYpaj9FoPwjRE2aa7CUKslxvP3XBXyhArvA21+0E+1yS6
AtcatRSOjCJY2Q4lVcvNUOcM9m3/mcaCiWNEyHzJ8f1NtIpyNzLOq0Sfe/0C27L9
4obWMGZIYq5hu76PSQFIRpzdsyOKo9cOZmdlgO7zuXM5z0eg5Om3aNWuRt80xgYI
7MeiSq59MDRg3b29QCbZuvONs27NguZdBNVwuK2hsN428qPdf5/meydz9nd+/npB
R76Hvg5YgWWF7cplTVGx8eAhpYZE16eb+u0oSg8h6Qk6XU2nWPgDHhiVfKkYj+7k
k9FeYpZ3yf32DIjm/LG2FPewogTfqQywYCBx3zoKB6rOb7DgM8aJ5R4DQ3yfJT4O
T3x0+FekwIkJi8xusO/yUdvNeVJh7Kz9lUeKiz6P3P4DWqWWMz+yh+Y2e8qapDMn
OIvIXmHSCWwv1wAmI7fmcEr3Pa565MQ7Ak9WVMuGPIYqpShQ2UqOKorX9MqQCVgY
FNOPIFijxW6vIyNrg4EV8wWqUmiYbfu1Acee2qnyPAO3pHemea5YxRweuwdlu1VF
o6OHn02R+82v2Hv2+2LPam58Jsl9LFonwKqCg6O/8YgjoDjl14mZts2cP45JLYVf
p4PR2P8nDFL76RjAmqWNyLcRr56y61cUzj31QLUKy7Pgq2BgszXJOG9792FfkTnc
gkkyXXs6fYvpL9D1Gn6WZt800MwglTUAnGkjV9zr2uZDmCM8A8Lsq2cC/TL+ETGW
enDoypE2nLPtlG12+QCsM1tQNLdOKFgAckPsoude66OOhQZj1Ba1U3+RTLyBcDqv
ZX8JUDKTjuz1dr+GfLLenMsA35UoomJwrSpOBA0z/0LBPbEQ9j4/Hm+y/TYDoTMl
CdIfcfZpPNGcczZZHr14RLSXetdND6/77oYE6ROujODHa4Lxe8fNk/AEACIMaiIF
gCvbYF6Z77G2YJ/lr0BS+2MdQEE33TGcRDw7TPbEGj/5Q9eUfHTG+kNvpr0l1n49
KV5v46qoEfgYYChqnDBVWkHJGL4uKqNLeye3s3+iBkQW9BlLQyZ/x5ozdxVbzXf6
gRjObC/rzximuLIvj5VeMlFgYz1t+JcUibonFM6tlg/uv/L9ZSEtonBcHviUAUme
3mCfe401/hgXlsw5qI/4JIaAp7slicLX10MtXzQ/qiTUxGOyZ1qYSGzn/QXpRWzU
U9qvf2FrqdiG50suNR984pM5iNji9zmsHSQIgI7Tq96FqHF+DPYO7KwQVMqXOUmq
lPSwqQW1h6urO/ArqgnNGVAqA+Pzij4GghyzgrbtpRUHuwYFudsCxV5R8yZ+rfIi
Ia0fqV3CbeydchasmiPquQXuxrTC1R2fPxUBv+HCfy9Q63mFZz/e1TDUCDYiAfXq
FOfYmWETxRJ8o2mFgMCop1OsHnxdplK8VDyAuL2TjyL7giJ5NB6oHVjhippC8AUZ
fXjmk5Td3wdhiDrizkUa/jM1l3Cih3rbAVjlI9TOwsKI+kMDZtQBK/7pno5nkBlm
MffkK2jGaGDmvkW0ZDK6qO/E97SwMOX4eh5Bi0HySirhjHCLAgXHDnCKrPQMZWDS
IuPe7cay9YPYG1anq2S8Ac9lu9hYyob3V1a23azn0B/LTOaAA/Jyj5mhBBNMoJ4Q
WtbaeHpqUs9vFBe3xam6us4QInuaRQsZ4lj4IzHZVtEm2vNrlMocluDTbHL+mqkP
zn1m9aVsZyAonRpE3c248IiU7c00aoe2I6E9oNx6nWg7z10d90EDUmSp14+D416y
v8yS47w1GY0Ibif15l2Vc9TmeUXzpOC3f4hYC9zcPoHHAdtEK25lespACPHD5ogr
0NrnR5pbM/tL9VF4amSWxbFuHSG3+w5UXDlVoJbY/MzYoICoQQbeSxqpu/GGVvRd
FGGfemXTu05PRNwkiRCIUU6R2JxXkIAIQPGuZY5bldMhoBnYZTT2u1iSBRnZ5+ur
EEBGTmSMNQIMajiyNVgj+jDwxc71bWUwGPkvdob87Q6sl+XStZidgfOdRzXtxH6B
cfSCMDDlAUf01+vN8c5br6542L5Z77kN2mv87+CLwq6llOMoxuVqPBb2niZ8Ltmb
sYbeO0PkjlG7LRBYA0nd8Gv/HW2BiGLSLdWHpE/HC68lQycCUTBIegvpcR+/joTJ
coLu+bpzte5IM7+J+M/ZQfWCoxCalfVRXIQuQ3JrqP3MiWE0v//T7OA6s03jNoiy
U71DwLUNZhL2jnyNPh5mQdTsxSzt5NjciTj/zSdH2W0ufehxzrPGWeAspPKHxgBa
KRTVCBWLk/6kuBBHGESWUlsK+4sfT1CjHiydPwWxKKJ7pAvW3ExB0yUnhZfSfGSp
Oc96ELYyC6BIlenCEUPANmP0LyBOhkJYwQyuc58nnFx7bS1VNkwCxPFp131EPS6H
h+xySk44g9KcQKMa5iK/sHMmJOajzgQkLiAc8aP3xxiLAIKoFbT7/2mD/BgYYYj/
b2gP74fJPdZKcvY4EV0SmYZ/SWaTGijpzUuKiQle/WO+e5IeUrgWkOMWjx1iitN/
43afz4GT5sTWhJj3fpm4Pe7cl93isOj4xkA1xpkMkrGVd+2dqheQStR3c2+034SX
V1l0RTYqN8NIkjljax2xiRO68IwbOV3M/P0XVXMKkjYQuXBL7MabSk61DQEBp66A
Ml1gvWS94nHdI92lP0OAxK5AWUUnm01WhGrui1AQyE4V3KVrxu5UydmvJKJJWyO2
3L2mB3236hdjReBMVMB5jMn8vzUbP2bPioNiieV1244vbe41xVw7EFi0ZyVg15hk
e70bbS+PtmpTAyS7v1ePvy5Z2NCmPxOfJW/WlKCBVdBBiN6AXJFWbdzGJSxbUnEu
PTQHO6fw/NcOyp/q74NEzrKLqRiU1/P8JbmtK3giKQLycGNLX0bDyEHfs81bV/jT
f28KgclZiiJXqZR/5k5fhBN5bd7cSf95fzYAJRkN0+GeXUsJ5mqrT1rmuT+Rcw8A
4hVXAjfwFo/YhyfBqBvvvuh/0xS1giK4m6uiIej3pZv3rAmzoVYgtN1qYmhPFT5q
vUA8Mb4C2wnlfr9f3k879D7jsjH0NglSW4bK3ZuK8c++PW/Y/X1Qz1hThdHamZ72
oE0mMaaPHKhuHcq9jJadBgPH0noPbIiIzh3YYetliToBEJoEryEjn3jsH+ZZbU9b
oJ6x3KSjLnCSzDfcLzeFPwGJczqD/amUGfHuLDYuLBN0mgy+zvHqeTZ2D242Z9RV
VgrPQr2o/dfG+ZpGpl7O+qoEcOjQV/mhUZv2HjVPCq1iDseegqaHm9w+VGd7M8Kl
JPC1lZZGeA6ytVMib5I9roWCUPfosga42nzDfDkcgHRDuiO+Kk5NJZJiIUxZEQJD
HELSueQofLL5rd98rkkSUquUy65cPo6R//WkCpz3LEOdYPQmAIEHGO/alc8IfjdK
lviCddtTXlu7o5Qc+55fjuvByad8tjyK9Clmy9QZeuqZAXw0And5TWiMTMyh9NcU
hMXsr/DbSd8Ppk/4WsLBe4NM79VzJHk5H2G4S3aiNzk/AuIAonB2a1DjEP68BEDs
dmEj4692Xj7Q2baC7IzyzfLTX/BJJ22tktiiYSOBp2uAv7CPWbyGrozNzZTfvELg
7loOm5EtKFQU2ZXxZyZEbcq18xCiv5PKoeS3dA4zAfzSHpLLn8l4IczmUx6AJmgw
Xk1IaZTrKLMPq4B8jr+bx4KRQYviIIu1whQWH15qj58LVM2ssgkFgTd0AyO3qEN/
r2HNIDRBpnUYGaKu+HfnOONs6EYNZXQ9FDslagb6vMr7LLVfRBAdNzdt3xTeVANT
BHXJ/s+TjLRD+MibLrVuVh+y42dhMIohssCN2+OXl0yzc3kGAveJhaUrkXqQ6+Su
Ch9Gq1UpEsVwP50CdDx3etJJ9tJhEi9BNOuQwY4n/91MoqUEj8mCyul8RB9RWLtt
YzFWwGvkdRoILdYrcL4FE+nis35wCz/D1pwwwsvkQpGf3QopnYaNkVKwksCl2RKr
cCASQ7lagIjueTP9toWsqcKy/M76BdC4muKrfosLYA7QLD+ymj+bvFUwIsxT2qpL
W0YfZ91zqd1mJqpOACeqanAF9f2ppRbIa9V7mdC4jcS1exuVEl+J7TEgHMqukhJV
P0zK9w39mzGlFv3cO3UB4jhMQkxWVBk/yKXiMuy2yHXBxrvE8rWXUTVH0FZE1USk
PXA8muhhFbHL1MjHh63TR8pZK1Hy14KnhfodhYMrc1+VgJ0HB1ir4YWIUnT7xuQz
IIcEUnfnTKcDYLMwRFarwAvHLpBTwOSdndPprm5WlLAeFubVzjaevyGTONxn8I4p
483yL9R5O0jSZIKBWpDZMT9HqElXmyO8tT82LHJKF51db51jwLV4cEvmqIMl8GZQ
3MryL+J+tGgUi9DxHHyu6ZNNmo8xMGP0nIhr2tHp1xgKBit3U6zYmjxBGyBdeVhN
5MmoFIrN34beAx3PK/nMFeEuTnNjyUbjjdyWOztA4eA32lQcP2lifWQ1DKLyJlsY
xgz1moH6YR/SYE2Swu08hhUFhel3t7FM62Ht6/npFHhzkpPiHiHcg9/foG3wpayG
yhCpjCqgctB1qbsm+CciDDBhbPX45jr1jfey0AlNAwPIqi9rP8U2/wbgbjOZBnXy
Suhp9qc9tdHkeXSv/CeuFCSca77rFSoIPLn6PYaArB3cZt3T3I2vbkblYVGbfrBY
74vuDqgT81rvI+P6st37yAeagERKTs/Pv9ceNeMunpREi1I9tBU4F3ce/s/PIW58
HtLanF9caCZfvSNAFoLTJM4vF5TtIaaA117iVEhX+JwnqWL0eTRv7O+zNV8J55B0
jZLG+jbAsa7N1Vv9a+cCnM0eIgJS8opwPTDsuZdCKDzLtXgc+EFKievySWXQuSkZ
QEsqCSV4Q7weV1729W07uscPJqeFSp4psp0sFvDeYKYPdG8eI91wTT1N0Nz6ycFH
Q0PIw1lLRl6z3gJkeWS8yZhOljDTJUWwOgM4Pa22pMgMyTJ3R01VkdW31SbI8kLq
387nGKiK9esF3NR7xi56pHSgRnoRpANWPIZqWQ88Pv77nhj9/X0E19EV8LcBJj3L
rpFvbVXJtZs1MN0yYlpUOrM22LnZW0Tl0iObYVzQCk80X5b8u+qAw/LqdLyxg2rq
psEnNyanz+PQWyZo4sG2jNBbB3DXw/wj0y9SnpGyjs0dlXmqwLDayoiWjnghcsQs
eMgz4XkcXxVHeBzTS0omN20jbBrHgpLGVdMR9V6uzO/qggmDdXHqaqWDTmJPPCUJ
inj0HnbDQtgLgdcwyjAFQm5BeuNEApHIFJ8LBOBT5lbcKBAGxxAJyqXyjWq+COac
/XN4KRX+Cn4I7+qVqCwOltl6bVS61ZMVKWTVTgZgHm3yMe+q1CheVc3IFP/uFHYD
LD9W6L05PBCg/5iPCUp2OGmYJ13NDPzHC/+E3pUgBKNsARexgjKhmoI85qdMEkca
xSZ+5gZmY/pC5Pf3h0z61uyILJxYnR6dPIcBEiTJa43v9qJ8spdXD3QhDqjkS+uf
8g98dKHcykbQsiZ9PTmYdEG+3Bqgu8yH2tkEMgBqhDezi7wzDRTJmPOBhVJb2boI
k5triyiAhBdhiIeZoWzkUr4yr6owf6kDcSNxlTQGNDohNAOX52aWs8ssWOKQNg3B
tW6blDtlKsyPxn2hSM9/V6dpNXhq8p2euy6rcsCccgcVcHVVwff+yKHSdA4nw49P
br0UN/jW8rbPzJqChHvDopYZYjqcXrBeF67ye1hDReegXhm5iKC868vMMPRJsPjI
yFMAe35ldKNrxS/cabG6oHRP8H+tOxzMBCH0zbeVAoHXpF9OT/6tETymP7j1r+9f
9EDKyOhh6eYWMxH23XqpSyYEwYFGI0/uMtnFEkRYvE2WvfLPILav+V+6rIkIvHAu
x7/4LPO2uJnHLwhM5jHT/Hq2K/bjcUIpKOdRcIWPx0Aq+Z+io04KWV63RLuh4kI8
IsHnaRCBRJ6u810r9tw21f9xeLB5qTaFaChjsPnxINhmAea8rTp1/Py9s3E8xrJw
ozS8cwu4dfAEr610tAX8Ygxpkm03wQ8tC8oDY+gnWLhX4xbf4zN1C1hFalpedpBr
KJAG8r11v07/jPb6VaMQ9gHQYEV4MzI1D5WEbqGWjo73R6L4lfjSJ8lWBWCvuttp
Z8xalYg8H5UbzTVjowcn+w7zJlqgsWSDG5CX6Plv2fABw3QHpsGROH9PbZcUcj5b
NdlmGHR5hfyvix8fAtgCNen3mgfdXw7v51lkoJw2LeQeK5tSIqAvSZwTKEQROisD
Mb7y3fA9r2e4Ba5rKdZ6TVGnBJJ2LQfynKlb34oA+AuMoLjJrwizdNPS5w1u9tM8
L7rkJ0qfMRQVIiY+N2szDNPWnXqz3mnmJMbjml9EgvEed4zisJgSENNGb3BC1BW3
05KPoll3SEa4HkGnl1RcgkgJ/WLWTaRa7S8cene/h1ghTMd6wj1KYAdwbX8qxkWm
J5vIgVsnBj+5yC1S6+iSdMuzhC49fKaWEZevWyOWDz8bU8fosUsOQ8iBu2nLjUpW
ntjPm6rQ3nM0BnxZDuEd9404przCS1ot4uQYaNPQN2r++iJYXgyJOH6W96yYEx7p
Vc/6+yA0K2ouBVSdZ9ZDagwkCz6Nm8Zt8G/Efwvaco9nGTANLXm5cROiWB5XRhzq
cVgFMsp7WkWhlKXktsUt1lFcYXNimg+aLDCiO7GRatsqdSCl3/4Z64PbRP90cO5z
i7M2HTRWMhX1W9bQ3LJiY5gJsq0cGClLzLAxDVtOuqJrU2H2Quhm6yme/dPOjg/v
+KmXmF+dXVEb6UA4aLzwyvPD5ql2ZyXZPQy9zPX+tUt+az8stx7LfHSoOrbh/HRx
3wtCY4wrR2e65UyWoiQDSWNuHh6y90k1hw+DFInjebBnmqPenOFJseL2WllUtWNj
kbWFS4lQIiu+loD48hGu0SkYEXy3phkXLWhjgyjHFkspvTBlehmFmBBSzgMubYRe
eVRTkBhDU1ZHknocwXeZUriPBIeuwPengZKb9bsD41y5bMWLD1hyhjgu33cKbMjx
TOZG6XEzpWjBXVL+vT1OaS6As21/cXcg5V0WF37RJWifW/tniQeN+qb7gayYrApz
XFDc/zu8/fY6y+q1dnkntDzgGJ8wap33xNixALkIO4dE5nRhxFeAJwF/XiKplcY3
+LPA+Sm74g9tsv/lBObIa3yg9u7Z8oY/pnU+srL31Mko9ay0aMXoqX9hjgsFRWJR
/MUR7PQ1bMZ8rwUAmOjFnOT8jJ91syvb9tvwhZT5JgG/cjIBEGoyaIMhWVHq86ct
gnqAo1tmdqqHzcflmji1f2lKlip3vnVoZLvFiZpAQbIwdBT4IE+ae3uZ+OnWfwRk
YSDQrzLO1NKvoseex1jf0hu33Ny6t/TBl2/NBNiBCgUpOB0OP/heSUXE64gcrvCn
CmpSQOKJs9tl8ESvIly3skVMkEvJVpd0kt+mxnLwjyJQsiWPh/ZV9F456TR+kPRE
5b+UoTs6YxYHQ9gy/HHNePY/HCobPLjcHmrmtt/Pk5v9OClTcFvB9+NqcMB0aPpQ
P9858qZJrmsP0Qx6W1AvLyXW8YKGXPoGTWCXOwDgB2/O/aNHiNzYaX/hssS5uE9d
BRCr8IDD6A4XgpB32FLvluZ0h9QwlDb2uUtNGH8dSCoU9AwTyhsrFb7Yb7FxhuOm
tahY1fla5VMglJK09tbT+F64lDUSF8mRFU8mC9ygh5I+AZ7bqi3zUcuF0BdWujjX
Jfax7JfWIuNTAZdS1Sd/XAJ2JBP3fHBbMUYU3GeVbnGat0yR+lJCVAdpcl9li826
2eZiA80h1JDycaKK8Yn7Ro4fGqfgjgnVsuCh1N6c7YzA7EVUlil5XcTkvZLJBSGS
81471HaClFaT97OA2KmffTXCfsyxXHMs3QGrxA4cVwt8BlRCDhk0AJO5xR0AQPCi
v8doZ34wyO6dcUr0cWjBhRIhse/cxpyDj93OJp8rPfsFidPw3boNNfN6DdGInwUX
uXs0dAV4MjBKwXt2MOPlcl6F+HexO81DAjmo/G2yY0klNE86MISuUGmlqf86wsV0
6JX8MOC4zrxISI3fWhGhCIGy961rYgZ5NxXXMEH6wrXjwvdZYnzpMWhKXsM4lApF
JEzadg2EnJ52m52FA071CqbFnWamGnHeqsICxVqchydT+o60UeJJqOXIhgUZ20jd
b0xaKbPzZo/imPzquayACTybhK3YTZuOtUklDxmt2wi5FG+927uFWF5rJcizopyY
QIdMfois2KgtQdakMoGEeZtMQdduUbGvHEHYfn8N92EyyAaRFyZBz+DxHcM8i6Re
mdw1CASnIAkdG9LEH61CrUiAGP09L38YoMZgimvVnFV8SNlCMxP64UQ+vWomvZeU
qAyUuqmv7SVtFbhV82zrabrsJkQsXtlu51JQR7yJR9z7gNX4/Smw7vhnkNz+VqkR
GoZJ89kaGxpAc+hHp6Wu5J02P5r/3fhyvvkoIYaBu9v1UXUed6U6f1fZHK+Jm/fy
JktOsixvxqkO6pYh7pkJxzpRKpQ3vtoWSXEeMc7yM2Kg4TIw7NFCZXQ42bdovc31
AjX3qHZgO1ztmVlghhawOhcIZZUqSjIoow9HNj77w5sdgKjBc0/xZQyscPK7CG7S
prKDoR3dNRk4zjnaZ0ZhP/5LyaeB/TSRs279N8rAsKMc3WKxBQ5eelUYceArvlSB
FB0wAQ8qqTH8W17PeJmcTnBtNJwmG20q8oGC6cFgQ71JcA/QRxUFHn8OUno/5Vkm
yKCHoFsLMbs1zOn2lYQNrL3vC86hpr41kQOTeZxmBKpnYixKzII5tf7WdNDx7tON
5lktYAYwxBEUYWlzTMI9cFjXEoRzQBCITsLF6aMlB2eo+2RHTMoyyDCKMiftwzYY
YONb7sk5cP0mVszwdnsVKuUUvgmWS0hGrDqsEwUjhPP7I/zmJuvemfvoul9je/HU
8ZjJSKA7C6oQ42UqpmMox3yuLKwLcUJRgURUrOCjJdmphWAL02IlED8aKgEJxU/z
a84+BUl1bY11/u1ZvkmQZzhLe/yToXcYwdmBrx1fesgeqJ06GQeFRIjZBa739T96
IdXCbKC1ziUlRhdbdRs1SX3JVPbkKcuVrIG0ChGpFixFtCDAT70LM2N0jyVM/dO6
h5G1QxkVe/LgwzEYH2pPlSTXrJ34hNo0F68vmAvJsSv3M9hVX6kg6kyVNzPK4RqX
HjOWmDAYkzTUvuRRXSnzYtIq+zWj18vfqSUIUunyHjXenPtH6yqB0UsBV6Wzl9Gs
Oqm5hrKexDsUESTRTvVfCiXrZtYeQVmNlXAz+BKrTRUc8KXjuLY+QmqBbl6Ho9KY
fuywnrKsnGyjsG8/eVZKXun7jiJuZuFkil6TwV7XWfj+Ujnz46c/2EOowmE1nVtG
/tjrWpFrT8UU0q9ri5ZvOM63Q1NgYRH60Ny8LSF50pfSUgjnlu1ZgCWKDtDgXf2F
oAquCyn561R44P4vA/hHKvpE1YRqibk5MTd5YxIgtJc0u1rF1l0QA82g5x8u4ZXX
wEnxtZKYxU1Nu6iKi8B2t/4dufNTtyc/XSVY8Rer+dPtPMsStzHbPJ651n6Xv9Wt
j0EgJolKY/CzQcPqDnBQm7DEXQOUzlOWBSMe0eIe2JKAfYL54dYwGp6bwjDaBA37
H0Q+OlTICM9Tts34d0DiV1ebYLfs8I3JsXTOEspExtxRSE2zGZp5ViHffCD/Qw49
AXm1XMVYF3Yhj2nSI1o4uCjr2QzqNQsbfAI0Vt1KUlKb+x47lbVL081lAwZSMRp8
+MC4SY0hfjTpWopEiGKcfK1yhOrl6UYDuiiTkepjB48Qwolj10mHBcFwaQgdyoCJ
AoZvIvu4b3cAC3teS3VZ3i0NGuXzdhHVz1e54Bep4a2o+6zAYf28YduOTwxkArMS
PJSza4vZe4kytavlE8j/S28CVkAJfYu+FoWxd9e3RREYkWkPP2pL8X8Es82KE6Nl
oAnDCyUzGuh91tSShM34/KHgK59lxRWVHHxKGdmw+zljVFGuzsr2Ms+aCGTjyDu+
iYDRk//qnWc7Nm8P2aMsZiQNopk/PVVdcrL/VJQrA+dqt5xM46NZNzi5DaAt9pma
iBvk9i8Fd0XTLaK7s2sMFS0FBy9DrFtH0OGG2RK+halnPAuqbNHpUsQo4uNNqOVj
l6eRNDsnujl6M6dxJi6lWQsOHDMprh9AoTiO+OAOAd3XOOdH3F3BMxGo1EKPCZK3
2uhtCUCEnau32Wu0IU4kg3ate2tyGanF8o9N8yiTvUprVkYQW/XJMKH3fB1G3aml
vcI3MQVnH4OZ5Cxs2UL23laIZs2NvOYvVZYHwcXnMBZn0GzZ/WZe+K7HDpLDxXsf
iXTvOOUVqD1FDVqhSRKAExuyTODOwL2dyjAOZmB/5+PE00Ofuq/BlhIn2u59USHA
GuyTznuLhU8BM6rGKQTKs3AMrV/7ReDVt2b4/Ci/a05aAR1qBhqLLph95dlD9QvO
mkJ1MThnDlfWSQh83Xn2EnVF0gYF61ucGyJe7wiVxNRTe60Mj/JvPi7ol/dtemuK
W8ltzyFpsw9/4I3iYUMzpQSJ1n/kpIND3UGR9xIg+VkSKz4fu3XFXCWM9CxKcQrJ
cKKa5LOqYZPMTBm+7dr97FK6zf5dzAB/i+ToGTogA5fI5xQbA24Snnb5UIVmgfRM
YEgwqmtDOYPo2dZ52fF+xqB7J3ajlnNuQKeiZZ8zre3N4GMgS3IpQGCN/Ze9eWWH
lqJliVI40XL0bBIvmu/WgPKN7plOp5NZ7GvsslK3CkKjdR+OsJgAJMHzZmghuFn/
JMbzPNnmyt/IvJrKl1EHAhQB6InErj7vFZSC3WuntuDtHHbMeTcBSm54phTh02a7
UWzODF2BOFL1A1vDMqeTVkJ55N6NH9rQs3IB7zJghbPROn9Mht+pqmU/a1TsBlf2
RYiX7KhIFj33KZs4nEXrq/UfLeRiuCdG+f0gzqdUSYP1DnoKKvRPrrVu7CpeO+Qh
If1chSKRf47+c/fE9HfBBPv5jd895K8hQMLAlrVJuB7WsfV6kY5UOQyH16XrEN75
0YTqv5LsM1VWod9dNngo5xV2rZb7bnoWiE84vCQ90ETZLIO2zfL8HVSSeS9aAWYs
hnhtwkqJA1GiDpGSW1RKFveP5Q0RidKy2HoyCebxxPlmGx6nklkp0m3VWmaR9mbD
MmeGxU48HhqmfEnETZv+ffMtfBw85uKZT4pccPX8dtOQg7OjawFJxdpP+5drqJPk
cZX6zFnVCjOfVJqqYfi7hi1jc7DBQ/PH7kuxkXgJbHokQUFyd9dXCPS6K0Xoz092
j/SVecVLVSkRVXmWF769od71TqsBCF0jj3uTQVTJqUgduAjt/coP8ille8JkAriz
bwpYLQyDRS3AiHQwPqgsRuc1oWgHcTWIKttqrI6fmo9GUtLktYxBzl6JpLdbkXNU
xu3YGyGuJf2ejsySccDIJ+EO1mW3q1bWv/xgIEwHSza57VPD4/jf9HoqxSCxtuRA
PqJk0c0qnQbgwi4k8JHVSLtCETvy6MO/aUq7XWwx/2IxwJeY8fVd7WMvkyCjx4Zz
BMN1v0mimEbwiIkMSpugiGoTHvajYXtoIDYfXGDFJcAbHskGZmXC6HsJSy9CEqYf
/C5uhwMWnyzAyHJycng+Ti3XNXhopxTHH9MVjvIhIviwyT1EXsyt2kww6KlqWYwk
HDkMRcFBd8AWcCwV3kl9HC4FfMudqZOL8cymEFRqz+VxlfYLEGeHGsMxaYXzZ7to
2woQx41W900HbKHhVzg7/+m4zPlzZg7nhhzgHv+IsfUWmKYBiGuQN35OtbksbT0F
K79t+KFH9VGIbU4ui4vKOQmPcbmkFRGgdU6bKemFU4KSQJU94hvh2uUkOTm/4zLN
Sic9wCeKcScUw2dtyWj6X4FG7Ia2KLbs264/LN9gRM989Br/AevZ2GoIzgOwVpCl
y2mn3vmnQVmiWrcZmoH/rHU6phW6CwmZZKh+65oiU7/d5UtwOWsFvlA7c8lF17+2
LijS6ehZrtFqHj6sZKDwLOMh6prcyArTa/h/wtewwu6e0psXs+hB9Gkuxm8re4o4
C3Jtuxv7I2AMxvtpZlGnkTUwsZyDT9YgaGARGHIDxjRQT8MQN5N3B8XMxUGvDNZ2
HgXlosC4Mpy5eVWnAqGY4Hivkav+YxPaiTPTkx4EJp/doNJ+lrEFlWGzq1EMvcIV
ql1Gr6BWWwBbbitjzZoK3CSWvocsRXBrGcul9G48urMN+WuUYJZrb06ienQurRlA
wyTQYjl41CXObZxt5ghoKJONwHb/MYr+nxH6lgAugWdGQDprguSVJgRUFf+ItquP
QtydNh9fhGTPdvZM/c7PBLC2YgAsSO7gTX4cbn7DmWsyTokPXIVN/bQMgbjqOaLP
2iv2rXeJJKOD/88xvYPGiXhp6Lk5ytlpOQL4Z1wazsU+RcQEA3+SSFrnv30MfgqA
SWNd6Cdht0LsNke3uMC+XhJ9a3aRtqXGkX8rsJ6O8MZbsP0/IFzIBY/W3lD7YjH6
do49zJBuXT34uTC241rwL3CXIEXQSKP+bCFXXDqAT4KrhlcwmH1RPJ0YYpAIoO+j
G6FQqqBL0n3lXlS0woHzjpSHQfMLfKNhNWbOrOmgR4V5O8g0yh/T+8QeRsYXsWib
8hJEKERC+lSs3XnMPWkPZrfvJKd34i8uv1WL+xvGiPbscU+YzBcflIVWL8Ylj+y3
hdVSa3IjuObHvjGoyxuDSubTCiL+9xz/ldAJH4jR1PtcvwNm0VAeBfyXsz4JUoJd
NDDdtlfngm7AXYr+L8OKjO3jwzPyh54+mtjAiNGcwNleG6OOPuQd8DWBXj1As/oF
pgnl2AVmm4LBsirzMkf+G5yDhsjIx5JzmVaFGQVPRFo9BNbxsVgcr2IL4gtgIAM2
iSGVLnO4P/fe8Wbp7+MkUg2FFefYoNkshii7ep31fMFINksBrXWgRDrzX7y8gg/C
nuD7HuLvpTxuQ/EC2BEAKlkIfGSLXkoe8swcu3gGDlNrJ3CLb6mkKqAYbb9RSMsZ
0YcgU+DuF1Z4W1GpV29pn1rt7vaWRkqpdL7viB0c6N8OYvewPDOhmTNAqe+P1RhC
oRJS1BVYA8TxrQwnhCdf/oAgI0xv3ecYTpT0sQqglOEyvGc7yB2qM8JeK2FKwRTE
Z+1jTAHBwjJJKUp7FypI6Kh+tONJW0nJBNl04fCrDrH3yrKo0NCdX1xcvEKMaHzJ
3Leqv3pQSsVXso4llu6sstg1s1y5sEIwKcvaTlK3fekmORqbS9V/qOh8D8PvFp3q
fxBlVmhXHfPNlUUhMxvGKpME41X3utkOc50qSyw4+5ydplKPQRMr5mPvDhwUVblh
/VmVpw/gNoGaG+fUfNqLYo+1DrlqkHmhinY7h4XiM59owbtP68yCn3jeILU/QhoX
hCPoY6p3qmiCuishliinINKsQbtFdziqp+ytjUHBRvKjGvweAZ8zX7vQOL0nwtE+
BmAYs8et7tm5DHI9q8djEHXmTnMVRXtJ5UmQPqVf+M8Yn39La4BpFRRWKU/oNiSA
MERL4W3K699G03y0yqW7vTXcc1kU0r8zNCAQ/yU2jJhqw4CCyx2ZyF6HCTUWk7OE
K5U6mbTlWnZD5Ml3ZBBZos2wAkZGbuRQFmS3NVEfjwwW0JPlvYXMNih6Nkqk/KZt
arxV/Bam/t1wY1VjuTMDpxaxl1MJ1BMgCjcyNpIpN7HO25urwqDAQ97yiVbXpaF0
w9olv10n+kpJuqHIoy/Ejt416GrpxWReUjVNUZmx2xpOIEjcZH1rmU+xD8zSZUgX
QenwK3aT/epet9fNiNIXIua2PAip+mRG29QDgaTQk0sScZo0XG9aZp9nEc5/Bg8S
cFtGL2xvvLkZt3H9P6D7o0rAWyqTjN3fqM3aGdS8Ry91/+VJ20ZBhDpIn55IPubC
i2My0OIXPHASGr4h2BpbTwIm4/LyTO9bl2pZUyI9POMTd505dmxyHNzSmRCeX6tx
/NzMt5azvdM6V2yjYFsNV7V8w/qfW8aXYSsBUL15YPhq7lXi3+OUIsnsMSLzNTY2
Mwh7Blrzyib3jXhIdKjBfihjvY9tq5gZdj4bbvkBhVeVZk5qnezVGYkvlZ5GJw0U
mwBs6cTbbHXVU8Z3emdYHAkB1VaegjPu6u6PcvVp1vsvSG4jPnVU+dMal8c0FoYS
gaO2LQId5VkOt/sJYoizVtQ3tOIK1QuIGLkkzFoasyC9PAj93aPgTPaN4K7xZU+L
3ogMgBrzT8iX80ETLfU4aJ43jX9/7IorpbXwcJ2yR2XlU/zFGWSUhW7jLcqnmoWB
dV11gFb3kYxE1bcbqADBcenvHwc2MMxgO3MDyVGTTMc4wyrspYiUrhYZh2acN50t
bFQmUnbl5YYFvhz+XxBmTpi3pVDbbVubZh0xUGWzP/g3PYoSPPfALWdzl3MB/uN5
nVZBWnbkkdzu1+n0CGljC1lVzqFkIgq1n3Ddb+Gxpoj4SpbFCLX84JwR5ktyMumJ
0RzSPvmmT2/y7fTpOM2eHEqimwTkCTH9HBSUc0U0aMFcMlLyqpaY26H6sdgxbvTH
JUc92cxzzczcie86slOFBpnYr1WIoAUAzWFb2ODWFllPsROaZY7JxSgBV4IxsN9F
BhOqNgWTEEqRPVPk3qS7ftAiYRikjyhs7CEZ8a22FzABBRGnFua34oUL0QKqhzPn
SYkNYtKvLl7/FSzCvrxjpU1Cwxs5fiDM4qKTW980iejzWVpReY9zsfaZJ1LO1GZx
4UVs6bqyivt6+C55pooR6IwhcUEanGrgKMExZ9UEn6155pZyn+bMVdwjM2tgIbKj
O1a7eX4RPuHZRib/lNnam5fJXLSEHfTcUf9fA2dtrq7T3hj1ge/Lf+CWqJ7Dm8q9
Et4soqkSpB2oTOMr1bO0D/riy4TR0ywZ2gVWYZE1am0+aSBszvbJsgzgTTxInw1G
bazuUhnBY68HcNJ8f+o0CsWq9XVB7VhwVar6ig+yzFaWRRmbx3CUo12tEsIlHNq/
JFEbN58ItMzaIKgwuxcjLu9sobYM5Or6La/Uynho3cEJtmLOKvMdxBLvlyat65xO
PRa3dxVm47Dib4T5aTDXUv2tbcqbiZLUBZQSwMhhYiyP2wHbbL6XsIXC24zx9vce
1s1e6QIvq8YA/CgeW8BRFRBIb7xw521wsNPMxa0+ywUdvnXafROWc/MVR5RSP9Ho
6oBD7qFy0+iB/LhHZzyeJSfe3apUlRG7yGIxaT93s4uYFxaykPZTL5hqgDaZYW0H
lcGfBvfFoNsF49i00WD7W/ICGc8q2WGcxljH78SuZFxsFUn9TFbkmTlqqFodNC6r
3bVsibrV6nzNsOm8ZuJFcOM3Lv8t83prqIBp6Wz/8Lcg9GBKjdpwGNzTvgpMw5VC
LtJ3yISJPa0OnqZJFnqBArj2VKPRGbbi9fkxVDc0EsU052ON+a5tQdnyZ3bNy3th
d023dmJzrRfaPJhtQv0XRG3jyReyx8dG4FtYIex4lxoAeFXVJjeG4FgU39mAnryh
9HrDenraj9Utp38CxTYURvyo26YNuvV+l4EtG+Spb+1U17ZvMPVBvDJWNAI5brYi
/fT3Ax0sFMaqPsscFZ1DiPGwZD7GmuIdU30CJI0zBTxzD4w92TvFzG+wRcqjY+6o
uF0vUhwCacxhRqSgewL6lQ8BCwLZXUFvyG5oSdpLcTV95d5YI0a7QrH7AXU5Cyml
RA2YFO4vMvsJpon6tqB8xO2Ap9fJB7H/+IItK0vjRfnW8fo5eOmS9cX3eMgtuvQ/
E4mUWZ/QRkYQF7DV+9XNE7DT+f+a/8TLa19CTlvQxtF7PBSvX17vLBz1MHu7p+1j
uMbjAXfO0iug5EuIW62aESypVbVOXQh7kt7MJB/PTy+xVaSRmlNUdb+Qtfnk7ZVE
Ggm+zv3iJeuSjk9YrQqHa1otLT+u2OjxZFE3ZrUTbDo8WH75jEc7gwMMYiRqxCFf
3ueu/Is08CNaYMOHAKAO0P/+wa2Vn2n7/c+FkUWPszZFnOnUOWqI2F5tnAFq5CwV
wvNviyQYbly9DwCxcOt/u1ApPAd25wbNptshPq63W+TOECKHlKMGC9PfPxRqf35r
DDHuosUHSNhjATrdpcsybUGIljswnfWY2QopgMod2PGkuDt3PJQIpBuKMtiC3gfv
+hZQsmS5+Zz2/fQ3HqkkcFbTxH+GEKzcQ7rDTltOBDl4l4rdqD+RMZ8S/RLaZFEG
aIOkr7icytmBIZN6w4sOGyPBboX/t7C0/kRq1kG07EjYNs/4wh5WMI4oQNlA+4Nj
4SJubj4nx9c1urr8S1VKE8sbm06tWtHVP0Wf/301aVTHNCPf9dlWzIWPEObJqpsw
JsMJ8zc0eDPlC8gitPB/4UlOJuw+GJT5ZTIwnoDv8tlbS5pEMxo/wBRw5Snbo1qi
FNI6lJJwLnGc6+jqBMEQ3hoL7GLAQvhzVPtgYkEJi0FidNDx7la/SoJCKkLyQyI7
MokXH2IXL4ilDe3GTURvj5YrC9WNLcYmm+yv6XISAe6l5E+70JnACUdH75gRvSYQ
N/t2O7kR31XgXyyo7gIPs4VRyexB737xuMza7jbV+pXNWCa9U02czS9pIf80NafI
XHm8MGcHHv71TBiZ7dxGKlw/KFWSsCYPhrAjo0mgJyIEjwYU/5q+yTSUN1QmoigP
NDXtnlf06HM8cjThwXoJt9TyUYnhCEf5NEuht1T0GxykwJxl87lIOuSxI3+E497g
RWYJ+fozQ0PKUPMVGAKWc6+Dj7dhWW1aFEJH9fuLNvuUuToOV7IlV4mGwNp+gnzZ
4VsyVaFvbq6gibhBaC/QgqtZ5cPS7eptjfiIimAsAlwcZA4CxN9ggG1Ah8vpsLqG
3SLy/55Jezvmo4wPhysSBPAoLBnG5X1KStSBD4AcL/geoZAHGQ0lTeSbUc8xe+TS
+EPI90WRxFKLC5Hl0D20LrP7TNyhGYNgU3+G8H5lbb6w4JHYe4WH87kVK5mWzRZg
ZX4HXFTOBkZX6Lt4LUdXvADMX97A7Wqlxnw9aKy6ZCooGEOAxGcEDHYp2Ew9MK/G
qmb+KHeY1R7dyScz+NhzIWK3iPLNrQd3mwChh/7Tav8rfjQqTcS+IW0sTOV1bC2H
AlWPhpqlktCy5VWmiIG7YQdf+HULQYWWshuAUUe5wcyQuBhIUM/sPXpyHND7D3kK
P3OlTim+hxGT8Oink9WVF+uIMASv+LDMOEeQsUhTugx8yVoLkF4ndBHa2Cynjxzd
dNYuBhPFDIK5vMsk1GPcXcORjJj9HdRmku9ZnbsQyFDvpepkIDJrZRtMDxflcDzt
E8ZvAYtDqvNyvGhKqKvp5frbGjPYxFr/8iGXDTBRDDM74mivNp01BNcYzL8Zwo4T
ktanTBoxqfiwRfPPTv5BOwoTsmeEhx8+71+GtPZvg7g12TyYfceCP6ngSMdTa8i7
KSjcPGO2ghSWV/cLI7mms9rVEZuKvrQogDqKRedq5vPZx4XCFUN2NpsnOMsmMRfj
k0hNCxHzxJ4Cj683JET+GqzWeawO1Vpw8q9aJ9CwCIVvrI0D1/8dMNeX5mpjTB++
HLYC/6wEm7/dJvUWxrHOPiG+iTwawFiaE2Ot3U/4i82NbvRmpCTTWvXz8MANpX+U
0EdkdEspk9U/ESmMpQao0XrVjsPKpdpMgKAnY0FKOufRi3LilZadB9WUGNr/zkPI
NZCqAtFgBbh+sVMa90ZsvGsw40QlgH++PgHmOv/ehfoOCGIOgPM9VwzIX4bJzLMs
UpUoAzIXid1E4Z9BNVqlZAqmsK3wAy9qQLVl9Oc3FozzJs+JcsGgGVtRl8ePpa2z
YBWcu2x04hGQ4SVUSn4JvY5/ep5PvdmsNkFZPmmVAjhKQZ8bDxr38YQTWTJ75u8z
U4ACuf1ZPF82y/ORd/AAmYbxo5Q7wMhKQj2kb5fJ9zXFjUdBSDcZ1j/79QNfJ9ww
7GIQz2V8EOJoxJiWYJCWZ7TtRysqtahnlqro5Tz4pkN2H07UHXeHtZpnmEzugw6f
0fgk4DHIE8TNYITtlk6xB96DB7+M8pMpZ9N3Ho4WP3WfR2Vi1Q60QK/GSzLUu5dd
J7dtsQCbpO9WzgeZwVroOigsXdsNCNaOnPtaB/py+ktl3QwhZMsP8gierB0NQc/s
yPN5iN/DlTrU0ZgxS2DAMj/OdoQO0dAEhAE9phHUHh1y32Z6CiWag54LRsx/zWp+
4c4f3hbxAXSglNvfE1IKA+MALSgpOYDZzGSee9wTsAZZSqEI7IViK011Z+Zchygk
Xgr8uPBTwL0aiOLvG24GEF8rQ/zeZtA+XqqCxYXgO4MILghgxDLW4neH5xekT7sa
X4q2jD+QxuN0dMzc91cDkgM9Q/3ac/kr9T1bhI3hHH2XM8n33QKsOhnz0brsa8ZC
SaFGu9A4hD3/RQzLFRY7Nzc8I4Br6zKDMYlD3I1BXQHZ7DdCXmFD9GplsWP+3lJY
j1c5PaZg7o1LguNuDbCCs4qWHgq+fJ5whFr2dqxWXbs7ktxulzH1tX1KINNrasE4
/sFW4y+0S7Z1ooG7fZUKWnfWIwMmBOrWVT6JZqliv9gP1vgLQqZTikmoi7zbE+qM
JdPUar2arH6uOQwBUrll39uTbHb6bVhXvhc3fhXor6mZeLkjIjo5o0zW724lrQRq
OywIuVY1zrpnhdIlgrb8WWZg3EeTPIis/mZDBwE154y+V22BSzeKGwmgnacZLSB+
7Zh0Y3EL9DXx5UXpQi6aFzs+Zs0DWVIUEkrXBuDqNTPMF7O82NKLwDcUK45RPo7r
Se26wNaoqDzm4a+XZ/+3cAwSG3rjSAMyvJ7pKS0EkFn0TsCG8RTGlo7igCiTno1Q
gWzjLn2fDc/eV4jqSP6JB+yF0Bk+4q92gRlJSQ1NOWxTakwGjcmRBOZkNq6AdmPH
g7IsALyYlMCL91oKmwn0fb0eEyo4sM00jiFFQPPEG6dmyMzzNjjCIpozebKe3Nrr
Fs6Jv3VgeXiftB5wZ2JccPp+ufH3C7Hi9F6FIon4iEv3+fW1xWy8IqJoX9zOGdQZ
Ckcu99dhrCYiyVtVyE3WDqyb1dp3UXPcWkezo1SxZgljNy3ecr70t43OrStYbVrC
oKETaadVzrODwTykJDRCjBJMW5HQlSBM2FuUmKP5upAFYpUTS0/gFMeZnN5JMwZK
OGe2JNYhFkBOJkF3RdkS91k6wPNLiU+XCuNaCfPmaCdKaXhTV8qVkgFB76YHUTKg
5xPhjTa/GkrAYG6ama0wu21x04gd5qS/ub1eKxOXQjVh00GizxedwAyHmTExu2n6
qaasGqB2gJ+GaxK7TGb+tI3TGqncaXHdudJoca4mvcUCzHGQ/CZjCsvmDnmhrat5
zH1Dk8HHH9fgGiQi2/1//Xhll+zm8mCfeCRGivlwKlnctlTd42nH5okaKMlt5NM+
2Wd/Hu+DnQ7+s5vrxciqlCYJ+tYYMznjVRQZ76nsfKjRinAnJhzCGoInFoQuEu/D
cpD+QZkJutLFlcKM4m6EU8JIrtPivxF6yUrmRL3zMaRBD/mLmDmHek4jKBxr6oLO
hQGVeAPtWS7J4JZt4SE0JbKLdB5jzryIewJlvygo3uRgfKVbO81ILlDO0YmKMO8x
ZmWuL4/q1tpxqLcIUen1xfwZ7cm4ugrxrmrRGp9CR8kvBNCZycxX+7etjUDebAF7
y9YWoO1fGeY6vEGrC6cb93jOFe8nPDCnQGvCbJzQvhGLH4FeiNfdBkflVHO3jdF3
m0r9/FZ+eP74Qp0OEISqaXAZZR5MqGU+MWpLCtCy7WjSoLqg2qS6iEewMPSejuh6
Vs4jPyoWzjgJveEpPT5tKZ9vc9BMH7tPWUuwPnNfLnnL6M6hy0Lb0w/J58Dk1xEO
TdT02iDsxo9Ib9rMQY1kJsb0iq3X09Rk/iNwhlagB24rj6VjsYTNIsBJ5vgWpNEv
jpKobassMWya8QPz4xW5KsIUk4giDAdYXf1QyA5eTULUCE/HFjEI7ZtecNOL/0Ce
2feyXhpZnVK7dtbtpIFCsSFfBHAvAL/pVdzHJQMqHoQ35BdC3w4IFlem/VOTxw57
dpRepfR0IdJVMfWiKKrXyYosrYBF/m6/VrEYEVw+EcGcNRmzYyLs9k/1zNCW68dC
Xwb3ob+0J55vuA8Mb2nlQEaKhA4E9Nsch7kI/MXxyHQUYA+izRSNwxvwnYf9vwXu
ne6VKcr1G1B3cV7XnmH5+W4rYSbz0i5owSe4pTBaajQUrrFDJIbiMurq2PC6PDQq
cvwLpcCUx5+tslB3QNxaakZWFMuIHi6IiRK2nC28Hn9vcHwCcHJJ/EuBc2VA0XpN
MqNJDRAss0DFvItFTmaISOrbdOjVh+69h4G7rwhdw+5j5gf2EwvGyBNjlZ8BwZDd
gsjKfmS+7eQb5XUugJBVEoRgoS67jKgC5NL6XDy2iMNEcZeOZnp0fA45eJNqzx/1
JeInNJzAta5oBzs+hia5vMuc81aYhuAQqWqNh+R1RZ3UlXE+xxu6BoKnS/SdK+N9
QjZeSKEDFanquHwSqHVmlJ3eSfWn+XfsKR5PU+f8SUMDQHBFatphTJk+xwIaZWoV
dICYjaLxl8rSP55SM60/ViIKSeoKueSf2UWXmf2diL4DUS4RpXQyhkHXldMrR3jS
6GonFZZ7o/0ReQtVVzbMzEPXrc4G4yUI83rqyQZAw85JGgzLr1DUsPN3Qjy8dkId
cr4AYXiTMgkG6GcmrwlYMWIa64rF5BhEbcwNFn/guAqhKNBLEXduNt/JIFaxbQRm
vH+BUWrcqoX4Qy7pSqp/+vQwSCpi9FL3rN48TM1eeSOOhYUky0koXuzeHehuYwDm
Ay9h+9pwHOChgpI1TD15qfYIOmIj9ZaO1RFQghMcQ3V2P7HgbiQ8vMk33Vb/F8Ql
+YNhTUAgnOgBOhqPPysk2Cg6KMmNbS3ujV85Zd6xMwViIwjC/55E/UVilTIanoHf
EJDsGkBLVEQPoEEAxnkxtk+QEG/YtsJf6bxFGTa2ym1eI4fczMqe3W0BrZjPd2KA
dU60K/BoeX1ugpOK4Is7Kh7+FlXZSK/8eDrSe3Vzppe3UxuROdBYH//XCC3TcoRD
nJNMcjl4IsGiDKsldDtyUAXYPdNhTMhFRPz4ygatsoiTu4JFGL1gbAkqYSpGM5K0
TF0LDDYtJOdHSfR+Vfo7s2RE5UBScOeubN2UecwYho75xsHS8U9hapWD0wBARiHy
Vy3Lwm0DFoKsOaFnQqcmEXF8O0U5bQiqYnmg00E+Fk1TR7zeoqHBzXNFaFDqxXXT
3+TIfSpucJWnQArKm81Ah9MS6a07lrJSFpATymqZuk0lF3Jzqy4BBXivzAwYMn8V
pNnopbvQFZ3nUybMnN/e/Yhimf7DP1zzV7kjG5wpWsmDeQ+3fe/bbEKSrUVoVbTo
tzm8PVJjQSd5Qg+Tl/1pROYeH8CfN5FrhCcR0Px8IeJZ8FfV2oxQ9L6jNo4GF8bI
RVKPEI+gWWQ+E/atGm/NkOaWz4M9U9ZLKMC8RN7wEhW1N4QY+F/N41uXjBQyXsUT
mBagXPQFsqoeEEjzqwCaPplWztqRxmYtIWKdoWTqaFBwzNVhImTniKZrxSXuJREt
9FCHMvJcwERbx7OohLuZaDALb1cnLEyG0lMyPvTIuKyPeoxOIz7w/oq1NqGQQEX9
d75C9GOKB4uSShQQoUJ1+VgmwtEyrJ8WtMU6z1ZeX4/zEXloYh0Di72mckX0ddOu
JStWK/sJRCpYDsZtapv+cAq6ET+/Px9ja4ESanidP/rCw1N79HpVzUXbtP+A1Ha5
zpTNcvj6usdtUozyq/8pHyCOLqufBJBwdeN7FG2KfZosRBfn1MDAz37uC2rUF16l
u8H7xw68yYkt/0YW+y1i5tWM6PBcuMlviWd863VvQJxGWd7QWYfSA2BXARL8Hoc7
8ADpr05R9BiGCqNDD/6oqj7GL2Wd5ESX7GkEGiD6Js+Rk6THJ0oV0LzhDKIU26XJ
zTzfOMMoaK5z8RbJQGxdfyVsww0yEpmbBpQ9KLdydAChdbucd1hEEjYilh7pO6WB
VxF52ihNL56LbnVoav9TGD308b5dFcYI9tRd4ktUIxJ1ncRg+Knx2vcdN8rqEO+p
rx8CWNp7YkTYDQsGtJQPaUeYjWx2R0JezLe5fSLvl0wDwg/M6OciN7DYmu4tIVNH
lzpulzk4fAPrHYIOzNR1fEfdrGpgSJBc8wnT34V5Z18QZTy0Txzw/lKaifaJwWDy
8ILD7nF+shuE5rD/ezfx9UY1ZAKMFYJITYtvb8KvqOgxJxXZB54dOOYQ4YoNuXky
jesFjSAaFf2wgv6skM2rHvEyH5nGnwbGn23m0L7zAxK9EuSUwbXI/ATgqA1GZCgz
zZ2JNgY3oqA8r0p1TQn+orGcvIEsuItDT9UrQyZigvwQ39US0JyGnP1f0C0jmpcH
lUu3TpNJiKhJLBK4Hj7VJMSS0eMKD/abRyRudM3YJpAuAvc66UEbd7m1H0aXB7nV
B63tYwgcOuaBkuzW6rma8nivKfLZx+vUwvPYU9IJzjlGVlKC4nr7yHakOVJmS1Dq
5a4zem7DV8kM8VPBeA+F9DVl09njjdm2NQZkERiU3nzsomSbq6yLmz9dfp/ZX25t
QLI+JWd3z8Sn2DeeYXNewuDx1kfgezo2gmWkTazbvUaNQ3M8Ob6Yp4XxqeyCVWNw
emztFeN9dQhCUvRCDd06iprNry9AKe8I1qfOtqfqeItGDIx/2F/tzwKeoIosac+U
CKWFzKBDI6QumBD5Zd8TZT2ruMF3PoXtbnCpePPtqlqO2cLbqCD8m9bquSXzBNOG
gScoUPINPBwMoUNbl0qw1nKYcUFRnIgKDpK+6J2rAP0zYWMURNVZAEdkYh/2oFdl
BmfgBofxP1Z2fPQ9ZGkHuVz0bYIa9PptzqDD+Muog7lNkrH60dGprZ6NS3+GEGSY
vNgPtMdtvxObKI+RZ8YVGhjdia7U6WQ04B7cEin4OLciiTXW2KoMwTJ1oUfYYtij
eSF0si7Z+n5KhxiC6jp2bh5vRlEsHncBSAldKpUKIie59FG6EGa9OQE4r8f7Wiqt
gOfk4RWo72tp62PXMRpAxmweEUKuiXiMo0bBDM1P1rHpp9/nUumKkVbrzm97Xznf
+SCEphE+GKavcVi5unMtkG7sTcGknfgMRHWxNoTLkSmJZGwUp4/8TOlBXfULSjLt
xZdsgwHzh3sD2S+Uo+7AygO3syOScgJvwCE2bATxfm2g51LjBzj2aOfHRumdSQCv
OWEUkRzXpq38hQ5/ZiBVlnGiEVDU44x8c3t2au2QdDmDCvJTDP92hpElxx9C7Zu/
UW9gTeLXPetqn3qAuftm8iqrWk7VUbDOCJHvm6YCH0uze7QuFNzokWHmQjK4GlpZ
aRixJZDsczgTY9FqCLRs90mi1fAsVLglK3fE7+02QX4P/RUZIGtowR0/UYWxsCXu
3etko+PTcNm+QOJ4HSswtuKPvRHNukTQ9bAjZNi9GlHVjUdrv+4vAAR3yeer1WI3
P6jcN5Vaa6uGL+f2h0QJqSLXMsYD/ss3mOQRvGsxfl3EcwRMZ77jv1dgcyKLmxTL
IKbiXH36BBrZPxuTY6RpobxGWub3JQ4rZ994cgjbnzc98pz4UEriYBMSKog5i7zW
jSB91mqNvgXM0TXrta3WTBr678JN0lgwRzVHRjRr3JGZlcHsbcHfV5FhqtNuIoiS
CYKqzgE6Tv2WIN9pOzoJNlACn990T7e/BiWk3j4ODUAf17nkKBIOM9th1A58ZKrX
jC9YCs6RTKX4R/AIHPx8lx4Wmzp0yOmnGHsbN1114nGg0yRg3m8yCKAG3aScqjQY
zclNVofMNI8V3zSzpUdoSd2V5jNQTPAaD15VH7r6KHIAUpE7zcpp3ppKqfr2c2L+
r83WqIg5rOAYgFjpcvl9ji4fuyjPEn356Hj83czGA9Uje7JH7fVXQanOm4XorTUb
vJICGTkiEkK1HVYW5d4SxGqM/T94bd+o/bzYoI/ADs39PoYNPbloLZZXtSKtECIQ
VKoVaTBV49sRBQuKPCTHRQVHqX3PHVC5w8I/xgh2b3d9rfUTE2k47qzudyxMar/B
/xRqdw3ESrAhZW9T6f+fxOo3L20Vnxg4qP7sP6ElOr1DypI1sGMHa+8zOVuDOvOk
SrJwso+uxYUdezaPos4oGzXBhoDCR5VzM8gO/z2Nk6dUnJSEhKmzpuoezmtr/NV4
kxB2B3d5iwc/4/iM/gNJTYIIF9BDKqu3nwJczyJUFr/WnwpKoN11sP6ktJF1k4qy
WzpSIPcQQi2xfEfeEtRwZpIsYKTWtFd0wnsE/8VrrBgFxEcQNgehldMuo4WFgkYK
Q+zlZwcnc4Pricvit0MQKjm7nRr9jBwpTK8SGGnwrXw+drjKvp8wnjy/YGh5Y//X
E9ockP/I/ecJtCZPyXGUiWEaNYx8CeRkOfEg0+ks04VZOd4I1ss36AjCNfuf8uPL
rcjzB34P1nleBYLkBtpEYWNM+dZ0VeP/v5VrvfH4TqX4zgT88UWJw3Efdgz6GXlv
X5fYjT1u7+80kZBwpZMl6zwbhQwekKP2fx1y30eCFKKIg6cDJOo5FU0j+inGgs5S
3rLOp9UbPn2x3i47pLxR0kf+PGDwbCLv9+Ui/yWgn77f+Um1n7PHMLs4C7Xh0hbp
LOHqejI+26ubQWJq5zcBTV+qEAid/Tm+c/t/Eoc8d6oIqRwzi3JB+MIrRzPSIV2Z
iVYJ8sHGzewHHGKq1feeEe0U7X3rr/UVI5iw3+grQbn7U4oqDlTsUpL+c2KjPCtm
+JXOj9NnHoSveqnTH9iLQ0Gl5UaAcCEGJNuN3ux8aF5Glc6i4iexzCFap/wHkZSP
+tuZIPcyuGArwN3regijNsTwTchCvkM0MxW8YvAWjGIg8Bzpe73YKM/Etb6fLxeN
kqOHysSXQMkvSwCc1t7jaM7SfzCZrFKYKXaupZFmXcUDTz0seVDUiJ7L1oomu3Yp
srH9iNAWzvOjjt7Kkstnth5dMGKlwMhHHKXaYI+G6AP1QFUGERnmOXa+cVHlb8cc
xhvCiDHy4w9BMxazVvWq8gDSjFmmJVqrxYqO98AGIk5ohcNtA0ZKB7QErnHmj3eE
9tAFUwadc+bDMMN0znpGjEP+rNf1PL6x5+9ceyiacwFRI0oRwfJH2OsVI6qsdhIG
vEeu7lht20rSpf7Er6IQTGkgyutXKOho/OuIYLWfHDYS+YYv1PRNFi3vgKbhxYox
Uro52ypoOjhMSReGq7FgcV7V3pWpgEgj/Ws3WnZKa0j8DFeRPfXza+wJGFjYS6zN
uBTRCVCYAza0zTWsWvAqSF1iGGMvlbM+VvVDpNT0paxJrQ2EZGgEH/0HVVBeNWep
fBjFyyXSVDMEGVUB/+w47XSxFyoCj1WkA2qvM0zrEZTO29jvLtaZkdswGK/byQYm
6XAaSkqf/B6gkMtx5DoC1u7mNZ2qPEE7yIQwIJN4v2w4a9jz2Y9m+S1Y6+2VNouF
HhM2D6AjO2JBxzmcvHMQAN5WHH89E2p2JC4j+ULu1cU+vUxX+QmBUTVQxRYl/gY5
1cDnwKDXqCplwCS7v8HPGycpRGxw2B7jAjI2j2pKe4EvEnFxyeiFuLso7g3SnMbO
9jFELa+UOMeh0H1eRtXjTKsNE7A71eMds4ARtEgw+UconWM7USAx3WfUHFLGrovy
ZEN5iw2wELjyD8HSI7LIier2hPycZoQRz3r8ZJGalQFmSZaZkoe3FfT1O8a98mVt
do60lIQmew8rmbquxv6GWdl433qGwBRgeuJidP/SdcHvpAsxrQ1KAabASmTXRFSF
RFz+z6Gbf8OBuS5ud3ps80DVgwnf28SKknih/i29w0LtTG2VcZ9IG7qEiF7DWjZ9
WQIxTLTvrI0eJK9alsJ48ESIDNEDisOwVbuwu+z7sBO2mwoueBCYV3mg2/tYNDGR
Bk1ucF6lC/JZCl66A8C3K0PxGf9u7yzZFsB6Gw6+DIdxXdtP2Qa3Te6Dzk4tRQ3S
UuHqy3CwtqWxQJq7vuDxesXq3UIc1u4OliN3b5BB/iOot879amMe1DczKMj95xMh
UNfFHiegZnEXSMXedq+O2voxbNQgyNbedkTlw0wVK0C4ET7Crr27tJTivHk3+NHC
Oa90zD71u4DLN2RBqwOdFgvv401mWh/THFogShM6xbKA6cun4yUFO2iiPKLxzqJ5
jk7U4E2yjfpRpjWs46ioMgN7Q0VS7LOH73Ab7tMx7PtJV3ix1b3G/2s8PY77EPWw
TNNJDF80TeSJMN8KipGH1nFBAPo2zgeNKWojzLqlD/pLi9N+Xn3uztCaQRSCNnWA
dG1O23++42D8cOnW0cOVI0ZpupIlzH2iMpT5bB27Uqa8oUrA4y+B9VULe+4RRCEC
mssbRSM+mudhUhf8U8PURvjNMeYtdqqktUS5UR4k62KlXW96M1RsubIF6iVUmIos
tvxXal2kz5vVPzWWnUMttv9UU+Tqybs2E7AX5yZdfx8o04LVZuTyGF+iIruDJ3xO
T1lwfZqMRI+OofCdu7jOmrQ3MHo1ME8YShefY9Cr2jEgZXkhiyOAR2q4T0s2XuVW
kbUYKW5eFm4RqW/EwhMyLi/XHw2U+hPxzRR5LN3Am9VV5zRtND7GAGK2zo6SbkB9
2RnRcChezafaVVsXfPE/w5wy5Z9caKq7iTAm1idPfXo5Lv3m6cZ8TmOh2/EI6rP+
omrMPVJ0/PxFQ9QikvQ2DB1Lm8tuD8D26/VCxPntqv0ta5+x17iYHBc8Nbz/soFg
JUctgFtvLxM1mGWjef8uu9aqfRW+dQ5DLANokxsCtVduVKhBC3BLWE/Uth0q3ZoQ
WpyUhak2ZXuJYam6zRfGpbKQ24sGXD/E0Tkab1/zznUBWeJOt214CY9sZ/fYoqmt
JJAF5HiMb3mzlDQINJdPeAaemstSqEf9L3cO4zQnDKF7SfPsg+J8cVrEVDb1WDky
vjOxAa+tBzfd02lBPDbW5vbt3fH8Xb78neQl55CN8hebXjAloKoKTvYCtVR4EkpQ
T7ArF8QX7G+Y5olKglwIHlkqeaLQvKVgfxrz8q4mD+ef8vWrYyicfBeY3w7yQ0fV
5UzM6vzXSaYYwOOmSDKHdEYuOy5PL3JPHIObH+IVDppFHmig/r6d5FCiXp3TfPZe
GHKaZbcYqL5an+iMczvAhXY/5mjyirOuwls4UbHxlOt+OxJJX41pZD/sqDPJJ/rt
Fp/pPeZ6inXKEzzimwsq2kF3ESjSWvAyDlKm1dKLoB54Y/sGwDErcppdQDVADUBf
fURhIWjKi3nfTQgAw3OIwVAAxZUt4DE/z358DpgBFS+8Qi42yxXVM8dlh6zvqUiH
z6X4DqA93A+nB++pO856NDR+nQZZA4vzNojg/T6vtbCcd0u9KyM8cNeNF3/pQUSH
UtTcITlGtKwOS5QlniLrQ5kq2Dou8c3teas1jwaqBFPJ4E5tEaoXHztXI8lLVJc2
fFOticm5TCR7J5GscKCudfsKdwLF2yy4I2+neV9n8WXka0uyTpjAiq2BIwaGzYJA
NRpQ6atyWyCvD+tGgKrpLcFtAY59QVYJH+sOpJvHDd0+5X+mA7mhWnxgsOkzl8z/
4P9KZ39hGn6LVXmj1CjAwgG+5QPCYu6IGclFsABPQaCqpQm6uLRh1iHk/Sn6McFV
yQZAmbecxpPd3ptWBlH4wI4Q2jnpBTd5fA8KjdUQRDSnhNf6BAUtqH1fGzbpJfQT
zIP/n7ORkT9nXimwY+LCwFLcGhmunT+GoV+PJ/nXKqn0tA7WBHNlvTlt2mWPYrB2
U7sbmzcTZ/IAUkVAOEsznJR9BgCzTszNVK0ZP8SKxFvbpfIhwtxv69B3Tkqv31j4
LzN4atuFAyj+UGUbAQZsyqKfVKItQX62Ywq7wUnzea7u2mSyUBIwNWfeXH5YY5Zt
Fb5VA2VbdhUiMKUn0T6E/U0C0DzthcvIbciPZqKYOhiYJF6qRI2psYzdsinvfHBJ
RG/P0RFZebbbF+LglUQS9JQGyQNG6+i6qBQmnU61g64zHmeWs+uGzWAOQqC6mki7
UQkP1s/8XtQqG5gwNEYWHBlq0+7p6EKPgAGXfMFK3aLVrpxFtuDIORyE9BhZnjJf
HsR+S2Bh3CLe2utvTKUksi5+fAqcxQebQ0jhF2HZW+oCbt+uQeeN/nbWabTiw3n7
NFzj9oPC3W6+J6smMQFFvx3OluHDZt63BN4AjOJ4OiXhr0XcKy0YkuJ5siDKFy0M
3PdR3kX8LLN/ga1nPOQpR7n8sXBQKHWGuFe6iEG2dMsqyd6zism+V+FSvzYSFRHl
ZEMv8nnUn8ymZocVKhfBbzQQg0unk91W3hoyABrVDs47LZie7UgBo5Dm320wapO3
MLkKfawwNjOoOqQ3YcgYVCcFggW99yJPBn45Eu9kejFz4genoYYsLITRL7GycvSi
U75T8wmDaARnPC0XNs7OS8k/9/jb3AZixAg/G4Bt1yFsghJNVmB5GIPhO/NyyXpp
d1q8k54YgSMFKCKsgYIbUCn1EccRIDiM51QzzlYlpY/1H/Y4jTRjPYvPTZrIXOy+
27X1EUZ/pQRVHkWMlgnSUdd2Cq7Zn8ChE3QLr/Ht2MdgaCDpeYC07w1VEXIf9ztP
/XPPPIOVcaodkU4u41MLrlizAwJbLCXneiJwD4C8KyKeauSTLXYBqCGyv2/kQHYx
Dr3G9UMhLPH7NzPHtUBvhMPguwJChWfwU/CWeCZq4M8KjNBCnMdWd7TsNGm3I7l5
uZ7uRigk74oFX3UMQapnl4eHS9Wvem/y5vhKUDwHN2/KmiiYGJEk4mILtpz5jVLE
/A8lN7R/C/mfm7YgHHniznHHqs4x0SDUnKtJfjtQ3NaR8ThnYDQUikk+pirHcBJ9
iePKS79lEnTah06ElSE4VFgzqonCxp5yther9SNzWQYWy7m3E3Zxobl5J0cGQ//K
ZMgNVOgsGbM3lNA6KijJru2B0poaxSLXv+PT+vxNJ/c4oSdHE5EB4gHnOfy8YZ0H
aYVV0UKsm/tqBcSjFBQngEwkqMrRGcnijB1LMG2rvVAJ8U4BJGvLaPOF/EJdZQNh
TE0uhUFnxO2irHUVF8vZmFK5CQ1DJClISpswj+VueZOnYcTuDHH/uAhQgNUwDgGt
WXwY8U/5Dw1+CEhh0tKYlDVvIKBolF0M4b613MAmIe51ThnLVoGWjENOcSl9uvxA
GyeW5eQhNk9xYkwnhzJu1SCfGAJ3uYGVPJY1ZJ9gOzCCkPK2Vubmo+VtpmRYlB3o
o2kKfeEctNJ/LxQwpqtEKe3ZkwEFdRPvTnHQryKVXVLFCtqwW6iaDpWSf0I9IQvL
aE1FGncMdSKPRHIcwsgZ9rmt5ksgjCut4lSv8WVyv8SsmleBycOrhi7J3FnIcO8h
fsMDqUe6sWyWw2+i3kiNdMTxvMGjhpeGANxuC5Z6q3f4NhlJu4peyj3Pn2dd2SvO
ntndVCin6rRZY3CH8nN+ANk2nIMTYh5ImKE8LOfeGwYx9B+GjHR3f5xcGUVheoci
E4pRLE9oGVKdhQ53CI+WmpmAluP8mQb7vzODBCHTRgnaU/fnJ7KNU8l+CmOsFMzU
4kPGWnOn8oNCDi2U9M1vwD7O630vhoMlZ/8o2a7GAq+lFxynH8CSszRzvRX4y44n
vuws3W4M/GJh/sRl3TP9m5tqcrGuCD52hXRgm6qRhfn5WVsNTqO0vEnyt9wawz2j
i2F6mKoNBGc3w3twCTSiOGOw91HRn7YA7YdjuVixngkn8kKRvZ9O3vlgU1mf7l6N
sAvx6JRbTJznZiil7HF+WtNmn+Cb7zz27MHuVQAFEG/8rZ+hvIzpEHawPDdMhjoO
cVCiUAu2yC9mbLQ3jFbPBdkqOJijTlQ4w0dII7wVQpXEIZAPoyBUm4gI+S9oqyg3
01wxkuzjbJyN4nX+2SuiLm2ylrWRrbUlpHiVZtNBMFEZoDAqx/uqay2bihzfOmRt
BrbLWCVqQsqlztNShDchuuL+N1vaWIn+f5X88N1gyEvwmY99RPUfKzAvbHgeaqxB
R6X2PjMiN1d0+58JOzggJPVcbZwDpnyuAARUMWWHLOr/zba9DjmFPUayU2iGfBzX
oUOnDPKitCpl4/a1BzzRtDUgp+EpnlakQBW5hIhqIyytOo14JhjDlwPlqiq0Jqgi
XESyvDgSvavp/Ukhj2zjV+nVKDm4kM0jrAgetmD/q+EngA4i2DrlEvGWSsPELMNz
6cMLQ09FyWuFoebKadBfTdGbV5+6L60nvbK2fvrASjjsIFiWsehc/2WINSLatdO5
EzVkMxeJpgxCsFKKCQjl/PeI6QsXrBpJiaJXzCDs7/ePsSzPyFNjE++Wx53EgFz+
YQsNiH/hBIW0GomAza4RiI6kpMEROEEOgS3lnZnGCSOVEHsYC5qC5ZcFXKgp11pD
Wod3WcMC0OXkAh5BmoTDWQNNhGVte371yBUSKai6/iO/vScaHSFEI8U/4T6JjIj+
nd66b51q6UrwzEQymXP6uiN1pWImtGc1tf5zxng6xPwWvgcKEVC0IWutdwtw123c
G+GFUMWFngZpm1f6DlogoCu9/zZ5srZRwRw4nVkmGjh79hrOcHSzQ/IVSeIc6C0J
eeSj2KA+mGEfTwBYN+irlZoSNj4UOcx0FOyCd0pp881lYslSvkD42/XFwqlMsQ8F
iTN4+EJCUJ0I9+OdlQd0PXchilDcCbUKxCwGqjzrkRArTsItbB6CmOaErzUH8Mru
gsHB4OAf/csKvAIGXepz1iYl1DpyiQDoJyaTF4+9Rz7WuYnslYClr+rtJeMWCMC1
HRg5J8PfTwOPASAreyA6rPiAGvnLCe6aIM/V2ffxDSrfvrfxa4ve82Exo7pqXWN0
bL21gzVaxDbEjHEqmu38yeeiDgl8NNzpEkTHMsHARUhDVWsos9ljL5p7c4cFQWGu
EgUw1UJKFI9DJIF+hp/y/6lZKFeWelJ0J0l6eND8HfFF99goUw/34mQnuh68rZnb
oydfw3DUeg6/rT5zBeY9KLpwwerKUeuOfbt9JGcH/Aw9FBLf4pQGffbMd4qkDyLh
0goIjwDEOGVAeTOJ1oMjzaI/hHg1Qf2cuqU6gk+dQX+Jo9pne8Af+hmMy1p21eK+
PZb8kCAP8sOJEw7xKk/pt0vOO5iA791gbh4RQVsU5CJ14DrgVHU28c/XRg49nbKO
RGA8q2i0xbU86+U0EBDZ6SG9gDz+5P1lCwLSroeiwd7jzdG9GnUjt7HO/pUQF2QV
WEn61XTRFXhky/Fe0sH2iaBqsHXd36JhUHQtvR/QURhgLGARGI/zkvt5MNUboExp
rP6g5u6M5a4B4DK1gRKGn9CYR713Zm4j9Q07HhZFSzqN0WyF/jjzsN3Ky94wkzy1
4joEB3jF3jTErVdMu8y5QeegpbQ9uLc5X78Cb3x5QSJa+mKj4604VuzW/u0ZIvjl
fIPkkI5QBEGV5TBc2C0v01/VxyWK2MqMFGrJNVNDla1VK2SkSMzLkilYDBpzTevU
cqpW4aL4WKIyT8wipyRidSjWkoqH5ZMxsDKMcKDvYlhFTAenahVWrAU29e3231D9
dFV9z/gHL9d3ss8gzyMULnN7I+JMIDVmmPU+bQT4SZTRQ2Ji2ZjGpX9DZ54YGhR/
rtFEiZzZDNjNamESi4gNt5W2HQF3nBhWytBdSst1Hi+mM9wwAlHpZGobtIF4JEJw
P3h7y+f+T/Ne0v6zMfzcE5t0Ppktr6+6J/GFWu8AscVZcmEPuW21R32PkpMtnmVT
pTkKvXEnNY/Y1Ou44BB8gTtkGAatcPqaGE/TdfSWqqLkZWUtv9WUWXu/AVteWWbH
1BtLJ50uEGgEH2Km98nqx+cNuMuYCtBSA5LiAoAi1qHvEmkwXUbMWcGCcNd/NZNR
vkvq3Vpd2JbSdgpaBLsdL5+7qcVxwwEQs8MZar6sxmmIZZKL41gAutYKlya1sHYh
FBsu3vAdvyBezjhaLhakEyZeaJepqla5h1J+HrOgR07pg/rnx477O0+KnNZehGua
yEqPWTWEo5MYRkghAC5AOGVz4A3JSy+t6bLP/FjScuVG0Bz+KNQFd1S5XA5lPUZ6
vUtaXArc0FFWjMFXpdWULRbK/rZDARKvWRHHlkTsvnbSB0z0Oj1+CGxWseY8T8AQ
XQrPrbc4LSdBh1B6L7bCXcLMcexAHD64SP+s244hMhr1gdCSyWAidbQlQCr5fRjH
0dDzl5FG3yhnslMInsJRUgYjUOtPgeUTknckGd2FRGiXNVJIEkH0j3PaqGhtWbKX
DiPmNL/G1qP/P1gP6fvzkX7F9D9WHksP5Sfgp5vgR4W2dSzOs4C9Z5HAdOhRDjWm
pZY0Bq1y54OaXqthpqVGAw/kxSX8HwO5y+G5Pq1j+NE5Qm64T6YD1e6PlRypVPVj
62+sL1kT3gbL0CAIBlk1bbk31rpn8gbahuCG9FlppJtKwboBJv2YoePbMJ6jo0K8
hD7kkBWzyjyIv8cHo8ndwAh47BSBzey6elgxYjyR3cMpJsM0YPC56dw+EWr6xd8B
Rsos10bz2ig4D8FzzqFLuOV1B3w9uuAI+44npGw27UB0HhnEkhNYqq88P9z+JfmD
86OBJGIou6TVVl4uWg1cnGr9c/4UsNCM37kq2vCTr/YO/RHS/kpFf/IjHEarmUCJ
Ak4jOccE08XKDdhBEn3Y1lbXR7ePMclaBdOdHislH/nFFDuogv7b/grIMK8HsceI
8bw27q0qITN0XhFGLD3uxU/lTU5jOmbXsXJKT6lVNpEgwPeZDuASGZe43xQNyXwq
s8OPGjDrFiOB60WTnF35hLnG+xmw5euIy/M5dKCfZ+gfGyzrDVwdt41+fGzc4jfD
5PhGqJdGDVwjqnwroXskZ5M9rFniZdlF/hdMCJNMks3ckFXKCgCQ6rawDGepy5ot
e7ci7915Ep1uAH/RrWhr9rfdO+a3ifWhrDzgM5ksbAF8FxPlzXfQCuxnQb7XipnK
y/cnRbsgRHJ1atF75Lv4TVQIn8Bui7LKWTYdeAauivniksn2EZ+Li/8P3on5Q55L
JONYIyQssxpqsTEzOi7mSsDXQSLMQida45saBG+0fqtI0IqauKPME1t+MQg5lO3w
FZ3GwkxuKXZ0KLDVirp4ctnSxrkzfl6CqxxfgPb9fjZMDMFKNHYPEJmQDUA1+Nyl
Sp6Bs6TQZTvG4lTyw8WLWnwkWoH0zyMQBilVMcxqXkFN994Ilocby2XYGobzVrRk
JHXXoN6jfNgQkLYsg4t4Mf+HRvbdzbat2BbcF8hHvYDB61VKspVWY2M7YARpIVcu
Dj802wuFxEhUGslkQ9stKQyVNB38wj5D0VGc6ff0HiXMXv8o3MTblkNPVdi3M0u0
2/OSZrZ/crNjE9Q5wHAI2RvgQ+LAZZLR9lwZOL6hMB8Hi4BLk1l+RDJvyRhAHjaj
47dnTrtHFU2nV6yq7E7xi02FUF3U8vegKVpd+E2+2TNZtgki0xYz9dxjQcRaw3Hf
MW8p5nrs/GTJgdml9VxjdtplExiePCiIFkBl5Cem6Yvoul2aXvrAbL+xTVlBO9n9
3cqVD6tbwHiEavRnQejYS/jz1Ui8kjFFbF+EV88P1bknXPdYx1NuCj0b11XCBOTf
HsoHdUv1Zs3kd01gKNqYB3wEqziwYtwaYb2z3KVJpmUTvA1sPZMjYx6WD5GaVift
ez0Un/kwNfeR6jtLcTITY/rD1Ru1apfxYDWmxz2zA2LCUlm4bddSSkes47PF6Kn7
o5GOqFJe4yY+qa1JsxsQhRe+xbeo0tpsfl247myr3Y0wkuz+mqHZcJlEDa4v0bgm
RjdWkP9hpywuMQ80XgtpdP5vqyIuj03SUzlfYvhj+ib/67KHREicqVkbvUWqFSqw
Fjp+l7kTLqTHwNHwzGCX3tnuaqYhsUoURoHSbzQZHjmSZsec0kxDzSwy7do3WyuT
ybYgXvTzps6I7kW8ibR1Lsz+HhgzVW7P1bJ49ZrsiJcVeEWzdOn697cylKaf03RT
eYN8w3+jc5iTHQTjH9Uh/BajxgOoeOmKXkYf8XsDWUjAEGztrS2kNWj+1hnVtmxJ
Jz1xMfGX4JHC1EQ8H3hh3SJIQN/+f1MuugPWwoQ4hv2h171T++lrDyiQNL1tbKxf
ddh5I+yWVIgejPKj78l3c9YkxpRrZmfEm0+wKOnSovdXi1MKpluve43lRC3gdQTW
G9sRfzWYvpZJwPlTdfx4+D4C6EVWLLaA/aLTcashSRhVWaSZxMfIuiYC+WPDI4b9
9RPTk+l8CAixfwBlstfii4rFlfBQCwSiIDSBnoKMroQO2mJmgpYsd5moQSb1rRCR
11AYGqbkcl+6muzZTt6xCTvZPs0P1Su+Zn/2Ky80tfEXTbqLTCd6a0ktA6gWZNet
JPxmIsdBl5KgeG4j+UImKm36t8UhWEoHEyq4I7d/5c1+SDXURiLw3Uhe+fS00fS+
RVZMvnnV74LdtCUurtRFv7wLr0VOXdRUglZIk6/FtTd3w75M43aoUHFWVBM9UNDY
GJ8AlW06QFrrq8eJp/N4FDNIunvcTZkFgiDyme6v5AFj/joyPpXHtkQr/w2KZjW0
kOWjJz+/7SA/Cv3nF9t+UoonXq4rPLfTAMMJ251qjzvu0pcbyY0n/9IuWjcFHmz7
UCMjbBLuW0qFsA2Z/djJzCz0jQ9hQGx8tIXzmw/H5tpIj8LpBF8m63/qMpb0vEIE
9j/MMKaINCLGzZaLUvHOGdxqEPf2uZyrnmNUW5itnK3ATtzqZ9XQCAeTR/A+7AAf
6zpayegL9vkt6VlWXt5qzgbiTFig3qZipCMFg3y52eHesMjwk/Vo5UnsjSShOLfv
H7muV8uCOPzzZRBM6jG9KRtgual+oajObTPM7p7/O3oQw2OWYR5/JiLahsv9TB7q
Gx2jHJyWAq9YMzqiZcvs0XdRr/Dfvmsbs4wS0o39Fq9dgsF3cCunbzWjfJ35B7Vo
1ccYTuRLyeYOe/xnvcs2lst8uEVtzWTlCm0Jr9omvtIgjqN7ps0fkwPo4iQlEWti
SG9nT/VVENA0i3wmUcc3h8QvrikZUt7SFA5P8zJfPtP9bGPpwyWkmCe6nLMuNzEQ
7Fe7K6LWjwpW7k5ra0+lGnav2pJm1OZJasfn8tZn0gsQaF6EoFQIgPs0AZ9AxnHv
/riSs9wjX4bpyGqGTMcLh8uH8SvHyfwAce2K8hk3Cn8i6rQgFTiCOPnE6fK1B6PF
QlaudWg1JCDfy7gDE94xXE8K3q0ZCT3wICeUpN61lfRXI+WgBoGhWhXphB4HxsS8
9LGmI73bpmataJ0K+8u4KnOHER5o0FQPh0xPx/SD9k0P10HLhLD24Yygfa78Oish
O9iqp1etG4VcLFV1lFpIvOZ5YeGyqher5xOAFaecpQL/AkHT20UFbRpFwwjgctiO
c2m3i6MtsmWUNNsAD6SNDEZXuYwYYsY/tdXJz1bu7m0mKyMSPsgEAe8IfsYqthjG
yNw6Aiwy3mLx92ekFdhIwMFKWjG9NRcQZRSmVOsEAgvkRjhTwBrF0mnG0XICBxHA
Xdt8tqaV0nUnN2lKWVCR9SjUdkN3nV4DgtpVGU1t3H7aukPtTqVY0tdRgCxINmO5
/w5n2fagQoiMhskQv79kUxJFhmoY9a/P8mLZpoGtoITrECeuAwOOEapQ2ErCc11V
MnBHPFjnvQNgWrRWftW6j3FI223whdI7PeMUN/c38JS6McOFApJOqiWHpR+4bd1s
ifsdw8Jlb7g3cVfYy2ShsLCvtzVJDg2IElAJpJG1f5tHLTTeEUIICUCBYIcO27vQ
APFZMhvh5YwJh7AaqN8NLcRnuLKytm5YkDvoYSbEg4klLYtHztvfQFrDURqRjtw1
AezOt/qldJnUDBFF4tZSemLtE+J/BEfS6y7JcJiWuWWR0QxEqp3px0TVUSA5aIKS
eg6x6+uH5QEHh7JAponTEgjmy+MBLJQgf+uADJyo8XNJA8IbyHHBxS512yl/Y3Wq
2aKgmY1X6VtNU4y5FWXr14LJByP2H60TS89IudC13cA2aUzQQBjKBMg41Xm1w1Mv
xhlydWF+kmuVDOcdv+B6Sb8HBcER1oI41hiH4NSMk6TwVdQ7FEwVYIjHRNYvB4X0
3U5Ls9DWqnkVQr611rINnwEEGyS/zwOPmr84rLAaeZrbja3GfTDBX4Z0MwvSguzf
r8WNBfukiM9qHyUsbXhUKAIv1CpuiL7ckPSaE7eNoOevcp48zeZNvidCi4JYvXMu
Y6N0UVB0cJSKQ5cmggEY6p3m5p0XJo+hrXlCZANCFgTXJ1mCJhrh1tieVPo2OJu5
BH4yyU7x41VeKrh2vHREJJNrY1ULUN3HSCvYgOJuYcuaymHjUP/JoDD3IvFQJBKq
HxsTXKHz7+Z4KOV5CbMv6a4VwTpwqlCSmS6If3pTb/9cP0+905lX3LyVhEOAPKL/
SgnYi4h2161OrF9kmKbH4kNjxz5rIxXsbeiDByt5KPa6ws6as/JrXIXTKevLxnC6
4INyWG9fqoHnTDbkv308hRqVwXPBbKYZ8leKzYB2YQrcAUEWYj78huxrVrKusjnV
q0Q3gZ4jMkrNG3bRdFDGH4lkt5qZkbz5xTqUptlOgk2M0yBhV296r2jjq9ekRjJn
X6E6TAHG8zdYFypYbJK7AQfuYu32qFj44TERKhnzpjDxZiN9LopWoFs6v+/2FyYm
pKXxELj1xlQLnEpuwIKp6E+tlmswbo+LAYYLaTs4QCO/iWUyFKyU8kabzGAZIHaB
2hAA0/gflCp636DbPwRVHA1gyPE7JPHMHNi9XffXF60dgK1ZJejtv1tuDNK/G2Ln
jhIEIk4QNl/ikUSNPDQEjvuXPo4+VB5DSwGp1P2g9j2W4zaFNFbYUxTOKQZ3YNjS
Q36dml6YuiQcnG2xSXnOdUE3TfUF28TBs8jQkvs0Kn/Xg5ak7R3XfkPKUdL//oYg
eIQXPttWaRAhiw3hA0z+yzb2FwzgbQCshabpft4ECqQx5/97gIPLow9OAFlRYTDP
RYjM1pgy/z0pC74hHLIGYs7mt0fFXuuUMOka3uP+9l3+k0o96IZwz072jRksT3nz
78hdZTDV4q1DebcsqTdmC49Ol1kyxFbHM9ONWmcI33fIKLtrUUt0/W5l6yoxcJ4Z
uFGkgKAubuYsnLJXakCdDDyLS1bSsVLX1lVrweL0fKzoaGRyy+9xMlYctPLfW2Hk
MAX6SG2LZOgt+drLCS5UI8oVQ7xWgt8K293j4Zr3PkOls3cYTqTBLCUNVZONdhP+
geumqFPPEA8EKQL5tvynmAcoZdGMUK4Ka7Vmvxf/7vcMx81ylnd8LF7TDLKGa+bH
sOrr6aprvLTBn2ep2orveQYsbQOe06FoW8e1gM1AVPw0ewH/zYAPWCo9FiK2i+j2
/eYzPGeNMkovISrOqX+/arzMugg05SkUOKJFDQ/XkgN1ggWrrkwj+DqrpxvMSE3W
/97BS2Tb0wydQ0J7aYL2LpZ+ILW88GDWUSY67U4phA02Vhy1cSnRGSZOTDPp85fX
sICCQB1fzqhhAvBXEkyyO9NWmxDWXSXBaT6lcbSyqiciLNwm37seMiPUpryuvDSo
cycMSHGVXs4anygo4g07+dPejHYdK80NHyB5fL+BGOb9y0ruGUDZznXKSQhktkMG
0laLORF2imRe6e/mcF85aFLsdLcMsaBHR1X8Yh+i/cC3RFbtk1jjMCTCZIkOV5WT
ntJuedDC2DdnOQmLhrH+rPQtRb/JycmzqK8HvBcHsGwzMm5slASXwv/HHyXY1OzX
HdVGJY6Tkr7gGgcuQFW96TE9J7q1R2S47GgZe9MBNfdlNBNLABTXmQI85w7YL3KY
M1bwpz5YBVmgfwa7+exPaU6IMu+kC9b3ExsvSEdq95S9gAVDfRJ3SamWfGD3udTk
6MKn+amd/VEzMnA0O6zMnQBZ27tny+tJ1LTqA/1leX6Buht7SE9RNlM+Xsu89hW9
LaL3EA5qphVq1fTmY9fIWWH/i0aBV6tEzrsEBNWdIuKbgB5M7bIPUqRyD9mo9CyQ
aUSchHyX0+LiyydW2ddwU7E2nq3KDsqcwyFew51Dcl0i1SFrOlIwaP2LIIIuX11q
NUAPfV7rFbS04t0TWJE6ekIrESYDtYrgJaZRYdJ0nIREIy1+BSoHUb04f3iTRMwA
u60CUJo3FrvK2ZzgiqUIfdQUa+D/m2A4Vfpz3cVwzXZ7rhLo352dazU4YKNY0NNk
4dy4BmYzKGu8Vve3FZR9GXF3oVNhOm6eHQB+1pwW3aLhbwEbqld8Z0IUTegYIBK5
OGRF75vCMc/FuYgTWQarWb6hnwW/iLLr6aD65AgL9QSZ1FqKlMCEHRvDpfaijQuX
j915+EBMK359Xe/NqPmLVg83F9eAVzcnua4eZK9Q9gAwLL993iK00vpMIvW1EoMn
kz+nQQHaMxJYQRGLX5WM8Q1g9K4/D3nzVSSuTju2KyDV/nTIbrZp0sBlurTl2q3C
4PrQFySBYdhPmtQcr5zz78g2FVfGJRiNmFU+LwY8MEVQqWD4FNPdGaT5qQOnWkuO
XOlTbDMsOBO7PH6JlHLWvbIQfyPy8XSy+Ss3DPVgEC6YnnFyoKaghs7j7/IN1IMl
WoDTEmICOiVSc+BRbM8MjBktauB4+SUvLJg2R8VDN8UrsIi3Wgi1PS4LMcDqzT/p
RyQMvguxUHgxFb6mvkVZM6aVGzKX/OEc8m0BQPSdmP+Lp6QhEd38+XVoyNi15uuW
Nr5VyiTw3LajxjDwaJEqfEvsXgVXdr9SfwLxab3kkqYwxIKNuMvKz70a7NsNYA+m
hVXlB0njgOtJAHJqHqSpRf2gU7F2HtEqNZ+3Fio5DlNtqA2ugtWiUMp5Cd5acU9Q
TfaFs/R9J1md/erHrTWj3RgOdP1P26hUOzWDS4+exnWy7YDqNcWfBugAxCFYxVXM
VRiN7aSFflpvY8RLCmVWCqmt3H1XznkQKGjK4VgBSV/nDVLWiQj+Z0bGS3WdT5Lb
C/WFf7sfS02RPn16a9ST6tAwIBFAieRab4QnFaiT4c8wt3EeclGJ6psWzjMmrXiS
RYdhfIDkMqhtQR5aPUARRlvG5bwGIYS6/+SMSPnuKZdjvEyXoGyeRI7DPzTNY9Ip
9a4KChdJBJ62YIhUTbvT99tUxuW3BhZUzq+IH5i9fa6BosAxmWSDmPnK1iGNgwR4
a3eEbjb9tZWmiEY3PpeensHdnCClHF3+SVPYwLBWL80z5fQo/otEC4f0DKBIQ29y
udLpRBJMIAnXfUWqIb4Bd3Thq7/cbN543DlowTiy4ZYlZHVJ1Sph74F6jH4Zh4vn
QCXCUycuF1KqXxop2xYLqckZi2jGvL70/W7B7/2gsx1BVm/tSog7uKceMGsHrSq9
Djx2c4jp+oWQvlh2mro3vHrAkfGX84YizJ13zbukmqn6OHjiIJbOnBrT98pixfWm
74m4Pit/jA24szp0NfwVKHl38HvNhm8O7daDxiBjF8k2ZSi//NCGmEke1DkGHFia
qVi8tPyPFaZUA62yn9ruH0lnIJjt4Zt0q9scXSK6N0GI1jiK7QYkrVV5hwU2hgN+
dv2VgX2rPrn7nRmS4o16SItEs//lmROqIuqGm0aEwRLSTHkcEVM4n+xvfZN9lRtc
Srob2sbTgE3KvroUs+mk379OfMxGVTtKhdoBVj3OCQZs1QpD9G7epxq+AbkvgA69
rdop94/YsDyLDhBhXcdKdTESbgie5q1QlcIp6SqVFm6b3z0nNw40mWSmsl81+lAe
sSZ8qwEC6wVdcEyoDNO4dFIW94oedhWOuYqthBeZ1/59OobxujBBe2LVns3i92W6
oMTdU8ZUePjxg9CqcUsU3qie7+tARF+TaigmmG+kCB5v8WYTY5273PlVNtat0AIs
polu48JR9+Sfgkc7dWF5N5WtnA5okdFx+ykPx3pEpeBOje3FgUQso2+2X9S46Xi4
9j4vVALNkmZSPvUnj6GkiiPATnnJXctv7qcxVY6pcTgBLB+hf4mmNY2+pPbmPc9j
0iz0PSNsL8+AxopZt9QWTcwvgW/XD2AndlZwV2z6gzY1oJdNi6bF1OFlVcuW0cMa
bIHXY6pxtA2bl7i+aP2RL2nVBlwKq68sPNLADmij9gSMBk9xNw/qFylXDcJPZQrG
qC3m6HhFd3sYvmUpEtrIkdZc7vr0EdThE1rb0azut+P3Gdoo9ipCitimuDPYSRKU
rDvHOgEW+xBaw6ZdlpZ/gdV6RG6qNQxrVrv9v/2v9KDHDhikMoAK8jqgt7f65UHL
F0/9Xg7OtexW5gM9keB4sTCOKc/ePTzeaSg1LvUYMQdk6z81jnfUfjFe/TlCK3Q6
phd4VM/ud2JAD/SR4KASoSL0zMzbor7ux4DLCekoxE0Rk2I1aVJpZ1lcXSmGFkNI
6F51wVmkSl/RJ2TVblk9+W3/Bd3pyflX2Flg8J5WgLvkNsKJv/GaFplaQWYgnzGG
EktrxP72GKifCsCR4KnNm0wAl/jIVE/JGVsOBzSecjZoNnq3QhPHSP2MvAyrTSJk
fUQHw2wajCWWra4zZPS01I16s2GHChYhFfUB7esRO0HLOofXxyDqMba+9R6x2fwC
u9G/+OfnnX5GQ4xTnJATFRz6g5b1QDfKn/PNvOSWxG/yrpC/m7fs1fwK9nA8Hu4G
e78wvKw7cj1oOLCruPKJUBfnmBMw4VZisGL7VahDQfP0DQeEblcvrV3N3q+SXug/
44wPo7pqbA9xuzj1mPjqJabaQdt8F8MmdSm34+v4VbP8v3rxc2OZREoD55BLqHAm
4M5mzwl0djOXkFDK+tpcb/4EqyfwCYV6g5z9Xo4pCJY111ALW6ANn0gEjqVXmmQq
evNExDLGTkrtFJLXh5bV06ciiTJThU+aV3CdBRa1qg99mmpplZUt1GYeoxUs9pU2
CYAWV+3QK2uuyHY5B1h4dZ6Tfr5AaGD0Vna3U1P+WwCWOmL8szGWD+hc+wIBRSRd
i4DVh4BMKZjJkU6e2Fuzn0kWjnWyEN38c0cOJwxUfd6+/0HBPXcQwppQOdYtJJ3v
Wv/ZXyecbUbehGqjHpynUKgQsZeOZ1Vn8ey97y7HJG0PUjHb0hmy7qJQq1cjpA9W
ETdUgOqs3/PECX02iQS0WJbBSj9pQz8Dwy2MGAnYAZXLlxwgus/zQM9sEFxYpsIK
YQdkArmxOyvCmJmQnUPdeyJMpBQhQ6Wy1v4ypR5tGGBVpdAJtWpQAOiwGWWlmbWX
H6kEQ82AN0cAcIlce7blYAxi6paKqLdUZ0zTgZ7a4AeW06sR8MnUms2FxXj+DtwU
13KW5Z9e4AgQAa1OR1nSZlqAvFlmODyJ/zpLvThPxe1tSyToitI1J5EFO2k3B3YM
j3H5TH7QZYprfj3n+ENkdwb/33ftaSkJg59CZX4qq34O4eRMp/KFyijaIuOK4pgD
kl0DGGizZJmY37qmpYVEjV5i5MHVpv/3PmSWNKctMyQKyviuqX+ivxB7iDN8rGFt
k33+D3lNz8f4QVgffKTgBfiKgOFvjomaElGtHPx8ga+mgplV0dVUFE2VMTalRO2Z
oHNaOIw1YoCYBYXXap2N6+kNcgVgDWYEFvDYECi9aDjUYC/6dC/E3FRLVR4Jbih8
BmhkA+C65j2k3KKQQKKREKfAeXAFwpzm5oef2plkBPI3qlczuwmUiYSS4lZvkVov
5TS88TSDzhYK+0wFfACYaQCDti0+COwWKDdF9Xmw8Hkc98h3SVOJIRXLVv/D4ZOM
/slch0SUGmGooHYe++ZGlHr+MyN84gzrXokk3/S4BlZC8xhJ3ar6lz1yiDOr7cSu
JzQt5VPayhvCHpttCFaO9hJY9pTVNQ4yE21yJLjy091pbvURo78uUW2yHxJiW72J
EVAkR254OVbG4CFPGAbaxjWyLt4WgK5tVX5H8I9kWlB5EgyMU9AXOBIT0IaApqHN
NE2Vozn2FW25Rq1t2ImL97KADJQN0sjMusKgUQ2aiBBB+xwXE8V24ZzPwChbhJ1y
7GW317uC+LdSB+HwgIMULMbXxyIykoY5KOt3nVrnY+iJN2N/10xPBfWO8xgrfTSF
5mlVtQ7PZ1h7Gc+jFyqF7pWnOoWwFA4aQhJpmtP0e1wydAGZ38NQqxoOedcdtPWI
PthX4m5Tbs89lX5a34jRsR3u9vRLAjCKfDg1050fqVXhL0HkpbWFnSDIgTSghNSw
NWKuV9jg4mWf3KNJYjwwEjEr35LCB7Q6F8Yndm0mxd56wYNSV08UfTsvwGeMYpv9
NAxMZwObtDCGD8JVHFIe2u3NIj3vVPl1SFOoctFKTsmAdYzFX/CIOzuT/PPF7T0E
e65uZzxBuEEjnkrlPMrrrw0MGUP8f/F94yGPhnKIc/DZ9adeZWN0P79WFE1p+pRN
Tqz2J1k/zgnfD9lX8vDDDbHca+NneN3j33CD4Cym6tEo2vXUnbMi4k1gr9W+k46/
ZHJN5S9GO9GgENsW74mhUrjXCzLNQdnBOougXS/tcl2Xu1YMKDV75T5kjxv6iaQq
GEd0uUHghEwoXrMNp7qao1l3Xd6wec/jeKr0oVR2maGAQcg9m7Hz33EcKFLfhJ9+
v3MYsjsI6gOWTbHcKv4kiVT5bS9Pi33a586HdSioqN+1LWtQXBpRzsrqu1L6cAEq
sH8HvIPpls/gd+x0V4MonQ+Hh1L9iEW6UgYbYp4KZtUvA+evRQq+r7rMzjQymY4k
eCm9ujp5LXkeyidrhJvPR+yqjHT7PTOQeM9qFHr+KBAQjkMuvq5Zl6YyNItqupI9
rzJVqdTck8b0NtbXTSPKzMbiwvFT8OdzZ7CptknzKFtWe4R6cPUPEZgGlWFBj1f4
YjKJ8eoymN0+sgxVTwrEDk+q6B7vM4t28YS+1CzJXSLZNp8BTVeUBUgpIKuaAlDQ
xGV8hJZcbC9B+FOFjI/5rukUELz9b02rJ4lKNwBHMie0Pmrqbv/krNsZ1zThyq94
xxRQ/5Co3YP7sY3UeuDNGiYchZQEbpjJPTeTBKqpMm7V6k6p+OHr56EAYomf+7Fl
g6kh4e246t0ZsiBYmYTl9RHx6PKfJ+Q6QvRR28deOdtVwj+jJnUGVv/eQD+JWn9n
pgMyOYEwzZU/36h3BZch1aGV9ozfm0gQXxugSwZJ+HXG9jmmTKuydw1wBf4xpoNA
SfKFetuFzg5OzC4OOHmGvOWvahMim6rjFokdJZL8EBCL6mAPbL4G1hsSr4yjoMWp
9oPYo9CiAkZRmxpFavHlAZ+p++OJtX90uw06E7Jx6XlxxuBaXeBR4MGn9I8jAw78
oKUxAwOENlakDt/799wZhd2pZk2ru7Sb+QwcpRjQ1PO9sXAKTgzIewcO9ndzKswa
yI6FYpPyUAMMzy51v28jGvuHiqd8p8Cba6455CMVg445QmyQaeFmnkThVMVlAvAq
mi7gs/7HcAO/RXryn3Rp8cN/BUBckIpzHGJMtGgtSVI7f6Ai0l6RdTOUuCDa7Crx
fN+eGdKFD44SRCjtH6OgEauxBbskq3Nqi6ycTEgsLO6jj/7i4UasBxGCpUjvuPAw
SA7YjjVlnhEMRXwRzXC/eB6CbFfcHoVMYNoKZE/VGm4k9lz8Qoyp2oGhMR+mqAf8
9342gutGDEYBrD7kNiOpT5Lm8bOJJlLbcuk6rEdoX8MV33QbhmyG7eIwLH5ubYZp
rNVpp+V2ZvlHyU3Qk2SquYZ9BNUdZccmRDhPHFpN0IgYQ4ObBdOVUn3JiOPRy4yB
hKG+35xWAwiRT9QcB7YgysB+4ukZsY56yOyaWstJHw3QYNZ6cWnu108ggu7Oaary
zXtc5yPxDRQ8Fnso9rwlIBiKJjBXhdL4iE2CDirhNLb/rTHe4ixwpeGxGsoGH32B
4Zyc1pBtxpoS6AHmlwoJnUJKmt2K7y1gEoxecfDtQZq+Y4UPA2kRpPxBolHZgXaw
kFXqUPn/9tBQylkcgsZdsa9rOcamB6QuqyZ++Sdy7TgYC1qVOO7ATv4wkazdWeOd
Y0s0hIyRSA2xuQ4cc6mOVWUrkfnGG1DWaGrZ89I9n2/rHeYi1mbqFHo7eEOAkQW1
5OI9/Qq2KPcR07s0IaJYsWNMXQhgMaXMqPXQIzJPvqQbkMSxvn80XFdPBQLbhqDN
t4y59JAY7LOSLz4EqQxFiS6Bb/SOhmsj+7vHiBaBBs5xCF6T+pKLF0r0i16G71BQ
/bbaWlZ9RIPm/Af8kqtrCbDDr4o7rdQ8AmWUISDl5IfSWpXuG9Rkf+SETmQ2GaFQ
6vmjx5JIVzHXrvHnk9pwZ8lW07RwM+x+AUCGgoc5GJbGafBM3MZaDhhcBh3amtzY
jaWZFbm8HGdi6mbWe/+2+sevGzBmIuwRqTb0pg55tl2VX7a0H05Co/kIf8WPuAQy
/MzqVxpr/fkTrJdTdA22IT44aqg28bcz7BFdm6hVq0GnyKujX4bV4kgen05hG85n
2Nmjj5Wt03mi7bgwKRLEvZJK3A3dYup/pH2BKlqxVjFQXloj6V/6P0Y44QzYUB/A
wy/yskTTOPlWCG8hVl9DEUqI7jT8tP1A0bn1uROe+vaYN6l49YBnTjpwcjwbh+dW
WyIQkAYnOUPqoJJ3EgBNgqIF7L5aye6xxgMivOD7CTSDwfChfkwxBIIw0G5sDaJI
jjH2JwmkdDcIpuBj28nCNiXSZT9GHMtd6tUrghnHTIYBV6PZGf5gT/tXsiFfP5g0
MzQBxJADUrXJshSZ7FqDz590xpeo/pY0z1nkF/K1V6pvwbDtj98S4m4BwlMUreC+
w48Bl2nJKH24He40aSRXisD9HylFzf42xVxQZesIhCDLyZRYu2BF/rdW2fNKPEp0
VJlWQx5zY2p2pwa/LvVCZVLuYqSqZWuleE9hKL/dfmqxdpSd0FZCBQ/jTtlL1DL9
GPSnUQfyhnyibI5YyMu2Y0uuWfHJRlhHG90b6QtNQ64y19+LtBXoMSImcmxQuJj/
UMbtBjr6h6kW+L5M8D5hs2ktCL3XsZA6pSqCEhpNXON3AEeLSa+8OjDJYPtE/6aM
BMplooytUe4icYVaKLitlanGvx9qoj+g9PNQvE9/r50TjFRNHc7EdKO7+dMrrSoe
FcjFEu53UjrAeFk0cSgMQk+c3mqvwvZR1/g6EUJbB9+eJvmf56BPFoRzop6kYzNb
zskyL0J+QrBLF+j1KTIivjwnT6BwrEQ3KnBr3McpPjz+FFKsDnXpcpq0vZxgyths
X6Mu/rUXBHhtNp8wA6DWV5frk0ctoMY41eX2Gc2VBrFVE9q2j7vmulEwutW5gnxX
lUBUp1PzbIvYJcsqnKN85DyV4HQp50QaWAm+qd9hFqnNZdI3VMfxF6T5vDHY/CRB
hunpzjMfxXijg0EKNPtJPSRYuKJLt9zq9P5F2z5j7/WsqJ9F9Z2OksmFN39i0nU8
Jk9XEcYx3ib/4EeEx0X297y1RSAZ95xVjV0/bxWyB4tsuNrF91rmyqWlaCQwemgh
zD4ZAmUXFjIPydCMTGfijXpdN+z+sCnVzpLkEvfEAV1q0I8xAMwiztHPr0XPMAP/
fTIKduY/Pt6HK79eRpa73+QlCLD0jMih6kDBHHZ1cmi/GlYMYkVjkWNyk6q6GeMs
0Axcni+tuqmDdkpLWTe3N2Ph++gpdHyTD/YlhuOzUB2+hxxzuqFoIQXbPPA60V8D
afBBrT3utvdxv2RpnZsmUIZ4iJ3jhO1mVfD6ZsOGzHycL2nwoudWY3m+SRaS9imc
qQatistSCy8hZC4bHM0i3A6Pd3JsPfo/fBYuxf3quHai75QZjqA28Ao8ZmmKOj1A
Fr+gDM6QCVnBFepN4Dvumh+TfZqia8Wpf4RHpLhYvkNGrrmIOAOR4B4dvgvf+qYF
EKMwS6mYaYHeecdIt5ltmSxYZnhPjs0bt/YrEERQbwQkkZK607Rwobicj2HZ3VPP
YJaAmVIEl0jm7d3b1ms601YxKkzO7MRxbpyWnkRYH18GdtD73pcO5K/dKcYCNjKU
wUCbAimlLJEAaI+7u6cyIFi8t0VcFVftpIaBGXGSdYkw+tDFSvu4G4AgMXRzcXss
HMqRnLhgZW5PJmO5S8Lb2jEBTPRrWV+U+tddu/axRQsDEGG0ZEJHzUlXF/HmazC8
UgZdPlFphChN/ymSHMmlyCHkj+TddgdsSjQy9/Okbim0LGXOmphxhJClgHGu0QNd
MEkczNLFnE/uDoqMkKI1qm1dQAZiEumaiHp9pWrjsg6X8QHDE5+qWCb/PWTprHXj
0ywU1z28G7CQX4xbar6HNggHvn09OgAB+q9sPeLItR9oDY5lJmDdEKKeqng5EA62
5lVnfd3w+B+6HVgO5T3mF3+qBCMCiFSC75vsM6xSJ2sjSJB95YECYbikAvk5569k
/G5fN8M/NH4m1Mc48kLgJ8SjRXowSgTs9kiKi56XFytrcQSQzHiPrqBKmzkr67cp
UUh1OsXjlvlmOfGUAjIc9wVmPNCPzsh60Ws/MlQdIk7Ffa2h3X8aKnl2kXa7vmwc
Tx8t1ijWY5aejR6SJQNBfN4ExuelBenbTbjhZgqvATkKSKRN7cSA4CxVwob70uqo
PMtrwGs44r1wdcgIzx4kyrDSeRiUwbdBDfL/myzquKXkSA955g0BwC+G3a39XSJr
7iqiO0ZG7pev5d37/WH7U67sWJ3sH9KuoBAoKY0dhgNg/+HAxFVMQtHHdpupZ4hq
xXJAz3uRRFOsetyrx/+Rn0ZDOuKpbCQg/Yz7YMqPvNZsjMil4GQKac9bAMNtu2eF
AtNh4SwUK7VkQ8ts90ia37tZjsj2YZlTLqwbubqXYYJgskDDw5HH/FtBaEDjMKR1
vf9OlWsWOP7qvi0do0gnE9iYG7jNR0Q3v5PFVuol+/dQc+BjaD/B0PVwg4X1WQoL
sNLthEbiINAHrQ+wJo45YVgLEnftnvv8LdrHep0673OfdqTqmW+odUrQb+Zb5xyd
Uw+rh1t2Z0ADOU3WQt0mA7HLTWVMvYCE5jdMFjaHwtMsuFhayMX3TW+bSEbPeRmm
LdKMlrgWHXqz2ux1oQNNwtVdy1ZOzMRvWeaO3EZB/PxQuHYFMDx2HAip5CRfsr3k
HskjmhZniBIwLRELi+dTP77VNkWYlbEXk01nK8AqaO7o8aLjGARSats99eRDVZDS
btqzaGDczNTwKJWI/LiuRSOakxCu0wj2tAIZiNF1GEW0ut4BlnDr0dNN7B7jeRSt
AqxSRzratBkohicFK0D+In+CN6xKybghP7knaMMEACtl66HQDO2QdSKg3nxZ7enN
e9rs1EMCRzgcdABxq9f3aH0QRLupP9p+ZKEbI8OJCWXnR5AWApHixWmr1Op/PDtI
K+c1gCZro5Z/MZGS9ALtmCQO5/Jt9tva2g56XHNP/vEu4+SGZddz5TxYgT9dGDCR
Q1wAHWD02aetdlYWELcLpna8jc5KGoeJh8GPT9Tc2/whdXehociqGJnfZFf6dqLs
2vaG6jcZPI4xxp3mOzvNY4neENGbWhaBPXRwrlJJJA3JRf7UHlmpZiM9DMIWT4tm
e+u0pnFaYbMv9CJKN69ZSrN5ocBDkmXiF6DtuDHBK8G1Q+ZFnHUJgaKmT+iboSsL
ZpkKYyiyXNLiMj/N4ia01QoQLOHA7igza5hfuoe5XQwxgRLpPbj2sGeMcKjDP7v0
Y64h/EyeY2OzuQL4TNVBf1toX9JFwu43g4c9S3ZD3Wq0rAH+vCtkheiqxqiqVmKV
L2JiGo48QdmeCJ/z1o/wlJOD9RkU2jDSwZAK/ZuA0eXVWgTZx3R03FhAY+ZVG9Ii
xvGpJqN6zOUUWg+L6kv1GBoPza3FWXV4n6eWrhpBPWdcxT8cn7E1YcYzClDTPP9s
bKdF8DD3zpiDdeZ+GvHhtUT1h/Zo+KII3s5WiaYxxAP2PHtaoRLhqq12Rbm4Oozp
5ZrRlB+Z1uJ/284GxkP+SyQuCe1ORirWFMmJGpKWw1/lmV57a22g1oLYZFL/rt2X
1ZbRXI2r1uRUUMCAIHlKGMasTODqOweLNsnQ6fP5VOILgUpK488zuywyc9EvqLfD
LJyXZ1aDtpDvsSntYsl2mUHNjfOS4DwXKAcLFJXRaVf+vnMDJN01uOi67l2VMMXH
d1ievgtBAlMY1pD4nPRxn4Rwk66VKU2pl4G/GOHuiAn7eD5M9/s5x8p44v3i/RwB
R1VwwUOzKcdqcxSqjoPTEGUP9kMvvjE0wI4meRKLjRgKNPVZpy1AnP6Mj7O5W9R8
Hm8FIMkvf8N9r1AqtzXkHLDQcYjQs18VMFNz2y7BYFfL3TS7GqxETeR0srko9Zo0
oBh021kOvDfZk8oFrj5HNBZNPFM9GS659Hb68RSSjKHH6CHpeM5q60Losk55W4lH
S/S5PZxAuZEC8273n85dKgutEh8gSQl2xn6+N5ZaKn3mWbWB1UqIrOFwGncYAMoc
MArULARDKq+7WWym4mwiVEyxH9IEYPuEn4gDwPD/mYLP6Sp8evwAlcsfHlw2Z0Jl
E8azcPZ/PlF+/+WEOIgPP8Jp3ZY1FQwaAVIUJ/VFu+hVHPiwVW0ObF00DQxj/9uk
578h3IeNs5W5+TaicyrPQmR1E+91DTDXni1gt6piCKJChgoLzdDIyOX88Lmv6h1m
ZjBPde/1GiP0DatglgaXycBBnB58j6lprwjujV2jQZ1sRLqsJHnaHZmKPlMjpaPN
okDREpttsYKZHxO2008Ml4taBhNWd6cexeRU4nNbaumRy0Yl144GuZUNyBgIKCbx
+xekxX6Sn2M9oO1LUlinUxSygGLoc0W4meGP2KLDDoYdAfH3eKgVgWO86hyItP9G
vERm+t5o3oItNyKsfm5FkJoAdyaFbtagYcpZbUxyX0gXcSRS7qYsQK6b1usxQjPe
XjaGyDF13WqkJmxDqb8govxQCS0Aixb3TVu+6JFG4u9ehBnsys86cipOGK51zaTX
zlHUyArD7GHO/IiX5NAu6NDIU+6omqidwK8YtHJtQV90n7C+D1v3Y8M7Fy4yWty5
iUZMJ17Z/7RZ9VVz+6RMdnhcGt7+miaEadpaMekQ1eX5KR0mYJns2IzooXrcX/xi
wv7XFsNWY4brqLfjtrQblW4luxTb6+YFpY6KjISUQ0siMX30XoHWUCqvzqKUqSz1
vS+UVrwTc/ormm/oJJE/rGoVB3kT6LEcsOYMcnD1ag6FfPpF1N3V1zLgHkmI6BGz
YC/CGnuNFdsiaKlIyRN9XXb6Brg53KGl12JZ+nt3z6IkFuR19Pg/ATn08RdV+uBy
vqiBzJ8ovFgthbFKAzeLLN7K9pxtSj30ibmXILUy+/W0uBcTtTZqt7xHmkmOtAOR
DsTTDVOqZmvwSoL/ONdgE6d2z6GWT2viGfCyGBLwmt+Y7DisAoAZvTJWqfCKbzGw
DgyzHmP32mzXOxDDXbENwOkojQZkbxgxsnAyukE35/4nuZfE5z3OqjmiSxJyDU8k
tR76h2wZSdW0JiaPB68EXz+1cVd4w5rDqbNoSJxAPosjHc/Q2exCmycgxbIoGs0J
eEf8EZTdGS/+8dMnQIthA/nEMP2MDR3G2B2Dqt6fvH7AjBUBv+GR5mtfozn4Eeh6
BsUaMFrsigccLDXwXwwWPCHGJKIR6ZKNqq/bfFHhe1nvaQBHnwPw/RJJ9UlQXnVc
36gavFJAiBCmGqIIpRTMfap6iJepXBSGF1TJzeBzIE9404HyQBfIDARRG25DHTRu
F6uQeu/Mw17CiKkixC4mq8ckEJgqxkVSttEivLJJ5ejVnRasaJsfEjosoKnAYwv0
97x/FVSxA03hJoWVR7w4WTqW3fD7i3SRRqzb6iS+nvWriWcbitAQ9u/Jjql/tGej
AfKvL3ujpt3EeovRJvwQ1yAbe9Wha+bFvbdympJMxt6RnHsej/KK7700ugnW5Uh6
vpqJOF70/vmYPwQaaE6kak1h9NJjWmwKF0d3PmnoiHaXJszCIUCrBhHdijGXAax8
OKoVe240IEKkWQLU4vgHJr0PIawNgHwL4idQ0QMwFxtLee2FI2ip7eZ0JKUgk7iG
UhjJuHBX8EbeCyK16vLe4164RqsZbR++7h1/SFaKF2g3tL1RzDmf6hmXGIEQLPCo
7XVYvgKY7WC+rOLVPnrkZXPCdUcwEyI0/cflt/CTwPW6KkWPuEcaniz4sRf6D0wV
CWvvei3aQQLMzc/p9W1cYl6Z/P9l1PdIu7OYNSqPZ17Vhn6+mAmw7HDzBC1SYBTK
21nXYmmn8EqFtn9DpuJTsRWBtN/loke1JDoz6hvls6YMsB/I/qmzNBPM7tdFKQcB
1jmsvTF2ZcuBKxIjMCUQo44rllB5zO+DLvQmPcmvkAtkXUI7vRKapLTAneZc2HXi
yJftGFNLVLAScZP8CHhdIf/70nqlPKv+Mdm2P4ayHGrFyry07ZvdkB7k335+nNlW
zngrPcIKcJzmAko6yinvhC1YcEbjbYmAX6q9U2U2cSV2Xe0ePlSJAQaZa5czOAy8
fEpglZtTOtPT8X03brDbAeaxR//I4loUPUKtGLWN9mqCUpcWEkPuxTsZBGe555Xj
aUtnOLTBFyg1/vqgU1yQmAsaGic8T6/tvWEJW45mYFxHAnjA1XcypcnYYZ54Uppj
rkKl7+M8JwB6CdeSytOiSB4gmBFMWsYF/7NMMM9Nxv2mgrfbrIoQ7SijIECLkLrv
sBvePzMoG8TttTNTgNAbS3lH+1lwu+rt2HFxUykaGod5My4Fuc0FtEMoE43dZthM
r9EZn1IjzjSUhvpaaD6TZe4ZgcU6ApFIC4buMvAAvdjPqLWBVIbQyOKNiQ92rHwf
KDXIFmaxwOQTu+EBl17ye647dCfq9bVO0KR2AzK9QvjbPH4JDtlQlmeQRAqRRlUw
kEYvT5nGAiCFIHzC+N2VqHabR57OQnkA5h7Uvo2OWVxBaorX4vtiP/yakBkjWE+r
Cupqkc1+kzVDjArYdN+OwYhaZGj5+hx/GaHKFHo3WnKl8Lw7e4F+RuY6ThRf/ocX
nDHUi4vnDwSjOlDrFfSCfGvLOWXY9rWaJvxhj3vELkV6eQ4yHyNoXOlMFxyfUKoB
uWhivJgBvbA2AvYua5+DIQIKhOV/OGfktKg32baVgxycP5cOsf1NOAMca1V5XMWj
r3qE1YE7pxpzWbtt1Rp9DmAwBHBPwdyuGQTEvVF0IfULLuzDITfBnNu1gO4hxS4W
FbFC0xBWw4ryGcwtIzB4dMVAfF0NiursbmqMUEb/qVvfItE6rQZFOGQ30xJwm/cK
qW2/gaf9TqHOvYpGsjjbnYHp3YPNUeQfdjGfCs1PuIYusy6/9jQ2EZpN5MjNJtG/
8J+KbEP/Wgi+qpr9YkDAw5y2DKTnaztBU2pmKH8xZdSjpaYjNYCIOVXBNAHeU/3z
WHV9jnkxfkq/DLkhjCLGP3eXYIhmsBhve/R80seX2ntF8qKt8tKoltViCvbOoLJR
/CoqCmUlSx8DbpqfUpq5SHhM5gAhksHYrTOj1dow7YJ5SVjVIJfCKcBoS63GCjqZ
jzbWDvJs+J1loR2tU7VH4ytDDjYT0S/Ea7Unf0O/I4tgOI33kFlqjqr1f9PGuZs0
3TWihL5bLwhCf9vWgtsjkp+Ng/tZEiNLVeTfafa4bKyfDfmcLKZwTshfMP4CeMZ9
6srU7tJi+u+UJ1SP4z2V+6vmGDlpsBJkL2S/ebZ/spYVMp6DgU4ZFgimrWFW+mUd
iW7fnSeqmhKtEMj+BLTLG2j68O+41Y+Fe1uKRAAyj5vYCm2j86aJ4xUXBJi6DyTD
0Qh0VqDFVjJOV7cEeCA8bN4GGh1PJaWJf8msqB8+lKSKk/KVhALTpuBXxIx4PtsC
Zf28vz6+R/iMUkjHeQUiVnl2ibN+ynWCx6J3wCsDTm82oqE6XHSD72T3N04wEMRh
WJcMIsOp23bk9a0RfGbxE+DzrtjH11BlluR2jPw8HK2pCST9QNRhE6rRDGmwQsgJ
T+2hwB9W3HLPIL03ijVO2VpwSdd2ElA7DlLsuJpwUfcNkhhFW2Y43d5/ROxtGvHa
4Bk/Yd+q+dmKf4O7EzSA6AKrw1CFMS64sc9OPx0DqD7IGn/fawHKlj1Wqu3nKshb
WttGugU1jlr7tZx5ehhECI0+I490K16OezUcw1aNgdk47HGo7U9Qt0U15tNh8N7a
9nCXvQnqwWommR92pLD+06aFBXvMPOMlK5jjYhz4v6vqLcGLliniE/DDYHBDGK9j
soj2G2YDPFVP2pxXCWpRyLK22BdyFkSJ5oHlZi6Ci+T7SyoSHai/QyWsmxndF+Ek
K/54eOFpHS7u2FLCY8a0+bpOghoOH1HXITwBwJmKfKkpn9HpzfVL6Pb/bSFm9yAi
ZqNSurj9adkS0GnvWPSqDBdUVyRfAA6RnG/Ccp/Db9OI2Zu2wB1BNCKVPHOBYRM+
iqiX734bU8E0WdleKYsHqbk3vlJpbgo/AnYXMmG5N+AzUbN3aN+MpLsoRCBFydV/
RwovmyxeSNZfWPIDILnJWvE7ATC+hHjnJ2JyST9GvL+hpmyjVBLRg2oMziW9yJod
40DfdXaJ5DSkI4JGPifVZ4TwzWIlM30K5yq1R+KqKOjMYzZGKzYHpvuLiYKGwda0
QTzysv5NgIRgMD7Jeg+1tn1n40qOYwBWKwLs2c4v9F+fZZnVaneVEBKaCRYc/DBO
v9nEUTWi3+nJkFdz5KePNZoB4uZS/Is0K3McMlFmbGdcm3DneIlp8824+i6oYurM
csr5UmbU7nh32dmSAwVBSzegfckzNlwJxqgShpu4okccUbkdkgC5Ub0nAtZmTQlL
/2SbA2bzyguBEi8QiaaSiLSxCZXhF7byrL9w3XrzV48+QlVfhZ7kF3MqvNf1DNBe
w/UCzSrfzR/T1NH64XXcNEMBSW4YyOZKJMw/itfSpmTs2rcvz7rh2zeB5hr82ni9
i5c+y5OSPWFxjdVR0NUWbbisSiFCuBsuIjP/vWINZnZ9IW5RjPwscfUflvNAAVkM
PspwISTUdlTYxHdyMQdjPonc2XfYYis/GyRWgY2fUHrfwM5UQmLiiuxXIT82cMmL
ZBAOiHaYeF9gGwYXJb1T7+dtodSkMGn+8LA5v9qNjg/i0wzBHjPqZureMrW6XYbi
kjaVekg+Ehzqv+qVwT8D0U1qrIONKa/jGtKThj+SJEKPZavvlnjF2i8k/67US44y
/v1fyj5KhNeLtjouFzUnkCZkyjif3JgP6j9q9NE13A7u0ZOnzabmbfAEkce6jXq9
Gty0OEbWbPdKwXBa2+pEOC4hbevfrJFwVbVreRhyqonNTPhV64lvq4F/006BvpBd
gPYG30Fu2Rks0dmcBaEnAnjUL4AtjdkR+FUD/c9BupDjQwVwAiHlmVLBp8JAp2ZX
I7T/fkiPfRy1I0LdO8HeXhC6kWlRLayZIbEX51fMTC1Eq3KJ3NNe8zKlclbc4QAy
gX/7CtovvB2KhAoj3cy6mllR1nOxhSKY5he080gmdKVfIpqNGeI5f6ogsoxk/13p
FEqPoxiFpI5JLzi+N0FJ9VTSLfIkCM+nsf/bnioMwHNpzTserudz38nuYpPMxOhC
cjMh2dzVYR0dbTU9/yKYNPPUe8xg13AnNXnqgXzlNn/d0YuINSBQx4Tl0i1jDz/G
lnfmfB6IajFT3f7TVd8NYAYDWcM47hCmTkO7XjVFalL91jKh2nezAZZWQZeoKmdS
b7n4UteqrxjCi71vtxzXgeAM8QLoQCCKqWTUxoYTvTr/wF9FO2PahHrL16RNdLso
chI7f+Jzlw0VTx8uEpGj9vlByrEZ9sUzuOS8yiPxtUZLBLVM6bD4Gzxx1LmVHnPx
PhEzzWMbbmwp5ZUHUtmkTjSHL1O8GrYo/0dwn1BE3ZHX5jrP3xII5oZdMTQ2ldzg
/KWnWASM5HiPf5pbo/oPm3CTxFYm65plnDgCbKKrZvILooSbSWHrKyeVEMm3GN5I
JbXk1ujWPnjDztBzO3cs5wneT5FMTuNtJdI3ZWjWHKdaSQqQageDdzS1nLxUidgl
og4UVSUUbLyy9CSz09DcrLJOVqn1XC/dG/QGoYQmfuWE4aXTwwk9k2w4pB8yrLLC
tNtWLQHgcorbhEkxJvHkZr0k8Rrw0d8g1tT+qS2li7DcQin4l34/SZsuQVaYMTbU
tCwP3MdMQXvZ8Aex6O82iTOR32mrMQq4J76fu95GDx4ObZ2eIovSFYNNMXzjkCHv
7JWC24/Apve8buqr3dVblj7ZTfm3XSAxoJo3NgA7fRphwLNQoQD+JYC2NKexelcs
9j8cHTMKJSV8Mh5EUBFvLr+elTafU5/ag7IeefOrjldBPEthfJ4CuR//ph+H/eTQ
Fv9tIIXq1XuSZtlvCW3LCkh4GT0ZxYPkGiYdJfoqOSGth41kh5N59ZH5vt/nl0T2
68OYuVR6fqzOt3yk7e2Rcnpfre0va7z5Ig2QrcWF2rnpu0r0KuViV/+x6lYG+Cwc
5BPsYS++ZvQms/STPRjTlbkrAn/yHDyrcph8bzOdHfyGTmNg1QzOD5UqDwCtGUTq
ny1QiP/Js8I849Agv1Qgb1I35c9Lw82Ecgutk5r7MdVAIo8OIdUNX53NXndwwZTa
iMpb3NQ9bSG+KCjPma3oCe2bpUJM2woC6cHr7C52PQQUHwSMD+UBTXsyVCTMnxE9
Ad1ixHNkzuOZ2RNoplV3OOTvD0Jsc1SN4JkedMvZ46azBK5zKQCLkLzx0l+tWsq8
lMLes2FT4WT1O4tiN9wOaa35+HmLKLW3APzcwq0kb+KTwo9Zm5LUCUQI9KnygT91
qAX1hOmjSYKKkELKgs1zP1/cGgJLuTHiW/pvWZG3Cs+HjGHIMg9Ns1u1Z7hC7zMi
KIcwM1LHSt9GU30ScK6KCgUqBvhtLm3Xbada39/7xAvNunHMtZT/wp/oT+Xiiiq+
tPDniRHapoLXnya89OYsKOsgMn9ZuhQNnQMEyO/Tv86uZrsp7H5zk8ynPyLUV3dC
KTVZW/hXylDqsEn+rqxSTyJEZJosYmYgHhXMiBH5le1J0f5ESrXXbk3IlLzG0hgN
7FKhKKnC/L/hb+0jEsS23xe7aBKTTZ+DGwGNR6UaBCBOXpCCXMq8UWs5LT5S0zkR
t5bN2dhCBvQ0yyl1iApptNdHWipElLBhOe66s3epRaeJfTwopWZJDoRv4gI6ix+j
kJgIfXpHUKAQprW0UcqLOgJxt3QbF1Ek2qmJqfx8J/M6Vuh8WCmVNTkjPpOjL7is
2sHAQ4cXAWa6uDwGtaheSTDGQ0XBYcJY3a+Yy8tuQ7CxJS9ebnHHHcDjnkl8vGLP
wjD+k1zLdoNSgqVfH487hWzjwD3dg2N3sVDqMbyFZ1gX6yb4mikXklPKaP2rwqVI
H5Sga76GTRXFJPtLFpg2J82NDPi2fLRw6cFmm1eimGb3GudKGvUKePkh6E0JjpYO
Q791iC2X+F/aU5UUoCLS2SXkAwtw7VZKBh+p7gr6R9wvP2XCIFd9O0oVDBmVSY4j
T1zDUAxSTxBj3ImhO4uM6xI3/5G2/U23rs5rUuOH5tAcL3MQPl1V//kVPZ3J8gPz
/BRyaxHueM7cqWJRWDfMpEx/YWztzXLGvlccLWomfZQRA9kYroMnz7ERU7VfH8Tf
qseZwXpxXFkqk0mbcVKHeICfKWL2cDnnNcBYubsmGVtIIWO3xPM+vvBHgKYIfghH
YPNsJAPc71oEOlX6//t0omDsWG48r/8pFidgx+cazycPyhFOpikgdeB573u2zuEh
LyoyURn1WbmhSHd/UL/Mi1Y9MCn+BuuRCTaI3U9UbOrRY4ZsgIOzfmFw0pL5RYxK
d3Q+dOOCenU4WTR0R5F8qdJ8eY+KrHVeHpiQQSipiRFdsMZduqbJ6N6MZCC8GOkA
0ZMVkfjXP2jcE9seP26A0HAvuI0INttOl99+Tg1CxuGTOSHb9l1qt8aEp/NGEwaf
dZ37COPtlfNsl7Ur4SMPxLpHAx1xQA3Nqu42jFXtne7pwS6zjd0TZoZlz4hJepyv
P0n/tC95qDA32iBlyGf0XmIAhXA899VOz4j8Sx1r2CqrdULWbsaIjwXcGmGjnVj8
JWaBQJOmHG28dcN+x//rcUUpY8xleCD3rZXP0COON21WKFKw1lDdkyPtMgluQnaN
jwH/vd9EAv+tNhXKVwMXIvTOt/cssZxaRz4kKx31xw7ua/O3O2zW+nNQCdUYHijl
hwXPnBbJ07N3/J6M7N+ztc/s0f3V227HAsnXQviULJKzzh1Ixwm1FLd8jRMinYZR
qeoaT3f3Z0NYChChg0kbiXQ5oLw41oi06HQ7vW7Pgt04789OHt6mVyttxKUsGeh5
xFmhauRg3hTK44U68aRxBcGJHY31AVTewmpBU3EJwrX9U/U6b9luxXn2XX7gAKs9
E+vcIjiFIvKTdlpjgOiWV6aYyCQZAUvh85O/5Yl6uKmTY4gAqU8ofMTGoj/gGywl
qCTKg+RH14bJzYKgJHI2QJ8X1Y9W7Ak7Yv4PvyYRHBwWHVMi1T0f2pRc1g6YMNJs
cMVLzopU3zRYEYqb8wyAliUWclRCCHkfE7eysInjvoM3nldmTXO7lLWz9ggYW5rw
VgnUaseG229408sc9LlIFVK0EATjWVwkP6LxNByyTVNWc2VAQDGPlaTTeeavbG3q
ZwiD4HOtpGlUWmrsV8BxohNVXlQA4mXC8YzS9Jf1cqrNjOLzMUpxNWjIUzkoC6PX
3rXgSPVaPLYxmHOpcK1WH4BoZoacjzJuIkqpbaziyEJ+wqKkRlAYRGMx77vrNCWX
5lPsCddoqDVP6BTO3+rxyp82QUl/8pXe4P02tjjSq+YT0vdgeJs23lctPPxLzuEh
FxD9RIlTaVkE3/QCZqGcI5hkvAd5iecHE5xE+4jNLDPSj1aiixqztcJFXK/Teuvf
r0qJJBFKeCNuRkTIkENyWRmE5LQDoCZqwPXu3/DZUrcqQc71b7jRY2QJS9xMFfR7
ZUGKQmpJznn7FWGbuesIs5GsdNLiExgyA1o0UgRJXmy4yV5e+7IrAYbyfStVs3sp
9anpgg/8btn6JGOJeh+QjpabUkUHIiHe0VXoyN8b7lrdPHQPZx2jHRVvoXdQ+N5E
75cekuWAZpAomCVeXc4dQRESErYsT2IynhaK/x2BUht8scPHsESp6S/8Fp91QzUG
L1BNRTvEiz69W2Ak2Xjm7W6PjTGZb6saDpIUfYhb4h700/k8C/sHVXG8/NSbTWjl
7EDcJpDL19yIeeIr/UHLCd/SZlsN+JnrAlArc5xke8iLUHIoulT/AbL9sPt70EdW
IAr7O508GcjP4+iKiDNk3Z3Gc0y/q4DbSN9uM7Ispa0I2MkztoNZPXdT3OoCLiw9
GoRerrFZKNZ1++yP2f/uHkd33YByBVvXVVoIDd8IOx8ljbuQ4S/STxlHub3gEQcz
ouDmX0TLDQ/+nMtGokhdDRbPZHo9LHwZQfZpplfPTh8RxksYUH7gI8FOOlKi/CGy
fxF7mcigs1KoLS+1aXvEAm9c8MHwyolYBWRCZ/uDAsiouGm0d+anqmjh5/zO8cii
69BkxNIXEF9+aePnPO28OINEFqD8ruYdULZELtTnFdlLi3+8NkgF65tVb43PqEvs
Kp7qnanbDBPnu2nS7S/MolENAOCTiHokmlY+Hx6/c3e2Qy8EVDsTE7WuLvlK/HwS
64p7oKAR7q8XLrLrP8q4L8xKEWsCjuaADAFSI5yEzZnDXhfdPUOsruKsAdFS3GnX
g5PPvY0fw4nY+zSOCLXkVQFw6OH0UHXaBw8vyT2LbWSEzLhJYIN4A9KDrDvyZTY4
PAmst1jwmshNenrd//FVPqJgL+d213okkBSx/Vdz9YjKoVbRoB1y3osRsoyjf/h8
vYrtipw3hl6sQsc/g2cXIp/P2UFu9onVatGpVd6B2TBJPvFdq+29MEiPqNSXT6VJ
gHW62V8yEAh24K3enqf/IatJFCzdt2TCnONlBhQl7CGwB2nrL1uTbkjCT/9GU7UZ
KcKiuTXmPhAyhikX5v7NbisCmriIpHBb90O+Iny/Et2yLzMRC+iAt66fIs1KHGdF
YqgE6XAbvJtofqpBBo8o18sIntMm+f5GMebASbaH9sbwggSmOwHIw9qF09oPslae
t2xd2CLmpI/Rptqtftrt3Z6o/FSZvRz12boz+KRrxFBxqtDrq3XQQfkj2R/LVcpb
Qqy1s3Yr9ZErzhTLFcoWbPynDDj2locck6RiY+HUce188x94PpPctfKajJYyYDd5
6m52GnJIXufQZ2FmXHVFciCxdCzeuBdIusilIJOIikNxHgv/erAfXr+KKq4bRY5R
3REFnJfB6vkdkObjR0Go9s+7/qQYx/IVutRtsedk/FQRtFkzX/+dl6uuGfR6R8CU
M0/FmgYn/pQePlp3lGFtrz9UWXWislE9ijSln/zOMuHxP/ALS6KAcr2zG/b/aonY
F54164wWcd+LyK7Rl8awBIdQrCRKh6WUIb4ws1DZzkAJvwGfv9OqQ6dWo1L5GYca
9DWJUwCNogyGPeEh5/4SmhxdVop+PWQ0361JR9pWgcmOVRu4L3CxRtvwR0nupf+W
3GM7Ieggq+xADoDRRPORPr7tuPV3oNOYYrYI/6BbMIkoDe5j1KQKxvU4MgblIlg2
SqQTKZHuvchdnhbVuxleD/Fsq0U+YqeYamOaxmO8u/Fa9wRnbZxBYT9FWQrh7y9l
OUw6EmGcF4XWmgZXq1Zms99CERJAWQuZZug2wn2bR99wmUnRYiB74Y+iEjHRniRh
K84smsZInj4FcVpApUAWMya9O2R1i2SDvQMQ6xSJw1saI6StXRvtokUn75mdFPv0
/t6OpRa6H8vrwqrSN8T2vQb6wCd0qzyCgzpPf5OvGfCb+sloxeATVFHXyWhQ3iMG
k6yYldIFGOSZWxeMbCaf9Xul0eTqrcFB7XbVPOpInM6mfhvo27KNNYYocIVu7x2F
7S+TNBk4cocLJVTwnC1ZaHgFYsZBdOcFhI5wBcoC1tAnxi2Yb59ngUyelQBko59N
BKiRqwKyrMieDFteXNUcExadDrWtWBuxGLxbyW6N2g6fY5pxDZCjzrrDuoQ7STgN
0KmcRNsbJSINbpzLLWIw+HWdLoTZffx9oUJ4Nbe4ChVlpQvKqKNOCKL4QEHeWFvH
79D46C8BilgdFX7lTfpaLcicRAiwo/KNGUEzxd95FUq0soI3jGe805OXnIHJLYD+
hyxMasmBKsynaZXfXPG9nHU+WijfcfSk0HLwwMvC0M/3LcaBiDI9gTnDPGq054HR
PzR0NJRZ3yzKlT8Vp8D6epX+YOGRVT4JoBYeP3lRuf2T5wsVYDVSNHGKqg0D3i1+
KZgQwgo68W4TdSoh2EzHcgBtslGl5YW8sSf4I7n9/EVwwcor2vZB+sJrMqhvaZuA
VNGZWWJZNOMq+UGKso8LUAP0OHsxHd2TonCLwukDjtT4J5OgvmCD4grkQjtSXSC/
Ghwoabv7W8ecJ/v3RF2f6ZujTNX9iaLYVUTGz03+uAUkcI2WRcRKW3CjtyUQf7Rt
oQGSu0Q5i/6BcNmevWMKAJzlKH4aY6BBpjVCxqaLI6zN0smcQour1jYTuy+u8+r5
Z2Eref1h2o+stMFJIzJojgpk2NatSRrHEr/btdFJPM4piEZXu6WdCOELu0EcHCOH
xpN58M8zu3inlbLxB9jb0KiNTUzZeMADA6nFYrNYIrrRNSoWNvV9nJN8zbG5kmmZ
w8SJ50zaSWKWe8lNAcss3g418Y5CbJ0JrzqAABRK+kdqBkl+d4ZUSEZPLtd2vA7j
CvziJSOTbMl34JUyLLt0V9PXhl6Mro4FgTpwg7rp2vAESIRW3Nog1busoFCDXI0Q
eHx2eNF83qJo2Rmvsx97DptXrhDmMnMh7t7t02w7wmohqDDUhrigp3CRb5zfBbFz
y5AtuwVCrhjdh1fma7Kuef47DrCToVsQqj54UcK4fDia/70C7jDsvIDo91poWi5Z
hfkjvYXCURce7kG5YUkcYvTB+aTjLIzMfOgTNQ0edBCzr19GCvM/lq9OeESmOfoW
GOwRmKdShLkQFdjSNtKjj29oZgf0uV4kKjjt6WyN8Wzq/tvyRYTKLDHaGoHR4vtA
eLZGmkfbBjglHvj0YEDyYHFBS8fyVJHVIsQp58wrY/JUU162JZafqNnfw6gwGhOi
HAeFopUzUFtMjHSlEPjpylK+iObmNdVhIrE5pP0dlgOgbySSe8R0DNnX7zhGL9hS
o1T7+PvepNlAQpaQk271RE6n88ysAO0oWZLyUidy/2kqVR1rc6CgusI1KFRG/tEV
V37YCnHGIswInvXadKfouseHkO7sqD8b9pYeyiZpREhCxFM5/+WPgjPora1VCkK1
Q6IRfWLCXUA7erMIsmiQ/MeK7qGaAfOAvo6ruvWpbBc83kovnmRJayQOCRt+FFBa
31wXvk1Y8RLWG4ghni0eXOXWQQ2Zu115KQPbIwbF3ehHKjBi4HU1afXldNIYNc6k
fFlJ5Q616DSD+7OjoSBcpBaeG+ZZ9kuRv2iT51dzsVOQ6+aT3U9xxQ4FAZwqNzrQ
o/KFF7mMGhhU/yHcM05+vSqt9NjxLXBVU32mCI6eSFh40PRAq0Z3A8aurR1U8UGa
FbXbLJUZjA7xcGVeiApcFizSRBP9q0wCnPX9ucDWqr2dPI5WURxuBzkCtRGT/N8K
hQ1qmTFcZeC6TXgzXp3hqeRsC99g17bplae8H/s6WgKdk7YxTMe8PM9swOweUTqH
48MKl8JcZMhUpoZ7Et6lqJYPyORPaea/CsPsstqHVE3Bg6l4HfmDfzyZFwZWM4le
gRCOlFWSSm1hu5DUZA8Ku6BaJtysP4Hk0XlBz5IRw+trsqI+e0UBYLThvoPar63Z
Rm6UnLGWBs+nW7QLjZbYIyNkAdnBYG4uk/ncsmM7ySw5WosHLBtga6JfWNXKOadh
KfUDW5KWoa44Tm2Q3LSomsCofHp8ZTd2JUPKuTJGO/zQTJcn0aLBy9yX0xG8ubcN
s1mDaW/uRECFBmgHCqihl63oooK/X7HdwPQkEeyLeej8kqikSDi57bynocd4J1cS
MnQw25FCxtjPa+GOJUdEWSlxq3ZG2qNchEvNaY0F0sqf/YwX3LT1NJrK9U3A0Wfv
vYqaF2xD7Rc6faXU6cG/BIRZ0BJXY/WtaRjaB8dgs5IY3QQIiLxuw2NADDHz8TJS
05cHMhXsYBhExDbXmti54pQqgL8JV3aHoZiKczBMT4WjiBlNTsDvsMedckmcRbn2
/fGa4xEpk5/tnnwdDsLLJooMGoBZBZ5ih8mKJjThXbfwjZG84Vk2Jfg4khHhTJ1G
fJITNWPcbzXEZrHyWcluwTw7gvwnDtcYDrfBTlecligwlGOlxVYMbyDtUSVqHOFU
/MhTh4ZaC5H6C/wO9zjZWGHG0lt4Ton36M2efQWMOj27qwFP/nfNi0DDaPPu7bYO
4bcfxmfFN4hQns2qTFuxhZ9e5LS+uNOg8ft5g5ZelAmrOwjVTcAlPRL0Df2LmoTN
MHo2mBRlMYVuMg5bVz0iyhQRbPQAy2D/pKdze/cLRjAq1tCeqRVM1fVN9zXh2SIb
LlweEpsumbZ1ald0ltiOC9MXwHCdBqWo9Ul+tbnqknbHvd+Sgr/lkWz8vG0WvhRl
mnxhbcXBXkRqcyeZ7b04I1r+/JRXW1Ntbz1mUPsmEhiKwhB3xbLndqBmUd+wPJzW
AdiO3hxNxhUhDAEDPXIjcwEatyGlaXQkzoDaCkKQN5el1pQ0nu/TXlZd/rUR6BUU
ZYTh5lmhyd1e0wUIwHrqKCe6WB5KW402sRgSFHjkyi7EaUFnnPBLd/SQfZhLEJXV
4tuqVSzi0l++t4HypwADoMhinEdgj9oPAN7dCH7kDAYLF6+IJwK5eZTT/CPqrUzQ
uhREcvDX0y/ZcVIT1PJTRnmTYBLPVB4VsYCdIE6Pvxuzrcbsx6wnQFG0jCqpXyrS
ins7T6hsdZEXQgWCOS5EIGBs7IfcyUrncQ/kxJ9EWvXCkFFIFAAtkXiym4XXl0+I
giUcbKNziJZGSYfZRrghqFtsSfHaFZrTCr6IKkhJxcY0v/u7Mbq8KNUY58k8J0lS
EqcLwYUiLcld9L3pGk3/bheU44nEnM60lAqCCNQ+cpm4HHb2hJMpD6FZ8c4JvB+g
QwxxRhkFb442eGQ3YxmjjSMIem/Ss94UIu/uXwxGe1V3pG00TYZCWoBCYM7JIk21
1L53I2erAmMQIupCjEBWb6gnoA7GJPRwWZloctcHAhoV4dUhwWBa1Xx8JbkM48CA
57G3iCadoIPSsVl+rm3Uj5N9O2qZI/mPQ36Y4SaKgEhU0+TjA0MadZrjA0fhz8VE
veFyrglDYqsDfABhiTTb6uMDLA7NT4LV8ISIuocHG/eQ/mVGzkKFFunt06DIFkfE
fUVCuGLg8RHQCA7237BuQBe20Awk+1xsnR2o9YG8a9MSukw7DLkNLuOAywhKV7f5
iUmL8orzoidc4yY3b6MKyPETOy3wTyeEarpn+e+0XKAv9D8DzUgzpMtCnfs4moW4
El8b6GCNi1pnHHFVK9z6iWGkU/VlbIKtGQ9mij/z8KQzWbNexgnFk5DGX6vGI0hV
ECNnTE/p/awYAs6woZJijjypKrUpu5pZw3eiTai3u9atN8t8slTY0sftuso1XQSW
UF+zFXoa77LWAzC++UJ+HmZ1iSt7ukYRsrglxeWd95legE2HqQHvkQWi3mfFdVj+
ss/Qmg+4dKOuCzZWz/i6RhvPowkb5H0B8k5CG5pRilcszJxvgExHKLw4rdtdMX6S
7HjicGTjRZoZihgC7DEMNJCldo3J9vP9qG8Ffh6tUgdIYK7zG5vR6M4rfftDbBpC
aq3FAs26HnHaX+4KkBCtNZwP/IfynuStKB0w9pmx6t6aBC715C5N4y3FgFtRmsl/
WPkAWIgYLPypgWsW7TE2i56Vf15qy+4jOvvJxNEc6ryWxYlUP0XYUXRfk/Os2IjS
ZxZ5GtjqT4fHPsfNcQ0+thqgQxz2K2XG1Jh7RYcFR8PH9ohui8io/+yEn7Ah2I+F
+rc9sXnBxwhYxw9c3Mf+cIauB/wyp0hrFFd3TDxqLI6tfygG1t4GSoQgTNu2ghzg
qSIiMBy1IjpB9FOpZHcoKFAICetQEPvM9wefkj3H/p++3wgtRcXKOpQQ1S4CX6AN
umNq0dslunGLr6hFrLW4AcokTyskMdyrmmXGLOI1JON1eTCYU763JqYhU7Dz8V4f
awEcSMDOzs/YiS2p/LTOdJFUCm6WQEMpR06k8UA0VKWHqVJ4HFM0tRaDU3YsJuSh
xY85ujh4iGu5Acgneocp3R20VICAGSk1n2rqI1JSZwGswr+OStfhF+8kFLfxy1Hb
q8r8wGyvK7F+MNTuEFh7q++8DkoWF92koPy45hB08TdvBDgZynpx4oS3ROly75+9
vqXrjAnk4xczQQsZLBzjEhrDL15nPi1cxQnPewC2x//iW3f/Zpmi0/jhnHq1yQM6
bEcDI8me++7dbQmfIaSdKDakStYaHP6qdFjpGCvq34tjA1oW8G4Ez3FUXM0QzE+I
cY7QLt0lRl3KlAneDTA+lA35JPgmSUTD5A2N7bZso++2mzxz8Z5yUGIaKfEn8Wj3
97i2no+UnzR5WkZHP+pcRQz79XoSAokd5t48Q/DRFz4J4WAXsSQa9kRJL1bJ1fv/
OasAY4qYIehfH40IsiCVhATwB6CtYRAvs5xlEKQ/XFEasMyqppZteL01gdF5cGnU
Yp1xGSc1PL+/TSP4TnERM8hwa8sdD16MSXFgWevAzWIEgK/Kq/jaRXAuLfS1bNUn
ZZ1QdHAa9HP+gQGUrn7U55cUxq7U+uhDIRfvQ+Rc0KW9WQb+YiFDsnvAlYuIVp7f
QLeNDPRRdqEq3Y4ZMv/cRJ7/jtpJIt9Tkvnl/eprA2qX4rRWrpsfUx5tvzSh3hxq
N4AL6Xz/Ipzpd+BAuwlm5UvqURbRakyeUSq9BTIkqm2ElPSQxcb7NX/1WX6mpyec
Q4dWYuNOz1RR7vxAy6tQDNwpYyaBVPvXbibTv1Dh9RciI/jbhmoZ4xakCZScMgl0
DOGn69uYIr7xBdfpQGwQo0j5FYpull+SGJc1Ig4VhqqktVjEBEP3OMsbcPRimH7u
3o82vGvibecamn0YrVnw3SqPXudE+REswp8LbwjiyvmD7q7n+UbRidPJTY0KhkCg
uhOS+NkSyr4LZeotaWt8pnjqnSNuq2g/+f8YMVIM5A2V6GI2rvaURMyg19MpwXs4
cf4DRxI3ZWVC9SkFdatWR2K61SbQUvq70mvJ2OJTcws00c8t+PevvTJybOEP6pz3
r5ktEVfySrWsMvqQhZl4S9GKrWKCt8RXYfvL40/NC5qcJoM8EnKOjgntGNAWoF/W
eK0w1AcJtcdMTDc84CV1Zr0bHaM5SNKVA8s5VgZXyw2D23CmQLVcvKo6IXyFEkuv
lMpier032HRUOVaJL/EeMsboeBWGTM5Mk3zP4g8i0s1HJ1cjIeVCRJi8Ug/4ogeN
hEUWQ+Vcjzp8/GcOcLbE+LUpwE3nTTe5zA5TVtLI+l1dPXn/wpvvX+FQTsX8e74d
vuM/c73+WHQVHiQxEMkG+YIHvpVlCZx/txDz+EdIagZVJiHs5gTqDA6a5r+8CNEu
qqR0D5XHzwxIjoElLay9EuWn7LwyeJxV/wfrlvGnGUnlnfjAYwhFPP9CL9qS8PMh
SJ0FW1IV2Wgukoq3ksh9J9JW7E8btzN0sQa7F4rOrRw/bmm2maBkXRSke80mNmGa
z9LdB1+kCqPNIczobW6ObYNB7IwDaWMTSr3RSXIkv6fynj2iiWz7efzjVlbfhlAn
MNrY610OxMJSgPDChDYRQI6znHlsjHqP4RImJa/j9QANwEtJQXhxb8Q2NkW2B+NI
OsKsK7DjKmJENK7VxGkY3n/gX7/XCXv44O+GXgxSiOTccWQTXxwu6zKAAtjXJBdO
N10g/a3+FMjkD998fHx7Tvy1GIKwH0HXlcK+kcJVTRqcim95KhWg0/QN5iEv5STu
Hq5r5oMzLolL2pNwSSM2uhdWaP0FZG/pN8Nga5RPngsVDvRkRORBzjJ1oOxe4ygM
auBMTakdxKfhwJmiRl8AW9gGX0pTU2O5MwdLw3JflcycRnE5ulj9Bubp5dbD0c67
U02tZrEn3BzHgtHi/2wgSs4RFbcEuPI3m+ysMIiAmg9M3X6DrkCur687BXU1Im5Q
CF3l9gt2RPocMkJUa02SABhDEs6FZPeZTkztzMi+pNJex6DKkZ2rvkTwXxDjfK1T
rgKgEz3FjnLVZHxwDJ5fPjLgUYqN8vb7LmciEZ8B2VcIRAboI0i0ddcmplQWUems
aMGlqrLd048lQjM2gGemdbsaTxRLKVszf5Uv3El1A9Pq8Eaq7XtqR4BMU11fBD5h
aR8yde/0CaSPhjqFzwlxzipO8IToo/iDFl6HKJXG/HxvPfP0YOW6iS6MYVc3a0N/
gPM4OhnfUsr+t25FryPbDUOoXAFMLHa4nchtnt6KUvkNrs4Tdf95IGrv3cdnOo4M
lvKyqGsusrAtY1RV+6B7n6WbuSD+s55UH0gUuQ7DmbqSqQ/LN285sR2fDG53S77t
yj0oXeHMtUuwgFsS4I10dl8LrCIyNKMX/vTNvbv9tPDkVvjM6CZaGd9EkUA3MDfx
fY6fcqwGcmmtFxnTLQqXeaCr9GjjPgyY/sDBjoH2ziQ8jD66XgSHNbq3pvF9Zpop
QvEDuOt2Qv2ro3rTnuLYdxgkRGTlZOgwBrtByxS87cx+INzOjZD96f7WvXSfGyDc
P+oWyamgrnL9xqCpGzHJA9EcKOLQvyfuYBHUX9H+8ud5gRzwkikULtV1+NgAFuXi
LR4qgwvKVIYF4qBpQpG2O9xzWJdsjixIgEHSYBtwYfdNzfKZuYSrUt/CQwFfXa6p
PBSx8uHsH3A3zorgkJqR73uw7dVem1wHa03eEFwIxM1b1vK1wt5s4XRWIZTle4hT
9kJVeF1oIiuzZmjb0Q80oDZfb5yYe96PfPmRPcsjC6B0m8YN0X+62ICc49u2d4gC
RBUJg9m2Ui/lklHj0NGEQjktbLJecfzVjtgoPnPSXSSxF+9/Xdc88SuOYfZ/r0HX
S8VvrvXzJ0o8iQkWdyPfY+7/bPbKt4xyVg6IzGYzosDvgKol80Qp2tOBxv3C36Rw
kb1dMb/jsSURSMURk6cOal8paE/0TvwG96+Su6HvUcOLsfOd6OtcbNQB51G/dSka
hn0AZ43/Xhl20GesFt8dzaxTD4dBe44DddiPLdtJwEX3LBYH4WAgLea/N8IIwGmO
mCqP+tPD/KLHB+2ScmFrtedKk14gMHoKAbqR7yElb1pb1ZNmJ3q85X3Pv8Kn82SX
tM9VYmO0vpyGulcwp3jJ8MPU5z6xq51lKddl5BtBXz7nznYdd6DCqWRLstEOo6Oq
XYcAQy74Fi7ltKd0O4RM1nu8YgTPW++I3BTViz+QM3TSLMySmEADwswerBGzXGoi
ANUxi4LkRGpM26/dwO0ga90StaQP5DgUj8lvLjeqzd8t1S+WBhIN8kL4ClDUZcZy
3qciaanRTMoc94BqRgYW5AR8d+4NgEZZiv74etKua/Uw6D4kKdDrq129oDKuXhYN
DygZApPEQz0Wc0z1J6Uu6fe5BOSxYbxP8FgCf3bF2iLYxvQ3uh+rj5zvEuUr9hFn
LcmKU0GyRPi09MEHS4OOekKMaQCOCfymydJVo6Aem8dDBLuBri1WkmuBeBYgAAor
S73oDtZ6U1eNczf6jHZ8GXg9NRAafhxRSqeE/JOkw6sy6WfOUmzWxe9HgxgUW0oa
Nuk1m1sLErGVjZ6kX5Al7y++8rlmTYUDpsUsYf5XsOpZ2JeHv9roD7l47acJoewt
Dt3jYLQAR7P8yrvUDWrkuTo+sF0P73b82WQGcHXGTuAMBgqQ6UFzk0eqOB+baN66
qzt0ivayGWIazMyvybkvklVUHl2N8A9PW6u0K4brDh7hnzKNuo2l1Uuk8GYhJe4w
Vv7h23ocTnKWgHUCMLiE9ghl3v/5FxTCXQRbWgIzLZ7OVEl54U4CTn2IYuTBoR54
3yb5SeYgfVY/+p30HAxYk1rZw7JmxTDe0/5bkq5GUhI/ApqsSKuu5VCST/Oenz8I
EVMk8nmTBG8lVa0zn1O2Vz7tuWreeb6864ipqsKSWqUO3mrPmen67DpM9b/+7LM4
747g8SMEZ6UEI8/ajAJt5YUZIL0x898PMMuu21rOV06ZvLeGVK18w3qwEyEBrYLl
x1LU23qvBV0cUSHvEkCCvkWj2fe+UPAqELZYzvFrc+XlUUqolt9NGtlqJVFmweQI
z5pg31vrlywksO8vKC6iBpZqIp7NNM1If82TCGlKQFsMXATYpqMVv/i/YF/CKcwy
YvdeXpWVrClW5nNKWuocSzRjMhKYb0RbLv2hoPh5znVX4VqD/EpzMNaMYV1oNiTW
yH7uSCKCLBzOUE4iAF1I2IKpOp74uOddSv9wes+JUguHKx4UG+CKKoyl3l0uo3Ip
yxQZ+/3xalFI1ROxgvAtnIL46i40xw4b/40k2n2s8mNpIVseO/DGNK0RhAyp8JKB
/3ztEZ8WzSG39rxNv+YtSHo5U0nEdk43rhLR37+MAiBk1whVcyrGpPuUc2q4yMfw
cg/q7bwE4OJoJzk+qa/E9jXNnW3L8M0vmaYcBOqy/73F8WZcbowLN/P06+rckmVj
8p/3nzmhOXDlWqAD0XJgBvJnquYXswDQb1TBv/kgLWGmbzeXVMgfnTMv4SGb7A77
lg3jUl1ieRD0n/sACdi2h0rwCgIIvMVNtyZ6QUz+D0iWNVnwO8NEMa4AJwZVefyQ
PShAdBZ0eIMkLRfZmUAbf7B+1yhX0FYrqN7P9guashMrvGXF/rrKyVyLGNLgNGEl
oqrWiz2oQUS1sgnzKo8/++F2nkK24+dIbEgnSv6HisIHQOSg+8ed9dpHYyoajTvg
v7CojhJprRbPKixKDt0ERvtyvDZkBUTYPi5m6zYchRakhKZ5oO4dzPhLXa7QfDBi
Dj7A/v4b9gSqU4P8wyikPeXGX7b0ZAVb3m0Pph5NU38gQcF7LeQ8NcV3ZGLbektV
EWQrDJVNx4ZYWQWcipW2iUM/rUC3xJMPnkJCz9qCOaj/nuUg+MaSuxaAL2e1/c6T
U2zZ+3LPd303lnlbythshfzCnzMeO+9te0fATQ3oqK77e3Zrm/SJCpxCs4hP0Yq6
9vFZJivTb1GLOA0sQVtYY/taGSH0cAPFNCdqH8LWaKZqy4MAIR5HF6x5N76QaMhX
hNbqTgsokITFwdH8Vft7u7jcL3uV/WeOfG4r8VGcmt7GQziYezPfvJy65N9nebr2
B/G/28tkvUH/n8gDYo1IZ4WGLiGyBadjxObhwl6qdt9pZFZEIMuHx8+4baYJvPAA
wOWbABMxnqh/vwF7bohPWTDlEJYvWS/4ZxH/4TRliQAVG+d52m8PWfBh6LOFP3ON
SEnG2QWkBTPu+RL3mKEGQL53D6o2D3SwaFQmmZUfaS3wzXwDNLF/qOrRkXjvXe8H
VSeeUV1M4csAx8yI0cIPQ7CtqxWUhRExyNSOfM0rX/smA1k8f+iM4B840OZPSwxJ
MOjGPT3koBAs+iIzgGeBl2FDUpwuFsSkBMFJpCcGjNCzQI2ZKcoJhGiW1fcgEdav
3e7umRKgGe7IwuyfTuNpPE20CIf75cuLAskLsvfC4653vWeqZsDy3zEtsO3gv7cV
I779Di+gSOtA02634reLSFUuRjgFec5kgBB20wVv9pab6VtjKrlfwGNJx39ORdNN
5hMWYZcAv9lV69JHK0sJRgP3bNrhf5fG7oaRwhRyp+DXow/B4W1KZjPf5IFwuIrn
xnnGMovjjtsre3U3y5//eau6F0rZY7LNXVGIB51c82dJitk66hXezzmi2FpMCt2P
rb3DemQlxyZf5dG2jpby4duE3zZFa6hXUL9qQYwxCSVoBcF0yDwSjkkajGzt8Uv9
ETm3Ro+RY7oejIWIhvy6hqWfdFPER0rwNp4IMPFbD97I7ZCnQnDev2fe+IblgyMb
affyRJTu7+aXz7AAS/wWLYKCxRf7UlEx42V/CrrnFoABEkRARX+yBG0g1kHkbXRZ
lkFXpTsDyl8w0YrZnHenHgZSY897uNLK0vmoc2nAY+hFzKBrhD+bNLVuyGGfgDT2
CJh52mRqt3w1FmksUvnAZ1WieoE/0qUZOMAvpzDdb2u5TIuYHabp4gU6WnipI9Ie
XzmrCfaRlh/RpVqxgKhO2/nn7nZpper1pAjokG/F32Z1Lm25Ksw8+CGlz5MIOdSI
kBZLeKlWibEI4+cRtWgUSXxsdIDTpX3dU9pX9z350VqCIyDoJKycESwyCpbSaG3F
8TXkflyZ92j/s0JdqI+EpD/SK67WdJxcuZSDyOcp8LfHQ2FDpf0ZRRYg87yghyRT
jJtAQnal/WN+0u49khI8nsReVSujDVspogq0RMhvFqhYulOxFn1l9aBD50uSqEDk
PL0lbaJVp1Phml3g6rneRHJxk6vRzprqsuwBIpG2nVQ9X6bc4127b30OtP7QPxf/
Gv4LLvxPH3if96OmbBjCeUIPi2W1lYnCzcaJwEwXfDOfIqM5R7XTC+RhBuqg1/jv
MhcVBjD9FJIzRMFQuxs+0yfiWWiC+NUBCnzeGr/e1U735eOSFbloaTNReYv6z7R/
6BlC9mW/vUyr80+J85e+rf7VONuwTHPNUWQdO9f6NZPYLuTVznEDTD9TRKqCBKws
3PO+KXnYEnX78FsaMSSHASZhw/9gRv6DMsO6UGTj4dKPc0IvH96f1yyrBe1VEXdh
cBGt24oZGpcHaVmMlKR3aObDgaORraJotMZweUJTZm1LLe+Ps/O1piRk7nGKfF2c
weZTzigoNgDF40T/q5qNtUPwIiWt4VVjkz/EcccID1KdfZ/b/evxkJYNaeVLd48X
u7ZL9XW3hj49JCO+vvS+2nA+xIMEmEMZ9FSaPZ5F9nyFYjEC9yr5ZODkZlUDgmUs
zRBU4iXeBuOvhk53ejLucqSUCKZI3lslUihb+IU4erRpWiObGkj4W0XUV23W5a9K
Gmd1//CaJyahq86b3TSJhuSQrpr95wl4EeY3xMcXgGi/9I8JnlQnNuUyyDwPoiXM
ZK5m1bdyRYQC3ly2XE2GNuAxG9qfDz20KsMv6Y2wvcpSeaxKeNXMlNyii0K07QaT
Iv9gxJiYKNWN+MP6x6NTdo8RypqD/7ONlpvkf4I/e5o59JtvebscSTTra7DJ4P7q
LF9fFgkDNMjOZpTC9KSzYweGhjLyhaSnJi062KgiHOKdRIY7S0A0PuNowWA8Tk91
FkGMCrxR5Xc5/Z0tCs/JT8btVcvvAH8KGxQkdIoWljWO/VSwd1C74if9JNwunpzC
LsIkEFcdQKpMmFbryNO8QkvTUBpp2hfu/OepjTffAhODCBr+CT7nTOU+fXN45aZT
WTJdfLvHN5h7szRIr0+7sU3nC/yzi0wACHrIwBc0Ob6+6zktHvNgz0nJdmWuVXm+
KFBZfaVtHkZI/ZJ85qWd4udfpDyGIYQ68F3qcWQViTSWf9rFq7WsaxzcJGYqMwG8
E7zLYzzuFSyBVhQ0qTtIhjOsn/2Lpmo3YfZZPE7Hsa8L/l2iMrVK3hGeT7JkDzl7
dDHKzmn8FZeVMKCdbKbB+6rP1ulMAWRTepa5YLrhmupB0nNXzwfmgWFTqs3Ok8EQ
SIiGGfueu5H0kLcPxn7evKJrbBKsiRMsHl0egCmqCtsr2og9zGvqoXY7C2C0+vKp
/K/CpPnPU/WoNXjgt1/PfKCk/Wg/oIYW0Aljo+nKXveh45GquioK7SQ96TWGTzNA
s3OJeL/lbOgrhKMxl4huvua0hgZ7Z3nlnCt4VcZFotUR9c9ZfcnL2C0wEgxueGaT
d6al+lxulA+YiQvGnXF69sberOZ4wUM14vFUn8l4NuRGXHD/7OZZ43O830TNz9TD
L4WFCEO4aTtM1BfaiPzaASJ1OB5GvUVCC/ATygJnnrYllj69gPBwEl+2Zhwatz+/
CR77fUuHeKFKXuN0uTlOgVQ8QzGbSXqtg5bD3Bqc+l93g7vFoZzXbyGqadlRDscT
Iqk8Q+M2O/99MpQLLXvPawN6VDoAfwf4a+rRJv67h7hcurBZwoWTEMuKAlS6zLTm
bjpCt14tRxAqRtPx2Z0bRjV5D9aF1OG24SbmCcXam+TE8sT9g7QzlJZOOqi9jFkE
iMGYMK8mR+NWzWafvyly3mZCLlh+YNyls3hQTKBC0mwCbcXsE718ewPOM5HAWRsY
sjtg8wS66r4Z7un3Fur1VUKb+rs1+dSWhwLEALryU4ffkoZfDKKQ/sqwsKQpcR9M
wByAG2/c1BgQpUuO0P9udnyMOIrzEhbmlGW2H1YO+XHzhYY1unA8QSdhdFGBcrHs
lc2HBWFdkECA/fKj7YAPBnSzQAlJqmpTRlRNhn2Q49G/+Vm77gw/cYY/vAyOYfPY
WczT+fosHgBaJmoIdj1KH6V0xt21sTs21+iVMjqu4d+BTe/U822uQccFoGrqVSAT
UMxT/YkVEaHpC7v5dEQl1DrXvIhBr+QQzrymvp5rZ7un1Nmm39Spe15Q4XAiHOsk
ZRWh2zc2mq+oM2hFahDg9y2wfCDCZ79YYnIc53N6xR5Xn63gtna9i4QB62LNR4TV
7kJypmYqWmEm61s00Je8NOV7oor/Pt0MqJsUhJVmmATAmXJpjZKgGuwrTcQ32Wc7
7jVSDjB8cT2oU37ohAx+swKyny4DKGD4Vxh+VYibm7W2uujvoGHlTNfrJfcKIuPD
notCJMLdg4uiLGvPu0DLAWZTio5QlwzkQ3wf+OpldpT3ojQYUcGxzFX5jUSxPcnW
sjmCsmDDGhPhGjNS9iX1elOKCkedCBZ0Rg/De8NWO0umRCkvvviBVlcUJU8VPjWW
iuPLWlXIEYS+0I5e2zWQ5gI6fbFEhcRClqb475+ho1tf3+Pj2MqQYbXv+J4z+4Gu
LWlXzysy12gvUwcVzA4PKmkNUBYGfOaEjergMsWKw035SGBI4FubstoIV/nSIKP/
TH6Fj3mG+bKvN7pfTE90digkMqtUkzLvLy/b2uAA2JuS6CdROrFMiR5LMQLHuUrS
3VJE4OeJu1p8m7sD8ORN1rDfwacT0KXUIyZOPOIAlicmx/+K7IIMPflnqjlk8lvO
VGNz/UzDFgjCH23tX6SUnJQKFznh4+dsIFeJXYt7H9Pvjcqn3/NDdb9CrCGw73vM
GnVMOCNKMLYq14fBDzAYGMj/FSr7zgRNUkxxS7S4X94vp6+IAt+r8h9fbmq4L13D
WegP2QkQEHuqaMTIYAxEBh9W58Cqyhn4PEzJuG0lhhx6IvZ3QlTU7YftnA1InHo5
IUFVKbSIGdzK/1hFvBI0m93/UbgAMslALELsWTshOl8FqMnoGbi67EjKgz4HlqyV
uUViX31M0sU0AJ3MqVfHYyFWn1RGFYH8OhA0J0MKcsxZNiOraXTPNjlYzFanPysU
ExCnIaYyGvjkm9yEhdbwzL04wbxJ+biR1BYYU9oJl3mrcRZ6ndAbWb4N4nOtjF6/
dmtXw2ptID/h2DhMmge92qNvgtI3dKOfo/0waqlAJfnwLEcnqplyRa9vgFIF7vV/
uNCF7RxAs0N0SdPMtWNtRj1lu3KIjggCI/wSABVAqfXf15UXabmz9RPA0p6NZ6TI
e0SmmdXJFtqgob/VmmsV1bhkhby1ECKVKeDsByDkY589hL/6ltbmxqke5O6xUdiP
Nj65yvNcD+Cw7um+OoDH4Lb8Oc0Cd1a4X05TTcSm/gDt9vBxolxauY1ntq0cr5pA
h7qa6kuwzeooyTqatBj7Gyn9O6U/IPplB0YFK4pTJfK0Evesh6SFITlI2JJUQzDs
q3KOQnrwKlYgJ8rpcFGL21BHye+9PcaB6JWa2ie9a/2K8muQ956AND24xzT+NgMe
bAEFO396e6ux90lVjC/oFgaBYEm6oay5MmyHKBsLz1MW9deWsFzjU/EhUpfmrKb8
vximOnllp7JoJCHWl2u+LWZ7c1AEBxTJXrGFkEzd6n3qH9FHnwCaSnEKTkix8rrZ
oxxr5jgbzBQ5JXYXOsf/E8pg8ccsKcU5ilfdw+EldnOhaAbpu9ytzSeSNu34PK60
8NdcWt4GVdwbTIJo6Pkxqeeo8sbtEp4ehYBglRcq3LFse/8ru8qcz56qAIitrI1x
kgOqDfDU6IOhO/vLBFhHDV3RqcAatVvTQXyiqFbIlxiqucR/AjYE9xpKikIF0o0h
/7Z3ZpZdCa92/8aaYFFfP4OHMuCz/fltF6+OemEEFwGFBA1EwW1Cp9WVjv7ZKYf3
By9HtIW1dn28nLWMQfZQsw1ikqsBQerTtifHWBpYIgtpwdvwnInEl7C8Tl+cc35t
mYJ2WKulSGYvPpXkzRnUB96kExwfQ8G9GtXBVx5ZEubqS/g26y3lqYrV/74rbWBw
8rRCEv3FykGTCoagZmPhXO/KYP/XElv3TCqqvdqCbOulEOF1Qf/Ireq9HQKgfzI2
aVUGTooeQ7KvUvWcwBQ8D4A3ywgBgSKIhHBTLAhWluYBzQWOc2LvG52QuRbmktw2
VwkC+aBdmE8H1+WMMK/EgljDFnx8WYe23/7TMkHHUPHnThRbL1dzAwlLaZ7Wy6qa
aZ/XiqnPB3T8F3hQZVwY9m3ZMdzl+80YpqDwC+HbUH5F8Ih9kqfgnZS5aETBxFD5
SRLo6A85AluzN9boJJBsA8p0bANlFeAhmLqyVCzsM7YvP7i1tmALvOSUUsANBZ+4
AML84kl01N6/o14bjOVgIGBZwZPxqjwsoe1Alvc+NqdLDfdqvw1CcNJfDjFXFBWO
No9mRqjVsQApxImV7itjAltp2MOBhkToqsixXdymRPiOy9Rv6vN70lfSteYM5Hp5
/Xg3rPnG93wP1K4iOigHjjn8HjS18SOL1PWF4NsBH7cqPRVMhJjySxASJTBVdQDt
y3woMbbQK6scywc0jCinFsBtg3JazaXNZ7WqbADE+YrkHckqYhLM2K1aWXeP5DhC
sSjmWMSlaF9oV5aNH2Y08Q6DTQWs11XneFM0j/vw2lLnioCyR5UTFO9Y9yBjFSB+
JEJDsAHmO/8Rd8DfhAJM+bw3NefFytp3bMPVBEloIWKNjbi2v+gmlXHZVK1cTg0T
sh+84xkd3bm2uxIdydnTXy+GXEDLQ9ZGGrMAZLBU4Rp3XeAajgQvljp9Jkd7mjLY
M/UYy7HnC+TifCup49Dy/n2e5CEF3TuJ8/bkg6ob1mFQfPUxTqUyLHCsQe2/V3zv
AAeQ9KD78oSBGwCiNOo84MLWqisflLjnTHwmh5PKUNcFZiY7LomD3WpPag7rgxWo
xwHeg0QTUuQZnJ2i8aUj9/mJexV0fskd01G55R/hYEQ62m4eFslDF4Anoe33H6ME
eumLaQm0iuyYNABrJnm5RRshEhSu+DZwJPv9u3W8i/xElVi5prcbEC9UhIKmw8U0
E6+5LUziG5dGuMfOzpBd3CKD6m5NdDwT9/GnRIGPuTMvpx58eZ53eN3m9uSO3HiQ
XRWy8357L7lzsezMlNuWkwT7ID4igHAZ2JLyh3c4rGhYZ/D03jeuCQerVL/9cXwB
bGvQDk725GPlUsbQNYPSM4S5+f/gr5fma9kGzmV0XEyn05xAF9uHpdEg+i27gS8j
0PzowPgLi32GQh5CMO/7h2QceQY9OHEHx1U47N4CHKh0JgRaW7rGm79CIqhxcyh1
K+r9e2mjqbo7SlB94GcJUu3+foCiwy17TgFc3AYu7p67GpkVo2l8qxBO+6JbOOP0
R3Vb9/e+S7ZZVhAhFqob3o/Oa9wCs5/AkFmLpc2K+GMeX2uF48xDyonlbIhCIciL
KEcSoRiTCyD+Tn20QX8El6mS2eLRCUir/bALExHYsJP9kZMS5aaf4U27MasVjzTs
V57CFxb72KsfZF10KlJleYhw369rKHrKIPwrNzG4ZVcuwAa/bH/nTKPz1k+PIFnx
Sev9nA5N1gq+9qf3DmIbn5HfiCrM8C4KCxaINV2E2im//VtKqWiMsn9aibh9t2qg
/OrQww/9uUjMRx0dO/clzIH0GT7QX7vlAGWYpUpsYeevyX3TmwMbvzMgxnmwyJHm
R6EC7QP6QZh413MXiykBz00DlNPVNgesoH0S7j5Ljl34kH5mjbtFAcQJaxY30rU3
Ld2nR/4l/7cqcNxc9YqmbxrJ4tTrWz6JpnWHlQoxrxWs+IE5Ya0ForOnHZdYbaRD
8YMIVjrQry9uWkaLOdz2gJst3F6rRHFD3gDbcEcDtp6Os4Gl1q2duX8SQrEJF5DY
4Uamu8wLukPzTJemT6/8ApXZiWLWokJQEYT8BoZ6qip244SBtefLN4WpGOG8iLlg
hKp4emhOzm3pm3LhUIzzP6ukzyCt8WPv2BY4otOwieV3/1aA1OX3U0uLIHmotO0U
p9m3sf/efXIGeMJID0Gs1fRq8piXvM/11UZPjsQU6CvHiuF+mO5DRtp2VsPzsZ9Q
GvZGjFW8muXN7MwR3JYjJixquCHYMcbKmPvnkAXlDFIkdEzWtCe5kqXvYSvLFOwJ
ddEQivPuINRT4T2tXoMeA+LeLsz613tkvNs+NcuMMniT7U+sq5iJ74phJf4iFPqF
XdWsVYuzv6LIAd/rp2w76rXtyKaGQceUz0XqHTe+vSmVlV4/lFqJLcmPyoms8yZX
CjtB7axFXqP382aiANeUTcn94BcX6atSD9dYc2ogcaDPQlGMR85jizf6MwVrHZ8C
OszCmyJ/DAlGoehLjO5fd0QdYrO95kOQ5HpLRrFBEHt2Sre6kWoEOApE7Z1voh/G
kgiYcNXm2HjfO/0DNrYULj4PJwzxPqNbmWk5p6IYez2gaOxxPKGXHvQQIjFelKzP
NqEzru7t+8aFQIwdjyfEe0gM4iviBgBCbEsjVOvVwBpcAwneSLE9NTV9A8G83szK
gYnKj3nmLuQdI0G743i+UXuk6FvRF486Ah+CLEHNJG4BHw/gi6Vc3TZCo7k3Jq+F
O/BbrJmVSw6pUd8od1n+/h/XibI4erBv/tKG+vHQ5Q6GcM20ErkMuU0r9CexpwG0
+cHc7wJrg12M+RM2Hu1IxJ1dwht5w84RiVwSCTDgMc8MBJSsE4nlVBp6UHvBJdeC
DjRs+2F6XarpD5444yBIiEPDdwXmEeYGYRPYUzqXc+gCsm7ZJHaI4udvwswruyCg
YQcdFFdww4TBQRqHIck5Oxhex790MnO9pCbR5dFptKbxYJmU8QsTBsRrctJX2JT0
duQSeFqVLyltQwZWHJi/J7tsLWwgFH2OyME8ydiLF7gXUbOXkh6wU09bUgoZIJNQ
6I+4icIz7zzsnxeSm9xuxWo2OFmqcSZQUdbsoA0JuB0Bm9R4nOG3bWJe9L+Qdu6J
qboaDgHqZnbwDQVXrubxKIR/HsK4xrZu3xicZA7bGMel+9XpftLwzX+LEQOfeS4p
Elz3+AhZ+dBYOA1icRww19EuataDfHnbOwPKC/wIUjcObs4r5tv/EjAuAc0019QQ
4FhBqG36Dqg2et9ZdAg4wmhHEoZrGonvvpA6YHvo3EXw+zoR6Uv6BxWSChqyKcyh
83dIlTprmQsJl5kfQboheIANHiKRiVdHhCKacATyMrrg0kkEEV90MU8bJ6eU2+ID
rJQP/nZYbdf1VZbABZPbE2qfiywlm89lFPRl1C6TvHO0kitjXkB9sxMraLLe13hz
dbS72ZhdklvMlGZb++uwcXxnA8xVjX302n9voPF1W4BccoMgpOkLLChiS7anfdsy
2FwaifbtKPnSnMCmH0PRF1VqJ+bG569uEtDAuz1JYal+tXz0Xdgb/kzRqMssl+e3
3CD/nu/xqRo5HhmDCSgoHB239EDm2l82/AUp9FVPQZEYvJEMR+ocg0W2jZP6YtcK
112i/wLwBKsoGKyrEkk65kFm9uQjDY/+xZAMIgWm6GSID1lRIJ8OBP3EqEUwlfxM
nKOF8cVBNhWHrsS+e/B/VrtkkE3h80L+ajuHIlwW4TX6/lC9xqj7++ZoEWzDSLub
WQZorA5R4lGbIiMY0EUtsUCE9viAuDi2l4hHfZZXwB2ovN5XZgkBima1dbScv4O5
M6fZ/k9GUL7Lrrbs/oEBOsrARRA3fkWPVuuS0HmBWm2CioiAftfV7ZZqmAC/R0UY
ld1tjGDFYKsrskpW6UMbukMFwyihhKeYnAvsU5wj8D1aUv9T4d4n/GQBvBVVYLNn
agFiqqNv9WwV8BeZXVZSwR2W0He8S485f2PQ864mwkou1tLnXVTOaN5O/zb5pqxQ
FsCKxHBSacDIZHOcW26wdZjRmvv9ing+ro8+gtAg0WiktPRUyEbCem4d+CSduJ6B
qaq0idf0bQqUR+YYtVppNIMkwbb18dvWpceEpg+HGPwetsSISulhFY0yzTAUTS/2
s81eEGAdajwkFUkkEVcUyhexnRySqISef1NeD/AEIOT6G2qpQWimvYst3u6CZDUW
rF4opb5Jov8OLrgj3T2KZ5oNPPYb4GgfAF21zNttLot2JymR+42mFpTLuyxulft7
ybwO67texX5/DZfh+eRQnzK9K234Peo/sx2LqtHtHjz5+NAeLBumLFvOpUpku+x9
Fv792BkHURbimq8PKOjzUpwbxxGH+UY3fGGPVBUlf+jTN2nUcpPXKWgcbLVWugGC
Og36Qfx++qWOL3ObUr/9rS4SQvRgcD9KeMz1gsKLInHB88Wgg4dPvi6/qXivCQMA
jej1Gubf/0g3eMw4GP8Gmk4G3t1kcCACuvJi9134w8g29Jk0FfVbWeIfEsCntVf+
Yy6KWV3asfj9hqv33cpfImYdOQX9C+KNHzgrNiHkjT99dclyO1FdaPfwkatcqvk2
snkCF90eAt+0v3YICrMEwquNVRcqjkcmDNUgQR887iDTtu2tkhVEW32cTLeqTNiF
QVz421Rg5JvdfTAWzxZ9XfacE6RtOl2n0//6QMsC6gC+NMhL52UPUF1n/MjC87/c
yxF+VnL9I5xmsFU2FVx3JZpMhFFPlV3InALgxEsJ55BwjwTt86ZFuDdOsjoqRVA4
Wh0yKURwmsrFoVfQtr7M+kxIYjxEY8gmi7J2OEIDbbZ4DYOQQy3wMXVfZqyMVAn1
AzqUvBQcE0BAnPmFqmAo2/87Jk/bf8ELS0FQ2mEf59Hz7uHt0v2C4L1F4j70jnLk
Xu2hW4B3tMwLHWCsNxzrymQEBGfpTyOhok8YivB6lcZ8qQ99mVzRrvCKV3+6Cn1M
i2MPKILLxjOp4PL0Lh+LXHVMQ5jwGP7MmtTSRHdQ9OYCKPrS+W6br29FP9VXxAYQ
ASKe4SE9a9oJ5Wp8M8AuajwWInxkehU68cC/SgVxTirpsBB0+DcmsmBpvVEuqW4d
f9fLSrJEM3vR9FJNFiLf2cpOT0s48Igg98ZarI4TXCT9TB14xR4PTAoaUHAvE30j
6XPtGdZI75jt3WwMUKj/sFbKdnMhIhJWaWfb5eFO7KcKrvUWQp6tYl1R+7ozqrHv
1DVwE+OZyhv40iVCieXWkIpIkn9TxrGGCtN+MIH6EmxNv8ZbenV2GUi1AP/xhLfZ
c7GlHUDd3dnouBYcDi0QwHjsLPEYaaK1xVJUg90KCLd2Dh6NZzvRg2yZkFWocbu4
mvsnGvGf676r001Dns6fohe8sCF2zj40lAFnymeh85IuDUSHN09QRcLPMtkVE2oS
h2D823DPtdoMiJ+ZiH7DaJhU+Nq1YpQFPHWB2ummdDee2if+GOeAqzVQZLTGcQuS
vNJ/qNTqItKaZa6HsR7RZ9yJmWJR6vdAdykQDcVkT74+JIUxJTT5a11O1EcBnK2U
PyWYQpJHP3PTuBBLf6hZ6lrCx2HRFWbKtmPj4cTTNBwjKZqeRXbFPCXzRlNdOyho
xrDxkZhcSs3kXX/QXQFZws2M533TvodTqygjqwhhrSvuKP6aBlXQouaS3esyQR5F
Zdn7As4CA35jASZ/Vkp+Khcja1MT1Y+YKPwY9/poFK5Cl54FpLEiZEM8i+rp6Ndq
xM8NYo1DQrVh1ReiRF4lxJRONavsddSMNOrWWEOO2KdHDvHS2o8GbWt690tIMOx2
XZfmzZDl0S/jSwiuJTiv1jf+va4csynUI/1yDV+HcnW9GwlmLJtZgIvgiTpX7CPG
pSV20oisPd7nVefkWUMYWLn4zM9XrvRpUey4KYDGnIqbMaHuZhOLZqbiGmxQX3pk
GfAQbSHUB1E15qkg+xYs6eTt2CUKCfpKMLjN6oAieelLOqcLTgOU0xgDUJxndfX9
6QMupeKdulp4cuOjmWMIzcyeDDOe+fawYARt615HHoLgnH3JgoKc7YrsFta86qVZ
MELtb2XulE6J4/7ccYe85DCpyW5JTrzMwLrSVR2ezXb4jrmihwcEn0I74jpLrfIY
Uy8r07tqwpUqB03J9dlWQhXlLe3Fz1RfKGOdOjcbsdi1wbEPX3bROvdhaLIJrxGw
2vIVz6yh/fwfxwi5LPhuRpzvktl2yYwX1BjBxCAyQtDHSjslRz+gjXTOEH3pC8Bn
u7K/bgFCYyLDNMlHDEeOxC0QAFH8xfSVy8wWCYV7W/sGOTJ5NeVjitKpH+faxmuA
0FN7DfC3J19MSRcychzv+NBoA4nzIrNrby1eS1g/a8JQql4Z5wLFrZDUyI+Em9XT
V/RmcStdPukyebYR4LwNWnVFzO+f5r9ZKGhRDpH9sAbTvPucQYDMj7vKc2tiTHLR
Ii/cKNgot5ULxoux/nJU6Rtw2XF2WqgCeeo40TI7B6jfYA+uWHtYzgZ/dUAu09dm
pid/c3rsBOWJ+Kcq6S6PpK3NSasHxIMPeLKPuC/Do1077fxxpheW22KSCAhaRmsD
2ppRenPFiDTOml0f2O6WnyhRPYU3RLyQ1CklqjvZkKfHE8v3gzLUI/4jUESiKwaX
bJI5j4Lbsp/ggxCLgsZT9GDDtP+J4PsG+FcO3zUnh02Rdy/SuV7ZXeDaTPQe673u
YjIBA9qLOcQ/C+iX0zR2SxjtlvzvLOvDMnWUQdeYKzoCp4mfFItWG6lVRmDgnPNy
xobSq+JiZKUAtEUftZr6hbjEojpEKlXSbTU83zd88bGflF6/PmfuR5/5glkaHG3i
ltY0P22jYb2efRe+qRp5JG+8Zf8BNYV7jP4iVl4O42FvJO1BXHZjrZhWXTzDsTCQ
hddFccoeKdr3TbwgYBEGsLawsTJclsNmgspjqWaHYtP9FUsk43PSJ62ZjwbJ7GN+
vPmj7osc7LeONTTua2hs5+hwX5QYp0n48mNoLjf750UH25uQ6BTw3JJx9oGiGxRn
GsSe32MtgoisKGlJMwxksZgsGbhNDZpkkDOnX78GZfbH14Q44MIQdxUc5tCTAGsS
oaVHwx3qKRVHLUo0x4SxzIkDv18dBem9OOyiUqrICPB2NtkLVjgyXRLWshtQob8g
JVNT151qC1kyfUKdxLCFcRHsjQcLopzsFPR1C8R53CSa6JtJ+85q9BAFIxlST8rp
9PvI8d4gssqPiPnVA0wFxOdd07gW5QbRrmdC7mjrFuQo0rbtxZteZB4YxJadOFRf
BpuRPN4j1ccBEaA4mRpEWSD1VQ+UcUf5o0HC8ozX2UlujnRFfk1ON0tQ1sSWITzH
K4kNYvNL69dWiBPhLgxC5TtTHLG8jKo4ZjD/PKWHQFZT4ZRpU+oHi0+prIrvZyxw
23MpAIeG83mSdrcWpFbbDgEzvlDuszWKpwHBUdJZMw6SE+O8NX1oE/depAg30ovK
8Z0RpKQcJcmh04d0DL+BUAp/4Q5foKOzIkf1F52+noRK07ASoM7bgcuZOOdRmOil
aZRtuVUDIBKqtr2mOQcPzKxOdbJXfWiALgt0LAcFYiypqmvxgV2ufQlIGJhKbAdK
/REi8tBNRxUMY0xHMLqp2XJ+Yium8oDbTzm8yknmnKZTzCPPblg5XaAo78aTyufJ
AiqDvoTDJ6zfLoV+9A0uYvJPuZj3P0C6FjQqm71cxKnktyYdZ5cNhP4v6YVFhB8d
1zGSGKJVwVLnw9QlNWum4T0oJwg+9mLpjAwMADlm29MKEszwlwy61QStxtojgaYW
mnU/3cCFosF9hIOJGNzMtXiQKDtA5w5AWEL5BMR8mkyqcOLlbagTf0SZx+dettmK
wlWFFwS2v4WcVJJcxClaZD/pzAZGxogFLNJOPNRGaeI7rBCZL9HhlaYid1QsKoAr
58js64zBt7wkQG2wMFmhbQRLyXAIBCNmhCz8AkwHCvg1qzNqXd4Adrc3p94VruZe
Edgj82S8rISpUo2tou3fG50LUMEAPR1XC/jcCv9PtPqfDEigI+8W1F4KR+O9ArOQ
LexZdQX6lGgAJWh8Pb/JAeg62B3TBp5V9BJgknSr10hQIE13aH/N6H3GeiDF3AOI
tEr+VAQ45JmaUd2pJZU22pCBYbK4grEDUCTnw/hHOE9bXQ9RSn8/qpODiWCyryPo
bOwQnecIL+Vk5vR5QZ6L0zL6BKSm1bwhdeIwe1jSwFEzl56VSYxBzgmI9inIRPyY
YMYDourvCUem8n0jbhesGekmN/zYC6reAfV22uxF6QhClsJhG3L/YNS79VyDT4ne
x+oME2K8zBhS62RklcznlJc8Pmq1d4LDt9khKt02hnw+O8wMg725Rx0tPzZ74OHj
bmcGj+XzsHiVj8y/0dgdzN0ZkZl5s5xBWJuA3aOMcr7AHA3R0hz5IymuOtX4fh7v
Zzt9SDMl0oPPoqWYZxWeeKrWKcvkaz/BJ+6Eu/PfF+D5GvggFeW7Shx8gfMw0VBY
DwUZ+V0xnJALoP8DW8MQbG6UzuhHKhpnMlvZd4SkkUsjFfZ2/wl5heu3V82g/uVG
gvv5wV7MAC40z0dHyA/7HQqLu8s+bRdsLEEhYM09Uh0EDBKcbPX17jPHoAqZAgdq
4TxgjaACKtEuCtIBXsfmCwSYIb8Ox5q/P8AIJ3UwMmuFcmrtCD9fHCqxK7vM14Lk
UxyuBFWXKFYH1s0C7XrBVaDQF6lh+GPNcuVdKjI0z4xJWvgbnjLC0C/PtmK1oBWy
qKzQ38yppQ35LXSh6C5QbwZOF5yoAuMw7RyhngIz77wylYptrrlo0jiSnt661IRA
pcF6nBCWZ5s2psP2zyi5EflGqBHPgjoYT45KSrAszlLWDPq6l6iwt3UshEe95LOF
vgvjzu7sV0s//CN2xdZqOqhjZ1jAQM+8UjNDSItXPx+GSNxKFnaKZgwhWtrMI0me
fDQnFO9QH/Yo16UvHBwxwVIhcAEKFUoHGYQJl1QsxNPHzMrPohlFRa75AMadcm/j
XQ9YcEYwF4qtTfXdTqDiSxQ8emCCMu2U0sAhh4adIFYUU5xDYNkx34Q+hJ4+NCjv
CA+QXyK6e+TwWkJo1fXA5V6C40wPSp0+xDFQfBYY2Koyvl+MqK9+blgqkTKNXp2p
OYETpqP1ELREifJYEHCoWNl0r3FXGw9bqtZS/QFEEPIVXl9yl2d2Qi8/rwN4vm4k
Bx8epYxpLW0qBuVpFq3YcPLSZlx9CCbqrLCgLV5ZK5CwOeEeBv6dFVSEp+ef/Of2
vU++hfls4PJnshXvvMpe3fhppoeGHTkjou19eJrAQo0jTkaqPIJgkSP3TzIFP0sV
QJbKcmUp63JRquMXyGg60MoxwyHb2xqO2lEqwQX8G0gx0ZHP6nX/iOVtwhrUcGU1
dDmLXT3eeh/xYKBEf8sAixVCrD8ryH/i4rJBPqtPHjLQPmxvck+IemQFj5VImLcX
8vUdHEsmvmoZ3qkERDGI1ROpDqjz8ufQkbaHge3V520CU9dSHyTPHpvJlokHpS1J
CTNCtzlUXABYrpgLDktpbmON9/xRHYu0Y/le4P9G2Ko2HOWHK54N1vC8e9hwhxqJ
enOKdfXMakNnUElQjJ19NyACQbOuY8F3si5ybgmCCZXwyYthtYhJ80Krcyu7uodg
106EPeY1vONzpyIVfYvUkGv5BNZ9MzQfgH3d5s2tOu+745y1b43antIvfqghL/5u
PtXeIWgpmzjkz6L6EDN9z9o/stjSvDYidEWRW+BztSD4FoL9/TXorwxY3ZGTXVD1
l5JgCKk0I74zkr3XTVYBw1ePBBJhpqbgIOdQSTeXRRXnatYKUKx6IjJAxPUn71az
bUQ8pd7B47CsIHV+o1NPQcwpCxW7RdJQXAYZe1aHJwh4TTCMncp4dk3s0tQs93tT
+4mIHAsruCoFP5xUGvvUhozG30NMLB0ee9+WEaOcKmo/yphrwfcTuIi4IXVtiRJY
egCK0xfxY76fgb82cTyDUZueH6tnJ5Xeq7JlDcWgd2eW1VMrZF+qFwLJMRrv2zm3
dJ0euH9i2QDcZNr6q2WRFdXdqXCCz2I9RJDEC7sCWdu1FWbDZiHykqMZoD7KkUgM
B5eUNBWx+pjfj2Y22P0AnYmxa5t2vgEakeoAdd4LRowqQ2iAAZzJp1EMoReJU8t2
dBLAJmKWkztRBLHc7/SjSs5+AS8qIZeMtXE5jIbnh0Va2UrhSrwOIrxVE6oZKg/s
S1Bs3C/MDf3lUblx1EwBh5V9KaKXZeQoSbF19wUqeTzy6/pKF4Dz4Gf0Bj57iX+0
c067oi6AkPsEcjYS5wF45zyPRdGkZf8bqFBtyNjoGV17Q6tNzG8eC/hedU8Tr5D9
bEUnYBiXLeIvAhEG/scRWmgX3wlP6Gxf0goBeaLxGz+G/rNIW9sTuZTdXvelxOEb
SViq+NTEjuS0nPcpygFYPfjWWPbwFNTmltCq0CeZ3qv13Y8hXRl/AIC6a4sdMkqh
xM+jP8DoyLp+by172PCj851M6auv2MIAQpqTd+KZwhGjBVt5qfWkJghrPXOt7JeT
3U5CgwfdbQ3IRTBkl3VRW3A6KSEq+6Lsi2D8nEvZ6+qDBjcYRKCkE+8PPc+gfopR
6j9Q8yj6NDyD1sABwv4/5eOcHx8WJZvxwLupIReS2GZ1UVAyBMxsO3BEZLwlLSWx
o9R1l1fYTJBibV27zLCm1LeZM3DYdaIHDQRfavwv2SQjHawklw1rO0SxQgLBtxby
kcd+BTtt3WmCIY6rKyG5rCG3nvhHtGGESmmZKlI+KqnrgA8/Dc7yuZ2zGYD/90hi
d/tr13c1tvU1D+zngk/IKjvZ0GQhZU7A4soAHv79CQ66ZBt52zmVvK0M4BafL+sM
cBOtrZH3TXvKPKJFBRpKlgZMGk8+wgQADdCS8EUvxUUHptT7nrCZSpV5hl1lcko4
exjTiQLbEqeAUa3fMltIkO3Po7XpKzvf1R66FzPxXd5SZo2kwUwPpeFlJrneeqpn
5wANdtukZ4/iCVgUjIAt4bXIZ2Yr52tgvN/mU0YjLqAZJ2gXl7BDjvOeNEXt8T5k
LelG5Rv4jWImCoQFfWvBWdzqC8MPS2Kgk6BsiII+JMNnOkpK2EZMHZ3ickwX4pp5
O2euRZmp+vzFrvw/FxDQoaGxtfFyUg9aoA0w1dHLURBhGW0ztLIO4hjFPawg4Vu1
jm4u1iCXnaptdw5q5J556RkQhCmpfkZ6620/R1thSuiZSmPYD/tQcaiZ3t4by/KZ
MSBWCQRWsjCoRwoZrDvALlgyU/+lxMHJINUoWEUcOHvRwD6rl70B99SuaS2Umnfp
hajosMjG4FxJZozu+ccrygShLfC/lsmrDZwao8ETH4z1lUE1aFmqc0Lwt+Jv2RGV
deRlq5aglu22+GlOUjzkHluERGApsimLKDuTlxKfqi1JZNJ1uJhCJ1oB1VTEMTvG
taURx5bEiQRLgTOIJuPGprlAVcFpq2sXWiwr1O5yzdM+fcokXnZnWtHzKPrS8jrS
VzqaELAikuFX1FyEBpDXgFIhYvXP4swX8ezs/10NRfo8deJUoGfDx5ObngcPLmg5
ci7afvkakbtsPiBEVCa5Bj6k1y0/1yUOajifOosmlb2HLdiwpnxY/2P/kjj3IhuK
YpsxWWwmhjaZ4k/nKNsZrkjFwYInNmIEnODS6r+1S9s+omBlz/bIvQ5LmWjDMDNI
hOkhGg+Hbikj+ZL//L8zgMBVrqBrL2UusHcHEZKsZVAPLQD248hV7FySvxfCgF9W
v7tPXNQH19/WN+ghvKZEgXCHuuDgfFmqrVZbKjMsZBFFjOGO09QQmDWAxSH+1Nvr
wLv+CPoM5XJQVgobizsM5KC7wfqeucA+qc7V1oTNE4D70aets8evN8gERxgQAM2z
bhU1QC001TU/YZM1EaqpN7dE0ZvKMYnkx+HHxQ4AaU9K8cL2QHuIW3ERBwuHoiYR
A/28Q/pponNbi+eUJrpHmeeNUvir51PyDeKdgpi8CSTmOePAaQUiTvBKqroa7smG
9QlBjGqbg8e3GkSln/ShFN7yFEfrI6PDHL/KLY/ozXuHLI5+T6PMx/fijiEEx50r
/fJJiLYrwLRE8Hrso0U41LN5CuVk5Fqt6rMSejFK+fE1rGr5qqZ9InDWjpTQYsWw
uhvWInoE90nYxX2I9CBIPT7Ve21eC7YklRulGzrAZECEKnFCu5k/6kOrI2OnIYDB
so8gf6FwQv4X7AeLo2cscKBgbs2CBaXutTeax9aermjVapubF7xWQG9FMeXGbvKx
vXiAyfIxi4jbRX1pnuyKDTA0kLELnqOmSIrIi0YYwRR6/rezi3sJ2Hq+KG+uOU1J
GgdqOE1mpQ16PRzTM1uBopx8U7UoV7Fiy9FfSUJaAjcDoqeNQz97VvqEzs33N+p0
q/molbQWFgIeG3rhQiZC4EPQjupaqzS1dyYTxd0jxlMlqa3K7l+X1XEp5LGVNDDP
MtGTlCfiONVSvGpJxWCYBnMzPRmLgCWCppQSxlP7D5m3ZyFGIFdk7v/Jk98iGy+g
De7hgKMHzKuziZFsifOx8+hmaSWq6hI8E83s9VcRFFe23642me+GTwU5i7rJSYvJ
CtD5EjAPeEdX6Sb7tXGCpjDcnZbDBGvYpk/gaWU2X59rDA7QqVGiWZfOvxl+QH1K
sY/4Evz7KXkm4W7A8lyksJ/QrT4kkD7iiDQsFAQcDH7qmQ7qkzy3n12xfwkGmFUv
qUgrFl1Wo2LUrBoMosnGDDMWbMOPPctX6o9gFqB7c3YHaY2sHCNx0qP7b+YR8iCl
U1Y5o4ItSHQaa3ujt5dF0QoC4gxxtn1b/8KMxgrVBrT6UTRYFCWjmFQCusWWVAGj
3O+zEY/jW1pqitzXge/2SUch4HYsNhX5rUAmwGOoCJ2HULh/xPdte8aYDXrHqIhv
84B1QL8we9Gq598qcxbOQmtAy2oRCs05vXDrC2Yt+53sIWwBrI9N3/3O3am9lSQM
zr7SVs7tJM7uPjDE5VCrLudXfiS8nzqCtHzpqDNgXDAzsbsOHSaUcr0ibr+WddTq
dOCTUwDW9aUqJzIix9pRZOpwZHOsl3YEUzzlzgJb54dOQJo6stVBW6ohrnRrL+wr
jBvFL6nL9nOBATOlswSI09jWuuyWCge9po19yO+FJP1Gp+xpC31Ej9LrwM+WCw9N
Uaat++GG3vJxI3oC/coK5S7+zZbXcQYZ+DkxGI0q5T5+iK22jUOl0kGQq9FDqrzO
Wlh2p3twumfYTEqATPcSrEvTpuI64hKbvDqb8ZFZYR9XUwZhhIKaTaQVF0Ul4GI4
wTBd7QyC1gHf34A4F6MHYkt3pYUuTimftJqRhba7WAA0fIX06NYHIl3uCJLxNot9
bizIwXIqpy6IpAV26w6WMlWeb06ykYzq/NhekHzK+iLI1MfEi+jeRaLOU7sAafMA
d5WXagmMcmMJYBgecXRCGRU8zQOKp0+8VJ1xTO2BNEnbMwew+8tMZk36x2GqdmPe
WA6D5fyHwPeKCF2uKgxmjOk8niKCLamhqhkQHLQvsfcipN95JmKx+RUpn34N5c/P
Sgl8jpX8KOJpWqLxCjb06L7HAvgjYbNWBlc0V+xcNEcMwWV+5fXZqncpDQVqmiqC
E3ywI/OAzKmbtx/CGPSvCkSXokZUyt3nhZ42lX6Ba11y6lR0u2UCCQaRmuGzxBrR
8hgZarfl6dT17WG+ZameZfcvnt8SUaWk2lXs8NrbTf5F3QYll7srJLJU1+RlL+te
R7VLujt4W0/ZpLUejWXpOFcJZZlzFTqTvnoePoF8cPRzqd2PC/FJ6edoxrR2Llc6
44AxYl9AFVdxxF2N1/nwVilIVE/okhyZKqNgWfnsygZVCctF0b5kgllew+XqkGFS
W5rPJAZ2MbjFeCjxN0e7JpvKyF9KoppjYVdF5evmFfntvIIyxT81n7B+Jd9J4zxd
g9YmmzkkPmcU0+OJfbc954kqqTzHUECsTDleNSkcHih7E1jBo9ZtW1OzT90ThP39
vdRnfXt6+h1WgAizvhoVpfY05cP0Cej9l4QhsYcBtDtliGJA0aHjbvC4IR0vUbeP
XoWv/9qChw0KkPtbFom+iY7YVYdTa5ZMKNtBAPJETq8k6IUZB2j4geUwoOnjRzFn
oXmoMLCNB8zirSKV2QvwVnjBW1suyK4/5QUiIOIpJ/vHqCovWC0giWpXnNdVl4t7
HYhnkOOUNKXloyl8jhHUBxkIsQuYnFSYB3rYGoKA03Fkvh3BwKpxHCng1RXzHfmO
VfOxo1dEeocXdTMyW2QHmHe4WijML3SxmcnRbJMo0eNyvd+VAWFQk7nbDMnCr2k5
1GaoL4VMwS08ZKH+RChQpkrYCdWxPM1df/+XyMrailaoTGlhpmfVa0tFUJRmsS13
ntKIsieXxnzO1e5EdQ7jQzqXj1Jvm8bvx5VEbVeT40mJY0v6IIRWHW8LsuwXINhQ
dqVhhrolIpFuzAPgQ57+TRVblCoecNRZa3XxVW4j0HXkRtFWDUR1VvHNeu5S36hT
af+aC3543h59ZvPLgKl9X6Od4oMKaQo9d5EC3xSIU0/nuWRk4UTF3YkXoxNKwNkG
4wNLtwaoWg2aGtm5CBcNaazAg7FiKoqebKosdX5TOl1XG5TXbc3HxA/MHgCDL+vm
o+N+ObMTpVmSXlPqW54dvdTgYCim5m0WHgnqLnoA0iVaLpnc8zKAJ+p5XKHCBiqq
2UBbPs4qyHVnOQFsRSF2qGexW7RRfNaKtv+J4lnQiLYCj36WuX7ZeaR8TThkbthL
lbFcDv3SlWqC5ZtSSZzPZWhYIdaE5H+oHYo9xaGj9HLMGHMrxbB/6gO7Mvv4FI0e
0tbEinYxaKnbV5OmIxbqWitVhilghKQmCX1OSCsQZa2QupzlKhAhvuF49XfXMenl
0lZMZIkDyBXZOVdhrvQBTpkIXaKzbiKKRgVbBRs/Hb8HaNdVeuczA6Gcrc/UuYIx
v/EE+w8JuJPuG+eG5akpLV+7JunjMvW0IxYDsN+vrc8ZyqsDQa6F24ZT8zJcwvz5
OkArWCYUq0mh0pT/y+pbHDEebKsKxGyW0f2OpYNFsSiyaXxRwktJVOc+ZBA/WPdl
qNuu/WeDwbsF7SNoMgKV7CTEK50ZTatTIB72AbLrzfXmBFWdW3dJ2joDfwZHh6Wb
dvnErxfq/hz3kZQb5vm33QHrZ2A6InebHaEbmfxBQKu9+7EmPCFPEI82i5bBiczN
chWQDwCuk9vjTCfHKgKm9DN0tHAqKLOFp2tyqxBLBEbgke5VHAkOjjAMGvzEAT1/
5iwXyNZyEgkm9eI6b1kksazvrNYOleJE8MLeNqlDXtQuZVrA/WBamYWc/IEw5mGx
fPASEfHDt3akYa52dl0+MHTBf9DVHH6ulaRdqpp1rQ5BvvfdROuhO7fwVdjln7/5
A9bMBrQMQ+UUkNop4T12d1Q3rnDGxd5d3pipz7NHoazm0JXjyJ7yjD3AHhNyuuHt
aM4Jr/dMCiISUgmmLN/HbsdQ6PoOyDSu4E1SZE+qKgDPZE7W0MiuYy8xvTthG9G4
7NOfiozVOUBWpzo2wyEqW5tszE1x5/1enCAQb+cdHmh5dsLB/itE/aLFqeBcyeD3
Uehxl7SCVD+XRgK+6Ahb4UZ+80QI34xn0EbWb9UmKy6m0fSQQwx6BwZpj0JI5Oyi
rI8SZyYf+oMd2u1gIKJudeFPliO9F+Ea0LgwdN9rWUFfm+bEKh/08hbMc2t/sf6K
lU3E1fIL4WM+2df7LCc/DBbg8fNzkJaOAN4495GBNViBnLkm41IPlGQSPYMumkSJ
6PhW6dOmMM6x036aWbyLcIfqdRIsi45LMgnOo61B3kWwKolvddIedr+sa/ZMpCcY
LYaH94OJSKPcoURKfBvhOjPDSzGZdGbjNLMG4MOWKcuOyhHPhYFtEQfLcdbAVkrw
O3q16CTXiVYfyPed2ItTTfHpkgpJNPf1RaXV0YepJsGt5X7ycYm4DBDqFwZB/Ixz
gmx6QFC71OAP/gYiHhlyGhe96MZg1lQKk8i22QAuCwjWZ7Sub0hDYOQj5oDy6tGo
MFw9FLbmuy05rb8ohI/N1MKrNqN+jirRUKEPsJmYWlhPcq2dmZVghwG7Y4QsY3qx
cXi4cxkr0hm59MwjSTIl8ddTI16xYhY3df1rZuzc1PYSvuaaG3QsRD6y5/OlfpoN
tUZpaLfP48zWXMBGjxOKe4HCYQTmdLVqNirho0SsiXLEoYOqedxITwP2vbAskUuP
IXCQVOmvd38smLJ6BVEPoxNMJZBynWEEmkPjTIV/wZpajHMuVk26yX82RMVZNb8X
UO5QxUxazVlTbLnW926pLmcCWYWEcTNAfNK0ylut52QBaUEGwnbOVJegnGkJyOnI
cGrVKEbu3jghJK465FioOeyUSYqo1REkfeauZQKjV08pT1uaa6zpgb2ohvrzLNL5
zju3IETnAvP15FaTL29peWE6fSpVGmyZQ3Z0YeuOKwNi5AILWfMgYXQHRjdAvK4O
ENMaq8czN84qEnVuWGxFbidttpPVxCdIRN4I/liECpl4AJptRdMPI7OMIHmPW5Z5
LK8gHTeiNmStX3pJF5R7bkBnUdTJ7y0bTKS8cge19+ALbs72x6G3/jQAA+JFrBKB
yvKxN+Wu2r5tokJH9dsUvk3gqpi3K6b5I11r9gIlAt2Aa8WN+E819CSaMbH1TL7u
qhefbuLsOZuauSm2Fmb8hAzaCZYWDRnhMB8+qRBtszNYhmxLYB+mGglENZoKq1mD
VRL6EOe1XQWandZi/sH44SVenE81aCUiLzzKOCVcYCVKrjKUYEQi1w+ae7nNjp5A
9+fY34hCLds0IweNS4MxFMO3nYlrSRqqfiSrQMy7FZ/paeso2YsXrnMLs9jh+W2W
QyoiayeBRQVHclixeZhgSAvJJA3P3PXvZx0XfroFBWqBIsJ/7IGb47fUE8hhVQx5
ku0dBoTk80JbMLYpD3fzK3YLMtP5IiYY3p7oGi5OFrjafw6LSnwnODiARjoXBH9v
wHP6hmMUXpE+B1uf+0rpr6hrc4a766Clnaiq3XP72u9CJi+4sDzyruhJ+9Q0wmNo
mnDDfYVFB+8FD2hfJJdk+jOeeyrtq6vehtZBGZ/jPA5urR+/Tf1j43FszJ1/mW6b
ngMnFMT90CSILKfDN2JH18/KeE/yQNi9QhajDX++EHhqBDIyfBdWDirmPoDMuZkh
CwYnQs5aamfk7GD1kb5ACPl7oSql/4IeqYliTTCq1R8zAmtTPSjTIJarrHiHQE9t
fgAqGtkvDPmCXqnOmEUJhKtaF95FdOeYr1GXvCrBqMndXrrpv1/1utpLfht7jeOt
WD/xS8874R6MvEHrvYlSV2RNieeZst7M7yVY673f5cql2IYraGAUu/4RrtQkmRhO
2YCQF/m8N0mE2nAlJhKwLYtxwqGMZ3mX+dUn0AIUEXPYjPxF/7GIvRSTiAhS9tVm
QSMTIe3+9wH1dKLk+BQH/NlNLf+XiJHNBsbsBhyScq6mZdpPvEJZ0o3kGOnncIff
Zp5LVRSErmg3vh2+7RMsA37iFO07JLTwWrsfw9Xvk1SOi51j8S+n5S6EImljdgj1
zx79iyrnA+uT3JrbfkWr3eWBRaT+n2ucgaLU6+hqZ1KuZxPmwgtNUWBPuvm33Wmc
Ko1ysLRIAYRPCUqPVwGHCCzlC6CdzSgwHCALouP2xiCEm5uinvk2jlLjR7W4GJqv
gHgM98u9IpPJ7Qe2ZMX+ZUqpVO0CdL85PUxQv/TaTQmNRSJYInkom70xQgi1erUz
Krxrer3XoU5+JbWOyvBt3lQqQ+re3Z1dW3KhoqiDoWnGnjg8zIHsX4grzBV92s+p
/qARMseK2QV7aby6iCJpOX44HWT2wAqwhVMgzdVyw7hmbGut1eCyg+USAoI2tadQ
1yacTZ7654GfHOcXI8PHNvB+y9CyGO4q8hNMcfLL7bGxovYLAsIms041a7n+lzT0
q9qg1Ma2ITiuijCHz8yuH3msPeZD+QdtCZst5OIFeDYL7otF3NMLKKQMHgBZmR8z
7zCtBCK0YAY0wGlNIf1ZDW14GXh+pWFSv5pI5WneGdhtaHVGlpspZSwMrRwx0MAF
pjKkOET4Nrop6KfWKjk7NI2L2CXVrc+3NCQm7oMxnrUIlTGeyBO0Ce5V0aIynnuN
/jVO0QWbq3m37PhEB+ZVkb8V1ovpmebU2+pVq3UTeAPWIxuy/1kNUy6USjbacq5A
HOcgj8OyvOQc6jfaGpBOEj7Fi6RNvboeFkkzwYI+7HgGId6MUg6MWtVHz26C6Yid
DdxKVRwmMwRL5eH1bznJfmAOnQ0Y9Gii6/3ui1rl63kXRYnIMoIolfo7IEOsuF/q
LPCT9saUi+zRZD4FzfAS8PJT2dov1afTZryBZAwdmnQXdGJ3qrGBvWHVpSuqJo7i
6LZiSwgTDNyFQSb0mgfEcoJqaV0TCGpsleFqlJXq+23Qw7jhWYxSos/oxH4jNG5d
vIndfHptQehMxTNwFMRj8TOZRojJ39tWGZFsj0N1Mp57P2b0L91/AfQo2iV4uz/N
IEZVPvEunH1OTPIwFDjvYvLrMZ4cFy0pwtojX5x+e/2GhsiKi3akrt8dszVvlTnz
SG9Q+xfakSzLA9/Uw8Z1Yvpppc7dPf9ePDMMKD5PoMtHAkfF5/Pzb/GStlFmDKPJ
8nhlKAEoPmssAGf9DNNbCo8t5y8sEbnxV8cJaM+Ea7epxod7kshqoWkaLeuERxE/
nSz8md4pV1+unlmLRkDyDemaAMIHs66fncSuwVgvM6kAqJHAONNszxvhNUAu/z/Y
QFQ3+eZVx+jLflAiOEi8l2+cFwX/xoze2g/APJso5bpgMq2hCKe5XANLrTMmVZVM
XBQAsQ0XJxmEa4kP8SQoKnZ5fRip8oKih8gjVEp3kh3LOTZvFx7mHBXackkPi+ET
9gJfZ7BTUx8mNwFZpcsy/OXquPhkgBWIUY96a2IhXwjXJNJYSR+BFqpwS941phv2
/Nvb1tQmo/G/AImfZEiiTTQr9K/ZxfcLzhKzPEh3QCY8BX9HBouif9suuoShRsyS
6QorYnvAnzWJecHxAPYyLLy4Z/kOjoUoalLZZa9kXT4UoUetbAoUd6HOe8YZMCSX
6uRxLAFlyhR+IcE+4rDDAIpgQQh6XSnq7NLieKWcixc7lNboWklydH/b//ebQl3+
XZhTEVY0BW5hHtc8MwqL/+zanSE886OxjDU1HUeRd501mNLq737NEe5g/UFzxr/f
L9YlBbfqa0vmt62voRYm/y1USInsx3QLEU8mpsvCPydx7ptGYD8KvkHTiC0Ih1MK
lnq2WH2Ow4aGI6XTn9nQCvdR/JR6IYPtQJHCZnhTzfEmHmJ6m/R1AhYeXhE0Z3OZ
4ixwKuJOt2+3gZmDX+RkhxEGaqbPlHoU7eWJ+8EvhxGlZ2SxOM3xg3DN5BGUsIKJ
SpZPiNhYr8xI4lXekAUFWff5/bbRlN/JZGr3O5kzY0GvK0rQBG+6tJcawIPEgm9R
+4j/jCUbZZMTnd9tp0y0mV9bSElEWCapiPdXIAAXu6xxuwtScjipsJIjAeN5WZzV
1W2Kskvkt2RLOHfsR6juXKFQ67v5bwBupCG1jzQJnBpjF3EqdeWJ7G6474kvwqUp
0AshAtp4RWABDifnwIE5/Lhjv9kJl22JEegeS7OnfCWi6SSPh2A+Qrr2LLya8dq7
iZlbqNZERgd49658bWWrvEz1zGHNgGhpJTGnd9VcTysE+zYuZG2TiN4GonYKymx8
Kg69dot4Xu+c1a9mqxUFyyqyBIM1EyCbpuUCLdseVm4KZAXUxgkBOx9dx6l66CV8
xu7YBCXYDY0RtzlTqQjFZkHWKpxXSLlaQWImshn+JitwtxmGCJ31X6C9iGDe67jd
UaR5GLkOxgH82oOuq9d8Dbdq6qJpQd2AGeOHv/VMdBXEJS2t5NXIkZAV4yAcgMiE
6fm5SDdhoB0xzViTs6+Gm+XB2dq4ZOE2QglvEAyfyyUYBW/raPzyYHJXzGax2Mbc
WXTeSReXfQfUSivhVA52RU5u4FZf06620HuAEXwHDktT48RIQesVFf14tSwyY8O5
MfB8r+MNnUxKbGOOqybbHQ3+OjiKnW9lpbGz8rotaTBBvPBeeOas4Rh5xZY7oS1H
I3vRP1geAyIRhncuQKptwN7nPrbHgjzg77W7JCQ8T950P5ST5Z3R3WSi0kAlD4FL
fnpTKTm7kiVVdLn9hfP86qF85/ysSxLtn3PNAAsljCHsWnSuU394LbcilWzcXN6Z
0zD1kbhwU68EIL3nbCxZC76cGhQfPz9L1HsrtIHreNik19U+VTZqanv2fMbOlWEf
7qqTq5+5o2sQwduPAZHpRzszF3CgZh4Gi8kfCup1i6Lv6OvaloX9482b9mt+mGGT
SG5DvXa06HnyPjxAeoDjRyvvvJDDLjeq4Se97hl25p6s0RXdE6/lM4WyJlXR0y7G
BJ1cAKoD90qMlOtcWyBpi111bEwpPgwFBBPmFF87eCAH9nEPlwDR/YsGIM5/PrA8
RNw/LRSLFZ8QsfdQlzFfyzY9MMFSth7VEiCIKrWboMxAMokbJRK1CVwywjZ7L66Z
aFikCGxRxC6C2vt6DRa7xiPH7NSkb72NIffZoSXG4/u5oc9Vo+HirbCl5no7zsxr
O5HQptQ0irAdJMXyDS2SGKtx+Yp8iJLgLV0WHuibcCKQgD3aNJb5GG+2AJAjAInG
cirVq/pFMpCfKX6HBfj+gWH+yABwqSbQmU2Qoh46d04o7haFU7CR3Ls3rSynNggI
QtcilDtVI88P+LGFv08mxXI0reAeBxxlxm8zRca3B85Mzdd/YHndGaL7thrzbecN
XfRHaYDHwA3l9QAxfigQgYt04gdRyaaNGsgK8MF/ZfXQo9nr2tEvD5OLJrg2zh1F
th9uPvKonmjz5dhhsdJTdDeUdx/aZQwz/7Q8/8AbeWBxNrIBnPDSNNdexFR6y9fq
mILkUriK56fToHetl+DK0N8dkMHU+vowlS4G8ypc5qBhIW5UGE+io+3j7ZQWQ9JX
YgWNN+7gdm7HqF3ccjYBnK0utgNW9qE+WM1fs4cHmwe1MYQ+XVLYDQkH+rUK8dfS
NI1oyr60Y5GWyvAqIhkzJMR72Hgsx3BuTiGLdk7MZLTMxbtLDZU1ydFFihBrP0R6
eQYbSpnOeHaEIRTpVV1BIju/6Dn/Z9bt2wIba2n5rCcQ92vlCqCbEnswoDnUqePe
JXtxR+rBrWt9Rr97HaRQADgRZkdMz8047eeLV0xJDoeFfl73wmozUfMD5FEnWWBJ
6ZUE3jbqVpfW9WyylWgC/NEgqwaZpY8OuEWVQyyNOzmE3s5uniK3M5ljOXt96jY3
Kq0K9RID7j0hapBjRUPcwJgJyuMI34qeVyovb/tpf2FO4/RHPGSZ/mUjF4wd8s5R
LV29jordeLiCUu3bBczLlJrXvanYjS/IENWzYmVB+jsF0kO+trCKZFEggfN80PYD
Z4AjYhsiOX6kkpn/Gvaxj/9ZAbwXsWYXOoqoMy3qAOD3ZprVaoP7972xwNnRyCKY
xsZMvTVlaeiTEGK9DM/lidWIgQ9qzd8fukOVLzQmCS7R+LyAOB5+IwEPf+/R7FUf
/e35VrWslK5gZMvQQOsnXQ1oMjnr3cvVvThUATZkDkc05sXIU7GqGxhZ+t0urLGD
NCi0H7HN1HAHpWrdtPIPhk84Sn3U434pHJf3WlMxcwIwx+KKYFVXvNCLxoIGl29/
vdjF0/CNgnDFHXxxl3UIZRb8cxp5IX3tEEUVrzRA6114roSsBRBDziLq+s3cLI4c
WD/H5nonNQfB+n3pN7oPEhktlAaRxyjGydn/GY8vsVw35LehQAoQVdvkUlmqvXGM
QTCCbOrMzBo+v+AleG+T/XKfSLmIcbNOOx5OfRMByZPFhfZTNxD63oxnbXu2y5Z5
lzANnqrxXWzeJg3RC3Yget64UdHs1pH/MD84i4E6Ex9jjgTqrp1K3W/s7efIK0Qo
aaVg7qwo214oxdJF5z6gcF2f0j/94AGxxZFjWW5LRQUo2rzZbtZpTDpM4HeTYumj
ZIZQ9lAmKlVtxkZ+BQXZnlrHwDxYNhlDemW0B4BWjBRjfYNMXAbPTIhML7k1Yafv
gs+eX1ZZ2MQfv6jasfFqqBodwtQy7chyFd+1scQMzF157ZxVVtrET0Cq6HWehal7
GgE2B6H3wSyYGhEKDkq/oDtgK6FPwpOTElFY/9tVR5CQGKJMsSUsQOkYIQcpTVik
OtnjI5wImrYs2GunOUQpSrUN87WHUzg8piXnfffoONpREuQnM8rlTDqPFNNNFVVq
IOXAqGlSqhLdfyM3XhSuzid8nTN16f+uo3K+441yhUI+E39ooKgr4f+Vq8LnbHEY
ZmKY7CmGMYbKN31XdhQbGNZBbOwUc88cJL30E6N/pKSeVQIpZe+NM2WhOOUMqJcU
DgICJEPeza2x6VcJIOcQiqYlpw0KIb2g+TS/mkb+icSd4n7jZyybCOL+VXgV8oyH
3n2C2eHxEgpZR53feBRat4uGjRiNcm5Z2hnD076b8DxzFC+VfHo83n1Ep5AUaOKT
yEMKBdHzk5KX7Z3o9T9jqpOcT/BqwZW8v4daPmERKdcCPBICqIzdLfcZj8wyP7w4
Sb+SLo4/XgddHT9j3KvOeBFQI8odT9ayoVYQuJwg6UKvMXmJjBC/BxiMV20Zs9iB
tt3B8mPohj3Fs7F23/RUXRQ3zPr6qJFaG0AL2el4OUGkk1eaEQrGAaWXVQISy8c4
5cZ+4g1+To9NVod34AR+HHQ5vZERhQvNbfHRcuw0gGoJUj4Y14Fz9Wa2huG6zoUN
atxyu3w7J/VpllaWyIyX6otKL0eD+g1M2F5KhmUr4nvlsGBuv2ybHStZ4L115OO8
yXY8DioWJbeu5mKLs4TBiNV1+iFr94N0wr0RP8aLORru6evT7U/0zi6tVGgJFPlq
IxfTtXMFGLBrMAqUiYKoDW/+c/IJfaS03bQ2OgfIab487uMB9LYY567uq4NxhM/1
Iq+nHf1X69ohR64tPfCakBwu1lvdgfF+rYQuYfuloE/W6RB4JBHY0WVlhbU3R6/f
d9+mEkPUAZcLtZLKvsIzbB//Jq/5ma17IppwwuutjYu3unLuFmTjyj3hplffaw58
KRIJZdunsq34akQ+gnl+1qHsf8Dj42AnKxgIhr8jXV8i0CWwRQgUq3AIt5/0tgHP
CF6kJ3AZwSxOLlF6rPHCjY8nSuC2vFA8XU9w5k9xr2VX1NdCAEIakLBJOWgUjkP6
PNSEgqYG0kFKVzwEl1Xe3AL7/pxHZ/uqjMJ+yKhW2JNQ/qopNl2Ib30sDlD3ewos
kuBkukyiMdSNGlcDSathjtagzrG+3XzoAeWcbs/FZyaHNGewhC+3yW0gGUMEF2nG
csUguw34bNu5IDROS+d9vXF1Da0dIvaCHX8Pq82yXK8qmP23569N6a40wICnJvK0
/uEokn8ZL3Bf+AcTwllFQkIIkf272kWd9oKOJ+bALaET6HrL4+7a+JrNLgChPw3r
hJ+0d/TVos9SwIGRXjA85QdWWOyDDUuzhTzpkoA6U+uEgdFfFQuw139d2bt/Inby
ju7euzlHjHKp9/DMNfocFvB5MffRlNXoJrZFwokI0cCGDwjItiZXQwgpSqtZIl70
Pi7vVFUkMurOR59fovoUaVprWi9Ftb2TUmNPqK6F93TxnwRuwlNtDDjMKnjLmB3o
XH46/ELgPyT+jtrOzP6F2xlxBiHtWNRUqDnIFe1SE6E1KEQgt+vdyJvJgtTI5nBa
d+r5CnJBJ/DLGZmvtjh06bCs+q2Y7flKoWI2z7HSKwL6VVJQcZf6CGopaFc/dI52
OoGgX6DWOfxErCRMtrqFRrAboIrByq4niaxZNJpIvRYULVz1ayzrh15yCy371cGi
LIXf8a4UZTSY0aXv35Lq24seh4fmDpqSSHq0SGYQTPcFXdzoETvnxFnqOU4vbbqk
lFc40DeOlA5GUV6VKOJ+UJ/YK0i26Cwvonk80euEA6XhgLsI/884rGPLRsVWdk9o
/UhKCUb92BZ8FQaJDnChbNLKJUycjTiTrbLnJwD2difJA1oRDHkIA+8Dx0Rff3z5
hb2DUpd4GltJTsfChi8Jlj7L1w/dB66TiWqsyB9N6XDLVK6JtIUqt0d2gSip9plK
VUtiO/YTV7Tb7BNvGNLKvccxlFKZq++pQPOtQr9BxK/UjdXX3fodoVofYc/kPE83
2wJNLv30GWAu+0uPm6ulyA0nJQELtymuC0L/vwRHt1dG2T8JwTIYU736a/ThwZra
88UzgFaE8I4bK9xJ2ZF+Ym4VXs3zgcbaQHwmC7YbTdlLZPe498piHKHsSXnOZbKN
gPITP3cIrI8uwGVHOUYfWlKDcMlmvjrYDu+pxXJP9GkfRHhhiwUmOl5/MTd0+E2k
psDuYx2GNhSP4NBRCYjkLlJe0/qRRQjiAiezHHcolw9vNgYkbaL8Z0xgEtPGHlV3
AMo1zNJoK9JgwZrAe54pJmXbo3nBpuZ+8HF3DaSQFQk2JX4NZpnvCDp7DYsOfUDu
O3Oi5wEpcaKt1TxCEBotuevvdrHCuZ9XWj0Zx6talDSX9rWfhh8fHf1WDQI0677V
xUQNEFkIo1rK2yXht0RwPMftGXDo0HjQTuArIX38giJe2Zek6Q7jOaaWbYHQX6o+
txyZkF2ObQyio6IPsYza9FG9Xo9mMlSNDQP0ZEAgCJnhAcE1cmrlrKMQDZxOgAYV
GKKbbBX0T0YT+TMx7gI51y7GB87gOIpgfWydpJIGnRlGQt9ZA2Z3ugoJPT4XjVXp
BMX9/h0QooLMKm4XYuEJQ6SwXCgMipbTFR2sq3mmZS6eJHL+L3fNLZc1Zd8A/WWe
jU760ZWQzhhpnyX5pXGwFpYd/TllJnAM+FPIWwiv7hNBUZg8iD/mQBSbvdbumcfs
QM/804CZOhu5wzLNrvHsgm2mAzMRRk4+zVK5cGB+O2aTZQiIXio0Pnl7QGOF1Sqz
R25O43vb87tY2d8q3xUxO5BIJJkAvc9FHjPdlyJ4Y8xjriEBDu+ntsCcIxCkuQWr
hiE13cQ5WeXUSlMbYoiFPi6i13InnQxtrxhfv53da3D2Hyn6z95n0BdBxlnSamVt
dqjkZqFVy7M6IcHxflR3DCwsna1mBl/p+DJzHMySneGMrv7wSNHcZoC8juVcFtgG
pA5ylh7ECtyj/L489E3GNXhcOHvv5hFlJmXLdg0YkxwrVNLiNhtMJmKv0my/aU1e
HN7s4eFphNSsUEzGscqLt2eLHW45qkDjUfxdC3l9niMRU37VgsDIkh4HgRp75C5S
8aLOHeBr0Pj/vuFAeAtQYuH4UfzKouIAjeRgiul0JRVTDMrGyvWEjZ+UfQU78bss
Z9hw+5/mwy0qwJkkH9S5oEXf/soA50BSf2GHY3CZ7UE3DDVEL4GJvs/azS7rHWkh
wl9isSy16lX6mGkm18D5pjQQUduDeN5QSL+sTU/3HLGp0bz+aYXB1lGOEWqPox6j
WGph1OdruOuujwsZIF7q/o5WFCtk1zAB89Ep6xB8KjWsTGB2LQ70VM71keweQoZ7
lR5BC+nW0pWLSX5y8juyyrMeclsoeH5pFeCX8GjSaBuTTI32KaUIOzy1k28JgcQO
Z3yGM1/LDb3kMygQkUIcxM1A+KqU+lqwoR05294f4BLu81aRexCo5Hvep/GwIreA
r8ni8lpGDQ8ZarBizQBKVVrip0F6yDtBj1ABcL+zGYxQqOzE1XwTUpJLXzwYh9i0
QpijYIl05kau+PhakIcFchYMXIN8ZGpC+r9KIYBBkJkb8v9c0Np3kheZkboQgID7
0PMX4+Wnu/QcvHyM8y8E8geef+nv1MIECLqspm2Nnaz65dWp8TCPVcWspXK1cU4p
inKQEI1Q84lku9cINIA8VciFtH6q8H8U2Cdmz49cCXJeTGDmmIpdEXmSPFwUMSbP
837hTdVeMggFoiNVu+oW3pRECr8NqnFTa1AxbnE7/tYJM3YHJ4k4cNX9usApdlY9
S9tRgBjca1H+v1pyXniZqtaTrID4mJysLtODIl88FAjcvJQRe0NMoa/WDDSwJEjb
DmvhuHt36LkX1wZC0rV/7CIJ9cqhJx1kkR4c9MOjvFqfIK/NYArA7dPWpXtfV0Zf
LmW+cr0FbWWHOXTuzzqsVNPgEa91C7o8M7+S77Gusu0nweA8APeFX1dzH+yFfh2z
Rr+UW0yhC0SxsdSB/mrjxhv3Uq+kYwcXQzhKtSVERFeMA6WvXeGcilGSBi9rIF9z
ty51ifwHBAu+Q9CePRqci3cnhNuBOMVp2fpn2lBz40Xh9bwTTCZpfkj2R5DtDyjC
r9UH2gTmtIW1y9nkfXsnq9CbHbPJKbfb1mDSxnLFkFlVuW5e5/VYGB+QAIgUhoFV
k67YGDl2C6E5IKQ9lcEaKwX10AZ2k4dn/a5lDCh6sL2x/XdY07NPA13Mw6E+hoQE
rZf0dyjCQmYbQsdzoNBvo7pZY6/Aq1rxZFQh/q/+xvFFLRVlknvjn7+g2+i8Mm5D
CqHbDNIEVK0+FdVs+r3BJrFQDJUfXu6t8wtUBuBdLJCail/GT7cZabm9fZCM55Pe
omN1vlOnhngnrpcCwWr/6u1xu2bcEPXY7igvhMdZUz+S6u65l0BJIzEt0BrDPfVG
LTrKzwrhfK79/xf5wC6kix0Yh7l2CIue09UmkU26imyMGDxjvPJSvCjNE4P7jTMw
v67X8+Cfi0Gy1+oS82his4EsxEgZAYprHQ8n1kVcSMWm13YsMPSc/pQT6mB2OSDk
L0gbH5C9yknN2T7zmkb5VvCjHfT7u0LwIsRaX0FRPzWASxWjncEnxTkh1VXQRjnS
Hs9JUh6f1SBtsLNVT+CTwhQNDB9DCtOK2e939p3B38Mha0S6FlHj97aIWB9zwa+u
fUm2EoPov0hKF7C2KQeICB7Z8g6fffju5EzNi1Iu2+qFh3MQXqpWShe8nwofVCVo
JdkJbObRLQe/BC04J5eLbtBC5r46Xpz4OfQaQbANxurLzyf+kYLG/5MGerdBtj/I
8VMm+0cBPFelp+pA9HfDoT63wDkrBs946KFGZMnxd7i/JsluiIz+hkup5dwXjbOs
jfkcl4u9j+shyxtGYdbRqCTLQCC4ZAxUfwWkS9Uy0hL2PiT/R/r4WUX28BMfVt8k
71HTDihbS7P3oChLqc7UVa1wCukaXKCYnqlA6qkGcymeHHNn/FbMPQagl44Mm4FZ
jJduH/6uTpclW1vAW63AEb+QRIeZuj7dZQdj6cuPniMxa5Rci/nL9I4SFhdqdSbc
cBdXGz6QVbruR5BHuOa5khYBJViTvv6/P+cAUfyv/QgsQq4w3Wwf4sCsyt9quV9H
ckA3DGuQVpJLPneiYX3jJrH2h6x8Vdy0Cz9p9tmQNITWLT1r3GyKtU9ZxouTPj5I
mv5aYXjgX54nTyDgfL7MiVsABkeEnNw9kdF/0GqSCrSVquCx2KEmZbJ+kBmi+6ks
PUbMsL6i4CKr9/Ot0OLJoaASOeStRBEhihUPRuJTCXX/Ku55BlNVmfKgij5NCqXg
ZlWaWjVhyrCUVGvUfWq27pp/P0rLEasi/49Zo0FgObjpWlicolcUvZ8DcXlHv/4Y
eoCSZSD9ZGSWo/oNIBtdqR6VvdnrMIZ/QN55eddWRq28qjtDS/pxVprUfzhYAcny
+1gsLJ+sYQ4kV6BKYQEiIotnycsdbVHAz4kp0jxrEu5948O26eWbD90S4gUy+7xw
l7QMYdjx0mfHcMY0VzFulWycddqgcZtcf/lufajswZZfb9ZRxkbpAPMwQ9VvbLeV
px7uNOXsErhhoi1VveXd89DCwsoyqMZ+n1w9kJAhbGFeaTmVvwrPFhbeyzP105Sx
1Y5RgNTStSLiDzQ+720x0GIHZI8a5pms4GZOqUtaiD/u5hW2XbggXDepl/CclsmU
tE/4hc4U3VbYl/JQ+qUvvv21mugenDjuVs61Hk+Jyjz+rOxW75uSxmAzvRadxtmb
yOOORtmj9UhqAR/G/eW5aHKI4KL/McMtNrZVynNF99u+6REcOHYT7H8F0kxuHaXe
Q1YBB08WI6+6HqAqNxsPlo8nZD9hegNuvULxrdpxz5v76xuiir5avIOVxfoLWclH
jtpqp3RYgHUVScsywm59BQxdMUt/+Sk51JoOAfGlFyoClNQBCeN96d5X/RUWVghv
1hM+Q/vSvDjj/DTEIEf2YJ+dPIH00bMHCK2re9bZvH1K5fwIag0QHbbHF52NAza5
dVQxbITVB35ZFzzK+jDFk0mNmcljUdhb5wln4cb/2UzryYz0xCvR7Bsj+k5XFRcL
X14FA8xC9kfGUu+pU4U8jn19rbZ2JLmaKlAZhF1WfAAkNnNfkJ7GfRCCbrVadprQ
hnTOsvpEC4YoxSBb0/dH/Vnic/ExDyYh8kCGh1vLv+cJ/HnJyGVciaFER9NJPB6M
a2AmijU3IHpNIplCcU7mm2W/+NvL/Q0GySJX8PIgJzG6q8VDG8bg2v4j5afJOKy4
Blx0X3EGIGtH9JyZICJLaaxfP769qJnOFiupl5z8UJVbXmWRZokLlYtLMlqyhByE
zPaRszx522MKB7jt3D6I0VuYPJdGTyvm7G2SziiF1KuIMuZ3NQV9Tcr6Jz4iU/B2
HlPj4YeJXsvEvr9ysooYb8vzHTwDwIQuvnbo945jHYsrPDiZ3WKr9SwxA43fRjJr
YDEBMfniTbTN+PYq1HEPiBDjo/R1Gn2qKXpKCy+EQpMG19PgtraR5++5XzSQOQyN
JnOle9Ykhh2O+jpISN1N3Vr/GwZTjvUAT7IvVaUx2GmVgX52yNllrsC8p6L97JGo
tqXulHFOmgHzWclhs7oElWA3Wef/ytrFIg4m/IqgbdHDr1PCYMuVRSD3OZ3PC+I+
Ta79rlriAwZpw1Lajkpr2pwkf1LWPSQDa6ZukuJDAhu3mS8DZB3QkjS/+eRPCgQL
YqjdJ8GEChHoddVRk6sCsby+AjFn/RN8s+5LO6ql1Tr57JpThnjABfHko34QmHY1
f5ybA6f0iU8hkCUfAqDucgo0NL2XXC+1GY/d1SyRpnZQuCMYZUHW2O/4eNavXCOJ
Oz+PiGzzl+cq7NhstF16EV5WDcWcrud6gYgcsC/7ZWllO9Vcp8dGbw9v+jNNW6aN
xXPEsprSFc/rpb5YOn64nQyi5a1QkB689UTitrXrRrVWpAgrzdiNFeMN5vMGT7QI
rmCZrK5VxoC//11I67bAtNWsz/OFVxmAvm6Ad0AauPA021cNe8JDTnzwe81vSUQJ
XcwzxPo6F82gYpruPF8qKTJzTYd4lJpdW9bGdGiFTgqw9JJFegoNiUjv0ubnJUd+
ZkzF4LSHlzGCDoN49RDYGOSuAbCXfiqcZThT5fLuDVOwV/z0CSNx5+JjkpNo7uGM
0VlXo5LOz66do3Osx2m32ImddQFwgYXRZys7Z22hiD3Vcizmzoq5/i5BkDjBdOR1
+O0czMEmq9b42H/mhgbril/vaW7EiC0jWjZPKrvJOrG1JhOIwRWM462SpoWzmYWS
UTbKVeaUB4YitEOPkavd0jUly2r7rv7N+ujtRgDeS5hjfnIiOKKjy1kKaYllgb4d
iWShoMHLmFN8GdycFwjBt9jugvD3K5uZakuqZp2TuMPUy0ZUPvmBkX48mS7jI/A1
PXtOeWu/7aCbD8a/EGpufAzt1vgtPjDYmY0B/0LPl67AOFUrmYNMJ5OMH/vn57Gd
wo94IDAkBwg7bgqFS3IwZdcLozmuLBdd9HUpAoLwdWPG23v/CyOtUMEZdkUCPAYe
SIZMfkwbqyblDR/dP4d4LsZyqr74qYUDx3iYhtQrkocK7uuRAiOjoK9ipBQLQZA0
Zp0MCa1IJRStC+1f09t93j5SEW68cnHsKpWF1iXlftorXKMplWxn8KZTmBeb56jQ
vtR1Amb2jIDmmYqJMzd3QrZoqVYFtsXPsXkTDkjA86R+nN2I5ZH0xZ0IEfC9t0/Z
URpKzmKbd3AOV7YC3fbNjBnjcWPogcNa4D6HHDpXay3y2DoF4lS+4v45NUhosf3R
qYsJ6RFCs+tpuFqpow684C6hoRNWY5SzLGcGqMgcJQOII8VKnZdGyPPtvJEpJhaz
8v9Q+VRqeoKlm1QO9FSh1XWja7xhTmDvCvTCVT7vNeOhqX34hDllPXIevbiyCQvq
vlVffHGjvUnx+9Y3FZW0Gw2cBx8nE/+DYe8ZqH5VANDAGPtru8XjVe/jwaF2pFs0
h2iqQ0eBQL3O36VuV+5DAtBbk08WhDD5fG9rooL9Wo00Qdx+J7ZE/t+4xX9hFtqi
KoOiclqHNtIshbLHD0GjPwJ/JPcIrwFjZb2yJr8M9QMhYquOOgvOkIeIBnXbRaSG
sztpbIItgAg5RSDx+BeKPP4/FF30af9nd4Po87dYJ5rN60n9tXFZwDYfIhPJ2L3h
fxRDlaPqMmr1dMSNaAWl9BICbmi2DUb7/OJx/CGUtqS878AH86TSsj5LruOpTKLS
fnMfgMJ4qnPJt2If9I4Fc6BA4qSTHVMo2EMjzAxPvUp+IWtmU4fDH9HAXqDMa1JN
rSsR6f2fiKghgzkHOAz1a5CThtDoHHzhK94tPmQErdTuu4SCoAsvsEHOvEPF+yTe
JXiHbUMhwAY5tCoPdY0tFAMQdxRs8/Ab7CbDs+zsOj0HHRDrIYrqXsbDPBjzb5Gl
pum7uhxD42+LsfnRiP2HauH+3ABxUEqV6dm9grNV73OT35hZ4dMhHU4v1VMlsbhw
euq+iZdZk1hIavOazU3TYTqztVA+Zf080Ua6Qz/572sXbT4qbtg/zUBDYgrYion0
uxrcG+iiiXYWIjrxUfP6YdKpJpTRiMFaRTOR8ddWTxN26jHMXa7vaQAfN76pDXEs
IaO+mbHwmK8Ar3eJGMysn5rPhao9i63tdMmIVdInPtGZ/3xp4oJrf8qqFTSMrA8I
+7uEtzERZJWgb5BPNFgjjLYRDB11yqQ7l25kKVl9z8JjJ3ibxS9hClSdbpVbow1R
XFhj5GNwf5xGnnzLmMb5rKUZaU10fc0WDCNGfGlEn5HNR/ExLjHKdd1BXCaf/IES
gqmuCWzfF7EV68TAjw9+uxNUQG2cNIWm+JCvmVqj0J0RxCr0fd5RyCn9q0yQ+LwR
5Hu5AyTJcU6f7w+Ew7aGqAsuAhIKWEZrZclmk6rNXsizbkjBsqmGLwT+NxIfb713
7+BAo+KnBxp4GECAlGmrxR0TpNScnzyFKO7xGep+abaUaBsbTnIOdb5cSPhurhjC
fOV1F10keABD5wouCl++9/FwOZz9xaHPQtLJ1c7L9POd+xwKva3vrPipdgW0Q89C
RRqMh1/0a2LEbKxrEz3D6Gg+38X8OM5/RYEdjXO5N8ZxRlyGX+iZlYXBd8DnCSIZ
RYiTnN6Cvchz/cDeMCRHdz4zESDTS2Rbb7xQgRjOsP4dSL84fMLN10Ppy+sSQ0Jr
M6va9eW0LAzEOtFl8iGIqdz9sMThnptSak1aJNZLEN1YZm5SClaHgntCiMT6TfKT
DSlmOwsdJn/S7vBPbxZcbA+IRGAOuxZ9CXcLi6GaZ6ESLJ/21J1BVVhQ/XZx/SES
rsJfNPKMdRJLPQwavE5swg61EDooq4Br0D5u6A3Z3zB3SV+Rxo89MMWGOspAR0wR
itftqftMoi+1vKU5/2kaWGtswsp2PnEvPbRw8+qBNxZsD/hbLrYKaUrkjle5LsvC
4mIStaDuJ/ZZktASdGPBeKTG0Ku/4mbyqDYmTWvLyyeIhxYIViLruUzh9F1hWEXK
72khCjj5aQBIm2RYL31E5L3i8WLnDFxi6+icQpJNj2NJpsYt4HrpyvsH3JOxWJxa
MvS5GTXMy5Qq75OuBUXJcMkhu5Z17Br/+Vq43XN04OK8RAJalQzrGtd+AhfAjrCn
5MjNbbDgFiLzfy2AlL6rn+r64iRgDJsDqWvtF3anaF1itEC0kwdJI7tWhDFYwsRP
13cgJm9Sv0qVMSsp/d2JRztp0flcgyCgyZ6v3gVJtAu7SIW72A9MddZwWqVeHu8j
KkPoV5iktVbnXNLHDPhqGYNa9uGaEbQwk3SiCKXjNGvuyhTaC7QSFhvr/d5O7+pr
Ilqx8oaD0TEHNKm9urHSOjebU42WOAU8irMCETqAEGcudUS7fK+3kJ8xAKFXRPif
rf7mZDsj2jD13WDqoN++sdaVaPkZGQoTeDRHxnRKSoO2K1pNytRJEo/ozZ54ovS7
LRBd6J3Jmc0WHdSGNqy2SrpBrqyL5bJaJBxmHo6GWG6H33nSaa1DZV19CGFJZx4n
WI9/2Vl5KjZJom+1KZIBVA9P1wSX5guav0wiI/Ws7p53LRnCg0e942CKdzawolUc
OJxzzyxl9eBEr14M6ikkJY9LbaPkbGjHu1IXFUPT9wdN8QqwmQdyoypkPhmwzYis
XHoQYKSW8LoFoTrAXbXL8Smph5fe+fzderq713U7Z3NCD9KAQfIvZ+XnVVEtSqlS
36wriPv2WCzP5/nQ50niHCBGYbHcfWySHPjvvkzt13KulNYtvBkifM322PpbegN7
Y2sMsE2ZiRWTEC2ctWNK6Uj1VvjANmWK/E0Yb7zGZiGLz2aTJHO5ao+Z2Jw8QUSZ
HGs4wnDWsn6UwDSXcKSuVR0lIuKbWQBcdWo7AIyBf2dQ3rNEzHACK7jk4ieZPzyX
N79DDLV898Zgn/40ioR0Ke72d2DJ97HNvxjuNV7pfdkgj2uxKFLR6CgHTof9HADU
CQEA4p8Fe2F+zVvlGY4IczjCivI9+JqQ7urnJMtmV9FNR1QnZT1jp2RGTmBSBg6W
wxTPcLou69pQu7NrDzLUDxbBCvtNbcARAwdollvhp6fLXS9bW4x1SsLma1E/UK1J
BO3Yyyu9WUlO5fau48FgR5Nht5OBFJlL6V2KWZtZ61FDNdlP+BVlZ8Kx/JOPddgi
OXENbJdOF1WY0xO0JwtknMJ30+/XM4QlSaDdlEwnO24sRGBUW278G3fS3t1NoomE
PtrpDfldzct52zplDYcNv9cJKAV2whl4iNaOtMGkHm4jsVSFvaF7qiQPwen0SdX6
YoUgSfEpb4dburoq2kZeB2tCB3hcfhRMOhtQAv3ml9+SQlT4+ER0YAcTPexUYI3D
YeFnmTgIG1xPG6RKM+K9uvhnvCYpRcvAH63zL9KJgiOqEKkaty7iv/bc0Y72A7B0
I/UlmNWVQob1ETxiFshWl05y37o1RHLodcrNkwpa5W48mRgJ4f2iGNb9ZPXPVsOU
Cl/FzKUfOnVeMlozKoNQIkNp6TLowvA7xJjlv6pe4YOToMj5Ca9P41fv8+c5khwn
jVpg4z7EWp7PhQbGgcB581aKoVcqxUuEB87LxccgF02Vh3dcef4ElBtr78xi0GlC
s3dzolP9kIJWVpCr+gU5UVjPhwpo0xKhD2QWj2DtWSJVcvd3+Ayu7caZ0i6tz47t
oQ3S5rbr7mibs3fCBHwydlXPXxcF7dYquSZc/PtKYVbiOC6YDn9+EilDDNxsFMV/
3X3OTb3c67TJ70o4QZKRvU/jyGUOa7VJBLZqElPEjeeLGV7vXVXRpVMysUBa1ygb
ACkH1I1DqGuO3H/h+Ifv2JBiCZ+wYMxviOO3/0P4DUOIkeMQjYp7FUUYckpcneht
WdcAuBhSO2HNyl4m5psYBiZELAon0b1Ln+prhCPNhtWBREdFhvIOhjarSD7LvdtC
2AYvCndS1r5VCYModIAPGjgwYAjPQCyP6FUK3ghf/9jyBx7NDmc30zxkGqKDPdY4
UIOw4kCW2ezKk3FmQPu8TTXH3Jotz7ddBmpwIhjhmV1SxuJz7KdN9F+DXPiM915K
ixn7Ho9wiccNN8IzSKMaiah7wkbL8jqoK1piwAeKBqjtDWXJ1nWs6A+oYwEDLvxn
qVPYPsF1n7FYX7y/5i1/K6iYJ20LaYhoYXbLk3xiig6Lf0jo9UrNJqB5XCAdOvSM
ludAnaBO+cMrz3dy6A7Y+IYFUOO81oWp7hGIxo2ooVhoo9a4uvbpYkBrC/g87miI
fY6puN0H36ZbrLuF2MHJd+0DrPXPPOw1JvTOmLvbaFf3KLSNRyqpizd9G+cop3n1
EylDSAhi3Dy9VI18RKpgryaiVNGHM1jFn6Q4CUETENwv2cph1H74+jWPkYEUxcoP
aHpuVlImvpFDRv/iVeuPPxC6q+s5YFfEzSdxsJiyMOPiyEGsLzJZ1SSYbLquKqzx
lZeSy1rERy9qaI3VZ2mW8DRIWbeWGVmtHRVaZJrvEOhh3YjVsBcYLPhEhJlI9JL7
N95LFz8AidiiA56y2PRFEC3jybMRZ14U1UrN4FtNBV0yK3zUJa8WIEomrw2stQjE
t4kaG3BtKJdlIWW1Gk6zAqhk/vSvPRRJPyaqI+54rP07NOR1N4YcpPSrErzKSSwi
PYtbYgySv+O7jO5BJWAcgRpAty7k/JtHUVyA5+AbOMdDl29E5cTMHYzL1tvdalfO
H5NRgz6KYHQlBeJ92yX/m72Ii6VmRd0kn9yNkctcO/mVPE1QWIz1Attv+nL5wuYW
ueRzscRgrljt80Uq7PPg+WZfJBz36a0bQDZxUP5YYSxxVnu6Ovr1sCgsClflAPgv
vYTEbshKwmR64wFhlkb16VE1NWZmk4IjbX3mPbHOBUSogZI8QaHCnf4i4+EPKvTw
eZ5WUzlz9ALN4v2+Ae9JLcfMgr+0HkHccCPyug2nmbiWB1WniiaFSW2YndvAZTQc
R3vAQmvnEE92WfrhnjB4ns4cTwK7fdczexyzK+M+xEhV8V8LXDOXZS8fhlqJkzeS
YSMD/WftXbHTBMPdTzvPK9Q7IAU5g+WS+5biExu+/4WeGP797exST0X8rL+paQh0
Pf4W2s9Vf9Rnpg7K5sVH8BXS34o/J7pNRB546cVXhH/w7IYibiojjq+L8SzBMuUd
3YKPbMUCUvyf/hOh4cD/gej7ciDPi4datfcR60Y0jbEJ/e/12s3aofd6HW+ciQl7
KmOEiEhUS+4MAKXcr5iljof7LIkFyMey+Ihc3PO/nnAmwInnP31MeyFeq2WN/EuA
LCENNYwAjcTB1S46sfqugRXcaWOr7k/j3thvxZbmez+qnDMY3pn/yPEaa3jmQD2r
p7UuX1GsU+9PHwngDlR3Mt221u1PTNY8Ogt3Dibd/xY7EllN/+0Rwd2Xo43+6NmJ
egWRH9+s4INf+FLhwyBXgJlHhNT2WvL1vnx/OETJksnBVGW4O+Rsc0lln6GE/lPv
puDPTsP52KA6zVno2wQ5Wu4hDBCK1JSnh9LRSocyeknWkQArf/E71y4w/R5WG+Fp
VpW6vCck/44NIEBelqxpE3NWzQTn0UOFTClSSDRAQgNxKsww9DSr0W9vhhx1q+wn
+xRax5jcvvb6qTLuFZySKYh+0b+ekfpTk56HBCgQPu6F0MtpX7xZlPouy22poUCj
UZHXS3CX5Fd92rLLtpqaXbRfkzYYd3WYUcJfJ9HjQ5nSnk0FnzMrXoYXH/zHpdR+
W+gY5tTkUfwTwBQxCP1JTnIIIuhJW8JNe9N3tikeIfyT7zh5DpU6VVkFq+cgLdJE
CJWHSUoAeSbMzD00UPy2x7rIzWRErCL9I/QZSTKgRqGhuqXYOXxtWqX2jSg33g9A
wt4iyYWnfddotvKRD0Y+KtEmDJE22ql1Y6wTPV1dRVuxxomTCZMYvLdhW18NGX7o
ydsCjG749g7WU5WRrwlu4i1WKPrApURz3elhdwtZXwatocjzwR1mf3fxvrxVxNr6
uPopU2AUkpQmmA2gfocfxMacyCqM/lVjGDASkDERfDzskaYYfg0di1ADMrdsnQDn
9LAyYJ3MMhhOaQLhYglMt/faWFWb0RoMwBHIg3EcJL1PY/2iHGCDMHT+F+iWHvTs
C7SG/IH71FfK0D8aF5xTxYR4YdTjCnICQyDHX2sukoUXmt4xQR2zL7sT/XKc32XK
Y6ByUa09NIcmMN6lCug3SOQ5PJTZknwvBz05oA/coQMAjh41SzIVTQiwBeEpLDat
M9slz/oVuy6GqrgJ5ppfVzElGffodVP0fSK48RkFK6NL/fpmk7vDb2KaK4AQ+Cyq
9UJPBDkXO4VE+1hNr8WWbffZxSmxKDRYWn4Z67ZUGm9WGxNgH1ddnfoS4hwVvTT8
ezgZ+N5Z2XNQLs8TF3Ckd4hsSyoI8sR99mQgu8NZzWAQxZ4BNL9mYoj871/a4lAs
TImxsR1ds2M7/VdOxWJWqXmNnz/MaTr2Vt29y/cegZ0cQmguJ61Yl1WYvn7BuWOA
aNjrIPzmfHaqqlmsuUrcfbf1M8ywSPY4jgN3Sshz/HchoDtns+lt/CqtT/oPxU/5
qf+52lZr73Ye+iMebmHPR4XvWlnwsaG9uov0OqSL87cGnpb7AmZ3FhOVLSfWGBot
HWahkj7WiCYOe7iqxEt3Ze7Xg2ldHcPpFpVbStCg1aSEvQUGcwGb7Pd8LKn/kKSw
SVkob0JiYmNFJBtk7FaedavA9yccGIKzYTkXugt3sMjFqUYbNWLCozCc7ShybXrg
F3DtIUAce0CR0zF/F40qihblryPRO4RaiQQ8dsq3rHil7V9Vy0/9O1RxC8x8RryR
o6KMgkivnp7/WKPwzWDBbpAcU+k77pxTI8bPsFv4cvizMN+mTK7DdQmslgOxeG4m
hLbnVWRj3KdNaA+pyg0AANThTifHiovfOZY3wkaymgrWEGDCQfabx6cUAJKE9zFz
2oY/U2X+ABFDJ5Wgv1r7wSq+GMOUxb6hqMb19z6b7OtCGeE8HzG7kBpvY2ttvB+H
5FZtxBy0epM6o8eMSWBORdeFq12zUAvbkY6cKUvDmzh5M7axmprVeXhCWAzmCDA2
fzpU3CGDqTEEHfcBguTVUT8fke0PxvuUU15t7+NrdlvZsEvUBrCUuPWKcu9PWFAG
lBMjhWjMTdNm4Ev9E7PzmaZDgwUnpyeSAB2LvuxTJrGC4q/mTBs/2ARXk/ExS5PX
YWbhscZ+YIRheXjUNtUK1qN+we9OrnbcQBhJwbLa6sk/Kmrcj+GTbSao0gaO6l/p
vNZmnWWWTHjzgYQirL7iPRXnQhmicm1rHdVkWV/loKyorhLageDdAeIJ75qYG34U
j3QrtsbJAY+Qtj/hGkDoqSgTep9bFx2R5rxJptp5I75h+ETsZ0WR2vKhtKqN0IGl
YbCCV545LYjoNsl/0RNrHvRLQR3C1EzhygoHBc/ZnDeSgCE08E5ZZqfPC8R8QAiL
VnNHI6ew6WmBV9uq9ysNsvBqoS1GB/xuo9uRy8DMhWTJ51KlReXA/thd8KyJNfyg
FZAxuZoDE47XXeQbW45xSqMYdVc/FX4hcUF6MsT1atQBTde9yc7hRfJyTl6T5yoh
k8Jp3wpO+Bv4aVamTQmAF6e7AWdhIsMxTjqEZ6vxmmsCxO7/R5y8bLmvy444wuk4
sMK0h8ef44DAPGSscXHfvcOVjbpFF0ItgqRdOTYExzZD7b8TEUEv2OfEnBAOkQkg
sRKIIk97Ndd//McqlWXC30yX2QFeUlJ2MZvMvIvXcOwz7+eQ5fA7PHS5pOLz09Em
ykl+GjJFWX4XXONX6yG5zoEqkoJ27XEttfn4YI+hfCf9p0F3OMdSs/PxGbPH0BAo
UlsUwqUqipCNpJM6evDS05wXLwWanoZE0wegJCXPCfrcq/gjfPV+i8/W6nMc7TBa
b2I/2d5GotqdVE+jmsataEybZD/OzzDJqy9SxNMb+ut5rjsB77550Msu/GTRVlL+
E/MrMHD959baU613fgxCy74dE89+Ufp8SIAd0DTxJQr/4KroOtSLdhExRYVg1F5P
3z/L/rY2m8GxqiltixlL0nBWkuOnc6OTaqIi72reIF0GVaXKf7i6WG+LxtBLwtVI
eTvN6G+kEJPrIXLtMC1qh0UIYbr/aDVSFEEdLw7VWFklqZU0df1Ed1pZXFM43bBf
+ML926QxKuMVM6mAySTLPHXIGibOv6nDAkHPpgQg979xAmdbuIogzGcEEcFLQb5h
ivQVNU98ebaqzzRNVYqX571YylmA9mNCNd644TJ5G9/DXFwu3lumWmM5QeFOslAr
G+fGPgQnm8VSj6x1EfIaXw2XixOayvHnGiT6ge15Ncf6X31a0LDJkmO+QJ0Bi987
iy2NPp5WzPKI72Qe2r99EE1pKYLngDpm1al6PcApE+6mL7sW4RF12Vy5yaACCcYb
53OqP6EWTxr0O/43OgVlcz8wd83f0gAO0Xwmh8btLGrOtIJKEkE18eWASen7r7y7
8AWYJF8Xoq4wffyPdfzFh/8N5bEyBteGlswcnRNdv+4rdC1iAZPPbJIvYr5AhVDm
LqNZqpbqIx1XWnmQ9EyzlXMsEaUJjwWlb2y2DUT+bnvjm1+WG79sTmNviSR/cq7u
/yPV6BE8/b0DGWUMGNgB9pcdRZtW0bqo0S2lzFoqbQA6FDwbBOlSHYojtpkypaAr
PVrDbTdSJ7I3KYheRJb8e+wOsUwEEwzOYdt9XG/N2bs54u6MERibDKEXTT24aQ/D
jKwn3GhbNtnBLm6Gh865OA0Or1DsvqBIO9dxqzi33JAfk7c1U0Dhb7zzw6TAbvkd
CEocFhHeR6bbywiRfBsyUK/imvgAv9BFCYpcz02mLdegRXonK8L+zQNEgkbxw5FL
rnCiYcdOwYDtXGeCEqZ8xbW0ojo/C6qHwx4JEJHLq3ukdKdpz/7GWI8+M9wyhBuO
sTS9yk702FWA24xvIuk2z/dO9GAgXo93Nh/G15ihjGPaNzX2ZqjXtb4lnmDn7WGd
jXTtuq/ayWFQ6LRqhxV8p7LcXtKtzOCk/q/7BXT74AKKEPG7d7Ejt/aJE3FYpwfU
fYuYP2ufdd/XBoHk7GqPGfYuGiE/8mRB2LJH/6deyJrmxUGtWY85djOIJk/CSK6s
rEIZ+ljUUuXBvEAuFIDacmPCr+Mk64uFHmjmA8sXBukHVUmdUZFKYhkfsvU0Mzzq
Hl9vH9uSMbgSgt9ydIm6wpC3zYMkTHon2xCZek9153IPAnKE4WuDf4VwtYD6M/Bh
2itCIhJPb74DKOJ1HFhFBDd14KOjdolItQc/wdac/OGh1aq/h0ohNZY126fxiEnk
31FfKkqNYaa1X5A1i7jUtVY2YFmmzk1TV+CoXiB0oL/oAUZD0anl5VpUx/OaxaQN
qK3/a7V4x6QuVRqKxuhyozE/3mWZxUGw6InDC5jr3ulN30pU4lPVKE6zGkHVIblv
UddwqT3rMljLaXVr+Eu3WU5N92ef4yhSiVf8+eh9KmVoHYotxxYrSk3YwNgdstSX
wTL9kLwjW0+tgrgi8FIEl8vwRaKu+M0RE55hfwt7WIxMoqsjqCEeki6NS0dbCEOg
GKARJtPboBEAA8d9hwqRmaIr1jREpt0OfP1MlroVJOvfdi9dcPX8ORSdXcHCixJc
PKs5KQc69phLbL8HnLGCbqIr3oPDFMDRiUZZlpkslhOaWwfz9FIoN4F+ZRNGaBt6
dMCYBoVmAGzpV7f6oH+SHzvCTtrt3rezWsT9DrfpmEzq+hIDTUrkwKhvIYl//I3h
BancfujSOzl/lxadGzMIhN+7aFK+b2fzKaiL2BYlUSi5fOzmQePxLDuYAy789I8L
Qs/NuCwb4+BFFP8jNpb/6E6VUsg12WoIQ7vBPmbcIt7TIqDCTyQp/GnQMnex43ZV
zRBazAgEOhTnrAyC2CQ6KZb+J8/GxkqZArEZTpDD4g2VPbGQikR7u+jeBvxx7i/S
P0x3m+D3l5OVRbqrcF0oA94JtEAvjxEAVdrNB+KKQZFNrgpMvKFcvsslE7mtmcnf
RMJRnimOgaetflOGHi2iKTHrnWG9CofhigBXTavxsKS+g8+brvU48DgH8YVtGt3b
R38FbgGzO5QKypMggwnafq3JGbNAm4WQfNeurylF9ElcmOXMRIFzLER1Yw06innH
oZxBt9u3BJXhTd1vVg8Jm8RYsLJj8udTaskMMjcNDr/89IZS4vDsMgQdNYzJPYn1
QvIij4wpshGWdkL2C9NWFWN3YxT916kCfIkCKtU42oeIvkzJR8zJWFj7ymvCsj8E
Ay7jGnNH10XZCXD4Qlvw7yRgasKBeA4clM9WcXKmZo/gElKv+h2K/wHm2NKgt5LR
fOa2ipIUd74XFrRJeqEhZYFNu0Uhq/lVzf9xb6CtgSF6ggzACdc5doGt9ZROmo/6
/QEwU1LqpI4s1IE8v46e/y2XojsoeP7A38iVtKbWBWJ4OyxPIDwsu5hEXM6NMGS+
C0efbeqnGoLyZ7uGZzEIUanNBAnq5YOffXN+n5FO+AgONE7VDGKCnXXkxP23EBCk
qUg3x4l9vvKfX38RdzkSAvflZdYJ2stTZynwc333ZXAuv1xIufTpYeF4cVouzAxy
oX/BDM/T6YhmMHSW3YXJs1QtYPzGD0tUp1LLrK9du3bOTYweqfvNhUG94/nelzSu
uVne/wc+tolk2w9ThdF3Fmus2dCsG25a4n9vGFPj4A2tXdt4hmXhfAYeVO9uYuER
ucWoERYaC561AECSfdvAb8GkMCpSnaY+3aAr74vQWTr248W6RW8mWHSL4EqEl6i3
uUtnhHF+s14I3UqNRI/ulLKCIolzE7sXjBGbFaY+8oiosiQClHmC3R/WY6TvIOWd
0VJaSC1FJIZkij81oo0Pvr+r0pHsjb3Ux7JPX+QeFDUAIgLt9hEYNcJrzzsG1i2X
47/1zBOGfRGWblJCI8JCwvaa4Md8/FYywq6DsDsznv0BKWikpGjb8eKw2YWRBkyq
QJ22y3ytkLnv3eQNzd56F6xe7zYvTNcM38iP/c4rEH/M5pMVEigTwzLFHHGYG9xA
+WUac45NztY3B4R8ITGytesdz9C2DViXlQljY1OernGghDkH3G3CJuthUutX0DOQ
7/wWTdZczP6QdUib67qV5tUddxWaLbqiiSc723vh3XRP8GUPjeyl6wufCmFJStEr
CmNYQxel9Wk/U2I05WA1WHA2uRCaxxNla423r43x2qHR5PXAGQSBvqvQuaUmoqEZ
bXRaf63TkqgoO8rxtsqxo/uZaxk43Fbik1qUsAZ09nNzpWNtCj40Zcayqd5ycTnj
+YeZKaaRiuz+Xf8K/TlBERVXu/dgH+lEpfw9NGe2z8lxeLHIxLViAth/kT4XFsa9
bnC2Kb9UBJggGIZMmXbXik3MTbQAbQLXND4f31s3k1zw5WotYes65c/d5YnKJzbA
nMBM6Ud0ugiue0l42RiMuof7pt8sXfXoKSWjm7/wULBVlXfvQasn3eA26RtypbSR
IdRHwU3hNwNDw30KIx53I67rztyZn4iD2/ztpixXI6RgN21zOGBtONTT6jMwQfKs
ZkSPJLTBtyD04UNfvQd9thUB9izJlFg8fcs/gYR4/XB0nEQ3SUwLNHwSPTD8ZEeN
3M4Uq8cPROQCbK8fEmV2OLeT8tUWrIVTTMnV/Xymqz6gWTUMiTnzcHgmQmUsDv30
ou6/fvfuNKhVoNyTTN0jkNE+K+Gf69JwBTeN7dzCugsk0IeCQP9M0Xf6Yij4JwEa
KMWCYSOq8OmpQloqfoP6/tRmu6nAfckURthLEYSC5PJRxctkzmB0Cm2olIaOZxQE
qdpagyPWzwWULa+Nm7a89CEtb/dTXa5KpRgbTMuVjDQ5EPHAwvsgMgFlvZuFEpEL
I2k6hcMtEQK9Xew1JCYabzwwrDhaI8b2n1aEH83azI6xOtviNIInWSdcGmGzTEnx
d32xQsZ2h+nlR4p8u/gdHTgeNabxE4wSxQIANS/Fe6xsg+pmh7PDZcfWusWcA1zI
u6j4QMX9POcS7AWELP7Daj7/djPkrnW51LKfqsCHVLV4dQsHyMmN8CNAWPj9JuTU
5CQAAHD3aoAprXlnKBa6Qd57aFNZ3ADbQthd25hCXVVwXg8i4UG9zsL1EmoLNPS/
vdNEoUu/JRqPToF+yKGZ6tI+dhREF3KtOULNDmnRva3TIeENuC6CDt6p38+IxHkV
ttbivtRNWIwbdhUcPiHO7rknuEg0dj6BvaE/UrpvtD6cbygl+tRromOrj90c0bi1
bEj6eeqmk+R62LCyuBIPTcgGkdzu0YQDFGOkQMywViuZEcKG3C8sMfDuH/DAuhx9
aD9KynHfeombaIhbpkjkb97hMj08bTokz2d2knpDYTm+Psik2dtNU+H0v9GbA1O9
MfmVQy0DgjDv7gLSA86QyNEkJdNV1nM6B6OEtmIBZOKkXe8VnhIaXtkQCGzfzP30
pfHoT+wxCSCSwldgqFDjh0J/IFFA1ncwN6da3i7vtZkiGMVshVoMK6A0fHS6KKaT
oG+HjwNeHccBoO/vEHnbG/h7vt7t3HLQ6U6PVSUN5fClSW4Ds9O01pqDBqStk6d5
ym612syiCUbrnMxT9wXsS1JuR/vTb8OzbZd0BDRQfHBZcDKAkSbUuAfXPSodsWaW
iUhQm2hJC0uXPxOsw0Pr2BW9h0SB7FQtNMkkPNcR69qvpybjK+yKJU7Uoo+ExFoj
5Cv12eRJMxTuD72VvnETjR5EzZp4daFSeCREP3dqxkp8DEfNC0/qnngNvmuW7tAp
diFUGwUx8/+xqpZrjgLj0iO29sNHgFC1Lx35Ymdc423KuN/hqwNjufwHpQcb3IXj
MHMyf3cj9AvC9sS0aRnmWzKvICTU0wgpke8UeHHjnSoeEjcGUVOnQAJc+OBXBXnQ
rZeu/Q3nAXmpxihu9sYzwp+y2djLe8gJ5N4pNjpDsoizdzfAbXDGTDUMgzWA7gfF
XMhYgrdtCkZkQUKFciyajU7CVP6W8DpBAwLCt1ZutFss+WZtIIeC16TVH8CMirlI
GQ8RxbZbw/tj+N5FoN2yJ5GLJc0b7kpAFsNH4ryQd1ERcPC9jxMllp/uQr5YgHpu
+5yjektv3ZffENG+KKREnTxD2aKoO5ulAbPlXlwXuPlpM0XL48Vulsevj1cU8RGK
UorR18hRveNsIEsH0dkuUnyonkdlld8xGDNjMBayHoRwkQUxZqb52QmvcTGjq5wm
ImWZPM/c1lCLb2OpVttpWiSXMGzMv+YkCVs1s8wZ8OQzLvJPBG9IxmJyCpMVYOtA
365u1YK5WlnvF7V+3YfUZNKF1kmgDNRmFfnadnk1HJEk91oFdDFOnmsrbVOsQLBk
Szj3zO7tsQkpr+t0AZa1nNE7NQuYAoSLUwAVuCkTlkrEVlxfGcV0wGJuc1v+fM1p
vFDQcL/wU2fpZlhAnh0U1swpQyWc5e3ZMO2Gig6braWgjK8Slrji2yeNnp0/L0JQ
sCPgYpJVvGsMjCHi5DPwSEvayYXjx/ebPTtSpdaomhdfxz2jN9PyA0xuKGbrH3ka
Kx/4FGuCatlXCuLdnODu4wUGUFy30rCOEYFXd8X0c3yJ5n++pe//57Ysh1PO92hM
YaGFyYhw6IEFpmNJDF8A8jPXtware5nbVhXgOwQLjbKLKi+Y0GSmIIXLii5dHBEh
pZt4pyX6Qfv6RWDHG4awYUMajzK+eA9TxKEBRACXq02PuW/tw/GHvY0etpLhdM0U
iSUfat6vyDtddNTM22+gdFwfCexlDyh/kDAAGtTRVYDMf90Wv0eYdbv9rOBGehZt
5+M4WGpvWx4lX610sG7F+xmGzTla8eElksBhqf+i1+h33vN6hvqYNQxaxI8TFJst
64gAgI/wOI9Cq9euOgg1eSP6tqF9fsXL8NVyfAkjP2mL7NyY+Rx1Q7JXjqZqBuRt
tegPfyB/U3QVAfLSf8y5JXxzf5OE4ttmuJD1XIo8xPYhc5915rYRgOID7QOey1l1
E+Flr0e25PTdJG9wsAhTR8KyRl3VxCJ8Z+XjDuqvV/3UXeGgcsM2+mAWODNRGp1+
vw7A3L/dcYOuXYpFfSbFSH+l7cwI46sA6JiyIxpvqW/51tTZcAiMx0FXSGx+49OH
O7KTzsoxqZ+2UUCYdAm8ReMaYko8IcWbSG4d3W8CkCJ9FY/dSi0hm9tlXfwcZD/M
fOsbNDBDehW3BELrHhixE/DyEY3GvDBmaUvGymbWouCyBjuYgnN/kPeUkPJRwjjP
z2n7erGa2cr2qDuq+M5Urn91/L28ZH+DatBMPuhXwQ308GWzT+0vJ++JqJ4PUEWm
x9FfiZVNQuBzCmtuJqvAIn2x+5XDxnomRHgbb4F4oKGwQbj/f6+ijUuiit1LTQF4
GPv8muuWe1qk0JJOLPZWNxfRWzHFG9mx7A0v4IM4Qu0stoxtHF5rn3O1XGjZOtlr
XqS0y1rPRXCGKdeuehvAgv9izVvYLITI1eMvt0ThPVHKd7BXJGBoPYYAi+peXihK
ej7jtx1Am7HiyMx98odN/qwaIA5mrHsoQNnhlLVEvMe3kpat5gSXDHyLVEFp3p1s
2DoOmGBLagvi+uyZmF4LDfNI+1IlcoDuvv28K7dCC2DpTl6a3BYFl2E2nxBlnfju
zhOAtgBivUIpFr2y1JIGcWJxTclBcJHHmKPVMo7OaltfOm5cSONtrSrwz8PjDWRq
Hqrp77sAdDfbWElsP1VbTJ1WI8f/p0DMfhDiPr5aLZmVzj0FisZslxTHWSfdmdki
KvqDp2YMUuJHWUahdc6fWFzWHncSO1+xJlrLgm1coURfgYLq2hzZO8vipLjvkNLb
CFBtbaBXQOMzL2VGn+4EaW5ocU8dq1Y2fwZ6B3/IcURfO0AfqI9+9xOieVSM/++r
9wdBzxiGKnQsVByX1xCYgXBiAIlEadLfjOAL3kObZ1txCpKIR77yMCqbSeMYmkeM
emxhkDJXWthDJioQh8k5mTpo+d9omNevq+HnajfOi+njdxWVFz7GJISPa1AvtDKg
pQDrWxO+z/6Tknet1MENxJQPlHIdsvIP+ILoqE7/hQ6BXMsz632WxTKwFlEK4z4W
5Y/EY++hTtEkrzzvGTQzaGGEzeuBrj9D1LqvvGgKenRbVuj5zmPupIWqQxlEVG80
kJKwCef2HiS0cfi537YQ2TCek4nnjEujsh5LOWEMTszxOmPGBjzl5AB2BpNTsmXg
mfzKqLDrvKxHUGoT5HI2FxRnCPPZfMMNgGK0nV5lG4939JDNhw6U8fRiBlsXzHS6
JHd1wBlWd+fW/0VIzTrWE/tDBN+PSTMdEI6Q2en40IJI6BAibOqweh467U7pnBia
Nd0aFZT58G0yvoigZATDLRj/pe0BQ8I/EkK2XztXq5MK0eiJbVvglfjDL37VOfZe
eLNDpqqr85vtTW55dpAs88m3GL/FFkzgr7ZIMTgxMttmPieeUwejDPvd11rl7nwb
0jnYVV4Luc/uWsvrIh6Q6c4LvGhVMZAn6+TzgNRZFObVOeokJiiQuhGMnZNydEXQ
x96CXPxQt5hGtrRAWnjlQSk9nyeuGpMBycFJ3+jWLUXzYptosb6dtYfFPK19WtoS
2VO9/Hka9a/V2Ls+mNoWwp1I74DOrclvgLg4tHaT9jjwSzLDc1TNBO4jYpU84GJ4
GXtyM/UarYZocS+/KRZOPmwA28qRawCSuPULh1Gd/yKwKml+/K8VIeCo54hz/2Ip
IPe6dWr+0HYEcBtM6u3khogIo8mIpuxJ0jQJBg9Cd1NGhvzMScBK/wECcK9FWb8v
4nn47mVZSNde4BjaKcQygFmkNXRXj4RmkDyJLxqJtd88fIEEC0esMqWD7vrWtU8w
b0EyP+maWuBsu+n/zHbunL69qFpbR8rAeb68YwlC4VSLv6soHAOjELCXQwvLWybl
rRtYhwPbbPEBydT0ECEwje+yA5UwnUGbby7vtwVd2iZDAxBA/SAat0RyouLX8WN6
YApSNsQ483jFCWbsXdIJO72LYeSebN2qOJ+3mGMAp7CdMM+0NK7CxcsbwlpVs8X9
+1lyYOnlpHubyX7HxqqdQ7RcCjdsCkFHA5LsYhYimGrNnNGBgAB9L+/CGKfiUvWW
RA8H6C/8jHxzjvvyHRuIjt2P8W6fYKlG0ANpQCnXBLp2xxHVZwlQPn+SaVjPB0po
TBCyZ9Z4DH9fhqyLyJxFeLvTUOlsoLQe4vNoAXvVheogMOB+Wm+YMhb8aBcafQla
9lHpK9vVRbFsIPHnnXMM3+fLZ/ijHThv0OSawot8LAYjJA2BjnlEmhLIzvl9DpuR
oJF4L3nJL2j9wal1FCK10gH2GE7+E6z92DhhbjY3lwGHUdMCBczpZKRC3rH0poDN
bA1ZRnR1nGffAjYOBVLs0SLhdTykgknpCLxB6qm6YboSF5UI8RErID3fa3mZkr01
qLZNex2n/B48yRWI5cT3gH52DbLeoRyzWCGGGYtVgsgD+757S3RLsUArkRMf5b6Q
yTDBeq1hDxzMcYQ4P6AA5sbH9Q1jkNwKVgCdcxtfid7ZANoMkaGlNSS1dXRgWgcm
Ck5/cTz7Zlil1o2wu2NnOwDlhZ6hV9FQv+VLnjbUZDgzzIf/rVbrxvTT1qgQnG1d
4M3bpEQh1F93gLdbbbP6tgQcQo9WPNabtvEuchvsV7txwXW0yRVy8drPBYOUzpdt
D6huxMRUQkxHNJikTLavuia2vcV7a6NH+ii0mU9bVN/eFn64H1mE4m+67QV/9ORg
UukQ8paETEOsRbwIUNi/FNnfTUSAcuOunPYnlHiKKY8puviagNzA0ygbsGzl/I5m
mniXgHal9INJ0xaHxu1ne+XIYDUgD05YR15pdJ+Ww5aHjqktGIyWTmnILbBvo6cK
e9zXwHfMJb9FMTuC1BCoA9hSlZujhhJDF6GKp1stsLE6cNVzzlf8jSCl2y1U+Jbk
msn/dCJCz8K7BnXviK/4fsSMBljw4QaKpfbFgt4cxyFE05BtpaCF8bGYszxVNVuO
/FXrt5cCGl7OSDApN4FRa/qun3Om2CQhql7vpPZcUIRgRbRI1ZcNgGusuRQ3aXtc
tqGszr+XHusEReuVQGmc1y1CYgrVVWo+vPqU6byuqOQpGp6d/M2dcro50xEyzFUz
jHkTbN6nKn/rgpnQGlLKKI9SyS1y5f8qpiavraoIa6Phtg8yh35QMAnZ9ldlF/EP
gJq7qzcmmRc9vUM8S5xyWV6Rj5ZS4UXw1IiIulhvdbdayxfffBANfXUUYowYCJRi
t0vAo+guzuMy7fNIWTkYKxaMSw6c5jvgH0rRgilwTGCXAot/LR45LS04V7BCjtjY
hvv7yJDgICmP9aTiI53wEScq1WNPpa9delX7z+VYWAdSKpXYvIcbneTmAeVRml60
u2r5TbgUH0kdVRWeiOLFPTzx0HB2E9dk6elJyNeIArHxGvaGLyPkGw7rQlp6374s
rnrcpjFfBXrpYweDY3KlTGvdwjETjd1iMSb5CwhCS6fb5MEPtZKUj2I4La32QXs0
W5eJPjMkVoZcSvvOCdVknMX8WTSOdpTnhj2FCtWkV/Ta31vpcH4zfxlMnRJOApGD
bgroy+wvTsBtYAIv6mnyw3quoNbhPF+X8eXdlL6LZtZ8JvyqJG1zhz5LCDZAeyr0
JmxIWNCf7LGC0MzH8SGT+PrMZLBiyUnZ8asVLLxll+3dbGg8zM4sRiZy6qRCDZd/
E42yQ0P6mk6Au6IneoDfFb3EUNkZZcloIShDz65iiBg1r7YfrUjL8k0L7Z/xO3zW
VTFTC1ldL5XxpDJuwL8W1iiZOTjr5hwzbwLI7RCSw5Cfr3qcyfpLTF/Rdj618rUR
xKtCbZWH2mX8lWbLcYJ9ww0QXKaLlZMtSrPkqhmhKbMnXL6uDdBfBSa4AMDe6hdL
vrwYx74lM2yOJALcTO+LGrNy6fGIS39GBLZzsbRh1ibbno5k85uHvF1MC1J2TYy9
vstVOiHx5IVfvW08pTiP5Hxn4tauwiUWM2OxfN//U8LNfrxbWs+lbxcOkiO3Wjms
7Z6zNI9jpMIjnDsLH2QHpbx6TqKBZT/WsmGUa0oivnQvI5JZ/0d8ekkiFIGeEZXD
m6/wQytVf2ISg7HJhfGPhSZivbsn7hO8Ik76iGcByY7BJzFI7ef+F4FxXssI03bw
DAZ3HrrbgjAjefm3RM6c/RsXKeEqAVN+7q1KkATgcah7cuRBnQmonklfDI/j+kdG
PYlDkiugkhqEyHJjvXJppTEqS1dE5Mk3t1487lu4I1OTWHi7u66l0feCNxcDuYLE
vXlC4P7HSduI/gQ1MDUR1Yvg+nMaIEz+88OnDwuO0GoTF6OuTBA6QE9Qvljm5LQp
ESWU2ogj1Whtb3VSFHUW4ExRmCHXLhNej3slol5V8dsF37DgKWbIZ/gyvlH+ZuFE
k7fDrYlA3HWYG+bXDi571kYAaJso2QkwV+q598tDTF9bLDC6JCEn1keRjwI6xkoF
JQS4/RcVL+8PGU50GxKUqvFcmDKzsxUsR10+6e58DXgZu+i1NH6s05wzuhUHjINg
g+95lEDK8SpzaxEQr6lFVQjT8HEylCMC3a20qLyAhW/xNEXhTMy+QLOlNtDNXXa4
s+ydoPpLtk44mtiFoc5YuA/GSAinJ3/tD/Zj5XPNeAGfm7w9Z9sJBh6GEleHNS4q
/ib2QuIO6bwQpbH5j9ya9lCvGzk0XJBrrZ8Z9sWWeCldnJ8uNoDqlrKOIoJXpK0S
5Isjdv6wxM629xYsbJFHTCKbkHoWJan6QuojY9yaVKzjp4ONO7GZmb0BCQOWeIZZ
21WzC1tKDWGLN9dGQQLXSrqwm3fxQo4K1W2lwAoiEQvydNvVKQEBOGPgMpMcjK0G
h2zCElRJmIeXgulhJB0OOpOjb3X+5Jt3Lh/2G6AKouEQRMCZOaA3b0V5rzStHoU/
kAD1Q6He38uyaVcEqvXCKQP3VSo0sqyFPPcrK98f34ZnPA000wYyAU1zkVOXAp+x
Q1OChT31bU059WmnVtPhOgtzf+vK9gLO7ZfdAR3uWFCUMh+PZ7Kr+rQiB6ggAOYy
Sw+Vsffy4J3eDiTyvNlbY1QCiNj+GAqusThybzmethYe7WWtwiLEEhtn8/YIMYVi
2fM/JyY4tcGWnzPW6ByiVCPzZniZSoVXIRi2LiBhZ5uJo4qFpDC+bbjRnOIn3AHu
mY/qk+lqVb8G/6wIe95hYD8d0cZKOixRaMGVUfvpsuGJxpcyyfqN5XicnSny34C0
tFWDBdmihL6L1PB6zL0Z5IR4Y/6nowNdzJ+lo/oO0q8hYR9QQaKC4spoH0qghCUj
8LcKXkviPH84HsOSGufbh43JkQoxkJhh+BlrBiHl2rsHcGSxDUCUnbm9nv+XZQNU
lOFM6EhO7HffAPBm19Frt4nEiJRnuBJMuGI+kUVvHlJUUsHqf/P6pVQfkz3WXHNM
KyIsA0lotmJXKbfhuQrC/Qf4BRyj3+CDJwWdUEMt0L5Jyfi7utvHnxZIV696rTbh
kVNml42s7k7m6N4/9m9FsEDx3EUkum0PKlQV7VMdXIA3Yhyo3gGwiJZjdrHIKTIR
RmzXd3r8MWn3iRCa2NZywlJO/raNTy+Hp2jiuHEiQj1J/lUbJwIH+woN7IBSy1VF
EfEo2Y9h5LKPA7CxsDoJnR59JlR1F9wH5wniow3LVmaMiI0o1AZTfj+n23GJ1csG
piO/TjX3im5i8+wOMKFjbwiMHHsJ7NrXBHYjltO4T78gHqAQuf2UEq+GPYGpuHhA
06Igz/Gn1xSxPv1oZ29ANQG+m/YeP35iulR/ssVlBEqpoue5jE2IJj6am6sdAW8e
o2wp2C6PBQK1cyE/DF1e0lhAOCVfummsS1DP0D7KRCd5QgGHucIaHAiH8QbpN9Vh
lqF3nxpVrp0+KJRD/yWOF7hhesPfIyaLJ9vCmgDfQKtR4IfFDqZkF0w3X1bhZmr5
cGoD1AOFmHtSpNyFGWEBWNSMXBPgzfu81VlUK3rR5ZrNyhffktpJ8MRzv68w04A9
31y6B3VAzwB/xwIiL/hazoSh5CoqgVjdnDWzu4DwgFBkRsRn3RikX9+/ZLKvgsz8
un1fNcFCB7+sVrZGykKXFLOJ23JWuzOVXdZTlZi1yrFhtdj9BbYhIJyVWrCm+jUm
i13U4R8ya/2tih2EM93ljhnZR2W8hkmlmORL+AD48wHLjsFnGVBpZ0Ml4Virvq3U
g78prgatZEW2axQ8rV5T02H+lqNkrgY6e6hsVX1KrSfizC1I0I39TzXyxaFjpqwV
1x/oqciEK84re6KRhgrLUoOYWf+6AZA+VkWhJnWMRdv3yLMKYBJ94xxSWRhKCXWg
/myeThqlSn2xXDjbu708xYv/Lak5bhHGguSIq6B1GSVmy8PHzl6MgK4ErcCNzW9t
bF1NuKdk3blHhNXr5ipN46xK87IgDqR5UXaZ2W8SA9cUurKMmhjsPETcRwEWORJy
QyBL26P+0nbMqOge6i1uswyKI/5LCwxONDyPZ1xp2LIxDzfmZZM66lh0y9TV3kdG
u5aPB4ZUNxvKqmqRqj6MQDWcGoygpG34fLfaC+OEuLTWjyy15ogPIj6KJMnBKH2l
wQ93TsLXVx4TjVJYbQvx2WQ+OO/1NahI5+HajnhJBxnyJ31DTDK5JULedTzcPf0m
d87EeCuCBM6H943CEoLweIMli9OZFkmOqrpxKtQ2hUT6z6dTXrMPfOiwGaq5nZF5
3DrapdZJbOD33/0QQRHVVLoFAMbc9fPn9KedxU6u1oA68gTqkzMO7fbmNehfAcsy
Y80bnQ7OkYbdtuKVPFLWV+F8x09sGeGelNfczUGHnY/iurlwz1fFk6S4WRfANXg8
gvPCzNBJmYaJ/FutW93onfZnHZv7EzBEbtY2XCe/gLi4aDkCeq2JW6dD8UPl22wY
4cLMsgIyIGKh8o8Ediz5uyS2uxYQ/pJpzV7bp3VNp3MVcKsDp9+kYNYg+WjHQ5MJ
DSmcRoEhwmI/bK9F8QCu4wXuB6mX5i1KWUJHVD+2UYr19fk6YtJQk5swHS97wate
5toZvFMEXJdsA6ZYejLc+mB8PR7K4UUJ5jMbtuDFxAaqXLZwlix4qi1QnMRBhOus
WWxzmTFgyG1A2/BUoRrC+7BeEUYgLK2rX0mW1neek1MEpl1XIZKYDuBcmxJRUCr1
kAADDd76MKGRI18RzrrfL6eyp/rZf0GBMLxN0PIzFkzQcZ9ttN7snHB0fYfyLDfs
GAw5IknJVyJFwMtIAhRcL0Y1NeTfNH3hNaF6bLp/9LMzT8d+BmWjKtOofrIOyLVD
Ml2SRQw5EjFWQFjzS40Yx5ki8Q0P72qnNYAsIm/Uoor++LIjnrI6M1c2q3ksQ8sE
vOvlvyVsZludl7cpmIKU10wD4zQMJz+FNtPVKY7S35wJVMV+9eZ22C3oLCaONrU+
W+2cGfQEeYWwn/xbKDsdVSwYDQTOXPlZSnJWgIOn9RUkwyeBoh5yx3b4JbzLgiO0
q5KANwu8824xm5dSRfRZkCPZxmItr50Mb8yxncdy8qKe5ZKVY+UZXgyaWAuWv2Zw
9ytioS7xJPfeRQuEG4NmUTBOCxEBX1wLs/yB1OH2jOrb2ZeqzX5EVgbKP/eUF+Xq
my8d+fE2gSIN8uaKJsSHhmd6GXGs9nL0Is5aobpFeFOyFu7bO93vyo4DN+hW5lle
CpJbhMUBf8ol9KnTQzbjepqIx32XyyX1gsYQibKRgtNZnheS1BQHaTEAr48H0ykT
kPpSVI7Ki4ZlA4zHWbV7pjukt+tyb3ZW+28iA/4H1aO5/z8PGYXFSp5wSCwNxmP8
UhhQt/R/bYJo98WChyteMcJDkQi4mlcn3VN2Rpnr2Rf+wV6cisfpLwHfSKh3jmve
ndFjcMnnUXUQ5GQc/C475E8+SG5eowsMl1gk11NyNz9eMb5JUVdMo4oEF5VPmZCR
xP4182nqw3T+0tJzUwQbyWUqwnNK0sPrqIzv8oGsO9UZiyy6xPN8Aigi27yzCREF
/XMhFFer3C+LuLD0H8N9yFPBp2qSA92Cd/TeFQ9P3XnN4cf5WYODx9cQI3hiuAhf
yNWavxRsp42AJi6g9VbaQwYcpBLuLeIfMKCcHdZJJm+LLb3eHiDwIbrboWCgnYmn
E+Q0+9kZJycFdzpgv4HzlvlFOk8yI+OfvyN6Jic5UfEhXVmyK5cxEQkjy7W+HFF0
axMB0hpnkazG6IOf3CiLZPmqYjYmySe9sgg5CCDB+bZQJ9cVz3aQX1BOuzFqWbL1
3Pnu0jXB9KyZ6rCtWwOcqTcVuhMxqCdYQb4HP5jH48vVUvkM7liZdcydk6llMAZL
hoFZ7Te69Tqzkeiri4jAO9sRZcXCQCbrhq5gh7r013HlKlDxjlSf2xpiOmbbRXTb
tsJBJbUKwvj1rYgVz0Y7/YLoELqsNqKIqYY+rau6vpIOyVHxYwGvgM3XypNGoMZk
COUAlboeLK6U5lNA9rCbS9OP/D7EobZh0elHYOBZWK2xYNpLUdEl8YvuxAGkFGuN
yGuEQYPG9xXzZQyXG+dfmF29/kSMopqRy8SgWFtRrF8G8mJf1QH2iY6jLSzYa4oT
F4LR2+mqOyT6jv3X3R+53tZ8S5q98R3BQeNL7ueHB38m2P1ynmJB0QfxtrBqSDa+
IGo831xbXlYXZ9oQh/qeirO0ZGQIiWilgR+FHxl9eeN7/3FQ21XCcwESxXQYLOWM
tmQRD6dRi93oBVPj2PhZeYd8ye6xJjxLRVkRCYbwweywHOrgwnpOwX67B2D2iyRO
erNo/nTC07JTVXnz89gmVLNvo3RtcXHB7wIhMTLZKMAG3xn0H6jPWWNLjEOH0+RH
v2dmt3z11jfzFQlWKqdSWNmNvHdgOo7gkH5AyPnV5lTTa6Bim2KnKsLKc6dyiLDB
Cybe2Cyj902bI+Dp0vSIIL7KcnwXPCEGLQWgtZGtdq4VKaH8augQ9fMN/GlI0qJl
D2TE4Qfg19SmUu0CGquJLD7sSW9dn1gwk6b3gTI6Vnr6LSmiTLBc2KAjcaK2+lTn
dcHqDbiYylDUiKfTJv1zM7eftUEjqBrNI9eu/X+vLC/bBkYU64SuL8QYE/MPQhTT
wP/W5Wb78uv3j9AnfvF3dl75k8lD2WnkDOL/W89w6MYzEIr0D9lAW5vKTW9UtPIn
70Jl/UuQYqho1m2kVD9lsQyoBU0p4NwKrDyldz6z8O2RpOiWQou4IGC9Oev8Dys3
U0/Ic0AcYfmgV6m/1V4G4IR0S0FSOASlPEdAAkigPuZoF6isaSSz6koW8UMHDURt
YzRib/vWJsvNiU2zjB0bJgwRZWkSqrSRh5/IBIxSns5eOpqGugsgp0ZcRNLRdJH/
fYuhTrAju/h5u133W9bKBzsuqTTZe0mAtJFICDKJHWmSh9pIoZO4j6OOUf4K8sze
zL1gA5EhpodQ9Vgvr3bFkYMEwUH9w9VHhqDjcrU/PGohTw5ZO9+kFUpfHFuARoOb
VT74L56Skhf9VP3dUUi7/asrU36vSJAgDAsEckPll77ZF1Obw7MnQQlvewVrFECi
I7lN0zwqHtH7wI448i8c7BjV0c2hlLYZnOds23JZo4p+V6P1pIPAFYZzJck7n0gQ
M1HHbh0iv4J4tVwtJ8eo9LNFimsiO0h/N62fC3JxQeOdw9w7VGS2/szWpws9/okU
slma0ObGb0xnbaiISVF+fgBel4mojRJaS0sgh4pjhCl7dBSkF/OivKJ+KRL6whR8
mUVnyeavwWLzd8trgxzCYHiHvloWIBZtuAKrsyhHRWHYIyGtG0UqhYFZ898m/ApB
11MIedbamL8+99NWQlKwmUTvgqoUpNcgDg6nT2Pa6Fay5viggrmnJBZ4jPYy2/2N
Pqdx5Rc8dleqwlnYiNAmK43dHHF9GNKsxsF3BeC++VccTLZpLs96MVfBLSYf6bK4
Fc2C66slgH3lQll6Zsb0WiepYd8FxujJ3QRN6K7Z0SGOvPv8/sWVx5Vx3ZDiJgLk
gUIEN4xqG9ccRA+55TAdgW7sV+mO9nuVoNlQo530W79MpYv1g3mosp5aRDaaJFnu
dPS9PXoEo2p5TLHBzZs9M9sWSD0JdtaVQvGDJheB/BeGyMYh5vsH0KW9uX7p15+E
/1JFzaa5iIsAWpUkzMIHHdy6oCmSug+u11svYlP3aOXsHYxcZDsuvke802axOsET
rMPGqsMsM79pINa3K+k0TsmqGxbWa4/FPxadirTK3dRiVaFJDkcodDnedCKNIqQB
Pa9mYjkXHL2X16vXBTkmvU9L1vpKix7IKXeUMRL+Egh6uH1Tbzq9mHv3P1lgBLhP
j1TKmVYtkm2FSXn6vkj3Nhciw1c1ieSjFLcGIZUt/UEI/ZrlmEPFqLqXuUKnKw3F
/PCMnBXph86l14FC06EixUXXTQ7OfbMsRRgAeHOZoJm/HbX2ElUpx0SFemxUtjgf
PPn8InAa8U+Ou6p8Xks125X6JOM6mcgfuHrY8jT/YZWUhLUmHFcctF8XTLZBArvj
f7pyI56C3SVYsYnIqbgD+8tAs9R83z7+Q9bKXcwjuoIhg8bGLlo1oneljnjm8drl
qKZ35nEgQYJwzChorKG2tKYn+S8CCOlmIRuBmYJeCc/g71fCMNFLziOQ3TXaqtvs
FBWMjSf7N3RI6418IEU2UAz2Xbwnve3EIxq5JOaz72pqBZdaW2g3HMGEJ2sARf+t
HEmLsr7scuM1DPXGcqG64WdTW75LsltG2nFsK9TOhmH/CQ6yhjQgp98sfSH1QihN
w3zJ1LO7xTpBc6KXc3g0JHZu+z7gtCr0eo6zB8ZT/xlMdbR+LouhSUI9pEqBkgvg
W32j6gs2N6hPWi9HEythcXstc+YjU40E117ZDA+8S4Why0R7qmAJKSupJ8dwa43N
vvWeRHOGFYe5O9lhn395bfKCklWv/n0XZe/RwM5ASEUnFs0XjieK9InJJ7XOugNQ
DniPLaGi8802QYMwvlSPh94czMKVg4S9//6mRlZ6zqm31SfG8G3mn2sRbMdTzv+L
UJ/kU7dXfxxBhsUJOvHEsgm2a7/dBhMV2fsCWm82ijTUY5iMseWU+4RMTIvz1mS2
ujlAijjii9z7z0gR6OweR+RNCxr5y2kVMyoNfvPsZpLtuZesIRLqOc4GbUjG3g9S
u6nzk4SjEAJUULF6FOGmmBr45BEmyiG4mxfIVCobbctbksdSDMbj3G1PRg4Ogoib
/jOnlQq3GDIQfmtKGubu0OMR0x/5Wx9Uswn9n++hDLQLjGj7lr124xXvhDdLmL20
v/Rf/PoDP5svMah9G0QWCxqOMTlHHPIOX2luxYfIBAa7bB3znPluf+Hnnh9PFWRt
I32fTRluEClow7GTbqL/y7aDEU6w1HlpQg/QpvZpgnVGOyChT8MCE9lOYmeESB5+
3RlyI0ZoMl9Ae5LNsyDNmP7IJYzfijXI2TLXNjTakDYxAPbT7oxED+++73TgE7vM
ASqPx6ejcvAxh399zEFdJqC7Zf7zScige1eAEJosJOQT4LsELQBNZ0XJ9a1ijebP
ejmO4PRaPwEfl07zpzqR2il7V9jthLN2rFkgIsNn+YgCcv3flsA1BIITR/4/pjxl
IMXghkpVok024q1Bvji+fAeJ0K+gG4BeydhtRAADnRHtwrww+4WqNtttZM8oHywX
bTkpL633qCjNlmXpwjUaqNbcG0/U4uOrbMc6PB/z/K+/8JVcH86xRdipQiAl2yhg
isWooK+1Ushfx60wGo3TOUMzrIKBgc1alO4e5mM7FolMqFp+33GF/4yTB/gZ2udN
fEaZ1FLG/uIqmzfG38QhYrdOCmnu1oGxuuV5VX91NixJFs8/nVs3YisUfl4X2/cF
VkrlzynS75FLqECiDv/gY3cFrBy7qXcNeLwhYug3BZlnwx/cATVxeWNR9A2DJ4yo
hkkN5pA074fGsEmv68n/1nyh/rq7Nx1Rcvc6cTsE0p0HFf3CCU59593DCh/6i+vD
XcAp/zosdnFXqCxC0tsXuQtdHvVkJ6Th1EqCFD/9ZdGtI3ysnLRI5u0hr1jceo9z
WczepIdNhYzFnhaT2O0gKYdeF5BY5lXmsH8ZQUs8BbmJUZnFOCaYn66p2stcEb8o
pnmNvmHrnDr/3AgWboe69bq48MT72AVMy0B1Hf0M1WePhq/fVbryTqrOtS9N4UBn
JLGnahmAq+2t+/w5fsgzZP3VJ/2DkiGfghJGSjHgPkXa5SUAsU03rdyXEGG/eW5k
29kVCA7cKdbq9TvUKapaqk97f1/Ir9v89Xl8U1pU3IGHs7uOWC4sJStAk3a8AApl
T50DWyXQKjbYeOFm4RjswBZjK94TA5N0hY9as3UjmY2eT/GYu3dnFPo4WOg5ntMV
fkfyueY9N3k/Na/QEaOUSvrTlBrWavvVRRWmN3A4GtsZGCQUZg7nwWG08f7O0nsX
8K9YHN7fclj7rA1w5unvWtXpm7m6mOvwFgwtPRqzaTEW4fA2g/5thF0y1ZiueRRN
TR8Ams/HMWKVgcpBQJJeLT5z7h4E73og3mboTfQP2cmyzbCPtz1G8jZrdgKoB2jq
Ii1+jH4FNF8sb2bc/xsqspO1VBCjm+uCZeRbEJyUrTK4R0foNxbD8uDE67MXhBew
ZGKJJNitRUHuPLpTISNnHiuGliuSrFM3h6RmVeozAteeNQRSlB2aibpkO9ExwXm2
Q1JmFiTTUptavfoLoZ/9zxDeNefFEAz/af9deZ6DswhXkcaQEY2qnf6RlQLzpQqu
9lM6lcxvhS4hIuiakhYmKnjqFA3xXtRJEr9Ca4PTY/oBrA/bfqarFU/QvI8sdVzd
3ViEgy6C/YIEH4OtBcp2fREEG6S7Nyf28/Wveb65E9q1OdWEE1VbTljXc8aTqQgx
zq243cFwLTEqVhzWpi9IgllurzRayEd1jSAIT+mTz+p2pZSgp3mhEmpVvKJZeCa/
Otk8NqvIHtfKr1eACBHBv8hfxM4ZB7tjkHZZTP3Q20wadqQpSKqsvUn8EIPpXBSh
sbF29kUAqHVgvBi0yIx+HGGQ9hEQmflI1sN80T4kTDY2xOw7a7JbwOl8nf58W84z
Y/wzBVdeyB67pcqIkIz0PaZCiIEX9/ni/Sc9qjjpwQ6hu2sq7KDsdHays6yKFOI8
uFvGEZvnx43mQ4pdBaKIUvcscGHFySGH/RTRfkA1PiMuEsSLscbPnL78hiclVCNy
lMdn+5Dgyj9jhPepv6gVrCoEb6OXwHuMR9/HP6BGa8pTwTBlCq+KGf7ChSdwfzRw
8wXqLXu0UrSfk0o4SzHucbFeO5OmXSjFVqdL2BWUJQnmGSKfbCRlbFhvIvqSbCmf
xm5pO8sixrYqlv0lJ4aJl3Esz12RbgnOJjuzduI6BJ1dNnkSJ559amDh8m/W6B2E
9vPGchC8F1qZsBX6crtMERgtVBNnnwd/hU9Y4YrQJdGcpFh1MLX5vQg3VAr4npAi
COJx4a+rlGVQL2uXgljrG3r64erlNXDLidgB/VLm0zm5ifZj9VEmgCYUY+qME4hf
eXemoYx1eWd8a4lPvjQuV2v2VK39OI80pDe2tiDzJ9tb8e1wfv8en7fnNwKhxloV
EGZqjJNcRZ8yETfYvaZqeCdFBR8/7IDyJKuAR+gD3r1slK45Ev55uzDTX8Guunjh
8jWkLIXgaJ6mJfbsmNKDeCQNMRgdzl3i22iNz+T8fl2gV0nnntY3oVqn5PvycYDC
z95t8rqI0bqGYjivxxGGcEL90H2QCIwfOx2irRGaZNbuXSRaAtJXFpjWE10bA/ow
I40Xq41o5/cjG78cMyo/5IdcqWiTWZ5AjhsUwmixPblD8A1meNWO/8A8cClyak+h
ws2SzqbW+wCf3RKtiwkbuyOjcuhJNk5aBCXTzdTj8hXGlymhUo/xAhPzOeaDpJ9j
SB5lKUEkY8HcmPuBtB3xztpXpES01hPLL4v648wjilDfvakRpPJSjbc8Mcxpuepa
4gCeHkbel1Vmu8c3IrIgrD1wBa+VjJUHWpi6SxlUuMOF2RQT4baczSHAjphtbUQD
kmPCgxmN7M0GEnf/vBjHDMRX2aWprIjx+MpeGw3Xs09pp2vmu1wWxADWxffk1/wI
nkyXYDjra2csL/xYv/OzjsebRlXDsCWLV+jUahGs3swZmVwDSmXmUEcsIs9MKSu3
NB5mEJYFFAtWDVgAs8ZY4UoHNQFhwb2eUIZ29rfUxkaTxqhtZV9qBhPauwvpVF0L
LU4ehlAhGQsMYbGvA1In9QLy5WRj+Our1Ux2LDADOKJdwYvY4zuTjvCgexNlliqm
B/J/EuWvR4TQJajr5yxCv+GKnpA/Uf6r2eaz1XjVSzhoWds5rksx44YNOmo1agNu
yXk/2I+Y80PmWuvKbb1NVSIOmd+2TDrGehOH0bgR4LgoX+5Thca5b9DBmcQmipkw
whpEfe8237qVPYlTKE0HLhfi/XBNzwTNMFO6rrvr39vAX7M0+DTqxxXhqo/KC0bM
QmU20aCJAnm6fVj/Xwo0SPKXSFI1J/rand998tedsWW8kE7Bv/jXlxKMcnf7BSxe
fzh6O4pUs2pTsEvIFnpU7BIwOxXLypP0lpv8Ft7xLsWnXL3jQiF1bcokPs8YES2N
mEpaKfrxfgKWSkVVJApaHtrf/KTonn2L0DkEUxfA0rsvCxpaAdmsjxOOgd4eVzfU
0L7QuzG1saBkhDJXc8typNt8nfb2uFknocMdcTEUufln84om+M9zYwwrzNYzms8G
/3dTyq8qpjjM/IDydwcJpXMDT2Yq93DBIUmr0V2BMPdQZ/6d5FhGZhv4OvShAUxa
QS0bTrYVdxKfobPCxTXIZis68a/gq5skuJSbIG7Ds1T7CKGxPNAG2rsXe7U/Fcv2
TpHkM+CMmVu4XC+tDkR1/7Cf5mtykQ+fC8wwBW1sZeGIKfk98OoxsHeuoJ9DsHdF
SgfLTq2bs6RxNqD2qN8odf1lJBl/uh21MJpK0cRlWFjBgtS8Zl1ufoF0WD6JpCh4
n7IjAv5kUf2XyakeKDihmGAS+RXn7S0N/erwwUrM32pklXYqQpwb6lUMPNY+1yW0
39JGZScdju9aXP+Ih4hXv46+4Ojfd1MeaWKBkthv3RWcd/2CAksWGQlLDb2Vv9pA
wRqtyRS05Vo/F8Lb0svNzjSh9PAyaKsfng287yYthLr99i4m4dNcMOPTOcZ9IsXa
Uhr8DdO+zj/i2trM5dxvs4WUlCAvXLW9BFeBZ5KlZLu3sEVDgRoRIWc6JULdjWRK
tYcTqgZ0BpRb5dkEVWl+eiDhYGT4fuiDEXc/uC/rDDmnB2XBWXYQduFS2cIBFf2Y
BDdSXndbPQMTtS1loRjB/mxdnkUKy5vaD9PQie0QO8wMUOYA9lQC+aTATnq/Y4Z4
INGxsQpGJ5SBvZui35LNSG8gTczfq58pzChiK551GVNXxuQgJF9Dt59j95TkX1Y4
iw0dgFpvBGPX4QF0S56wTLwLQ/eZJTkndN+SHC30jQCPcMS18VtcuMqljuh3PLy4
XEWhIOFs1vddUthh+Z8tA8+LJXQNuyj3IujQV3iOlnGAbwIv5yYcROkMwzeE8meB
AUDuOHyKCIh38iKQW7wNk5eA8Mmdci6oN76AO+awuZSuIxIRXUmBTJB9HMpfwGet
Xz4Zg0QITBzjLUbjCr1fnm14KIRORWovMkE5aQRD2HOuDIKT4BHFFow2jD5VdamB
d1gdFr3d0StGTWVX6WMgAMnTGBt/bJfG2tGXGS8kwVEcbO1Bl+KtVFtbwsaTlv2l
0JbpN/WvZHGoq6ElVzbWgO/ZXOy45UsNoujUMoPNnS8J91oOTkb/bEM45H+3npSV
oY1DxHGseulYSzeD/PZcXVURnNOU43HFk9q6jmljfYK1joCLrsf7/BADBG8gsMw7
Katn2RaXhMyrx4TYnSctoKAyr9ekMmKRYnM3/j2LpiK4WgWxBlvztQEZ/JZMd1QL
fxZAeFdmxq7eN3rFQ7LReYzR+kS7djiln4nHHWiR2ds0uljjJhzJ1BzvLgZ4jupT
iN1u3fr0Wv1y9zMlUxtxx7Zja2zcD5/aituga7jonq8+vapKvPK9egN+V8Iyl9m5
Dc8XxXO5hZ+iRViSj5YbmtS43YWDXsEkwB5SxkX46SsGKAExjhmMLUy6hjqWWcRu
NOgq8iT6lPFbe3l208iSwZjEZXfD6A+tcioOOm0Re/VZMe+DTmyy27nP6H6aRJC3
t3i6dyY9VSTk/Io+D43e9u8jtsTyEmPh4iPwOee9MwWIouSzNgFgjXB6o48xzyud
v2rbTqm0M6Sh7BWXojPBDJRmTMROkwpiMTyrVSlh+pgoEOQ5SwAMuuqK2AlYp+db
T6JoryKyNIbbHxJx8GmxerWr4ZZB7KgfCfSMVDACwsDABathppgorZxn/5+/2TN5
SnR8SZt17L1Oxe/H/JSXOHkc04/ZLiTTOF2ybRe1LK78zk243h9BmzbMPxqyS5Wq
mhsItNP1VWHAntHSZo1zvmeSXdqQJji5xAbQh9IupZugcrqzDK9QB6kI3uMGjLA9
Ol5ppXXxvTGyxOpev8xK+fEDzobsL1Q+geDQzgtGIfrq9C1+GS5vQ7LYXcA1Ay7u
ormJVDQyYtpp77vVUwS750DB5YiGPfCnvFWE907Y+Yls0XDgbSOsdf/xvfuRCVTi
7aQyb4lCvF+ouZcauloTOt261w5a0bxMXNfO3ksXzTUBkx5HPHtyVkpfs0zfJp6F
paGq/eo1ZarzOM7E1OjH6VFLY0g0BzMc9rDfO++DIXRM06BTV2Ys5hsbWeI+sSYF
dhEgxMEDWI588RDcjMFDiMDL8ZthLvTK37fDnM4ezHmKArdUoFwJIoDQ7Do3xYWj
DNPCuDG83N0c28WKf3BEQKNUF0MosOzpJZ1K89une3vFWoGUmCk9czD533nSxqAa
WBPXGlQfTSbznap+JcoJIGLRRBAqHLEZS99JD+hGWHcDvww1DK9aV4sVqjN8tgaR
DEG5ancN8dDaENZOhwHo/9SSwSwkQBhzUCHBWcntn52qkcguZM/7LJqG9RZcq5ed
zFtgr1fJwVgLPFjqQzSGiUC82zN0sljfkog/IQpwnseXgJ71h+/0z6sU1IQlyw8q
07XHRV9gnvGRJoWIWAzjPYxUxFEv+DSuLMMRi0u2xdc7aSt9rf2YJfwLTXFNZT6M
32qfV/2DDLEOqWE0AkS0mySUinEqIP235X22ch5KIJiXbEJkt+5bCg8QahJvwDlJ
js2KavtsqfXNzt6AQGFgEa78eCzXH5f0R81PkMAB1EaechPQJpzpiV1HyScox6Zo
nx7LJ+Ln8TXMK9Ol9WRbSUDWHuoLTZiy9TeVLHofcKDiDYVyd1/K0S29w+VDIC0w
CLEDNDx7wZ6Mj+Xtmi7ll9otxTq+pwxCEn9qSja7Hb1C+lwH2RD3Z4kIK4oEuQa+
0Tx2PnYCvZWH9heda3HBZ9slnOoE2xOl5ARrsiFRfLwK+6Ip8v9crDm56IEma/pU
wOMsilGY9ZowDeAuEMnrUM5d2urAW/a2XKsAL5eqIYo2tSFG4A4oBJSedJF+zAAm
znZOGfkPBqyVMovE/3Iq0AOGP5w5IsfzTY85WMK6dc7shCFiK5hb9VdKpW7uKzPz
XJIa5CrJuZHHSMJj85QXM+5KU+fC31GFpkzerIlGp2mmgF9/qFAWnuCWW1FG3NoH
KXTs4BHE6uEZQcm9hGDqg+hkD6A7Sw255c8qWo+uMja6KkAE5jxApC2s2cHRXAqC
kwCBlOr3MgbcJvI5UYhGe8cKMC2okom3za/iZIKheQUXnpWYjwzAiKzx7SwBF7GS
u2GN4AAVzwLDs3UzKNzYEpmXqh+OCIW2r97ZMrAbHeUtNgUaMY62kAQkN9eDuCp1
q64HFN5BHhYgdNv/0da6D/gKqVH0wMyoMdd6lm9ydU91zFGNdRWCpUQ9Dq0uneMx
bVJGX9id9O2Ca5mxphvRq73aSFY+6Pnxhoz+4aJqXo76Y88NvP3vEEptHPopONtJ
U7GlBuC8YD47nQkaXxtf1yrldJfG1hixwhrd0Zy5uAsLJJMS2j6ve8j9V0Kj1N2e
SUVbH1/Y/DDOG7F+nXKq9Q7fhBkNvv+m/W8nW64pbAW0iSNIFDKb8GxQ4ccxXpU0
6t3Nzp6eYHK1sVPySNivHM21Ea2vXNk5k92zDJMT5b2QCHjjGY23si2YStYCRrpy
C7qJAonJ45h7n9EPISjwlZ8SfvdJ4nreVvWoQyXSACT975r4KP47zafyNsBalV3M
FcZVxkgZVSvrv/nLElrnNq3SW+N3s8x+fH023mcOQqUeQCOk5kjXS7/ylbcfEGQG
nMKcIqSbbquG7nyMtE9rt2l1I1RYQD7zxhZh7Az5MjMyNZx64OzZF6Bq691TJ8j0
6+x1691ucI7NRnlNIlrPUNiXvmKTv9U9ldVWDfFBuNQntQzepLh3P8Rrv5m/CK5O
h/hAGLHqfOSr3V0Ma+b7jT+F3Yp0PdJ0aqT970GytMcaMHOMtTyO+KiXsneUamBk
yfZmesRfzPkKaM7NValB+GbrnqmEPx0gmx/LEy7EBpXR7lIOlAP2VRNZfBykivM+
EQmPVtT9s4KTn4U8mMW0Mo3A3sstzkA+Fb/jqc6mURFUPIbMT8nvUvGtVyujP/s7
yvqg10MZAuWJB7LMv3bpm1P3tp5e8Q32PoA9DrQCCS1QhRr117FGGZL8XUmBzkqp
YlpcM8LB8dTYZTOPYOhFkXMMazzamTQY7tpBoxQP4SBxMUQmakDJ/tk/Vt9mKtmX
vNJiOlEQ2UmGap4BTo0pX1L6cu1SV0y/VmKqRjVUVZBhKFOiamNABJeB/oSweIV6
66JEHCPKmCakhRtve3hesUjnTcZVtuADXfQIO+d8neS9tRll4LktnOyExF7zoBot
WAb/QLHGZzbpAGSyyQnvPMjPmjw59Pjcjsl8qik/XYDKILgAHA0SKc/AKqWoS5Pe
SvS2jSqO1v+9TSQ1jT3OeXKsvB3F4RtDgFmTvD/3ja+zCNDa6aYNQ0Nm+XoBtLmq
DuPQWoCDqfIgxiW/LBMPxWp7Fz83m63V/BcyzqSl7IqtRSiyR83hU1Ze7XTk8qfp
dLrUR/XLTTS54ExkXO8luL6P0jwCX9qGkFgVNNPQQ68B5FKcGmb8eWEtfhKs2vOX
C7iHnmKegWAWXs5ftaUFy7b9jWsa20jAVkV1YBPtG6KBx8xhpY8GG5zIiHYIpxek
mEyET/gwgRpD/fviRcKL7ycwPKgBDn+QyjjrcmTfK7p8k36OblHZlK2AMdkFqPyX
qtJiCeh/LVdF8WAopNoMzWTliJWE7eIL4LCnIlej5dn2R0gjaUuULw9wWQcC43+u
ufXcWLlVma26ZeAa93DUC5s0csRRDQgn2IUn9aMUTNuB6e3vb+zcC0fSY+wCI1dd
hnDlr2ytc+HXT48J7qXSDKcGbWt0+KZn8pwdFP6CO6Ygo96LeFD/iViskJic8LCI
O4P11qdraEgxZhEIwEP5keRBv/KDbKubd9p9VhfX/4aGHC+TlX2xscWNUpEn+F6S
ENT/zIJuPJ0V8hWv2i1d6o+c+zLhA0Ub5uFIxHVgxlQAWNXRESD5n+/Jdb2Tpw+g
25C7kJnJ7KOgNzpJf1d/CGTZa3J6aFoHzHZYVFiHDbSsAoq/yylKB9Pc2U4t8IO3
pxuJQT8eyQoXj/HmsVFYXkELOA4LaseZJ5iTnHsssgybcprZuAEfsqi9S8A4oZxP
l+ZKU2hCrpMJndGNZD6bamkMmxybgBkRm+Z3DYRWClKVxR/HwFQIaCoCcj44WaNw
PJpkU+xD0s4hDRY8DM3E/h8hp+GKzHbZIXOJY/1bfHS/FN11PeMGOwQWr69UP71I
4d886+SpJPm0XBNgxG4NWGO0++CfV2C6ehli3tP63P7yI0hFN9JjaLm19ggqD/40
Os7vfsa4DG/WC8DuiQLkKGLJzI6yXJIsTHevky2E7a5NkCutMf4ov9DjjipNwSAG
XuTHOHORN++uqcwrELsz8qvSyf7byKLvGb1lAHOGKu+jAPH+GkDIu/2TZ8VGXzDt
L7TGEuUCOTOAvlDSpCUNpILA0c268s0FQIfdya1mEeGNwwJB7gg2nmhiXg883spQ
mbGHzoC65jojeezU4XPRKSt/xc8tA5giEg3rsJweqThNr+1VT1IkbtuhvfRYNBP2
EsKgKvwk+0+5uqQL3Q7niYS/1iqz7Vxjxm/MEj38slht4/7ttWj4WwRdjqpfI41g
yGPaxo75nNeq6blMVStnDm+Oz/MN3fmWT/aYWLOSnJs0lJWWSHPCqgBnZ9ewWis/
u5tspdx+IUOsuBmdZgj9Wf4B8pJP/VXTMLnd1VA31UT6mPCmg2b+69ir4+pMTupK
IO0gmMpaaH7RVjxBLk95eFGNI3HhiFHpBDFewZyIwWUnQyu4q0bP9ol8adceP2vA
6M3xK8Iu5/TmRTwmmDPT4iHhfwNf3E9aMSEBJtk5GGQ7XOz/Fg5+Q2PWbSM0P7EK
yvShLIcCQmnXDIQZJAHpbThgPScFdwyQ9YthWsdZEeE0IH2bMyY3eeQ8WzZKhEqF
OfzITlWK0PbRMiYTG4MluL7iaUdUr+x6zDg4V5gVIVTedynUOvqHoVa6w+X7xDRS
YpimEWNhH6ZXq7wjKLDzvU8HT3JVyVHIDm2v+UfyJ/dNkDbJ4DKu1gVFHc/pHGYE
nOGRku2QljM/Lj169v4eoytMQ0ZJJ+y9pA4CAWUDbW9J9okx9+YJJpFp47Vrk+9J
G45PLX/8mZ3hgtvvoSkWfDhsAzLT7mTRabON1BigG3uXWFrzpW8CYGShpGXUKiZl
gH3ED6fBldXjgZSXQ6SfoW+6TUvAzJ4qZ5xpAyMiNPVPi/JRg4QqybHZk14chL9a
WvBkoZVmVI9mm5dEIj0JM2jin6m8UOVnyWgec0o8xlCTMB4W/P682pdTgVHd2Zic
07oGDMhWtixIuhRNR/xPeU+K+Cdh0ySAh5ELu8ews+rYTmZgOcNpzA9gh8O/FOsc
wHzPed+JSn1ky7q/+r8W2HCEsxnGiiC0Wouz3zKya7ElwAuY8EDEYWhMNKhZVaa4
a+IEQUlcpJxwNdfsgpBsA11M7pBNb7jksTVZABytswkEePbFv2qYKUr0xhT61kui
SPBTTyovdeQ+v2+b7owDPeNHEXcMwAf1uq4VPeP5n6fxWeTMz64UEcZGDlu9EjDM
75yTXAuchS1Pl884M4GZw1e4nFsLLxq8746+3XIT48bwVIHbpVWfAy5lE924YY5J
/o7q4Gp2xFBsv6QcvQ0f4R6Dc+ajekhWNAMLblyJxw6bcRMDuduAQONPtzUPBfGy
dfbyDNC4cdEiYno0OFyMntXD0Qr1Jv7JjXTe4CKRiZZkPbV5FsiDJcMXcI54u7aw
bYk5GY/WAeICzMt2jl7rJfJqkBv+NI4hNmak25WvJRx56zvauVdoTiP9JiIt0Wcf
DZnhQMzE7+oiudZ9Zw7A9jDw/YMsQkVjZRpFuujE3qtK9YaQW64pAfeuK0AJtB2J
HR1B07V3Qk/re+YOGayHTPAxsWlZ19rk7exrBz1l6+omD1R5+fccggPhTHkEE5W/
xpqg4O+Ify7pFd8CvVfRzl0PiOhScK+kY40f05E2K+V4cuI5xvy+ti343tFxOIob
vlBJv9OjoxtGBERV25rAFCGBHzQy4irOk1Kp5aOawNWV8qZAOC7GO6nknshjW4OJ
sAzKCNfJs6A+myHbMSdsivGBFYMCf/7eZxHqQP5fBbiDzfUD7kgnWtrJDt8ch5kW
T80KXq3KTYSZyfn8M0dF/GJkH43S6ML34tEZXonT53ojEUg4D3+Jz62bOzQB5pcb
y7bjVuykoi57RSy+Fku9onpmM3y1LzNFKzJ0CeWV2smucVY+Ur8aGiX+zuOQhvcW
RXYFnijDbDR3c9xC7LjcBociF/0hqLluKML9CmJUqdJrgAUa2wyTLaNeCygbO9wQ
I1+VXqQMRYTHHzDxaOnDOqAOmQK1TjTPwE8NbkuN81cN/oINwvGIuDDP9k6JzdBP
ceSIE/D2OAAt/ODTsXB7a3qQ+1fuoJlOa74vF7/Jy9jicbcO3jZsXwM8USpb/d0t
akdK3QfSk5vBrqc28VOLnMjh8jzWog86ttZMSXnYqslmZZIR13+R5yxvntRc//Ds
Dj/SBNV4gfKW81woZr5IZ0A1pbLv2qmBR4bkMMcFIKw6iUKZgLkbwAtbdKgEtByp
skg2hFUQVSKKlyE/SowNW7tNmc+ZAPcoNOmdbKGXtLofQyg0zWuNfjrkyGLN+L0e
mw7I3r579RnA0qWSj7mfzdckSMtw0MppEvqReFb1pmFxR/tEgNUvRRvUc8jkfa4+
ZjGN4g1QYQDzDBsB2gJKx8NXmuHcUYK30YNCheJF7/zJU3mthPzlAPtnREWJiQUV
mK7ErogKPUYbOWCyoQEWyzdKhvRkrBE6qiejQejY87qxLsliGfmiTEXqBDNBJGQf
j+1WM18ZASK2eAiFxoRAyHgsuqp/wpRGzHrXFgPpBQYTDV+RKJKY9vV6LQFyyMZy
D4FbSMhFSHKO+rGPOxJfxWFTl7hrHohXHajMiRiMrA3PzdCYF7aawNjIoevjQEcl
mpwpw9O1comVDoc4Fbf1g4PixAAHmeA3+0+Z+YluBDr4v5JrabXqGtSgS3M00SEy
HQ9r2ISdPtUy2UR3M6TZO9kONCfvehUMFCik0cdSlFclSrVM/KC9V4Gk6/JiH0O9
A3n5uC7kjupHyNFggsZMiE/CEAVtEz7uPedBhLSD4DkgXSg+Q8+HwPzlrviH45kG
DXI2KOYghKgARiwpTBI+q2iqiqWlD2P/iqgjPKyVV32ltLx7doVLdETCpWcb6v6W
l0t7J+26g96y4jqE2tEnbeovvkidW/E316pi7u7Y4uZNCP1tdvQow/vwa7g85FaI
L3bQUfXIMvAmgYDdY8ZVMGlh9+xHKG9abAbgsG959JBvE7inDGc0Td5TlXQZtX/z
+Bh5ljtVasYWBliQdygHV56OrlBk1NTjTKR09DW6gk0Y0xw0MwwutcTw9DEtLd3e
Wj+DkfTVDHzY853pb1sAK4VwsIZerm5mWh8t7TCMEhv7U5o7d5R51vwt3Wflxbpa
/rZpOAlxGGDWCHZFZlB1FS2T7qnVr4wDzHKjqP6T8s8K1jrwDxWH5azQlR4lbpOV
xqxuqiYtAkKBpJBy444sLPlrifsgNcUiRWjX9eIiBH2XdPpsrZPDR1IHNO/KVFpt
2upt8W64+VapIWwnyUqULEOgnjUfZP3VoRBtCaBFjunMjQC8TSlcJH7kiBa7vjD6
yJgLivCrmh87fYRSmwx0/euUXgIioXJMmpdwMnUthLv/0O27FqdWHC90hpkWLNhM
DFo8+lG0cc486cHyV1GFp3nTtolmakMCPi83JW0qXMnAayxIjtNUxQ+FI/hXAUp/
7TMeiR4MuWofSvfXTZgx3BU00xLcKexQQKC+eNhlOcax0W8Y+sq7UybyRFhcbnJ+
wmgNTl3jLTrmhHpyxcEXFnk7ZddYSyB6dT3ldirVkYTdimt3oSQZs1IkZqU/5XWa
/ArN/sPhHFWmB87Faih+CbSZDLuH51eEaCjGzB6VYfVc9VqwMjZ6Ys3EGZVcZREt
MrWuKlWFZWM6SLuz/xBCHcOvRs1EROEyHr2cVivbSGqF73Q2fivk8xDcDAeYYBlm
w7r6FiRV4BcMKfvDptRSC58PUMUMBzkE3W1UCRqQlHTH4uA5rxkYXgVTq7CCB4uU
jvNWe63nG9xqqOPqbh2WiujSmlXaTRz0SZLtlmpEDuhDZWTP2LS56rRgNpkXit9S
hC7XYdXZA74ZbcWFkRgU3sxkS0EuaI2MvFCjWH8yRR34wGWqgxqGqThAip0O+Up5
A5TFVo6qLvBAklg6PD3xMfGoHQRf/3pcxREcfqSRvcqGGO4qFH/sNgX2ajtm7O3L
fnTTDh/U5c69TvEhHK8N1MVGND4aW5+eeZxfitiwRExWkXtAz+V0iIk6J9cYbUbd
452ZTU8dqBJfJIXVtyY4InMLzptLTpgP9kKmWEn8sSdUOAc1KehnaLSVbu7vz+c3
jEfYbtc3OosMdtRbBkZ5+rROvhY3IsU1/Qep4IJ+Vyk/4FChyrOD9DedBzzt4Sle
S5EzEoD+QmtVR7qWEfQh/Nfo6MAZayBCXx4B5CeaY3/2XllXQa63bd59FBDt5wyL
YVlkl0gcx8uoAzUZuPwLWt9pb/m4tvS11mfZvXdllqhWvApc4N/ZpC0a9Vv0wLRh
l9neB/yx6qjntATB06298aIIXqe1rKxKPcdHRS6DOIZ4rr/FJo8l+lMg2j0ZbAsD
r44IVfUMjHt3VAbAR3qQQMstvlfM7puVUZtt/JcFAGrvlxeE0rbGbXl7Uu5zZtud
kSeCZ3w8uNHwkgmsApsk3RjmEYhJcz61Yu4HdyerYNj1/4ctzY3RJZeWfLgMDMHO
apMBdEdXS0G/p0MBNsVhyB5OdOm1ElopOTULblZgE8tUqk4La73dioPFBJxAuKeN
PP0uWffDMQryorajDrEBIwNRMvHOWrUVi2I1ISB1xeh8vdHrb8M6erWa/LnfKCCe
s/1XUCbIW/XPxMI6LL/sYrgTUjEQVTFYwPSqaFN6uWsKfn7uW/gEbA0ue2mDMgph
1smwChyR3GCMrquirbYPe/qbSiwfEaM1/yvJRonbOlj9pYwsBdIuE/Q+o2o4FMHk
NpdlfL5JPCdKRgNzjB0jJtx89UHSYtaixp1w5Qayyj3JtdzCqTzB3g3xZsjelFqq
YXNARWJafnbAH5VJGhRkf7P2v6PLBKIywEMmMn2yqjPUtjnfpL68EpCSjhSL0PJY
EasN6xkyVjM365fDHebVZLvyp4rAaTaB9gVwvIWdWY5lort/8RsxiN170pvPHIiR
p6XETIM37zweo/V3AYkt6MqeNirategQ5tYn8XLY4dNQIxpkCWX4Ymai0NX9UijJ
ttmlv6T8v6aeFaScl57SoVnE/VVnKkw8BMAPE/fuXBXFsL3/hrctmhu7zmXSh5IJ
DY32TK0dMCF6r6YPdQ7dRw2oxlXFIVFFK+DSqe7rPdTjCMoTAuy+VjDZERDspVrd
IZlJgd8+fn92HQfFnpDpd+VO3z1B7vKNPWvG8QZ3T7JKoYhJ3XdhFq+/yjuR87Yd
+zX2h0zKQmdXoXWk2FjjHbPdXDSRniacbvpMuxnDU+L42SjN9H2KoxTEMxguh6re
e3KZJ4fh5WgJZzI9iUzrydig++yDMrGJA6Fx2bZS4QWIGllPWOIuvWhJaq2NFJOU
1rvw1C38SWNE4aGCQLApowAypAGnNiIrH4LeUfBHXbqGxxM1tpiGn8GzGFsNFjkx
Y7x2XyKDGr6GJZ/ImR/mJer+D1rv3hvqJUXqd4F95oSArx/SF3+WwlDuja/IH+ei
YBKbD6KO0+6+WF9QFYzxEKGg2bd8oDpyFIo9+5FHj7d4Iv2R3oDuY2x2cN9TeNHE
VdjTR2wB2LagtVRFei0tWqsvZPHpGYTk2qw3H29g8bqw6LpXYXkl9c8XOjkahkew
Fji5qJG8M4TjI2UwIpYBhRXXYxQeiL6T6bGv+zOiZqebplYparpq3bX5NTziYxKA
nsSeHLT086LjqWi7ysea2ahx374WxZ/rfcLYPXdfMnSUIG3rfvDjziidC32B7xei
PWqT60W7+10aJemEzhIUZZVrPQRwNRFlKMHFvdameMrPY683Sva2C4ralStGweC/
G6Nf0JZYCYuBdPsqClO7VjL/i974zPn2qzr96PKXE/YNoYUeT3dhtsyhi5v/gxE2
Z+ZRveZoJKk0c3a5O19dBTYXr1h4YrwrQ+iK3Gym3BYH3IuRbWNO5OFKJGgthnOs
N1wk7g0OEbm7CxqU1CkLp08Y5Tr2Au85rN/yY8+2GvzSz5aDjuT29mtlBmWrWUoL
JN8yVR0cO7VdhBcV+ngtimpmacBsYtBAlgzrSo6RDO9D+YHmbc13AXP0sCAS7wO9
p14SaQEG74wLY3mUnoaQfqThNDbCM1BUe8rQpytt4TfmPnIQHQvqkZWLxEhmozeu
I9+TMQwt+jnamdEIFvjFrYVabIODGxgHaAV01NOP6811ftWc/qF9wtbvwFaDZAM3
0I3IcWLX/2257kbLL7iil6iH5dTaovgEdB/5OXETexlc397PjfpI4cP2rlvd9I2J
B9M+kn2E3aiEPrWCoBkPPL36V6bZdvwkZxp3C0THfwUTRQtE1U0G1IIE+2axxUhy
yKJBg+MI+XvUwCqXZ69btLlIJTcBmJ+fht2x8JK6wUBvkpfxnU+zmwELvAn5/PxU
m+AUQCnMFQnKPuUx+M7wfl9Eh5mSO+bF+4rYngU1wditQR9onZOq5Xm5A4sfVLLt
SCjS2Sa7Jhz9etHFNdyzjZyTaJ/slDWD0iSjpQ98Mf+Y3nit50c5ybjMrz6TOTPm
bvIhA2kYJTY/AwUQrM3zy1G5Ocx13CH1m2sWmil5yoYjHerWX+f+5ezDyZMxVn+/
Y6aHmoyr5k553+W9Z3PdvHaZcnog6SRsC/JQ8doSlKPuF8gFPIvTQbCyqKY7KyRc
1lfqmv+PhKr3mjGXz+N0BSsuf7YXgwUNwzYu5zme6nnNMbI1baZ2/FW8aXmAF118
7urvgo4a87Tvm+5d/AUEX/uATkG8yZ5aC3azWfMzSBabiEWfvW+nj46e80YQzS2s
fviCaFkyeuNholKrZ0h1v4UZPZM3JCm2hRXG0cimkBvsUpsn+Kd8XhbrUlnULIpO
E90NesMLZ3mkIBMHYaQRPka7Sdzroo2fWF/XK7IhMjED0B7oePrRPfMHEyIJSWT4
Yet2HsFbo0OKi9U90THEtY7F1oaQ9pOTnG6vWq72ZjHcsD9E6POM9UKolIT6dDLh
FsnZGyUmaSqADOC6tqOsinWO97o6UR2yQwnNuF8/lOo1CwCfia/9dNRpiMVZtZ6D
X8wxqDPYoqxRFMCxI1SU7Rjl7wssVUBBgxubJwv9Qur0FD6Qk1B08Op9+kLa1RH5
gzGo5wNv9fv8mBRmZMOrWkPi9KOxxz9R0KX58+Szwe+YngP/3CTBvpuKo8ed6d9h
/1a7vKBajgiCw66SR8mE7/L+Ambhntp6rdZ2z9/mbp88IQ7GPFsRWU8YA3eQjLz8
Sa2JW+udbWjemLHMxvSqgtXU4Re81mZ/bF5E8YO+qK2PuuILI2mcCTuYkcm7vmh1
1/kH1h4KF3ye48xupnzWO4AqI/QgMnvl4xniD/g4eh9YlSj7EpvXr0LBeDTrHOdo
nhZeA8yVqPYASR6Nf1Xfi4yXsm14ytvkqKx1UfcorkF0H8qNtFWpPskbNhIoMq77
joE+Q3lspTed0F38hGD/V8BUjF5GuPqC2sTSyWv4+5om2dn6dHjQ0ugPU6kBdlMu
zlYNsAxf/twlMsgdIQXxVU8adGCpDnlW1NqLhSN34B2h0RGDx4YsOqVi71OnvEoj
v29zoz3NuSETHaH+bP0vE6MoLxBQ0RDRjQPIAi77Hagl/DbbG2YnwV9I/eDNADb9
bgO/haNwny7EpDjCwnPtzbxmp3PYwf65ZIauN8wZJ3WWCBboRwWmiHW3gBxL7ILl
DMBqdFFC9g9dJX3/z0l+pf4gJN7y077t+Ckq3D4AaZA1w2X5Doz+F5MU1F9g3tfo
D/G3lVFtimkhJS/RW6WH8LRbr995Dcucn/8xvAn8y+tXx9pvk9Fg52tvjl7z5WUl
TGTEDJQidGt+gyhdA5ocl8Wj5LxbkUPHwxns/qdgqYdJhPlJvo48WENT/IulzRXF
L8l42jAVw2OEENeJiNoegVmgc35s02RK2sBqGHwa5O2VjqZSJCbYiNS+iLbrt5OO
vukN7Sz7EBVZaYclAoyPmQsrRlS1iGQ3HK/Rin/SHwL8ewWljVLhhkXfpbZMcuN2
mXbzWdQJinqG9DtJ5ORuAaEWvoVBXsw+hR4UKjEB/buOkPUXTsderX/GWZ9nnw9M
+NEWq3Zx3wSLTyUR5OfalFJJocqVFtM8k0xTBYl0BbBFQzILocSFYukaOfDT6UfL
JcyhqDpbbYDvMjeBZsYecrcMBVe2+KlLkurG5zXQeBcadD0wdJOg3xmb1nUe687X
e4erc96hwM5g+MImlyor4iYiOfTZBAH4AVuUqolw3HRYcj4jU7kTImhNescARACO
g0LlRKoQWx7r/NkTf3RIYIP2G8FKhwF2+IwU2sYUV0HtO4OqfbXRevbHkp3BMZoc
7k2tLhJMeBeG3eNo+ol9KivpJK5hfqS7UL1pZjo3sxB07EBzLFqmTxzKNtzUwYQf
f7Zbq1Q1SD2TbhxRQlFohvzj+ASEz92LIKFwv8Iw0LMZXM/Lcbn1c1Q66xFsuyiH
6gO5TuePk5jJkUsFzkVYbIYOfqqE8Z2c3fiqs2gEl+y3p1KL0TSF5GB3z3wimOho
9WZhTrwPX6poDMSBqSfWPYBd8KuzOonLYwOla154IjFzbibvizgQVFqLCM5yoehD
cN2ZEw/34Pzb2ED6raQlleSd+qLUiIXr8l1IYWZcqJUurh4mL1xC6A+aDLsj3dlP
DYHNHf45UpkxelAAvAbT9iJWktBrJjS/YripA5VjHELiN0YKIHOmvgM97qDzwvnP
vVb/k04bUkd/LtkmyeThDjO2zLunZEbVMriwL9BOfUDND2f0ZNQ09rj25SQFMlG2
3uXCJM8mCij/EGSLywjtdrugZFic7qGRovOpNw7pB0J9UhTtuqdH2mFfWgvIH5D3
9hV7OvpZyY6TgJ1sN+i8ccMAF5IHgQCEDGYx1laeIhPNTHGjW1oQ0ycOu0V13XwB
MEAVRby7mypNv9iQpdFIvDS+pgSFoZyk2r1+Pf58jToxFgxLXLLpGmVR3zaA/tZr
1uFOlK7malfVi5zKdkNBuUDuNPtSOLQDi9b5Im/wF6yP4La2Vl8y0q8+wTtdyyMb
WOuRglRjDaccuj/UcOV9yPm7o3DB+ZTYe6y0xA15LnE0CeuoP7N5zU16E3AwtZOx
6b4+16uT67OHx/iQqCZcFMP+Ti8DS/7fSAfZ26F62k3Hx0NMpPl72MOoZ7BlsED4
rq9+lOoWOXE9D1YGas/WOb+ZYXMk65/mnAgmtQeIertffGOo3DiAkXuvagJ13jnI
fylhG+RAE8DL1HbfFOcqp5/XBa0fFcPXiGfZeKwvto3Ml9ufQa1Q/TjJ24vLI3Zp
mFlgjVzqTHATESHxhU9AlO3OeV/deQc2lXRRRAXeVCbMo3DGIvu3ggD9gCgAV9DS
54GlJfISCUCqgjldejGjhYA72xnNgw64ASZrdZu+JCzKuuRPuWHWadDJ4AdBLm+W
aVLTGiTJ+w5JievbqprBdMYfZCLAdhqW2UdarKxyJii3DIMtlh7O0Mv6mmE994dY
a84+2kXr68eR56/9ihOr0eFieiSqZ6Jdz/ZO3PdktGmFNM2oWpy6uiguTlYQlZXW
Ds+UsXcupGshxEZ/cKLA79P8LgAxbAHgYJniuSIRBJXXBd+3kW+HYqoyEIecS2oh
SPIqXYyU/MuGr6UHzkCQCdjlUhIUi5Pv7/4mXEfqUsEWXuhues84nHiXqu68OqdV
fUO9JPlf1zC0/9svsL6NwBtvJ73DX3BR+kWnC2npyWgWspeiBIMCCiv2vXMXd1k7
kVOoBcpuE7cHkspQ2rijAZkUkhh9o7eTo0OVrTvgTy+Da6eE3i6FCdlzFwRrfeHg
5Nk8izFaAvV9KKiPbABbP64xV79Ferrg062XCBMxp301sms8Ky+PghMkTPV9Beck
ZCU6Qv72VYNqg8Esa6d7FUQoFvWgSKXhF9tLLDDhf89pqbajLqTeHFqHx68mwqVz
MZbKVtDdRnJ1pQXO0NaL101CCpBKusCIXJa2hOauIWGmV5Z25Exxzy3k/F+I7fdW
ZHhqrua5FJxFYFZULBNS2IcmZFcUPEp6fjroi3k7r+O7tLeoLqMlr6fEeQYrXnAG
Lno3VgDZsHyy+lvFZRnM+ZQunl0UZ0HNxtwPoH9XrrqZhsQVeIOdn2PYJTD8f5oA
pGQWdnaBLeOIKftuJsJ6XQpMDKCvWOm8kjNH4mY7AB15Su7MeEksDGN0kBexzx+R
AcaYshmq5TX0ug/UOl8zI1zBT7rBJSwj+N2IF4hk9ollr4qljRs8Pk2oadxEZ8MN
nXVEsnV0dcR38a6XqVMiCDEu34cYZ5qYxsSz7a5/exhhnVTFPTkLMJbkvha2hafJ
yY9Bm2NZLbGHNvGUAQ+hdSuPeqW+ziMn3Kuvy6sqyuJzKvNyz06B7BqlH5nRH33m
eiS4Z56ek+2VJvAl8s7AMtmGm/bTuwXKcN9/oEtS6omEGhV45TF2vQWiCeJOFSOQ
OwZJTsKplSiK+My1SA3+frXMkTwdjIsoFJr/347sgbCMb2MuWYJNGXpti21RZBVh
MGP67WY5eBoWkjSs22ikZVqpaGC1AgroRvIndANnL7xxUlM/2BQAlqMxRp8Z7NKP
zvMmmZra2N7d1Ps1k06GUmfD2pd+p01T12jFzi9c/kVjOqIVIxrCWaNqkZTcOa+G
IVHbvx7PItVPx3f80E7rZUeOA8cGUivn5KdJdFel3s6A7OXrQbw4cAg3HjOKS9xv
t7pjnpKaagR19Eh9oDGOi9blO79z9520XKPOrtdH83ZT69ZIzJV4nCqkftruM+sS
Lg7WGm/JtyzaIRUcS+ifp7VOdIiTaAGx1yOEkefR8u9s6YPBcVCT5etZM3kTz6o3
z/nS7NVYLHZDn0pSDj/X6QyOIo11gx5N9DHCiYIP8opXUCJH75wltZ/qSowvaE4K
I1jsonCX5MzAjsZnz/gD+2Sc0F9UPDOEKk6xwOhSbWrhjV3+oDQc1c0PY7C47Viz
yo0uKzYQjy8wFJeXrHxM6NxUuLjQXyML+35t5grjwQWer0UxKrQSX0jZq3taFqZQ
pyQt7ODDMhsIMTF9pGQYTgv7DPtyKNjmcEDFGjvykMAsmg1+/nNX+Q+v82qP8lnf
rtNTGmmxdE18C27X21uHnvlyug519siaOtSh571v7dSZeIjSByod+uH8+o025kl5
++TDeePOWpCy/MSo0FHcyqlB58bCG4mMgU+72DWp2NIc+dTGh6eaghz1aUrZTeJW
CAoe1vEsHFcSAuhVb6ur3qDDBK0RV5G+DSMVaCBw3I9W43/Zh28ZankVMaYsme1O
SP6UgjxCCpzO5nkWO0qsampOJWxj9J0W8v09AEEHyEREEe9TSxAVl98Dq+vWkmmq
y/fmPxnzNcEFNby8kZEoWi8EKA0cH0z4JvB4PeQrYJGkVX/Vk1cF6s0GjLb+a/Kc
40ltlBWBB55QAHCdDYv9WHUo7HQ1PcsgW9toiaCluE84AQsBwC5Mhak5rhF5xlOp
WKibkCnYQUy0fUes4OOi07SLUB9qpqClb+tevXhm4QTKDQT16oJhQRKnX3IoaHLC
TCVCzUyeTMhTeEgOOEwTwemGXKdo6dX1zO9IIYMqMzoGgwHWrrikBLHYJxhdk0Pg
3g4WSqw7Uhzft8DJxaNszKgtcaLOP+mxDYgCwn1B+Wh4aHsbcKZRPGUnhOUM/sQF
LhiB+EuneiQYlmPwxerJ+7haEeDCfoLA1QAcZFayuY9SM1Uty0P1LranMh2hGXM/
6iy8x467Hw5uI1fElUozcOqtOdTKIwR6nAhVQNTWakTURjEPOJBcsXDscbrg6S4W
re3hyrbEbhgbgE/AO7MkvAXVNT0bx4YKxnQyeuKcCEOuqZEoPhfuaP7swkPoXzMv
Md2B28FPNYy2PMpWx2zpeN/si0CYO06nmSnDWaKjYcUCnyzTwNIlbX9wbNpGTRaU
zk4OF3BBEZNlM2eriuUwAUMLswDKyobnnMxQl99hbj7e04ZCXJtZ8CT73jmBzdrY
mRCPbEvWrXaAyuT2GwG9q3H1zzFM1QrlF9k7tgRf38Z8XMXM8hVe7J+/zjCl1vxl
FyYNq/SOg/yGxOywynlaPRHbZtKIAtwlQk8JJ9eLZhqJRhDWzJhmWXvxUUMA3eWQ
JeiyRAUzJLLv587syZlnHC7WE1fDtiwSRcdTiq2P21gW8DwSQZokG7fHQ0T3Cjpy
1thyppaDjWeJil4A7QIFpC3RgJ+8EVTxQ10yHT9FsquBKttcj8ObzHWjWcfKZA57
29Tm55aBfjzz0VUTaGaKOpxztmaOCM1OGB/SQCqdg+g5af0WRYUoPWP5wTJfT2sG
3U8kq+uchOWQKKpCzF+G/IR4KHmrElfsJ0o1UUedAqET1Lt9AjX8dDHL66SAtHvD
PFwAimm3tKtoxA1OzQj9gC/nXEt9kWvZ80x+02Mo6CyCDBMi7P1vIVQGqpam/dX8
qus9nlsyIw8ptN4SvT+sZsA4GLlNwHJycJaCZh4xYZ4baRCQqTlwk5gdXqGy0v3g
dsaXg/z0Gjdp1H+1iKMgYxjZXJNK2vdqUxYtGBC8e5Emy6yeVtWmp6GGhZEE/Jvb
Z/ADf6v5NgbNa7VVBO3WrtJA/02vvCsG5D6v1MKCCTOJIRdthbuhRRevf5ll29w/
khO+dh9oOZYE70gMfxLy+BXxJyxocW5dBRsX9FA7O4n2fgh2vlTcDt/kTpoepx25
c9Gui3PK0isY7QCJa0kJD9B5Ud9CM6SkXNqbnTUO9yzPxwgbpOjL3XsLJSwj6lZ9
U4xZWfhr/C26dTbjH8+xWvDFOJwBaFdwm5JDKUUUSV+TeN2XMKQMO3bGqFeVh+8K
benyGxec8fOmo21mh3/mjC3ZoRKEKb3sottRmTwsZUBnna+jRtPoSXmVpgeaa3lI
JV3eWa3F9z7FA7fvcH6JSDUDlzAXRkCMMOC3A/dqZFZ3yp1k4Ig5wGOtQEwMKC93
TOPpIWytT3q7S7/WiiQmNeVygQ2hIN/RUiZcrlGy2Y33ttvs1l5ODmMvwnkp+ofF
bjae8VlC/kQ46ohEn/C2rkrcSisepbYyo+R0AJGxi9IXqKRDVz7oRlnR6rxf09Mf
lJGQ34JdPLaJMcomCY0+0oLhvwVJIUSWapRnhanRGz6yOYfGc7m/LLMdaQXk8T1f
ppwLqdLJ1mFN+ZMUXUVQSnL//xRywXJ1APujSxUp4blUmmtNNjsVnyZ4qTYvGuuP
acZfO+sxfKXIxjbC0yDeWLg43NNPU6gUM/NjszTNoJ4WsMzLKlLHG4RFLIfj+g7E
cRIbrzU20pZlNCGAZnOD4jm+Hfi4bc41j8RWzk2V/N42N5HZJfGBWxumN1CdgwqF
gbHcfsZP7wOAkhTp1M+l6LwR9vrYbcBhnfVkPjR//K9SdB2LN/5FlixgIj0Q0OEH
dpXPmwLE+AAZZCXo20bwBqEZ6YZ9tmY+2S5rhR9EdSyRimKbLgj7p3/RX9gAza9n
KfSeRufjHCEjbKU4OBa+MZCltfgCWFCOndPaqPpfCxk4dH6nVhehnpdqpnptWhOb
I6+RYskKMZC7+oaxzmXtw32NHQBihcA5z5BeGmPVhQr5+dbDRN/aDYIhPip8YpGs
Ncunef1ICkChtUG7/kHGcWBqQLAG2tX3SEil/RbbCVjLRanmfeDT5FWDCxXXllu/
bq01xDNIPu7V2OH1bWyrZVRGth0NXeUS7d7/ApSn2mJoA0Ep+YeIAwxRsvO8lW9f
TJ9sy7sPvkLzg9j1eH2caDR324ThMht+frffWkpn3vNC4Pnsg4Jf0DJ1Ul7jCVol
BGTSIELOSQjgLfJji/uG+BiayTCzh59qxkyCSw6AoUkKinU51GIJ/mhrY1IspUTN
nAVLw1TYT3bDPEYxb+0IDnhIrGmc5EU8oste9rMuBjXfOKGG9poG/h8HIr/tYcwD
vqdPbOR+o4jROxsVlsH3sJR4NWNJFfs7IjUZJjWqnGRh+iPZrZ1niwLsRPyPR4Lq
+rMenaJaqhZR2jukWNdHSGnadGLKSm+GtnDa0Pb7j2SVKP9l/aMQh66sdgo+Om5M
65fB17mTu6c52Lc1NIp/3lyV2E0oLScaM+ZdVTbE5GW/JNHzqffZXRDNGVJXh6RY
mv4hK8Gzd7F9yXIEL6PMz4Nsv0R/Duf7zOVLrzG8uB+AKPclvqK5+n2RB+q03uF3
0xunkOouinsBlHkbZWb710hXuE9GkGTbeO34HMIzankYS6PUrxOQ9qhiuNq/bT+N
vY8ZcIy9GMteJM498cMxgAosx04kypUECUCs0Iav4ZCJtjKxo9vL0dqfXlhMcmbn
gzM+1UBZn6js6tbTwnZYQgguhxymDOkuK9AcvieNUzSXAw3tDvdJMkPInYYD3Om0
YTGzy+wwQcD3cFto6c0zWsHsNZa4e7ezWsM2C4XsPa5+EfcCa/vPtdnjlzlVv5Jn
3+te05peXIQR6hDOUvP1Bgx1Z/MbJLyUEODM4f/GGeIu6Ufu3OYNQqlOyzU1PjU2
fwVZVmsGgaMFhRsLFQu0W1UW8hq/yYpUlRrnlLjyJwErk6LyXWEwuPK/2UoGRzP0
YEBMq5hUoMDqc54MN1KrQwEh8GqWTO9Pujhpoy1yPS7mnuVh9UA3ZHMbDhiP1KYn
vzNfhp/FhDmX50Iy2x+cZ4BximFbxs36/iU1s2UudDZSL2nqxp1XBq0g1ocax7+n
pNoUmJz7JR2n0Lh59BKh2tYuRGUStafjqfIdia+vcSST1/uCRcKLEJN+Kbx8HA5q
pN38Hx6D4sfSdSrZhqnXB4xKCVh1nZG6e1I49Hk1aZzhOy1F2YyFQboS786yjmqg
lf89Ssr6o6rkZePBkzl9qHGe/KMVLt8sjXlXnB0yDqtwkGs2HRPBPZ7wokPSx8sB
DRpB9V9bfs929NcQ1IVEObx8Wn16KcM1hikfrUhKYIgwOWTugeBLvKwz0wIz8PWR
Ivv4jBJPUR3IauqX+zsqa5K9kjsAxn9xLuSTtqN/mI8/s/9IYqjLCcyf/j6PBNbO
mSB35zsAWcEH16eaGt1dtFxziu/YuZk3FtgWBZeaphfbpvC4VETbnwX2FOrzk5xd
MUoUt7NZWlVMW/7JDLvE8ozgkjZSTJzFsHETh0jt9jegvwJPWA27fX3LHiCtwMNK
YjBX+Tu3q1QkRrbbYOkjYNIX5KDdP9+PpFAT2hVBESqg9ov71Ob+W/ediZHuTZRI
uCz/43CgaBYNP+0Y6uRVoGMy1S6f2oIPr33uGyriswxDvatK0Veowk9X2oF3siOm
swuZ2d3GSx2fAeXko4c97C0pJZiaZwXfWa9yud0/iv4FRAJxkBIKeD7T7wLHBalh
SdyVWEdc55RMK8KV0XSKdH1iePv9KREn1umC+VN/a+AgFY4pJeV6hetXM9Ps4hqk
gjvN+iCZmukTmZEuiub/J5npmDM/TCjjPrbNt6i2bWTuDcl8DaRe7HZO7hMAZ62M
0ESZhHFULIlRPiWBVXPxPX1QfqEE1YO1RUGUBpNziUlg1GbBlRcODlgYHcSccYb+
Gq10MasBrFIEeO8OitD7ECbZTxP5aNoXEyS/Lc6vgyNbVPBBLHll4tTUTYVgQrm6
iK5r6tuALBWubkkDTdWRJW8HS/GQuBYVMSma2mWssngtrWy5KANB8+PV/wGfJuK4
tWoWpZvN38nCEzJwCh7E63cAXgIWU4g/TOzTEeuyVCm/WOvGh8XpEz44UYF242hR
KczfYp77OOpK8VCPXB+aT3OO4V3UzpU8XkEDf3VlPqWWBpV7kWg/8fJ6bS8d9TQ4
1pGnmabkKX+18KU+ZpJjWNyw304/a0Ba6DLS5zU8AqZXhRsL76Rc7LKhp1gfQsIH
FGmORsKO+fKmYLnwf1Oj809z5MBc28iICX2GOQa/kLFuOYdShIFJJ96E0i2xYvKF
ddE8pEMvf2SpTuvKo7MVDtgYNmifRQDb3HWk+v6FVcnNPSClkq6TIRTQM2GqFzwg
8LApAmFhgnLVZOF95c38XAI9DQNBp2G+vEJAlMvwvnkgQNcMRlcmvmmQPlfnt4Ir
/wl1DdHzBvS2iv4zATimHa0QED5e1l/rcMDmGx5ZB9KXq37+t5sgMBwTF7MZppmd
Io7OYMCeUWarXTsxNnyXhn1Nq0cAXd3qCxloqERsgYq/4RzSZXQXEeiCa8t9zqb9
FBj4F0y3p3U8z3+dhNLkNT02pkH+jdBUllVRfIeIiXdXwaVxhC0PbQcZg8eReG+M
cC0VpN6tkDOxz2Yq0I9QJIkkqLzexHYz5456X4N28iU+6uJT7qU/pJGwLyR/ak4f
a1QQeQvnmeiy/MXl37yIFCTd1kMOhVwSO0gKEHMO2/cnex4yW4WMO5VV/DF/9nFR
vJ+sVi6zPuzWsEM6eHcC5GuRYnn5hFuFLHltwLbRgwLPgcveR6/1RBXY+FJfpJhg
6Tz6LhETj5zy5wOn+PzF7CNCgX/kIt0skBHzZQxAj9zSVL7hJista7mkU7OLF8bn
IroeAE+SbkiOnBr9u52QezBQy/FsGGrkA0GJXFun7K3+rbi2WuGXNPo8Q8c7uEFe
+dQ6cw38d5ZBWRa2ClxHNCzLmwlvyFLOURHCJ7yY19i+ypgYTvAyYROBKZZw002q
Dvot+RQ+2Z8dHQPV4w/veZP0LIDvJM+Qg8KU6EFVp3mgeWCKzJKajD91WRsR5ozu
MAkraytZrm/b8+9MJtg4qySMz9NqDWJurldr+a8YIfECw9sg1hbkLcAzfu+Tpx2+
5qQaL65BNyMPRkAWsqgc4NaY8C3nTbn9cDdAIsE2Df3ZJYBOM6aH35o6d997Vlnv
SAGuF8jx6VCI+syiQLaouLI2c77CC5qHuupN0dKW9FYDYKDmaTSVWvlOHbzAqzRb
gU6uO7+gcWTXxRZ8wISqPM6khSQFNhWMM/f2ssZWwCJiEwM8wJGWkROf668Juuop
VxuZFWaXFCjWn+HSFQZABtITbuWncqS3+G4EoeMyZZXu6cahmrGakmIkvKwZM58A
ePVeS7uuNRmzlfRd75RMNenRj5C7fnLvOu+qxoo/oJBLuPsaHXWtPOQ+LopbDUmW
fI2+twnSdBs32knOlNlvxHPGKPVsYD8V5FKm3wiiPquBvxrv8i15Uj9gQ2fnWObm
uqr60xkorrTzcUgEEGTk46x7TPSNM0F1LbvW9CUKtWRZEgpGs2ZQ0bbvOop/yUgK
m3paACMl9KBOGDUkvz/mIGQkCtOLNRcDOR3PttH9fkWKu2HaSJkIQZG62y1rZ3DK
VpLMO73Xqy5PdU7tIm5uRZzvAb+ZMkCwyTnmHYcunQf+Eeqqs+bbmVJMpb8zbt+G
kYeznfcHc1SI45Rje5jAFjT3mwdSF6AVKym7eG/aFL15i9030jspfUkx3rpkjOeb
OkV3ZMG0nTCezkbImVg+2xnESYsvUyoPdUsRqOxMli1zPDef7LNfVtoWzu1tnMRJ
iW/VnAduPElKgmrHWY8YahsTGK8pw0yywuK6DPnAOcPFNRtfOvlzDsU6ygVxlfsB
4905n00soxRcKUtONPbp8VEBrmkoDtAioImXPXNrgwIEiO25V4MhNXW6Ta4AbJc/
sU770Yw1HppDFvINVktJbDbT/p0EYff9hC6y1WAUnWNcxj+SvQ0MV0K5prpoENya
mi2hXHRACZXY6UeRu2xVnfKlgyL1XDmedHrIOFuucu/7hTTC4AoSLSXmvJ4rke6c
GrIvkBUGgP9uRoZg0zhn4rtVOK/BE1SaRntNIxUfxI9q2dpFaGJEYKzuctCzLWfb
1J0Cmg86p1o2ummjEk4NOKQdxVgEoeGZh9Yd6Wb0d+r/GnvrEWPYxw0ozSp+V3gU
7oUlWmOevpO2pIa73FPE/li6PrAw9euCOxoDzhyDwOnwbmhkQ6Jq0d6RtbEvnb0U
9TuShsmPzIZ7CKtxTZ+P22IdbaiiwM2HishHtjHU22h+EZ4Fp2mhWeE3sjDTjRpb
PpP6PajHbHBoUlzFTVGGklhAxTx+REKKJ3dA1JeTi7qn1RQY236ze0mPYJb4EJD1
021C8WqFDG0xQiw1VxuB+a1cRwJG2jtNBaIpwg9O+O+A6Bsqr78tozn+J/Wt1PtV
nMWQz2EkU7Hs80I1RczeJ59COBmkonoTu+Gnsqw4HDdrkB9r4ShFLANU50IBf5Fa
/ZwtX9sfbCAXte8qlXekk8FHbN9cMwwfKgraeR84eY/qJK/J6nUCPinDl06+Pbsi
X1qCfve+JPnSUN+laGwPgB3l/PBXwjhpWY3iN3wXf/Z3J/szMADUbpCmKvnexP33
76Xt8/lubV4ni9OYn3WIIOgcrMOYQsrB+K2BMP+jxxOTYE1BzqWeEKVhmJWiYUZB
D+UluH4Ja2yfTmmZTa3FXieW6ZIFIe2VV12q8VeaJ+uB0tG4EDSBzkBNLuSKLwah
ksCt+0Qeovg6/bSJBoJ+D6DbByAbBNjy0SVcApU9KMNpLZbSzEBHPrj/IX254jNy
WVWvW+JoUmYgneA1ft2SGfj2OSI6LOigB35GkPtTF7iKZ22omACRgEjJIz4n0mxH
HpERrsyk4qvCGtHDQ/QxyF2pXxxFJqmPpSfZ8e2Q+C2Ovacc4P9LPp/e2WzmaM0G
Kr4yFntwX1YOyjUCYDR0aXCjYDGGyXfU92HmQQRyrg+/xPuAoX8Etw73JzvhQD7y
WV4gcSdk6bG3uufqbW3ZbtzoIuXplfEXluhpF2IpPblseV/xK5XrXSwQy75hewFt
Q4/+j2OZNtbz0EI5NyLt3GJOl9Vy/Oj8wApk7GYOWZIheGoAZAh1nXqxF4m5+vg5
RxrkPD+cm35DigcSbGoH9QFzKepyjRkmZxILdAKohKOPxgPyZE+6E7oWKz/Jqijv
LYJqw2InGBb0TmhhriSZP2+ETMBHnrX4lXLi+4dDhmbTBWsz2KXh8iyvZRaRcTdL
E2XcCDmiRt2n9K4maw1dcGYcbi92OMHwhLoZhPwtqv1nYIZbsVpKDdE3di3Hbxv4
qmr+CZH7YTc/Un1w4TudeFOju6IJfA7wZG8Bc33YBUE7CtGuk7BegtSBVET95T+3
UN/zEb47J5wvEeqNstb9FgCWeolmDeTTrkCs4VlgX2UISqD85PbXktMPxyYjzO8v
cgrtrVgljk0t22u+2illKdHGoNCcmfiFleGwT8vVK6RcNKOGyyl8Xph62Ty4Ntgw
0+GOg4dq6WQHTiq7q73a7AHuSZFMmcJcEuNR7IkPgdJOc9CyP0EbB97WF+Rc80Ul
3vTeoO8bB1X8GJ+xmdOqX9T2wSwP9lGNgjpd8mQqkY8vOkWwTIYD2jWSg/IRVTJV
4Yl38MxCQWB0YbEH+YD83noaoCMxWnCvK60Ihb3I3cQ6BsnwTRtUIE9WTp+WEjjF
f2rLvq3XKlfNBoXCbW4jq1lwruK6cnHAIKG8NYiG91dXB/nWUDP2XUphOUYPEtrU
8Ww2+GA3oSSbnmj2moLFv+UroobaYoE8HmHG6orfPlFZ1NHSbeWC4wPjf1IlNPG1
lNnxneZCd/U0mgpbbmKxheoNejypzQTXtlvmnRGYMZLBub8dGtig1emkw+R1pWbE
UoFxHOmnMsfsAzzr4pOVYFdVLWEwOCGcOApjk59qeCbEnkhjguyP7VK48m72VKwA
kw3nzG/fA4VMFm986YDgm+Fy4B439DYoR7n6jpnfqcnqqamftl0Z+MATu4EjW+AK
C2aUMlpCPlLvjl34LeJD2fxpTo2AYTsBSur8AkTeOT9Y33nLzX6aYDXdjekUjHzH
cyvmJDhTz5arS0BFS0NucsEiFVz2+xyEb+VQLNqJAnCmHQ1VKX2nahaRnLIKeqDw
yZUPfziuhBQ+6OmQQQawx38wj/fVyTqEyUaiui4ZTx/vDslpaPj0RXVhB3d6AesU
s3mhSYLYv4JYPKfvCTCjyiXSm28YdGhXlau/K9QBWhyE9FdsOEa6r3pVWyfcNrq5
8Yfx/jpOr2cHA8rm3yKWNI0Xz+iDXBnY/gxd1DNzPzhwXttc3rT9RUGaxLpsoHpE
lFYKZrVyzoyJvrGh/L3hWFR9zblxn3/btL6xbON2lyYqMZG/3A+//UShi4uQcgkj
zZy9cdbOjz9/04PiAh6f0FEKjKj4R+boLnMrqcVioSqyI+FkJdYtsJhCQf2RTcAS
5BYVp9Be3QWp91wPYN8/BioOd+zHeSSH3K6IUiMJX4dPv4bxRm0lT/pttNbe67XW
CBn3lRNKJu9/l1Pc3Vg0P/XqzuEYuNk/dDtDlrdvXQ/ZAr+mBz78QohKjea47FwI
SfOHkRdbLC4kJ0LZpqQI6exwdCzvzN35TKHM97W5oNj2o+NEBuYxsBga8HQ5HFFs
FZdgiefBnVHH2nggnazQJxuvKeg/bfjfuLdMb34d4R/YVrmzOGIcSgN41yGlgZ19
DxF6BWlBfVe8qHtXh72oeJ705JJ4ZtUw4ubFHXTU5D518Xuz8g44b1yCScbh8Dfj
ubhFoC6hMbOMG3Vnx4JHjnHAOO3/bjU4zwf0qc/jXqVp3lOgv+UC/mh7niV4IqsY
XeFQpRUfNm8owCzJWR9TjPiewxGcnZrpnzF3HpSrB5AFPKOQ2zHnLqBz7NgsSNf1
pBol5uG95bj2Csor2aJcFCfZt5aYQfyW6YObC3zBFmm6IcbKg7nCQXkvwZEIT6aY
Y9cMo09QyF6rAaVvLd2CN3T5kGF7A1pjm2OH0MsnydIoonlsQLrOvCSCbLG+t1Kl
52If90fNZkNFCxfRiDb61SG9+L9uIMi62b7xzpvhSpykMyE9pboPz8avJLYekubr
kNvwwvPXH7jYXYCbNfrcp9vWqx5gbA3pZz7wIfDFqpKHjqvIu6bGdmdhzuLCRbfc
L2zGgRzqpHCwsipWi22/uApy1IgjzdQJ+iHWfWoAA49uk+E2+NCm7nzOYY8k1tIG
9CqGJs3kdfYjSv5N+lfnWUdPFD+VX5vdOmcnBNwv2e/M+/1shcHjgs45D8gMkhp2
J3c/YQpT4WhTZuTIZ1KV9fVWe+oMmGkxGYzT2mj5VO3QkM06SRk6Z+WQ1m+mebPc
JWBvGRti1D7dxxusnDqN6xv3ZkrdvsNirfgtt2/eD5sSe4uIunz5Jdm6lvaBx+Mg
1p1BKX4Fbs3LXZJQ5cX/WnK10YVBixeh2VtyX7gj6qPI2Z+lBWExE6gaA0EZJB5r
BPyN48GkyDioo8sm2UQEWM9y13VQ6tC+1+qqkhSltNduDCQugdDTVnbx8rNMIaP6
A56GeYS4vwF7jWa2R68Bc6XhanaqVnWPmlW4TH9+u2tqT9jMiEQdGLFA+KEs84fO
OB7AuGIEX2tkO0zuOSr/mDlJEa7gPnYj69C1KpLkyIcRM+Bl4AoiPDVQpmVT3841
dHBau/6JV+bgii4cFmpNBjPBg4bEkk0THQfBIhKCHEfOW7zi6Cl1NXC0aSH5zrj/
+opnqMjQdv5jYkZqGPjk0pWT+lQQ/jhAUmagBtQzAAED6tXM/taLPT2Z6la3SKRF
kUIk7P/IPRDPZdLzApXttVXcTiDtGaiG8XK2ETrrvjWjjYZDhoo5+ztwvsArDBzz
JXBArNsu/lLfEKc3lq0xNHF8B5+PxfKmKqB4I9EzzTYfc26MjxvZfzVGfv0LXyFo
DmpJHtNwbxeUiQDHyTaXLMsjtz5q42V0MclsH0md8F8UEnYPBmwXZCUcbHag8edY
rBUMIj/nqyidyq6B4huOxdQgptpdygmQeSUVshSWHXPa3uIq/eZIkX2/wgVmwKo4
MCq5qxmhzYW0q9Q3oX1Sr4jbdES6qrqPqfVcy7UzowUt8PG2moNVi2r0bJV7WDOA
Sux1dutG2USo/CSQaXxfPZd60MBvhK3Czu7Fa74kSqf3WnP54NEbBhCLRTgeGCl/
7I+NiAM/brMiVavWEIZX/Dr21QrI/+Z2xkK9hOhOSf4hmOcUOQPeU3QM+df4DUN9
MuiL/maGxKHbh8WwYW6XNBF7d8ceGjXJcgXQ37gLrryOdWfmA8i94fH2r3R1aY7F
3Zcf9uDsWtFLoN5sVGN2hncjzlMUP3A25VaSvlQwnYtT9PwnCunO0PVQijSpDukW
QQSqAQLrbt3BwJplr2fjJa9UZo1P3cO4nM9pqf3f6Aq/5IznM+JDZEDUNMjp0nJL
8aDOeOEmzQ7o5Q65sPdghNHc0ClsWsfN6DHmcXTCMMAv7aOvB6exnemalU7YaRwO
yXI7MYGkOSPBdlBmmQCzZyAxHbyJds1ATNSYO21XOYox4p+RgToQ9B1KmNlsbyjj
NgaCnP6B+c4ACPBu+PtDwnHC8hXkN0BNl7fndY5ufg0/Cbss/HOmrdO7FLDSOigQ
Q4nQ5lO5hDzrwbk9NNQ5cuka1tNmaY2zmo1m7B1uLxh6UuuAcKO26Uq2TZ+kEBOl
LrIyIKLqd2vA0HXlUehXvdeWZjkJCvthZK2DivvBa1anBEvqI07B9S31xR0iUSTJ
yvh8cto1sdB5/gUScmQXhynpuZ8z03R/RChUUxYpz10KrhTMY96pgMVttgflWa3x
c6ytKjy7kSLBVRbCY1peFeBC8OHG1NLmL/o68MLbPO342WBLy9wgp368+yxR1cxK
lNXA8QRAhMA23KkyG02HV/sqLcHkD5Iz9oe1o+YApoHQXGEQYoxeBlWTOHrRCybW
gHGARrTS/+Quda8TVZryVJ32yyH8GQRTbIcQqjc4MzxmySjgEOJiFy6uhO/gC/KK
YIr58eqKTa+Vkf8m+M7KWFTtoO/PeghjdYfiRTvbm8mBExjUYP0RDI3vEdk/4S02
4ZUX+5b3RqusaeRu9ZKBSBdSH7I79+yavJBjXlC4SAMg+SmyYSuAelDAwyBGE8Y7
2DyIsDaOPU6G6yijq9zvGr6yiwKcfVYe94TRJJMMy6BO4b2wjltoD2keYTrf7686
Ev3KsERNYGWCU4O0Zam9n8ovBejhRHNau2CnN3tLqCmrn+dgwQZwSOMolUGT4Q10
HFmB+IpOPqfOx0Q/g0Ozqe7b2GCiKdUZLWjixSwE5NehU3aMBLfcru9JZdSpWlZj
RFp+zuZoKJtXCtaWpDNhB6rth2er+RKtF/QvS2cAZpxll1TrmxSw2ZYeiLPUfgCr
MVVrOr6o3kj3gnBhxlYtgyZtT9n06DWZRLfGNkpoLCcQ4JmbSwBgznK1eBZq+0Rv
nO7nuZJa6gQaginKXCXMDPFnbaGZo3lkx1ZmiWodjAcAr1zoTU/T7fC/LilPw/Sc
3RK1hKgVTM99zKasspZiZX+iHj/ZrgEZB9xzOiPKOGkQgXjWj+M995Mva+sC0My0
N4WbqonwsRR+2FXivLmM7j1aL9GiF0l2l9gR5jn/Mw+aJEASdZrKFT4uPbbi4717
fFc5R0kiSg6EKUbuSHnmmNobQGmdz81yDEPuLg8Vg5au9lwUf0L5tlTwVlZS045A
gLUi71dq2ATuqP5bEGLqOPgvj8QxPkQ7q5Vzk3dYGaSP2pn3kPfnyl3k24q99+Xr
P6GpxeUzSo8ZSuBubdqJKkF6SlBW7pJ/MU/eFWP6LIuwf2/asSfrdyBfGincQwVZ
ckLtJ2wPguJkjs8B0AfENxZlh/RCcH/Z68rNPykPqDKBAX1cRxBWWv9o9l9vwi3B
ulgM2uwtXSgOXKnjiyC6FqoWZXGFTN7eZgDr0jtAPg/Pu5KGrXkW5oW7i9kCr3HP
Wx4LJaMWuiPN8VayyDMLlVQjR+TplUZJixxMFBK3BFQCIGgU/4ieMs/xOVWFCPFI
TaC2TrMpH8hHLGovhBKfRnsHlChBK3z7jX8Eu+Eh5FWfCzZD90mYYITF+VM53qK6
gIWmMbIRnBPJYraNL4aCpTlQKLn1Uc4mBZJ0eLkbCW1lEwNDtskY5yFsTclS/ftk
EtPUbRjZMBYO1ycnmrSdJTPWcPcsyDHgT3Len9LtmXK/6a/EbaNmNb52VdeEUVmn
t8CU5aEW1yoSNcAxWAfXxkkoZYO9/1LM4VSOG2tjYZ6S3HyRFRtN8xpQXd7PDIRk
6Qz5qOme/1eva/nLJk5K0xMRPFggbfKA6Q1FyOiiY3xsgNmWcTc1k3xnKm6t3iw9
1K3LuqDoqN6xIIor2aj9rpKdOc5yj5QcDEzneysqyG9pOrr2zKwu9G1zyXmJbGBE
Jdr8XDhI+R+ez7RoolYKXVTcP1RHgcHgH2k4Cl7P7f87jFLuT6d/3R1WZ4P5fu2q
IAa/mQp1w50XjZXEHrRUXKcBuJTulbPTQzierOXyGimr+ClZAat6zHrBCYG+blM6
RJtOW+Vyi4qcmOEeH7ggkobhXoRKuuDiiB+YZ9XiEK/uG8QmC43vF7dn7kMDaqpV
a+pMnCfjOX+AUS5QJuFWrUbeWVJtqJ0ko6x3myAoldwpoEefUfd3w6soHgOMAzNW
j0iBmngmuMlR1UV/n5ZqLs019S1QCbA/JaXaLyzKRNXM8OfJrTclUa2lPHs9xYgi
BX8kuBvmfiBmGIZH9U1h3/xKhZ2gl1beFKAHdIgSXybNBWmwGlSCg8f9P5iTFSrT
nhJv8KqZoQBJByFCetBDJ5zsVW8UZe/L6CX4BVeFc9kX8py9ttRSl0eDrkjeeGUA
RDxV+ajQrXruZQN5L7rMnSJ2CIRG6KDftrJQ8ul1Bqm2pjp384TBEkKBrcNVmeDd
LJLdpNLpfJrpmCStCMDRifLcWFXfDXo/UtzjE9AVrLyY2UAWXlKF/HK1wRa+r3Eq
rWnvp+MVnnkjBGvIxOeT8SCl8eX2K3QfeSpJn+ahW6Q/aZggyQ1RgiaQgYCr9N5I
hNMTN62eFIWJ+2egbwBlJu5Zjigw4d2Yhd+4UYS9AL8nwjllJgOqLvoMSF7xUkdQ
UC8J8vVJDhB4OJEcRF2m3fwZCxTmTQCrhRVcfIy8enSYB5s27iLP5vk/JesAPlhp
/9yHcotfqyQ4ipyIu7L3tOO0FuRK2ZAo8KSAEL2YUJR2OUZcdwWsgZ3Mrc7jcTAr
QHe5PtTGV3kEzqVNhXg7Lil72ajAMPFdYExRTuGoRR96jRfhnwWbQhuWasHn4BzH
phuD7MSkbzBCv0hyk8uaPWbI1QvsiyYZ0UzrRx7utCCxiqLw4yI2cEUcq7bKp3T+
sMRjoam9IxlS2KJ6SlN678GVlQ7c5Ycp+49Wg0c5YPXaPftCW2ccevLocsAFesFY
LIT+j+MjcRQ4JpmxzmhP0NInbfKzjtdCP9OFc09eUv0X07gmh9zwJsY5w+eByttc
RSIjxWCIMBEwDQlocU0UV6IY/Mv77dHPID+H/qqvezEOu4IQrA9duXL1jBzXhSfb
08EfwdA9jASXKiY15s/I1gqWcls2TDghfZHXQaxmS70Hfkwsj+3LjImobBHfF1xH
WMRM+PF3veFL7V39fHGjygmXCU+nxjc0jBEB4f+IFbwics3tlwfJWDj+HD5LyFEE
3+luet7cnt/JjXVgI/4yJbAQXnb64TWpviUOXKjonBemJiFbU5zUiqCWywM+xWzY
bD8DdsNaKGpfBtG5htLcLFcUBJFjMq7NFo2EmTHGqLEMtTAhVYq5BvlGFZoMScnR
W8qr+XVJNTXrMau0iTh95rWe43RwmNVoUetW9SW+66jhtWtvPfGFtEq3rwKxUhJZ
dvAga0HC8tlNQQfDhaNMcZS7zqSgMFuFHjZyd37T5GrK9lz98enMCTZYGT5ZM4bH
hzG5pIkyXRGAPE6tu4hbuiboA8fvllBkbpaZv+BRaFGJWaGnZNjwU4fafp7mYmvn
FJS+lISDFlQy2HzrmQIn+58s93g6uEfL5Bd4B/+JvVgbSboJn4yaTq5czB8AzRWS
h7SC4a7e1fr1uoGXNwMdJzZ3Yd4Q4RHNeTZ2wzoZ5T60wHmAW4Vf2xmuNXZZrm0R
VFt/YZDMwr5HKh7TOpypaaAjFBC7kLNQkUpRs+znxEkkEXZ8lOQQ7tPu6P7NT+8p
9Bv+UjKei+i8qOpY8tjwXamcmAVNj1ps46Ot0eQvDrcrRq+o1ZXvT6DFSrwOdReI
Mr1XX/qcXqw4N2lrPbsuMmszylWaf46aeJlIFvmyGgae+Pgsjsd7M7dMDID7d1n6
2MCcr1AaVMhwqELj4JZAfY0nfsJD5K7sr3dC03No32mMdAi3HujHycITiTnFSgBJ
jOaSXcjeDBbphk967wKl+9vYaQHNuIA9PILx3HzjlynWZFchJg8CFomVllvbYZGS
dAdu+AyY2itZiUJQHjm085jdDOBuWArxno4uSTr1c11arzJkqUDnt3HRCJUeXaPa
vLR7EtIliqSafz2VflDMd/S0t2hM8EkNBLQwG5B6FK6Ep1WAyyizUoow4qiKhOL8
BbB+v1MvTncMSIWOhcWmiKb4Rm9rO94X7B0XdCxop5eUmu9eW5Q/z+2f22MSJWRR
n9zityOvk/ngdiLT3dFqxowuZjVsx1ICgoCrDM8Gp5PA/jlJjWilhTSlEidKOrjN
AwZMu50rxlHN2sORAYjgSd4WDJkynpA8YijdAL3mvjxEPi7Ie0Or+cPhAnpANdGS
uIeQHpd4K9bfdKnbdBGFgMLn0/T2yroSOulcGIS45jsrU7gEIf+gQlCxiXvHU9jZ
6wOxDPMtqE3tYUgV2s4p8ursujhUKTEq3XdmnBpjhYV61YsF1GSkWR+o8HjragfP
GV3Kg80uwh0NMaM0NFnpF2Px851sxuByEVYZaI9OxxWC/BVbkYLTuaQP42nuEpd7
x/5utar1pGRH6OTh3ACsW54k5H9u5iD1gDOn8NJIMViHOThP61JZmE1WGS7RcLFM
l9XXaxi+DCUvdv+dgOIRFT5wtJ6TUyl3wMKmoK7ghH9jAn1i6Wz+ziXdCdBN4UZm
33zalCGovD35WIwAIvtCMPH99L0tGUAbTq/rR/bedD9nr+t6rb5zm4BkzDc4nj8D
KmAzgrIXR3kklAjPe1Q01YixfYSCm2FdvcBFPhZEVgjLMdp8vnqedWog3AoyqHsv
i6eIE9uHTwTEVBy5H0fC7tUfMqX5zU+wVvHdqMb9XOCjuE4gvG6oL7w5cb8VwAIF
Kwk3fFeHehbMpL/Vb9ecCKVcgk2yCgFbhPgwF4Nctt09Qf7vxZAAxk2qhVeCycSM
f1GYj5ibAxD/dstC6PUwh5cjgqtSIWlxV4BZxfL2DKzriG9cftk/CDufbFmlzK+Y
0xWCcg4Wn3pAtCnlSXhpkwWMGfwgh0TJ3ybOVp4Pmf8t0Tkc2reIQDQoY/HdbhUF
fvJooBZRMFTIjXOGjzRANsjWwskeoIqj4HE24mhPyuZFF4k7DwlCha0QyNagM8OR
mbpCN5AKzA8m4JXmhLxL5oQcabXnd2onBVcD4zUORTlPIP5Z7/McLNLYj164aicI
1Hh1R6wF9dGaBfQpMKWGGPlFSaUEVHZbtt9j3PtpaybcxU/JiBFQVOoiZb1A0eY4
ooxn7JxpAyI8me/aBH9aabb64kGnKATRqINcNh8opS3lwniszQKuO5rYatM8DoX9
afstZPK9MLwiC5MHfNqdCRAzJ3685TGJz7LyV74C+w7T8i596hzHZ8hCb0YruDZG
u83U6zKLn89s0bknNoe5CAYJjtS1Bwf23CwHRexwUC5YPCR6HEJ5vKFOIA5ZhmPF
cwfsY5h/DNJRBd2zs2KUJWA6upAFTnmrc9il2qrTqQdCSr7beBredMxx8sMPZ5wH
iRi5aWYeJCWr/62XjlgpKUK84u/gT1jvAXHuxgA0fFs3Ia7yJxn/qqE3oD9NzxYp
K97KziuX5at91cm6aQoEtNfxQGMFhrNY+KRUDRjWzFdq3eHZ/4odLLw0ou7REnK4
GB5hTlEkpTWKGbNZiR43hwLVw7lQAh/Wr2aUKwRne/CPmkR9NjmwHzKzFRb4vwQK
hWwy0SOjxCCrmoADBbRQmn8trBF5v1J8uD8aWcBGv/EyhQiSgXhKYls44xeLMN5z
UTMHtMQMz0jSgDUcKBShwP4cY9nTbCNJGJsCO7724Mjwx1oPUDke7fDj+yaOPT67
VJqAKL3mxD72vcPZ/+FBy/+Fswnx7PDJpShKQtuRRHKuY0V6fQViJ1JiWQ1kQtV9
Xgs7PcPXkh3TLuyKT/6Ldj/ZzFBxyKTpmZKvPubSTWD99HeNNqCqdu6TZ4jH9phZ
r6GPsdhCm+SjgxXqgbzXmJSis9b93wRYQ4lHV0XlyW+V2POE3FbkkbgEr3ToGObr
Kcphxz7Ey28yck7e5g7xV95foraRIeADTlsMDl102LetybfSSrg5x4G2OlOscVof
8576/PqBeOEqyZKFRHkEsRXcWoPrycpboiHvbbl77SFPdp2uODnnJ10X+e4eVyXs
9dPSGCB5tBMJnI3cQ1ZZKSJk5jwYX/qAr4ei7D/XaZc3fdwLRmwAmF1i620f6lZM
a7wxIoQZ4aHHKuj3KuH/6uT2M4Fw4jV7GuRSagp0n1iA2e9+Km4HXdX5YjLj74kU
+rvCB+yM9sEGFOHhvkMJXazIqFS8/Wgu15pQDs1Uq4mq8PLlB9lTkhS7j26SaCtL
U3lydirCM8duiR9Zm+6/HZQXBUQZ4p3ZqyotVjoAf0i0MBVrJENeBtIrD1kBgRSM
eAbk2TcAmRod0TvsF4fQHY0XLdyCy+5aCN8Q4i0O968MQQ55Zm3LOPtOZTCs/K6n
NO2dhDKWON3eABLSFD45RAXmAZ00FVJstt+YfIXY9ozLMSG8ihmrieghgvhwnvq2
CdsBTS8jdrfryp+4qcXgXiBpq172yCVpQaTPuHEQl1q+Qjk0kwjgdFX0/aie1p8T
ByZQI6roT30ezZREVfskqsM4hnrC5rrkTlDPi96PmC43KQ3y3iR8f9FeDjTfOrSC
t5ck+zlCE0tK2Boqjlk/1SPcGmwzMy1MWSuroemBHTvSKMh6Yhm+6umKlkQ8V0ei
BDkMTHNW48AcfWb4reySbdQDxftyUSPb+1oYr2ZhajoVZsVW8P8aLg9dlbNqlkvZ
5wuNecELdqTQudGX5b+rjNurLkBT/9eBM1Wl+ZXtZ1McMUT0vv/CwZws7+hqIoKa
OumXYewCfBHM9R6pHyHO9hntiO8iUziUMWIltf4EJCHmt7Ro8X72O1nda7jg28ey
UR8H5a/lM5D2825WknPNqJKoDkix/StVpfWGX1ORjQ2heu3y1GzqJZAuA1jzAZvt
trqc5iOzrbBtrrWr8/B+hGKax73ll7KXmFhQG17NPR8SBKIgazXnh7nXeNqVZbWk
Wyx9Na7v7W96mWn68klrFYIH+6/fjUaIzwM/W9ud0g3yo2KN1MEk7D1XESRQKZAq
NFwf2IyF/Be+sEvA1fJ+vtTuNg4QxlYBccN18AOEdd00gS9wCS4Gd7Kd+7kciJSH
JXHopvg1OMfHxvtCud6c4qRL3cyp2TmtGlzYIUJjjSmZ99EucAmrXritbsIe9MO4
S6hsyOUX8Ymx55O+KAvcsE/8mrwFnUIoLPPxazpu/wyhE7MjJV1beCE6JvCG8LPM
bg+BnPWzaefo6za6Z1qnSSlVIZIYJ0jQJ3MWsBpXpN2v2BsINMvOeQkXFXIAUHs8
BXjfffBYzG02njrstlfyoY3Vh0r+XtnfXLM3aAzn710YNqHj+sKTCXR3la8tLMij
YAGBUjYynMe5aAsaGqQxBJ1Gx/u7+eoaZYUfq4HHLkwtIZu8IdxnA22w/oi2ChlM
XzEl6b5n2QfDul32SRHp+ID49TbkJiEj3IumVg7C2atIQjDOFZ9Vku1N+SRXdPTE
bGtMkACQaNI0Hv1B0/AJ7ljMGn2eRrn8UQNUSWkT7Uj5bG1HRk4KhiFGQbx91jVo
/z2uZFp3cb1W/q1UZuEexAaiaxKMLA7LG1qBdyMjH0ECclZeWLroD8lHH5nG0mBV
QiVek0gUS3xtdXysD7To0YpbsotfzakTSKZSc+PLAUNcVtkx4iDth/i1WbAlvxnW
oeGad3iDB2ZVyEc2b/AReUzc/pfQOk6wrBPElB5G3bCTnONwILcyZkQpj3KZQhXd
EQaZ7TQeZsLHZ+LfJ0ycXlktP3r373EkVyU6vep0wamkIjNvaZD4FXQ8LVRjs1GC
ubV3PoZGCu4OOgJ67GlbMeZYPS5Zfx07a9VMeMu5/2AqH/eKKCM9q9zrzUaMbezU
7KHeNt9qsRGZLOVgRbn8s/gWTR/Dl7l4ppWoBwKroWYeLaygm0gZjA5mEt41xJj/
9vSHqCKb37jX47cai0oBWgfnSsG5fj8w1Z5z90pE6cZuJby9W8+KpjfRXubgjm5K
0d096pJqL5y/d5xzmXk56BPSk52oP21bbbv/CU9HLJjYeD9sBvlFWHX6dJSzLSyx
ClGOJDIs/4WdL93+tiypUdJ+S0k/PLg6/UI9GMfrxGuj+7FKESjRunxlK8ZL8pPs
sbEcZwZfjaWit2tu78BPBaCau26SaMV0TGXy1uUUT7HzW7TIGMa79UcDt+slBdTi
V0OY9nxhWI0k9y+jdFXJuutVjfFM54jPXUnwAYW3nlm4fXJ3ovc/0eImde2Y7TfB
LesjJzKvY+ArguPZvCiFTHVF5UUZg9dfYX9oIGF6AbN1fXZqTqU+s5XO+TWc5Dh2
vLcx7P125QHl6+LfkItwOUyqKvlRFRYaL9o/I1DFNwTxyCKsecx+fWGUmj1sAS0n
RAB5htiapRsVNjGpdyKosSqTjrW8e2vWk6ADd2avOq5XKdG866s2BEQkT8mWyRns
0ATU7uZKUJX2PPEOJraJuUgi4ZKcIx9QggjNoNpuMuMStbV6Z/nnEIiuSenx7TFX
+8N6+B15yfcskDEc9h65nIybO5LnV4e2FqsGWC7vASTwx/OQ/u5WLK/LCzWn4x27
vdURVF0h58aQVEh9BjTQJoldCzfLe1+wsKALx1X48cor769QqJ+FdBYV503CxgFu
aMyvHrVcCR2aj0WqqFcQuqrVp+rUR6qOebyw2nc+0hoe6+2GkaJYwr9BTcHcay1r
Ff3pzy9NiMg2njGNUEULzvCuS291nfM5CnH25kxgD7dZ4WiZYCxheKu4NAx0447H
IRGKJ3h5YBzoKIp1F42QYq+HD6D7sXyUEks0YoDxURxL0OLkI0ld80i6fnOnu/qb
t5zpaKIuEzIBX+B8a4z10sLwnFEEsHbo9B5uVlR0DzqWnW/FldaEUpvDFIzQm577
C8LHfmVBDi/gsuLg4vaiODPnq478S7ujJhR3LgqeeYESc7vOxYB6ZMZGDoRI9pHw
uPHbOudb4TpDc++u6TJWjpqPLAvRXYEK9H4JGRla2SQnApxm6qR1B3vk53Ssr+Jc
nzyi7/dPIDs8ym+NpxzLeoeAuE5RYmZfIBTajBBorvkaeT9WkEJh2/E2rrydjoYU
eoLcZqEpvZTI8NVtq7/b4wkCtmW6O7JnAZZoeM/tNuHsSN04j3uAvY0vqX3wEry0
YCkAXx8lGtK4n2hERXh/UbpLyx9v8zes8ahsE7FTBAUrcY6Hm3kN//PWnkcptBsH
aiMLrjHJSBSsVn5gnfOne5SSi3XPie1YxwRv8uZCgUT3FcPXas1eNIHanaJHcxNa
5gIRpDTX/uAQ6m1ag1MpKdJSVeEc2AL/qvLGpGWLYaWtpL0Xt95KWIyitEc4ggDf
aFu+9lSPIhjugjdmKq9xr+GRfIQIz4a+t6Keht2tzkVQF5VBOZRyp0Z05HjprKzl
mkTAf1GbQ+C6NlMB8SvNJz/LYFoGaDTT8Wle02VStA6enT2PN+fvAoX8cOWMofgL
cyuENDaMjKdoH9m3AgictvPq8J3qAe1EvWbobR1V7C9WpMfY/VVIpN67ekaZbbfP
gtDJVQ/KvINQjHJHezingoVkcSevvnzNAfTFoXL/YiPnsf8ldwbmv973akiM0vox
/GDDmk0Q3x1S7rrPdzONwk6EU4/3ox3h8igPpaRf4kOe+gbBMjUvhr6u32VK3FT8
MP+Uu61A/28siRDS64nDDH7EwoITaZzh3X55Z/DSOrSnCMKMCPYIgewQkBUT70/f
na0JTV1930LuT8H/As2ngJHEZLnjeNuqlt99YGkcKTMwjfNr8tN8pxnHePd1NiLK
bJD9l5JNKmIaTYzzq6+crGC/MDcjJJ/XsoOshak3KKDWc5silBybVetgYZgCPN6S
ZdIxcqZ0c11YyEFCmxqfJY6gwA7xmWiAooV3kOLr/U93Gy9/MD3XqTcy7Vt9Jdms
qWclDf3x2yzWenE/XdJQRxAYz0XcWAuedqdZNIztaXmOiNSqUwZwqsNx6FWXuC+K
zceSVzJJ/VmqaYC1a9KvgTtbjSXWZ8qonPj64Mfp+udo6dyhHliHKp953e19GUxi
KRajzVvSRhvJvDWYI833Tk8yvaPdNU6jrq2DkY9qpO+3kxXNAkZwCRMgqysTdjmF
R3m7w2bRY8FG/GKVAuAcX6eq8RTIcLMMOEt5fae01l51aFJlVtbcmLlh1ObD9XAO
Lzi4OB9fV1OSs0nKKFSzizuMKe5gZd85mRzG6o0R+NdrV1jrsGupDoPJbtJu89aj
eXmklqpBzDomDIrnvRJCt+awL04DA6wQOKNtUzs7IOsqj18CaFY9RVF3wezdVwzw
bU73+9jdb5wgerO9ZwY9iKbj7c9WSE400YwhH+OHB1yu628QWlsm+6EPsrbd45BD
nyeU2Bhv7NEoO3vipQaJUS7YMWDPNJsPbByJm9xRRM4Gfdd5JhAiTaNSOQ9pDgXE
Vp+VNHRTU/fkqRozG3FyDalvEtPShZ4FzGXEThKBGrQV2ia/edbQwvUwS+/n/xtU
L3baXuy9C9t9uVHABz0TUy1YvgFP7104cGnPzoql7h+A/PjfDT6zcToJ6LzxaDQV
R+ElvpU90aYaSQfxxM0wwRlTD8sSSbbSunfvBXUTjZUZtnjHjay8YnvebmotbZry
4J+sp6CX/3vGnbm+bS4BO7HCD239lgo6RWTibhwOJ7kXf8riYACNdLTB4agFRF0u
jaAz65cgADKDxgMnyHVEJCZ6ssaLG6SGqtpkiXZNUON/2iWuyWS/c7FW6ZYEd9yF
8aCCCOUCnKA98zZyv44Mhe84NCCupCB5poEd49ons0qGBQjNPvzK4CAYN831mMhr
l5uM8iMKSBCHdzTzi0gKcDveEoVLBXgNLDDrxIRpmDNctX/K3EdLkvAKIkxfIA9G
4/kPJJAGYJvAq0Abk9/0RYlQWVAorkmChdRFcKHqu+WhH9bqgFRz4d7dFJ0olnA/
VaDgPKRPms/rCQw/dFcLCMGyYBq9j57Hb/7liqeBHDEms5aTXQQKcsT3iJJWxROc
NFxlVA1z095c7Vp4tW3vjU1gYv6EYXqfVFaWSJtm/6QRMunWKDl70nxQJkaP1SHt
JMFwSTWyoQdPDdLhMfKl85EB3t8EQDNYVq3lYWa76XIKBtUbEyzVNCGWbBC4qLeR
llDEk2xwI30u3Sz9sDXZkaMeQ7dwfzkQe/O0yqsXo0R0geeNiNMLhk/aBq8+55Vs
raJq/ZHGqpWrIxr3hlrjAdPCzUrOznJiJHxnM1T/TCWcCt/22BKu92FyyMX785QF
tNmo8ozB2ulcLpjA4jZgAhgIoPawibgEOjSuU1m3MewIIsla4e6tT5IJ5GPse8PX
Afud8UiHquldeA+sqJnvanLeBCcdE4h2Tm9mhOxgmNKUMx7AuVxvRGP/Mp8D/fWH
q3fEj4Sog+T8/nn0auZlCCTvs0IQTmM/JYboOK72UpjEGGQXDBDUvT0617KX1OGP
2u994vYCodeyAXsR3YPn2wiGX5DVX7bAjBCwtobWSwtkohdOSWUKDReJ9+g7+onQ
RqVD2ct6yMCFYdkKFp9FoF5cGFbRSYC8ejJLRhtEhBa1gVEYL07hV4yGdFrVuh5K
Iqq6xT+jIFS3c+LVYmTpHwBqeCSNfu9i2NL+gs5u+aqBSi5Yoy1RuXhblzkt1w7v
SfqEwn8VUcOqEXYVBFuKqIUezFBKHebxzCNrkp66Q+0Q3xdBoY8NaBT8ggCzs1S/
F6rPFp+1QFGYzS+UHlIkr72w1EEOLKbaD/Hm8hfadLBvyigZSdlji8jNG8F9gzsf
wkUKh5LZDMFpaC7hjsYdTjGDQd4mGSrELTsrDR7mz2aojBgZv5MaS67UfhRemSf1
3o0A9eDNwmPia13g1DgDsrpb4U45FLpJQO88UUq+Puzth8t5xNuWQ0sWNKh2hHdq
JgSCYWsu0R6oVhj1ObTR5p7MbJD6mZPRk4NsJw7FhcRT0zjc8GmD0/SkNm3TbRft
+T9Lg9XYpeQAawsdaQdI+sBURp20QrubT+AtzuFeLHqbYsL06zJcQiol4Ixi19Ss
jzOc7MHeoOCE+zUNLae4F7l29qGcfZQ2KL0l9xMWGyx+Hv2UjvWTepA0F4u274gQ
Yt5sWJWP7UG3p3c9dub/sJGmix4GYvIzePlFMiopsEUvYxzYMNDBqHa26bZQCBy6
+4QRQcyZN0/n4497+cqpccYnc2YSIDmcQR/fM2ufPR2SKohJJv7PE5f/2GbuUf23
zhT26W6BeXK0obSDNh6jk7e/7SJEVEiZVEewmP3K2bMX0mu/m5BBYr5n5e0bugBC
xp/dPU99KrQe3wMLIzB5rGcD+tmNPOKbwJSbZuf6bnxVEifbw9Xbi55DOMwBZpEa
jlr9/LXO+BSdoQELDELLyd2T4h7jAQPWNcXpN1VM0EQU1aJ4hWstyOTXwBPncmOX
otRGfWue8kT6AT0e3Qu5Xu/FXn7iaUxRrUIWn8Wxh1xFfuEYkwGBZMNpPOtdGOR4
pkK/570I357I9mzx0xjXWTofI/1V2mQgLIzjGPU+JqXrvL9MuiU+9RV056N3dmJ7
+W71l4UQIOPcxxzEJVv/fSy4DxaMfAsr/t7dquXrZS3CiL0Nz5jO0qDZPmz3SAcP
8gt9d3zGlHHzfQl5+otLR45islaYc4c9H+CBFA4OgoeVcCYzDU8LKrPWcxHFboI6
XG8XWLpluQUI3fC7mXPDiFz/4GW19CwNjXkTyD6JAPckk2ckKksL/maIpbeeXIgo
AWxDGC1s7TVsvMxIHn42h8iTLHdLGkzpFBVOhqkffiN0KjSmJ8Fn2tpG6SlS+6tB
6vo+xI4EHRSPhwG0c3XRxNEsMk9obmHEIVt3nKzRnIHgV2zDzRFJjoi9JnQJHhC3
isDj5ae49Xmg/962dGZkc69PTS3YTTNS5TodlNdXu9uiRqJM2TjiER2FeZmRUVSS
Zxy8gqGLmP6P7guOD7vZno1IPcfuZZ/antvWqkFPiJxmu8zFSYvj5hESsVXwY1VM
ovTTBFwFeNooEIWwJW/RTWlNKQpqr/Miw2/1npOeLiVdSbSY0iMOunCkSIJjL/Nk
iYymKb1WPlLeGtD1LEY+T4YHZgEmkxOf4BoRtKIqT37OP7bnutKuMSqu7hSolH4p
WUjJujL+l8/48aXz8o0ajIkDNyDgQ/sDPllw/QPA4VW3KRvkkSS6ynNZCVtn3SyQ
JGbDITn6CMPXLPthbG4KOxF1CwqTl+0uLRJrqtw9RTaBV1mUPK4/48QB4bWdsOSj
i7e1M6wl+8/cMKd7K3NfbZxsxHh/mHmWUdicnBT2JQ9+vItaj3eQZIo2czwA/NoY
BwJWfm2Jnc8gNT0hCO3J2Tac2Yz/t0lhoPyni41ZuXV+LuwsDDVa9tnrchjjG0OW
N+9C2zDDn4+AKdk3eb0qyXSNbBFAddVF8GUh/lCm0WdY7E67QKGPToSKkL8oE5jU
hEPr5ye15EpJK0RnKBFAKz+LLXCmRbuuNPMqAu7+dX4VBV0HvKDSTi/mgNkXRVRP
QzKH9IdjjsxCz/ENTxgUZgJB5OBfm1/hSQNJ/tI0xudMNByBGXBNTAUzFZVi+NE3
SH4upcQsOp6HH1JspUBRHNq5s9637Qirx7a6CQMX2lw8/eiOvmswGeXf5daVCXrg
xJDVxmQ97DYBw05s81INgCaJ5NLGQA7BaOwPHHO8MvPQcYuRbmdSHtqxpPmXbqFp
SOjsYjws8r+f155X3aOrU31rJ+yazSwrghhbJPaIaict9p5YHo/G3h4EdgHvD0IF
Mo3a3EnYrdRe9F2BtmVbOBi+Ck5Kyj/TrIPn6qtXf6lC74BkhiAj7J5LAVsgTft/
FIEC7xir6+N0fPZdudRk920VThZhD+4xOjwqYTXTziACKreYUTn7QQXPavFQVP8r
cZoxNycqC3bFyiLFmTU7ZV9Kyn0eZMMktF31pqrBHbfX0SQVeWtl8cNaHMm4oVFs
iuALNErQMdXlslGx2WuGjD+YOZVzoykXWcEa286U/BlE2nfzUaLomsv7yCoJ+ZNN
PQNwXk4A8mJ/tWgPW1gmr3YxwSe+GJgABRSmms3hV3KPWOmhfH6sYYl9dqF5StY6
w6vczdF0BPWlkig+qG9EwUL7krZ5JTHIK358/X/EH0zPjXdIwRUSvMb9aX8CFxML
UCVAakKpE9JzGy/5onKoxiKlWGpb4gdHNFYDD9rHS/mGqiykLfT20vFTuaBwO8/7
c6wZKJZlj+jellYCD3xnKFpYvaXJxWJmKszvpf8T94Z/oxe7n38P7Hg4u5T6HhvG
5UMzpUGe5373zF0JVRpYhUCMRUK61sufx1G/lCDAhilGgoAqpUZnN1zaHExFXRct
sAMa3ueXPC5yL41lMgUvjmjj+hWhfwJPKAakzG8/Ln4wJbP3aY2rAdmSCBJRR8wk
Aw3Qwrt48jr3jUqdSfU8QaTHy0zsWtEW+g8Y5F9Bkt9qUgUXhSXCsZfxqt8TaJYo
bl05mJhpYazoQjJGcyN3rQmlNVrV3lEotLQp6q6SeM0S/dQ+lizHghMkXBd29pSL
l38S3QYBRW6UjvyZLhuFgKUEqAm7wjP4NypPYgx1pRYw9RBSCHE1LLKWl2c2QAjk
WOy9P7QIfaf5X4n1RtmcM3o11euxrBPOUj35SxedWrYISHSo3DRmRD8RI+Kuutaf
h+Ru9rtpa3Sdg4gZ0wh+1DnGRPhsh3SlB04G9M6Dna9cf36IrRkxAG2qv4P7Oa4D
sInUkO+G1kAHO618yWwI+UWa/oWNxml87oiIsOS6bUzgzQ31r3SYrL3oOQUZFv/b
9tdE16zxJYDRyrOLkt2cLsyS6sxKL+VvRJ4a2IDIgXwvxaOTMk7A8OkBHFE7kPWh
MbboilKiETiJaX7PK5gknFMip4AHntGAT0e4/dCpSjy392XIztYt1uPhweOWNQ7r
IZAdB0t98Y8/iK+OXNq2nDe2ccNjWVqsV8teo4Q5x2MK8R6p8J4/4fp8qg//JTyi
cbOJi7hDddOlL4GVzi6sdy6eaIU1lMZbKvdRd2PgeriehQOKXIol+a8k2yBYeS43
ZG8WOcb3edmjHtGHmUvLa5SWXnpfFbE3zzbllZasaUqbQvT3kbx6rYsDv2hXU/51
AcIyHXObo6Vo+muNcb0UKAZmX9t0BBV31qPvm7zk1HF5FZYLJ5j39tAB4HO3UNk/
DiJ6h1uLuTBiiH+BCdsiXjiFtGUsITq+eVv7Y80pPAzMV9M5AW0Tpq8+ZuwGh4VS
CVJaUFcAFNTGOzLEiTlfvaqZOQ5ePdCnBDVpoCJKqGP/ajDn3pXqPeo/CUwUF4bO
TP01j11zJgWxrqgtNHq/I2u0jxfSOQU5q/+JixC5goqx1VaEa8WHKzUJNY1TlNpg
Iz6KlzVrfAbs+F7AHcwHNNrLwZmB/emSuzTMXVjRdUdYZNZGkvHtkF8gAhjatMJr
I5pA5R3ZliUlRAumOXX+qBg7h2xXfOF/5Xo8KnkJrmk4rddTA9pqtS3YxPwSjFum
SwCACILcvl0vGAzMT+ZMSRqnUeGTK38BqYN62ZwpGEgqGFRwbGB0xmFCd2+25ZQ8
OtJcl4u7XNyPNFfPzKDH11O3xvMIPGF+R18qA6I824/6KZ9d32oyNkNF2lxss4NO
QSDJyUELNmhxtLcXB9TIwx4XhpxFxuCVQ5vAxBGbckE2PVP7LwM7UlsUgfm8U5Eb
8v5PCFF/cGSU6zB7JtW0B80Karej1Tc69CfPnOuiyP3m4bbNrkZ6ljsprNEAwFnw
pRzW0RZv/SrDTJR5QhWsnDIJ77iBXWg1rUkLbHgfXsjo/YUlqtLOk1PUzbT6Z2nD
ZsdYAJ0S4hqGlIorb4qqEQuXckcj+xluGY7K+KW7mVaXj/1BR618KkIkG59QlJ+Y
+/YTZP1OXOsu2zKBqA/HwG9U8/GNQhma2iAELGLHzm8DVXWnPI2kQtatKOCqmY6/
B1Ul/qHfxgY1Gj4DZCqsC8K17qZ+zNLLWnJjHHEGtAehZhdC1T1uwD0XuQB3BDxL
a3yxDoMa3KgAQn5NCeOGNSRRZ39tfLSTxzIEX/TdPSg1DFg3MvmxK+/XPiQL1cMU
YVqkmZ1B//tBMx2KVkroC65o/gyXFh7r69UidIahYdLW4it8ZBtbMpW3CIa+ax9H
dxzDij+gtqNfJDyVXXn4VgbYX5uF8nZxO5wIdnU5N4yyc1qEcvk6XiO4HgyldsMU
LmhzIX4LuIBbopXXs099jOJJFqQjZqbZn13VOIH7vlE8vjYnoNNmDyqfvYTRmFik
16z11P1ILE/TAcL4kjrQhtcLUS9khG8/ZZckINQmMbs1t3u8Ofj7eIhmv3d/SN+E
brbO08Pu/3LKzPcxzuBDEkPQSY+Cw02m9XB+spRtEMgHZBtamQvqfp8teSObbrmX
3AhGWr0OCe3FyBCpCIm4lmqQUa7t55lX9wlqAX+pr1JseQgjlAeXRU2DlUq595W6
0O/kvS1iJb3fG+urh5KfZwQBflfqGO0Gi0e6Qk3tH+EP/2rKZyOoJ1QhY1r+1bSf
OBybyUAEmbo036qywtRYSmBLahVWMDBLdn0rRSzrXdyu8nZQ16mk/uUXxjDVrCoS
TPi5/IAQWU9UDJTNQZeg2zorBTWjqlteayjz2PX+AAwQVvKHq132/ztDazuuf1zA
3uyhmFGLwFHPVrzDW03zndACrPBpBJ1Nlpzt47Fm9diTdzfFrR9jxYfpdZZ9bce8
pyUuD7mmb6yd9QTSn4m1MtUQ35nAteCWV/6QMeCjCMRcppx9Xr4c7Av93K9YuNbP
3J3hthbXnpVZaTewuOI/NaS0KyxsuzfLr7TWiNvxU03ruFYc2jcQg3RKwLqa1OsN
55l8LWwe42MUU8r50snhGWE9tNL6gyJemOgFyPFBJtR3oWPcxGfErsdxq2qAqajR
96yyX7Rkclzjp7k/IyTeP0UEsDbrZFYwKMzdNWnujI+BdY7FXNUzPJdCxxubPJWM
G57kPLZ+bo7RcLwtz0K40rtrGtkqW7PZJAUGvlqOMX30OJu03R+h9CTfDLqDOuqz
RblfzZAC6dF6CXUJQF5u3hiRw7jgwTftpSCBmxpnXPN4lzz578A7NtxbQ7shkAz2
850XCUxfbRBSMr6UadDOhGTxrzgUGRuf0On9zKbgHts1sAEKaft510LLtFwF0Xfd
NIydB4DsKCdnPBx6GzRFJIWTCa43uKjfh6nogFs+mAPCPlIJI5JfC2aMxVY8q/ko
ZrGcjtoMza5dtWVjshHpO0lnnFMY8VDp7gijts8hnGXuctjhVWZ6suyk/rTBRwmm
s22FhF8tRuEAPfIWnTDpDQ6YHLFj3KiWrEYHsYmj7AlYxoK4uveT5ohMw5nwVGiy
siginfYhAurxae8FpjzNljyPN2TP6WKYy3q1v0qebuyFOR266OyrxUjsni9QXc90
qi2CUuQkIzs74Uoz7kHFRb0z55i8V9ZfhGJ6E4suA/JMYnto7xGTHXMrnu5HZZLD
naZdlEH96gltEVXT9g3jw/QMuABvZpW0u++XiPW+kBUgdun/sWtt7z0etes5gghC
PUDxFxRU+uuXp9JtQWdHDDkYII7Xkjd2A3EiOW0stH44zlF3ibO0QgKzn7jFReFv
TApIwdvwhDyxvsxfmdoCOoFVBQ1qhwMWcFmwswlmW2eeiiwsR/hz5HycBYHEWsU+
P4TNdEOLswXoLC6k3y0rJsuUmIp7mnD8D0XnIhxp9I/c2PvKvvqkP9ecoVBqu6j8
niCzZ/BXQowSlHDkwO9g1C8auK24GTbv52yguNu+1GAmAu/VhFI61yedZh8DKusq
4XRIFQv6IJAm3NksQXZbu+FrLmGBpKdooV5rLH3sd7euyD4ph51Mwg7n/lciuQJ+
/GxUhZeL0rrlQZQG2rERXxxm1yaKA/DxWqdt5i+VOSj9i3rnSK52qEXWCaoYFd9r
ofPvcMrsxTKvyfYvocTsgU57UR3jv+Jj3fMv4P94FOKoSoiZP56suef53dN3RMIM
1a2pXig5WW+Xdqiw06YCGQOtSlL+K4gANYvy1S2sXEtRa7F/R9FIt0YymrqFitk0
U81ws0rURH4iRh++nNLGdnl9bWWGQZg2ZK5uUKg/4LxxQbg9q45SNebTLEX9Mysk
oo/DIs5WZLtxJ8EAZZn88vpAkNXJSdMbZi4GAdmEBbNjwBB49P3oheTtr3uBuaHb
YOajEwaubCiSg5OuqPBoqwIq+UHHOWUZoN4PHhnkyQQFvZvwkD74oXWw14S2Qv9+
xVDXB9xQPuOXMlfndwfWZ+b+laWsN0he3U7SZhm3HFuKx8RuhI6DyomiPWGDmqzc
HAPnL7LHA3w4GaHBvymrhiKqe0nRHT2JrsYoIJha39INGpjpvuAXxPJMIW6vjIE4
aI1CcxDxsDSDzpXVYJPXv+ajjVSsdFBWxMOxCOmPxt7jaa+PjUTcMccBAlpkSjCg
7/irvAGpzJr4BwtZ0uxd48LZINme1fZ3l/03qskOszybL556KXmkPgzRhEBvoLYD
M8aUEtbrAjv6Xw7XGgoDX9481iaxk9/mqrrNIIBnbnsAbb0MGgnu8hNt79xajaTf
e8uvEFvf/JutEnOvYBIVoLlzfTLTdbssxKHxOecxp67n4hPggsuiYTwcqzz557D1
K2hEUXjaU7qxDVb4scPjy75lwRFAygynQEqxz2kt1i0695F7hPfumKXBnq5rry0O
TD50Cy++RU3gZsCcOQwZ3w4PrzTG9uUw/2kajKnxmC+WnAobvPNJ9tAL5tYs8Gck
+fdyEIBVmGxJpJl4R0Fe/yKrsxfm7KPL092Q3/+mpJgASKmayLFdmj+jSPQl4aKX
UW4FHsA4fUH7Kkybihd+pffvOs6Mo4aVi83+eo2XdB7mo1BvVo9N2GZm+DUutx/r
W356wZvK5so6LlwdJPEMxnYSKML+H90tKw6AaouMIoqoJoVTCz0cbsqPk1lykOhd
McymAB+4shPCD6bIKrcWoXIwpYzDQ+1W3fMViQS4Qi5DI191mfMVxOU+KE3KCLsZ
/f8k9f4m/4yGh11mX0XuQFwJ80me1JWknzsqzv7j7wvb3E0VbSj0B6gMzKpTlgAc
0Isn8M9nW8Fw4XrNUgNYdXxFVQBhK54UOaXZ3YErcXTDDEHoeVC206wZh3sP3vzf
qXIThWXnFZl9dJGWr69Zg4zC7FC+jG67/Ip1QKMDecEM8cH+o4JBkwN4Gcn/mS9t
B8swspxO/Gzy9d+xaSZZN80fiY5TXmKP85jqcAjl70Kv8MWY7v4jGO+Xmw3vGOMl
9j1D3iO8i5HAxiH4q+JIJCCBm7rMsWGIFDonRatIXOgkUdkkx088ogodq/9U5dWI
iVB6oFwSDm1YkjEzaFENsZNFp+XX32HRP6LgYFVpbws57IYis1+Q4cuoiAvUvWnI
qwop9NpEWMfiDRsuMHbyfPqzPmVNl3mfl/gHP+rKb+XU9ragjee2EXMMv/N+496z
29m/2j016pjDsSRGRPcsNprdpf3Ht+ZdA6Xc+QZspIgcfEXkNxIwRxAJb1mCiIaj
5BofioHZYpzne/DbpFYwu9ZFPtEwMu4hYk8Zm2vvjJ1jdgy6w0hwC1HBe0dXYOPL
p8qp9+4/aMEEtmlH0OhI+9FmRm/GVeavOETOhLzA5xdwISPrpZOWxbB7M0rpNm4o
SCKwNDw/VJ1Lfw+751r64y8rYVsg0HOvUgDZsJYtflCm12ytjwegCbVGwOL0t0eR
mBCwMb85vyzsXdo8Db0YuFfdeyNrqfh1oEs3QtgICC9z5T0OTbchgbdDBwvJSgh5
HRrmWH37b73I7UcpBnpd+Cfa3Bqn5+ZNErC1Hdy9xlfJxRNy3frQMgnPOui7BltW
m23e23k4ZRo0bKjH/n56uBxBmdK0Q0uXcovoKh7/Tp4nzVRFdk/cLkCvxi61VymP
9fWgN7MityH2QTKrNbmdTkN8mrgXX4rhEXGKP2rjfL1CXT8jyQU+9jQha3XCaHF6
mKGVB0ISFvxGKPqkmFDe3pnuhF0VQMr9LhYTG+nKkVD4qGy60M1tuewNUV1bgBaE
vYz2Dv7Ify6M8V1lJx+XE59ub6Sr3tc8VTm5smyBKaO2HXD3KoDHnmYKKtIngW2H
78uFRNJKTsE+2dhmVbX+mRj/BxuUqjRw0n0yRFP3jpBEJm77A6UVwGd8LCuHEiOQ
jbsF1d0jgvVTs7Of8lU7HaeSqiwxGpzRtXhrwxuhTWHkn8ZCj970X6L2Lse26Sdp
tNJd/1svkuSXMKTJuB6eZz1Zb61+T03CL8OVPe2YCBfHaBFOtDLkkkwOU//wjKkQ
sj5T456fgGkDNABXWT2nYQjTS/xrL8WzWrM0XDflWVZ84ixqzaF/yCkhXDLhggjp
/AFbSXqtc0yclsRf7OBuyVMGt5kEEVxK2f4qIWRxh0Ml4nQu/KHKqE+/UB9S5B1r
ry27sNYnm37FAU2qTVnavrGWEhMwsoTJauZuXtDFpTcQuCLOzfv6Shp6L8EClv/Q
gK1MNkRJBmd1BQFy+3tz8+LIzRe3zInT3+ZwmX+V4jdQa28iRMIv3Wh4rgDdm1BY
qxoWe4k9U+U1OQ/xr9/cv49nnQS149oHFKrCqEhn/Y//RImHMTshNaWOzioccAVO
lN6oNQ4tIDicW2fTYhLC6Pi5wBvCtKso3WjKfdVqoy0damraNXQA7lNeCfr7AL3V
EguTjUpsRugpJNtftfOt7XBWgdQ6+0LJbd0BwcCyKYhQyGT30UY7ljxGdOfdeuMJ
5erwaMX/DP6Y3AWlT7Fc2bJYbMeiO4qiJ9QoGhqovE5UAYP/FwoKYyZuc6uoS2dO
5FYAOorkppkkk6Z7mO0fDlZM8uD9+cUdYnixINq3rWSlCVO+r3xKuJs1Jh/2hGPk
BcfNNFhY1kxyQgjroFmuT0vBwPxTrmO1EB7vPJnahPlfK5jEdY+gzY8kunf54h5V
dIXioXb9MtupHBxSrnPYeVrFDVSUljjxVjJ8LT9C906tQ4VguEfaXk14zHEVd+Pp
AiCqZfTwgyt3xKuAmsqNgwdCNTPmkJYewZQ+DBvWI+hxTOAn4uchqJR6AOLu903k
HW6q7J8f3qBabXkvo4IDUUF81bOsoJ7hoLjBlWR/WSqCCXIy004uqFiSjluQfBvv
zv+w2mmQwdKd2W59k0wXen8z2NbWR5jf9gOjgrDgJyJQNL0kLXKj1r+sHRkprznb
FlatkO6oyGTzA9h1YKD6ugy1i58hNbwuio1Smbvif9TFmsYIj/AxhvamgCOfAENy
D/95a2Ks4EXIYLzOR6AlZpoR/mzmx9dePTeGn9TFQ1Pg03/I6chuG4PId/KCg1BP
ug67qe8lDRGj4sr/IAr5qM0wIr1MkweDPmsog1RIPgr5BJ+0J5dntGlN93bWQKF2
fevXLZ6RLPFpZG4Mfu6sDA5Q/mSNNE/JkfQ+xJLZnuNOvHXysBrObh+KLGQNkzUT
FQ+u7O+3GMluWJCEzdVHUE8qRUgeGFDSOt6t15ueIfDqByGpt2oCJ+qw6PT9M8jl
aOXigbuZpUWzrgFXnTnMo9A5L8GDkRe1CX243UigDUhiQyPWRiWT4qcuuOEoAoEK
Sz6/2OKr0tsTdSfhbYE54G9tEd+77CMOPadbwNg+wzI7tHSYu/tjGqzUfvxvLnPg
FMqXgO5IiOoY2KnmUHO5VN3CubH2GfVwnVXcbdsRpu78uJSr2g+/wOLNodHZ4kYD
qJWIdJrFChMc9La7bgjYQLvVQ1qx5M7h86Ni9KHKqz3sONCfNFP9MNnT3vZ9fV9K
4OsgBG7uGGpxcfrO2IXvnp+0D/nT6p8l0udKt4fr36aKUvkLKeCrl3rwTNO0d+uu
o/lkQJJ5BnUxtS8X4wyAIJsA/eDAg1OE8+WLfOP7B4rmXnCi6WEnH2Bop+Az3nvC
sPx0eFHPZP5UBrxH/seY1wallznz3+GJZRUG6Nizx3VsxRh/rydHGQKH8MyhfIzQ
M90z39O7UN953sBu6+EDye1wMRP02HsfXWdjnUruwCwJQwLJPg86UqD1KbsS6TWx
2CqwWy5Tfdk6viYYhcJZRiP8EoV7SJidy6MQ9hGCtzdxqxqk24MKX+IDMVjV12+L
u5qfj7CmXTRrDjgHusN9E+ILwHWGn3e9U9cRrAGm+I+bU3e5+3M1KjaoXP8/DAcX
oW0DR4ysu5kc7sAs2eG6jAEqo86eJzT/ClQNLGxt7eZJAiwh6jaKazY9Eul/XNK1
rP92VJE6ZArNuBdCbjjMT2b7G8HP+II6gGheq0nFEwWmn0eB5fuCx4rgiLzn9aaN
lDNsf6Qc3oMQIBfuYOZnUv0OA1HzG8jMcRrkho6n2IPRKYJCxwYy6yL+pWk+iK+2
ImjoAoVNYt6y8O8LY0MDbRZoNTmzN7gKgdSmvFCOVgfFIXyQBpHvC0DPqzjOPyOS
J4VYty0Ql3umMQgSkmnupTCDMiO8hj6x3oCZQiBYFkTiP79XbTwhDKAcFMg3ogMk
4LgAV5AdRRVzfD/9gO4fYaq8Oa8FyUC4nloyuFaasP54AUZecTWD5+UYVN3yGtGE
ms9Chsjt/8u/4Bixm3T6O3PuB1wrVYwwSwQuLBiCmro/2CSazJFQbjpYAd6fInE6
mT384b1IFDY9hr1vRQh+zmygWXSX7qbLLeKpqbrq19SJhMCIZjrp8n01tcSs0O4a
pifBLY5nIYFIce2vB3Sm5yvBo8h30bM9MTz8KLPeM9ZmbxoyixcVRw41sdE4nmVJ
Und9bThF8TsTv8tmd3IzSvZhSFJ7y9YPy1J+S0imOlCvjKGv3m8oOSYVNaAR8IxM
W6TOts7zwtT8u+Me5jY8OPMVtI8Btv+gadQeCSk4BxhVOGax1hpC0IivE3GTjPLD
IkjeP1uwvbH5zqLVQuRPrrhOSZSk9Ui6Wc2M/fH9GLnFlQVLoVHl/c18UMXN9uQZ
pOcBs6uU0Mvjz96v/9kXDEhc+8RKcJp4SlrMHOTaMfju8vqHyIYmeKoOyfWaH+Wp
8vlbowwti17cd9z/JkAqcpGbzMdYfUPJ5jQk1TRWYeSWu+M6t8HEqB6sIG7dsIbx
BGhGrmh3YbFtFfKAdpmZjKNi4Oe5te+uFRDw7GjrJyGv23UwuDnotSYiwabjtlbX
hShFi52mcVIXpd+ce/WvtJYhQpDw2m9+TwQwT7KucyK0hj5OepURNlK7aq7FvS16
sF9imCQcUXlaKmty8KIsAzXGl0JNRrSU8sRXm5TplvGfwCcO0TthpGxfDRyqrgsY
0Ptv7JhCvYHf8W5rFuas4VnVDwk7bxTwAsxN6SrGXFSOF2mhpQHPVq3QhVj1CiJ0
OCf8j/+CjVyallSmHfL8b77Cb2AQU1TzeUMNMXqSMTZ0ss3uTbORKRoAWE5eXne2
LwICw3FoIoULJu5Z/3EW89XByX7l1zzxP++r0ZvUu327fkWRokxajFOtIdrto95L
d3beKy2XTY2CoKoXarMKbkJsaq2S2K/ILTB4d6EkeSBZwaKOSS94HaUd4eZipBBn
pjBoC3NR0eiraTbP/o9njxZH2/EPLblWgNZ5JhlQ4RNAuT7zqqmKbW9QF7pIwLlz
6Y3x2mTpPqn+0sYaREyIBHqAPdB+R4Jgiu8qX8Bb5iQdIYU2tXy95GbEosdaUoGp
iFGz/C923Ez7hFSyPLEos+DALtmE5On7n5yHlklUqJiQ+E3OoBqTAYVKp12F4OLS
MzrS7lbpnGxtRFwi+grrHmrtCDOWBO+i3BonXDR0zGTiMn4fVzWNf9Lq8QGi7cZk
pwqWmfWXUJlaBXbmd5Yy92+X84JNBXKreqGVIimNRjaQnXwjF6+8BEc0J1uJuLiz
Us2jrU0hLZR8mMBrKnmNBVjUkCeQac4rWa2aClrraXIFA5TFJnuBfBTWJoRKVAyS
MpB6VdC7Pb+d28AB1t7JC38t9TwK+qjAqNFrapYTVPvy1E4qzbghjuM32gOatcQ9
5L8kVzUN48QM7VWSNfkuBH5PrF+vRRdniL0lU/wDYze+NTSwbH1dInR3UBduzfLz
tG/eE5s9Y/N5wiJtHiJcKae7OKOLXqE8KXFCqxGoDZVig56FHzjKMusaufdPFwd3
RdYAiwkI3LynKF6SwE/pyp0k3rFGOBc1r5Sh3Zung3vIbL2Nm5XR3LeynVkl2LV9
Xg/MJgjHtUChxi+pA1uNomEOKKmNhjtXIjp3DL2r+D18a4KVZy4G5h+h6EVwsoMK
45ZOGjCFJr6w4QR/1/sx5I3L5Bab5Fiuphnkp5KWsPiujDH+2yQw7iaMdgnATFLu
Ysrj94NOPkK77oMPs4SV2XVAHxeSG+/eWTazXpW7lTHZnb71pWyEBspVtdip/Cpc
udGoQMrKY41YasOMJkdqHbG4DnJCUE66WCt36SI8yFLGG5TEy2qqeClywES+WgwT
3FncmGGjh09wDjZAzjWrS35i6A+sPuqo50K7WE9CvSHUcDG/pzP/N+cB43CSxHtU
AqKGjld60imRvW1RzyKMKotcLoczce+NluO9BKj5zOMnOfd6z/hZui3FChyzkfv+
6aE/Wl3dj72Xa5kPdxmaIr9xpuStBTL4SgnP9t+5GpdFowlMOCboByMR4Mi83U86
iEOtcfQlwPM3Rl7TwIaW2oFqYh9X3YeFGJxT/ADs5XVNwtqf+C/7gsW751fE8NuS
Seq+jj8+LisFHWc+GEfXaI7Ws7ulQKXcslFfuum+9bh2cE945kZo1n0/T1W8AwcJ
03Z8VY5Htu6gW+M4lUW+wnyZS1Up+cz29nkTlenEertKcw3y+UaA2pyxUiCXiTE/
mm/7RHAvCNtZrWab8HMzsF4HSXqiTFT1pMSow5dmi4BrYM6t0xKv9Z1Ea8aWfNgQ
a2L6zudP1/yd1Ot7Z+epv00EPbOKPwCPjmp+2hxDeI9IX0P+f+w/5a030sAjRpKF
pRaSD85I4FyIH8n54PCLkWKN7cbaYd5rQUX0MEG6t860ikW3M8UbeUvWhzuQC7is
/iNmsvvlfCb2OxtxmYDsMlM6sHlk3G+j+O2+X8UnTzZhAJY0OGeyFRLubqNeF1d6
nNh2eV4UyiRM+b4FptsWzm0CEPi11OroAlchVtGU6m9kYH96rzQVhyigIuJ8ACpJ
MxvBLKzdkWV3hJ3ALzYrR/v63D+R5VAM8kbOYZ8sDqAvbU47lqZ/ajTRoR+i/VT1
+dkSDXMA6qYEezZtD0WMAprb9/V0/gN/Hnj/mk1/LtkK4t17YzRUP9p5ys27yPR/
4mMdINfq/JwBBjn800Omq0bHpvAsbRckhP16GhXEaiBVhtYWwDRNcnSQGAoKMhem
bxelmDov1FZkfDyXugDPCuqh46YLgSXKPEfp7ZbuoYLLz5l8ZWX1EMCMYjyP/bVi
k/HQ0Vh1lDEW/Vrm+7wIWpNd59SxK2/Hb43ENaHTKowLP4DfUk2J71K2LkAqMN8K
Y00S63pY/1cCEEXap4opGvzDA3mv9zyJeucDgne/a32p76bR6B1LVs7zqMbD53n0
v5Ns7hswef4fzX2bswqetfxzapm2YA1PYrRjj6L7Ed8KmywtsWqJiUMWUixpt9ye
fH5uVi5xeK986Yxqm4EV5aUqZBhruBFfvsXIKLJGj/x2HplDX5LAp/tFM2v0aPLT
PYKF2/JMMgUlCRVPMo67QM3cdgqEHTdO0p7xn+WKGRGYYbLEeavdCqpmYGks4ZmP
P6e6gI5esJqYOShj/UGcIyn/islZMP5MqcHkG/O6OAu/JwFuYbrMiFe8R9K8HHlQ
O2ytDNngOLrkNeCrUM35CUljevZdH3vlYN9mnKNWmgA3Yq6KW+NhDJjmGEgYn0WG
afqHnMFN7cFfZ3Ezt8PPMgGOU+fBTYWUhQY87kAdfMYudCO+ZnOYGq32GeNp9UxH
VXBDaRMNtNpzajvZmtJVYXCRmInnqUQ22ZUI9PwHkmwueeaC8eVMNwjyhHFtt2Cl
WzGP700zD3gBZbboYwfysgcxwzB0tMLD70J1RVdvSQXLiNWTEqMiRhLYrZuWz0aF
/tj6zKh2md4+xGBGzwkwS77h7EMUT46ebQbyFNCfJg9waW392gRhoGIPc0X5bp6H
X6njoDngE9frENwj1LNh6XVlwFIzN1PSpRhhLBCLuk/iEAfVbgECDbp0dlZp3Vpe
/xMNY6fsJRqDjSho+BfUNNBU7PIy2ZBw6t+arjS2E5baXpKEgfSxXukRUDOGaX6E
pZaQhGjS6vbajHbM5hH/D1f7yf00UBLuyBuwhiaSK94uO6NeXX5BEBG/kJpkIwDk
sibWPzbdOPOqIrQ2lylokYHDtvYS1sDp++PER+2Dh7CysUbkOWwDHrksfzzC7j6T
ULZOiCPNYYO52MDxoKKcA3RWT0UVGRWH/Eu+yHudBrXPXLoYLsPKbKCFgR3diPXy
NF1F4fI+DEYa9kzaCQJPFqV778z5R6BXscLp9bE0xchAvtO2qd1pehG2mQTcbUJz
5J3z4ABP+lTZQXWtljM+1JHUa21bBjbR5EQ4AOo6iZQ9+dgSytCDmLNV3yo49THv
lTAWC+4LIEGIzrCPNbknkyjbwu22avwiltLRcObFtAq22lUpsBcx91yLcreTmRFO
9gnbc+Q53jGB0O6Oe/6xYpIR43PZRARJ+03w9kKYw60/bMDx8HgMEtvpCjCWz3Bu
GmVCR4VUitsrLMZ8Pu5QhlPX/QLimJJxKlXwfjfTS23sh/JhvL6xMetXPGiQYak0
90UWrhyK8OdtaJHt8UVigUo6NZou6HUkBuOz/blYfjdQ384Zqnfr1LqjQCCpQ13v
Y/rHDZl95JHnY/2J00RQODr/jNOIZrPrBmZNB4GBEiFk0BA5Vs0Srn8iOX8kzR09
kX4WzBBxrecziWHpmmZhHNY/PI3Bs5vlmD/myupRjNxfOXt0wp4GX/viPVvyHMwI
KJYCMVaQTleElMWm0ldjAm6+cwLe1P5LG0hbMMmp16uAWzJ24ruY7qkDyW8MTWS9
5/j/Lmx7rDU1WR1ZbIliUDbSS3i0mVsEuazQ5eYYNvgLmWeBDUVQnw2q6GIO0xGE
kYt0M0gt1NRUWpJUI8VRhvp7RM8PJZtufbbuBh9UH1UovNi6zlaRo1MPsXl3KZk5
/SyZ277wjjgNavE9Zr2LxwSuEZtMnZFcif/Zo4DPmG8ykCnot27JFgE/SVQCGaGf
K0EsA5DVg4vUTGowgOb/ynx+mRt2uyZR8z7Yqr2w6ufxqFsxsv4TPCAebsaZA/g1
AvmZ4lndIkqLAG3NSGo2oqKepkP8r5mr2z7Lx1hHsI8vJ+xxJ7aSO/QNZAZyIPPb
5BGeu5lNKBq7qVBR6EJU7upq060N6jT5SZwZAcE9s4bxSDgr6pStamYj3U4hygl4
5F95dd26RiTH5R4jxR+F9CbQF13jr/UipKk5PGKdox9odcqexzl9VHtHSEDa1IMF
uN4tIfs6/DMEjDNGXfnX1oflGxPo5BGMCIQq21W99gaq2gSoGqLd73CQHVFpRbSw
qI0/M9sUrz5/4fQoKiYxyl3Sr3ceXgaL875FW/eFjY4z4UWZEf4DTEnI8fRPCdi3
TbGTvJOyyaOo+PkFIiSgM4Jx5fBsC0O2wAwu3SW2M+SIkY7J8qZS90+Rew1c1d5p
IIou6rMF44uHfWT/7oEd45DUncC88dvmW0p4ddQVdAEf7wvLxqS2uyRp2fnsrG9g
VzRDJbYHnmadUOhfcypBS977NcGUUm22bFsnIkpmCZZFz1uDsvTbY5IDujidZQxI
jjBd5mGlxscYjgBAmmRQnBcDGzFtgysHKUYR50CPBXsJxzusVH5ZDrrBHZv26Wz9
/NQzUvlMWGXd6nouDNKvInK5N4Tqm5LF+65VIcrJQ+KsByaSGE5WccxUjIu6feva
p5KXP512uI/xTJX7gbN6KWTVpx59Bc9I6A8K1imlfAt7veMNcygIeNfGCzKYKYSu
lCyCLmWouBQhjbNTyd8CkUZwLbxGTxx3lYITl3ElzYSgzsIQ4YogdJbkwTliP8d9
JBX4ZzahfVlwx8GJHUdq/gW/XSWdwQ75KWvmv4xIFv4WOh1FZbFaQeyomudy/RNw
ypAV8nbWGKNPQYZgzB6xyXaXejd9GazUJgGtZHPBM6LQm54GqlM51akVQBWgztLF
VYM+hbFJl2M4oYQImeZW3e2yq6HUpZmQlG1KhoNUJe4vrLElhUI9CglUsAtUSDif
0gqo8xonW+hXLPVcnTjE0KY/TeqGhGyLzXKoLk0OUlSZuV9Kaw7b9TKXCkn7mpOp
ptqImELcOO66T1vhMG7AwQ7fF5sdr/I61cED2z8rSe9EAUUMVoWFFbfSO+7ocdVO
rNOdp4fzMRvlMTUVfHX2Y4kqOUZirNnapSXS5egU9YZqMx6wAwdZgCqcScWc6nZl
rtTcKWbmYMIlPEdfhzZe+HnyHugMzafblhAmAKGkfGdzNVr5lT1S9qy2VdQy5ud1
2T5tVKtMOhpOvNaeKbHKv8N4fB+xvcdiYN6uT+0NgDvp6PsWzoVtkNPvM6P9tmet
P9SjjseGv0Qt2tnlzZxHi85XtOKbGPnBNmxgGwSi6mVZQo7TuL7HJ1lVJjh7lt+C
tdTe2CyH3fWYwc/QUR3gvjRT/hZoiGBfoiOpe2dV1yu23nznEnmEDWQ+I19UzlBR
u5ckO8aU4kJ0nerZHNC4B6a2ddz7D3KF0JGU8Ai/lgUFspXzpcpi3S2MEByEr21l
SeXI5ajZPE469gB4fI/Lzrmd1YjP7ufWlS+EUhsiP5ic2Nwhh7W2yIBgrnL7fWEN
RIzYQjRdVr/BOjKlK1yE6d3wDDPHU9FM8ifVO5052z8D09tOyKnrCXmW+IwFXtCa
7RPzpoYOy15MieJo0Pq3S6kPfaTWVxjmi1wZWxZHPkVIkJK2dV/vizlrI5526KDY
D3rt8ZAQAs31x35gV1Ds35OafJGrRECJAZT34XyznvhP0xfeBrcvMTrbuL6S2DEd
m6K1WNoM7HhpQ9Cgu+Ksc29/wJQtBFal03SU3yv1PNhSeSkz0xAAunHKXCZUaHZc
RXZHcdb6hDn9ZZsVHAILnYVJQMtBWPCVRU2oZER6CRWUrhxULnhjcXNPiHK5n5TD
+lgMBFavlVLFTeXrHsRjhSac+O4+C5xg8zKZCwXev9Xu1mDmNJEIu+py0Ii8KQGa
R64YLeY5p+mvQy0qasNnI3DupRuPhyhgIm+3vtcPy+6v8Ie51kYrStVZ+O4dJ9VK
yoHgS/XCkixOuu6AWAXjA77cSyBHk8xlobkIDqWISVPw1dQkAL2jAaQEjYTr/7tB
4njNQG4Us+u57GpFstOUvY3BobM7SQ5FI+DdR5kAfv/KGAGlybtS/jpv6nPrFBag
lkCK3oSiKoDo0ouCDjRF6tDpA0+2VWKZ0aCLna8GB8HZ1dAsu1HYMjreF05hRxsM
wtl2Y3RqUEdUeNXCeXwZuNtsJK9BT1fI1nZh3Dv23QLVqGxcFLLTsfRQs4/7haJ/
L4y8MgkQCiF+oIyvX7lpS/1ReaTK8cJc0ZGpvN/iZTYBJrK0Jdc0h+yS8D+7K8Nk
xhUUuH09QWogkZzrTD3MJD6IXCwEfO/6b/o8BqUyOfHP+LjhfYxErCvdQShv76cB
Br2UrQ80r4f0v416gO1E85i3xAQ95sMXfijtfvnc2XzpEK49WbYAkiJusVyeXt2a
X6Cf1Uwj5JMp+QAMYyZey8M4ddpGqxobx2QB//0Blza4prGuFXZpVfAdLEqgVEc9
7z56EgkZCHkK3bFFAp4tQYvXM4nzFXA/UVK+HmHFPaz64BoChPmtVYw+RIHVBS+W
LzJDEchsn2DE5gMB63dH73nxNfDYUYyS0PjdfSKDa8CJ5uJNnoiadMvUHUG/I4cR
6mf+1tJc4+KY821ZZBLoo09QgnSgKoLZJnVg4OUmkriK9yW3bMoi6toUjh4GRSi7
V6lAoPt4jTRXN2VaosKWMkp71ePaIj4CBryhJis2MPNffqUSLj54jj3h+EZIHljL
8dCFmsn6YVZq1nFWjQNenhUS483Zsol9+Ehfzzf8av1bjZUylne9kDaRiAPgXr74
v5SdrrWBR2gUoUKCr3G20tlQFbOMrYmp5QylcbSCLBFanP1wg8IPN5QD5zU5Jhyy
eMCWhl0kptuyNGFgQF+AHgxAWWdDlyMxD+81iLq/ezdXoAYgpfZVpilzqqbnrMCf
2fy18nEwBrHImsMllVttVTZdwZtM1Z+bTKYhbYVWWQmTULvO+Wih3VA2sBo4Zjmz
LQz85tr4slR7MeNpHpkmG68q8izeK/xVrD1MeaQxwgDCxhxIwmiJWVT6KvRklSrD
ehfNYmbNpoe67vGiMgHhwf8cdOuEkda4N04LQYWbP1IS9JbUfwKDb/2kwZFHh3t6
8/t16K4olTHkbphqiKFNOM/BcWywVdN4nmnCRGDL+WTBIYyLQa4f4vt4hF6uDCMC
jTThBfjA7BmOdrWvieWkHnfjzP0QHqF3kqBUY7BhGHEyfrTrNiGB2zYEPbF2EIC/
Rui8WbdiyjQTPS//A552vc/HNjnIfEWvI9BmOmXyGKY+QcWlJ119C70pU1kQOr57
WszYmbhOluewuOPLk698Sfei9PYJ1dyWL7HSEWOP4naDkqcB/uo5eSRGDiJen1xv
7owKdNGHGFyD2i4crL5cRFWOZ4DvF7CqxDpbHbUeUeCElh49wCkA93zENEno9pOC
M5T0pv62X6mzZFo+Ise+RqaWdS5/AbowHAkW9BGJnvtW7UPHmmCO9XdtACzS2N4E
FdUt6tFIc0fKdhMA1mtGSJaGOK5VHomAkDrKijUKtLCFWaVNrYiXduOAsG2BMD86
QGRw5ZHKkzDB7AUoSE4zSbih0CbJcByljts2odWLWDAmHWSs1qhj07gEnaPJ4zL3
8xBBxtEdNgB1NRReOj6o0vXhammRD6D5WwItPMsc4Bq+PT1R2tF7b9pxeCjdbeUW
pCyn+JVzSP6IsOiviSX41d3hrDa7jKV85fBocXghzn/eT3mkNJs6vHE9trpiH9BI
ydiXjxDYnSSN11LYuHKdpNLHqqdSS6RGNMEeM8pOjsmW2Tq/Rr3sePnBY7KC+xhv
r+L3mw4G7+nwskEcMqS2TID5B/8EVhifpFnns2U9EceNFCO8sAeIzh+vK5l0V6eZ
PvsCwXRl4NsCfdZA5qJZMMMmCLtP5+tlw9dYS62EIuoSYxsDaEEXvi29IHjY5Fvq
H6IbUpZcm5N2rtQCSYYp5KWWRTpFPWMuDCdt9n5qQ9j3uYo6zG6J0xc8w8AFVvt0
aG9eoBlMfO8aPI1ewtTKIn2zLdQCDkItJ6a39SCvZQYbJdNj3hL2HThs5foBBg6K
HxQ1eM5jopBFiZlZPolXLjqAEx9m92tcGQc1ePRUtbc740dPsSxqQx0oDTPVluBJ
GH4VtHfBMVmwVt9IyaJ+8mU2rKj4kFlNgK5dQK+/5D7lGMOMfiqZuW7Ocp/c5HME
e2xrm4ruzD0C2W8kUC11aZVabcvoAtefuHzdo6No29GwS/ypKWO8pnI9yf8nIP3w
LAllKTvoPrE568H6edxETtwQyc/AbNhdNfUgYOQRkBKz3U77mfFOJE7TFxmTfRVL
tvcd6jPUxb1TMMHC/TQXRBGMk3v/sKWJ6/rmgAffSDwSVBW3VtnHtACXZXAb0CUQ
m/sexu1OxLOoToY2ePaueZim/DuExo/0lqtgnVdsCsxrsKW7S0SlYDWUjJPaah2n
EGe1XbOoox5gvXZePqYBLK4nnGkTUceDQeMCOUkfvRxaHCboNDDIiYvg+9DqOgvw
atLcz7Q8BVaXOBpJDVENMPWa44MaRAZ+oVDOI8ztFvAoweikyZ6cI3eFPVasNqVn
xW+nahySe7uO8KVkqw9v83cJUtHTBjOGOttRltATyvUP//RGp+ArNOoT/M8nnhQd
l8pOGVI96BNWWGcr2v1zyKip8CLDTzsgnsMhSO51fRvnWoek3hq6idY7X24vR8kP
IZ2t+i4ysOBaibMk/2um1ayMFlitFbFAa8PgeCedN3e5BDEwUJqyIwcGArwIsT3k
ZVTccsdKPR7I35mZPAKRCXII0v7V0LbeOE6qqiwg0BOvKGHHKiwXmiAVNmCq1gE7
HUFaek4o+TlCjnIK72xZ3qdP8qZpwxoMOOLq0cmAUfGnBPBbkEGk5dLkEkdD1pyf
snso7/A2V7uDOUgcNqib5ZQ9/z+py+85rDl/ucl+xP5wklUfKaM95mRnrOeWiGH0
NshE5sMxZAyGPVolDDIDn2tEvEoE4xOoys1A8HY/9BZYtkDtE/qSnJ3RtBABLAm6
S9CirN5NqA+jtUd4Fw4Oyf0v8svln3D/vb+wA6fpULKh7MJtMqx7adfnEPSj1kUR
xsqDgRvjXapqHjvOtjh/B0ukho/2xCb0Lb4q9H/nnk8mF8FICHMQrxKHydilWMVU
gn+Q0JXHFcm4ElBGY0KdJN8vgZy01HPm9XoBBfjLf8nOVAHBLV7BA56y/O0IGWZ5
V8r0t1i4N5dFYZKCUOVFmIOfxxozg9FHve2x/C8JW4EvkUhcIlnEHxwPJk36eblP
3mprgXhQEDz7ZSwo3WaNmH4l8zseI9EdEc5GSv9lJ6nvw7COacsXqhGS6gT2Rhqo
FaBzM0WSCXc7MGWPVX1sPpy/R4aXQ5dk0pWd22bdwG6Z/flA6WysKyWwDQP4WC3Z
uQMlGB46hJCRRyhOkyG+JAK7bAye9F4018ycQyPww9V9bC8buqvpGo013obsT+PZ
TDec2tnvWC1iZiCPbAVuIErQlyOB1FUtpWfQmZuBr2tVEUsXAq2mHeiGV8ucRVES
RNWVRf5ueYsSk9//lJi5SQaxQYR+iTak+KiML5Q3euY6cyQ2qOigUr3uw9aQ7txR
z9tNx/oXTxwIA/OI4QhQ3NhOOeIFz3ifticZ1Yc5DVNC1P8igGuXO+c/U2Tmj60w
2rzr6+xg3MP28v8sSA2gbESNyfPgymYc8yJeW+RurbYBkZqlCJwpVprofbdNdJ4J
Mi6SghLq6XPC1u1adizmHTOcf6EuByG4XW3pBt5O7ZmChxDw4RX3SYBc3dUN81E9
z6cnTpU7e9z8MgN3Kf/mO2th9xtEyQYuvIWIdolKZfYBrMShW78+0/PmY44RNyMi
cZUBrgYwWulUhFFGaA3YT8JisbyH4U8cGKlRBRVXYOAiuECYIo7G5A1dxpuRFJJg
GHYNzZRQKqKbFceGBUVed++v4KFQue+/jG7m3G6d6hmBwosRspdMbC4Qmeo19aar
ic+sQ15n8chKJJSBuO42J/CTjFrwoE2/jchtcEITdgq/rL7IN/PpmCa2DCHCq4eV
RvqD/DDgP2gEeWAy+0RFWxZVZ4wkicpgtAqm9VJNnMBm97KM/nzsgj6hp/Nm9ACm
mQ7Ibs1RzsU7f60Uj2D+1xsGGej65RVsg3fVTRmCGyCo7+acUCP9O+/bHrq/vQ0D
j1No6ZoH3GZh34zsGBLkWGx0L8zKsBAyaKqn0Kyy0bIg++crnet0z/BVe2Tmuj9O
+gwNe5LMlLFERDQ1jwbMOdgXXMftjEQoZ5bnceO8Gl6Fzs3wJc4gcA16GCw7RguJ
YHuN1nlgjccN80xHr4K2B03h+ATgr9beQnXD00S05Yp9qqnPydMju5x9XlhUROOO
PnBiZhzTDcJb2tOXeUmjoo9mqypLp9ROiXg4xhURHMzdZot6lvHWviwCZRWGdsvp
r9S9Lw48XEnZyCentTuKWGCw540C/xBAfNcOAaRSIj3aOJ0XqQL1FcRsGQmzSoZW
aFUpc8Ba+leqH4qgb0MLsgq0vJ5aW+2UNTzmNc6WT3JpkXHTQYL7tJg/gjfydXqs
GwxSi11iT3VZMtG4NgMKGFJEsZ2ydAzTJ8I64es6Lx7IJMXr5oWoRWb5w0dXADYv
4PSIiUzehzAIKQi2KKgaBvbmB4yh2NrDPok8fQ6+VcLCiTLPzalOGZmJQuMDeHXt
zqXUBcnEsHnfAXzfk6bD/3bnX9pBNdmM+/MwC5Gy/Ymmr6XbEJLwQLxpsrL6wk4a
kSK7HR0AQrqRD42aIlSNdoAUvXzdMl+TYRVbBYUqjSJ7u0Wi4Y+KB+U7fQnZ4cxG
CBiVZWrbAP8Z82GDQrixSJ4SFZrL6/fc+LE8S0RcjStezmFeiuD2rDv+MVkqYJsf
uxi0MY7g/cVhGskM0lt8qopPS0p5GpDCy5jgrjRSJGGGB1Y7E8e3est25d795ObF
W8thps/vF1diezBlm7nyp1Ifd/6jV9nOAJjSNSBjsGwyBzPMJizUao59VxMJCGK/
GvMhjaWrbNakjEPYcbK2eDhCBrmTtbvgAB5thqakD7vy6CrK+oVnIvPDdsHaxu3v
Q8/5z/2X/BALNxN6Jjo5MrwOwQc14oPyPsre2h/fiibyqJUoXk7btTKy48MW2P/C
zGyPmsKp/Qq0UMqm+8LQEF0bPjQj6Mr8re6tUmkKT/mdcOuH0ahmQf10t36Nyxd2
7IaYED4KCAPqzwci1DW948DSqMWldyFlSdSKmwdqPWmcyon8fj0JHcjOIoYLI1Ax
q0KpE3Ra6oR1V0wzqezon559FgnPdpDDh1dDLjpeLHUQO6DDE5zFExEPjnsse5EU
6usQ8ZwVooK5MR2793BFioRITX69Pks6EhL9cUsWYl3LuDJCon0HDVT1C6CwStu3
iOfREKSmrZ7rlUcKWh5qsx9U+RfoMyY4fBOTmPCiC3DZRyCxNMnigz4b6WYAQYj4
kNuYtc+Fwo24tnsAAzXwlAUqdfXzO4cGgpeCQUvwWwjMzHkCMOPDzxuyw+B7dW9S
WpskmmkcNjjJ/HQQkhCCPFZuskCoVD9yw+NRh6P+UWtoHvJQpg9xNv4jpT7G2gw/
rl8pFDVFgoDNCOiA327iXkL8JuWL6q88WmqLqse6eewXjtm4lJTFL6286bEqJEhL
fMThY8BcUfxa1fq1cNOLxcra/9jBqjmu1f53cW2IMynoBuyQSlHmfP7Nk6XzGB1y
iTIYxqhvZubRavjs/o4DHDTj2XaoUYZkbquKa4Lz7xEwrIb/KHf3T4tgwHPTH/XD
WX/FEV1izn3ubfjB5EYRxeURaMWJvGQnYoqdA1VRAktUO4yJ28yoh5V/q+lYAuqW
nAKy8JuhwhV0rZJO4k4m8cro3SUWbxe31M6h95zzN8eb8NBMPwozNnaF9tB7xzMk
oWvzqE/KbFGBf4A/ZjcPKdvi0TbD1Up24vXjHh0X6R192Yg5HQFemPC+SMpOEi0K
4YK/1EW1gO44ZFZ6NMT+PnmRyK4vzcackFEcV1GHRSk0cyDwiOdY1RTMFnQK+8yC
XiR8TiApszR9nG4ss+MP46EynpUGFDSqXrPE8bgXQR1VVRBfiGlHaGOMdkGnJaVS
xIm9vhzTvnVkjoFTh6vJWkfMitMNZicrzmf7CijpXLb+TAK1EXsCIW8sUDU+EvG/
r3RjVz7QoTGm0V9mHOvKCfUP8/WVvDpu+5CjTk30cZwMM/dqOkrZSzMD0JfVbjmK
Ibdn6MnxFEJFayIKoTIhK8/k7S9jrJ4exSUM8k8HkjAt1DPCoS9jVWqyJ5aWmjzb
KJF3Ug/r7yRKu51u+kfKl9/Xi8UQqZe65LSVRMRWPQb2JufabxMHztp5JMRP5u0D
XQ+0XHHtOycFxGRgbcVAwbAqBPPB+shFJcEXjulXl6Ntn+ogHOLFugDFCD0JkhSL
uJmqE55/kjWqryUVnOA3xh6+Dmih7LGM05ckTUS7VQ3tC4CeFAnDSXfvt/UhaXyU
JHhCS25eelwh67M2ZYdpvcbJbq2RjGOLwWtk3MlL4lihU23ePLzyq1l575tt+yek
idYF8/xgRk+6bHD7S92kQm//d3vK2Px3tsNOH+VpAnJkpbRdGd3N/JdfwXKvU5w0
MXwdO1k4eaTkd0ZHA1RYIjwmOV7cYqsjNiyv7s86HAmzyIysccIsB/aqddXVFOqf
UZirVQA0H081Hq8pnSuOxDy/qcrQjkA9tnb8dWQWXF4oWNC5VSspRx/7TzajbZdi
90JMa9k5Ib1p21UficIGNCfNIQoEPH++MhRRES93tso5yID7dc4e2tNM7zNk8vrn
KMp5nVUVPWE6XPKbrDq3ZVsOJ/V4sTb3XjMtG72XnBMbtQ716QTr9smBhHUSSQOn
mrzJ47vcgGDD3MrbUgmnvTeTMpBC7RY9kOtF0tzS/BveF0ntbHz/V2YnMbDACu2r
31fXdOwVmxy/JKHPZXjaBVmdvKT+oEqQ5HTAQJsr59zEbu/DM64A5XV1RuvhsN/H
W7BokHGFxkikIzZ5W7P8lQ8dMK37Ds0Jur48b3TkqsZjmmuCAhsTOlAyGKEG+I8B
PRjNFWhO6f139GiVgZuNNch4t3UxGavRwwLWqGEPilmszowTS2sTnYae93F+eazT
lyvmEipElGq+iIt0I5zuJt2kRBnP4HO5lN/ekIpbfXP33+ZgrbU61oUv59mYViXb
j/8zwAchSFK3JZLNOS32sfG+ZgdUihvAon5JuJo0Vxvc38kM8aFnj9hRCOGer2dn
eHWFWxRCqykW3nMlRUVEsI4Cgtk9t+xzIbmcVjCF2EySrYdEa8JgrCO2IGVmMwtk
C6VCl3F6S5C/LTz1F9x5d7snrfJgz0+l9s3p+eG4frYX/+/s9vEKgWlx679/84Xd
RvZoaYotEDGgxU6WUXx2NgmTExdkHSuvVJThkX3cY3p644Ig7ohihdqmE5sRu8eO
dgYuNNNJ3/vajyD24vl1xc+/Iq5ptP3Y0Fy+cSpUIQnrEE4RkGtS0U71HzFyqCA1
BpGBetrRbt8fpfWZq4H38VPOKn4/RNPBHihIRuomcOblJnapvxAj5ABwPwdKiqLG
tAErvRlOBrT3KqirAEQokkXqz/rQ5Zjp+I7cYs/Sb4KgtyRZ5WfKRxNB7mJ1X/ss
Ch/Yn4aKgRWixXzMAeqpevInuDfYi8KFwcnmgxYxJvfi1Bvoc3kV3FAgwgqtypqX
ZNtw89lQR8RICJlhhPwlRmn+u7hEWMUDSfi5schp3fD5pMWOnNVYJAW16sDMd1Zw
Ptqw5JJdsRT0bq/m5shKbsaMNCELgYGzS11xxQIhLzscNe3x1a+ijhSknlw3f3Sw
PpCSItGoSKbDW8Tlswjs/yuGh73PEuJyeCL40TNVBPh2mKDDXN4skmSkl1q6XXPu
EZvbUbIztElffGS6nRjVWzrxqIEmFNl3tkpCijw2o9vdF4upOC42rWz2z/C3ZdWh
Kn7sMSZfeQ0bQS7CXqFIXEMcZMxV1YyrVtqPmAu53RcJO6iK7VhA+fvMQmPGGsT5
ywd6zRKeneyy1MsmQJs8aSNyEyytD6VFS1GM7RbEc3wUJQytuA0YXokJcnypn5E+
T0v5iE6o/+DiepU7+73eBmGVr7eF53mvYiYEIatfgIhJvOycauUl6zgCnKwb7VIM
RGq0P36323iSO9SF0tjyfT+QWsJpynVjEgyUVXmwXAuzXVvsKGKnLD3hMq32SY5G
kLSHcohKXQZSrlEgmCEU0JGewo79ZEqEVdpvPQ6RL/jhMQaMXPRWiFQME/w51vCm
kifQ9aw0Vpr5uyOEeKgCuwX0Zbn/ytus/O8oGcMH8fRa4xZhw59u8LgETb1NX8QT
wsN1WcumsEsSK0SEo+0c1+Jk7HBFnsG8y2LMeuQjEjK7wa2adLQH6Zt+Xo497rOH
1yvj5Je9CWeRodg0cH8hMlHwP0gfIcHaK+qFBhQ5tTGvdelEog8VJ/CKalWLYN2z
mg9J2HLtyByIBSTrqTTbNW+EWFRRyVIH3hRv3soqRS4OF1ADmepSkLnQNFu0W7us
hICdL3SwgCfx+P8mv017o4LQI1bqLiuXeqJ5dbogtuSAnOY2Ocvg4ugkNHUOXdbi
mcqPoXInCyMLjhD5le+jDlQ4Z1STe9f93OkVER1egPWjYC5uPk6HCLAjD/4n8CBd
BXwq2hhIdtc5Uv8NaP2kEd6PDdnvC+se3dlYihLnQAnvu6RSLL08nuBzEK+aTW8k
xnecgdVZvoqsfe8TpUygF0lHgKScTCwGCKqTkWMROLNKxvYvrNfOqITde85MKqJO
NRcJkUzDEUjMXlZ08Vkpze4oHH1baEA25cwf6gppsz8g6t4or5jXwFEOGOFbRhwY
it2/v3FplfU7Y4sFurDXp5MJ/TPltUSF1V0+PePnT0Gbdl9qw0t/9S1wnHdk30PU
OWiIxFzsDf0RmHE2K5Hi7Ew8vdFm5EKdZE36YvRb7EeCjSQZhoFkOOqOsKEiP74v
DEr45DylDDA2RhUrx1YZfKTOjOVBLa0RK5bI8M70QJttNPe2WPHHaF199V2dfvVt
2YPEYDv3AmhmocVzFgh9p9wStsKOCVUx2hikBSZgbjiTE4pZevyH01mkcqUyy2kB
QjQqYChvqOvuvE8FhBktG9r55Z9jNLbBsrfYEWhdl/SVrCRMlS/JySTn7eKttM9d
Tvn/35CityR3tXe/bkDehB8A5lK/q4HRMT9X8vcSdeZ2kKXswOk1DkWJuB5unaWg
Dh+COugYCaQgVX9IL9eObmV2XWOg84DgkBvrgO4o/cm++JGb9tNHRZNk5BPsgub3
FEu/afROo7SV/4BejkyBkeWKB9UwpA7HH+NlIwphUN96ZESqkxpfJMsI6+YRunp4
71kbs2YU+zsr152WSWRe7ueytQTm6kSy0pJsUwfjUnBui6uwv0QrU9R9YXHUiFaF
NoNB187/OJtKMMbcKhKKHy2wb3NLTtbZbRlEI+itt0tOx9XZUqWwCmplLlW6eYLG
egWj+cr9urykAiAASQi/G6e0c1uCTSHF6/o/E87WvyO/LFi6nDNvGiMppPhRlXgG
MRVf+/eILKz+OdpSvIlEj76H/5eJgzEFobUZNcwmH/zOMDYL/cQE2v4JEayErbWA
S9xJWo8toF9oc1G23ERHA51/lQ579pUMQY5ZeJTpIGlGe+62dx+8pP1tqAuUmAJV
dDgLcAwA8Se1r12ZAMreXxjun2O8z6kWsBQmpsprDd1tZjS+Mh8AAgSFNbFCxvtB
4IJgHX+wTIrQJ/QxRwEK4TfYitnLzt3PVHqT2i2QVBempouGrHUqZcNY+H2cvx/e
NFSmCu6JKfgLN2gZb/ML2B3abq3ArStnk4jHsI+qK3cWHWywuYjRoepcSyuG+wry
uDGF4yvXgjATf7fD6h4I1ye1B6tef4vieP2Y09m7EV0eBKL82JqKHgI1WDEHO2mf
CxyWvOTisxIKYK0OBw0VOVEBTQD1MewzIqu9Y+IUJi/ikQvBOVODKiWqMbdDCybV
z/GUr5K919Rfwb+aLVXsGJsKb+FRBNhB2dqlr9tYC7eEW10wSqeqPdhXxMx6MOqJ
H/A4fQjOdRbt3XzzP2FwtvIjfeA7GInz9jPH33/gYMj6+kO6KsPwmvTdsXgiFYWC
5A3pgqLwIrmBhL0ma0rcmfFHRBxQxy51fh3kDhb2m1ydF76Fjk16U9uniJx5KXgS
xwMSR5p8eRoP9uR+jOPo26NlcGxu0keqlhKmYxqhHyNEvFmB6AAkk3dY83SIa6Wm
cU4ZIpkCBQwrp1APUM1SaSfAXQsTFSVyo5mUX3WAuKgBIk/TBO9NxcrB2hfR/iN4
zG2cp9xnyghCzQ+2w+6Qb4bXX0wrCHEHXd+W4i2Uo5gDqtkkpY1vLWzZBAV6C8Xl
z7135Qo/dDawNrH8my8nuxF1VQnwTIqyCycG5RttF4WHnyrS6c3g/UPvnxinsmc6
Il+QL/s2INjRUAMp1eZfo8SNigKTp3upksFMzaz5Mcit0LPCBStgh0wXV64A+lvr
hMWwBBJ/T9P6myXpCFewYQyJEAZs6kpmrFArk/ZuZHI9o/mXbxNfnGyDlH+/BTvM
Zj2ymyy5NdbEqqzA54EYHLFPtUM6K6nInPF488shvgM0dmNQDZ7qB9M4ArIMoOiU
vbOYdZ9rvnYgtW3YApaYo8kWQ+QNgoPNQfTKPoT8NIxKxHg4b6SSJpukSR7w4r/v
aFysi5Zkzx8RhkPRyvU9Zq/w3UVCjiVm/K1JMYBJWyUMBOlPeQoeLiBiAB4iz1ZF
+ywPe/qWKP4OB+5uOTZRpBT3iVcJapbQ7twcsYhox4PA8QLMarCVyyktzzLn/li8
vgrzMb7n3pe3LY8D/CNy5akpQ2sBUTusiYUli9EvS0p9OsblSp6kkNrBt5eN8Y+Y
7ReVvIVjAhgN/6pRTQlj67pXn/UJSBujfILlKQf0vbVdufimWiDzJvqXbocBh4Zm
VDCI6aNxIQodLCdahV68Si8Ilu5whij2u538Wis8gYH4wxIL6fyt+SD6poWIcWh3
zd9Ios48MJ7oRjBWc+AVNWbvgk2jBTKIQeOB9Jo6pM86VhPxnzfwmA72s0OFBzsv
iS16S0zcgc/jH8Ape1ts/707AlFlPwc7bWJb4aeALFSEA5vDoCIY4wQ6YxaEQdwl
dFF0XMnof3qY5naZFdhMEX4JCyWJAXYOwGUlUhZUaf7Glt4Qb34bxAv6gUrruYUR
Z5vJb83btrPvqiJI7kWuNiAJlIHHxPbkVNQQVRvLP6Sbkvm0+bhULhu8G22OooQ3
xX3AtJ3F4+SaPiEAni7cGOwttmRXl2JJLJh5wnLJ0JfESynzl2N/d1/Anj/nRkLE
5ab2vAKdiWzXs3L19IEq1XYj+yrYI1ITxg51xgiCS/4GfmTJKEteDOYNMV4x26MI
0WsSK249kXWsumA0u/DXLrrHkVhxqsew9WFQsG8yZNC+3N73UBuzNYDxj3BE6a5Q
9KDjm6FdZ0gzi5JI7vlE7W63X2vLab6Bkjynkjv0Kjb3g+qcH3+MSniV5F2KcqKO
5uqfZNXsXTPqeugDwqdAX8kOSUj/2N5B5PQIDhap/TUbMg6e8vTqVHw9HrI70iBT
xCRq2QtY53qNuaKTc1KOs8SLXyZYadOLlq1A9NcwEmWwx1nEoyMtLufbzeNEP6vI
jaNKBiq23eJ5pBYWM8thLXi/9hbBu1semjE0+tU+6Cjt0GfTJ7vT3/0u1XG19CD0
vH2w1eIeuOqcmACjd2CI9GL5Tnqq/Tk4CFXmEBhZzuGFNGdA72q75mlkW6H7RzuU
NnFhsMgIidun53RLBYSHU2d0pr7kRysj0hIXszt/XkGssijxqU+215Xc86X+POI/
OqvCD8xKIe2Le06PeTcvDDB/tC6tAFbqT1CES0hIEIBBWcBch7BS0NPxvvIZjxfJ
lKKNclstqkvGQdDWybqhy1FKOi1hZahC5JMWkRYpzymT8en88eMLwPHO0wKXvQ6G
yivXRRWJHTAlKnc94Ze3gEoHy3VZmGXc0zUsp1D6nJH5+VFcKN5Yf2orCNhjsOnX
pDIq/+1GxtLGQzzWVPj2atYvaDu09WMoVD5AfzmjWPq1sKvLK0Fr4HejYitZVVMN
QZFerDmU+8QCA8DdWdJa1HsnjkeSbTfPnVV5ny+Ivqueu7IHRtZkfXg0kd7f0AI3
6iZJ80Z46DZU9f0XBSu8xlrce9mA/SMen4dRZxjWcLkgM/Ve5U+EA4pc5NmgMGPy
5R/btoOXVWKXlnzALdniS87l4m/lzkJWZpzMXUT9LlMhf6EQmVBn3KbuJ1lNdQ7G
niZHY+jdV+kbkQSO9x8huypJGFI6Cy8O8G7B1KflTDJYtL13f628JFFwbtUSevt3
G5LCk8DdP7uBPeunOVwqq7TTJrByE1RcULVNIoeEhpJZ5Zq+XSolAUeoviq3GneU
5cwPV+0CcY35b/NriOoKn3X1FnT9Jkb82CrGewKj09z6mK0Tf/CU3RLOeRjfxdlP
JYLCYXMQgl2K1ub2APxPF8G2hN36umr7VEH+up4xf6VufEMCcr5pCAYeFFIYT7/K
G8XgnUIK//KTgs1xwOCzyew7IljFJlHuobbIspd8l0ZvYu7ZLstO/ZRNHC0+F5Xi
vKwYkpP28a/kY/v3U80jiclc36d5tdu6hKa5dp2zKvMI0cIGtGwmQpUBE/jq+XGS
Z734VMbjQELRg2B7AN3824c6nL3yzTprH958R1YkYDx6gZ8XqFMWbC8vVOA2aRQl
oMJUl8IypbZD1fNEH+cnsQBAQnIADdW+CE6tH9U+7S02ymBVe7fXba3fWwpGiTFE
KvZBJFzyCN7Pb/2sZaGF4vjFMeIJNOxwIHjW+1O4sJxPqf+KZzb4Ol8gc/nweQ8W
CB+qCelf1Au9C1BlOBfIzn6Nvn2UtT8dg+3eSQ6EjS00/NqCzwVNwgVAaJxAarsF
+QBKtkDVRmniOuJ/ziVTMX7gaXAkkYGn2hOsho7F+YOhN5zw3nMmmfTVMMqhf7Hu
iCVbc6BEwOEbI7DbVhqUsZKqjAXY+9rlaXTM/AmLCkP/08rHkqg/0o65SP6wDnuk
u7hWCBjABUl0PfOxFt07dpVixKrbVTFm3/1PjbaCFc5sK50ANRsWKm7g3FHgaohv
eQ689zE9PIc9m6AYfF1uTMr8CKujumducXiMGtulnkYkAsUPqbRTMlHNIU1XDtOQ
PURLpYB87bbWQAKi1bcs+r0RmC2QSs2BFuSSeIFFZmyZIew3/8f9veGQ//S3PuoT
SSDkMykXwC+8+FKSDkvcpYZVGsdB0F3y19onr09PBS9/itXunOQT1AirfcocxA3p
y+KgR4zoDbznXieKFHS3w98fIInityHn9G0UfrMu4o5hvknV7hw7sgotdVaLiG6b
KdPI8pru6kjG8AiwrHRG3ZpuA0s7nqiFs8Q6JQ67oSG9MbnyjudZ7CFmwtuYMLg1
bT6DswHTEwcu9C/95zOEV70gOK5xoZY2yhSZiUgef2uVCbowV6N2BFanhFOOUgTM
V/r+LUm1CCFWNBT9HqlZjYpOqrmz3ZpxoK5F8OTCkhiMLCQMuw17ZfM9uAbtRr+0
sq5tylLhtq2/lVFcoPLfzmJwH6a2uFPd9vFmgPoiRsC486oTlZMpyTLB8bgMRxMJ
3BgCencLzv/wVkGire5VmcyKwNjkNZr6tIkmu7twqX0Io+l6kKOpt2VcHc6ZaYRH
jzV9fxlvFSor1zZt7/7YCnmZLSzbenZ+w+2g4PTGDVuJuk3KzTVgPHSSWtFl1doN
c2+EPQZCw76Ef0FyD4471nSUja7QC5xayYv+bkbh15V99SAFJYsmZAiq5BeVxeUm
aXJ2vsNKn7g5bKi08AoI3Q/0zmr3fCNZZt2NjbBjtpZDDVDgo4juO4s/uf4lRALL
jlM5kQWjnPu/r9DUg4UWMqDJCaSVNtv4y2+qJ91OqVcnh7wXs0iW4F5YtJzSjrVx
ZaGHW6H9lCGiGgI9AdnH9Pwg42r3B5Oy6IthNXxo3Hj4rhnj5YoVyi1024oGbYwt
UK+fgY+Q9X/GM4xe3ROE8VefefBHbJ2e+WbSjSvNELdNlGHBhkheQvNHbtsoB9Pr
0vVV4V122t/lntcHlp0mnfKeS5QcRJmpKlbnkL5Yg278nAQgZ9rkGDkiopNRXuoB
tKDgC+RWt02XqD0Jx8F57u3XHgxFsyHxYqVlBFQyGSnaesnyciLRviTPihDPlasG
lVerwC+tcxUYdUOdFih94o857NTCBqs3JGkYtk1HA4LAVLaa5CqzCHinKHLV6hJ2
Lf516yICzDqUm3PsbujLqtnDbeSHf+Sp/aa8uG1LHqvv/RLsKZ2HXyk1+zjTastl
l4mexIdXgufoFDKXYKVtpIeadAsxjT8aN+Ly2y1E31hJrFEHQML9x5b+oizCeKAO
sph678MrbjQ8Exm4KvOv0eJxQq/g8knIqhMITsivyzJqWrJ4xsAjivTtfskCYOHG
/90HJYAIymqbQMa3MhkCn+7DXIDII8mwbRSPfkZKz/BXPQ2+czUugHEpqN7GcX6M
wyt630p6Pl8JmNG/mv0gRZjIOUYdoiEmPx0R80fkcTCgE0cliBKlLITPD5WLj6kp
2jHSO5b7ZBWVyzewenm01D6s2pFexc14cG7kyh8I7IYnZxGAmHuBgzvT8RYaphIL
0rzWnczlxCVTI6+sLurVMsR0C45l1PIVWv4LZW6ULyFrR4Jtk1fSqZstFWBRK7nS
kxX1NIR1837Z56BU9tN/BLygR77P3XFb4n68Xy6P+9mSjgdxlkH67MkWIF4AUzwR
fqqXpXSIqpdqzmnSSfu2PghnpDR6mrI7gEETxaWRODNl6mATbqnYdPHCnj4TsWz6
zgCKeRI+OsVOulT2svEUp63keJodQVs0lb7vQp5xyYyXLCoGCsSX3PedBDGOdRyA
2yv0tmNwb0fLEa4KZF1SUx/xrSgRugtCFKboa/Eoi2Kt7aV6fUSv/wZZ3YPd3bb1
HwVFESjMVRDjr1JLHEylVrnsdywKTjGpME+MRlyKJ0zmgaPBnBzCCin97Er9boqU
DtyGJiX7hSLw8bdWzN0sG9k3zV+KY1dTOw5G23Gaw4XgQQ9+tODfFiPcX0zJ/Uui
ju+HoeQoJGlsbWonXme4Ag0kCgPvR7/LhLetdo7linnyU9LhjyxCu9qaZbCZ7LCx
S/VAFmCanVqnwq6q7ciQuv5IYmlW46dz5Kvd5QyY78SDKZ1OJjrYciUqiqduvCse
Md8cn1B5jMTul4/wHbUpI1vTVgvdJCNAttBwWXzIW79Lma6xCcGan17wl8fRQTSc
cuinTpgoTRjsUhn+OClJ791VtZN5BzofwhEaE3LVIn4bP7VX7iy3C6gaB0tVm5c/
aOh1ojBL/LlTuNLH5YYLdnPDOxldKcghG33DRbEgmfqQGH1s+2qg8RUQvsA5EYwI
zl4+VfflztVBNoupNDr2Ay8NcWuIfKgu4GpfB62oN3lwyUh6Cgm5JPmrRC4fYqau
nTFytiZMIzdV09ByBzD3OyXWNyg/eQCX+/YTslSpiifSAXBKBWpjvSwXrnbYKP+M
Z+CR+4r1t8sxlGOlumXbrLmqbIfu0diwze9S6UlIhzQkrM9QgPe3tBH0nzbxIT61
sOo0aDTwuxVgTX9KVUCNfcO+F77oFzaxve6R3MzqSZ69nCNr7NYmIiD23knwAFE0
XYEmiVKeVF/PJAJGZDinda3h7eJViZwV4q7qZqV0qJv0q76oen8JT9bW0ZVZ8VHo
yZFGawISTg0+JL52XfLf0EgKL0nFz5vnsvi1KYUKHHtjst4SGCi4tYusdbU4psj0
n4HO9V+pxr+b5KzEYUZNV6/quC/nZyi5gKoQVg88SrM9ihv+FLTehQzUJAMPQ8+6
idMV1E79NYzS7gxg16NszvyQsNy3XOuMHbsYT88pXp8J5An7KqBWVgoxrBxypEh1
Za3TazH/Arc/CXNCppYtkgaJgkP9LNWDq+5kwFQ8gMum8QBiB40vhoUxuM4QHLxa
7upgVG3IV1602ljK7rqrwF3JKUTH2vKV8Ku+0n5CNDsb1jKHZyhaQDvZ8JbeUB0A
jU3l9gEPk6kgDeojCg8XKWDyB+W5VcMdLpSJr5aIxxwvRn+NXlpod226UCxdocbk
Ia99RxEEYA0B16Z/lZNRQENYKjcfjJgUoL/zO/xE7XaBMcvv3WCAxmoeLesHEJLP
8VnHyFnR1DviRhqFuQTjbHyvOxoEjTOLzGcUtrCXwt62Obskvg9W2ydwJjeK4hHw
nkj8o9jWmS0pdYd6S41KO6SiDZFFxIrmJTebv5JlRr1Ilbq8XpQSStgv4ozOf2TI
6o/hPqUbyUzsnS4QTrN+OfpTu6qsack0vkGLiTwi8of5qXEoCSVtQ/0HgDTcZwk+
F/lb/MgPTDPeZAa2VAi0UY6P4JFsUH5g6W1rDIhSPOErYIlxgEty6ZqB1wEAppSy
/sg2mcP6jcqgjYZPI3QQCvNAdhQIecxQvZHfzqzv8Y/nFX6L8HkEp9pNXCLhpFNf
d3IalIXOgfKo0EJ3sQpWMdc+5rpHm2v862q8R8bsXUmoCuP9KHH5jpNqn8ufgcnp
Zif/ljCOp9/4qfW9HHqHzQW/Kc2wvV4EpIXSXGgw3kjwC9VHRKXQrxLw2AOQZaug
M3I3UvIojKb6VeFrpE/xM/HGN0dd4lFA3W8GUlI7xD1EIA/S+jwT37rPbg1hfvgn
GbbGPHWVZp+7LFoMR9nSO7l2avu/kHLBKS+74kaC/kMCu7O0VVHhYENFhGHavigI
ds151Gh5+4LdLMEjYJKIzkJk649S6oYWOjIfNVCa4MK708UwJwud7xghjpCCa4Fu
sDohtXsf9dTc8lnHJe3d2GXgwqlshZAIFoOkI3WJcVFC1ZH6cFAeZ6pETGMvLpI7
LzVDXuCwFQaMDNGNUxYchCr6vBwlovdC5NcybMaM1S9F+BrimWD7sdUrvksIL6DV
Eh043vMiZOZIIm3aouRgs6wqW6pSHejqe+DgX1wnEooRcfEb+CaainDdGTQRlZHO
X/hXW+ILtkzNkOwOuamTjETm+QW1lfVcO7z9rVKttdgwzzRgvhI73EkQrLNXxS8T
X7eR5YQyy0tK94DOTIKmYEwV2p7Tu/Il5gZnfpeRZpxqmb+HbMQujZ/oqDW98LDz
vjDuD7UfTT25Eenv8fOgQJ/7WaC5u31yqkbbFg9FTWJzG/WauneFRQhN7e8zoCgf
JvC0TjWijUqFQsFiTlN2YDeTSLWtacqzF+IxphRqeuB/tih8k8HXkFLtHF4sN6M/
WwbQp7owcCvlB7zSA3DuUpVC8AG+BshfAO8kZhqR21liRi3m2gFHX4ihHUaDTHeu
QNJe6bCFlhYzIs31qfNTHyp/4n5V+UuhzjPHH2ZG13Fg3ctBDpvbua/KR11ljmdf
Tw9BkfOr6ITq9r9BBw5fF5GYNp2OgXv8lARgzcl8BHu2TGzefRtL9DUz4EKyE511
9Wkt8S2gfYV60lYBGQ3cmpA31bHdrG5ZieReGiYerPs84r3CH8DTsXn5h3Rhwost
LubVrorUAoGVs6+1kNX4dCFOeoK84zEQ+dtL6cy6wqZO795usswR6YtiMsisXTh3
LbJLazbt+QYDmaAhncFJG/mEB+rXcvQX7FO7vwPNHKhPSYTlYJLQkwZOaKEk9bK9
L1iHomHEM8ciWnSJwFBVOe7bKgDkTLpyDqIA1zMDCsbk1h2NP1ACgmvDOTfJ2iPL
+8CYrExelcqEo+3yA0VD27uUXHl01poAoMoOlDWkxYV5Tg1/5kqm3egsJtr2U+pe
eIypqVZAE0AZVOCjZSepIoYVW2M6SThNUAAZ8ui+1tkSFqDlkHpJc9lUQMBEVGqT
pANbpAFT/2RGmnZaoKsFQ4jxcB4zTXsLQ8HLko3cuQZtfM4ZzI4MzbF/9arhD9p4
bfx/wetqCh2JYe4zLlrAI0qEb4ahe5+VdQP/8TzRzodwqbuWjQ0nK0oLFrpoV1V9
jMmCvoRoMrI0hfLG/S2wNHNIgKXsWdcJhVhVliHr0hAbcWBxwz1EXA5KUnji214j
/IWw/XzWQzH56OYEoMuHtAmZuqFhcHbi5VrT0JsklttnjPu3Xu6CeaVyRVjaQ3Va
UwbHZUuFqR7wTbPha72ypOYzf6aU7d/cHPuiZ2w1VsI5QPGVyIOWzheXO7pBbxer
Jpcn7v4qk6ngeY6GwpAaABTIXcusTCnGXiwB6MJdfhsTYQvMAIiCMoebNG2EVNli
ACd96rThpkx/XyM/qNTe5Ld5aXygxSb0pTxauWdMOfdfe5602KIM/OGsC8m3mcil
raNKfAqx4IBH7subsFYXrJ+kz7mF9rELftcwHp1d4e3E8CLLKj1pBwSxTaTTcO0W
MchYgtgLW8NuMryuDFHRL0t4ARhusVtlgqRtw+MvAdnodoJP55z8uUwPOkqn2xDq
9b0y3bw5JWDnmSKiWxdB1kaeEiSaoRzskzBJdN6Rhdxc9M2HGbwsPnw2PfzNAvvG
NuP3kvIZdLcTP9Y7546v9Hxg0YPcjbjZAhNRLOSuXUS5DJpG65FbopPC0/KrU+dP
i/SMebSIZxas2wZeEbFXR1WA2IrklAD6Y4BxiPNjFtzTiTGoYyqpmcNtFbV53g9e
NdRmXIl4r4GtoEJXs55Y9doxvy5EbByIBJbXWc6w5XDSqeBbAtiJ9/02ZC/+jMM4
mMCbfkv4nc7nK299zcgsXLawogZoxtk0YsCk01GiXVjq/DUlCMZa8JKMc8GE5COi
ZzuD7+T6AYI/8qUULDB0CVT/hSA9mkvztX8/yt5zCRrldmsS2vydudQehu8NkVYL
r2JSQJxcfB+jpYu3QlH7dbRxu9ORUbuid01RN3+K+QyhCq2J8EOfK6pEpvq2dMml
geWEjR+G1eVDMjnGmPYlpDtMwIDYx7VCR8p8okkNG93HfBx2/aYsXWDq0sJH04Dr
w54PnoWRKcPFzANhOGEMvo0w+kP9Zg0irfRyx4qoI4h/mkyJfhwrg6YvazWt1rnl
vvruVcd11RcuWAEYl+vYmOvCgmnwD1/VMFAh1Dq9Ja8Qq6gSr/5fSYxm/xYg+O8P
ucSyKo+Iy4liUun6bg5UoHPjiqfgp0fOAJwOzX04AWeFlWzbaUGLXv/itb26FTxV
nNBuhmkvsTQBcZ9gvGUfpguph5VuMxqwoEN1BPf0hzL7E2g3BgZvkZSZvG8tPosB
+VOtc4IIAIaQR1usXPeBRD2k3QzM6WqdZMemPKwgkOslnA6uUbXp6aSJUmEx6qnQ
cWKNKbv+N412OT+yuF7DPedm4O5aX8JfTE9k+CYYlqIjzR6y1ljumViRmyLPRXAG
GFBDC4YekPpddmDdutj3sSjuQHzsUljDbDmVqSk1Bjqf7sG09Y8qPHSQrXYn0MpL
riFbnj51cL972D63mSMlgnwwe1pkgbVPYapb+oyPwprkIv+lpwszWSJGCpdVUw3l
Pj62hi8UQaSNh9r7LSgQBXb9qDih7Do+1cTmK1cYyveLPDZgpyENVtVT768/w93V
U6owbSBHqGWLY3WaglcVFddbtEqs5n11LMP/50ZwCaQGH0O/YGChl4aJfcw8PpWs
dV7qfWBDmeDPs8X5o8APmPdkIr9L6Mg01I94BrIK7L+UkiMlgHVfE6Ak2aYAJyjq
3RGKO7Ny8YlvfYz/AC7me1giGjHKKLL7brp3u6UDlTHT2OAQisERvNMf227jFDtN
Glmewhp82j8vZHKpzsMRSeg1u5cJ71+BOUzWtXNG9y0hTEx3umVr8vxgmRMY4/UC
hoylrzpQ/PXN/nyf1GaORKyIC1DQKIKI49gYgmqCpHzUCyJYWZ1b9G4eatVGqhc9
IUbgtqsUjujgF2LPbXtMhh7FVQe5TWnpra8QwGz2+NSD+RNWOWs5Al1SdY3iFrH3
hKfYaJwNVogqdwXPc2TGfqVpMdcuOzwwKx1HJ79UrKaIgRUgtgFIzBh+fgJ/e6py
FiUXVALxB5LtrWBPAXZyXTUeMZegtNvpNPadlxf3EfIM1ExYik350s4EqQjx/Ej/
fhcyB/qOi1+ebcFMQMtifKwh4HEhEkpMidLNkbxgItJr1hKvTDdOv/ej//IjLqMJ
Rs8rETWvXEUvhsn9MjUdn2ctV3ZgRYsBnwex0KyPw42x3EsmamJidGEVRegLvwR0
DR73NkTeAo31kbYgsKJtKej6A9WIK4GRuW1zUM/5yHLrJ3UwgmGvRxBQ9whQjF3f
8manCLpHQrrfFDCTr1UTthDXVnQzXBe3VK0vaUgIjQ7PMKRtnS+nMOoqOJNiYx+6
56CdOF+EjwkltgPHLy3aO1awg1IS095T3NjcT2225NaMS0GSzGO78UecmjbAZjm3
Sx+vCeHsG8J428zaiQJuFkvf4lETGcrpK7FsmMZSpspLvf4WYm1X/8i2URX2JIc7
Yw0ETJ8iklvZxGiB7O56AX9C2a5WLzqxBfJ+2/cdo8N4bpdCj9dnM9JSFjpj4okf
NDMgDAxaYAM7pVOjunckG1Yj5yjSmlFR0nZOFlN/g3WAo5oACQD7ibT/oWoqp5l0
1kglLA05eoRPXNeYQI5bQ0N/zEdf2RXLEEQKdF4hKcJivIDS5/yd7maW6n62628N
l862X5KUsaOrcTCGPpYSAQToE2gJoYPr1mNOnRHwq39V2u2wneqn/WRtiDoVR5Mm
vdr/VEYok9P1QhZb2BHm+lAk4QC6cFY04v1vxE/KWGgCHg+rDnnzKlGb/0DjuITf
R497tg1iM8x5z4NWLZgoCU3iiEWdLpWp2xaLpyTlkHjhUf6FlpqFW3RksOiHbyty
uZ1cYyh3VRp8OYVYr1QyWrgBuJ5038hBFp/m+H57mBOSOvG0JghlTVF4FRO+Amsm
HY5nhn5gedjNK6em2BlnH1OFVXAA0FyyRo4lQD+vF4s8iMoLL0xnGkHfHxKBdihe
wn3fRKcrRfrHA+yFDKAoOJIY8gzDlixDphVwBGlF2aV+hiw8kjJXNY+H1MQ4gAsy
SmKgtRMK+H+J+MB3WkkzwWXQgXFu6miSKVC8R0Y7LiWfhE4q1SSsZUjvBVMbGfeA
BySmn6aRaZvUhPY+emUU4LAc7xguUjVEs3ZgfJTIDwcd+cqsFundGQO7//vbS/0n
XnUh5aL17/H6tNzR8VUSCZ4t40SWYNGQDBhsofE+8+YccqZMfYPb68Qd8t326Glz
xA6en4XJVueFJdayNiHqnkpDBCIg3iujt60/k8G5x7QDusMGCIcp/bSV8ro+/aS5
RtqUFyPNmN5/ILFke8VybEvha96XOGYVS2984l8cUgQm02GOBPOnnM3fbU1ZCLJ8
WD004ATpQNjW+Syu7bced1tlUryBJn7E9GUs4Zjq4PGdgMkwkBxKKwzc0+q1B7Ac
AB4d8knh+YWFk5+k8spZIg3XszAggc1s0lYrtdgCCI+D/KYpxNIMMpx6GAJdYX5o
R8K8gXPQIEUTEvEzrq8ik9KNB02n5jcHgBQJnXDjUAleqWNYXI01X1dpL2AXJEmI
IpMenm8uzqZxEX9QTff0k9I7bl5ERw7JO5GEbEGUEHcGkuk09cq5Ntbee41zB4BI
7wKSOn/BSZsLEVeMp5MycPt+Z5qFsdZchEmUsqQICUsw2CQwxuhyGUjmE4U9au6I
BHldM7oP1gI32UBLJOOjQ0jr9aHIueZmVODtBz9sgx8keWYAxyBX02pMt3EQ1owb
eoSJvWSrMI0Xy//3Pnvqv/g4+0Ti1aUnxnLv0ggEy4NI3IQhV0VVrwdnLJ8GJ8FD
fsT7Np/9I3BmENQjQiKcnfd5J5VFABOjQnvLd9dExonoRKQWmqI8V/NGj3o+appl
B0or0SkS5ji3vsLKk8EUTwVTnouk50a6QuFpdtinoAo5Z8g20moGA6cVX2rCXn59
k7PypYWgxQ/wdFTyt769QirxKc9C6iNB6HhXtkcNGn2elTEvDuYVxSUkgzdX6d1o
PVh6TodL9y8PxapLUenXyLVDcfinEmbCqiRa8mHAwP9ujKWVAXTH6+uSLd4Syoda
YDrHwknxSgWpgf00D7NgSrDc4em0goh0009i69yiB7+MGlxFIpAK8Gflhq6BaHMl
0WCo5XXz/eB7NEDdViWqG2XYbSEgTRG/V+rk/CPeI3oObGxVkak3gqxh1kvohuzM
x0mcbCKtw5P73nLrCDcxHBNA3Krmpfol5tb+Bor6jLu7wxCbadukYnB2YN6QFuMR
QcS2voJDO5bqozX+ZhN2+P9kQP3hYcCTnHlcfA3y1N3nMSPZXaQePg5K+izWNoXS
xZMDAoU8PltWwnN4ws4LqAWmRlHDystxJjlqwYTXmyd1HCj1inmR/tjLrTwB5QBQ
RYblv2qrSKqBxAEnUSqXKIe825RQPQksi/43sdCXOsxSpvcefveJtOuiMjVZRboA
s42EjTTuNn9hjsEgF3IHBiUiUd3GjL6JfZfctOols7d20OAc5XsSJ+U7dl39qBmg
244inx8hGa16kDv86wR2CCV8oIFxbb2NMEq76EkCdioXCDT9vIlAdvPLOcWAPFd7
40plcmytG50ltYpCQo0RQxBvu1G3e7HERBJyBdnlxBJpDlnHi5hIPnwMRNQK/eYZ
rM6j+UjdvgMvsOzt43GTqJIKI0zW+Z1zbXgyWGqfNB45wsr82dZE9ZoXEdlj1BJW
GDqE3bDRIKa+nq/RLMTMrM7NC2CduBp5rRKJzquL4HYRmA8GZIdirZgYLYrQGlyK
Th0vlA4UxwUVNC7auASHQ5eXfKhVQRRvc4kOMI6/rv67MXDbJIwhjysWMY4yNph5
wXmlEIiKaJC5uon41YFvSqCCjah9EXLS3TmSB0greWl03HcpAqaPKxHVk2EUjQE6
24GW+khHn4s7nFH/Z0WBWrrsrMrwbIc778GG6uc+AYHZEHU0Rt1w5eveiR/Cd7hu
blF9EKECTLKLmuy2AbM9FEVSD02T8fYy5jX+tjBG9roBosFFpHW/gUJnD3/g8YBi
ReGIYMwpk1yLTRQVWooSjivrrba4qQ5q6YBzMhA7PMZE8k13A51Fl43dEvhn0oLW
k73tVeZDoabmMe9F/3sigIC4CxHdLteZ4cETnp6L9QgjaCYqTrkZPUNXIIfyAPKR
lRzs27oLn6jhxnJDq3VS895Jv0sO7PDlwNkche/TPZIai9cZd2pV8lwDF0z9HSJX
5N1x5gwAA2pRblzAsqpWV55wxHCIl+hz54/ZqPi5WNiCUrDQonwAB3mPHl63YmKi
2f4HBN6jse0zhzW9MCLXz4mhO1mthMZZu8JbS9OVeLWoDN9/mfe3AYZ/X65adaFY
BvGX2CYV5xCk9BpjW4vDFYB2jsB+YwwTGnRSl1nm5A8BJCpgs206c8jEllOW41T5
XEhBODlklUe+5fs6lVKjtLMYjCCsZkqLMdi/ePQe9oa5/pqufhBdiTipFuaTDkGX
TDxtuB9jKomEmHxsBlfId+NNYpjWFzevP022+yUbW57Q2xncP6ChfqvRueuwxkjb
jqnJ8i1Oyr5B5YJPcBeL267TuTNQIg1eyiHlrQyHUKcEh+nTDOnYi0kcUzxrJMcz
hHdGXSdfQvdyGuTKSqn50Tn+I4RImJJ173ej1tkRpCy/cJE0L8xJPcl1ra5eBvDn
r6grKlbXYaLCwq6D6sRsNJ6J4piKP7PSO2YblFNW/yYuX8SvxTPdEGYNr1f9Kog2
ZbCNktW45XbfotZu1YjKUK3GIlqNcKmZ0njdw48Kb0xOW1R9jE4ZulDNNipH/7XN
ANTw6HRt50EkeRez2QQXO3yDWoBCrfUdLELdwhIIHgSwnT7wLT4cU2/GtJ+CG0Ye
P1wrZX/L5MuH3o91BW2LsbYLTTyph1fzwVw9yTE4z310NWf/U4wuxLBQA7gpkDER
haR7e6igxSySyGDG1X5DBQDxRP2C3oCD71ODBNhKmWvvB6ni89dZI5Zb2cL3txJY
xtEmFML5fw0wZUvd1zi85uqS+M0dz94B/LSlvPdUnbbZszUm43lSJREs/sPvdM6Q
KZH56T5kqQrMSWfL3Uz/BPG92Bnvm0uEUzk85MlMEqmiTvYJ4WdJzluwazWZbKnz
BekDuTBSwicJAdhjPbQdIGu7en8sG0bsIUnY8E5lnWV2zDA0tq1AZsyMSL08Q4/c
/2cIobXzR1CSh588xwPPnz5Fi+fQjxFFZEggOevDnUer+l1B9JdbPMUBEPHf9UK2
mXyltnuS5bcqyiHutmnq3eZzxVTWkXjVjg1gWWIRREUmbDpjBCXLsNqWpOKdSRjf
+Uezhux0rXoxoCsZ3coMBcke9E4Ars/AkWwdSPwZe9OiITrcaes3e2RgNMiHuz+g
O3TUSyY5JNfE55pw4RwDHSeR7Eb5H2mGdBNHu4dTHGznWQVANhmUi33BKcY4wluk
1NBdoC+WKea5DRlStPavgQRIHWg/hn7pfqta1WtS1TKemLV1wapM80IUsD9yx7ed
xqi0hmrSPwQFHX2Lmez19Y6ZFp8C3gVmGEM3VBwn7FBtiQqrzCEWNPa2V+cqpoN+
N4nqyAsGjcfsQcpNIGHIoCxv0oQM/LU64a4FUgwFW+tHNn8g7RdtXQ2KkVCCcgMp
ammr+aqa+cnPtw2di7bpx0u7V6kleUSsGBrgjNzVLPvrXrG4rhsTv1cD2LbmHfci
0CkNUCxBG3+5VJ/wE0jfLBMCpOKMDXfeJPu+/VGfKziwhm4WkFqG3byaBLiYowgQ
LZxMffrOaEEfo9fuX7vGan79OplFQnJ/lXWY6Ge51Xm1yomKvAGV0RqKljhDFvY4
bIGuUdJjfg1poy7JSKmiSWLp1hHH4UMHgNwoFZgZVb1tY6jB8XQuwW4fa0GwVLSL
qaBvHrd0kFrwV63dUSmIck7pWFGQ32tCbtuEaxFRrpAVt30TQx0SNQB7RKRzHHjB
EI+W07J6KoBH86wDFi2LtO/gyV33Z3zat7fE0rxbQzKBk4dXUVWse5GNy22KEzoM
4DijeLv5KoMKFWfydGpptuG1ksbVMWuoC9vITc3lBotxBaZ1+aA9rnt8URXBlq+0
og/yI9TSa2KPbfdYviruMAeLL5fcn/F/FSE8VOuU/qZ6VjB1V7m8e3hwzm7XT7ek
Voxuh+EmaqjaQ0xAE8gAGx1arogsKy4sQOI3/0ihwTMVkJ9qmx4GZDq+aLszJdXa
BtzxBJdlcAnqA7yzsT82hoqL5+1hD/PpwpWGobzHqBUqVeblKwjcQT4xc4IQf8Bo
l033enwtyix6fLTQ1VNjxk26Slr+t/CobKquJDZnSwOliJnySXAmVr6JhvWSSeGw
NsRJqFfM189vtaLppqj6dt2fAxdlbH7kv2d8U6NWKTP9k/xeGoFofw/2NHebGmYd
trIGquYvl2iYqwB1lfjVZYuQG1LNTV5NkalWZ8q9FCChUapmpbhrsOo+bAxCajdM
yuhLoram+ebTwdn6q2nLSDwgHljC+KGSPjO9N8tRFDFBkRfb5D/q5o9nJe6Fozts
x1PXsp/j1CMfhtSVTawxVbS2OubYctROG0c0M2Q3eU/U2+Gn4aFdyiuF9Om0aYQX
OhE/JWB7NVK9RTC013HocEE5mTyAkg2n7I91b5PyVXJrckwDnQQwBQQeGmRSJaLH
92aDj5jVSi9lXhWiayNSrupDO6Rctxetcyh6iDtyMe/Ca5h9s+4gzy9l1wc7O2je
4cng2DDGOnZuYVTdQhMoJpAze3+25HAxUcLA3aq5c617PbN+91o6MHz6tWYaP1oQ
+OBBQLnoiTrrY2kqlV8w78VjpxN/CArNwtXnplTy7d9myWJLx/+qVseQYBaeNS3f
1Y4GOSjbyShpG1lYby+51D/+9dFvpIXyVHRxCDmpCniYdY6Q5Knu59rjuSPggSiU
/V6q9cd3+79TLwqNsuZBL/zavq6meTVyvQ82BwsGDMJxlLbgJfo1WrrITY7kAMic
VmKgOUiigsJrBYVG77WH4siqPNsv5OaiRt1D9/LFBjpR+6a/aJhuaxjW31FyowHL
AwIUvqX8k57MrmjO2sGwZ1hAiWC6qhISFJKS2LUW9EKlPqf6Q1g35xQyeP3R8lvh
zRgY7QLulsYJR56Hnpi5mnMuVTgGBAI/psaiKERKkoBxy7wvXSIj+NbQBVkgLCuT
CtUsbzE0vQR7gf9/cBKqiDz3UK1Q0uJReoP0A0ea8VLF/AJr+K6KVt+F7up8YR/h
60dPAsFtkE4MsATZ8Sex+FM25B/RG9pq1vZQHVg20BdU1WI0k0LMJ9ad/bMPjhYB
0r5bLqisv4meLmxFAvn58zHFrH1ujw5VUuRpNz57c6qgXx1WD1BEmifIfDPsXwnR
Wh10I+ipU0TJkYZG/qM/2LDUb/G6pY5RXNxoHHPn7eM8wEQZUHSkmhT9ECUG7Ilm
Ml0bv9s5PfbLcMbt8UZ6Ta7a2ezbo6f0cGY4Bn402GZvLPBtIT+f81nVgVT2cp9F
PVLW9RDyzfYWopWIwmkTq3kIK5z8BO38qz8v57KcxlRiZIb0JFusVF6nupwBiI6p
4Dpu/oihReOdxndTqCKHe+NQ88lQ9VT6+1fTK248fxzLbvM+3JGiXfuNUgGOzyL2
v4W2A59oui4iFRCy3KzWKzN2XT0nqyszKIEbLuD69NlkqDK1KVvuyAlPRAuFSaVl
fLoVgFpN5aoFjm2ebQfzj390O2tH1ZoykmsjS/EzgWGkyc+CWro0gcfkwefKmdUK
yT4oJraNcWTFwUtDQrsyLG2YaEWZZHIHotJltmhVGaKstidpY4CJd9BoIBSX+CYF
zJFuA5MMaMaOMVFNpKCWpaHlt1XyW8P9g/0Jj3k4GZsFoeUbtbKO0GJSXjoUrJXi
Q1jAR5eIPcOJSzffQrWfZxjAHx0uG4llztB83esVlB/9s4wkEHYy7HSW/QjDwPW+
+4q8y0w3RpE42/akOMEjXGVKZoiRFkFyIp6K27JWVzbMp+h0SaqtUBcrj/3m7X/J
nzuZ0v2Z4x8S68WLLNudbeEj8bT/M2VFBOtskSVNea2YrZldMB9oLNsnUdjiQXbP
fCz8haF54a4RzVIbdQc/KdYU3TVWEtGs+KVT+OD6ewjj0sH4y6Q0fCT87vBoG9fI
QLyIf3BntDfiqQQkOaHD9lhy4WiHgVgRs/ysntPcXAY7SsvndItjKp+SXGj9nQp/
QqsRTx0+HlNuiHimuU4Rd3yx0a7wMzxZ3X4IYurHbKI+jiopHjxgmMSBn/DuFLi2
3gMhp0fGN2xVjlDdzX83SMdxSmcCssyhPMcxmqViBS4NcCsIh4kRm7XjUgMFCGQT
I7fp+8tToHXE+743s/Q41xTGtlg9GOIP3BtuIWodCUk0yiqVItCn8AZTt1I6ML1e
sGJwdHRSKfQZsP7HRNJb5fk2KfezOMMNcBColmd1NLi33vqqgImNfguuMAOS6dir
ZOoXX0QgM2aoVGuA+tQf0VGyxrE/g9dT66siqbra89CwntN79Di1oqOESPw8b9CD
muCytK/9eThjc4Bxy2IZz6scekR/P8F17jFGm30l5H21K2fCb9DnRMROn3k3sF7M
Mp+0GqPyKSJx8V+qLtSrtacGn3AbOFsieQOlyeXYCQetLtVdSXMcjs1hG/liVCSA
34hBbT8Eb0MrvPqt7uUelaMggGGBZKhT8xZlHyXBXej3/ZjTXiPK2WOlB+oJgYIK
gsXh4aSJOn7D4FAjkjcrqe8Oz/2m2bKu0rWDzw7oLF8aQyNqgHjCA2p/DT6GlwB+
VWqZ3RrwwXnpa46lF2JnLDQSaAwxfH5Sr07QFpsl/L1eD8QxePF/HgJl0YeLNkFB
xcqcgQuV+5Ta5cNN9G3TBMaDiQFDNVQecrG6kyh59WK+PVjrgcnIvwtOmG+ba16O
EYO7sqGggmfGr63amox6OLJfjdmvIDAErRs9kOQfRVxKj8yh7in+OWMLBcFBID1R
xg59b1Ybb+VK7MWWZ9tbPu2zRTOpFuWnpqsu3tZy9+wwhxaGeVOFevUy1WiPecoW
aP+boolhzPj2epoiDvYYrGYBNJDIaNF6p6w0v9DB0/SxXwOEDyKWS72Z5jgbq7O0
cdGq84aflya17OQCGcHScGhykm5SRdK/pEod9HoIC21aJ9HSbfUpblS2KHYASRX9
Y6Dzl0bC3IiPfryd5+ev5Q8pH2HPPLelVYX1/h7ISiHv8doL6VG0EWC4wUFm82Qc
sGK3D0ou4C/6qSqqV5R6dfXHuXPg2X/TPTAY4ZBFSuUU0IMR9skHaSNe78ffpSo2
bYnRrIfhQLXti3XnNr2orGxnD04SEbAkOkLT4u/XJPrIud4tELZh9rQH4xyYDZtB
ulbM+ISfaK8COtII4XlMMMoTSnOTwy7J5oVs76kQ+y9hQK53BAh/c4kgAlJMRdUY
0XijfV+kknipyYQPJffzGuzbUi72PjlhdE1sax6lQFaOppkJAdNI4IJOUIrM7Rh6
DHcsFO957NGzeSdgBuYG+ivNkQOE1p/GZIsduVEzjy4FfVbZ5SSQvhfAI9edxMtG
JK+8NEzkSusoHZc7jZvlUbzhiY7NsYvUle3dkvoff5xYIAiWOmH2FE1KbBqAameK
yiGZZIDb8p4U7/HXw00ha46lEf4OYyTgOwbuZuOkFyZIT3WQaUbj9R8z3rSPhXuh
mI8wOA048H1MF3ZJnGy0t2WmTaivX/ACsoLzi56qs4piMi5uY+RACAV/VAxFqtS3
usTkmjx/XIxvI4RhBBw394uyW09ITlNtvLBQKoa2slXn3yNGDS5RmEQz+yJEj3Sa
CiTfK5Nt0VCDhX0G4EMxsJpuSqExHFn1csK2wFm4E7C3/GzG63zUymItIggrNiIS
pf7pFLrnxGVqwETBNCZcLZRxhbV4FRgUjfdx1YvALEaY/gqdkU2Foa5IEktK1CVI
HmF3f3GVFkQWApa8GXNqR/mazTt9ZlOEMO+eAM5Ciz0nldvcnAhZDwk6NBS4EjWq
+jq6ZbnHG3gYctYyN9Y3BPMNkKUYImKbNSDHRu7Nm8IvZbTTLu2F9b3DsM0O0Wh6
XWXuKfq7oZCSvOpJf87t4jfex5jdlJ9dETDEGGSuivL9To87wZm2PL7r2Ko1KSAi
cORfGVhuPDVj5fVOFcImufJ4KEtt715QSlQaRvXR8B9sKaFhHn8iAayvZo2GCMTZ
v1GZhpEQnyfgDUK6KwvKT9sk99VHe1tiZxysPKZcJ/PvFogD8r9VqOBzv0Eb3i+E
NotRKQOAe+wH2I/4gJn8vwqo0BHcFLtsekd2g8wYmfsMRjsQ2CUwtHNiuTSdG6b+
eytFqwhvRVYB1krUQXHBof5KjJUCE7VogmsPyPUKz5TXqaQnAq04giEIQ24sI30O
pIMrb2FIzUzQMVbOvybf2XlfU92U1QrfGJrSiD/a4BknzC9xrr29JWIqp9cqfJyF
KGCaniWRhvlu53ZWSvxSPuOvSQrCZ7DuzPgAmMpxLvmtTebjgpwWv6yWedhx/M7l
iLWsjBv7Va/fxSKIdiqWkg9s1KsviNj6LnxG6+65AOcYrPKQejACqAT9lA4Hi46f
pj/Ab+pzPb7csoDPNKHTxKGJWD2bvEzdCaoIww1A+f7wPKIGyaeFnL2Luisi7zWo
1JBwtm+cdeP2RYnCktiY4QeNzI373K87SzqaPnepdu4RYc2+EStweSFFtvYXvAvH
JxznCwZaccLMl014vlo7dSIo2riCIHrDA3+OLQES/CdL9DuLdXkTj2DCTDw4zlqy
ZkydEtPS2VaAboX3RoyZxzAByGcmpRGqmbhSP1JqaGba8/jM5n/HfccjPFlasUjC
7Df9kh23xWSrs19mFz3uf4pP20PutsC/+O1Anz2puPow2l8NyMnIBwErgLZYDcsj
ERFo0V2aCRf+ezalFk6qiVrxKa7VcaIpOjBmnrAcWDZ82D6Qfm2EZFE/aEOxs1Pq
RbvRn1ezTlMCKzUhghiinT0FezZVhHb1Lt2tIeU/Qm1uQjwikRCg/q8OytlFRRsd
ItEIxBF1yhgt2JBITHvhlP221DtDX4Mf1JOiT4x7912RaeymUna/jW8Sl7MlKfRo
V4gT32rHjZHlAbXz83T4u1fHvr0fjd1mN8350/oP1hg9+Jq+3rSp1xJCGmSRa60h
cogwJktaMSPiZ8OuODXu5DnKHa1DSlRLX51UDWWfe3kbWE7JO3x0VBVw+X9iaRYa
d4cMJJe0eyfn0jSdcgumvuB9xiW7bnU+shvVEjSVa/d2OELTFwhLf92bMLoTPw+V
q32Im1OvOwQ8arvQ1sKWogDRGhG1v35B8w+smmBOIwawlZXxsJ+M960URk8qo6Dg
JJhjPjdOs3LPPSmuWM4JvvkvVqpsrlHrO0IDa6dk3MwJ7lgNYGutY29a2z2O5EtD
GbvtrjjpgLhyayjj4lXgsSOjAXOa6FSljFXoexvd5YdbnMmMNH65BLzkG9cGVj4s
ukkE9NMO5A9Lg54n4FLsV1jkVZ4KJBI11Qfl8vkg44me3x6Hz+0OVGiwBeoz3qOh
ZgAgRrin3QIA/CbWYQ9Riu3qvaoPNU+kAJeDxblToxPLZgoMRhdfv5GSQuiokzzj
5cz3VXDJF7s3kDJHkYJXPpX0GzSFfUUV4VoxPCxZLUe4HJgIxZFMi2zmdjVJ53hs
JimGsduc96osnlIvUjx+neFbCA3KMXEkrpH2TW3L9sf2JuF1Do3+Wj0KpFrZ8Lfy
tgwax9VS/u8ihlRQkWQL18xCnbWHlEnBgZtzpbbBH3lYKxWQKhZDrxwX9t48mGII
FO3GjK7L+mFSvPO/Omth4LCSPr9b2GG/W7YwLfwVDAAA05jaWg8i5hWPmatQhaf8
Gqmci7edleX/zwsC6bR7rbrxJTOFcE4PKSwrpbs8O3ofUke2EOPRz8pP6dyfq1Hy
t/G28RxjLru2bPXWD3Z/3R5Dl6J14SbZ2ayHYXSD16qoKddHXEnO3tCPsUV4R3oj
sGB3MgxvQz8dHMpR/OsT3Z3s8El1rYZ4QX+oJZCa5gKpCRz8VsW7jbFVDoB3yq0n
8cgABNRLwm1bhbZO3GHH6TM7bAhgYC7h3OW8nqfaZgI6dJeKJPz1HrfUEl7Beyom
eKcjHsvpIv+Y7NYzvCOqK/niCAIFtB4lO3Azzk89ZtCAH0Xw1pKG1cLoxhLA+Dqx
tXcWDEPZWJ4+uAsx2A1uiPsgs55ctEtTJkjS+12I0iAeTJXrZ5S8dX99BjqePoaQ
CGyWXwv29wTnGZi3jB0N5JjZe0o4R/LZutBz6jXFkl6x2yRspk1Vx+Gmni0xkQeE
rcEYLuCdCJq2fgv/cgVitUz+k5lRf5qS3TcfTYsR0p2/XUZpZvY/QYNLFXdL2zO4
dVECCVtWt7I8jzhPQEIoEQpQ48xmA8ETS9VyJNXO+TpL2WnTWgU0z2PTedmc/CCn
pzMJqPelkgAsBh3VbQd959U7vEGgX/8oKOWDWl21sI7wR+Uexq/uKTgB5X8180SD
RwKzhlT0kTOK+xZ8+4WdhayGEXlDQvCweK9Quq13CfIRP93fL+tQAzxWONvrGoWg
rQ5Rvi4E/Uj+AjgTsOVBptZ6P1VFlcVj6kGUTGKhv+7j8S0e3qE0wWzbVQq/jqKd
KEmENILkgpfnxh5TKZu4m4n4G0N9z6+GVRYk98QHJ1xY6dUux0kW8E6XjUEKduoy
1AOfIX3S45hBBo4CWIk8ZSdm8v2ppH6xyUUsCveyD+f7yyajF/AMyP+2aq3AbsEA
RjHNmIGq8RhLbFsr8kAozsSJfsQmIDCOemECkryb3lvo6nt4cLAkGmvVs6Ng2I3y
4D7CoC9C8RfzcKnQvNd40yZtTvX94/frgSz8bws6PNvOwTnxjJZY2NM6q2kQiXoN
dNjf1T7H9gLEfpYhu8yyjErtJ9JaZA6tAhbSItCuEGKXEaOsVY1CpkYGyUuxOZg9
hZR6rnKqrel5krPsgSzgSwMyY7FwruFM2b/9Pf3CeIk1JwWHrdyGH7niN6GWAV8B
ZOvuDMJ1FqGUrLhjDqG7Ft1g06Rj2O7qPRQ1X3ALjSgsUifdTEj2RPUUN1fXRNnY
BKfXE7U4IoFqkNICNi8eA2cvNOfmtfyWifR7T/J8SndHobt19GskgGWNrZaUnPTj
BAuBBVaNQYHwSEZMssKvyArERG2f+d4IQDbEeJNtLEJUBnjvGrXaNA9zPRJQOGs7
Qcbjl9QNTMglYMHaabDNk++4BN49BxwPuiVv/JufDhCBkKlRGIRYwB63WKzETK/m
HpicHEmBS28cbN0jeuvvT0daFS/CfvaLVA5hv77ZQtpecRLnmZggLTe0SY6qNdO7
QBALtKQsp+6RPtiopAj2k8wsjkM2yVP4r7bUyBoOG7txEVYjko/dIAomQaV3oOOd
He6SCrznFmNhz16gM2aV5+ZWNY5Qf5qi6fY0U/QzzhhDy7mxyBVquk2DxHtmREQX
B9IMBKyYJxhFkSY6MWZKrlo7VYOfeb/a8KM36z4S0rtnbUXydZ+2kxcxEJNWiqTa
G8SpgLLilq4Fw4gtJwWLasTsCihhkma7EhxboGLUQwSS3Jh9iCosy53OpL8yXSJN
jTTCIsqGw4v9RkYVMHToj5DDakZ1Y6cIwclLEJkG3ZX3OENKDjm9viADwaAYJtHS
kbYxsXuKy92aX8WHh1psuD5E594so6uNaqu0woslvi0n8SM7D9dRiW4AKheMSfam
F3BDQ9vYtUJeIThHSTXJ2RTP5BT36U8m9zaqr1TPSD0PMyZspPgmWfdAd39TzALK
c71qsZ4KzRdiutmbsbJYIy4coD7LPG+KxXatNN16gM8zKUqm/lTbfCiqDjjt/iyi
kUf0cykAxwCKyTqay9r96gORqJcYdfQTd9XNokfC6kg4xWpe6K4yb0IrbNs7tuW7
vC/l6dNWuAt+P2QJdoVs17oyL8lviNuHk/6GrXTifb75TF7nwSQDewsX1+BuHh60
saqPjtAIozFfDog/xJ3dIaadzQhO6uBrRlxOk9akHHOtq3fa4dpo9VEK2Zz1ymnR
OYjj4Lcwkex2asubZ4MYplUCIVWC++2yxJehPD044fufhDKxuZdREj8219ErS04o
OTDJCqGu3U94FpxhHsAV0x02nhAfGerEsqcfppCaB+rJ9i0cB0MLg+LsfcvC5OGT
m9ENDS/IQIhXDriP1IlPiKPIPXnj4r6ado5qhXHfvN0lHt0qctNYyZkYIWZznqH+
JvR6x14UXRVzd6KSNjhTw/qIz/BWwYORCYHY2j2znp3FKwR+H35aD8SkOtDzLLxZ
CfrjiMXqfEHgVOrHZMohAX/XmiCvKm8ZNZ877GttN47LmJ5Sz7hPFlM+IyWMeZC3
+89CNt2ofiK89e9fUGe7J8nfKIY6qplhz2esBcV4OZ/kz8bkOINCHvx+LvkviSYI
Kq8YoLmUdbmSNQpZnRb2PQQX0QmQtBhCUo3bpCxlbS+Uv0K0QbjUeI+WNF+stRgn
XQuAU38nzkE44ebGae3rL+zW7cMEzDlPC0mcwuD9eLMwz5WS/EzzvbAtBnL2weN8
mCA6Yo3o+zl/FVSmQGeG+so19hL9rrqjg5B/TssgGDPi7bB90tHHMVoAloQPCySX
eua0Wtn+pDdVsXIm4dBZAXSFjK7BB8kcwkU1ZziVs9+gCrHNHSNU4RirDUx2SNWN
QjxnipQQzN+lE6413ozGtivdKpPWbn2GbP2eRiamrKu427p8LF5NgeCydU3RPoSi
bpDAeyGU2zYO9KkmNKPA/I2yJgbQN9etGzIx3kXUz4Vn0lHpWHDgV6aaHkxDgO79
xHFEeyYDj8JaAXtZge6fLJedeAdiS01rMu+1Nhtbxo7Jp21SdnvzRHBkhRm+72vp
vOWgry2KlX2mVyIDzcZc7Lj6TFJgHXO05NjMgvFpunWrICtohxKbsRjSbvyk0ZZf
5icvp4qLr7M3nvqgtADeJpurRvlzhytC5bVDoilfU+JqT1IHjjTN6lrX4JdpjuJo
EZRN5H6TiIGcv8WBSwxjyXVpLSMwKbr/zHqCztOQjbMVWrkOG26MilFbQIuisQ+d
ea4sZEdWbXJIZgkrxfuV2kxvnbGtAIMhbPmaOEngEV9CRJ4nFpR/aQuRS2mgYjh1
s/6SrzFTqh3k5a8Q01rfxFJ/SNLF4OFcBTfKITYvkXcE/1KIwriX/VqaBIK8Pg55
UBqj0phGmNZQtGlWklexWzEt5laaQPYsXUHoj84QXvqPe7Zw49eaVe4pW9Ksv09m
widimnv0aalNYtZZVjjMI+hj6txYNX1a84LyJ6KW61MjWnB9v+rPiuTBkdS0MSOM
4wL9GCcLoBVdY0f+DGCl+Zf/09hd1jCFvy3IW9efm+mxJsfBZkq78pi6fAXApw2h
7xvIaJh9eA3qTSpB/eHMr6GKRTP3sQ15mIXUxiwTgs/g/hGlePmqVWtRILa8N1p1
TCykXExMF15AclE1sjzK89e1sVGMIUpNIIhQUdpHRT0gaCl5Sqa99pDl0W51GG2e
gDKRWdhAsnV4gtnUb/Q1dCW3NZihTSEUaNPL+uQUSQ+fv8mpoPMUgHhXcOs0D5KF
pSl4NXowuk9pPYFfqJ3wSZ7LGlKKEJWgyh3wt6dj3bfa8aXXe3HTQCUypCqpphCu
/P+ipJ4JIK15SRTC7ZvB/7Mo9U0XAQMwKlJtIuipJDYwlIH+C2zAnz7plWCiGSK0
aBhwTYcGP9JbVQHck82DyUzADv8XlL74jZzLS4fb/D8BlFMqYQyQFrCh7KyeFxcT
chYaAHi0zOkxEWuQplelFT2kAQ/okkDlZditMIL3jr1oc1o2PrE8o7jh93gDICPv
WSFce2HEzRnTsjz8dCQ9B+qHObwr22W0okOFTMwUFAD5hjGG33JzzAvWneOOhYlZ
o0ukXjkj5o+Gie9F+LTSl5ncQ44w69kVtfcNBrlT2TayLooUPzEZLYloOL0PIev2
Yb4wnI1Zh54lbsaLIJpiPHrY0K1vRXe5ESlao1Y+dwvH7/nel8h0qsm1FSw3TkcH
yvAOoWicTHpYCoqrbQB24wS764BAGoyj3K96pKOIIuouqw1Iqn6ezYCzCnPVUEla
8wILvVVgRpRN0AKkXAOlF+gMZspAQNiewryP3cO9puk0C17VJoQATFzIThW6oifY
R40btE5WKWhgcXe9fCAclDZzwG2ZyfoZMg62p923wdrQqorQyuVxptlQZ01A1eys
9clpKoWX5qAJd+3qibzy550eB9dJcsBmZB0xpKN53Yd1gyrPuHCMYHHh6PXo8dkr
tq413UDsSGCRMiNri0Olmg9ZxLUNXoPcoKDzb+BZUYDp+kM6imE7a1G+P8KBWIgl
N0TrvXVBOggGYC60w+olZ1kyuhBpYo0mdh6L6y8tGFXBsNYj0C03JhC15rni2v/q
mgXh0SHA8u5xo/mFARDN7hylGMZEfYYFo5MwsN++GYcvRACoRipdtExL0+1PetJ1
hmla9parOOabPfoJwoWTbLW3Jj9tdaBbwttV+XbwJGJXSFs+6IyU6tylgfZ7WbeG
9XOR6BgtjgGKXvqVSBIhE0Glrct16dGSf41zn51Gp+EaTXkqbEDjuAVmBQDHDGRy
rG1Qaj0HIPSYMD1iQEQxvOpGMEwBnXca+hqXqsJquc+RTPFtXsGwUPpN6WZaRng9
ufNf5sYhaFeelU/2OA2UX9Nj6P5mY9JP5xZzadBo2KNRHCnMuTHXUOuKY7kPdF6v
j0ycWMKj7PYo7P+VzJozwZ6nP3LFWpmnqKolVu/MsJ3OaKCU9m+hmNBSMjebSv48
F4fTyU1Kfd+k3lCkXdH7hG1czq5yNokJaa9Z6zq+GqM+qtI/ywRabb0gQo5BF9wk
3Uvv7VdyIzqTYtNr3anPoLU3Uvx2Rv46z5TJvaTG4TfwrcD8XZMluIeeLMbE/TkU
+pLsSVHoT8sJVU3f/g93ZCZXY3CE5eGZIH4MsTf1wUuwNi9EWtjb2fI7+fABumvY
rATCUVl+bd/D12A6n3JqbW8Y5PUHbbeV7Suh+S+VmW0d0sCVAqt8R4dQ2qFx6prJ
BhJadr6TaERdAFU31cK0cW6nLwQPYTv8raltqSmn7U6NEN3oZ2mzuO43sDq9v3xA
xeTK+Lnfy9CKlCXQ9wtxT2qWdBjxHhVsELEZQB3lAk0wuYWB6Bqu9oUFUwv18spw
Qlc4tgJ23Sa6rq+UMNEzld0cUq6T1zNYNfk1vr9J8KBj/RcPfzMCgeZp/DqYNvAU
lEZkAIYKL158xp8PDxe9d7nnX8TAxf0FTBPQltRmBkwKwaZn7Q+VAzzuKg33ZZ/J
ojErrSMgfDFbLyANedL7FOYNTfBQPTH2xfrNUo7XT3DReCb6DrzGSvGAaoaoVQZX
S2562E/cm4wNxtO4bDW/zNU+lloW9XD0oYvSekwmwzhfDV2Z7945ldufx9J1AeGd
RHIRdhKA5Nxb1e/hHgXai9m/2KW+kayXRyiPiQgxcXtlxlC2fw8z7mfqzOOi/UpJ
9cFOhK/2IFAcL2s4PbRGjGySHYrgg5HvFmbAuAFo75YbOZZhsW/k6FBvf6cN7Iep
Xq0V7uBiD7wMoa30ffb91QFAXots3a/PDOwpHOghievsleH/L4MbW7VacgufUO+1
UZ1Up2WJgqajNW4AiApQUGVfXXKcufPgYJmr/NiJMDTJ9qRTAeKjbb23mTpic6oD
+buyFb5/u9cfOCuvlf3unLSAM8mWsvRNL2Ele2FEie2JG+KR8fMRRXitdGvBoVEo
J8/YUZw/Mo34Ke5dMtSXmWCeLPDbwO/XB/1iyalzPxyY2AV6jlqq0PnVgNNks3r7
mOAejTYf2wvxQnGBkZcEmM5Bnpvzc5HKS27TzCZSDmjf94lCadPE6dYUX+9Hj7fd
gjHJEBWthanZSlXpOUsoysxsrDASz3Ntln9vuEer+M03bTNUbAz8oh8GxRaVX1uJ
lxeKl0HvTr7gLJvEI/p0Z3splpdItMCDV4MeSnLmdQeYuf4KBcHV0kJyBk4k0ui8
7L1VYxVk3O/nc7dD2l+hr7mp3WhCaTWA5X56kHK2JFdTd9If2HGJdI0zPSBCioPe
wc/6uapOkg626gdfG3i5RN6uPFAZ0XOcdn2W+x2nQtMrj0GDeAwmisXMvlLtvol9
XJ215ZGtmw4uiXjRg5euLth8npl/j1tRuP+ItHxFZoueYAQyBs5Yh3NT49LBizQL
7Epq9sqi2BOBEpsEeEh+EBzdLO09Oiq7JVFR9fP+IBYryiCnHU/abzrtbBghSAey
i1zEGYNsIjBIxV9vOuoFdYbHoXH41xUlOdrQqD+orF9gpPNIK4tSnCx83Yv32Mk+
6aqkdTo0hZZrsV68aQTdYA9tIhF3ZPp2ZXC4Tl+f0n6KegZcv/hmPG6AGYpHy5HO
HEBKCvf1brtWx8aaJwjenKAihRDNNrKs5WT8kxomFhqLRKm8iN9BaFB0VqECMH3e
pA4/nqvP4Bwt68lcGKiHuCth7qlYqbC1JOUsVb6gWFyiEl9jF/CFizSbXX5Ail93
BXhrkPKX1suRpKANLwYU8+anMW34elIE+0gYWz8opK1S76Bm8YTqgUAOnqfEk6fk
+fJwyCzJixPXFUra6Q9ZtjiV8CXLwu/uaQULFAiFpAjA7P5tUQyUtwiTmvywVbDS
D34URnI02KuPHly1l0U2hy3FkQ/Z4vyl7cuOa9zCgMxwcuhLt0OS6aWt6wlf+FRe
DFeVFS1Er/Sjn8WcZ89rd/djQOBu2xOpUTTK6FbxvjmCxbhc3NRCjEZH2hW1aM3f
PoweASgA5v7UxSh79UQk66uekxh9s5W3uavlTY8vrtuYZV+EZDJwY3qSRQXxTj1M
GKdkeWDknfai8388B0VhpYez13bYitSuebcZllCbxXWhDlNNqj9bwZ92ko5qZhLw
rO614+VKTtkGDbZznfP+N9ToMWE1wY7FQOBRqcN5GKdxYLUurNdpUzWlNFyBI2Ju
FeJQqG9xMr3jStTwRoP8KFscyMwpnzWVPDm+HFDum03cxtPdj4fa396TsxxKvRm+
2GoAlZcXr8VrMerq8uWhFned5f34Wa9U2YzsUajKPP+hR64chPRnZy4BbOQP7AYH
moF8u4MBmXbuBSYLB4BQ3GgzUwc7d9sihfPpRXIh49ZiJmJi6hMp1wlWX1lCPryG
sbIGQuqGzPHs4zJNr2X/WXh158KiuQRH9A/71EePGcKISUQD1jOYZet7Tw93eRcw
JsPqAlUV2+arTQPSb+ruxx5pRfMzDj5L0vrheeQMofN4EcNKbcccD036dyo1tTRo
WZav8J1H2Efv8vixxurumRr2T+9H9nzRCyKsKBj9RQcKNJ7A/Jr8Y/lQzATQ+07I
RD3k3FwMYyCf5M4j4q6L+9Gm3eE+4zD43tbArdH3p8o3ujRCfw37u7zRY5R0/5Mn
+U7y79HEI3mK/STYFAmozBmtbIi6CXIDHQEcxlh1+BMcSyjVa1dz7oMyTo+BHuXO
6owLERSERGDyIxxwiBfWQFNrIyQ6oPxWYT52PO+djqcpmMLWXvKE+GSSEgApEHAB
RkmVrqTdV+2Hdr07kGP55/nD31HcE6DHZw0Mb+PsLQboQdJ51crQLdOQMFyJ+L0L
pUk5t2K+1WADmKz1PV3kHVgLEL0Zn+cEvyk75s96vZYNlA1XIO0GQZHkLwVUERk5
mEMml2g50pA7uqsDAn71aVySqsvTFbvfjFTTcRDjdTZ8J3b4oBSwjp4bPQUZgA4g
/hlAumrced+yvMXbF2PnuGq8fWUXmjAFetoWq9iopHqOTP3NNcpYijS4MhNaOTix
ZtokwgomvPBOVMIa7uNWderMICLiCgRlUP2GTp4EM2TocbRWj2iIcFIKmt8b9sew
DxQzpUQ3tF7JzkaocJpiDydt2dMOp1qRTGGkKwNC5M568GaY1m16jM/FfkZ4nd/9
e8Gork0NJ6V2m0mtImyblpC+MeiYpGQn2hnMeAB9HH1fG/uIZ+59PI1gjAGvJiP4
9+9sGQCtL3SVn0zapiEex8xUsSNooMMxYZDLWuhi4QsKI/TkhMOyKrfgb7C73tAU
N3uXxJlSYKpU4C2IJCOAqqLYJrL4T+dVytsWar8GIitK37cFkL/VJHL+2bvBrBrn
2J57ViBWMCjub57ZbYTNBEjAcJvpPUszYc6Q0r4qCEOAcaooC+lWPOWKfB2Bd9TQ
G70hVFOTKHt819rGRFDv6hKxIGSHdILqMpzLwL5ZpemM1T+ENUNz7SfAOi/GV0GJ
mpkj0cwANXd4YoAb1ErfFixh8q/vflnYz19ZjGoqWSwBmNaVMbl+f943fmIAfEr+
qnYeD3NIZ6YVN8uik9vtArnd4htjJtpNzaOUlVbzHWjVKvwHz1nqwaqdO8qvn+2D
bJ8lvmqppf3xgNMhi9/4Eun2XFv+hIoc6JTq/PDrcn6VMhKqlOg5RG9HuP7Jy//i
k5M9k/H8oPQJyDFKE/+OySriHzYJpO90ifTlQAJs45pQ/4wxMlucEqKXsPBT4lXy
VSLPA3uagc+dBXklo5KW5U++hZBSan4NA6eRHvfCp28nbdjJnvCNTPJepInP70UX
Wfhc84BG0BAJ57B/EKoyADCvr9SF9K00rMmvm3tdvz+PYLt5U+br/5gFozs2LfXd
du3pT36y91s12U5ZSe5ZZ/4u2yhbr0vBokGGao9tEWNtG+VPGPeX8ATbiP/CFFgN
azvRbs6SJvUJIola7c6it7Ykstyrt2HRguG/X0scxLg5GpZUQzcxa9whCqu+1C/B
ZUFXh0SnIahKAm0kTvdWngHkrP9G8nf21dK/S7oBi6doX/3WBIPoCrXqDMsEPo2A
4dgVLnihOFgzoP9CmdUJombdQpXs07RXOJmZ9byAFEhkwNO+OO96nxtIwCuawFPY
WZNLQApycdqA1xtBfAxEzU1kVhMh1AGME7LL2Vp2v726f/ISs1+EnSnlZM2uRlau
3AXhKx3ZDBtyGeP+Dfardrglzy/NyD2mjIqQ26OWLedO5EQszgZo2lSESYVTZjjv
GKGZ4FxuWNFEKg6YaLJNN4UhSG51UDembxGFtCgSJf3fNIR6qFTNUzs8Hzs9yu7i
C1nq+Uj2S/QwtqhP/lCbZq7sn7AuXgY4LWa9Il8/OyHmJOCrS3Ufi7k+dGA5YM1t
+fwEy/0drnX+coswYblvFma0ubTQH2xYPCtLoNKZvrHai4ipHHdpoPfYYpHdohoR
pUqvznah3dghSYruTVwhkGGQx7HfaI1Mx8noIpjHvENCejlQ7PfEZExK6j/YKrti
3dXw+pn+LXvO9bOZGR+vHFMcvU7yPuCDcgvCZWU3e9DsQh+JGObemVEs48NyonA9
NKAfaJG5Ekg91l5veIEOFWf8L9uEgcjZv47TdBrcF4XAjCOLAC34Cv+z07MYruKM
AzvSYgw1GXNngOmX4v6V2EQKpfWdbMpCxas5IIihIRlmnYkJGIw7YidUf5EcOXbp
Vj7/K6I/sDuj8d5ePwmu5CpjGKm2HntWEq18jHVwqs9SO6lMgLWI98N/JhgOKQys
5Y3QhoE4r4asqP8qtJJ50y5744MC6WMsuSTOeorAXeCt1WnfuUeDKNPYzzp7tij1
MB1wzHZXpm5BYJccprBSVenVgCPwc5Cbx2XsllwtpKZQyO527RANbVHIC4Cf4txl
0qAu24hdRCv2XsjS3Jv3yO9Bwa8eqeewroqHNUFP5dGnaDCf73XxzTyopYzP2ryN
kJF99TiKLLP+nm9kSB0sGm1xk9wmCKo9anczJdcUjrrjx3KFTw/BNqFb4CIxv9St
gIQPuV6Rbb2/n4/+rDGdB4Y7+c+k0aeCTnDiJ9PZoH4y1qrFHdsWqi/92xl7k9IB
6Vti6mIPTwA/7ZVK9AWq7Sr6crqg3ksmy4UQw7wluxdlpQ2EbyT5Ocj7h8UTXbww
kO1UfLKrKZgG2Dq0ehsLb3c1QjHedLDnul2JKJ2nGhsHhqaMWs5thMVVM0PoXPbB
6zfX4UpVXmfxYx3QBnepgwsq/V0lIF+uB+YWkxlzRdC0B+q2zn0/0RkH/cCo1u8E
aCY8T+lX3OEvQNEUQXZq1Y6+2xi7LWs5vtkvrO5HYJFnBuyNRIhtB5m1WhkgdyNs
QD1FeJnAIAxZcX3DmKmjYbQ9a4MFM0y2oGEQV/4sg9+Qbu0Pe0WsGS9K2zocQ9Oz
WkaK62VCQNt/FBkbBsd95eHHVQJV0b2YZd921YgnKLM9IVrjufWckuu7s85GqS0a
kaq85wtx8aAKA9SuTakGSfdwcdiH47UJoGo1RNh+HckylmaWwpHdrcqN6z8+froT
96Zeidxzeuh7nQnmYZKwapahEHC5aQQzQ67AdQN/eJYoDg4qJMs9VvhBox/25jTA
H92OHL+NaARL8PBKjkIsvuG35lYAjK6jfG8MTlbqzDiUJhpgsvQhtYHKmRYDKXfk
8srBvm7Aw3T1iztlwaHjAEoTLQgLarsrSsK1ejtVIR8TBq+YYs89btllhqdLtH0h
qQiyYWwhCHo548Oe1OnCuUfHSMgzti6fgYDn1XU4P5le4we92gbZkObM9PzrUxsf
4KNSYxeweUyjplkHpeZjAOdF3V1p3rA8HWB9Egyu/+pKXx4eWcHTgdnqgmxrkq9M
JiX+qgDh/b47L86CL7aL4Ef7DjkN6Wd3Nob371ws5GY4oN0AQKPPhp8rOkzTw//L
XgsOBjW7Lo7tBjsuTNFWv8Oq6U0slIoTyJajI1NdBcNTDyKQPxP0yVrXlTKVmirH
KxM6oGR7vcjoVkaU3wQ3V8CZ4QBUaUST29hQAY4NmmRKqnt/33yuPidtPdb/IE/T
wKy+CvnFrsNLNTH2YZ3Kph3ijK1QyBPQAX8UHhW+twvquYorOMORUpHzxhOXxPZs
5qTWyTxpnkM1l3p5/dotjwR98jJ0Y3mdv3RbXE6NTIMgms6zMsZliSATTX3ok1Uk
QaQ0wCVUaniOSKMSeUeuO+Bnlyn5RqyJymI/D7RxPhM1yaIGHnnhYjtbl6NWtulB
HoD63T/U/NhqkIhD3bVdjoMMw+hQ7jruHa+iyLEfn8IY7zJoXrGzkOIbwpxJ9KaM
0flTbGYsRcBZFycbeQRbEuKbfK23WXGC6P7QcXbONWNO2rAb4AO6kOUepDkm/3pJ
TTk5JAzd5RbJPgBADDCEmlVGrd5tHxJpfBGURRYqWPnbdmuLRBfX+szuYJyu8d87
3BpYP6I7o08yjf2JVKxF358PVsB03NCDWZTEWH+xsq7XYeMSjV9Y3dEJn33xm58V
XVnLx+6eJGOB9dnWBsXX9/BPMmwxQh1P3akXplfru412JcVXo/tnlyGLmBhoo+4s
p+O1UWPV5VNNq/Dm1xgmcmd3RpVikI+dD9J1IVYpavUCbEN2OLxl8IWlZu7kWg43
k+VqvaOIKMZy0PdW6dSG2t6DRusHtaShEkXJRzQ6NLXrWj4GrLlLpd0Zg/lQ0rMm
NUIaVDFw4bt6j76pK7UHqhZ4D7SHKufKQYvry/hMtd+bfTvi0gPWNuT6/3oBQMUk
ty0UaW2i7aNY5xTDxKueJkyySJ671c3XyJ3v5Rynkf9va/5I0BKb+vbDsO/TMEgT
V3T+36+d43cJdr4w5jg7NXYl1Mcvzh337lwRSdR74GG5/CQAeYYh9u3rXG3UNSbg
ItwVbaAqpNoGacNzkwI4pVrmtCIlDLRI+3dbQq4dPRhx+6xfmZYkPIYXiojzNZdA
D68RnfLIlr6ltdb3IxF781xrsgPVeYr+AHhQ/U9KiFPPf9tXyt6Rf83JCVzsBIWM
1D75HnWXAGs23Osc6+cHIiRwXhzStx/Y4efqFJ3AeqxdvZRE6O3792lJfFdNWarc
BCyGkN4zyMTmrFka/9NDBQUQtjBaPRtoxGdI7OLWncIBP5q7nTa/r+igDLRhowUH
Fk2UF9fHk0OEpVLpd0e6VbPcU09ZaPNqimIL6IXZNJQSsniz2oZzinxscAebf2fV
gdIfrhQoLxBS9pPv9XXj8d98fj+qgrplFzdje8m6hcJPBNXu/y7kNVly+LwlN9/D
ip83e2FLtG6KQ32wra9qU/89PgAAZQf855A9ezAkzJBf9azNXsUvTtrI2NNpugkL
xum84vxWBJ/CuT3jKi1eTDhmaiwYIy6ZjBz9Nfbzwa4Sdmo9PDCa7EOOH8a1yzhs
0aLKL7dSzqaww05TfDRqfy9v/59zSWwqpG3i4tB/KqixbaMd5x7keK0EJDmHKrvb
jjI/AJmJdaDqqjLXRMjzukXLrs8fpo7kM2TTO3FDh+sswOwhDYc+/3U2hHttfJbW
JL9GMUE2pl7ClALx3JCqc2aWMYeIwsl38Is2isI+lNB6Nt0U+hZRH5LzrEIEQ33e
j391IFdjvmZJoigOilHc0tpbIT3WpA+yg40utvup0ZA5lhoNKB4j9v77gME05KX3
cR2IXn3/Qf9NiCbMkFOyyH4EUFlDWB7Ed3owjWJ7QP4dhZO6yLWkP6a5JnXlaHEu
Bi77NHDZwACUvRwQsXgQO98hDyZkA2M+oj9a+mwisavdc5xnps5pBRaGKANPVUCq
R7IiWaQxPm3JwlGV3yYeg/9hy6iZsmBvwtXepx5Dz7bh43FcR/rNQAuwTwwQxJlf
0Ha9V3WTFZufUAwa3COyaYZeeU+Ib3TrjHd16q1I0XqmiE7j4hD3JNn9TuYAuOPJ
D8Mtr4CYZOgwlRKkMcU1iLR7Q/7bUI2xbxqn4+fRPUxYIyCfxr1PLgAhzc0gtJK7
hwQyxADrA5J11BxR9JC5/72k0lkldvw3eSe4uxXGvDWr709pkayqFw3Za/4s96t7
IyvoWL01eJmKrexsqPVUC33z2C3rNOUKQP+3Ax/Or7kU7VSMrIeE9zRLXOkZqhDz
IYXXj6rIhS92uS2FkxVzug6Hg1LaFlRs0irRahz177pwJs0P2evCOGoofUbS6Ul4
BAFcf+td29IIjHD39ghSGBZyUgwzpKeI+BSpLqq7+zO0HMJ1qPJO5KuzltOs2tTk
MBE4uVTkfx3V+UijwgzAsUv9NXMGTBILRrATCmU9NBrar6I2kyf3vOMY72VAlEQa
QzKHmQ1PIIZP+KPYK7xg/FeeD89lrjCyXSyv1cTTJmFOxLKXmATQdWQBLz2J1rII
tIqsKNmEv2MwT2Q5bcHm44UbRe5qoTyZQ19tFPRcpmvoV0JZzXhUBSztS3+Fvxwt
bnFm1rksMueL3k4O0ooKTnVMf/OBceNDEgiHHrHQxo+PkkYmdvPUUFe8Uywvgz2G
ZHa7XAgB32uVIQWxiXfuNteq3nBUIDpoYCZiQEJ0zJZqsSJH88g1w5/LikIQosUk
7QneCsdHha3uectPjnZd3Mt23LwHKwwPp46UDLkE1ahG4RWe8DJpbxZDtzaxm4+V
NvQoe2LnJwqY4yrIFi5tWF3Re9zXgj8L5+cu0PhvReJhzwj9QSVTsJvkBG1H0xOy
OUtir38G5zx0cpkcix0tvkEPHeJPgXQ9cMR6oB9gGk3nLShV06dieTByeiP52cgn
ukxXwQMyhS8M7j4uXiVCRjaEhEgV+LsqQ/jopYfg6GpKZGqoeuOWG3BY/Fn8W+aY
ngAbLnfXDTc5NNZyKGwT4g+4LSOi5BIVb+4mo6RAl7Um8OjPH+REDgXb5SfRU2nw
Vkd6Qla9taE/X8Fj6D60RrV9g9hExglVlO/caJIb4UMpDBSgkeJgKfMvpinhOW6Q
bHwKJZY8b0sLO1yXMv5Qx4GSDpgAnksrHIM5K8PqQL46DphrppnM696RWBZr9RA4
mqB2sgCvycCxfUyssIehInNkTGoQH7Ls0MpgTdq2KqqfuOcsyQ4uDoVT1LX/8qpx
9GC/yn6sa8yNpJZuqXVRTDiWRibKLJRw+DVELyR7uHkG4pw87CMazWvr39KWu0qU
blFFQUGXkqAgYTD0Pg7tYRpmHV5JF54CwgXtKsA7aooyXOyGux7XBB8f54wc0Erm
yI9x3xyJBi7SIOx0/2Ppi6FacIV2WKzfFFWZAUJBLaRSLCCUiJWvk+iEgF4hGO5V
oTSHRGaAPPOLWxYLfn7PFE0m92HEQNx7vPGun+QETGNnQWWBottNvYP+4a7Tm0Ve
+GT7EMENMQxGxcxYSYSj+fJ1VvoTgjibh1s3CKgVg7UtMLsumJAB1rNSktt4eUSP
6kwA/rnzCfRZVjK4riXjRk8ROWEBQuUgk1Ak0zOyCW8WAeXCuPEFCuVp46OudAMO
YbiX0SAyyWifELPtEGCFfIV6pBsN0qby2YCj53XloNuix9QXDGF2y+fjBSbq7mt+
oh5LdUoB5ZP6qY6i/3hqwvW6QOV1NAgX0SBR3eNr+OaTu1tHfogmTzUzvX+pSm4J
4x+TrbgAsec9S069ZCl4YSq9iwS3sN1gc6GxyH3I3CblDgBOAwFbrJno0nmqFWsl
ny40+4Duv8UwckcT/HRsXKtnUPx/5TX5ewS0q2hwiNJBA2HdN572BMAwMylP2t7s
8E5G04gT1q4glopzrvZdvHeYyTB/oVLHzxTHlUnKjwgHkftff6uZfJ/dB3Fce2uD
bnU0d47NfVAzZMAlFgFWUmF34qyySyFyybH3tpk67qBAA//ZVykeTPbkzI1JJ+Xw
KsA+KPm7Vf3qIvRIjlYCSzuTyrG1liVoyfn6xc5cnSbTI01LswMv3xCsZgQF+qQH
f59YDhyWjBhNdTlEucKCAmVboxHnnWlPXIBJ2ZuacqXvjnhqx5V/QCLsPvnAwd6O
ClB2yW0wSxDodBp69HHx3dmQImMm0jjDzV1Zyg05np9TCbd3DDb605X9p8Lbq6tu
KNgUp7MMfzHpiICMN2+/aM5FjUYwmBAGriiLpCc3slX6N+2pFbMSEAUhoGS+ZP24
sqxO940I16JT5jXy93V2hbJ7EckhY6JOfAx1WvY5lUcqLi1KBTA+mY/zXKPEP0qr
g+HBvg3jg7ihiymlkF91gPCzeV1eHB22Qs4onojMlkqhZNbkUuAYyTPIe/9kfny7
AONTVqyEexaI0igaF1kB1S9nGkFXBvUWQshWont1fZ852XbskWvf2s0lB7SKRjfd
arrbbC8NQUU+d7lmOhy9iV4esDGG0wnSNjnt2890BgloxnHMEyAP38s6E+btevbo
7Oe25y6uLdj2bf9NRWuXKktWS16EGyR+4wS1X+WVUPDW1kNPBHWNQvd0fkvwDtIV
iKU6xPkQGQupMY0qBOkVZEBpqCC3pWL4TL3M5JF4mf8nBEMztyr8PSGeciLtAk1L
ZBlFIQoRyFCHVQLpAQSFx+qSCJa8ud41NajtWhN+H34iHgN2ruuUYufuY4e7KOqQ
U5oTst8iLCaoRmigW/QbhAOv2Cy5n+wqaqcyC7HtvrBt/9RuHiERL8Jg0eNwv/Ml
lleIZpSLPMCExipHFiLMuwdrtlfCqWUYBWVr37+T8p7UbUzqs3+2qB6vhs3l9hLQ
F2YIYUWGlWr9GInr2JAST1wRAFK+/hRyB0yd78s6e6P/DdQXD1jWkIuUm6V8vHs3
y5dAdJD7XCRZhl2SkMqJDpNGlkM3MpbtYnZ3lqOQkhanMY9UNpf5nku5CvhnnhyC
1dFmFG2OKoLWWW4I4dx2g+hunhqDEA31IJ3UKTmu8d4pwbZhZkoVwLj3Wk7Z1SuM
rzPgE17H2MvGV4bsUaJodlXWreRLfUBWo2V7L0uSaU5BMXB7ZvOdo/wjaQYO8rqC
C3CcuJw+Wt33jSAPOTYfYMC/mlyu1ww5cg+Eko1pwPoQagLZtK6HduE/Ol6M/bxs
Ceukg0B+o6KZ4KCh9CSzx6yo8H1Cvw6GE9k+owT/zKLv1U29WtJSaSsXb7MTgTv4
34gKWV83VLqpTQjBC4Iqp7+8tCAS0J8ruYL0wAjf2rQBuLqIcLgzV8n2yMpwv5Kt
q6M5FvwITZTBdkLOjsMZXlCMRsgnYXoq2lx8nc+6PuKTuiSTQ1S6QToV0uFI2NuY
mm36e9g/8AL3bO/2RD5CRFRUV597pfXLbubcMJ8k1Y9MhdxyATQJ9HGNyZOb5Mr/
AnMAiM5iwBdcLhyAXD+cvcDsVa5df4c7s/x5w467CPSDI+Sqs68xxyOApN0X9KJI
LZ9vMwajiASZuoU/LwZk7DRrRX/hCJb+3znAqfiBrAe8ojVdRJAoWCJV+8/OKR7h
BskeEYdn7V1r948OjkY6Xr+XK/uHdr+8suRDu82hUfHhbZK1giRLQM8ibu7xeOSf
lPYAfZPUx9AzgxKxjPIwZVql8n4rWZlMpk+nTy9MXW7okhXYN+kjE67JZw9fCvNd
L7heciHbe815rEuaKviP9/opE1aziMJAxQmvfCzN0hdH8Yok30yWrWqsjoGPteFR
JHdz3nB4QycPVzbvVSzSpG8fJ+Ma2br1Z1jEODmUNvNwCjC3q0CKdBz49/gFqoHc
vPLJ1Z1jusXKfP6KfWluVTD0+HlLjnpfvT2VaQeOg/b7I/yFVzcnMxgJz/fADEWt
zZFzp10SEXFsY5JxXFtuydx6PJcyfWbgJUOATZtpyB2atvjgRlxeC0a/WaTxRPvM
/0Qi/E1VAPlZfqrUepC/koSPK7zWZSbJtpi8GrZ/nnuSeUADXHAIAVgjOiL/Dxr9
n2nLg5KvNg3G5/G7YJv+bWPhnuV329Y7Yapu51f6bqbtoWeFvpxeIYtRVC2ckZlf
xLXkBNd9yTB1cRiPHnJ95kh5ionyV0k7cpGcYWSDH2TzwLdM9YR5TolwFU4qg5TC
gB3/B7kpga6H5X+oEfgCqUWo0goh9ZVsDU6XR6rJUtUIpLn/bD0xUfJh8lSE70Tl
UNd4qLsAGtkaAevRduTJue/4Cj8ep3BuhChZbiX0Qo9k6hFL7Q7Et7XVnE7mPf4D
c6enU6BInkqMduXXCtFEuOxbnvZFInqAJefYARIcoFAlssa6n6R94dILTdNsXykO
5beWPXXJax0h4wqzuRHpMHlBIUr9OZZoK6WsAX5dlZOSLG58/TGJ/DMEXJA1hjvS
Umw2ZVy9Ouhitu1vqfSN7QRggCbJNxipBnAfCrQBGSJ+8IOkPqski+x6teKvgSeu
Ftm2AQ06W5fakG/K9UHsfLo6zSSp/uWdSvzq+wg0esxkchjP7uD2r6Wle6kbNtLm
LttgVRnERQudN3t64zN+m8Jk4U9c7c+AC23UPNTKnjdLeaPZcU3M3ePKGAei9CSo
GiaGSO5agttSILhpSyb2z59bMBkNgt/bXsCpBfhh/ep9w+jyWn1TqtiMm0vDYKCX
CHW/S+HmTMT7ffVFz3n+PIPGIAuApXciDWxejDI2Be9ILhXg0J8KzedRyMeJmF+O
hdWXefbLCyhNYlD/EWOUnXMkCwcr8jCbW8q5htDUMIEFqVtlN/qT1MWtdul+ZLra
PCqZsbITjAt1hMfDCCyq6pr/+AuASlfiYivX5s2l3kDhEJR6a8EmZmjEaWSrdOlQ
HJtPmYDSKLhYo8tyYnWLBShD34Eth0ZX2SqPCqX9r5nvknkRkGW5SJAKSYvh8xou
ochleLDjUPAttPuyLpumzs3Xy2vPb61i1o5rqDUyWBtKTlmOBqg7ckSD8LrVSJHO
r21qt5xO3wNI9kcViTobYfz22aAUukNUW5fR1HyqTtwGzaJj7/sOpiGN1izSgYWz
RwwjZi5DmzPB2z82faUVzSK1XgsHc4cASNcESJN/HcRre0/GlhnvoPXaCCn/abum
fL+LldSdalspxL7YyvTH4hDfroBxskJrIvJ9SvniRW0A5xU5xy8qR0Ic4QII1jKH
uwjL+/OiNmrvzaFXSyAlruVAyuGeBMhXiemVC4rcyuRKdZUdsmJyWYqYcS/nU0CL
nsNYuvsVMGmwAGw8vyRJ9xM278SGlsGdVJnbWPzHdcbCMcgQB8DfMHySgljc7Llq
Hm4lLChAy8/BVF4DTK5yyWBTVnoXhiLhEY/YWw8fH9J8d2+eHSz185xvWtHrfgmS
JqunyMLiH0qFBfsEwiVjgd8jea5pI60IGbOhnw+p12xCY9s/ogV+a+U2Yeg+N1z+
v3p4f+fbIWQyqpQeDUxo701JH/Ge/hGdV4GAI/CutPvUcvnul/Og6lfUVb6/+vcV
0SaNwSo51GbXtGRPAQVeBOD79BlUsdYYWukixjqN7f7F99DJfvmewEMLrPN1DsCz
nqtgTJdjsZc7w90yfbHa56J6P2NXNEeiRicQs0s1nfI0/jVLAHCI6auvLalE8iXZ
AV6DieO9t4Oq/L6oVE9z2ohoSBKUFFej4B+F/zy4INxE/6CbgCluDXRnKTE6hxGj
FqK61KkEOaQArcpwVZCDjHPgObnoTUm5e1Kle7OK0bDz1cV5dnZ2OLV/oAMob4nW
Yxr2pKV9oGJKC2FX9ZgPENbwSZjDr6oObTn/9BAGEnO/POcZGMq9W6RYdvuhBpgJ
Uj0jMjroMSAtLRo4iMoiIalqhntVWbCD5yvnzGmimEi/4itJ4NRz8XID+4URO2qk
pq73ENsSlLFc4NUwS2WJFY/WPITZKQAAy9p28GMHOnld2s5jyuiRtujzhnDSkz/u
waom39yPZwCtf39Hcc9QhKjRNo2Gn5AwZ0MLMZ+ll9cdsL/umTwHrF6ngPRIW/cV
HkNzM22oR1IMzdZoBPi9oZvcOpi8amM8e8A5ubYdE936ijISrtW8bXVwevm5P2c0
yp8JKQ1e57QZGPcCQV/8VPwBMZl0asMg/vmTXa436xt8XAw/Ztzz0OwGuIrpR15a
x0hyvWdEPrxAX55EtW3vE2xD9dMEZ3aEcrbqjUNkI3sFWeNVf4oA7sC+wDbqnhWs
WHphDdbGH4mFGeFu8EoBmUGlyYrmot3q/0oEFO3CcDUMTVk5lb7S7lJ25S5DEbXe
p+fKVfsPGH0kngWnRZS0R315yzpZuK3FEgIgYc2ZJj1PxC8ZcuisgCeTSZFxraex
NAnm1b3oCQsDdccGr61G8H/ShNOkPAcy8rzb+7+qfQMPcTIYV8nMhp8Z/a7zAxWV
L0FSVWwoxSUwKOlz6sW0d+4NRlKyFLeLh7pvRG3sbb8UI9SGuRAYVdmxTEQL5STR
POn7dUeibf6C2Kt1mOXqfsA9/5IFVRt8cYMYWm5C4G8ZOKas/3YEbsxhLiPftKqv
d14eIym04rDXLJPtbBceST0EENmlXZyvJlRdiVIdYJbzEJaZ9QjnKDaMK4/KCm0d
GtXD+eX9M4x0cAPqIwdvqIZChWP8w/rJXUug1Hx24VGAH+a/BdplwjtvIJs+Xl/O
UIyQok+fZDCLfkJBxDHTgtz6Y7xbyUGROh5pwJ7X/VgeBFsDUOUD2HLLQzxwB1iH
EJNTqJdTK8OcAfto2HmZENExeLAi8Y6KiLwiiue+WHHlHu5krQDqSsIGVv9U/OEb
MjSjjS5jxvt+UDWGUyWTkUy7mGdI0WslLYtsLV7GQ7Mk9OZ2DZ8I/YNu60fbVAPk
IMtElmFlBoQPeBQxLMhuYr/wacWgbfUiAenPGIjzNV8a62TMvn4Wn/kPSVo9kU+P
n/eTNF+uyUc2Om0F1oxymECboURO90Jzn1V9S9oIu99U8DfWXFn3JEXDmrE+yA8T
ejWaMKfT8vCdDBfCO5B5Uvd46A7260zuxaitOxKUmcfNOnBHm8S+jKPDdogFq5R9
dW2VmnPWySBWAa/07c3N14EGRxuj8QcOqarXKVgcklfzTFmiT7eiVX5Triy3MVHn
6zmtFawDvWENiAcdcr3748ESoLcrV4/GCUmK5rQpE96mCR6wa4EVktUVvDLvcmGy
wzcNf7qeizIKlWJeOXbismZp208SsPdQrsdsPTyNOFFFf6MwkUrbZDoGpLUNv2O+
l2/ZaS2Z1DGtZb3cG9RDJknkTwP19JuhABiCOKB+KAc/fU/GSOFjhRXdaNVt6slR
6w/R6jCpNHSPh/XXa4mj3wA/0JV6vswDfsXEDJNNAK5JGM2AoQD6PZnCNuLvLHWL
fOs0G4xae3P2TYUkI5JLRu5CdAviVAK3pr6uRxNJDrb2IsVyrCyzomzYCCcZaQxo
44Hfc/iJZNtE8/9id1CbLgKUEj6GlMD2wCN4TLzFfR3yjwKj3MN6MDzxw643/tMc
HAU9sUh31DAZE4JwDupnieeCnHB8fKdByyilvu7kxUd4d0GJD+VW2deDrkuEOwA0
ZagH18STxiPPX1LiJgwxgW+KrRMCtcJDAlf9K8JEuNX9rm5SeGmJt4zqylZ5J4h5
OSBy9XtVDhbRVFE1YCC2/mf51Au/GLbI35Y8GwAHi3+Z+lUzBNycR72BkXT3LO2H
w9KAcdJkmz2b7ksizRzn6051EFvCoypdzFH25H3yoIzZmQEGvz4JUbBR7UqQo4Zz
AUn3w4s7h/oMQExHJisUzBQC7sqo3jilKJDNMYzCnca25YU4j+ixBvXFk4qf4Zcb
YqRa+WW8+ercktcncyLcXOngSVltdc0k7HWYXzjSq+q4ycktuGgM6t+UC1Bh/I9/
7NIy8Kso2kCMkJpK6cQ03Zph5b0qI0w29DhE0W8DPbu3QFgHN8JF0kVkoXl20Brv
rL18cVSVxT/Ibr+zC+QLZjCbz5vU0tr1vsZecx/S5zLUPf1ARmrXrFx2T/8+tSA+
zBAONughQtMfiZS8nNBr36BGjAF8eKtuuDWvfmo+VIcLxq5CkNIyX4KlL8N0iB7b
67feWWTSZnrAcrcPUM5xmuN9VZWUnNwzeqbbx3r8b9AA4gl1OYKIyeK55IFaoUXi
ev7ttJfK7YdchB7RLSjeKqesr/c8YYVvVEqYwpG1OCm+kWDh/v/1FpcsF+bDyLWJ
EuwBjIkhdYr4S9ALISXA9AFTw4R1HMMDkSrCSwPCH2lIhrQhtrt32h9YOlwqZ+/P
IC1AWBOyg5O6NbHjIzqs67ynRuAFuKeqROUIkNsXJ8YFFjoLV1c66A7j2twniQyZ
fNW0iAAy/D5LTDZaC4w3EhunRF3liMcXphuVpqa/oPc7kgM3fhlnaCo1X3c1scWy
yNx/3EpBerbQIkUFEulKMiyoSLnUa/egGfBnTdVRblt9Q89rXdmZE6nPhQ/WLWpx
O5zVSJrZf2niCqs9s6pk2dKg0I6Wsj1ZrykNUEX/Gx/YIh47oUZWIp8yaj+W1SL4
NwIM0S/NOz6cyS4wrPn4XU8K1nF07ctr0Z1FRdKgN/AcCaFxvLcS8+/KUbR+wBDW
zs8EWGH431ILW93ubwCpU+S4Pi4xToFE0J98YA/roThCk6xHNzzsBu+EwFF+09Af
XYbBDB1SXMLsNIARUliSUAzlGJ43QgAFMSwMfvjR6uQ1rWyHcNXaKNFKR9RVaHqd
/nC6O4ne2NFoVcdHcp0QiXmCEDOSpXKm2yUgN3r3kJpIvTEpAecYvM4MPqIhjSt1
TP3u3nj/B3LzVw2gYug0Noz4no+LG41SmDgQt950PnCCZGhPeDr+IhjrXAXytMff
ZnDEnrFW4jjErRjd4yL3AIUlKfCeU5pPheia+9EGVA95sidOXxseKseZ/ixoE3JA
INoSFKvxarvm8kbvwOl9h8R7KbXqAbyiZhJXityvon2fwgwRTisFxP6WP0KiCS8e
9Pj6fyNV2HK42ODdjOOvtZixT8uiGN1wbkkziY/GT1pGpnBDZ+4c4hIC4vxk5QbO
7axoN1CTSoIfY8S7/i1AwFA8a/TZbY93pODjBQriziLybntcmUL+KTKYwii+JtcZ
liRpUOcG8ax46yAFkfAhPGfKXFnY3Jpmab+T3Y2sx27Sg/g5wMr9NmrRecuF201F
11vUo9mUBI8v1Opxq3d4Tzpt94Vr63Ecct18tXc7NB6AiyixG765lU8KQXeS8qYx
iOCwDW0YKWaDAb6mYymkM9e58l71TY4hbjvDBD+wCPhu1zF0aH9Ust39jgYMSHwa
b6Wgx+oMPUxs7lVOHtR4D1lYrLh0CL7XqSU59ZDpHRjofLbS+ClD9SB24pOw3z3H
C6e7xqCL2JURwts6YqAAEX3fvn5PYsr+xDwYXJJpvSbxJGo9Gl18j7RSEz13qca4
YzLFtn2QsIu2yuG1gZIVQ9dsv9DKbqkyENi8vqyc1RVJ+yBJkkzkHM5YadGV4mgV
h/mGy3oDEV74wVYknU5MqY79cx+cTAnaNkYZud3BSdL4vchEzu8RqY2V1VhmrKwG
wBgA1SP5GjHy+1soZ49V0fWiIFJlu9ML9vrVfE79OdFmhDYKNVEX8s15mDNDhphX
7LXd3r9saScyBtBExPLx09wZK5TxQ5vA2+Guk3dDhjd8JcLzGQdaN98u7EYJKvOL
d3i2s4YHM3sqDtoV4/NvLgdyiiipjX+NBhoHYRfmcMpFu87Xt1L3PXM4v7vNdJm4
syixnHUIa4Fe87PmqWppD1VBhdXj0VghR20qEaxM93jDtd4u2xZrElV7ich6DAeq
wgMUqfIGxArXL8J8Q/zl2Ec25bRj7OfMJQI/+kzpBdiORJo2C05DmmqZY2ZD0rS4
aFR7mNQtRjvlemySoG4X5ZorEGtMMbD7sDyZPhFGWW2wEMH5th+1e4K+Ra3h2ud3
bGjY2W2BO1DvP/EmglDXX/sIkrUkPtQu1zhmkPbmLZzT0R2B7TRTC9TzFwmUxVnT
GVMrAWLsrjXd/JMAEftzyDC6xnn72hSoo8dwUlWoMcslz43egcTqLVH2W/08YLu7
fC/7xZsHzo/yRI/mjgChK/ymuK54AuPmHvfPv94zJeAk20Cw4KiwjXqadYgQMJ6J
Kj3GLf2balUb/x3gRcEdFehU9swqcJKkqK4AAJO/X2GCl5I0EhA1znZ27Cv9sdLx
cmcNBFzizRVvqLklYB+MFc3QH7fjluKLal+kMP3ePBYW7pROxvK2K6LHKLqQCcyM
VwNvJpFdxsggqtTGLDyrMKRhSwoQsVtTRJtM8RDgonkulXVvnKmUpvVzLFyIl1Bg
4LK8itcX4MBMKA2pId+KVHo4ODdCBbAMhAuXyko/7oAYVnsoEmBYNbSbwvd9g5g4
+wzOJdAjc6Lajn3hzHT4JlT5+e8hjDTT7ccJxLrEIdItihWBK4flVSqCTVnCuuRD
D1yYWUI3aOwNXcVC1bCTBr6xjJn/ty8iyzsnM2jQo4NND8ziUQlPku9zfGgfXOwo
jMfAOiIAmgm1NQP9k+WiQkCSYQ/lPMKv97SevBU6D7kcIbfQ5wUajOdAGjso9mqJ
LQ/iIwXkwJAxRKQtH9PuhLtjhUHg02jAB6xRj4lmlNhfPjTQqWRVXbL39PQ3G83B
jOAmMibeVwOxJIZcenyHml3kZor+qHeK62u0xo8KHOZoQwcOJ+RMTMHstJ1+SgLE
gbQwuBZC//etEBP3Z3cQohsU+cBuFEBq0Z6eCXs+km94Y+7xkcpO519saG5WQiXv
rajV5LJhq48CDxBgtIFprytgUFlZtfZEC3ifZlznFsil01KT+xAzlCt1bnW7HALU
K9BFURHAcnsHqE+3RH+Ed+C1Ef3s1CsZ4HcOsiJt6+5nJhCB440TvLn8nXT4s7Ea
zHfwng2cEe/AlGJkpTC+D3hwwk3sY8+rtDjZ20fu/XeKm0fl4ATFl8H2k8z+z/S2
VNnNJiQH9swT53uCJD2La3wJQjCWwu7ET6BkLVwY1jcpufcdWEwTs4c58hvewWFX
hL1RRjstqnIAmPQ5kxfPxHwHCIqMbof69LWRAdn3kVK1hORxd/7OTOTgJrt62G89
2e96NzfE9M7Wx+QnIjK8mPz5GTSb1kcRCxErcKMjShssvAlD+QM682DJM1+Az4ir
5TueMYizmVbk1iVrtEq1CYPSL9T3aqI3yZL/MOYmRQd2v1/blcKLp967ko443yPa
D9l2k3ZkKFpVFMVeJXacw51LKuS6HeFxmOrNFqX2aTy1f5xANW9KmRU5rF7edBDN
0QjBHyJFaWY4/nm/JKNzRzrWRlcTJ0HRy4VeQ5vJiHIshfwzLgdD5lmx6eJukEi4
Poc0byxtZV52L7uGrOJxZGvu+ntQxKAhuoNB2BrtwjNBbRZEhyBButowyeJUvyZ1
LV0B/uIy4iRSrUVfQ/5aMxpavT6wlHM2CbkJ8wUGciFORje8zWIThf4SxYTtTjQG
S776kv6pLulaNmMC3+LZ3OcmKQDR5fLS4ll3X23T7N5lpk+LhY23sRIWtGzgG6T1
rF5q83wtiG06cAKsvBgt6XUPKTgN+vqTnrl60xFfpar3LKH51jGSfg4GaOYSrwQn
irV3aISiVgsj0b3swysrd5xqrhdFXd+fK5nedt7MEfIp+lKe37/LtRVUMBacEx9o
uTErSYQ0H3uzFo88a37xdMJcZD7mAAmft0wc7gIJ5nj3kjVP9dVJ/QWbJd3d7GVH
vX2K5mLJriW9vptPay23i3M22Ca8IcaEXgMBynUNEtkoZkOPVKskg3yPfzro4+I3
o068x3NiEOTrJZjDA6NFC+vpgnhHTyExSdxGvG7CIlbccmxJlWMGuO32vaMKliyR
pv9U83t8+G1QiNkXQXHUf163dULbx786vCNgvMt6kEUg+sUXGY+wFob9B5Trk7zc
7kXKJQc2U0EOey7KDBQjXDrQxxN+hKXeHqF/VA3K+an0x3rg9qSKREBpfz00imr5
+dSEaQwOBoztxZF8dINfszVpUCheY/D6sv5ByvW9mobNpWOPRoI0+13OEELz2s0N
HrLZ9BnN5feAr1CyEILu8PDYLyD+lMebWqOrbC9s5nP9kDjdZNWt9gde1wJ2hoWl
wgiRr03XXfp/pIRf2L0dp9hnrJIwKnyJj4Wb6Se+nKEhBigPuTlo7c8H5Mx2bq4E
ndjho77Y9/QAguQbTrj45BrGp3UBBp9F51i+HJ3HRQrbx7rmxwHR+TSvAAvPKzr/
FI+hNZrZHJjbJqjkaCV2xrOSnSfiNKpFj1CnIFdNHkR/8CPXkHMWQ/qbBW9FR+vq
5qxvaPyCgZWMaVZ3dDb1mlJXv3V8Jzr0pV49mFNAS47teCMleUblB7g4oM75xYEn
HeN/TTeKt3/nubE0YXu+h9Gl1Q1FMKFsEHliEbpEtrPHEyJSenmUG5PQ+WODnBeJ
16WJyb9mUtvddbwe1o+kMhTxjJl8RY6lnHgZ1jgeEhl3Zm52SzLEv/FfZLkN4Qbv
F/hBxt89zj7bNKsyZy77cx6RAqlpjNDZ6LDtjaeGWWvMulV2U0d4FxQN+7QLe8sM
sgp3jgCuYDp/QIym+L99XYR+tLR/9AH/LzQQ9mAZjoBAnd0Jug0taujh3TbHOkai
WjrWr+lIPqez2wbdgL9fYNrcIcFeG5YLbrnS9X2Di1wV98Cf5t/Rd8eXqjTM/oSZ
xzM6bRdgsvn23WBAVrXkhFqMjhC3S3PBClgRCFcY1dfcKz4iiZTNB3JvFxNRoxQk
p9ucYPxW5mLDWSqjsc+R3Z+BI0/f5g5AYNac2qbRS8c87LpW76NZ8vC66U+bUNji
SE3J62yPNmxlepBwaPxJAK8/eV48LLaLTquqw6SsV3VIYthcT9NW7JZC2hpGWLHc
5Yzg3IiNJYAU+RAfGk8vmzZtP9SKHS+VT+Fh1oG+b4UauFO4mocqyqSZ+FEONnpc
ZtdYYcmsErGbrtJX0SufZqC+eFX7/s92YgBJjpOQJOwNg4nO1gGO+g5q/p2QjBw0
50BI1MvZ/+WPXo0v/nRMe1Kn/maauJ+Kf5vYe2iKjX9D2dhwmkiVMzAHptp2rA5d
NfN/YAoOSc0lyQff8Pk/6Ec/nSnffLbW8Jdk225ERuJSAowaR3XgeARlRFnyRDUb
LjC+qCAAb25vAXHt49hZWDyRTyGnLX5Chk5izAec/0+V38QaCoEcTQGq9nRig7d2
V8T8tu9+5E9CWR3cVQHIOgoIiCcaR3Skg8DZfLRCo+LKVS6wcxOdxzGv0JSdkgg7
isbDQWTepPMyrhZ0DvbL2vP0WjagiZxqusQmmskmFUlPxzk97JPI+h7/CnIMTKbK
VALPhgHfM33OJb10+cq/eEZ14WeLPLI88uus6jhPnVWkpo7XwGN9jpO17+9Rd6D3
/1niTPcewJBIaovtU0MHwAGiru3n1i5KT3k5K9Bu3X3eHz/5rev/HD9nBghXIfNH
WorSLj9c6uNnozsibT+kiTC62J995VGKUCUtebhNIjMvNY9B6HMQkuV8932cY3AZ
KZhkD/17vtoj7Tmb2qldqAGi0ArFTLmpyhp6o0zzOUVhR+TXgPwaUIpX6YXb0vfw
64rkUSecytuVkSW2KNBpMYwD7nYpF8H35qsvml1YBkH1G3x/QSqAjYQyYKqnJOwk
uZy9IGHupNXg6cg1OPa7fnX1dNFQEVGLkADMppydWoW5Kug5E+D+IF3gQ17uAH1/
bfGdB7oDhaA7tCh9RbHxDXnuBN6vkO7cFZn3aRuTJYGStBIEet3JiSkKdtDhIAGv
69o3jh5+95NlC+DaV1RtVKeDd3sM9H9oqrXQzMIQ/cgSjGusB486tui/5wssfGiY
1DSXC05atx4oczkY/wPujmLLchxOdMXIkzaGwDCdYnRcbLowcMyNB+QJzPZND75B
dpOGfXCWyf4FxQ5I8nuz8yhuzP+1uU/MYdO3GCKM0F4f4J0f2T6RNdjuXmpSY8sy
zZ+r/ZuWQPxM6/urzenLniKcvwHMaGtnucanE18YGnxnxAQgjQwRHaN1be8cN3oE
QiLQGb17Z8ME0ShRm9wU/IHzgxr/0s6N+k55YiWxnTND7GCr+oYW0pCaeZk+4HcO
xTKysmJd691LHHye5LH3S3FPlBpaAEUiFX67VHXToSPc3W6ZgME1zZpCKKMjj9lv
Rax9Q3mriJAvkcPRwJiPkkTmZuUAnNXWEaUQUr/ppxA0H9GquopAybMrHmQ/xPEt
8V68xla5iePMbZcEo67PqXqNKoW7ZuNyM3wLEqoGUolqIm7gO8i1uB108kXWdSB9
ojPD6qQsFeXBmXq+FxiwqM38DBpu5Gmp3AWA6GiIwYz79uXrXmveuMfUEQ4xw0v1
tvcajEgslMRdnPFouukDbZzcua4hiJRBo2MzGtHDAwaojrzrl/n2HaQgQR50ohup
2v5UknGxtKfjTWWjrdVc6BNQldfiL9mAet0moR2yP/eR4PiaGF1uztKBYLj2sEYb
41TlTUc+tiD9IIvkxhkMUzQDhzKNWvf+B/78DneeFrbnAyaiLH+vbLZ2y4G5xcgP
jp2YwUW0HXsY5HVWkRc1jsLVcduOJJrniY8kV8cWZz/JiwBKvg1KPbbSwC/+kVdx
nQQrocZNK5SzMr7PoVvtCck8X4fQ5JM2MFCvIYY3I7JYANCfYnjXrql4mPtNhKQ2
uW/MyRvL69ntSzkmTfy9prEsqaaBMbi9wTV9yEqJjogwk+OY91e8KcEyTryKNKkV
ixdbwFrzSM/qKFvQk6Jr7SEN6NV03BWBUd9m9Mc70bYUtaqf4hAY6zOmiglqHBUU
EaYBrg1Fu+J29wTaYaEVMt88MWfVqRS4WCw0vV5D7VRbszSWufXshmD3V7nTQttQ
AWFDnGA6YQBSaoRGOXPqoGmPRlZ688zT4GfnFG1/IPY+tp+XnH6GwhGXmAZVq6ws
0jSEyiawDTLXkhO0IcQQ9vdgDRG+01CnvJxxYbvrvauXJbzeQ2+nyIM/XJr4TVcK
5jOa7UIsEWzFJO9Puv6U2pc2Wj6hXpwXrXbqvgvv4jskedH1OFpmhe1ibiKYX+tC
fXlow6Cuy6ZKV18P6uCwIY3V9fQIp3TJ+ts0D0eGrIqPCkUY63UR2HBXnxVL2MRi
i1TbMcOJhPfG6FZ0mtz7obmj+HBA1oVxRryJr4omtj7T8X7/N5MJ5i4L1JWqDa+G
tvBKqFGGrMQOBbXi5doKF/BiJPtJNDegqbhE/hIBHst1k2CJsd2bqX8DscFnsjz9
NWqkpJtkgN0Z+MgdYbaD1GswaEWZ4E+u1+Q+YLECvc7f6NhZACW5XPYeIUDeY9pQ
CQF6dZ59zodbyybuhKo0IssA8EtI8uti4eNGnrtANri421NhB+GNP9Qksj1L+hO/
aGPtV3vRT5HzouNsxHqjALES6zLqEpjn/tnQyPS2MMWi9Qv+WNYGhgSei9rEb034
6f09G6X+wxK67J53IccAdEJP4jIOrhHB6/MtyoCCffFXUT9oljCe3w+Io6GqFuGe
yvojeoqM+s/A5qdqyJI/AlZFrbqjkHsh0eid0P7fDZTnp5QuOKmk2o+mpzhStOfL
6Y9m/8FugxUNM5mKWiFTcv6+BUuIiR5IW6dJfo5guGyzlM1La4SRoHVsd0INd7m8
ACEK8Y1nZ09sDviJNUU+LBZlN42bWGHzSvtNOHBg9fwaOVM8HNR3ns6I0yI34trz
C2saDoQSu73BPK8dIU47QbmMXcN6NmNTMly0nJUBDkAq9rtbRwd9gnIOdigDwPzS
qICftC/QCZRbvhKmgbntSOSezBaVhcB//mnBu3phMksZEnf6huk00JPvrEJAALUr
mfjarIYQyB2Y8MlsHfFUFuDgwX4dr2cSNV7eYFND6akKmXDi51hW5gBnTZ83H6uy
kpXcZZIBXUkNmah2hJoisdimKqfnEu/9rF77dggweiuSqBsIXkgWLPnywutOCVol
59Z30nIDmVOz3HlaBlmUtcSHslIMT7kUx6R6knYMJLM8ZPkoj2usshL77hkigQDr
pr64GLpBDIAL3RWRLDhzyzh1OyMyokThMNFKg+ozJgRc/IxIpS6nJSB21CvzsiwP
+lKQTC5BOFmmH/ILWASc42YykIp97DnfIwKUkJz4TZbHAMokLS68N3iD6IAyFsLR
CKrZI43AtsagOk6L5lSgzsWKLDiZpJttJMxOIbRbB8p1uRAJEUpON8Q7mOwKmR4E
fBE6QM8leVLp0q6YlgtEEG9dVAXfYawZHhOIQoitEbsJs0O66/B7xCx1cM5MAOOG
xbE1pca09nZWP0tDFu8tcB+Ex1JHPh7CJKIvqz7OEb/ZQr1eGgomRl4k900Xx5dQ
V0oAxgzmhQhonJjgUA1SMC/JtxMQz2fcG2F6G2NR+vzQ5USYtW3fgwsnv5dohtxe
E81w5NUznrjDa5M+Y0csxX+NbgRH8slstXiDWvooKutMNVSGNGj3Z9c5+BI/7Uyn
KJAswxA3T7Smz2pwciw1vUcd6diJx4jgkllap2CMgOMwV/tXrzCCIQgkj4YerVlj
2N2dxaWk0Y/eYyxJpg3fz0ygCe3J3snkuMpHSHIp7NTWv0Ubmx7Ifi8eFcj7NwNe
3/XCiRSMJcxGTaFoATloLY+sRd8RkHrdy/PgS1tQ0OOhOMhFyp+f+iK0Uw3EX909
K/yvjOdQGP+1AapmiOfa8+Mu0ysLNq2g/OubazQOUg1Pz4x/HbZ4Cf2vM3rtKs2+
2hE5h3wnjM3lHcCVSwSkN5l5eW2Q/FvevrCNPtS/TmEf3fH9+SpqXrzeqG4k0bAd
aMomAXxphgGyGK4fhQYi/ILfw5GSPrIvAGx7+dNQe6Yt80zkfkgdiYX2aLQOVPqI
jNWCBx1vCtlx/W7w/U75DocbYGBs6e0d/Hu2e4Wc5/qa7xJbnEjGCZqEVBBrLSMc
oaZMAFc/zx36k7BjkObvj6KCzla2pMtjgl42JNgtuFkpVBTw9++72x7PLzE+nyMF
Si4UYR3mdWnUS/+ME9jJt0OaK2BAjlFarYFUIjX49b4uC79gqPxn+YryiWCjlS8U
8+JdWgHlRCEkyvBAd8dhOO1WnhCQNwav6ZeeCKaRBaU4WSQ6NH8+mnqRNLKyGfvf
1yt+lstqio1d62a1QepsrLcR45uNgnQ6mZWLOfMu4ErPgaIt8HQcTcWV4ocQb66R
ZPdpu34vqhB1cSYLw6EyT49gknZxn8WfWegWoVIhdY5e/I0GulET3+Wot6cKT0JQ
y8qyXXExpKYzjk6mTuUAjP+tM4EhXt+EBjLx52vFxu/0AZWr/hbPryw4Cz0SNSg9
DJmdRMqvXvk7Q9BE6JqMVC9kXYwvLjEhho4Jn2F4p+g1d0XwB93LXik0PgPLeD+q
74Gl6jTn8NPZqtgPeU28/CBEmnEWiEQWLBwvOvJXkcQIhL1onmBEZ59rAvKQ4gy7
fowyIcsBNNKOMTDeUppQY6HjdJjrO8aV0bh1q+UlzIkoaFt50xrLTNuQDI1CyFbz
NVO5vcvZPHGuBeKeatKxEnCfy3gmLrMexGSOtWTDNVzl6rX7eq9XOG++Ze8lAjES
m6aqLcPTojprfCvZyBhPp9+DG6QCa+FNy6TELchX2mSTZB86dHN2vxD7hCmMdLPs
bz2y3J2HF9418SzM3oNG9w/QHRH9NvLkcH+i+0kAooRJbUXkB4dIC1P9A8ErQ5+u
AYVfPnNPqPR0Umr9v476L42YcB7nJ7FyWv2G2gNe07K7cvscJfT9aikpRkCH/fTY
uaY3QzsGgqnThVHQ8uoFGiwUXRJDO+tPZMHi6qjaNjMt0JPMCv35sTMYe/7uT/LU
xHalvnrjzOQzjpqrCHMvJqLzsOlOVFDKTppUj79lm6b3IpkBCAq4pYM7UlJ/Xtz8
HENRSBuK2AUtFhykOk/Ly5cUWPjfEDXunMdmoYQ25X38RJt7nLzLqhStIhl2lxWv
HIBJTD9Dj/mQH6TRoWAAWIXbcRWpEoSKzELx+fRyquPbXANb0+rgRC3Dj/WtOAt/
k3IKrZ+eLhyY4wDHSjrNvWV4XsSnOflZ2yTvDhZ/oW4oHU2rHB83MxFZiltgPadh
UbhI4I9ujHQ951TdjVwtjO5KF4KCb/ykMuCmTX2iadPHuqDmh2J6b0D9tVEUxoIf
82JhkbOMhe5sO438FhXlDWXWPJdOo0kYYZ72JUuO+DLmD871LaxX5q9b3jYPtspM
FgK8ZQQ4xVKgqoteO6hDsGcK8vKNOoAdBH/BlSG5nFl4qFtibsJkvI65RJuy53EX
pXMTIxIivc8FgPK31XWShTbGHbNhbdEZ7JX5YaTVnJdhsyqcGb6NCGI3gjatCjKF
UaDf4P7SGfhpw0k6AUOW6lBFpMl4v40FZXgI76pGjG7yHFL3LDV97YnaSzIWaosp
LVmoRDA714/UTzcUQxRAZHTH7SLIXFM2Oo3T3UpRkWGmESaASMqa2xlts4mAGIYu
+5P8IdbGH6eWhVwxZhZxYTmMB3DFg2q067e3X3Ga6+oslaneDRwHBbuIFazhTwUv
2/O37ZF9ncXtFphVGvNEDgvRyKCnyZyltDNRCujX8P5ojm+Ittt0pZXZIJ0se3ey
8Bz8VFicpzI6j33BOIwWDck78NRXDzMXBB9qDPXQFV9tLPfXE4pRZFHnKxcOq8EH
kyUyGRWvcwJBrJNvm3AvQGfwANMEARXsYdfF6/z8tNKJk/bqNtdABNF79Sv1OyiV
Gv+PJiaDnLgAh9JO1+xPzFZqAMDRNE7RI50WkcakuOJRzsZQdBKtiMy/tBBYm66g
hSOnrxH4RCE830F6o5dFyYgeIB8rhDJEtH10iC7P2k7jxoyiAJ/Pl91IExsc2/Wg
cRif4A/HRI/Qi+sr4p/o40yoIuXhBcwz/1Q3INuEgqIJ1GGmMdUBICmet/VrX5lG
ope5/ZAusqBG1JsRRKn0SekVDt9N62ZnjQ+KsBu5fD8M63/QXt65H6bKkZh03Qge
RzmHh0/VBDbBO7vn6H00rv5XnvFGETWvptjl20TVWFPAlwQv2/VSm+5BeQEZaDiV
bm3s98o00Ns2Dw+A8tJJ+CqEYw3HgCzkNpbDQIT6Gjh1CqKR/Yb5fZhIoUid9YXO
ng5+7WfA40JjKmkcx6pLSoc/DQkOYRJVBEd1ab2gUqKGMciHKSpeb+p0gF2IJgye
WwsQGJa3kakSEiobk+skUr8y6oBoe6GwikMjjAd4MZLI0H6vSN+4CORcmZRTfvqe
IhCu2Q7za/P2t0Igyvw7YzlunLlosVlf2DLAYeMMvEpCxvwRyE8z3tXO2DiDbQAJ
KbudIIDACHVeMpDzUMmZjAviMJA9C5Kr63Z5uDc3DcpHW/E0lP1QKO9UDYxxZClJ
rc4B+rr457tkmQgiqw/jOmS88nVWfe5z+PyTRMmQSvmJ5Ix4PeosgKaAzKn0fMeq
I2IgE5A8pqEIF5LDT8wxmx2lmJ6RFAQtm/NyYb62+wQsL50DttFJz1KgHemeAhAU
NZhyZ499cnO4BdwazCvKclCSfM2BW/oUcxT9wub91YsFTJfMyh6CF/MiC8wUO9pm
U1HQVldSx6vVozsgfdY4YvMtoFLvShINzr9/wYrsnyJXOh2ARg9cXqQM+RAM+/QG
mSqf2YFrNYRrt3swl0glVQj4QntaUMiC2OXuz70/5782hJ3OdhChF7j9uUMbtlPp
VhTitJs7Dbl+xANZ77+cGBMLNsh+llHS+YeXjaJjtri27oXczpX/HfQtAvdu6Fed
NdNJ1wlYwTgzvO0KhPP2fLQmAfZk8WLuKetvgbpg+ZfK0WmGLP92XgbE5Nk4hOL/
nUF4LSSrGqu/gN4DJwqn5gh+X7Kxlxi4BmiltNDqCUURLXx+CXSG5rNYRe3QVXqn
JDHu+jKKcJO/s8RQmZIoyDn3RB4UMQB/9zzHnqs1cQEFtdp3WbqCm8hwSmqnlw5Y
uKCvP6WyLQMWI4k6ggK1RfWfYlfgRFt0YGP1iQ6uysDql+n2UctDRMsPy0YepyGO
xnKw01UyfvDpgPuG7QF8bQ5svj/06PzXvyJLwp+k3KTYiVpkopWmPBy5QZYA4WpX
uOQI033U50IwvVfOZXD2TESB63G2uiUaTAGMj4tRZZNOP+UceiYp2O217t5FBzfZ
7uuwL3DeApGRMKEEOh+uN0EDYB16Hc2oz3AfpFrrkrsIrd/04ETEyFIGCdqoqmEc
V8Rnfxv+F1tObSzl6pkZ908NsXuKAfAKO74Oeoz3UHoIu67E9YhOGc0vyngYZpKX
D0G/dILpvxvKQgp8B1JfrgxKziSEsTJOMGlAw/EfQ5DD88UrzXmGVKorzzMlqSfI
w/8SDzbd74FTsA5m7e2I7uPJwuB8e5kZz+bVNAQ/UMw+LwMopgbESr2JF3fBCply
fRoDbNlsY5r3p26lQSleUExZf/PJmhtAWEtzcBh2+C0GrCGtQdbx+Ks1IeWQn3sW
Jf5UECvOr8GoH4UZUCftMMRUXA48HohL2n7LpJaxO853tq7oOCSfdY8bIOPCoMk5
PYuRw21xWhlVRSbaka4QdsNC9v+c664Gnbx1/jGJc3NnXUz6lZeMNZwHIt3RpxRn
O+avXz3y7wCcXliPuugpFJTBoFJaZQBXk04SMNN5yvYLaFzc+QlnF0yjQijIMxhI
wKzU1OOR2ZSqJdA1r4ri690OFxjiB24Yhlzc3rK/muH2Dfw7SqoxGqKsNmU7k7IW
f/q//8JnqmbkCyKy0GWktmUj84GfbGGs5xxpov9/dJrztv5cfNA5KdL+cmXdEY+s
WwzQQ7Q9OIxoqdCR6tcz24FX5jNFje2y+bBD0a1mKy7EWkZDKL0rjrPERA1sJJpY
8MuJc2a+k4JIxuuclr6GLRnXs2wtd2jg63mgajSwPuHS5G1kUghiYR4wt2Wl5A4k
8sIeG3f1iN+hdF6anxJnqsCVYBiUMFcai24y7Rd52IzCbX4RjbkKnmHOdevuIGDg
ufWTmiVKscwQPUzQYgijFQdcpTaBpvFpMR9/V594KJ5N34IzTco/tUu9qYNR8VUE
zCQJt6iKKX6fJzRmFzSaJMwxEvU5LKCwDipZhz15DAQsLQwBN4BL/BZgQO8ayMGu
ZJC/3E5OmM1iWOVo/4lvunat0ZV68cCSysYfV4jVkbRV/TVLE4q0D61VGFoVL8NF
HazHvTcXt+z4hrFuFhfRUrOvjIIkpqi/LzUytbJVergcRm7ii3bqVc5XY8IH4R95
hpbMDND/m6dl1XDAI614Q5moVGCS7Lk01HmEiI5p8IfLkDU/RMA4RpvKLh7Hv5/Y
V+wKqan7yUCTZIJh46fPHqP7KPSowXzlcnrYsW/Zd+UTSqLdOMlthP4D7ha6laID
fsnv3N2AK0lxPCvZj86GB1vlJNdA1qPAXUMZ78lB+D3huwItP3On5iaQzNL143Su
lhJlF6mLeR9FY++C/YjtiPuPk2nHH3xWEY7eO83Q/WJrbtTWNIkyDQLcvwSLh8Ck
KLyLIADmW6KlMwtCoZgTep8X5yBnwNYGEz563UHRjASlCo9qVG9Edwqln/houKP6
cL6V17L6w0ttLlrCbcTmdMwGMSGI5x7AdMtRvFj6CLEg3FYyb+jMmxtPc2ruUbK7
TUOhTrvXikQqQhjVns1XSfg9cmsyoj1j31hDfs8bN7ni1vWiJRBB84acZYps5eHa
sAaYZfUCCD9LO/vzrgA1mJzI0VTDAzL5kw+vaOIcKpMCppEPtlgguX7WKKniDtga
/fN0U4jURP0nVwNQ53mG5QIiPnXQ18Jdd9wSV3pGjbdAw4op5aUzRVFbW7/zG1KX
Ds1g0AsaBHCLVmzyYBhVCNL4ccZOMHMc+AkWlA5sHAzK1SA7XAMf2L2uCWfBZjM4
JCronjcrJ65aHnwjIqRh9vYPxxODs/560k1TNQW1ds6wl9IEZhpY1gCa843RUTM6
I0k2eWKW07+RhfvolKudRS1UN9lWQEcpUAdu5nDGbqQQ+GJB/HR2P5uhecJtK1gg
aBW86+9v2dEH//5B1MfPiMY+Peegqidn3jEJ2yfAzoVwnvKYzYbgv6px44xum4hM
v3MbjIClkHEmsflGO2LWXVKvXiSBNn1w2br7R72xjcNU/tFgF4UvZkNcZe8CNnvF
eV+JRDSZiPecSYZwAXWVa04Uipeok0uVii5ljIMq+D6UwD+PHpde7Nlgxx/OosMq
pe921sKfD34qXUmZJX07DIvmbPRRb3r1wLmCh04oSxVvsBZYVW8XMICz03vxwwxA
6CTABzdVbzE9KB3ClLieJNwfWWsSKYbJnUvx7icyZuZunptZxhgUD0eweQDTuEiS
Znb4f9u8/XEXjQ9T1FwxTUNd9kYLXUt9wC0ohKNk0w9PSL/xuT5e7b7lmSIfb0KQ
VL7BCQlzOh4VzLI0adIAWJUxmqnaWhfyo2N3YK/Jm2+yEiHUrEPPPES95ALoEv3i
DK+RkM758v7ERPJWheWbIJ15WVWSsQut9VUIai+aXQaZsWr7cqADokvuhu6vZIO2
K8JvfzOtsm8wB2xiINU/DFsIVJoIEGT/oBoGUvHmnEFcDfhhVFX+v/M8lKvw1wez
4hZGmO0eElJ1gR+8Xs86dEV8pLByjHAqC32R3ycV0p3WbxhFXIVcEFHJZbILTJ3g
XQt9XrRGTAC3d/H6C99o2wNizDJf/B6KCxc7OiiuKHwgVZALLaqO60n4+1JHmUgH
EfMx6LaDNtCSUdOsJt3JGAkusdzBjuHCJvME5Hx4TW+k++gcd1g50MxTJ8tb625A
s1j09aLYOr3KHVFm9iWcRQVIluwhZRJ9R3suZXA3K4zmSqBvq8HaNG5fpHRSdfr/
JQwsl7yRi2xBViXMRtycMMM8woFP1hSoeqDDcPFFuRL3Qf9VZgnjaVD/RGTEkPZP
GcOS79q5Au3p0OfPRGJveTRUiqaJg3FN7yZcuNfdlM5kaee/MZN5WWiTldmfMIMJ
fnewRRDtfYHdFQaJDOeP5YpaTsvQ/j/1FyVhXovWL+qqjduRlcJj3KbbLOzk2fvk
lJxZop6Jz5NVy/vk5Mbk6BL0x/idP/zEZiJ3RhXEgsLN/NGmPcrd28+AvsM/lvWF
slpUrug6KGvFauwtMFO3qka0vxKrSZE3iMBbzLBbtSA+rnnzJTqZY+TqJQ+u+vwH
nuR3nOlAzN3WbZ4g9sI9TvJXZHOsg2UUQVsV5d0HKkhZFMtYU1xuryidiNf4aSsC
tuz+sRtgoSPrUuCBmWMdWfEs0UuVT70BKsDS+iOP6WeK/d7BmHeJH5dvQ6HX+ePf
QLMarsqmjwng/WpqyonWDOQmP3MbcEgZfUaKmdSq+aBSVlqR4XSqmrh9tgPT6WQe
MN+X7c8MCeo1MHCn6Ng3ALGSNFS8GOKOaGI6gD8f+50kMD0znM/bJPtas0NQo1F0
5zzUNpdT36JL07JJHQIzLTyLNorKxEiJMlhYN+dr/iIN9KUIaHhiwU3RyOZ8VNid
ZvOFSyMvsxZVX+roiATY54DsV52EqyBYgu5cO7LgdVAjW14Zg7dIYQchPc0ZjlVD
+QQbfkDazsku3HRi9uarPqSqOMZpeJcOZn+Ro7OicQ3KqHPIVDuArzyWqgwc0Dkq
lrqWhFwDkfTsGAi9+q3O1y2f7aOE4ltwxEb3SHcA02zLikIm/CaC5JPuH6V+G+IM
x2UtJWTQhHuB7DejvXm03MhUpG8WPYKAIHKSH0V4M64M4c+rtz2ZhtdRGz+5aYtl
ODpzjzGM6TAcFFK5vmzMrzs6ynYsdlWb/7tL8G77hnllz6Nmr00Nx+/82jdkqcta
kIkdq0uBBmI3ej3eumdkROnnZEqwCHJYk22bJFSJMZ8hk00Ef2j7glZSg8KueX63
DwvZoGtOWdMebf9YYShQWg0LXZdY9i2UOUognP2+EXLIVsCztPGTrGPqcZwEvsHS
qCGjiPkM7Q+/Tkk+bJt6blznQ6Tb9TwoKmQ40ZwMq/R/iKBxwrmSLpFMClvMaabB
ywaBtRIpMf1j19ZUQpRpvElri1CVJx0nvEmstxc5OuZov1jqqDO1a8N5NOd+xdkW
f4jJay46DcaQqFV4kvGpqRk4iC3cMgJx/X2npmFI2GVVhXwcAeFB6o9tcewSn4hx
+m4HtSVeO8x7lcQ/6tdfs6ZJjruiBFww+dwISpMjzJOOZu/92bmTWfqrcqVyNLnC
PrcG/Zk1O2d4zSXRhfwnhA2m89lcnCEfW2l/5hn/cOE2D12Qt+GAqTGb8Q+yC99E
k1R8muXbYM6rhJ+C+pIKobCiGYk3kUwSG1a8ydIIH/6ZjMs9moiUW/hcaFoyQjvJ
+Y0D8h5F/yvzmIQyOSwkU1gcO/ICt2Sd3wrKRoA8hRgKTSl42wFK9ukvnmVBF/el
8/S2u+OqAvysg37vW6EeiC/eJ7rE1MxkGNfIzRb/TDQjxQ9nk13HJXqotfqG+YvO
EEWJzVpvs5UQ0FD9Djd8eQkS+XNahOJFawiSA6LOp3JOX15HANdnI9OB6HogMqke
n8FV7/CzhMSjOmAnTuQ0B/jPb3oMctUU7tZ9WlNeBx5zmGDK8TX5k0EDxc7MQqEX
dYurkwpIwxvILD6ydWvPcP5E61Kpb+KV8Ic/PDs8SjkXyEpyb1sY5YLMvdyEsqxH
vpdqdNOvjqW2ndAB/hED+E3jmzgQucfprCeiF4FKuMNJMJqzGb3Ugl8fgEY1eSve
efzqYXGAEhguaJ8uDQ5XYJtL1u5nN+YDfEaK5a5s/D0uh8nB1mvm9xFQjRLZH1XD
sh2ewYi8yzYYLvE/vGq1gFShLkRm6LKLOk3eMJDgGxbBSbQMNkyiGEXYHuFv4UGO
aAn3mVMsojxcVxl/3apCMqa3bXJDe0fjmeS4jdsHKErSFDlOD6agez5qtoO3cxxn
mbg9lH/h532mP1dLBdWmqxoS8Oir5NgpFa23F5tUzOWolqHZYfgLEMl1pDZAl7Zb
I6oRJQCkg1xt+Dt9XhZ3eywqgfGrFm3nsX2G9NvrW7kwX7UPf3XU/zfRzq3JyVl/
2KLqeWJhhLY7xFysAKgGlRBwTeYlctHGl5mDTmpegv4vWzXtELa6s7SeZC8Aod5I
HBIu7vKpJXkRG8di+cIqL/cnZQZ+HP/82opNmei1Rzmg2dakJjQPji0cgWYnOOLg
gYCVllXRpriNW3eyADDBT6bc4efn9s0HWlQlkNqcGR3iN23c7ErMMwlXqpWKrfNG
Cf4Zsn1zuAKk9PX5s3LJNe0h5IMIVO53hr1+KWFNYN9jS7LoYhx2Kt0lqYg/AJCq
n8RWOVB2pcZ8uRbr2HY3xksnnIfVwkXJOlp1qXLO8q0tTrBQEbFJ91RRqQiqIyv9
gwPZOLDJnQ2DnQ2xeIt8eSFnGI5fQjrPx9ZdYVW5Z1y7sRB7eVnn+/11FPgqa77o
mokCNmiEV4r8rPpJM0H/5HPoZPoeFfGHSWNwHEZiJWNAlvh0xShH/qM9fyCcVtrg
5hprcgB01nLFqAqgeirDejvlY5as20027vYrhXVkJA7WawhUeEvl+LqGZ6M93anu
JsyVDCXLHYCzDk+S5CFQzeZVIbxTnwEIKIYBGUsnWXVCYyl9Vg/FYbzzFSjY3V3s
w9maqcfus67gpuwLI019eA5r+O8F+Noesqig/811u7+95NEhzT4tL0fmN7zAldJS
fxoW+D/DPiKUjzkaWryIlbUfgLuDUan9VthktmlbBiqOsqNxkqs4i3rxU24Noc8m
Et6Q2IyfZoNlnsJYdhtCAbrkVNnTi+NlRvxrDsvVNKDySmfGCogBxUi42WPv1du5
gS6wvkm5FkwD3n8TeW9xqEQEut3xJTq9Zm/dVYsoFB1NncQk42uurx7TSFhLjYlL
UhjV7RGkKCe4fkeF4f85oukCb+yWtW+nSOrvrcfQ8AQoFqp0OR4X6YL8uI1JRUfW
hIxAACa7c4z9C0jMe/GuJUDy7f82BEFkgXUae1L3827VGQU43cdaEGeWRUSgaJuF
XQ3IdpU5DHt3OghQhClcnFszZaFxbAsqatBeXcxjDG3jceGMUzWKrysQCCWEIsJU
V7Q9HTrSKWTt0RKUCGpLbjttrShDYqI2Tr1+JIbhTaXBGLugCPBWnxtLZ/s7GFYo
xkT3MBG55hhPUv+gKLFrdEoyA8s2kI97EWJiSesLoYSepJ06aAAY6PQ80xIwXyKj
pKu2ai7vSsx58hnw2d1IyobTClXX2sYr6Qm9cjdrYnxBaDwv4m0hKNVBYr1jtZ2P
AQUgcayRas7c3+fFRSTFqBV3IrIZMUhOL8zWZkP4IHMVTKzaKBXtKtWROO4vJgQ3
xB1/7WL0taQxUffhLEkq/YpzSlCMGiS3kn1urMZNKLwrD1gJgqaAJtaALeycB1wc
ClQfpWFUoNXmJ6Xd1oIc1GxcixNBiClMMj8A0tMC4JEydNT8ZVpLpQw4EzAwIr3p
dfokN4ikClS7NeE+DRTAI/1gvnAzF921q17hqWqRcZ7clwvdhc69LV2/PM4CgQWt
U+q0Xaw/MBsRZgjQVxoP2699D4kyZZnBteQ+Lh7Oyfg1AAQHIDaU70H18HJmalIp
lWbLxH6WHRd/u8l+MUNe6HyTySiERGV0dIKctPtQGlp6H4NVpzEihjV13No7GjKc
BCQsF2UU0V9TG94E4zwrDF5yD3LJQKx+a5EZ+/krA2MKWsdXgFl4arNMRD3iEYzH
XFvuWyC4nedPN3SuJiPHnNX5DULW+4eABYfD5ZDxwUhbGFTm4yLaLSoXVoMY/Ra0
BHgkSI1DuZrz5K/a0qi2ciLieQT9oXzYFN880+aRtGtqGK5lLzcqmE88p5dL61qK
RmLXk98AIvLGiY9RA/letJuSrsTXKs9FB0fPAn788e0Srh1n5C29QF5ZUFQBHZIQ
pZKjHxg6S3YlV1Rc+o7XokPA+Hc/eZYLDrVkqm+GO8sNmI34fC8k97eqheznaxmM
dfHvRfhZ+QETKcFLPU/q3zprRqCu/keOzZKANbXte2wYQxOtJS3itsluRXYCkBiA
v5y9plFD14j1QnGdFsTi9wRN6GiZCinw1NRokDRBvckOr1myFUPYmi8zkRTDLVKO
+jhAS52J+j3tXE4g+MhPihpvK2nXYh4kCP2PTaa35iuW2w1z99KuiQZWtCIs5s77
cRhtyBM+Jxd3zxiDeowdo2gGipLOWQTDBSIBO2zthUAi012ip8oILi+e/cHD0RCC
vSidCaJJXigbou3H00fAZNQjlhea3OzEMK3ZqNWmf9P6WfsAC5ODfpQgfaJnMy2p
wjMU6M7euU39rQ15VJ0qFx7ee9oLOqvAbWHsxXwXxMY7fBgfmESSALK3JzInP4WG
rPQDyzYzp+8y6oSBqlNCkNqQodkuPo5KKhXB9pQuHQ14kLLPO5taHE5rUAngPYM8
c/O4yBwjvr0hksGxTcno3QYkOD/k9bUPOn48/T5FVqzZ8CK4YRrh3lqXuQfUcAog
2SNGZB/XhKYOwxfcJVzpglgZp/P8kWXVMQcafFOPi53y+peUns6z4rkHVKoFspYh
WEResvatlGdevtjVBCngG+UjuaEmydZKRgql5Qvhau2COQ3zayTHlBYmkG6FgVOe
Fe7Lkya9l0X/5RBe6m9DvBhNuFbLoiT18Q28N/0+9R8o0P4ekPhWSNYwPwrUZygF
G/jT1eOIrSjPJwGFE+b35cbGLwsjMbXnBcU3yquH9yCsQwEXd20OyF3Mpf29RpiI
22d7MJMtqXRQ6Jeiv5r/E2aBZTEnh/Jmyovq5TJoqaFk6nKByy2+e7fl/yLfBTne
+yVZEHwlWNjLCq1iUdSK5P4Z4u+DnJcakzWNc0LlQti4X9G+lbnO5uneT1siDJN0
8W1nNWNC1bsE1Wb49iKlDLh3OAobNIEKiziErEUC3sugjrbLxDZN80rzSKX99dkY
yzGPGahAn9VyoSzEZLXX234aCJfPcrgpF5dQezGvW4z21gsOUG0spAJAPRAhIzW1
UzOB9CuqwLo4+3odMrkZNZhm7lPtfJwheK2eBPRWCBOA5M5dWygGG2SBL6Kuh6jo
kkExQG4ZyG8TJOJFlrl+jpPlc91HEEm7lkLctMctXm1K0uJ5MwT1HBc0yDWlu7Zk
4gzEcd35vOiV29QzWGn+u91U7CQoLDa7fatBd7oN3rXffSeMHw4Ry6FGK7offa1x
K1HjXqD28u5RqzS9NX88KW5nkzfenOPJa9P4UcZz3yQDh4IcXon7cuz70in7J31x
811Z/CYjAftH08I/ZNKK7YiipoDJb9dV4d/WRONgXscUg+WTsjrXCecQK7D+7oQm
UULrsgkMoQ23SWN2E55mYh44B4EpnVnLe3uHvY1cG2krBlWZDqVyFXYC+9EdWq2T
yhGTusyuToE6lvDVttKzXsFtMzQgm/sJKHPrWri/pub21iZ1mqJVQnK3K266qzpU
DPnNNz4DhtjbXA59D6XC3AcwyB/EokkL4YQkp6NibXQaqVLmrbTopO2nkpC7usL9
PgzUPyIWCWR+/0hSfAYfns7vTSz4weF20s1s55TM0xfPSBv8GWxlIfep435r/u4j
Lr1VZxhxW258xNSBXXUCuBUt/UZ2YkKZfxM9TneMVFekEMQdY7RY6uzMoM3+iz7s
PIJ0axTw0FfvOwzSssJy4g19GC0Q3RrVZ7X0V41dNrM8jFAg5luNR+AYzWjmmlSU
wvoCsO/aPfFDaRmkRbXuBN8EKoSTDnj7r8OnqBvZtyOLpbvGHZsw9+4OtqkfRNVy
/yXAEEp1ordMQQUz5mx6NH7Zw+IovwE8G0vmd1An9RRgU5E2CoxScoksPvlVf+JN
KLgGb9EO87Q/mSRpSTryW6H9Af19oVlFUW35ekb0WaVrVQhiFfZDL7fc1eISuloN
ZF6QYAWgXpqyqSzkqx10a3xQFGdaPQR24I3Pet0C/oUn4oc00Fhm9dTl1swGLDnW
GEI9NMevKzFx9Dk2aOhAs3kNstmHuTqFpMY0iQchv7erZbC4FsZgRiljegJ1MNbu
DhrhBgaf55C2EF6Qe+ZLhJ+f3mcoa0+FPhpvCy3tUzC0IAc1bjrn30Ic8MoFimXx
bCRmDjpuqkLRJqC+xVAJ7a5Cq42qsDwfaZa0p75EZHiIJqrNz591cBbXjWa0VuqG
pgHmweOx42lahpcRO5jVh9SsFifk147DiLxrngjw45wdgilif8JTZeWJGx0zSgEn
N/XDapM7+/LwOBXvFDZ5NR1rKyU1oOWGi9q2OhvB+Z1PmrhL1vFORxIBKP6tqbKW
u/dRgSGyeDSL8tJjlyy7UsmQixiI3eBAdDQFLetgesrQAYksPwyUV8k9kd0S0aLh
02YDsYP9LF79Ebgjajhy8c3odTysQ8m3uEY5VLriaajRaWbmFF/U1JXkZS2wRX6A
QcQ0+aUYhsHwRbp9l8HulOWW9SNl/kmJjbEFnyV0Fwt+WgCRkn9VpE93EK2IxVRS
gfw35xWOCPloMdmDn3G4M5HaJTI/7QgihNEOpvK54hOXwJGxtrS392oG0tH0NoPt
wCBR50TlsiQBaF8YFPoDugFT6/xhvZNk1Ktiq+0n75usR2QqSh3oc8TIYFKWm3Wf
4H2UfylT/JQZlZT6oYRoywRpDNea8ee2xbzLwm2oSApgmSOneCYrS3olgiQGFikj
cfgfs37ANAwqEdfLttZuuF5W/n9l3TmsHfoOuEu/KY5zlvGF/VatQ72MTXuBxFnX
SvWgEWSCWuW8nmUV0BvWyhzYkKzIXt7eyt7eBaxxkn0fIq9Jq9s9xLffH0b2+Bke
RjRS58cmi6Q4QwLzDxNaxAjpAAI2c2d4z3a5A6fpMcY4HmZW249VoKfGjKJoremD
ba4GAqrlsfEhJLaCvwoP75OTh//N8f7RMoP6Z5kpKySA61Fyt1iYAPIL2GgDhVNF
oCxEYDeA8oMFRJtyZTG1aPh0pSP2uKhNmfM2BpkvEg9wl4rV+vrDiea+rE5q2AcQ
W/TnUD15SMJxGSD4dkYuWXDKdo373dOMfpCOeUnwivQkUHJ95pbcnofrmOJgnokR
4vt0Ij/j9cETl5I6r0trrRK8lgzjeAV9rT8QThW5wRZnhW5eEVT3dnK9zAMEeCzf
ZHyXqB5IsQUOMQeFKxV4pzGvJCz9hLYZubI4jhY4n9zw0Jz51hI//KPBh4F90iHT
jXGstWBYSZq8lSkE3lzjIn/I2ZavqUGGoZ6h7Y++6pUPfCKGKr+x72Qce9yqDprH
BVFJJb5ZNNKRHTjMKf//8Htlcpdoe7aIMtLvgFuiI6c3RJSFzeY0gSUDW+qu4yVA
zOvcVVZoYKt+ntSVe35brXpcJ2WIs62CwdU1GNoQ9OBDGwkC/lwd+p6ku0n5kPkr
9GaszOnl1OfUy6gAvx1N+7PsKRYFNYdAiM7KSLnZMRul4OG7kihCi7B2qNfayXF4
dQ7rDDVL4ULy498Kpbwnq70NchfxtNWOkAPQbLwneNDlg+ZUzabT2TNttgUqoA98
k/uTKmPElLoipLyiQS7lFeh11D7ixjfsDTzZPlOCAUztvoIYxOfdA+zHmbxxwL6J
/P9a13pnMjQsdomCwujBgrg/DSXpsDcnyHj1jNOkGxOCd7wKqXm5hKGqPb+WmM8H
Zj4Wz2OKr9J3DMCL/iqAop5yGuftHigBAPx3PzitYItT2NdRKfIz0k/U/LJubmq2
KMdISwB3Wb4G+ADM+wSxZKgAnCrgL55qyXIcUADuKo1G7PpYOrpAIYA2LVb/MnYy
4rurs/eaDC4Io4FocBY4L2uysAu3E3FK+22ySeB9mlkIyZfrxZmGtD7bkuPgRydO
Ntx7Sqf8TMwyT2vJU6SRNEXjXL3YKfW4t1mlI11j07r1jnFPMaGTDVbqTLgMczID
WW5URUztHIDJtFjP2wuqd5dljhUyQCjtwdhs/XfGigcc8xPcSh1o187Zp6xs+HPL
Wy8UAGweO7zHQTwKhscb9yPWSZt5LCNP7VlPvql6mpAwiCE8ziAfGXKK9mzcerRc
Oy8yeC9qdtjonNkuuPnvbgX1USVTeyHEJ70jeWFT3UR6JWYN2La/3X5PXcHKnNad
aH8qrFdet9mlpf6MipK+N37qa/T1M9U4q/r7ItXyXqaq2SZlFCfc8LWkrCNeu6tj
mnmY4ZMN3z1jxKthtlvS0O0LZNFnByofGFI9Bmj+JSnT3mBfIiU7j95QGVuoMzmt
aO7pRdvgakZa2acPSRlpPoDXEeCaoI73DblAxE8mmKTEEbS9WQoF/LHYpsHBQAHi
4TH93M1rByiLLY4lW5r8HB8VX93HRBr5sBq1Ik6nv1DloEUNJCmhpebL6ngZkNVN
MXmba8+sKPk6grtjMNXvQEuSY1d/f+p350KmhdR9mq5tr8OHyFbBolSEPfz1bDcC
gY+yDmEJSz6vVzMry3kC4xe0bACdP3VtZmMXPI7ArgmA5GaKS2Traf5qzDRAPpkq
HGXG06H5zFHx47rPhvqCynAQP+cI+EEWkM98LaderlWijHQ4OG/2DUajpuEarcsj
R5bENvp1aRQL1xk6njtWYHfHJJHJ4uSdawfWnvXC20fldI0tqhKeORgM5l0vQ/Un
KAfOIpLNWfTQQjR0M/5b1FsE1eyHdiH5iOtkyQkcek1TBQdiriMsJV73/RfD+pHw
z1ayJ3+0kseJJzmmXtBVhJDmjkZAZKpuW+NeZW3Sf10XW/DuPv3Hh0+jC1Xj9haZ
02GhqxLQh3W+nIa++AnqR0vTqlDcXVfMaFGyXvHp+sKcr05E+jd/nGh64JdSar1l
IrXd9gRqVGz5iZoA8sAJkLg443RSW0k7U92gVCi+h8RzvB5CYswJIC8mpK30Yg9t
Ef0rbEr6Ix6PS1xRDNcKjgVtWv+46pcyet7cILB6fooz2iGpMw4OP4aMJ0uMA0aR
Qknfu3N7YMzzB8Sk5JQ/lrYf0GoUVM7sDC4/TcCtl0AePSIU635GraTU/VhNmqsy
F2/sEExdQabf5XvZneunUMz6SVZhKstsYTKxrRvay8yJ1EAuRhdUousA91lDQtiz
6UF1rXGy1E6vY1z+FN6A+8DvETz/7f3tQjKG9YAC+2n9Xmo6Ks/cw9GnGxthfSaP
29GCjT14sw7BR/G3xkShNRGoQfoMWozdPbPM0b20SvgpIV3qtDoCpUm9Pbnfdure
qZ8sq4e+L6ynMZ2+cwJS+q2qVv21FlyVRQyGd2wB6Em7J17T9bzv7vp/JDmzFJ3w
RGRUfK329Y/L8VfGZYX/i+ePCIaR47eLdn+Gib9tmr7TTbSGAruiuweCTPt5LEFz
GiXjzhdKu2za+NbiNwsHxOUg4tGtUbjHFnCO1EcrVx4DpHy44wzKNNOHDKR8Vjpm
O/mloaOBlW26HVgNQgS+JK7dmaDbvfZhoobR/AE8VRsI2Cm/4qhI2DSAcDtivjLc
8e2XSAwnCesIPYAPkyxdvjxluGJYDUmC6hTLql12/BnhrgirFAfICqE3EPiVxyKC
M23DZ0LxQ3KTGm7UInT9tlkpQDvI/ecoG2jd5BDQ7yCeYs1zjr8hXg5st69IrUke
dqzq7j9XiThfr6SVoTbDNlAkDQCflDcGCv3hdVVHZCuW4w83hNrKGmOtg8tsGEu2
uQA6oDXkIxdkiyCRNqbKi4zoipHtTT2IJFkhhxMx6u8sNffx9Mlrj9Jr9UNHtKqN
YlM5exPsmSxlE/oRcacwcdjkhYpWUbUys6HmygZk697oFtQdl7NhlGVSY2xgJFRq
I+hz27bvcKRcuXGoNW6+TtzHZ+inmBOfTWLR/a4pe1QmwvqPykarZ62QNpRrUUBM
uXhOkYS8PHBqKQNDDYUA3tlHPbNsX/YlZ//QmHPBSpA3m5gStEm7EciQh8SGo242
F7jDmV44KDypQ0qVr9sWda9STwlmHcO7hQMxSStJuiJV8gjB66Qj/ZE29fddpjzi
i1kK77ufPc1YSD59tUaB3Tp1G7hIF8vJ4PnAGWsWHlv3OiSlnSz42FB7isnAYaMC
2cj6BU2kyfCygGuytqjtodNcvxZLOKyVv2+dQXTGKkV480MjJ6e7bVOwZhociOf3
NjF6ck3OspI2vvBBwAHVZMNkoAEAe9waLI7NnKD2dpkvP7LFcUFwS3RTvFb0ErEU
nzEX07eb/OlLVv8lF2Vp8GuKPlHRkIGR9M2bdijMOI+bY8U1eFuw0BeZfLs87cEu
hIgeIE+dffFoFt/Ms1glUXMYiFXk6OlSEm/gVA62PRULS3pd3ZvkoSWCMbylu6px
CfDJkOyuur11zj7siGFb0HU4PvmBjj9QHxobcGEUWannkCuP1ZvHk8y7xTOLriDo
8SJHU9Dh/ECO0jA71arFu+LdZhBEGZ1iNqXoNAtCQhBzp655YJ5LVS+CpOcdG6Ee
5l+tlOJsq/M1882/tinR90hl9Ipgr/ugNLofUB1iejJtr9DMdRCB6eIAxTeBBKtm
YjlIsmWrCb0Ujx+9n0RyXUMaS09r6TNQO5OZOr5FVjF+fIyzdS8wN8DZ1okk7JPp
312n/a39tse/VTTBy5hSaT3J5ZLE2fHMimdGRjGKvSJkTXrgsYQFFfd4zoDK07so
oP6Od7/ccC4388NsdrpLQhgL1mz25YfjzwJB5tnQpFkg9/J77CUhAA62mx2WA6xV
arciWnjbOBZ1Bts4fkUiTTAhlEAu09GEUJHbkZEnGFqzS/tf1oTa7MXu2wyebn70
GO5TpyqNzR5Z/szNayZR4mbsfsQ6yC+YWcMWdpl83TnpPWtC/BJ5LJox2/dzynxP
1eHUQwb1YSA+lu5DU743vXbAQVehQAFAL4WpLIFr7mpU4AIQ98PDFcJip+Z+ngeT
dVW47HXgkMMJOKU+cWKfjgA6BsjOrN0FfkL1fqLxdvH0FNNagyzWxGLejuBC1QVj
QDOVFCQ6EmrX8SHswGnaU/xrNKQTBan80KFhIjf03q6JULoJuhoS8yzuXLdk4aSk
+50BltgiXhUCMc/eXaSIzbhYZXHMJN148sll48xiH+h6+nRRVHlOewzVMwqNLwAo
iCw1l2K91bqA18vUpShzoieQWHKPbdhGcWshjcTI/e4YEAFfdIFxyVAJ0bPbP+jN
owHI6JU6UPjQo38UVui3ksOZHvPurOLPKYSBVX9xUUU7lb+Hv+3wgAgiuD4KD/TQ
MvbAOlF1cNiK+Rnqml61mNeto2+RAAQw1ppJkhL1kkX3cnHjaLXMhS2Loc1Wh00t
qwkYPawYvnjdP/sq94xzs4au6wXrM14e8i7Erb8MlRsl524yLSDulw92qsbkgTIQ
KJnolEcV/sUE5Wh3JUAMGXlG6w6kspw2JoF/bPoouSOmoph8BOvHJNbysN7FozPq
IYv6MkuS9UIW29GkN7r54Dxxz/AJyqmFfkepNBnS6xwLI+MUifb8asrnm/NZdHGR
PwMX9z4frrOK+FmtglMny6KJzXQ5+QVlDPaRBRe9dy1kp4OSlEGbR1vQBxCMDQko
Fi+4LDaUT1OCQTaw+Seg384Q8bPloCp7IBF6xlhNMk5QUR/d3z5ELphLfldHivqF
i83QDE61VyHYbkzIdKxJKPPI9pnl2kFErlEA1GIwsRJUn+w5Dt2yGZGRbqK4Nlbu
e2hTrbL75XlpKfAGp8qq50dSmarPF2fbYaRGw1466zGmHO8/c0CcY2AgeHU9dSDl
geHZbEqoNK8W7AOTr0oKyrLxNDSRZh+3Qw8MWCKmtQvKmpbR5+XcSv3071IXSwpe
1TRpPpYpISfqxoBvB4Y2r3RbrTjlqUWVGO7eXdbXr2ER1l7zy3p9ViL/ULl/9+Rb
ZQB6xvnbwhamkTEgRyv37bL4LbNGALEWKP50ZC1vRFtHil5KOiuL3/16oY3LZTbv
SLFDZPgwL8WcNGlaRnXiBEaxVhcRm3TiCP/SijT0tWoNOZEiZES/l+BEZHImOibZ
AlXwaikBYDAwGtyOsLMhGP3IvLRwsE7EeD6HVGVT8QHTxfUsU+JBTNiPDX+jx5A7
Jy4uFUkA6ImtGimySQHFlgbTrNXAx4jFmuplqMd6fWO0nSP2011/cbEXnAAOOmXT
jmyHVjAXwFpRLbpEt9tJtboesfHHEvlQYCqp35vTYapfd6urLzMv/tsWDu3uv/wf
0VZKXuZk7ATOdChlRJv+TE69ozr+S/gRsU9OzaUKPf6/w7lH71jo1nrDtpEbgRgV
LHJMeVw/TqrT6zlqV39MAOZcoEXjqE36kjyN4O0ZVnax4XBjINrYVggKospfLbLk
ZeyQ3+Hud6iZuoKJ9lWvOQzF8+m4Qk05s3JSop3eOVp64G9ikPjtpo0Kj3o0hs6N
s8piIMcuGlHu6/ZeEQ3iulndVxNCf7weKuMpm8NhEDky4kW4NshvshhZTL7e2LIL
R2Wj0/Kv239b9/be2ii0AdkSrqNLmQ9MJ5gBQNxdHs+ScZz3UBj4uKj6b4gUTbQl
Iybjb/Gukjbh06chjcCtxhyTfbkbThD0OdvbNODa8EHRK1Vcl96amIpoLqwjleXV
B/guim5u8otwYcqh/hfcDGdDhn7YIbw4jLUNQpWFIEWfhKvq394BVOwkLA4ss9Xn
KVcWXeebwjH95FDepk5vRrlFXW2yXQrsKjlt91n/EnrJxldIdGWKGWhtFkeabrMG
wZGI5PimEW0FfzAwpEDPaSesIc9v84g0oIGbxSiBV4E8WhghcabKQvDESWk5DgUR
Rjaj2amc25QonrSagQy9cZJM3qLo4jCp6A9u3ZANTEn8/Qp9EgSMmi/RdkO38J4n
It6O/Aq/YZtl0xoQHFZFZRJMuDnStPTCp5p+txJJDJXoW9L7YSZAYuJ8CxGE9Y8D
7dysCvmXdA3Z4KAXY3aeRD5tPb+beeldxmQzUFhJE5dKzMYSRJLhTAnJ0OO5ZBQ7
Swy9+RHUBL9ENHM1oYxvV2zOhqVdQhSCvh9KJkMOoeN3kprZF3fJUleKGl6I750S
5nIyUJO732LyJ+6l1zKe1q9FJXEO59E/ihlBcho/xqZDFXYmTXwWc7KvuANqSVHB
RgP2DZzxxrV7/MTAviVGy1wRNVeG0FAdY8l8zfEpJyBxMEwXl4Ad5LJxkqIUoe4+
HSE8ulnwPz6townONChaIHgP7R7s2qgC6mZsQV3Q5r1pMd31jukH0Do46EKGctI6
gKvuFfVcGLBOhAgtrNR1KcFf9iqIC4g+iDTP50F+Dw0CXrGGFUliNDYfga8yLW5Z
XHJfEHY0uio2M9RtYL6bHvf/6BdOzCIC5FG4m+8KrLqvV+4dmh6o74UXvDYWSWI3
1DWN6aDbO1+4gmCvo796TaQQ9jtTE1ERYbK6ZlRuSTDShlTy/vZTJFXA5MFyDbce
6TyMU8G22yYmrDX4TqdXv+dUL8naEdoRJaH26MkSjaqGsDSbg8gNtTV8KHB/zlmh
cF+BK4C0vjTmHmB4r7r0domlVuPezybNoAOM7b0qnDZAdBkEzKpxquWKnxMCui3B
zV+kmXCBENkqFsrPSpN0AxOOQ0tJo3YPdGiIE1i120iltTSzadtTW3hitlMDcfI3
4FMsC7TZLAUUyx0Xwn9Tk2bPBVqBx4I+02S3HTX+fC9zo2pOChdmEICpoF0BLoH7
xpG4Y2cLclYD/gdrdsmx1oL0j1zTYFLZ6TWDcE0EfYaCa3NA31wzB8GMxhuFHuc5
Nxl4eNAm1UW46gLaeBJ321j4lF2ayjfJ3RiAow+8v218kLDkO0opWtI4Iu9d57UX
u9ZnwmcwN4rD1XVReVepp09CFsRkCNesW+b9H4MME/4WZNK8tqePnHRixSrGOXIL
hlEj+p7wa3UA4x2lGWmdTbGlvMKQWWQXyi23ZXkpJL2OvYJvI33PK5Gs5iwgf3wL
GnUg0AkA7yPacA3nFfFkOdOpVMKgDsMz3PXZB8qB0x4qguc9z4UACtnD7uJRgA08
ed2//+Xa4s/lGATTpOb4bi8gELxMnxJTOAO3aqbeCM8E+rNB2G59VJVaxwAOKu/2
VQDZy4Aoejiw/KtroYBKHKPeS5Uk3/Rbe0p/yU6gzaBOOT455gCclxEf1j3dhdoT
X/Nn36v8GDC/7+Wuu+2Yx912taZkP4PWHB+rijxRIOBSSTggmnAf71sIxvzUJ413
xf+CBpQ1n+C60NeJojqa5rcwb1zu5HMCejHaJ1OcG7phC14yFluvlQKxfHmpJzlZ
GN3KGD0IiXyBr9z7gzetZOACTvVPCXg0dWvNOoiip1QCxS7am2I6mrUvhSDgZvMN
RdQ6SkhbejGrbadKvFWhA1iQQ3+RwxUFNJ7T5F5Yll+gU6wab/3keOdYDFV9Z7LJ
921mZqh4zMCty+gjKWKFiClaA+GZj3z4n0qMljlWalx8RI6pKB98kIWLNgJUEHpl
zRE1ciIilbXvbsZ4kxRgpVGRi1a/+r4C0YQPTSuDGi3OaMeD5aUQ0VGO7lJQ7u/Q
6hZ/E5tySATIkbL1imtfxpNS4+dcfvz5zZijUxtRvQ1UFAWHKBv+flQJEbKh2rEH
p9qhxi6dB89ljmzxJ9mXuHoFSL1T4HfaWgCFPfknLFaAML4bj1rbB63QNuvnzI2M
DXKlEVlDyzHYSnNfkscDhgLh8SBUjm91JJ4KYWKVQBnlSUyOu6yJZWMzIXE5BeeX
J0l8884F5dFKB3scC3ZCcwVT+9vdwPlACNMmq/Oe5RA55MFDCL8GuKvhXcLw7bLG
OTpNZZcaVxvGAWDPOZRsSe9EF8pD5FGCtzzjr9XUPKNl2BtyHWs+AfmZIyvjkSDq
hw5enpXKzBgy711FK8AmFuMztr7BWsDDNGTzJdRq7Ow6YInzKSfHNbZltI6bBqzf
t9/2UsTip2nU5ci1dNWI8GxropcRa3aTt5Q71J65wnDOPtbsPPLHsyhE+iYakDcm
/5ZzBjX9In9NoGUKyIDjXpuDw3ZBzMKHXcPhoLLZsjYCAcVas+Z3rbufWC24xr3u
AoB5+jHnbG586IX7ehWxoNW37Dv8AmF9YX9szuyUErGNs7WqKQQSCvjtTayCwkcv
MlSk4FajeRnTPKEgUVAanPVa5ZciHwNfqwq1Km5T7cR47LM/k9wSbT+bNrqFnIv/
BskBkprjf6aO9KoLoNl2rXCpFpDvRH5scVQJEptvjSnFOineI2dPf/K3WYQ8b/Qo
mW5BiYmSPAOOKUd05ViQOpTe7Q4ZksZKTMacXjreT3kCMqh7PZ/1F1P6dEm/M4/m
Yddfc6NAaXpCObdh2LPQF4cH9kuPR+yjDdqnAzquGiA61cFK96opUl+BT8nCevSs
suJ+2JPI5unbx4nScEaTb2iKJpH+Q6WTN/7yKsFBAsAkMa2S0QNcE9OcSrrQ7gvy
gRzXxz8exlSLyga+u6aIMDUUUDJNnW8K10SaSLkiKFD7yVHCzrY10b1XIZx3r8jr
fpiJNd68gj4qBtTTr74/y6dUsIDR+OJHV1Xr+AiRzDrumuW3NbmjRQQPvOJsGVLp
vaDjCxTDILzsrS+a1fRxLQVxOHaPn4vLR7ukV5UPJdBpLe2Ex4+eLbMFMy5GwC3b
cpZow3tIlnQb4grCPx6gn4Cvwtcw9nCZR4Bj038YCEHFLyJ20ko/yOeIXWNgAAIk
+bFHML//xp/t0jYbjA+yPDDvUYZX6oecW0VBr8ysJ1wYN/gLf9z2u1plDJtza7b5
AOPH0qKmjRHJIXZyZj+Z5KqFMiSV2d3bk+ptiQ3PIgT9Y5zotgOd0bwqEKJg53Q5
UgoWv5EVOHXUdwWsvGr4AG/z3z4rdQKv1lY31o5oqHvXjl/PD/K/lo9DiV4rO/xM
miV3b9hN8Sq/2JCKUDI98nTTPwyUcS1as8NPkXXVG1nFWn5fKqKRwODrmr/aXUeq
3jIZuUTm152rbuoHstsB4t7OsF/HFamjUa+xZeppX4N1eKGuAHBwnokYHzzNLjXa
JePGpzDT+qiXsB/O9ENglu56kDBvMmn76D9C67LUKz/zlnsHy7Jl0AA+8hXaXAOw
PWsfos9A5+ptBfr0YXpNL6rN2ofDBpF5AY2VMHW88osq29ta7Kwp6AGjdhTSVRG6
mzgcldlzISKTQKdwWJYVwzRDTaxL7QpnP8yNN3LUI5k9R7wic1KoRBmhlBG9nqOJ
YYvr7PTAt7rOyrKN4tduuj1p0bSRk0+Xnv1GsVMRgc9B05Oinx8cBxjeOLMBLx5A
RLtbKWItCjIj//l/ulUfe4yazz9Ch7UNTCzI53+8qLJwtKpLnSN4P9Ob8H9K9uXl
hGbYERrbbR8kySx/mmT/YoEpNY91qcKl1AL1qBLJu4fr8U4VpAuXt6z+WzU8sAmz
heJc4PQ4ZdX6zfR8QLJQCV4BvB/N4TQKJOVkrmWNhL1iHIHjPQtNolB+6Gq+G/Ke
ClKheOPdII6wh7HxR2RAbMnD+bXgwLN9Fk1e0cA6dJpX20zdwI6O+MBG0CrWoUU2
IWrAfS09bzm0bD+baZdxhoMLzsxsIqDU+G45BhX0dceMmZYOoBlDPAMS7V66LIeL
mmMl7kdmV84LYLgshZFuLmUfDpRZ3Eu0ysOZkRwrA0K03MSrsBaEMd5mdRsJuNwa
ojwc4taW9rRQu/FbXnKRtiSjZJNpDHLh+v4u+BjNxUm+ppvOxVa9FTmU7ngQgjWz
GDaCt/8Gf3dwGFUaDm8nvL++dWT9KnzvPX8Lx+dEgKbqWbLw/5BtRM4brlDYxJEK
R6ieOD1Fvm8OwJQLnKUzcBkEwdQ4RsZcteHytTz5o70diI1bwHPr4Iy9Dr8JAwz8
p8oMq4FGjs+TcySFM4RIXWumM9aeZfvhSLB40+2ZmAL6XlyCK6scXDDzcGB1ojob
Ft7hoFXkPDNdPcZ2s3JIxgqliCf3Rmu4Jvn5I2xoM/3AxF5N8r87IlpA+ccv3rev
T6/AQvXzyKqkGeYYyObD+Uc3yBO0rnVrorOJAanWWwFlJUUKZw7k/ZuRqx5WvxPj
KzdirQAJubAR1lNTP+zfAClfeSTZ1mZt3V3oG1ufB9U1QXLApRpn1WoOYd+OrXE3
9mhkYV6jzJfApanE5D3XcF4zv3vbyc868R9bfR9debj9wu/L+gBpzG887M+rLxHU
l32V7YFAYkMqJ2d84RJyxdoaioReZlDdJ0VrWW2wbmaW2FH/CfSgx3H3F8C7QMQ6
ftKtNUQ4g5m7g7EvsQISR5R75mk2JNjftDTjJpmHxla0a5zRTACJe1mTP6deyCBc
ONx91IJGM64hnUWp3zY8BXEPS3bIfEtipwY08Qiyu7mOsIO3xxMfCxJk+dm2b/Rq
IkFCA5LiYo1KvL39WL54wnRWoBy8YKYQJB58+0VsPWSbwLXXgrj47e6sgpyAQ/Yy
cseCHuQbvL0Sgad1q+7jltBjWtorPE4I+2ltRdAjX2DD+jCAWZhObxBoS3w8FEMe
CpahUBK4wMDJVisOzCJtEFZExlacR8mXPcqxMfnUVFlnuxhG+M8T5/GGWyzbhif1
LJyLmKBH0Mo7mj0yityxpKpbeH3rSnXPiv6ffpRycOaHbSCjtqpijMlEHybTtbqX
Djp8VT3Z5XPwdHhDe3RdwOBuMPx+04dUHNtoJYEKLOwuJEgvW1T74f860fOpOHBi
mPaAJ03OaW8XBBQg7PFkdn6DynHJDARfe1XPBe/ONVDFf1mD33+fZZUdXv3unY4q
YDq6AMuadYIvXCTy0ZYmEhUBK90Wocw7Y2pf5dl0hIx+SOkscrYx0tO20PHoMVRa
sWumHBmwecbFkHPnWYlfD4RMSevari8G1FFIaEZ4tJeUUVJYqAWW9e252Jaa0C9M
kXnTsZ95b0JCsuGrwBmoFCK+VxtG1GRvi9S8lWRhPghMuNNHscHVE1EGLwPbjmdQ
O2XuVs5O24MwBp4iwyfn6D/TDQ365BB+oFHGoFzFJryvd2UgV5gQLQLuapp0BIiU
+wBHed4hDK0HkCx9NcNoEm9DMuBoDWPTGJA7hGvMaYcl3tCy0VdvdlQyi87RS3jL
ijfuqFLQPiJ3Qr5L7CiDe9hOk3+wqDLS6GsH7NIDUyiqvY5vEGqvRjzd+Ud2/M7I
3ydGdrVRp7XqmlY+uxWYIWwrvIghW4rT3z7YZ/QiCW/Y1D3Bf31IcD6XNdkbWjA9
gWM9Suxpmld+D6GnmE+hznUipEeLUEo9jMjcyqqXApVEwCXKWvdtc8pxVOrqKjId
4sFVjxhGm81PzGB9ERQD1Ajoj39hxhKfYeeYjqOmFSnZuRKfMx7uy/SxNF08Ebiz
cfbFYKOUuE/bcUynHDsR1DPzcAGhxUZtA7uN19lKN6rDUCOdtRmhJDFmgIf4qhMV
ETCcq9ZxbKY5xAtCONxt8bQO3ExFLxDuX2g3Nqclrr+sjym6SXpISm1ouXIljlx9
XNadA8Xkb1OC8GFvDUQfdAtiBxpa23pkOdikLYkMQDi1EKccjAfHCZLHJUQSinP0
PQ+XATr7ptgXVgqYzKWxH1xWe8RqW3p1/oAIhAj8i7JH1SSawjF+dzQGe4G8+Wff
e3iMUu7vninPodXg+GRTVkjrcCfrIutCUwE0L/CX6frNECtuVhqnPOpU45a/HfSt
xRaXfz3dY9GZsySPHKO50avm48mGQNZE6tla4wLxxM7MfWxG4dkGM4g8Qn83sgVY
tpwFbobrkMCbVZ+ekX0WxOWpsPRYCgP/pbWI5LJQfj6/FmWPBvdIrXQR29ioGaEU
VE5SEm2ZuYNr95P2BOwsKZ7YqlYcBJUuqVl9myJCm9I5Du3vtXcYRbQoc6I1CaW7
vbHIA3C8OLcOPS4vpMWAMa8qoZxkphCxRP3Ca76F4id2nK6fDTgT2BM7y2n50JyP
eoi4T0BwtQxNv1cYknHqeDnjU5ZD9tyEXmNjPOqwzlS+2XyPRsECf/0YRNc5X/at
W2/ac47dxFRtg2Wv9//vGXvE8QINxwvIsv7NjLNzso+bzwE00Qo+Us3toTNtEd0E
x0MrK9xjq/ESmSu2B/4Pax+a+HxWDJTwKjVx52kN+UQ3IrJzMRvwOEqvBmVIJGIH
A7ViC0ca/I/NVDZAUHWx9eKLk3EKMhj/nEjfKy0VvfZiAgfAADgxCRR95dFk3NpA
M/Z5jqRAugc3R/2zxUspDIN328kd5sa9oJww4BI4ZMlcPgIyRQebnkhaeThls9Xj
8wRDAGuiT3LRYV3oCRcrDbjmk112wXnH7bcP3lOV/uhYM3FfBKPuIAowCo97YaRr
+Rf6SSr/8hX81FZyb9UNBlJeVzdBX/DBH302GJNWmEXvOvo4uBQYXc8U3PMipxfr
uuY4sj9MtSTEw5KiJfznTVybh5CyOq5Qxq1SbgujlBRPYg+f9ebPMLO/cefmz+/n
CvGE4Ds7Y6ALYzDjJaf/EA//7xGrKeMdZm3/5OJZL7AWftdKy24YqBkftpCRdc+F
3zP3wd3pZkor+4aY0DwFQD1+genFyJ6lEfGPoT1GgobHZaRqkohHQlomy34Vzlp3
JKG1o4Pe01fmAJ3ioewPVhDACJvHu3hpl4M3in5rO+bn8wCECHyJQSJ+E8LG7CT0
RTmvwsr84NpnSrMwojvTOlDVhrPbSESjxiRUQgti1dN0S+lpdUJ8k3YIBeTTy/kt
u9kHVHmx74OWrrp7k2rq2KE4C2HLtAQMVvph/UmTWEKwkumXxAMmpqfNTlmON8w9
g2sZw4TRZBd7dDpjJbhLuf/lYAEr2VtkFHQowHTkh+oOLg52Mdspg5e30jyVwW8M
JU7UjrAMsfSD+ZV0vH7h6yFP7X8gxIXavriDhYI67Em5oyIK/GSMU/0HwiM0oG0k
0bV7OBKwjcphD8c4UXmW3ihT6iIpe6viELjtY5AnB1LgH+bVv1qLjvghgWUXltvH
stMm/P03vIPDh1cnpOJ46dpq2lfAuQe+Bt+GeTQgF1aGMPc1hosAcfdcaRe4aCv0
7p3itdfIeDNFyEkkH8NZFAb3EYXhg/tdiL5U4+EM0zAoMC/EP+eJUuox5BZSOxYu
kTWz+xLt4kTz8d26J/ZLG0iU3cRmKYlVt2kFJ7m3iR4OTLOxBeVhOdh5i85XBI5G
GV9uAbkyL7QWMES/7Tyk1Zoy4wiDOEAW8ub63QkNGhAI4ElWPlPWxUdkntZewbBw
y7a20E1KFsztEvT3k4PR0pMJ7Nm5HPV9XvtvQxf/xy1MJh4Xqbv3OBAAret/Bvyi
+icgZgIywoMpd//oYtxX+zc6hFkMX/48Zb2Dt0+ItzsW+LNV/0//kTZKi2kJgbEC
m2Y6ePP7XYU844MVvHqF7mJIXSpaVWak5koeXYe2iTyIWEN9utTnwnXNgPBy4Zzd
CjxFkdr91jcrq/OydmY4+NdDQcEvBw+F6mjnaXJEguv8khe7cHgH2FZkqSNwRnn4
PbdiqgqYIKA60kGqps4f2ltayIHQ5a1z13LxMa1ygrEMgjrK5W7L+ASxAWJBU4Tj
4VFUallbCLkEOOBuHyQblgZHsJeSyaoMIXMdezH0dM+A7ZZPMwmLRLZH8E6AsI6D
7pp5SVbki6ga8JDIFJCrzkUOiG0MHl24Msj6I6n/HpY0L2Kgz9dHHbElqri+pRWN
EVjY2DbqYBBfwr5GCeO8wntWZRtb8+L7az5utCuu/CZSN8uRrOlrYZpYgh3EY2UX
PezmU97n4qfQkwiy4MAtALVEPxfi6wVthHjXJJQ94Jy0gSm185JEycPl26XTQWMB
xrRiA1SYzKLnfgacXHB7NQYU+Kfet5+8iSgHS9O7/a28mvljDpeQuNomiBpCIyLV
pHnHuROaOG5bdFA283IrxLpaSJSrRU7/jnC/mb0FkJcURYklrJs+myBoQjos0say
ooSiQzvT+B8iB5Ijz/7dgW5AFENkdbCJU0XC2rs+LA21nYysSSqWvQxXkIKZIEES
BlkLpg1EJtGv31mgSQXJBgqCbL5S7z12K/5v2G068MdFXbMHzwLXOC1OgrA0bD84
LL32albAYhO48+02CTsgivqg4zlXUl5itL//dQldD7v7srShgg8LQSEkfUxe2NnC
p5H5SjhxUmEt0NHLww6OYFGpkxHQV0VG5dhD5vkkJKchv2OhsJNpEIFJ9mEJNbA1
EK2XTIwql/xeoKQKqYiYxPweIoGYTYK+fGN+Ebhc3JqY7YIWTMq4DrqwOAN4Mbc+
RvP091TljugLABD41jBp8LHE4AUK/jye/TPLpdw/bDEFoOEIrjpYQH1GoQT59ops
mgFlQx3fTs8UW1uJaJHWDptN2KL5JjYYhb+j/pgx8TA+BvWZC8m9eURdHrthaEGU
ZYukBrAifcYn+koURb5mi9U3Mees6qRXV2KF0dJCIQIGBU/f5KvC6Gd40yN1Nr1I
7iv6xDSIJw93doytI9taGmcSlUyXCQE2m5aSa1qGbIfc1WpC1KrGCyv5l5dqTGTI
XwEBTBw2g1JWQCXp69sOJKXgLRhr4rTaLdRhPwjFsEKDZDioX3LzGPS+UmA3/IfS
j0ghgFcM4UV4Dyuqj9KLxDuOdKJlPFkS75CjjmivOCM+RMopQVaonpKEhWvvnnTW
W+Al4Bq666QaTCrszLcHx82tt4Yq87XvKgLwOMYHpb7DsGJA/lJzArHHbUhs8b6m
s9e7jAASz2sqWCQwRuZwBcJh0CgFZCVb3ESwp17XwH3Mj9scwWUztL+0wYpHFi4D
9ycll+UfM77pd/bYL1uKYy2nydHppoG58F3ZeUUz/1mf3vyluwgp1SP3U2+t2pT3
lnLyfq3a+fuhkyxK1M6B53dHfj/Q9AVU7qnDNCNEySHKCATTacD3BXW/8HuLbk9l
gdf1b4Jkrwe8/j9kfDcNA6RVlkvO/Xi25tk1t6+eKsey88GmlAm3o7H1Jo8ouAHP
RgJWIRE14lZa/QkwJ67fhhyxHr6uCdCiGWRya+8igDVotTqIKnvDOnhZrk9qAff1
N5jdjp9mUzap3sd+DzX2Hrw5d4ULppV1pG+uVN+abGR29TekeQpxVz0S9Yu+m+p6
UbQgVVwRoOwdyAExRw2IM2P3FXAEvDQGo3d5QixdIsXRp5nZOczW9Vx/cVbH7uQG
qy6VvbN7siwyOLDrelFOGFZBNMFz+uOQBwNR7As92ZRg+kVH9dOhg6CnuVuPLQ5k
0FnGw/iQ7WFjJvzLlqLCg72zP4atlZHkhDNF3TzHXjNWj0csd7Ga17E/2n8L9WZV
klnkAceUCAing+cdY/wYA47qwkZ8wTkpZSLTdJWdOejPlc2Ydhsh0kCKThdcag5x
aXm7m8tYapD5UNY4iqyoH9Pwj9IXsoY9DP9Q0Xm7hk80OPCS6TrMm5MwkxAVEb3l
HhZxzUhNzo5RGVfKnwBUpTtfJOpQuXHnF7+utsrav9MUOZEZCEUXFXMuAfKuoGdg
AOefeFz73YjM4d/uRgJOL8ORC5q8q8r/nPNTE6Z8eNhPYvpBMWMkozHCGWVEIX2L
9yscJ9vxyPw9Db7mn9HiXMKusvDYcaK6Zn2j3Kmz163OxU+5LhIzzdpgoDd1XuNG
wT+LCp7AYCCh+7PpcH8kuLj/ikj3t60IHFyW9xX5/HBZKMhph8f2PHWC0SHp31fw
zau17p9DaYZROFB3kSM4+FJkhCaukiCujGxjhZsfTT6cR43dUrKXIzVnnZgDiZne
m2QkZSHpCkSV0x4JeRnv0MOVBJIPtREdasj6hjO20TBguztvuI36XL6CBv6C6gX/
a9Sw8j6OpiJQXbSc23PHc8lu4kM9NutZr5aS9vB9d1+jb0vVj9Tokn8BAeekQBlZ
g4NLkpqAcJVy+CaIJzO0yBZFykwbgyDh/quiI9vC/+q3yaga6uvP1QM2upVCgvHf
ZJuNucVxgXonWKrqznXUoyYmSo924k25LzztENxulGDmAO/uqP7CV/2KFLUCRLYm
0z+JOPYO6w1SeTtSgwI1/tgTMBfZ50wHmfMI1mgHojiKADDt0htT64OLLJfbAn0z
89mfOJwMUox4cKVMfpLDy2qaXUYHlW5C0qodD93CDSmpzyaMdZYml0Z+B3uGZoGj
45FT+2hVPjSFwL1eKfbnM5e8FpZwoYegd7g4gqnUf/iQNTe3wLYYRubiYr+EWNGh
gP8TCeGz5YJS1VF0xkeosglKytAS9vQJpIYcZmnpGuOSM4KtNzXgvBPHuwG/nYMb
7uW/sxyLz+BykMw4YmGn5X6oF8ipZ0QWyXJjzlLiyHKzxrVe8JgzNKoN0Qow+m7m
QlJhjQZiKmbHSH+awLMSt6GdHITGA6JWek/UlUaRhDeuZYjAI7KyNv5x214rSdww
8o4+SlUghli90+/mUKzq0ALzDehpxr0z83gOsElkrLzCNgoGgVCPwcgEk1Thw4v+
EFFTqGiP4PEKtHSRdDvPSth3WIXBWrEZnUlv2rrz5aOSbIqtcpqxVTZm4eMbJMVF
Li9ewGrMJlZEHjGpP5Q0woFr8chfXkCMztSJ3Q5BiD6VMDWlJzDOfLtznT3Rh1y+
BGjXQtaRPfK5q2tszvWJPWsr+51rSMlsBv9Wx5CTiTZGP7i1f60i5Jj7PvokqGrg
zLjcL/lZEc0mUyR41spH3P0IQl7e0yq9OT2wSmgCi2rQf2+2elYppZ0Y85ykUWPn
/qxMul1O4f+iwtFCpRir1GCYp9CiciXmLALoM8ywy60YY2ooTZJDHqpdzTMdCq6e
E++02kIb2A6YnJySEULlRdclE1ndlnR5ihDwh6bmi+GuPOcgwWmyiN0QyZpgbuI9
m+edXf8sOjDhv+KZJ0icWah9ghaLE1mhMaLm57SPH9tZmy1nA55QyoJlP54PTCII
We6vUkhC7f0NkTRSoiS4k5y/QKlfp91xTGnYla96IS4cWeeAt9dnIsJEAdnffv+T
Pcl5ETM98rbHuNzxBeJ6ox+b2NX4mZRTiC/6rAUdz0YHnxk9mVRMeLRV6tmFIqfT
sziJ1f2hS6Bam9PP88/EepxPXqz3b9IT3kLVd+3j/ErTrBzP0iuiwDd70kiu7MTL
bEOBPIcqxchyuAd4boVZ4MSN2KyMImWxSvfdsyfNJq4gKDUIk33byKHNEo/0jhgH
UVPKomEQ7z/dWvbrgTRoHS5OoM2a0dF1mpPeqOzO3VmmzhGgv8qmuw7qDL8IdJp9
rWuSv82NC2eQEj9Y3d38xfRtCumSqRU8sF0oTMtne+Y61T+51Cpjhoszr07rLAIR
QxeV5rDO/U9feiwoH6M0bwpdyJIB89Kj4TW7Ps8BMXcfWJMyeWVseQDUGMwz4xdD
vHIPCp3Ul2K2E9f3VohvAsupS0PJWTrEd6iMpIO/DAyaHfmqLMMfwD901efqcryn
WZI4jdjVu2EiJjzDuVd7SmniC5+qWBlVvKe+bDheH+E8ERLF4YAqz8EX7AsPnFF1
yZY/0yz8yNle7PRGJioHP0wReA8fIJq7nfKomgrdpTUc2SIxKEItfwq9Sa5lcgeY
KDovd9X4esSrlNo4ToPQ8Hqbs7ZzV2CKfcdE1/bAbjjX8dWrrkYHtgpAwIkroF0v
urbfVRc1kDNCucpfdmxuVoA8QCBpocLfJF2/f9acNz6vGNkzZDqCJXyMXRkgOSnn
eplRkDV9ePerXiHlhoDnO2KP9ecAc/fW/dvM+x73/xaSYSQNQJghBsDPUBC/D+6S
MP9xrps0Zs+UWz2Yh/ychCoXmwdPsMNz8HNjBsSYfzEaEnulwYMyNAhldfX/qldl
0I7PCWjt/X/lgNbFlRw/x2P9DEdgm4U8BpBAxTqzAgSbSoiw6xD6XCkChfMB6jjy
K+rhwg9pMSGbKCPWu2UVlUdENjyk1qGQ3+kU8rPcuKCun+e6qdYqwkeBT92jadXm
PLlNgR3zFpWdEZ0xKCDmyFBfC72d84IhhEiJpgoApZl2naUf3W2NagYsFBS5f0YN
EYScCsPwzOBEGxp6vXed4YiU4FcWGjKfZFbqoCXmzkPo9IG4MUI9vUP4I2N3t7KL
noTFnwAWvK8ppKEDHxWyXjmF9qV7oOXB7w39aAQ5UH26o3MZFldWICU0CPsbsbOn
je5o/cbxBGGSuSJpVtyGIz+YV70giGvrs5jJg0PZXMj3mOirL1z9EzSJSG6tHAzk
5c3GE9RP7VbRhL8XhjaK9en6gYHt8nDHP0CtsCOW1xM5eOqpvZTXGUR55mCtvIoL
gM2DW1mT3rzj2IpubwuMOFhWA/1y1hl1H+UboczO71rztko+peuIsn7x3wlLKUyG
juh8CLKQ+YPXZqg3hRuvJ1DQShdLB0xUYJW5nEw5IFNlF8UIrBE/WUe6RlDNeiBr
9VnuMHEMfLTDMsd3DsDqECtqCIbQoZJv1Zef9dxleGC1bZkZ9DnlYrM+FmjKzbSx
0cSyqT2WsxuSD57xduHP+yDvw0/4BLVsDJNx+mpj+ntoIrjzvSKLLI1whucHoOwR
fPiLEygjb29dmeMXz+b8scYaqTtRo7GZ9dZLfB5u7L/P6eBIRTNjUrocF+vmRidu
wnbN1vJvy0lSBcBDwTqbqeVj4suDWL3eZY5eBlOAV1hZZBGxIwl55yDDAsrT/upK
d7xDclJSF3svp8GVuFf55LHL1sIa8HB4KXwq2i4thz16Y/5SLTP6n0OqsA6bG3BS
Gv2HPkbVP33EvcpLjXFgGBGaBpz0dyA1+Oaq3Vy/3YdYh2vWvLPsnSSNEq+zlz4b
ExWPbowY5UcTLe4irwCv9V+f35LyZhEddOnfEWdyAuWzl04NrglAcXNPEA+DyonC
p0NAD51fK11xGY76AL7zu4yxuaxfvFCs3OFwd8qnUC02xkr0PZVaM0WI6wAKxUkp
wE46M//nWB6/mWF7g1wRjKeNaK4/fhK/5zvckhL/EF+7wMAR5MN1FiBHoOxITPxP
h9VDIgGEyd2z1E+LhTQuPAVUP5BMIi9dMK2Gj3+KC5MIDU9EbEXiXeDfi7iNjM0a
mqn0KWZ/e7WV2/jtAw3TXKzX2B4NLhnsePicvr3YDIeW/2viHIFx39XtWVgn9HW7
aG3odarQ/fxGvvHkrj6I1ayAFSh81Hrzv41EuAe7bDVrV0G1hQ8r9ID+6w08YCPl
k2PwaG3PfGcY5P1vYAdBYT0NySwIQ7U7gn4qrhN3EaMDpnLuCfH87fjZWqj7tM7C
LfVxH8XvUvb7JJr07IzDLeXe/l9pBXc5tUjYpQ8bgHH7uQ/a+kYeraid4CPC4lDc
Z7jxkk7HaZ+8LLac9DXd+hCcOSvweU0gkWrrw2/8d6wHf46OK4PFpncqvUB0ttH+
0zrd5d/NnJ7gTE/yE8BH/gP+STr8Y8pgC56GpBPgMWo152XwH4s2llZEmt8qEIQF
OYhpyln2gUfZN00gf+LgH7ErJo3qt9EWFaizAfNpVLQnD+niKvpVH/CcO0wpsHRu
u6Hazs8u1kCMQpfHIHuvoB0B9Tu0nA2dUbHxc3jLcVJKVOraMzHgZXkNBsHoNSwO
NH7n9/twDYXrYPEhsFRl/77ao/mp6tU+t2gAOHEETI/hSLb4NBjdr8A2rQXSbKan
5DNCUvPdoBVa3MD8xREeJ0YuFMudD+5HoQnSsJPSX+mlZLnpXtT7SGXQx8caFotj
R1vTaqmJXDDx1BQzCQ3uNZzwDYGm/W5OUjfOnuZ2u6hG5dkb4wpfvtxmSjASfx6k
SCXCPhU2oE8mqwxiOvoDRhhCzkAFWVN7mrEPnoJDVM4jNhQ0Q6ZELXr77Y3xVaXS
g9A4wETgiJYqxkVjekRCK2cxFLabh+H6RAtsQuQo9mE7tslUVkJuop+/20zECJwv
86h39LyecETHEfijuC1D9ktBtoT7hid2bbSJAgYKKPHph2ti3rtkmDwnXMVCDY5y
dXxwnJ0kYZ0jIvaVxVtcwnC1UkX84sVEyS54uCyGSocTwDsSQ526lFvBjUqzbwkf
MoyUcX1k4LomCh/54rTXjLFrvnNtZVHkm4TJBr5ay71v6jVMDZxb0dQfVvWtXVwS
u8EuG1J4TAEmjI6lfhyUAhkBQwgiS3o90llUPvkfVxz3RelAxq1Lh4DoCCLPsY54
TcDpNJfYC5pWqgZC1GonNqal7A26bw+xR8PVZGotCYBdZYEPo6aiWu1xl+oP6tuN
yqfEtoVjV2BwEAi49GwpoKjTe46/ruMsRcU3IgBQR1pEngw3IgXKxv5c2vdzb9hs
xVt3FgRCy/M0gP9GNSZK4bLF3xj+hl+2zHLUPrBr1twMDy8+I0r1J9P6yxEF5KgA
Bnf+cNCav9QWLkqfXayEAM+PqYKO3UdIvRhem8IC55TjbbCfen/BJsjX2K19ptR2
ytix6ki2urXEMIjG6/bbWxDz3kWuK/xAOnySgAB1o90GN9FyWjQfAKjRsrfLvdTe
7gjxMyPp2kiBuBfBAt7CWrGE080nCM/KSTxEI3jNZ8iXVoCZmrZt5XSkgJMVDdWY
Yjb3hS922rOshzaeyok6U5uuDKP2elVoqBBQdRdsNaLgGfneh3kGUGnhAin0Gerz
9v1gz+hqHB/z2w/QGIy73C8m5rBf+JEVrSRBEYnKC/upG04r+MvTYt8WikQAVj3H
1yI7VdgcPdshZd0k7ty1K0OEKOZtmn0DMtZtZFV/cjtEhHURAOMLvpX8pAXZCNIu
DVDAo+r9wHX9m5ldf0LXoZ8cb2Sh29Ip3lnhja4Ax1zljuQtsuRtG0UWo2LUZSfc
KdOZMLwH74k2IRM+knBa9C/PYRrCveCQzqB/OKOBGZkaJWurgNQaNBGjEynXvaFT
V0lVEN89svHIqWBPkE6O7ExWfMN86ReNoyArxJfoUN4/eIkSeKw7Usf+/QHNeqp0
KaUV4x11Kdz5W81pAMSucCCNAvufNZZ4rlZeqcDeOM4AXKAuki7KKrqPDMMocnOv
DxyUSB/fqx98dT273ySfkUh3EH0XBevH+usBUDrVyGISZZ0inQmitl0xKxfr+o9+
RrTcI2WWKbEJW1+PHhVuflvg96DwnXBs/+jBcKQCVD9SJZvPouWf1MQzuPf0+wJA
OLCrBAVZ+CcbuAR2yH32uKj20T7UpbYDaP1e5ENAx6g4syieLrP49UGso4uEyDjU
YJHlmeg0p4kCoT5a/htXnS96HeFsP6s6yQn/YATUZxI4ZG/q0QFrHe02PmKMJkKM
K+3f8dxQCBNiNPA0ADuAkA/7m79TBLN3JKUnjbe2RaJsHN0lVKqyv0FB1yfRk/lP
neiYD5D3A7QlRobP+JY3rJzE1t4t7RA2jbnA0T8+prONoXqUdj1lbYUTrap7N5Mf
k5qfN2ELeFfs0PUeEnVCCk9fGyQtGui6g9+P15rVhg/bcQIGr3cqbUt2pFafxEnB
xF3ACAadKfCOKl6HGwPWQhe9+NpdEj1WezZOPvv8EUSraiUnjoPpfNR9+zlklcan
Gyh+jBl3h/7AZSKjOHXQeaRdajAxmhBQcfhjn+gbruiLruu9/cFzyD6+WDH1zBRF
5qdnNZWjSK26IrGwu4YiQRR1xqZZStjBEln3bDfdHxEV6DmKP3sPBTLCa8zxJyIP
N0PLjJZEEJOrOjj20Rn5z3riVlvIGPgeeAqwArge4YCJQJ39aq4Ua/TY/l6O7tQ/
vjoQ4TJFIrv9lXwNnpWOEv1fW0DZqRRNIPQ4ByLpY9N9hrVUcuQxjbT71eevsmFa
bTHFXh21Cf2ulZuZZQBaDZ9otzjfVdLN3+UaY4onbEjpdbDRdyhuJiTFzJVdSO20
dzVHHFuK7YvH2oCE908jc1E3MLG9nM067vp1bhMjMXmLO7O184EFWe2IBA8Uhdam
CcwXbPNl7bf6Q92AdE4jC/Zy1ab+wpmC7etzW2kc6uBvs4UNMNhTnh2OTNHmeZTp
O2qFw0lF6FceJ7pRNG3iPu4snNfaO0AGi/bpUuONCJteDT5uCf1C9vHxjlZfqh/x
ZH7Ni0yE4kjP16rGroqMdgNP8yMAfD414hVnUB8SsL952YnE7K6dz8SadA2/uNnM
tfR4xfC6x2YfRInLFIYoiTSBgtKINFli+bk8OILetBKYmYTErYwL4VyfiZqGU8oe
z4a7tlbDszvPuVRwUz0Hb9Fm+h23XvOl82ahpnOBI1So3Jv83Wqrlgt8ZpsVPrNn
xGr2eSaEeAPFjNnNQuaZZWuypb+/4nzPpkI4IAZ9VAPJuTgyxMYzQv1yR8VuiBdn
HcYJ1Lq5KRl40YpD/NtU9rZK+43GG3a47Y8uwukjxcIT8+6kCyX2XmIURHGXyzBy
lPvcTRUKwWW/cJcshkCegfgjMDYxmXwYLBhbIjQKMMXrU9f6btazZlIHsBdk4Z4S
o+aiXJEAmzk4NH05c0mU9lGXzD7cWe4nB6W+vh/X6a49mXjqzj9qYrS9dKYhbsNP
C9ougnAFPJ00FVw+gMRinwRnyaeOnut7CX4GNgK6DLQDxepiGY7W5LN0yo3FKnzS
uQBPyMyKCsq+tQUhI8/4+p1L8VJKBfRRp17oAIK6eROis5/nT9awG7+AHILdLovm
NqnT+nal46sgXqM/vk9yB2lqB+23gAJ3XF0wY6YuDRc7WRuwAi/QFYw45X0tV+o8
D4cBUW9592/CtLWkKHND4ogYEjDX5p5Zp6ahw+5MWwswOiakv3mbJykRZq/yBF0Y
H9tmdr2iwWQqvD7ZZP1uFGBJDbwLxlODkhFRYenzv8E0CkgkgO3XMm5gdeqHF31n
7YJta7SWbETJnNzUokuvN9nEmgT0HH0vvkzut2SRfuC1oZXmE4m8/BlMTT/9gK6Y
IGXswnZZNXdHiL4ys54+nNFlUQboEuAS0/Y0/0z2Zc78KL4sJfvlouKPXgnkyYeH
G9WxOA0bIBqewvwXiVMz2y+CjaD+HivHQJIaVaNBOa3HodQVjUAdWNLq6qNqkOi3
LSTAyjrKCou1URwe0+auXk8dx2bG23JbfdqXa3TyyrSBCyA5OgWGveU7sgCykf+Q
NZW9Ef4s2eIaHqRrUb4dpBDrP0dNxvCzdRYERkF9y70ee+D840QhFv+C0fdWe1eK
LPKZ0s3AMXzX/1Cc30e66cEn+i3QrwJAtQnBpcgs8SNKBcV47skDhEm4i80LLLXo
QXni2yA6ltkDzd4tXkYLBrboJTCzyF8iOVSnJCw3HPGr0vASQ8JRgM8QA4z1nG9j
ccKjErwPT57tfUnRmSoENNG6+arv4Tj3n+AxJt/sSl2sah6xTiWTPTmevd/hxmG2
HhuqSwAEc9Nd4Slw1T76HSwCEUj+EAI9qlipekORsL9f1pxGUMZLT3K8oMzeP819
68oGIXmAP6rSsepE/0B61F8pbhZu14y31PokjyNCce4fL/TFV1gYnJy66KKQcQuD
qWnBhLKSM4Hs66foz+M35w/1FkS1JXOQ0r9ZrRKC9+0qBQABei+4Q2iGCHRsVhwl
mHnEWHEkzB3Uq937wO4bT91+U2d4OSQIhwuPidXNC4X77kn+vacH75DoQ6ZK1PE1
0fiNSIh/giBlHF7Q0lu6t9Vm7kRXn4AX5g2R8Qu/MlKp6eL26rzDaXu9o2xwYJYW
auKRGQBZYcBZQG998fxA9+NgBl6T2Flm5OzHThgxOHWSM69fEUYZ40bfwXs/7tJJ
TkswAYIHYHKI0HFRR+YAzBRQaQ7QA9Skq9HcWrIqweiB2mkwuZI8UX3n174wWdxG
S9yr17L+exlB0N12S7i4Bl6ApR5E2nL1H+pKMjMKuwFe1qoqtht+CXWI/mOgfpfs
3LLFrIZfj46sn86hFSFjhLnox+d3m0wSsQvX9umUOLHXHR0SB8e16ae1SzhSNGCQ
BIrTF1AS1Voc1ieW/ywdl0Kc79KX6MTc44EFAuyDfkrB+VgJRlwbdDb9upZ2lJdr
+rHEqFTRsjB8DPZWfqqQKq6XYA7yzYcz0tW0ceoUHRJOGkTAX650b8UJUviOn0dX
GBmBF+iM3tGI2KCSI1Fom94W5tQ7uJoEHzixnRqDmiXM73V8ceuZee83SZhkH/9X
5t6p7f+trsdLDxsU4+fOXCiPPrsx5OLYhNJJUOAu9GkCm7ISQCU37kavrObU+VKv
2K5ppazpo4SIvCVi1ODenLVR0IIbqR7MmzTjbheBBRILwv2JzgQvpF8SJbAiJzsr
nzjuDgFxgi5HZUo8vhertFioFyntQ9nbUB2OhRbVzTVUdWkXNLHgsqtzrAanWj/p
wWImTEcQMHCiRLIYlSUWTOV2jHEe4FEXptZImeeqobbicj+KdHk94265YqzxEcQL
TC7+KF04dh9Pya5AyH3+x5ksa0XB5IzjW2xjekmz8yDneIQx3OGM0pDGc/lLXr+c
EMVX2S1pT0cJnYJvMiDp2OZDb7yHhcIjwqen8bH47mM28Z0Z4Vqa+idiV7s9Ri+p
rzgYn/+bV7F+zkvpr6uFhnpPSLD79dRjk2UkBjnWhX1u+ieoKOayhp4KPnOHZKkO
Sr9j74ImQlHrUiyAXOCeQztck5/bulll7B8duqWrYRNzQrcetJPYIqzen1saFGfV
ocT/apKq5iTEtisF/04qk7L1rrUL3JrBxpTLntnToakQ4LcKA31s2XkcoO33bSzP
3eRE5RK70Acm9L2Bx6HJrbxBxXxzDUZtMWWXcReGfIhfpkrspml4pxflmo5QdwAP
FeNlrFGYjVO5eFiZH6s3nFFE5JGV4184bWBiOTODAzCaIFvZ1MWKB7f0AVQb+5Wr
KB+dCT/HzbiJiZr8gJgzu65siaY1+Gw47ulm7k4gjD1s4oRDPyYuMbqM6sQ1hWX5
YooZr9eHtLdU/0MGggylEhbfxycaNRzn0oSb0vX9aTuIo8vDKJwq9PEJnphF2TT5
+dyo6p1NViHzL3QQSM4k/mGimxZqtB0tSY1nOOOjl7nDlqAdKelKMZ+7vBztlOBy
qlW2Otrdu6GnIeuFFtuNwDRloguuF+8sAG3O0ysEPiS88lVabDvzVpMS0S5WzNKq
aZow/hQ6cNddqeAdGCys0YFyEhi0ieNt2CcUjT7kZBtHmKQxrioqxuFfE3ip2Uu5
SvzCF0WBJsc1axW5KM+Zw5v7ERrrbRDPwbeKJhGSAO043/QRURhMGUdvJlNlLiOK
ShQuxKOOoUfS2QsB3fdInLMdDWkDLSDJaWv/tNXAlkrsoS8kN/0dFBVBPSNjcjN5
HFvvEjC3EUkU5CqpUFSUtukX6ptJSmOWVDLKFE/6N8GefxjudPV3WpLWNX2JEYv5
w1K0qc/HW4Mt5A84KCmg9Fo30X+PIAHgOECR5Rzdo0UGgjQ1wCfHeMr6wob5sJIp
Tq2SypeykuroHceHIx2E1sge8xd2cb+K/g5CeTvtgacAM9AFEyHywdBqCZB8VKry
p7snrlW8PshMAknHGJSC93LwBOrghPK+qoLAi2GNfTDyIpmPGSRcCszlOgex50id
V4xLxLKr+L6c4LbH8CLXHuembcdmi7MqMZ1jVSIVwhPV2hbStVHrtMSTMNjFyXGV
EN9seB4fUyiM40MZW2hiSU6f7a/WQ8uhRZOF6emKfQR9vUQ6gm/1BHRBhc9TVaJY
RIl643IVmA0MMSZ9RN4O6UpnVbINMwt9PMLNbSfNcMif78qJEDSm502mGfV4IYYr
oYkDfFl3UO9HlSS4HES9IXrojfC8HwzLPoVjwqOFn3uevms3TjMUv5N6s4IkWeQ2
GuIvB9yPszD3bgnRCRb5gr7lKvYmCwuxBj4hBX/3swLH0ASQ6EsNmUiaTCPA7Pop
DG0suwXbghfaPeJGzfCMhMOgQjp/D1YUmmORdxQ4mVzxuODI7vMgidyTjmkBGgZV
eBcxhat7ndjMyRpxlZ3A1kvzmeLTVzblLeLYJmwDOwKd8fP6q57jCellXhJiRctn
iN0fF8XkOz0knmJp7s9vqMGOP89QMdj5JW6THY1BozJ+B49KTPp+poLXIQsR/dza
wW4G5mfnh/JM3N+DdckexNCC6moHPN1D8gwH9F9Gm0n7WFxSiF2di1Hou/4Nn37M
I63ny0PDzw4XUhXva6PIMQM4hds80qXU7Zp2zKMLvjEs/Td8Dfj19C9HC0NTLw3X
d/IHEeWDRoDnVqILX0W0+y62U881fZ1uHXrx0WbgqQO0qf2hs0rzPV+VAmGcuG1D
y4ncgltOMDzDQUBj2P7gBXe3I0p82nSyiX1H+0AHbVjlWgS2C95deBNNeqe/aVAO
IhErstr6n0i1W+5fWHYcuyIoiUeJhqFDN03/m86TOk8O9xY+9fGtYGzIOkpdmebj
1IRIkewr1B/Nrsp6gu3R6ElHilsGM93/FozkuQH9Xr/764l6U+IzUJJBWGDITWgF
hjA0CrBxzS6BoE0tq8nZNPvNv2qRlf7mU5UTbpHCQs8QUXimeT0ivZb9CO54LjBs
PMzNo2Lk+U7IZpiVfT7JAIJbxa7JijPQjgO5dw05QEFlfdLXIPmd56wOWSoGyieU
g2lm13USiJLTOgxNQRwDyHOIipgPbJ58Cb3IIuWe3F5I5bH39gFMy0Ils28YTHkD
ISdFUseLKh6MDUwEjqGZ0ywupAn62ZsuTL/o9WgjPZPGHQ6wRf6/ZfJtMqkUYbhb
vl8U3/DmLrAM95hWHVP+REq9fXpWDmSgDtiW6LJ0HpLUDFhye4evA7N8rtc+G1hy
lE8Oa6Fcq/stCTr5eA8NGaRuCMxVkDILjy3UD6LvcI18wIvFmuoWz/LgPyug8phd
PXSGrprNtFaFpcM486pdoaUpLfeEGD6CaMxEbGxIpNgnn6H8obQ4fVFMrP8m+UR+
E/CbUXu+BG1cZDQI8owHRC8G3rB+fCEqS9cvKCn03W3Qi/csa4zkXOalFX2qy12o
LzuulAuaCXs5Q/+btkfRoxGCuTSla5bG25sLyfI5rwmOcBIaoi7I6rCR510B5ILD
Brdr2SiN2DagTGkviV2OAwpMWgWGnstlCWRCmOv4IStLn29q7jrVmn1fuXrZu2Dz
SREesUXMEfR1X1JlU59HMnO86BG3JdQhCZuAyCHUSadStiDMe0QCBECT/Dz3TZtr
ZA0BrPK9kLq1sQNeS1ix11kgDyhaiYl5uJ7d7DLSbDCjf169VosioCTxdAsW15ml
q1PIAtq0OzX/ulZiaSaWrWfD6gRQyPDhKzfF9Qk8K7vBZDDBdhgroAE5IkGGSh5S
wG5XRBZTBFqRXJLhsKcZ/Nfm9CG6EYi7zMgjgxka/pbmO3W2NYoYQUesmysWmFBI
wctuPmgVv4cUzLplVZHlWu2MIMmse+Wx77aFZIwzQSCa1HFPlXYDLBxEonSDWqMo
ZAzVr4TWCPqvFxNO27WFQzAyTHw70A1RjLVj87K54cwgEPVH8ggl3mlGMHINZQ3C
JYBTwfuD9qrNC54acQkxVfxMQKve59adHhVUCET2l2+23hKcLxW/5LQ/fhZ4Jof7
UxNKgPP1lNZSNXNmXGF+b7Dt+wyyouSzgrZnqaZr8n1asyG+01hoQPZAIai5h5EP
aZWuECpoxCIyesuPzd66GO3rOaSb6S2j0nANkan2wkgG8cQklw4+6tQrh2VTgTsM
2ZOCupNPMwuEaYZV6G32cChFE40yzjUL19ye818TSAVNl283cpHhaBKhv10+IGE4
XnAY4A34xCHfdCeJh6mkdvHC2ecJS9JlrmP7Lj1Sy52cpnBHn0u2eh9eNHOnzpY6
ILvNqm8SxJEp105YQrGqT75+8mZqgAuwh8GI4UVZWu+BYGPQOvPwD1y9wBhUed+2
9l0Bc6DXXPZ+YY2P+Qhab3bUxbfGQXCvcUmacEO0HbaQolJK346ZN12v+3/QjxjA
Fu6vK89jByvZ01FvZcai43dJBgvbU3ZOVxPVR46+wxw30xOIVXNPeyPOV/vIr91A
MN2HyCTfsdXQt8rdLsCxMGChrrBHp5BDYLvSI6qUlij8mEDrZpuTxylSStUEkHhs
swARvU89OK6IWO+ffEw2m4yZVFdAuEss92XYT8H3LNG9oEsZSOf0iLej1CRj0Zfi
RHuvF2W8XOdh6tBS8oHav8K2L5uPcF1P680p4xWUsJxBKa4vTGJEGIC/UorBlEky
Q/Yg96duyzojQ/d7x5iMFwj7vchuE3LxSYza2KBwAqGIidPRjWJHdbpIllsuV2gc
v1BiqOjRdWqEtb2sndvVpQUUDelURNtxHn0uRS/szuJb4ZU+Yiu1n7nV6PwjSD4m
kyaDC0pQHZ4wh+aKb55DeBQ5eki+vFXpzGLcr8gNyhgz3noU2iMzCzxVkAwIPztt
JE5pvAIkNFhKACBRFgqXUxf1VLNHNP6V1V5XCwn3xMZIsRM75ShCz9KAH9/nGJTU
d8FYl3QxmLt+Uk+MAIjBe9VakphwI18NozDm64HCAB8sVq9GQIQ57luDpojVBE8c
f35OnuwiDoVZGiU7TxeHlUOtn+MUVyrCWrKKSCZzdjB+/OAjfFY/xhljjt4AGiuV
uQQhh5u7DTqW9CNCxEpqwZRGhGkXGMcK1wYl1aU8mZKwi2A9UkKphA00BkjnUFhH
N+SutSCT1sak8zgh2p5GzUiXkeSPIYxtD9kBjNnXdSwz2iu3SYQtnd2pl/MVOYP0
+vOLGSyQR9jK7H2YD5wGbi/ebPY2/pp36kgvjAQbxJVrSM4ff3yPAxunvYrY5LpN
pMIXKvMH+aOi+mKDGRJWStcdJ7GwmvsuKr7Irs4DN9ZW269/bvvpMIXMRMAO4cvZ
TO4x5c/Go5LD+zblKdRN4HIqztJpqa+AXuRAFOWyaZ4OWozEPurvGk6mTaBqU462
pGcHqybKRdHFEeLNG9ygg+0flF72VYaVFN5+VYxApbIvsbgnca8fvy1LDGxV6IUh
AZQDksK8weSItP6I+I9vIhXbEguwwSyYtxD+ToSJVUVQg3QYL1DUY18yndcatcEo
alViywJVzhMVBmaXI+syQ4sxlqBcJrl0WIy6ZZGh6+DHSekIMvT5VPDvrX01Xw71
2pVTQrpn2AqKVL2VkX91mLn6jC48p04irbSTtZPIRai8UzvWd4sPwmym9e3ZpR1C
uo8qLQYcfH3ECcpcctPQQ81s6t8WhWzs+wIe7DoM1PPjbtdSrXawoJMxO39/zavS
OWtFShyZQisO65QbRi4h5nB2Rb+TpvXH+KK5OZJiSPUfcwu1BxY+a95Ryw7kDXjh
0utPMyzLQSyJL82t/0os9hKu7tTl/FvPUe9VydW19gxM5UjO7Bw/Ibrl+6p4YL44
i+wcQbIwyq577oGOE9Tp/1jaXsA6Q4Vwon1MjCQLPmDhudSQYOPuqxduFV9Zn5Lo
wEnVCpYFFLgYyf8tQAI07naGAPMEvZY0bd/Xxj2DqeRobzRuucabrs1UpzHroyJx
eSmkWRAmvZwp1t8M8UvuCVc6iV4cyDDwFmXsxvRf2+cYNTn5tzhmV9wT08V/OUIf
F7HKJJDqmTSIfFlJ8FfwPdUHxKh4bFje6njV8VeDZBuqnI0Qt4THAixBf1q9aeN9
xdebhunmaS+ACR8c4HwejxWs7BDfx2dK+Z+jyRONZBK3s49A0oRL1l6+HzyGGcsm
a3Z2CcE0zWI1tdfd3BaN7kmjrDAGj8KuWsDoqiQfTA6RgMEBpY2R3MgM+Zq929HQ
NPB47zcRjwt6BRAVJQV38PewALQ+H/NYO9JTM5HGh/Tl5u3p25HEMWPktuxajPII
Wje0x1UC1086BQvM8qyg4+lWyRoB7icAVNqo0vL/q3NoerXKwzmn6ZWg04kmce1k
nJ23Oj4FfvoehJ1kU/EGrD9gdjgVenV+akEh3Y3FGjVQnAsc6dPW+8fVn2QMU/nm
LbDvWU05eEuDhv+9jVeQSjVtBKHR70irnAsOazZ1F0VdBmCJXKSPmNB22wgcIEd+
6jrEFzSUtZgeNUp9KmIIoLfF/57x36RiVMCNe//YgBdE7F5zRdHiYdntZifMAgbM
3pTWofh5EcLib2GSErGvgs7u1ERdtnqKV/aiyDsd9EXRMBpJHAL+RP05+Ozz6AlP
umTGwLVMnv/9cjOCPvBcp7SJpFkt6DoAXNXCRmjri1rn+o6DaYOiig49mb29a8wa
zRVL7Z8+hrKfOjdKs7OjAyHm42EWlLHg9hmJsE2a/4u4Wn+tycR/sLrzK9Teg9vy
D/6toFk/4QXwdqHhilNqiPOkxI+MB9I7wZbWpRAmrm59wAHAujcdFx2uhhrtl6pT
JtpaMx9+gxolRsg+bU+jFKXmCAl9Adn+UEB+ulFp1Yz3e7YkY8MmUjazH8hVRWQJ
ovPT9k8X2K45Xa1r1XJI+bjSba5LwJphTMNmVbMBkxjzGe2ItRd6D5XwwDZe2II0
n0H0wn98GOWeJS2/MSTtTdnU6ysQNePifc53pgOKzaaT21qZloSI8KVTbrcpEEq9
ETIZmWQO9mNHyTzkkFeY5q//KNkMH4pDm//oh3b2quDh24X124rhvYpSVdO9KKVV
J8BKKco3wMIUg8RrsVXvTkGKE4zeBE2yA40dJ2/S3ecILmQupWOWmIWBmatLPY24
MzzSn6URPX8IXPbCRYljId4IlAgsd43KZM8k7WGkNNBgZ0dtErY6LaGepS8TUIRf
WAkGiNFcxCukytfcwWjQe6gBrpH760QXt3d7oDwRky8m4FC3vUVcTqQVpdWWYYn/
enwRsXDl3xQSD9jV/VzIszvnlqLA1SsxdA1Fk81UM5ym/lX99zEnH8RXSvviGgbL
BDhjIqbcxocKUjLiSvJBlys+G1NxtVdNB7CIFLnKA8A1NUwvoKjAxqy99Pp9wW+W
5ElvXpxiXD8VLghRtVowSsxi90sIhYKAXbQ1B8wbExT/MpvhrSYUCWapzh/yZ6Y8
PXKI/AdQj7CuZlj/1qTe5pv2bBM7DDBN3nQWaDwFeeaefGF/hpv7dRvSn1iiTS8T
oXKvwluh95o2xHqJcPInOm9WOAyr0l+/t0UF4kMY69rCU2+amksNPNyySxiN1JCT
iB/VIweOFp8I05NnSi1NMr/Ht3P+CJQeTHietNPK0IbNzr0ntTFborHgC2ei9M7g
AaXRlSKCGyB5Tcbdd7gaJas9Pc7cIktmu6/KWX/kO+XZ1+1ddllsrEDnyoTiHZ+p
pqYOTrEWZZlpzczpyJTeV/ktWWDD8k4MiT7fhCn6cvtgE/DwMNdtNANjGd4go7MS
yRDLjKomJqbzC6eGPFCqWFZAF7DqZkC7AP2bNAukFxnnzxcvZfzaKH5kNWY7HB3B
p0+3Y6+C2hmFCpls6NN4A9znSqrskMNeHjcGCweIGUPnNQJRzZ+EfomdN5zHI8AC
L15xteuoDTL4mj3FuOKy2R8S1VgwkspHWaPYSudxzXDSO7/b0nzRGOdr0FuGUaWr
HdwYMhCRmbTe1G30litftULVFjm7BAOqCevdlMSPWWLvkjViMzMCl1OTf0Mx4wOU
QOw1UEDtyd4jp//OI0aYDvh2NBEwiITqSze86XBAy7ERe+DrvIvtVxDQpWrxhuUG
PllT/xLOL5qFj19MGnyjaph4EL9qmLny9VCiWcBVaRaKetckfttY3B20DGoxAcI9
atg7RuDoppMnrIy2TauiunatiiyB4fT/SrmTw4pOE5Gvntn66ojAz9pn6VnUziMk
AtIw7pVFsUAlnirU0NS0jyTFtuFD2go69pJ5eBOiK+kpxd8i+4wcQspqhjicHSo3
WwfS5K4o5dL7CfONQGe4OrYVmdjlpqGyX6efkSYIbaru/NLImJAqpLQPzAk+ENWL
pL8V8eTnjMdQ0OIYesr+4gabqKhxoxuYzE9VQabEZCsWfSj6whF/+Ov67p0pZdNX
yrdFDLiu0Jn/0CnBe85s0SreDolxgdlr4j6kHSxjj4lq7md9s4Wz/5ENtwNyMFqe
UhX9Rc6qAkxhyKi1egK/46ZQf6p2Z7QMYg6rrBUtf9iG7UEFmjqLxsKShb6WG5Uv
Wsf16Hj1YjjJtOqa54WVMxZOSz2/ZlFsxkTWNNPjSPhCI6qZhw9L+5ojRCn0I8gA
CmfXIepcb7xY7BWvTUcwH8vKfPp8zPXTw/0EoPAsNTyO/8OFjmnOnKS1MYU1AXj+
02LN/qR+81QjL2hGhxWppdRyoiq/UakOTKyjfcby8G8MS3iPFJUScnCWeOWJG3gk
xirtuMHsEl7idDTcCl4gsCE1L1o5ehgttVKjrQTnTAM9jxPXrhVXRm34w4pUqaU2
tOi6aQk9Aj578cOk+O98jolAgqyYn6YF80QeLPIDpne5NMqgAZW/FRXhcg2fWtw6
Ygr1gyzQ5jhoqzAeKOKJ4JA/WbuWN1PD3roeUERWXKFCuhOuVPgYdrBLEdGhBxr1
KgWYIjAvTCm/lCVH3tJOldohWI4VVt9IKlUvqO6YePdSYxuHF9CS2Ln602JGk74z
kmiARxsnlrNnnD3lbgyEAwIGzpEHhorsZxoE/s0zsbaHJtQ5lWOLxmJmVnkApAGz
+hpdlqGYOJqG2m9q4g66g3rLh/pb81fY3dAN3ox+AWEEP5BO8t/zeW3FoGaalRMO
LxWGZT5tR44qC66h3jS+Qqv/tJhPwKYXG2EleyUjYfNnEE7Hh/mFP+MhIVUk+1Dv
15plwr2rhiqBbREjXuxuIGp1L8Za/dNSmEUVbNN73oypJnfo2jBFQZuQZ/ViZvkU
f92Znt2mpJRouC3QdFoo6b3Zj0kcTZKs8bh1WkZRV6+yxyJQFCV0GjtEGiCQp+vS
gXVtciKLEuwARaegZMiPJHKpuAngL1W6Tpy3xlLqOPgbkM1A2Lk34RviOF9telyN
3FoHRgsdGHXmj5J+IsA32Mvv2kIdFV5poovyneCBYjiGfjpr3Cn2kWxMT7xAdTKu
jwilhhOmO2/HQtc6dtGnC3JjjDdGLG2twAwmOziOJR0ngghs0o+UOHbAoCLBYhQU
dlp3+MLOkWawM+hXNcE+Ec8a2vJ+/U+jaFvZwdAf4ezpYvyh+FLmqEKM+oIwYPB+
FgHaa/pjP+kzs59P5xIJfbc3PH00HVCOxF9WvIUdz33klLJOSOmefKmZMyMyFKn+
q4SomWXJzMxISRIBZewXinOQhQxx11r0E7/CW6hG+OHLlYsux/DniAFPZa4Hx2vG
OZLlC7ZLxuCxAOqJLDxv5IR6rbLvykCB4T3GWtt37QeNEQo+XxNKRsHdCzNS/E+O
RmHaaReZ14MALQ5WkKrS7Q/HD6X64YjmUoIYZGHyC3GzJb0npraBkw95NNtIKYI/
hDe5VM4iR6hDBhyVofsV+7/YJMqAf+1elttZMuH0JPA+ik3LIxfVI77GSCArXcB0
o0BxX/vpOQPUISsQZiwmZP5bmrUAYBCLiUFSiZkVucneucE+YPhuTBMmubLSGqTj
PJpQP1A4LQJvYgqA/ync/7a5jPMJgKR+By4BMD1Ps0z9HwHmAIxEsYA9ItCNtj0h
WCmWaUkAzwN0HOOOJtEnLD7PInkdzvN3bFZhNnprIOQUt6k/SAO01BobdkI7+NRj
3nX/T2uEjq/4sj6LcNAGiEhn/2yUBiX44ktB2sdFqDZRVSe8FJKJWVK/ZVqhsS7K
7K2PNKARJDByTGxTPt22UdIC96RArhuFL99TgzP8p5E/fDq1AuhOredSWxVYkqhI
MlKa9bDoRJtnzN4VT37kX70W7eCNNrKGxk8dvHTAc4UoaQf7WM4qjyC1+oxBNW0F
NpnSkTrdxyem7N6LAij9va7I8nGKzcZ8+bkGo7T1Tl8lX0c9NXcZFfTAGpUOLh0g
ySZWDZwjs7nDSFwdwXlfE4yuTQt3SyRVGC0YWF1zHQcqF1WGsuAPl0aS2mT6hn81
gkdaGzH0q8ZzqlmpNZgojWTg4AiayyBEnr4WkBCHeNVN7zo1EKkgtuKn+rXHaXz9
2GSrpyCdhvZJ+awEJY/QeKK+LPgMCIGpD95xZ+SS1BAE3Hkt7iH2jYaYsIsl4EEV
w+BJFGTV2Slm+FRBFUBA+kf/5xrV51RUaTnU4guTLee7Duwp8/1Da5w8vLzve1F/
0dHrahOv6oV4uf6q+CxlyGW2CqXsdGtkOqxFr5J4agl/Tb+ZlwcztYdA7aAAhYye
Oxo1ECLXA9lzmrTQVNILJHhT9quDtSab2Eb7ybYomGAXDLWRXOAXxrF8h/vX4TBt
beP2rV3I576zYLLUzCZQEr7xc+qNaEU2v1lxSEtbZE9sTupz3oGffYYDTxzN+tmK
RTHIhCumqIoihbL+BDuvMxqqjAzbo5FUySBgbbYuBW2s+uBRV5FLa8cnSIzuh4+a
T47G3rhI/Y1qlkrwh2FWSmnZD42JrNLXnP6OHCINdaMv5vqzqKVks0gAy1Be7rAx
3xvQc1mwfpvoJwlKpnwCyEOCgPVYF6cCSOm90c+HgogAUbRXF/y3cEDiPTkx632I
TmVXq4cdFs/dbjOSx1Y70Bd/iGGcaqLxprajzq3aeccAB238HfdCbvjCoQmRPc6n
ZuEzRYZZzGOwppwQyaJluNgUXhKacjzbX/mnfBpHSAYDRrkjPet2EPKnRuK4uSD/
Kn8MFqVjD6N6scU4RsQUqCX1wHTDcoQH78dKJz+dlJUZKM7RnR6C6752avwujubr
DLPyJccCijoQfj+OBXFVBEwi9P4IT/8YO343ifSVr7chTl66BVBjeEgWP+Rpk9V2
rlYYs9jOXfHk86ZIgmt0DW/Jh2m+tykFq79QqIdCu0tVlLHp93N65P6K4LJA/Xhi
Jw53BGJ3KEvg5OcT84treUfmaOizVUwf894wX/q7+FSRf6lGNGAbIESfrWun4ZqI
ofgR8pVGuF4A1s5rvVHKMEAH7ZoX+0jfCbE2ZwlcCjXQAyCbDp3ioqpRsxm37lmA
pj66iCNl/z6bH1Wi+u4s9TClbMmcbbZjm+T32OtsZ8KcKAenCOtDXMqS8yuVzV9t
DM277P6adM4OaQc4fqVgGv2gMKt2W1dVDzxI+5QFYa+JLXL5IX7XCWqsmyCQOj3g
iExrzZ8+Ov+3IW7l3/sW/i/9lgXJZ6sXphGhBizEHhyrXXKlAtn86wu7QH6UulQ0
8kQJePybKaQIspE8Daalrn4V1XDgah3eqOp1nL+bpXY8w3q+RPRxOeQpyHGigjwx
zKOWZaRxyrhiG9yTOe3wGyZMDzKiXx27WusBBGjhB27fL6ENAAzCd1AY1TJz73cK
WqHhynwiTGdw//UJ//lqZrpt8z+eXoMimSgs5GpZjzX3x614HHnvB0XbtOMkQTn9
6tJG20UKSiJGeXqdfKNlqdh5xPyLeIT1URxuMhyNt6EZg938r3r02yINHhjIKRXE
atvtGwQyBAIGs5YTEHGDACdhv9oBGYmPgbInhnf/Q6mVD7TrzOLyBPCzEAobahU3
bESNCymX9jd60D4DQZfaOxQLUQiJ0CScjTutxUNgywffBkzE1ll6pYu7iL6IDmno
J80WdSPNj+SZCgUR/JKJymDW+Gdq3b4py95kfSln9HL5g7Y0+LbFrchhqDJrbEM/
aHFYyUoEjjO7D0usK4Wp7flGb/F2yY8tJtx9Di4ebduCgm8pxtK+1cC+o5PWuybq
4Q0YoI2CX3E+UdGDwRdiQ6YWPifLNgljijUvppBtwZh11KRg3hKUajNGW4hHHqDH
bWMkxNBupWvRlw3CxsdzJRsM7nXgT9CBNWb+y7JeArkxY4/6oipv4glG8u3cbMUp
JlNgX6Ac4ahJxuRJYeznjeKTeCoXY6a16bFjemg+DbWIm1O0v4M7mRS/3qsxxA8n
H2ZW/vuyb5GoE2q7b+KIAKm7/tjnMPQXsTk5g5CqhB8Mh2b1eHFJycXZ4ytX4a3j
I6N8ond59acQCT4IzoCWzoL0zSfXi5tN1MnF3GdYYw/s7T1B5kfHh6Zm5hYvcj6z
svruQk0LhhzBzbWH3bW70SajukYOC/7YxOHqHJsGdjQJEyyVoxVr7ueY9dPMNaQN
e3Q66yYBnKh0NzQslD3RO8gDoO59nVXBR8n8AvcNZZejroLHw5tDs8mptyY9qrwl
floWGUekoV0BHxUfpF6Ja8LLHHDAAQuT+fh+7VXfWHRcDoy+p8D4Tn6VLPAlwNsu
jDAu3OlcUQ2Bl1WYAGmo1yT0T5s2GCDhGSNpks0H2ZHL7VUj6fGDoFPZDeMnZDY/
DoGETBbPJod7MvWkoSxFh93/+n/FaBN/jyK7tqvABdAB5Je1k82D9E2wJr2kz5qY
5Dwzvdnk9VkBfIe+Kq6uZ6II3r7sHNjMjyEa8JZsII0rr6dOxQm5MojLegsGW4qb
QCI75MSAXDdrsYomH+x9W2kmsh1GrYyHJh2D1mQrCuWP/ohMIwm1mfNxNPsGVBHQ
hCktGcLOoffoXs2NkzYRo92e3MOPQ5UQf8iE7ocgNEwp4QPPfxMLdmuguqR1RTt4
siBAnKpR/3fzO+3vb4IlKIc2Fc4kXarWAF7A2lpzTGY1ETVNW2GXYEmcnDOlI39A
KSc8tpv/FkpdMwIdyaA9z+Bs1jJSEyUoprDp1tKk3OQPAUMgJywk20ayCE5ioi/T
wrpiJ1Vb6xyeMjGHvzK4GuVmLHE2d+Sptkf0lnBNK4dXY8DHF+gFr3oX2R/1g9Zh
tn3m/vALXluMecDkEmHhLfXVWVVcVxMVhNNm4rfzOlW+YAN5WjGnZ0oTMzxUif8A
ZYJzVIIv04KIdqFQeAPmUgNV6oD6QU1Mymsm/O2PqontzrYMf8Sb/Ax6HTH+UcIq
PnmqLcs3TB4EbW+pGyL2WPdFPYTQbxvKkfpwOepDhHoY/x622nV0oHa1BosQzD1l
/HXv9KjDu0xQUl6vnuMqpDhiDZn/hqeNMPHIwGnY0/rsJAb9WahMO5xmQK/KrYLy
B2vIdjCR400I4si87v5uR62a7p5D5oBflcoTceecrhimCYTNCfcFOv/NLzy8Iose
4zO2cFuoa5imwO8k2zVSureIt1Y9EgVE/kmN4VtqPmk6aMswTPckX2gdz4b8FU6T
ju3KxmVtxX+yWboIP/Wx4ZnT/uYbbktlwekgPOluuaKxq+1CZxbi2HeTGaN14IPW
2ijvy5b84PaWbVYIzz5IVAg22uJWDu0eaYBCbzNV6QFbi1E5NKsyyq39o5xquLG6
uICc3+euCUCv+0Uw/fei9QQ9qkJ6Ukj6n0G02dbas2pHtHQuk7G4Xg4mx2hOP2ob
FgeUnsIfVFYqpZIXfeN3w8HLUk2T3t4tn73c9Wo1lNdqoGo7Xl6A7ibU9azT30vq
qgZJt7Q+rbetFAvBaPQNJV3rCn65ybaZ0Rh4V/4Fj6gdDLDds5kD4kg8baaWwzqG
UEhsCBk81f1vrVaYVkQU+FfyHTwaGcYck1XoLyZKSOdm2dH76m46Vdf7Es86mOdl
LvoaAbBZnGa1OKNljaRQx2RyatpZsKiOL89lOiLRVbNUWFwsQKclJW/VXbP52L9L
GR8HyWP7NhMUcbByHv6JCzgWk+2dClqqhlDZubOwqUbtfBW5bO0jQfs9AXfsvEm+
iA/xlawZ9BPyQD+pgwRgcixmb61ZeIJILboSoL6L5ZyUTamtiMLVYKVcxPthwcuV
E/OzpXC2J3xCrDzJL2UZW1OuHnESYMkXqYYcX0OPEfGEgJssldiKe1NkEI4FitN+
sCm+IJPDexyJ1hIWorA+YSE0kn+Pfp38GdG5jsXuEV0Ht8PLRqY9kbEzzocK3ibP
fb+EVSRo6mM7VLI+hi5AzJIjB4PMU6yZRkNB/IiFXOf4M2td/Bi4q5B6MFw5aYTp
O8M+EGrI6rbhdM8svtoL7ioCkiJ4X0hLc3F1v8s6xPgyJ6aVKNXphOiL5st2c46/
3UJmVxET4vJY1s2GgqH6zVQUsZ4fzwEK0TZxvLe9eXPieFfY3EDd8O5FirC4cYc+
mrHvK/r56jYNI8RU8ECqESYI721ntlKOgaAgsvUud2DlT6URBDWwUvrHE3ajGIkD
oTW6qzcTEL0VqtI04VTDwUz8yi4/PiWALq2hSSDllQPV39dYQvWa1jEOKjir3gFJ
UYZtwnCDOBfNyJ/GabRkLMP32v0II7to9LaN3tGB5mNrAd7bCvurGBeV1Yh4CsTb
hR6Ib8OZatPEHeJ/q+TkQtONtap1iISLC6BcJnxmtnno+HTPRRAUGGnjRzU+sV/j
KJ7Lita1R8T6MoOEbAp5Lte9J75eqbZ4pJd8gxeEFeSBx4fqCJ0Xj6Yl0fDFZ1wi
pcrupEh4c2KdZFsT/wbJJS3FPG6uJg06MXTMmIRG26B5sM4cDayr5tM38UHz0r6m
MtRAtZss8+T2V/FkbLOe8RM2GOZYgIfTk2Iyhf+e66n3h6TpEIhxKselIPVesYO7
chpIUvVL+Q2+F+ENrTL2UNDABvmArxO61KuC0+7ffoYTahMW5t3p57Bb+RPk7zgP
EJ4WVaHwB3b+ZrkWTLagM7v6zcuyDR21J2pZJV1D+MH6E5xHi7UBrRgkY+wWeE7S
GgqoSZ7uvhtvRXjJ9EXEr+1quuXBlzauqRdSrGI8+Y1FpmNuJ0qDF41x+Dow9u9Z
viOblKYZqg6EW1KFpGGazOYbSMhII6dR1jX004OHZw7slod+ZedqDxGZORMArvRN
iu3tSuAMpBCmnUqt5ZX/3dsK2puKFua3SwkHevO9CaZNl7PX8HX62pOnRMKlTaoP
2PEtUNfqFpiFZsxOI7gh9cSyJ5GUp9+56DLAAp+JsIMbQQk463fkDFN47UjRYSJc
NAmmIlfrp3w0wVPD37Sg3bt9mUFuxYP8rO9yOIDOw/g+jIu5wFp8zlaTl7hkFO0K
l6VkC+3+FwTAv99nZ2wxrnAvVqSQZLC5uPZ3jmCb+8QVfJbXaPWxos06sOHJghkU
n1Sx+qIbzSWfaDNh65rlyCDA8aqnlp5MECVpyUKFjgTUXTYlIpcM9Z5HAq1Qoh7Z
0YFE2uhoGo6BsnN3uVm5K3PvYUtzMmWCDM2n9112+jxvWzNtvOr5eXL1Xh5OEId7
iolt4x2OH7wbKyfpJ9R1yqfh77aWNrc5w7+DQ8Mx2+Do93Lqj9sXjweHZdvk0Y4c
qLWYfHFXnAsi4vEfARX2fQPgbfwMLP8NKoTLEIsvp2M7ug/iLwIVn1OlPtoOl78L
hh66CX2CSGITN9JOcvC61oDSNzNh/jc5e2ycamRVpsB8WpGIElZkoCEVi7niNjL1
1ZrLvKmf5GSGZ57IhxgPvU9jfY17l7BMsKVuboboO3iTX0lmrgeg17FsbI2ixsWg
KlsZB+QJOzu3rWfTGyQqwHpZgfLhY4nb1IHCePtocNkoX8om27BFdlN36M8bCxM1
bPBmRiJFs7Q4xxcStei0eeur02c0RYzaKyNFo/fx+BnSxLlr8A/Z2gSSTM0vb5S8
IToAzZR6FTGmzovm3uOQjz4dzi4jLknqSIjU+fJmgTcLmcwk5dL0u2m6fLonuYAG
KvubIvZLt7XPQxhf5rwtgK3/Aynb39snp70AmdvuAiPKAPIBfJol9UwpTuUUhBgR
JrIQqMadEa7bBpiSEu9V7ljbJzymnSyqqV70KbgtcebTqwmOHh9aBZNwwnT4gOep
58FeUm3ny5rXTeRBOz+WtxooQTVQEEJlmKswh2//507NlJS2oLELUUBVXrkfKcXM
DMvElwjp5T4WJEXRT4k1bRy80E0WxgMofliIsF6wGCSOHUfiP0VADtSIlcBLEVzL
PlYwaC2V0nyu95h8tOWvz0d1KptO/6eoxsh+NA/EGVl3DXTAI3XNG35pCbbLP9Bo
Iki3IzRPd8pFNnM2O83CQHciqUwv6LznUeuTTdIB55LBhO39aYMozW55/zQ6k4yR
SvScG0p2jZnh8Vzbkc9WidAzD3AjEvlxRz+ydWWDTcRkUxaHmw+AiY0/FiusSReW
TzZvKxpMDlxD0tk03CpcefDYz8dfQyDoDCqU3T3HpOlx/KpE16sNvMfUWT8aJu04
U46c25g1lrfoVcFynVgFR3xeqWN9af9VMi1lJ9OeR9YzlkOnl0Jc22NDWvV1BKPB
T1kH7q7LmEtfhcXZ7gBjVlONCETCJB6HCi8uvwGopJ0fj/u2zyth5pE9FwNcDmBi
4VPmhgQ7V44k6Yt+td3ZAL7zVtlg8dvr3DWCOcLaP20GX6Dynhi3VUJMAeO6iKJO
5ys+aUf8G4wcuY4YQflwjgoUwZoB1ekgBwubTAOdUW8mvROVmQLkmuAWjr1JwyPC
BD9Lc3Z9Oqr96k5UGDsJ+30b0yfAzKDdO4mPrPZr3feNYLzju7W/tjqOzLDEsV2N
3jo8CG+cPXmoCGDX2wIlkDoUZlvTdWUA9q/ZFdThyRTJrCnOMgqRp/TRpnUhKTjE
MJSzc5VgHklUD0Vj4Swhjqj7POvJU2Re3ncVzLWDORQg04zxyzqKkPfUTDhSJPta
10n1KUX6nFVdhO2LTj+yW6L/DNyWikoi3xuUvE2BwXlYgg1UvgJWZEql7bC7326k
K28qxlDRDQyAnefyDdzy0thC2EBwjNR8saz1bJyYxIhoiTZs8MtR4utjDc2Y09P0
aFmEuirOloUXnqxQTAx1r1wqALirVBLFhK0v4d6YQkC3OeAcaQeH2pUVNmjOXUkK
m9mCBqTwCBApmR9BEJDm8dMPzS0t8DtGEJP/qg54agrWfHZSMpW3y/oUvmkNnBM3
mMx6ZClwi90hnqGb387Z0Il1IFBrqkmz2t6e9hh4g/M/LfrUB6oX3t5ntZxkD6PL
HWrDdIYUNU9DgNovkBSKAAS/dr1f+XUm1H+rc2u5H1aPJzCbKwj7w2+vQ0IPUw5o
zb9ra1URR9pDBbXhP1+sXSf7+rSyHyTJJz3EcQLicHS4JUi87kuiRP7t3Ded4sjh
XPUyBmrccNbTczAt3k8P+v4tf3Cgs0S1t9kHY5SnB/MMvtf7kRNaZMInNkbaIzHh
dUebJTZfSooosn5KqMCmYOvf6XHkWIlFVAyGH8QVmRsf1BifmyFDfAapSWoz+KCu
IZBNAF6r7USL+xXrq3ydthximJjpOsn2iRm7f1R4qua4VuKfyJQBx8RgsiLEW4t3
nl5bd6AHYy0zWNB0Y4wZ9fvR1MvjESpVTItR8Lpn1B8WWO0b0mfZVz/GHReP3vFt
QL2Pw4/Kyhq2+Umxc6bnaWndq5Ls6Ksdn2ZV82oRpUd69HEu8woBJtVNwqSk7T9P
B187peNDFxMIbBss2gOJfwP1JYyXDr3RKzXokGtvxHBeis4a2Y6bz9PhNbwFbmOe
RlVMtAIwVE5683mzOUdxTmaoJZTGMmYkMx/lgkL9VFdvEdWrfxTWjDXj3tUJSsJ3
V/uvdveVuFyEH4KMPfF+OrjXEcVTPbXoZJ92q6sGlBR54ijDN9bBMV8zJpmyWsWx
naBRP1nx7O3Q5XCMJ57MsG0y7BSL9zuNQS+7ZWRawOSE3/M3qVtMciYdMDQUNNTr
bGhNyJ31VnESNKRIKO0l3XMWLsa56HKL1FGpCudBtowG/jw9u7DslNj199ILiNEN
2PCENABzjrclmcKQQ6804IjPXsdUkPFxGs65Wngd2+uG8lERWXIZdjT2EpsL1RAI
DmHwTtkBQPPwR0OhIU8CjclujEZbOCV2BymMPR+XGpE4yV8Z3mAhSdT/2i5isyfD
D3k2v+NhMsBmcgbhKAPdXuwkiFhE8StGr4MhBt904C8ehB9RJTfzPE39XIqHz75G
MyiFHEySzwjBmF+cGEC2vV+A9Yj2dMh+ngjOwnSrtPOBje3BWrDZojf0gIhfjEIN
ZvMr+/Th2wUGJIVyVqk1eF7ZrmzOkCz/kBUO13zNHwvzTfx4PJQG2EqR/sKhDQZw
REXjrXdgA+Q7jgS7KmI2/GaQUYN+zuniae/l2BnDgQY+mm50NEGhEx7284d/OaAB
kGHwtTIYSZ97vv3IvRPOyjBneWIqflS24On6m31Kx9Sq1fofPlUtjpKq5dX0P9sv
yJ3FVkO0bgt3ozd4vWYRKj78IlmGqVaoorCIl6TtJqo67hBnZyLi4ZWiXAvr0fMc
5UY7Qf6WgT6mSiGcXVNi62QF8d8nSnCbh34x6hJLw6bA8GGrFWrLM1V+caSPR+kf
3wY0Kn9qo2GMIrc6yiyeA8RYuk1wr4/MeWjJONo4IclCscxVGH5eG1eZxWCw3CXj
UdYmdOCcH/JXlrFY3o3f5SGDWnIDzL6Bb7vDTqjKKDSiNOEnmU+Lpi7BQ/MvWjDK
ZxcjEtFX4Ab/CvQd339HGTVutN/BzqpVaJZXQWOTXuXsnuuMsxJo+32B0jOsPzBe
myvoBFnl7D0PglOcqPBRgqrPpJ8revCYNg016H0eUjMm4RMm9UFKsKpDlie3Sw9e
uVQLhZtn/wN3RRn+KXB72WgJRJFXDjrKMh9jFTuAnVaz+APQm0vHrRDoiS1ZYoSe
cDXJVCeem7+Qjfjogw7tJbF8gMzZIaxS0DqHbPSHM26FUKmFUItAe7du8uGZzdbq
d2VjQEMIyq+BrmhSMg+SfLOimm3w5Fkilb4vgPGNAd7pNZm9GwW5bRyGc6GgPo8t
obGQSIoZGw6jgjLTRy7WBs0cABtCv3EfndpO0J11ffFwq0LW12Bx+4l2+F0ov1xD
aUtP0sU7qL4RDnvfiZIU9egw3xjI5zIots+pytzeDzEyx6aZEin5MpKIQvdlOgh0
w3cSV64RvJxxWCy1wq1c9Gq17j/Z0dqOFKVQcV6C1TpVL4DdYmUH9A2Hwb+hb0WP
nVRxMy0xs7PdC9ccMGiIABqVzlCxZ0TiDPa8FPwUU1suv67hLaVmmT7PM3uweH2f
cFDiO6vzAXHkhHS/z+sCv4ODwDqYKQqUi/E1Ymdesm45uquTEpzADT6HIn7VdC+y
K7wh9dak/fpTU2PrmX7P7wSs+VwCvaof0W9NEZY+6u17nPWPuGg2oL7w6faaetYF
LGZCZ3nE4qUqCFcydel3mnPnBOEoae5CxPUWERBjpIw8lRL45luMPdAZZ/J9O0Qw
6rF9ptJkflvp6ou5OWz+mF/FE05PvOqHQzlc0ZtMAYnlA7ctDA3MkfAylfm2FYWT
Wu3ZzAu5mfEjtNqxML0dms/c6FJBRXYXbcxhmgy+v5bHoZg5Cnm9JX6CG//kze6N
pCUXSqT6EWkTUL4VOtz5GQI9yNLPK+8XAWrR3JCGMq34Et6YBfmO/51FqsaccJxr
t0RPOK1w8ORXGugIwWys2Gl6L1j7z+PlmuhqQmikwhTUus16tIztcfESP2eu/j8A
cnZo5PhvPHC6tG3QCz79ryzZ3PfVj6hju+2OOQWcNObXA/peSALIaIBXHiiqNn9X
++07k4pYxNcjs8OpPGthn8AmO4KOKJOp6RxBvgEZZbzfRn24H/zkzG+Ic+zbBLdJ
LhWqsmkDF4xZsTZaSVnqQOWOvAiI/KSjwHl1MeXkNTRdgqvU/7vNi0+DRCYaHCPw
Au1d0h0LCHw8dQAYWn1NTcGMTMwp0JlKoO7Oa4rBYVYvbY+3UpziXCdzqUrz+mNJ
QJsY4m9K2T+jAiWI1G1Otq9uNRAl6teXAhb0ZJg1kEs8gZoJYfrspnaxHzub7kri
IZiQoLQQAiQ4RLe/Fpql+LCo6cTOKCeHr4l04voye1vG2pWy1O15Yeh3nGBKkiHM
QIgyvtYI6b7z+MTc+ZJas17D2mksPNcjUdcITu/AfxBmJXUxHHaJJfldYNwvuC2U
v6Dyth5txnXKwyd2XvA8NvTFTrd8LUTHpi+s+UpD5QPEnyzTiYIMDRvJE3tWHLpu
hbguUhGr5ntCXJBCsuer9X+SWj4GxmCBkwx3iEAnceMv16PxOSB5EU6BxRrR4Zfi
tLyYEaHoJjTLSF8F8XUc69U+GM0g0mGM7kb8HFVRkwx0Yx54JvQGzpMyqN7Flsq4
XTizuTVwO8RTBKluKyhF25pavKHBVQenQxI4DPRirhMnMEEwnVubkKcO6Cl4rk//
HhN+8p0EKGw9RAD2aci2o1nAy/XmnVGMFx0Ki+bgbuCiXOFxH4VCyqpgy/bWRpth
csTXQe1ikYTOCJl32RhocrJHhcBNl95GySUulxT03xBjub7f1Pd34BVWZudoq/YA
nwyLBINnhX9VX9GM2Tu/rq1w4liJEuM7Zuxfy5ozBIQ9D7jhdkJCF7fPFggw+D5A
79HkRySXMb1atR8dmqzZITktyB+sC66/vSV4oGzTe1uESsjKec91UCECeI/SXlto
W5GLxYu/OLjzQ3oSqm1sC5Y/IBZHo15Gt2lIoUj+czZTIviZT6hAmpWCRwLrZS6Y
cpKkPj/4p89vDHXY4JS1jiP2rPgt9Iczpad4FYXRMY/QbxzqRnMkBplz2ySUT2pT
IAkZsjoG7WpaRvBMy40bWLKC6wOs+DUwHuXc7mQQJAF3XVkRATsmnpFKmRZiOqg0
9Sftr3mqiS16Pgi47V7up2am6l/NcYrI4DDP7UhwHNNhmfUFc6hwon1wMBzLOSe7
8ZdfJULJLrhD/aXkZ47+hF4s2+e/LeXozctPg2+dN4dChfX3k9K6QavTqj3ARiMh
jr9tGEb1d3nIEbq+CiFU0DvmXMWN/oP3RvK8zE936P/J4TBLSscRFwrOvKnTKNtE
D/7B+/25BxQ1iwbT7GPpFDQeTobtpBT8BCsyhEbiV6FEZX3uk+Rci6I/zHI233K2
8KyM0EJyhGmxmzIhd1bDqLCLghY749ObT5xJbMjokzBOPli3vYCMV+q0mVlH7pah
g0RyuIivL0DQkduYncaTyB4g9wLKilE/p8k7lL3KB/75d+niHJlX3VnKp8pzocGy
y8ql3gvo/zLNvXY3oyw8rjjrsdkjiqFipPqgXfAhN393Wm9/Pd4nCbUBYAlwLfbd
jp+NcxwmlQvxbmO98UYJaEy2cDySb9M8UNHBidw+j2E0gIR2CW9Ks/7JE4cWSr6j
6YOlgIf346WyEcpVkJSNrDDYYm6bdoYrTaqhRz4IbpF3mdNUPJbOq1og4eZHQ6pI
mBaA3EBLXhotabBmrwGV+kwMfPTim5uZWSc0qu4EMZA4Q4AxsXQg1nNHmG9zu+Dq
qVvZUN69pn4bVE+b25NV9wAwKEPwzXONVQ7Y/bgaiRokHhlq+l16LfqMeKX+XL7X
q/PoMPci7V/uAfgf2sAIr8TSf/uVzNl+c9MVkdLiVbfah9Vf4IkKgCPdlPlE/W1e
/9LOwv0bMbwRqUKcIUhyXh0USd8o6ylu8IlUD8HkVy5u/mrNB77ChhaILuRXw99L
3yrV56tDjE4G4jnD63qg5moy5YiGPl1EMaFPVeXKN07Zjn543hB9mQCf2eA3BgUc
eqL0hx5V/kZrQBHgaZBQYjuluhrQ6ZjECkzRBGwhkYQGtW48Yqes4A9YTu4BkvJe
FZ+W2n4YbKxrRqZwza2Mmi7hD8BZhE5epdPgB8oFBDNDXyi+PYgEXvtk0G4BioZx
hLFSs3hcLVbmDMPE0D/Q1hbynCRl1lnxSjTbCVsBzmqx1C4Qw3ai94o2qSdEjPxf
vGzNVLZUYOrlf7o6uj5INnmupHApcKAUbHjK7xx6NZY0Ipmxcpl0ZuBERzzm6zrk
Qtnpvlif3Xs7wAomPtSG8+9yVp1quyfy7AWTRs7Sf1bz33ZfgGohi1ZDukg00bLh
GSXa+rzkfF9KVkOeWAiZl8B+9h+wlRmF/Y3AYWk2eW4jW3XfA6wMKq40zHcxzWG1
c9X6NrOfX52eLYEbVp71WcvPvkIx8/a9lHCBiFqv3X9yYalcwzK4wuqyUoO5dkiJ
VHfOMaLuwtOikf+SLl04TRz6DjiC4cavFPv5m6Qu9VmQBQRzhueys0H3/VBnvLpk
ZLNoSE1q95OboiG+eHk6Ax2KNkQEGwVZhxuz7L6bBUSUFCiVlpvZkelBvgOvpy71
wIJ7ZRqOLNGkS60Ba9VC/+AxwJFW9fqAPl2ZL+1I3Jp6jL+b5+wsK/uv0NCWrak6
lNhLLoofyZEvwKkEyqajbguu95gKG1pb1LigdpMaqEzG/ObuUsticIBgMVYtt/po
9WbIGTRlpQpId4qX4T7NeBQuhj5NVJz/sA2qYXykTlOeSL0AvivAtwYbE4ZAdNdw
yTKFVA45/LVawYff/MRWdXxhuzswZGyzqzTazQZCEzIQMcjdF2iqvwC5ZhEUUh9i
ChLNKIPuAU9LXoBPGd6/vdv+LIaoj3O9HfRSepkXWaBrgKlHqEDx+u04W8aE6uVS
0LaL0jWhF+t5NQQzGnQal8iZjYuL4ZsxsXWzcN473YfH2nVzyRC28Uqei++BYpZe
zmGrLDwdhbqzhZWx0QYlw0wpC+Vz7Z929CWekrFM3Ot5UUbGcDwnYz3wjsFH6B26
nN64uuKIUQ/2En+/G318TzdYANzFKuIbbB9boHJWlwHV2E2fEsPYthBv8J05xflv
uKL/e4T0eLgtVdhNw1/e4XVt3TBtfHPCiOEBSf5xcAketjl6SXLGt5TSYvkNyZEt
2IthiwAi7LVzHkOa4TIOgjVuLjFcrtA0lmkjAPv/g0+k1RoBGOBkbE/jK8zta7mX
TJeCyaRuicbS+NNbP7pbpo4tGqjJ2OFqc2mSuGhqO4/cFvC7AGVpdtgoxK3iJSY7
ydBODu3a9JLdizht9VcEVMHDcVUCbLycSRxBRvoYE6W2kev+fSb+LTJii7Nj29+g
0sdWT8Gm1It0YKluJDzWlyGX/o86xSHzuAWyvDMpQGiqX0n042UlpDvBnlELp9ss
VsIwli/0t7Kb60jWCTDXbtTQtPKjmm0kDRNhtUMZMl0JoMsz7vHtAUAHXAkgsx05
Xg4UksJnp103vaSLts271IURDCUGsTYqxXu46Bh8/BAJAH7tJgE6pnL3/8IEiqzN
3ha8bMo8cUwxJMwoU1YDTGXX02K0jBySCF/pMvfRpF0fLn6UYliz0itlbUItY+i8
Z1g9zvgZoy2xDS2oGGl0fnM4cjiSLTwH9FQ2KavIVVUhlbuviIIPyR319FZwNR8k
Jl2DQC3O6FLUBnsdAkCLi7fhEtlGaTyXo0rb5orBh1yv1cVAfJ35PkIKf3Glvzih
ucAMd6jfWbPNcFKdhPAhBioyxWY96cVAOY1qz/N/aHjBWlKUputCL6A5HWqqoG2i
TdV/pIGbnxg+xri0TMOEK0Nhv/PMtXNCsgU3NOkOFEhsSkuO7+SylYlcMp3sZ/co
/KrYsJVSDZMkslHkOj8LpoO1eSh7SavXP0GlSyCJywBQ7aVPSUFqaET9NGV1YKB0
J3LY5ePNB+CFRBEVLjVqQguTV1cnVd+rWueilvr/6btPESnhZozsaGwmk6NiIB+h
3dk16Jd7r1HDjDgJ5Q1UNGaDeCTgOdtGNjK/kwrwXohY8SwfpE0gTpcCaoCmUHWr
JroxVEd6t/YSAx3DLBfcyZdW5LffMgjMph/KQzIjOAK9J+P21ak4YaesM5RLQRT0
BnqIzURlLTa7v50TCszpfYIvQKlXn8QVpoAXxaIpgq1g0rRijyVA9KRhGNhWhn3n
upohfK2PFlWXxJdluHlgPO1GJ7fzwSbtWmYWwq1cL9INa55SIm27fMrb80K+XH1p
UIRsmYWDiee39Mw8dWMIq5EfJCqZ1SuTmjjzoaTqpQYvjNaLgxTNP9P5gV3iUDJL
mltEq3KWs0qOINVPFgBLK111jGerv757hCY/Q/GKiZojbryJx4tD1OnbJ9Yqqe7J
VY5hhJ9nP4NefWYAZT/FHxcmr71vxxCV6qpH0T+1zObSfXY9skIoGwufNFBr2KHY
QPpB1qZ+BkULX/VmCtU3s86yl/bYJ892m2i6L8OKUZygvZDiurJKPzlNwjylmPIr
tTVmM76bwshJ2FeXWHQzP2sH1dLUbcFP2Ca3j0dDizOBRIgk2MSCbTklOC8HBJsS
T7J1EKuB+pMPP+GeWfUtg/UK9TnC2nKa+KPCo3Id9pcTIA9m4M5t/gynwhglEEHq
t8FM2viObBiLZCgW0j19y38tg0JrTGCGfqzRrQxW2cNuxt/pCKN/zzrwYN7sg2qO
U07xbkC8rhEM0iGMqgNoEO8f0H8mPJtK/tQpRvoCTLvj8CQVVuCJ7dZBBchbJSs0
0yzQNlNqkzITFrIrIxxXLMmlVaNtnKzyzi/qYPbuykqfKBUD/toa1RnjE6LpksFX
crc5rHSuJaKUPek+HJaG+lQCqyA8WmWxTKm+5iOhjJnZW5rWa2JDkQDv2hncW1bS
Ha832JsIX378CcOY8uOtfNrDannPWhaRokPryvEBt3+nLTi63hpHvpLLZOA3oCkI
GPezqUYrVebqsF2TAUoZMB1MyIWZEP8WTgr3vAga0r6h2Fhx2aCgWfusneTN2S8b
ddC+2ByPhBZSB/wcdAJ0sQzMi1gxVkQ79io/d8Y5KenKz52ph3dISLaoURa/E6S2
KP5NdML9sX3pcAYcZcIJprfEG8KMyvgrihZw1FRAfu57pXqXEMTdm6dkC3ZYU9SU
Kgq8fsSEM90vBO6ztXh0wBwIP7crUz0Waw+DooufKpJ5weTQXOeC/u3EBMLY8pkX
tA0mxToWDqK0iODRNtmphjt+FsiFSve6bZHttqlnJp3Pj61VMsE8trVjU3/ufC2p
E2U7rS/S+ecZlaUNdxFPEnONEZOEw0FmlqT0trGtWPNcMvJ10HJuA1D87gYG9PoE
OndVmQVtQoV8aZltXv/J72eTXpoEU2PllZIgiBiIO3m8GDS5OKOX+1Q63eKkeX3p
UvfcUiOTq1adUn7rke98wssj7dxvzTybjEsWmGBHTVy75ogUbKdJ9xNDzLwh4pPS
pIpKU26rU/N+7BDfqaBp9JosVfC+omwFzqSxAJQPvqpUDm6aeFjXudo+HKxo0lPl
tMeL0HwupLQVBuIwgz98N8POVdUXeToIfWY60c1xaB2Y6nfQOX+EFQ+OUv6zlwzU
8SsTzCxAjpxZb/g5DliMEwa27krT0DKzQbUxTdX0kjJbDWP3PJpQV53Fm+uu1pnF
rIv/yN63ih3VA0RVMxNVwKyP1DFX9ROQmU37ixnKiIk4jHvRagjOGY4/i/7CE+G4
0Cdq7EqEdWD0Zql8tllyVJgT/lFNImKW12VtrVm056hzzCHUT5yqH8spddqsJuh7
OASoKtekopwcr3X56Y/IWKOxtl78KsCr3c8EceELR3DyXynBGbtRTXUx0MWNFnSX
st6qV2WWl/dgmrcpkriiITXRkuoW2d3digLrJmWQyzl2+ObwXmHiDlW+IqTc3SrX
yNnuZf50q+uQFN2GCjGwiRTS6IQYBl7grSXii3XnfVMHKJ2EeFdXlAXkN9IisAFr
tyRyPd2Ur8jjyIcQwP8z+1n7Mq0Sks+YriRTB7O5BZlPZnqjjZnVawfrDXchVsie
g4IM0qPPNGL+bojPjC2oqdGxRT9uZCHDWHBN9rHvuiyy/HxCyQOMsUVvMQvqzogH
aC/yc2qnduQi2JZdpRFxgZahMPNlnCLe7SgQudci9z1d4kUPj1NwiTZefxGelzVs
MrAlJcgsvGJ2Aj0NNgvK1uz9ZR5bZaJTJ4asC2TdHjIaTEtXWPJXKxnMMfrlEJRP
JhossKQhs1g2M2gkEriZxl2d9uf2lycYYbHSU3I4d8QQOPJbbopadD3YRiK/y/cG
9AjaH4x5BT4Ne4iL7zqTABWMPPwiki85jIJIItL672THWRQQd7CyUlDd7byphiwe
D7g84n8+3+uoC+i0yFC+r7RdCgcHaHzukA8eSe8+euWcRSRMGJTq/TIbcOKbkT4L
0TnvFmOtOGs7ASyUqwrToMq5v7i57GaBUxZh2KMy+GGuhZvkjdstE6poq6NwMsiJ
EAQha65/lMIjBxwqVL4XTNfs1DSwcqSK3MvVqzzt6ZxE1TA6RpCGh1L4IAv7JmPr
vsFlcLIj+j4VR3S0F+Xnsg0GanEpvWjrh1qN9suLys+Gk8tZw8Et5NO6gg9lb++j
c4y2TvltQbTB31sdWOgIGiWZsxQdjIkl+45QmcCBppKVXojDbuY+kwcg876mWWAr
anE9+XstBItAORH5DnoRlOQyVYZfgFDq7w20Dtn1r2twXuEfiGEWg77xYqvUueYl
1WjbzTcnFupnxQ015DXHf/qLg4S2bhpvx9lJInrLA9/zcAS1eym1pb7buJD0GBjl
qn/7M6h/5sE/H+zLNlTaEuj+7ilPWUx3DZvHDmypagMEM78xjqpWytJNVFwyYKcT
Id6A7Eo4RFNFb/FKr/qmb0O5zR4igviwOJwSQaff1RQG6Wj7n/yM7PGruSVc+TlL
dZNYQ9icDKyMwnCVvNkjRpjw2u/Qpw80xOoch1dpW9e594ayTYwnszDsH1dbFFY/
UX/ZqX37CCDUJlukkixg5W3nD1X0bEgqbexza+I84DD71Xc+FjyjE9mbsGyavaRo
WGEBvg+5e1SC7FBcgl+OTi/ovkM27kU0l+n16Nlt0cbIkHelw9/CobmhHWI41aMi
ME3EmYxArNly6nxCkyZRaLPaJ7BPnM1F5a+N6OFxeyoLa5aBzEdGlMhgZe3tuxXg
mUODh3ocL1nRjbbmfGrRNrJeWhCXuFrr365v2lfPWrnkmOfkt/PgXO8PvM9XoDNb
zGD0LXMzupvbAHlaPXPmAjglUMg+dYRY1q6oVdwLC2hMh4BrYLnecIG0nOj2L+uy
Dc7B0TCiAjATUNVWRz9K+UU/3+3RPSFqTaxvkxtEKDW/evDIZMNk+WwDeOd0AVD9
Wycc/tc8Cl6aUESesE7wDM1vv/6SE2IrpusyNe/tcS4eiz+u6c8AXJ5Zh/CcEv8x
zyiyJorMMpu0xhJSlNnf9Ex3gEQR8psU0ECH1VKebrmXaVtCzrCj27FjKMjXuWGa
VfQNR4h+dwcPxTwWWtvQqdaMOsflvW/SA2UwBAaRhQGDQkTjXSOP0QbGdcR/DVc+
ivlap4PvWWTl0jo9BRI24nxiOLyK7io2bEmLQGH3S/KIgX6iuQ/t7ekyAhbMpcqm
JN1cTRqeAsoNuVKK6BoiaVFNt8KPFd3S172h/eaF8uJ4gWasCOf3/zifqCyPtgTB
NV9GMD15iMOOIaT9ZGPeqt9NYmAsXnqvMoIPsZ24U9nE3RUyBUvB8hvtFlY31HLs
ZugeFVpJpvfGlMbwgBuBcoDSacNJknc7bTgqRASJyKCCG1qu2GE3G9WjJjDJenxa
VEtmfqW1//lWm2WwG0ldyXhvd07zfxVO+arPqM+8003kPmwaQGwFRbikuY6S6JD9
gRyRtXUEdcYQoK/Cykub3GOZ5rd6aHNpLJHKMpRPkcwROBodK+LrszML+hKWeMVH
fBekTcWI6Y8nBIv9SiHkWwC4hFZQOTuEDXIWhNqoUIm0nrKN5pMGGm9FrbiLnEZJ
5OVe1uhw/kTb6xFhxqA9pYwgCrl1k/pAkQkU2XUPi1FeelSzKzvc7MmRxVj9MNt0
DgvlND0GmjgCbHBX/aFQPWq/ddxSR5u/TeXzeccT5TufT8bfvOjOdPu5Z/V7ItNS
ZfjBFmSSSrYjprivL2PqCQ+37bLCBTGm72Q5nSaqmjQgLXUElBJanCd4as2+v9ny
p9iZww8/wX1bti5Jct4ke6DYbnfFQmV8RE4VVcGT6358VGNH/tMZf9A80ZAu6KeE
9cS3NCOTTlsgm4Tzvj4pBqoQk2pygS4pVmMqJyj3TbGGMY8jSTRtc6hjkeI27T7+
H709fP/pHNp7vBrcFLN0PZD8cywfVEuDprvl2V839u7+dLSqw+1KY7/g5gABIDTu
eP8cA+dLAp4nTe1mWiyAq3keUJZEpghTPPWmMoA0rhrNuv8YCvj2FV6cdC1GwCs2
rzoJWkPohuuZdzfFvI9aIfbfp+wF5LI839N4tRQq/zaIQ3ZIF3n01I3hcUckuk/D
WX6orUdfUnTn9u/cx5uRxh/+bpz+b1JJ9SNStpfZVJeV8RRByfMD2d4107xEuMpf
jOLR7Qk0c6UA/ocM6cMH6KqNWLc73ypsQEmecdr1CoCImsmDg9bdAgDoDgFi33Kv
tbUsdTNU2RLflCmJdszVtdjEbW7cYoF1RlKnBgWs/QGMjnO6L7WQyuXCHfJPB7Wm
45L0YKpJtxZxTwuo8pRHm/rkIJ/fqpl/kTlUM8z1x+Y0LNhvrd5tsIY2ePV9Owey
lD/IysGNkXH3bF283EBf6y4wfyhjlyjeWs5CRY3HvOlZm/67oZFuailklV6xUU0f
2INvmYcf2I7U2WM+fCw5w2oiGP3JPiJk91UJUdrqiabfuqq6qIVMPs6QgND06K7r
sfathbloKfzcu2RXHZBJKcT3twFEHLfwzLzk/16RLcenrFmi4T49FKwTasY6OQiW
cU7LhF0olT2WcwR8tleWv05HbB6BptIOUkb+lTZ7MePY+iOPzoXyXI+a0+GaBDLH
7KIcTNz54pj3PgsP3Cp/dlWXm2m1Fd5ZZhmbn1ZjH/EI0u7re6AvVL0zdHeGontT
t62+L1Gw0w/WcPAuJxZuLtCr99HrDVJKUmBKth70/zOC30JaBJJ9P0VZNMQfNXLI
rsRxzQ5FTV81mJl6sKm/BLdzEbvuFSZeLq/3SxSgETXdrZmFNc20MknmIIDUfOYj
cj5Xa1HbI0JJYarA5Dduywwiy9ersYzwXp2lI7X1z5rklU/BY1gVBfYQYgSEOfDd
Ud8aifHsw93iqSWAGKnIDvbKMrQ4oMM50ELi4hKYmyFH6XWArRqoWVN1H8qQ0NJD
IvFiJYpKhVRdjAG6h0nbYEyev1dW0Y80zVPDWs2ENLJ9GN/b8cINa3/6RohZDsy/
f/Y530mT+wM/6wScX6EmKaAirPqPk6UayFqOqVgU79gsebhjjPfqzorrLyZwz2wh
sGpnBp78Ckj2wPySBzNqSv7KSHssor/QGYY3um8ZywBvcAO8VrYNkLm0/ElNn/dR
XgKJLC2hji7s9HoNYxn4P4y7TbU04Bj4Ts157MEY5EUvwoTxBTPTBV7mIK6kx7P6
lKtRQ+NZBZAVyGar5SYnoD5/zrsIXX9Zu/dMBVdqXP/oGsdO3LGk1rxMJD7ElBaj
hmN9xxE3V3+ncKFLKlAnqA+rH1ueHGr2tja3hEb+ZonzHRA6ynkYy2Hl1WgYllER
ujTTals9q5I2gvh4G9aQCWxcP0XqsxKvmOSG+LvPzBwHu5OxN8XJQXfKGpp6Uglp
f7Qczxg6vBaDz9LqSN+emWAYunGaQoqCWmmuiRw55/qCzpAxW+HWKAbn7DubJ4Cy
a3jZfQERj6YYCf1/Fd0XCMU1GMz6Mgp+eThloTFJNOFJvMDiMR8Bpj9PbF9ZvHSO
fyFqpyMk4mWTkELqXGMiiRyf0rJp3BPFiVz3zXrINCUsObL/szcdE93HCY5k4j4y
mI6V/GJhEkVU2aQrgK0ISo9Y8QQOI9HAVQHu0sK5zX9IdxnvksodGd3Jp2NAEaf4
+qSL6XsZmyQo2+9s+jcP6ADr/fl6ow2euvbcx17fTKddKOyVzlGX4IhyRK1P8wez
Q2soiUUzU8Z94c6KzBAMKmJ4CtIoToQkM1gyRRdS9lXqZ0le1ma9cLd3xbaRxQ9h
2PttccydPvstmq1pcD5XdrXRcudBzxn8UoTuKPmWnayXhaUgZpzkJy1wAYf4/g/o
o4MYvxLPtuV0DhVbsNpntw49qfkranIN2eQq7hy20J8arQmUWhSc+uqWK6s8up5b
/h/7DNGo1f7WRcKCjg63yg3il8m9AG2m9FPX5SM7aBCziY4guVXTWTla3RWcO95i
wg7OMwYDdWXhnbzxxohmrcZtZwYIm/Fpif1lkjAbf14fjl/+vw4juNI6tGcU5xn3
WKlYvFvsTOK8UnKGSSWRVxAQAH1uZYaVS4btzLWDtxxTiVUqeqwpbkehQOZI3qUn
FIwpmxxumt2qTJQ4+InddAkLLuPllGCW0afSWPvMinDoOLBRIsT4JFw621zrpsAP
+Rq7burDUwWs/F/2D6nGdgRhDLk4YamPl3IDKXBgTyTDBsO0zQ8UEvAkghLLjJ1b
fAk0YpIB1PNOKZDxA1Xm7sbl9EPNZXXdCFj8UOe96hKQw8SITMzgrvTMr4t7wcwS
M27etofb8I7rhZRfvKpcqpeN0TAQ/5B/LQgha0ogvzcLHOy9RI6BJXwK5V+UsLPf
KPf+Ct0Sy6UlY1eFEFQW+c5BAMtBecik6dqszm9mCaVA4nuOJO+uHmUxUbG3/nbH
Ehcn51Y1udewlfr3Qc/83XT+Ur8JVZnPQ3vKii0mAtv8gCKUtxv2AP7N0MLrEf+8
YcE7falINaveaa+xGIiMuEwQn+fd9skp+AqqJ/bfmB2rNGwcHXhZ6dLE/cjBujiH
aldDiLdyzWTwS8IOZdY7WlZa9blLx/Mhzc+u0MfoXS1UYv0vwNRrSmEeb3emVWZo
JCej/5kir+GYjCqSsGTa71FKwfRG6/hb4xzimzZg5Kk1IiTVC35lXxTZUAHK9Isb
RiIZ/rLmxI8X6Fp07KvGEyCuKjxf0mTT1m9XWBE0EPSPkCt0tDPPIHSunqyhCzCq
RhdQbxuJold+3lTa89nEXYWJoy18SkYNCDZMNriJA2TLUqhegyCTxLPA9v8LrFqP
dt/G/pJkTuZ7Nc/xwOUV+KgTdcWPsSqBU0BStFK1FvnSbqIu/GDKQa1mDzNwkSAG
ZUGozUab5+5iKWrQV6i0zEbH0gwk6zKUmqrxH1sJ5e/G0o7aOkQp518dTT9CLkDX
XF1hi1hHGnBGAK27DARPvyyHfamymOUr38uBS0QOR8UqlqSTVCVblu1Bu77Ssvsj
QJvDKZk3VrP9vuAxH26ha+q300r//kIyCl8LNqMVoMsDJ3u49kjpxaaFWlMfEUeJ
6ckpOCvrM6VEx1utVOMq4btdsYw83djGEHyI9PRXg9U5tLljNNyu5XNtDAhGTaE7
T8RnyBvlmtcQLPa1j5JPt1+d/dTpovjkl1BGwqrWp5RU+GOgLaWz1v1VWYDV5tRp
r2GZd+v+mTjuqyS2SZlVQPnqathhSEZWUQ3h3CDpGCLLzHs4/P9TUOcpKuH2uged
f3RU5c/XQvvrVjqpl4xzgSHVx5vQ9dWPhRm/aTumdcZe0y6tMN9gXlbm844kwVV5
iCoYiNWRvA0vEQdS49a9giYkaVTfC+toyKDzJmxkaY+eH0I6pmPW64XnpTSJWpEd
lhtHsrjGShwXEBRds/ShkNo7I6MHvZxjdKuj01hjyXdG0d5wo2kR0sy3qLuD+fTt
37xUUxPJRiiZamfGt3uaC4sxN4RMJMnZt5CztXvacUnnyHhHRKSVDV2i5fcXQV9A
Tyb0ddP/fNmiKTNs1AKgFIoAjHxzqGBdhSdLfsuKO1vBBhP0WbMvs+6HCdCu+VM5
P82MkeEPSESQ8mdZUR82PZhKzTiW/nwm4bkkuqdOOyDhC8ajYCzOXx0MDXsZMvBu
pO1k7S+G8jH9jCWBj2ejoT/HNcF7Fgs/v3aFnoVJkwFHXNMIArJjPhIrJ1bpgltY
Yv1ipHFlu5zvCDR0Cejz9nNQkCRPG4U31bLGabj/YYmgrUn3Tx2kIa8hO8P2LOj6
FzM1+tzE/Y1NzZwKZL/WNXRzioFeO1sMWGk1KWJbncrztFBEJGmuLhgpLczkqGdc
k18oVJsTdPCDlc5AiwtYcLODvPShRLMzOPs0dwkK1n5V7ZqOf9sqzTuEYZ6j/HdK
3XczYRsDzZj+kYuEPlq35V1aLsgEmp0S370J+NrDNTlgJ1DCg3Cs4mfDuUIrhrVg
QNB0TavFrikFLKVDEcy9XQMDCLzsGQmeWxLFs7+KWrPQtmCju1nutyi5Qkspyi3+
lFJV+paQ7fVvNeTYcIgoOaONNHQinTNtHuYbkrSpdEkevsqq6zHvY6mDJkL2hC7i
1GTkPmCtEstt5969CTD8Qq8MwjYcuXAIAf68HGNyxWZnHWjhkD3Hl59Q/128tTUF
UhXF/hCVG9T6Oc/pRPZajds507Hpwk3Ri8zWclV+Y1EFNQs7EJQb94IAdgzDgh2D
CV9zR3IbAJ+i/s3nAXBn3O/cncfWTlzFw4z/PloENP7ldIK2jt3WavoViq6jxXBj
XdrtgOBWQWr8oPBLbEc3RWOnrWl5j+1ZTjYNXtcy2M6zGpgMYYkb+SFh8+A9jhkk
M1HSJ3Dyb/dYIJyoKD70LRhvlqBBtzj2YqTGCfGarvt35yKW+6HkJr5JX+kls0Vm
v+o0wawBq4mbJcurIcauq5TkUv/8m9EVwCd9jhaPILz8dGko3zC7ldVkQwKwIG9b
ZwaALaltqZ7eagtQEXL3zMRYWGTPDiyHz+d4SkyzLyPntMwvBnJi9FxC+tQIsRI+
E1h51xkOMXa4dI6HvRJF2wUQSiu41cPM9eoPGEFheHCly8ftC6UAOdkF3FN9i+KF
2uwf41/cMWnIR4O6GFeWDG+2Fdw1boRBFL1OtETOtCzOJWn0rPe3IkglLV2s04P4
5kNoiQRqx2RpQ0UVPV69R6I06rgwlVkTvmJ0rlIQZohi7fjyKz7sgCOY/qs4rHRS
ZlR6GM41iXzQMkTG7ZOJQ8egh7+SQ5vY+2Hj7d9gymaqdWipPFOOsYK4myAkZecu
w+ATTElbs2f/+jmnLNQioLPdTgmEuVzxgRvz6LrSq9BpT/3gkjZ6NBY2FbekZRCT
FdoX04TL/qc24CvBwbeC+nTBhkq3fZ5AHwl8o7S+h3lR4z+ltuSQ8rpMekPGJXhE
fvWvpgpsYexRvbRtxeEwuQjya2OA9BUzyR2JrdzhyXdh5BPQoqLiJ7UNe/kmzT8g
ea8qB0nPFYkGf7RSsQePuEf6Mw41OSHU25lBi79Mbpfo18Iat/Tx4P/NORtRJNb6
rEaRGckvxETD8KYjuiZ8v9gGSKkgll83gcIW1i5QRbA1Iu0jlkSUoe/K84wlC6kA
do73rH9GWGdb787yQowGgUvd4m6vRF7t2JhERfwiYmcnJisAEyDQX7MpsksR1St7
ah/InOKp2ZBnDXlNML3E4Ppoe9Tt8GINesBAifaboB6BkVv3gy8b30VGwJjnj1qq
XICtZwSrPd4KcsqR4w7ymiXQ8/o1z723+So4GWE/ObB7UWh4OwwBVmcjcpjZex8i
ib06v6zLGg9vHhkMTmZhiM04wlmhNP8XFGxQAJLdsqpjYuVf2G8e80CctwaGkMUH
uBHRe0j4fFGffMUF5SiZfpn+gqyy6DlhR0JF4q0wuBRNC9Ry6yVYY2RrYV8Ul85P
qt4EtHOa/s6Qk8/EzJoBPRHox5HCqIOVbGwwQjlYYwuVeShzpQ55xtMI9PA8d9br
iJ2/43J0RAb9nBPYQJKkMAFn4G5rB4itU20icFsvLI185hOA2F33tQyrv7cFnBHB
B1wPnGcCXRjQD+tE9CML9fGFtV04zKmlZpx6Ueiqdj8Dk/CvZT50ypzn5SFQOaBU
QhaDVf9VVgv2lBcaUcec//J8nZzZM+5ab7WLQ4p2H2fBLRNwY7UW+8sx+U6S44ac
9UJQIaSqLDEOQV0g+p06CghO7yjMq+gQO/9o0uVnSpOOzgYGUlPWUad4zUNa3iWE
IaXEwxYtOXkpcXo0UAlYSSECuDdAex6+XQP3MZ1TAtI1fWUU5e4TMW0RrkYnkaZo
1tyIyrlYpY6T2bScgDDJL0tTYIDpNESOp7SnSzZjXPM9BawJawgN6/l5sgA3yHbm
CCYYUD5+OecRKxWRYUoG3L8tAvHErBIKHpIMPyrRURVg2vLUKBpziurC3B/9x9ZO
sXuqrWLu3fAWLb8ZL2cyp7TROAnYjy4cBUkzeg49WtPCTP+komyj9nOYxbIkIEYo
cH7BodWaeLAeeGGkAQGEPrnBPCK2azL3VN1f0850MkROxzfPiTnkgfVgPSGXcQ+M
O9CazNWNSv4tWPP8JXbhZxqOCO/Q8G2/ucV0MyX49B2aaF5DAGwBpkJRuCrilIL+
iWDxIohg8mBLO3wh+MtGWRjDK8X8e7Pyt+NoKKl2UQqhmG04s4I8ZXJNKUN/hOwW
QgdV3XhDJU1BP+csq28JfzUZztpTQqqccvQ/FerqeNFnKkmmKk2T7M3jdUlk7v/S
hgcJN2Uay0Lt7oXCpFDtDMFsGl37pdSz5WRWQ6nAysittmh8phUVzUxrkjesMSmt
txk1p21OYQYpcnCPd4Oc/1n+z1e/QUwLEkNsrens4E8bg7a5M6iYoCCsxdTlhAsa
GcU0tCaS1YbnoQNKleznFzJKaTunWHbqXldf90+qCzOiugxO+stkjMCBq1nCfnsn
9cz5LEHATv1YVjpH/Qkxcvo0sfOBswKTRXO8wyMNnh0jjFzFpy7L0mvtrtRbUTCX
8S57vfHDrzLcRkDLCOFtLbCLyZ2r0QOmnsBCYXcv4I+XKsEPzWLeNa3kbKyN2aoV
EzjhGXG8yH3nBthVvIWBB9uOUw6Q3f9BD1V6+i0Z056BsphZLJbReIprwJgvY6pa
+7A57teoW9ee6oPSNrTO7F0wv8JgTLH8gxaXtwm9DRDQTmcpBXxf/bWuwn72XhPC
gGyRssbumVNx3GNEfRUAxHPRWmDEQgjT6yA/F6ExeTR0Z/ftkvGdTf0g//G4NyoX
r6JJkmJ5yk6KCkFzdmJkx1IAu6VDDfwrpVhEeHQkH6cqFPQNKne+UbY5wSmoPE2x
mQhLL+o/Jn1wjgVa9zLVtryv4LGssfUuL5vqpQRKHhIK4pJ7Xd0LKRyoxW0+USep
xMVDK4fN/KHT5IifroxW+kHRhVvKxYSq0gHBNFmqZ5Zh8DcNBwfKXO0RN9IaKOsH
526q/R4IWRaWRiviwljFIu5nA6HC1MoYyxx+0VBoDgBODi8+SUs3Hy9LL7voHEW0
xtePLVMk9gBgv/EntaE5xqGa66zwwxPyyZQ1kYEuSRCr9XIWk0x+S297y+ej+ZIV
QkoIcwEPMih+84dY9+yE0IOfvHUiIO0x8zBhmWIX38m/gufFhLiOdKRc3SvABGGG
otEisKBRkvrdp9wPkvfkUVWgNHKGKyI/yPqQLKIjBsMwQxRywxLoNquPsiUfpx0A
Kz7xdsXQ9aHY5GQPJJPwR7dpUz9Wp3EqRJqywN/SsFcV7jofyba/9qRLMAlOu8O2
PoskH4y5P9mTEoPNxy8sB5ZXAHGiEFyZv3BAtCfFcgoXWOhScDjof57AHKFvQchS
5m5INDLostTN36Ybfegp0vy0cMZkGC44d9/6al1iaacIUspwO+8ogOA7FRO3L5GH
jX+vp7zk/rvgKu8uqweBueUEwQIogU5wWkxWREd6DYJGIZZWjVfFvkAjvpLEMimF
YOH+DdU2qF4dSB8POD6MeAf6un5hcC3tJtV9C3VzhOCWPKDQJlo9NilkBq+/8Qwh
+NduBEuyx/5Ncdx4yVZ2iZWtukE7l1nRENUtSDw8UXCS27HFFTyWtqYMdigRSPeX
PiNJ6hL2itjst4pMoSci4f1AvogwOQKMLs8luUEZcBbBDgWSJzn5qdpC4f50/4iW
1CjuDSyfnLXkVJfL/0AT/A24cd78Ky3ct6bA5pXwqG2xgfU7+LfU/ECK/51kgCZ+
aQo+CjxUL0L2e6BKB4RY1+J/cZWbg2vnjAhT1jYWiOTQChXSf7p2yTSpHfDlAEPw
PTUZn5R8PwSrJNQl85BUy1cA/BVCplWpYqTzpyiYAKuRvZj94pu7EUr+V3kGXjyE
3JVixp19KK0gMYOo+7R/blKhd/oOdilsBie/UOVPofkeSOgN68qegYmrRysqK9Xq
2b7pwm9Pe0+zeKNFDhbfaORN5YTNCzov32hyZwChF45PXbXxCMvHbRo5Y/wPVYgH
i8rvgi9r8eaCuVwYtNEB+GMq/95gFfAypFe77PTC3GuXixrXEmLrqxbdGeB8aNcJ
1u6ai8IGfOG7oi6BjmzY8QwhvXeb178pAb2Bsa7eDPfeaie+RWUuJCsEBqO/rXFo
Fme9HEx7tBFYaAi8eNqTSygUmvmMkmZlZBPU2fLQXUTDd/hUm7v5Javz2SkZ6bH7
etcWNLHIKkFyLoOVvXAyGzDTVtd9jRMoJSQs1YmT7xwgnsWbvquQ95hn9E5+CUqI
Zdeddo1zeEYgFz4cbGX4BSyraVj3c+tyuQZJuE82MOsmwxyDawq/E+MOHNvh0JVP
S2HjWFq3QHZXAmsa6zYdIk2ILrroTzzdkFUNFNVkElufl29tALHU1SEomdctx/VU
jzm2b5XIi7sGdM+xX75GeF9bM/iywknJvzVkfNCd2f/mbdkvtatGJGvZIMwZIQ9Z
pXr+4d5oOZL5qGMoG5i440EcZAsP7FrvZN4gvu8mHOUGVLpTJtUww0ADQp9FZ4PG
R09tVGE9doDs9u75ay0dIaNObwWY1cuDooXFW0FZfVURC4GWLBXl90XNVVn6dq6A
fCsJyyjRG+qFQUUtiEwOCVomKV0Q2lxWRYgPHht/ssrsq01pJuOQVza6wtFl/0C6
R8XiYgzFMHPv21Zkb5dGrVq/4oZDVZuuvNiymlHO/s8DKul9HXsb905zOFfdvx7T
/WC6CmtpWVVzfHaehg+VyxFXylvJCn2vIGSmXZ1rEHT/4SmKoEIfN/G1BjZMM/+K
FfAi/quglPGgmob0bCPJiM2brJghpQGOMyFKF9LHZkwso+c9ukQu3Amv5EIJvO6s
G/j8+1QUHg0KRaVOl3P39khl2GQn0lTeENqeLabWwrLNkaeejh9A5OjP8KELJLA4
ZjfNBQ8Rvac6g4PEcnINIJ1Kr2N2EcnCE5NPgB/yXB+XIKmQU1dbErwlEaRt45p7
1JExUfFqqCSp1Ts+YrLKJMN8+a3C35rbZJuGKaYYiVJ0v+d2Cc32sUNSULwmhwCX
loiDazovjr2d3h2Stv0S1ZFSTcPqg+UNt2GtJ1p6EehlyfUHrmbQNk4D0MeCfFLx
Elb04dG0nIri2P0EKlj5RF4/709xj0l3g4CFI/1j/z/p2ogl2LCY4ZYSy4zlGOas
9aDU558W0CRN0nmRJr/YwNnZqBCTuy67AcUnvJwxZgSjGeCDsgWpLsVC7+dKHEub
zvmUw2002E3cdc+84kkV4+/o5Ex54zIJWjN3zd9eztCQvDi/qp/hAmaYEh32PJpu
cWHBDp2JWxZCcB3AluteiPJ6rlNiQymt59KpHG44KqE17a0lcXEFaHpBJM+Ig+Tv
c8/zLxQjtVMflZ7TTgGrS9v6rrFi4u/fpG17s+oHU7jZu2Ioa7iIp75KF/j3TYtO
sh7IWgEoeXwKVO0G7M5fjFt/mfyxPS6IuI3SvP15J4boMs4gTUghop+pys6rOelT
vcwFyXFuKoSR1z4etLRupJJUdr/KPQj5albl2Bv59kGR2P40nGCOozZjX29z2/nX
W28eT6ZymoLd0lywglzmB7Hb5zM+XNUOH1MN1fNkaRAumr46r5trROEFrvNsjKYS
VyFoM37u5JiSR1MELXsn9ekU4vP2Jy72w4VUeKQdIi5jP0Zb1lVGB2+6QQisKaT4
Ehd4qcwtqpV3MYd15TQIwfV1coH8BAbwbGSTcPKb3eSfsEM4CUwhE33hj8N9zjLN
k6p3VzRK85r50EWqz3BDTu/eDBQqllL+db99OwQZPWEKd4JdgU9emm7uG0To5FXn
gj4O7uyn6mwhRT7Ba1GZ6bSTc6TujzWc8As0t7HaGaIU/vtU7dIUbfRJpPDpQ1o0
oDIq6b/4fPqNtDbE26uMslQ4PTWJVnJtg5N5N7DRWgidgY1HSAb5u6RJGpfj3iYd
Or+TrWYiEGANlGBdlUQvxtWCtnu9wv64UyZagS3MOe8NPQVrkq1tonP3CJPeGT1K
hcfUjToIX+O9B7/LhW6Lc23fQ2JCyCEekOp0Nz1UEEFIqdBjr6yUxIwLzl4DhjIP
dCcSIwjovVkl7VnkHFybHdtkwo09xbrrnsEDoLoxVa0UmiwU4PYPEAijW0BKhGVN
DbJA2ea8w07cNVvbjt9KlFvgF5pRkk+INMZinK2p/+FXVhlvME26VdLDpoqw8Yja
G9XWs2aO2GU0tezgiYGF6Ys9XwLQQxRSOqQ4pehg9xQ1q3/eqG8ixdpXaruuEKee
NJNPh3aJyeiMqA4lfk/0b796jdPbvPemdl1AaiAKHXPyMbMuKqusVGvrKzi76q6t
VUd0As/YhfGc6Q0yhUQxxEbb3SnTUkO7MIL3ZkqAzoFwpZdMjVbN1ZDEqCSVROnb
hYQ3oUQglWlgcgcqrP5ybJoM90pw41S20gruPVkikA6lns4ZLqDNKXghxq/wyn+/
Mi30tv+zYowoKtObsoPD3+L4C2Co8fnDEP8Z/Pc5t3WfwNzLz6ZdWv/aKBkFCE3R
vIo0VKYwqbg4NESVG6qWvjA9NWgvSBxaGU3Cv94Nk/mW3/dU/Luu8ZYrV4IYZ1fX
/pAKaft6agErhuIetyusqDu5rPkJrOauruPZtfW5LG5DXRyut4jBcsg7PIFQSQBJ
1jfsN/mPxYfU75u8I+Do19BIcwE28HdIraiC4Bd+SKhIv9Axy3r5kMBDQlHsFDSi
QdpDQxTuBX/PyMABrTREAPU4M3Qmy0k6Q82y8f8q3KBp39xkapYRd5dU/mAgFYbM
SHzfuMbXp52X582MZZwRLJHZFvwDWW37Df8Nfn1yLi/UAlT4WbK8DGP1I50Z4H96
BrMUqjqpkD16fZAIUbNr2dDtFMkjGSSH9k1geG34vtEGoC+3CMIWvHIm1Iv6JqLs
tkIuvmB8zqedtOugmknTCx+MCj0qE6akBIK2Tw6hgdLnlJQhxumz1cVsNgRC2f2i
S1jQl+zi+/r9iAX/Cfd/Gakw2b8PNFcbNuFgvOT1Uz0+lErP4Hcc3Q4Ojnt1Ov7T
yx+Vo6WwCLssVyDsHOeAkGuAWg2yJhN2VZSRj7nyk2H3qnupb4oRJH+CiyOYrETC
rC0q6nWE9oJdj5W17Qow9GQ2CkzSD9EdC9bwxhWf+jqkSMKXzEAiw/i3wtkqtNlE
CUrn7LK3Pq90+22drCEtzKJLtP8kwVqPuRnHeEDl66fm4rEJC9764yUtMv+9ct+0
vHCWfBfA4cUK8PmyPWxt8eNqPHDdheuExMXab/Rpm1fmTyaE/hNqWm4YTrK/XpO+
5wROCvxoT2eApxIE/N6HzkUVKaCaWwXlZS/8vSbD60ig8hdEvOVDXRFjbdnGdZv6
mrrCrQx9bKFrRD08l+QIGjNt6IfZIQPHwk7cGebpz3qRrarMmzbCPqty6zTBdI7Y
r7KEEnPJn2JMKxhRvRm3riBEOBTeGf1XgfgapHRvBwQV8KNVR8wz1jS41SNNIJuT
xqZZrxrUFSAjm1ba0vYXl2Xgwu75WtePGR1OlEC8V0kAafe/uCKiNUe0NAxy/L3L
/UjROmDBIqyI4gDR2ybX7maUGGw7rnIaQOZyECw5YfnI4jQcmQTqhPE67KOpLZG+
s50wjJAoTpD5/uHGBJl1poglqnfsIaXhlr1z7q/hUgwPy7fn9SY/PpMOj1rINRI5
m9qWHcrpnu/yVYh5RWBUmUlNps02eOZULeMaJIr79dMCLPlleb7VOeA9lJx33TNP
v4cOe36YnCQbbjbDT+rkCDibzl7QgZ0NL3cl9uUXA4U3goDEQm7RPvavGoOL8I8J
/FFBZl/IB8Z/oz0+qNDLCPBUn6NvFIGoYN0BZcZ60nc1ci0ZrxyfwucXYpcEsvZl
WG+k4buV20xDgeShkEAssg3fumBaIJFuaK3J4GL9z1q4Q+CBAor53SGpbLL6wYbC
d/C24oW6zkW5KmQ63tBzvHTYLmPhP9jP5pDeWirFt6DY6OiNmS3UUZrthjv7FlED
VJXRdhX/fTsmdBjmedFI20T9ceflVQeHu2sRyNi3JY4cDUlkMVZvzmQ+oyLKxWWb
bDMO0u8BU2+seXihixy0HwgGPD6v0C/nz5MI2rx7A8ysI0ufGsaBYLbLw8Y7c8pP
UxthujhMogYAniJ0ozK/pENH1mCE/2huPckJAUNRWIu6LYdb95Y5wLiqln55I+4N
ZfXKYk6HsEhGAiHcd7vCBLVaTLsOQLr0kVgQwuHT9vAjbQjJvot4zFO8xWhyp/ht
IMaMIg94Z7RnLKlRnXVW5zBLYTTM9TA5oxgCAaqBlwAv7tn5zL6ShqypImAtwvzK
Ue5O6MqjfWTmTdZZcQcXPgicKYwnq7DhQyqxX4JURnD1aEIj6wBj2qdTjxXkr+JJ
UNQUxLAfP2g7/Ywbfdju/z9GhVtcxdTted6T5cwP/uz1kikglDYOTnMtqJ8o1Zyk
NEIRNEw8eQ5N3NMgIGOAhiUzJ+866Lr3Bhq5SKTJ428Z5HL+3Y4clDDITS4uDbg7
oxJNt/8LFoqj7QKHeNfGI7WIurPGx5A1xtx9guL0nX+LNAjWbRF0/D889AlFTtDo
W3hWqs9EuXNWru1FeZ9Y6L2HHeBjFezyQD440BjEbtCq/KQ5S3eJsBusyH6H+waU
URQdKHXihowIfW9eEtFiJuz5jLVOvIaEKVxuQiGjLGo6glfvZylYYKkqkfBpzs5f
i4dbqAzvDpSW0y44vKdZY+4rhygNY+Neopapq9KojlZ9d9CQJkxqqb8ZX2EpoGxM
j4EJphMFiWvwuay8FTZ3n+7iIGDYQQhpgsymSyLkE8qlwb9Cy9KREw2WWtUhwIVV
KRk8Tei21/g2rPAt2n9YXxzJuX4SaV/ZRmcRjTjE6O4j9yu3s7DAMJ7d4FjQHQAm
nW9YH+DqQskW9xvJgT23zJ7FK5r5fjojHaZyxFzWlMyEikWeVhE/maXVxzGzw03S
cZfeuY5U1gJR1mRMYMXHjtaHTKTMseVB1Kq3Vvnf1jofCHQarKStUayovIX/HyaX
od5tqqImid4FIj/cuXrnVQ1ax15qUzXDbwvn+7hokhEfuYyG+2281Ip4hSVnG0JH
2czA4jHi6Hd4euAIAqOBK+CyBuM6PSi+U7+emdLFeup3wqHtTLQPqT/WifyoTXR/
7JhWTbtBAhsxt4C0wLumAQ4jF1Wbwqv2xmoaHwTEIvRfsGsnjfUqbFnycdSKa2sP
wJL7muO/Bu6CfQkOWv1q+rslzBsZgSi8bZXsxjNIbxB2DqPHDRtMRYFwl3UdraFv
imaqSZsO/FVm//yqE/Hmy2qPxmAMhZCSipFU1Czv4zpVKd0KNJgVH/xPdOjakPgf
p0w2KIwRL9Ic9W9vr8KNLMD3p23lIbqv+RfHBoRebn5IIx9Zbw/4qh3Vxiwin9Kw
f/FkPVNX4/36OlKR+k8rezxi0xPAQjKYXXjOF3yViB3z+UdGxp/nwiiS53hWw7Ui
sO6lbbZWBbfxitvyaH9HjXaMK7iGQMFUePoUDCzmoD0C+K9rV1ohAh1V5G/JcpLN
/ZD8CTUc8O4THnHb9dECzRhKwJaJpTUFouAEYu+BraxLht4BnAH1VLVsMh+ASF31
O11Bg3zD/sOuYs7eWt2BOmRCf7k2TB09BrgA7m1mqw5L6GtCxgltSHfDVTXyud7S
hsVY6V8pYB6SgBb3H0eEuoLqsz4Rf372ef5/MPJ+EFOA5SqvfUbRQziDbhhCefz3
rCjBwsdlwe9Vq5UTK+ryIafDfkcw+JsjHIBpEKh9dz7SMP3DWxBQSxOe9Ei5dmRe
tmcZxvbK5Ue7R4t+hOK4vaCZEBOhZPSFhxKXe1Sx7+jnBaNvLSeCIhSKiNRYxEl8
LLobyM7lRaItDw8CNFDHJvjRV/TUyWYu/fzmEK4I8tfNumsxbjkvmNx/1giiYGyw
5FRh+QBAe05KCdEJPQ8yoTP8iNHU2ydBhGddNGc2JAmpaLm1n47Lk9Va53KdJRsg
5X4krDCZa1KH80GX5blLmITsE9O5vc9qZN4tqcHgN6WeGNclBSDJ0aLJ67co2bgA
FezuWmXcYDxRg28IpJI7IUOvS/D7ut7T0swfCiv8mgccD+3dWjwxwDdRRqjAoyZS
DPP4Qw2diRAdWD7/pSlft1uYYi/8xprcDoT5QO4byXHkM+0nZOkNe4Hh8ipKOa7J
9qMDzpK2iEFTkcI5wrBifSFU/misOi/p05R4/h5w9jWalFjidKuW2nSXZA9WI2lq
CdQH84w6v9D5Ij3XWTYe83VThDDGXfC9IWq5Y4vyjMYLd4A7a+L/fttG8Zxngyrk
KqtKNpDjqrEYBt33b5PEJLLf347x60ggjN2UYXEOdce8taMTAyIdN0H+uZoKYLiF
Ne3m+RDpYOzVcnrkqmFEZbbGa6okiGvZpKWa2W5WTDgU1birvhs2HpQPeXltwr/A
cP11ARrxrKUK1vR8AkiRz+hBnTeKksPYBP7iLQn9IQAbs6omycUbJEhQI40OhbE3
FY7bkLHvAND31RM1IUzArFTZ3NznYKJc7XzA/s1TlWCx9/jpmVIIOFV0u9dCVJSN
RYmiy6ru5RhDjsH80NUJEa5vtz+i6pM5lbda9VPwfcRgLSUMgTvOtgvbactYEnOO
H0yZnxHB75nLA89ZYk3oAcI+qNjMqElZ1XJAqhN2/5NzBRqKe2jzYEsyp3xUo1c3
ysF06SY4WxDKxEAlUCQ4i7CIs+SkiiHO2TjI1RBT1Rp6IlB5X6MF+DQmnLhWGS/h
Iu2G1B9lbW/2ABLEpyT8A/fLFYzy7b9411hqtSK8pG3dtlwKJbsZR6ICFkua2V7P
N4h/Vdk/y1fxRkdG9PCjQLHpxVlzSmlxeofKaqAkO8pE1/dnt1w2AiA6D7D3POTE
k1StK1kHb7IWg/2L9ERDwr9bJo2eM2oP2Pz/qhJ662PSsGPadkslt7E3r5n8zqyi
kZcAyqRPRmlGl3SrvRapVagCF0eb3VKJ9VMkrjdN5D/XTTHcRz3/AOwzsH92IeLJ
aRstAUV5ScHFhQ4Yn7fXbu+c77lcJIfUHCMRSZ3IikuuhUUAG9AVaZOiY8bRY/sN
LAi4SrXTRBYiKN38ti+YqqCpmj4wTzUHKB1hRpFEQMtym5AzXHZrYmqR2b6afLBX
3l52LM2/IykS/DXRei8Jt5L/P4v8TuUp21RajtlH/1zIsdUs8lN1nQSleDLprwZ9
po1OHGO6MVehnFoatPa7nq7kcfPGPXvHhiwKhsf3rxGqHWuEkuGnOVexaiXi1CL7
A017DrNi12nqpOaCfGOynI3ncPYuO3pPrbI2N0l9YmjdfWqfFllr8ZIMsfV43WIt
kzFbUW/ib5SOmHWSYBwUzMSA09qPy3fMlnPQzkodKE7eaxWX4z1rFF+sy7tGiUBK
127BDvVR4G60JLKpU+563I8bypzjgYO9fotdoFNSd2S9GyQ1KW/PdIYShpvIHdMx
yiX1N+PcyyycmHhA3OJ1z6mj3e86YRpDK1CSWxItqeQTxgCZRI84X4ofrazASOcf
xVIGV5AHNpZm6b0x/oL5s1ZeNN5USFU+/10Caz+DZxNLBtjRoB2OKYrPhzMcDlwm
w0eQR+r/d2OZRePeVkMXcVLFphtnp/wvApvJOIzLCDDnIV3m6ful1RGxpMq6nu68
zIAqGClTOIt6RciUOv7CdaOvFQKoTrVTPCBxrZy/f5jqtOXENY2nnc13zb2/2K75
DsV9hLoE3oOBOhC8wQiKKQqgCD0XDkJW8eLFWqDh7ovPi7m1D4ovzWtHd13yzxNb
4ZBwCZf0w9AZt0kJBp0xOgjCdmvwmJOJO6Ytx1SOrrhs20n5rAVz2vQ/UMk7HAkQ
VUSv+/1qrUelQQbrseSUsuSTfh8fwp4YvMxvrCzonBtRGr+ywFYaypC70LdMnM8x
hQpL7ATjNpQsatirjNnsXoN2SUjq8PKkpeNwtg0IRzHCd+nlMiYjovXzEHywPAax
OA9r/sTWtR1kxgg/F6RZ4qK8QHlycLcCal5NDRma7x+VoRvvGk+6Hed03YpzH84B
8yzTbMgXbLVgZaL6nXkjSC5dtl2nGTLnmwPhESwBsD2gbZHHixrDfJSthCMhcX2T
I+Geka175+uMSC2lDCaOP+9xtdQrUY1wbIoMPgszKe8BKDMFhCMKKPucJ/bJKFpn
D+dvz7ii+/1quU/F//ZV3XILDrBiCLdtK+dh5dn+zl/tup+o+yU7gZ2tKeGu3fZh
jG3m0yBLEg1KQ5VOogmIcHO33G3QrRYW3QnVtdh91d39Xgb6ZnR8V65eQaka8EzN
xw+4vH8o177IBuIGVelfdChwdG7iH5uk9AzIkMRes1kxq7wG13iuUsLlzTeDDGzL
ZK55rkdGNd9154Ee4rmn/1m78JDocR3lkWEtf8mbc6k+Aqy/Pdi2uDZHsu2VlHjx
rFo4wBYzgyc0eYZESYUEuIVrrXMDkLMaHUsvEJh2g/j96zxMmMbWT+uFm08pw5bg
+OUuf7U99G3pNSe6KakYS/0SRsPXPZQidaRP8LLxg0WFQcWbQxW7yGIs4HcS9iAv
VPCyUx6tS2WkKS/9tZtebqIXKBncHA89ScSumqEJcaF1+XdigFg9rl0A65Ir7vE+
eV25XgJAI7ElYoZ1bV38MM3A+oGGB4DndkB5mArX1/Dd5X2KVgGmg3AlDi3lbxES
SSA4DoO7FrKsWm2ubeNio5eJB1iqgvhiEiprODjIWx1NAKCfe7KF1yLPzq/l9vAq
njx7z7KZq/6TuVuCVN3F2YfMT3dezoGpjPkd9bbgccpHoZrRbv+NpHWLPH011TdW
9w4sA50y0oar9UbOOtx4ycl3xvPvmluYSF1fKCLnMXYCzDvFrF1emc1WVI7ohD77
uacI0z8S5qb+gwi4TDEUakPQtzZVMcYFQfmU3r8Y78t0p01Cx3mLPxjqC1WKVkFx
wKxYg92lNeF/UNomCw2XpMekikGOCmqUKnDIozOfEXs1+A6sgMohmT9wqG1FUKSM
kSR32+Yi0UaIZpW/EwcXRsdvJfNiOInUrMkBhQmJkdhW+9SfBJ19J4189VH0f1WU
Wg1tT4nxiCL2Vm8dW0xQmslE3capl1/VQMWy5BgxY6kvZf/D+HM+vHqcpB8NWiXi
9W065PTWI+MFUfic5PDg3AkRVPG6juXVXII31Suo3GjWKSruop6ok+SFyoqI/ov3
XdyrosmIh8Riqduj2Tz1W2ZHX2rZOMvvlMf4NaO4B7TsRua8dbchRqoXev+nK/wQ
eLrCN4w+fplwvX2NHt1E2rd7O+DQXeHyassztpCrY4dO4MeoeJBqGB6CxqZ5kfgD
mzmKzGcHbCRBxpVWBEztK8+B40NhSZNiyOG+Lx/UNvBFtWaO1hd30bkNDVZbbraz
Oy+kt+jYkhKOW0Oy4AwrXsIKRABCRwiHuWtxTMFTKXjlMBLx9cwDcLUByDRP9iWV
iw5x8LtdUvNR1PGLzi87kTW9v4DXHygA+MODtQzKMZDxawNvEmRlmFfsMfMZGV19
x9sYeEpSbuPLyiwRfPUbGkSMVrz3q/URIkHm4RULMbCYkwu9g6ZClBqMji2v3+Ak
37nIufQmifKyYFdfkX1HIWLgHzGoyMsTmq6xVF7TF28CL9Ba5xekJck2zva/W6Zo
74cVNYxOO2NVW2WlbqvWHCPvQDanlwmzvBJaR/EEUiGddp/6XibBFVZmgYb3VKRW
j6HUJg+oiMgvfPexjzwsALgomhk0ZWZ4QsJdwJNvhpVGLx2jr3EINzmhD7+ePG/W
YOM/BrU8yoemk71zR3qK6wnEeN6KO+oH0Vso3/ElnbuqLSr8Mm5o9SPXiGWNoAVR
l4+Vtut85mCjcmLZuxr1JW6JtyazBtMNBD15uUto3U949lxRe6tOQBVofvENMPJ9
Ellaz4BQQUAYLHD111Ui9Tye9nF32A/VdYEeS1OeY4GiADaH+J/7r1tdemc1u78f
G6ml3JEi/rvNUgzD2VFGOKzcK4em/3LmG8AJFFyNKFbEv0DjegoTJHNalnpl330k
2lDzQPUHeiElLjOKY8MZjBZxHqV+DySMF9xH+wzUUnAKVjHg+Ap9tXHh8gOhOcy3
hczS/69xQQQIO0Y9OG/bVaZTg1Bv1xMM0gdavZeAGfZWxNS3y/9TRdHiOncl0OYN
qe/EqWQnlRdGxsJDmbN34XgWNJ31SyKfP9hUUGMRw5ozBAOlvhxbVUhe2mNFpw5t
a/4T8wsbAdDaDmVqIMCInqlXaGDPrxr0TBZjo2/zveCnsj+KcU4mYCEhCqqbovaS
old69x2kRYEV6IecB02uYY7OVfjerWUf8Bvly0WpBdIlWVoAj4MjwZO8kPVi6zYb
wOlXznZ2h95mf1P6ua3jqw3yKUgwT/mcIXezUeNS9w8Cy93oZJgKKt0KHvaDOGyk
lYh08NPekTszQafD0I/pT3kW9ZD9JdP2N/yk97tN4WHjpQfmWSwc5lgPNjnSzPd2
hUKV9Vvxz545YJZojCpeQhhrh2Pxknje0mHMpWELIJ3ki4ZhPdn1DgO20U8PN47e
vHpSciFYxxEpIHsrl22VjYhKc+z5xi6aCsbwmaPJB8FNVYrApEQ6ANJcB64Oiy5S
snXlNX8ZcU3XaIHiZhWu1WQbiOUT96KJ41BLxVpU4UFwfWuyr4Zs4XSScKDKkqFf
wHg4EOVpC6Oe1lep952fvdsFeZYoM1XUroFQrISUm25OxiMCv1MRoOgVhkyIHvhS
mUb2tUCpO7T6RF16ruzsJjlPwsdh1EJHbp7qEL80opxLti3ECuf2NbCAnQW3ksZR
BSC6GFXGYBIbSjPA6fz/0LS1OX0eidjnp5A6+oDojQP/zbhPWwwyWD3zXd8dmWlg
dxWWXs7rA2v/R9WolCxwg6Ygwqnk+dxNWyxAxFZfaqthj7fHVIBML0zIqSmT/s8u
hy/gywQQYGCvRhd6AaK/nNCsYBJh7XZLnSudWSklgMcR5mOdCwvOS8bEnE0CL+KF
47ZDumD2GlddWgzy+am5qHDM0m993zioNO1SaKb3k8KgO17rAoLmOe/JPnVeY5XM
S302ktM4AnbX/86XTDxwBrH4cbktDN2ezVZnxeGyWdKcbpfxcD3af4zAyuZCPOgU
xnmDr8Xp53i2tvJ+qhGp7rW1GLutjrjBAhWONq05chLMlOvg8+nZm3dItoIwdqcO
APAqoSaBAQft9Mk1E/7TbRQjI/qtndVNRSLEsAlSfPGuAESP1sjsA86CuRdgVfRQ
bs7lKU57DFIA7bbxmBV9c2fyutnXtLK19TRfSqfzTQ8ia69jE7mRDmYSty8Y3p2O
iaKa5+BHT9MULGK9qPcLUrXpolJSaaQJzExu71LX3SuvV9UxHHidqOqu1K578i2a
r5xpVBzT/h8ESidRx/Y9eJoAsuNFfVMa3WUNJYLc9COO0w2FnFYrXmF6HvLsNxAI
dRGrmHvAYGTS6nfqqUrAq8FyaVMNtMhYK5I07+qpm1muReP/G8KVa4mz6/+X3NO4
tsFHToIz3P+fTSONYu048HPNmnLBnT9JcNdABSF/PrWIvZv7KnL23FjoWWjxI7XC
n07PNiLGpxi6VCQXneERoh5kf1p5B2Rh6MO6EKR2PXy/JZ2e96gWp9JfjxZ1iHWS
380FNwqvabovqP7BhdrDO8+6ehkDF6sZswCCDTsCDegYxOSGI6uYtt07jEo4+OFD
egfx+MXmqoH/JNUNimxm92zqwZ5GowVx4aAqKZg7Ip3tcMe0ywDa+4vTQwvq3Pnq
SgKnwwmw33/H5+q+eosGEa/uwHnChHuq/0jbNmGdlZAl4ipj/R2gwwmhzg9rTVhx
FGvCZuOTp+LRv6dx4RUk+9KKP7OptVggwmvAIrX48wxLPlYAHvm37mXgvtqSBRWA
K64zIkJDJW/YmYrEYc0Ubb3vYhT009YsPUe0hsRqUAVHxNiBcm2omvUwIpxMRRlz
1K0jyi7Y3agslI8Gz8rGQ24d0x/KKYuO5ii7t3jNQtQuZ6Fg3awivBHzA0TBSii3
7Dgm7T7tu7fmc/2LJXDUptf2obKX3xtYbZb6tCOM800f0c34ja51Upysm/wqPanp
Sc+1ZbHhbggrQhGLNghX/QT0wv2rcAIL4zp1cH0yhD/wBYJ1BzS3HuAdcDg/UGUc
AKAWQtulLto321jASTebveSXf2jt7AhbllS6MamHkNDOTmT5VqYWKaB8bMaiCuRK
HM3pJRFVrVt5piaTJpumu4imoF6UrpxUstXuyZfPkpAKdBp0EXFkAXlBc9wDI9yv
9vOzwfvt/FOtJH4PQh/pwTzpCmAh5ON5D6losPhLetiHgAOmQn+FmbRGYHgfeN5J
yI6NmFxcWvz03vZ4mkd1vBpdbxOtlN0Rm8FhPBeiu6l+qYJ+LEt3NA1ilmjSnKTk
vzKHXwn3IDbmM0IJ55d8f036FIMno8FbWELFaSl8sFXLPSskUFGLSw7fOZQU2gEs
2e0K0tpHs411Eu7slks1Nawd5R1JBFwq/BZj6Ybcf1smDeYks9M2/Xq12Z0RopMi
mUQO1eclsOBTppnsPiRL52HAr2gyLNvkbKwwNvIp/ZdXHRi+4deqWF7bhvH+XXi1
BATZWpa7/3JQN7hdGtUDwcBlErqcoHPRcpLGKsmrzT28rNIoaxeekvQupKYtmvTZ
XtKZRDYN4bRUJjiS4dYGgUoBHCzSsQP/zZJbjiKdx6t8pyvLpizSPymiKJJKMZJS
LplsyVhMx3a6rv/kvwQ0qaEX1AUtF3uVAYg7HObZPCIdyiNUjxJWKnRXASu5nT4v
eL3zdnA6N+VCnn/kJ89ex5KtT557i9sFicA0cu0rp7nbQHKe5BQD5RUNUPu7pJMd
SLlOn2xAFPr0i0ZD6OUUExmNJto2SfgyD6wiiVSVYJViLYu97pnhqcNEcSOpZ8Gg
lE0h5QbCuhLQbTZmd4aRw9ZciHXSHDXVbWotG1UY1g3oZ3ymUF7vvxBxwo2Qjba4
5VEaLbf+XFWfwvbSwWwASrQt+ogZOyW+pGlmYqDS864/NbYd9BOo8cmYZtGjbYmn
Vy3vKHB5FtrXjw4mIAQr2X6gUFOtXe5HohSI7ooFoqKLhTCFC6fJ7HY153B9bJ8a
wEEc3cm0q9D8KDEzpQZGd4kSbOGkhlsTFF1F6qFMVIbsC0gnTBJEeNtyk6mJe+Ql
sicsVs78/AxCrGekw9TO5RqCIfinDkXewOUWH05vliRd8eSE5UW2MkwJRXKu83Bp
4Zmb4bJznGaU5oZ2toZ9OlCyIDHD9bFuEfkHEzoxiJ6Rt4OELx9Ie2w79GmB2MFh
AIO03mPden3I2HOYaIMcNnEj4UzjfD9VT68Y1uTrysJ+4wzXBGMPDJWVmnoKHH9/
z5vq84AjBY93/9T3cMgSwcknKGA6J3QDn9fECznhrqJeEltjvQSBdOTsNW7/tNN7
bU4QakXs2Zqy1FYZmedM4gj5reULzo1y8CT8QRJVmC0yTeZq2q3Hc3wFtyr/znV7
PXextxCCU83f5pYqzDlMxsTrd8cEhA+3JEp2Kln5+g+8Ucy+pd8tWK6fbC7RcqTl
Xoq8IpKnENmCNGSZ0FoCuy+sbRmTBgGWC/cKhu5Lxnc2g2H9w05E1bpyTSOJH+fg
d2db6iMWb7y64rm7Co0AlMepYPqXsHc/mc1q1qPYkjy17b3oeC42RRQrucR0nsak
WA/AaIvAFIIOTGzPDBQXyI8RIidvvcuazJ8u2Gc7zLJfjveykd5GEvUnDkJLOuuJ
3YV9tmpfMY/aBA4KF16ANf1z/nr3N1HZ/WtQTZ3KyKqN7oncUhwHxCyCowKHsJwY
PKT5QGaOyvHE4b/CrGTIJustDKTc/jSsbIq4yRFHUVRXisD3uJLflnX47ImMn4C8
kusIpg4FeI/NyEk8+sGas0wLtBAsTiBTS8iaPVDwxVhCvLzYQ4kPb4Vqd+SRuAEI
MgcYuSdwf1bwYc4k9hqPNGG+FU86QBajgeg25j+5a2EOYxp4Vu08MlLyWCTMPtuR
R1at//d1CEnPIswfVXDxc8JMho5f2k6LCU4BvVzu++GgTm5463jCUvCe5oxV+PXx
y1HEk/2tmOMP/MTSllgFrxOcKqLnNPDbfjMTfVPlFOCRCrx4aQ+4Jaug4CzejT9r
Tdu56arA/Su28Wk6tLK+qYYMv6Kv9mg+RiutiD9JN92p1VqxKsRtSRNhBznE2+Vw
YWdpBBwTh4lv/z8nEZ/Nok595zIsfYwti1ZGmxx7vqpJ5u9VBcx1UT/tk4A28PYe
Ok4BmEdNLy5YP4XuTj/ePQQgsinoGpqOvht6Rxs3Ss2F8dyHRwdJWodp10UKRcSd
CBb4vP/ZNLec5lBHQqJpDiBZR7TxT1+yAxcnfhOdLDE/J5R8vqmAq7QOWQMPKB8l
tLzIzX7YgW0R9thUqojkNrZ1Zeyn4g9y5ka2Z/Jupl5PCeQrqyMTpUdTwlzP/H3a
HD5fUxUGaHlLfnHOiF7RHXrYOcDFvYsNj4zTRkqspvoqbII652MyZHXpJ3SN4udG
kMPAmcfLdqM2ARF9sqEKJ+EcxZJbsL8t3i0UTCazV7pYizECzGh/Vb1u5esAP5uy
Uolcsewa3y5ZwTiKwvuW1bxiScRvDl6X2W+WhY3f0q47Tf6K6rgai6BRhObIQ0Q9
oGNKiXj7zdDeazZPjrPPsPafLWKlnzYnfNapzjV1OWpBTu1WHKXPaHhppPYESNob
rUBJ52arjhwqvQVGbC1Lt4xA7T1oBjnLTKmhJO06aXU13KhDX49BObbJ3os9qCKx
x3TGLVgGMXdv4FDJjHutKgwmyE3l278+se5S2K5UIkq1CAV5JJQDdSd+fU0CFsMh
pqUVJM/8wNKf+y6x6KfQUm+l61C9yrjqHZIIbNOEHHULfBoL5MAnpXbFypO+VMJ3
qb704rh53ImHrHNF684AJ11Rh5qpzmY/yetYXZijy+CUgTGppe66xRyLdZPFQFQG
iaM29Scw9uTEGDxFiZIueQ5AmDVlh/PMRaWXiSNxiTqdbryU2FPITnWrM1/XQqAE
P6L1VNKw1Pg2sIXVDcFOhTSlUcyH/174PVQ4rRy1LSsggzGxR0lV29huLAwasDW6
ROntQMBBNAuGAFY/pXM0bemRp9YAB03kCzTIoqQK793bReaOS+SHFxXZe15q6B9L
1WeTLUnlw0VSpO8v2Wj3e8wIA1ubl3ylOBYdqJxHwlsdHeQ6/V357XK6H/9Rr+Xe
k/IU6+z68YFZxPN/u1MF4O6MJ3EE48I92JggBxeRhTmulFq/7La9ZPhcZIo/9p2d
wIij/uPSWAa0YDDcZYbSmFqNK1EEoZS7froXNB1Bgw4yyILm+iTFj1pP7MbliVb7
bqrNvBa3oSberFzskuHNhexi3afSdOBThzZ0Ibe/LfdbphBdIWZrszN+rYOKh9dK
33ePMzjm63ml57jDeHD0JFvSiRaYpjAMcaTm9tWokd+V87N54LlPTUk2Ivm4P4Bf
vaVQ/Dd+U059xOIUr9eyhmxV4+4vTU0MMMXbXtJmcMWB7A7d3+fJ2p3v3+5YsOlG
MzId5Cw7DN8XKT2gksIa4lroMtqH/ML1rf23Kz+XvlqeQjTcIc8g78yHZO3lZh6M
jenXEZK9WHBYww6RfwWITcL6PXl4eyQ8sBBTjiMIyrGz7juQL+bJQ23nQoHIJyqK
ZNCdp5WI6udRzIuWam6sZ5qwDHZWu2J49Ptr6rbuqRYf+YKp6t0Y2/UESxcYjPS8
RyMpj7MfaaowlOHl6tvV8zAUuF2rBXmSTxWvZJiWogOCaD84o/sxWTDwCAH+vOE5
KmwOOIh3nRrj3x+myloxFbJlX8YxS+mshihAG5wwCaqZFvZFUUAxSh0m5T9ONCok
fXyGQC2Zzosvje5IRvOsZriUg3hX3jTHxaGnh8qfE3+/M3XLGVK9jERi+UCsbiVw
Kgz9SIDcclAnchN60Zfomfjw16czrzB8rKWoShczTu8zH0XKzST7XWBA+At5t18z
ZpP5v7uDydallZ9Zd9Drhn6vGRbTFSjVEwGoJ3Uig87mXFVjEYvVrDOslEfRD6NN
6pmZmAPVrMYtIJbGonjlCTE0xRuxWFJMPjXzCg9PLUe2yMJtOvw9PBgg8hbxPEKv
vWVIblq/aKb+HAiDov4VFJHKKZQEJDGmnaCUdDYDmzEiOc56YEC3zo8jj0LG98P+
lkiE+ggyK3bG4qIvgEY8K98MUoAl0y0hxiXwATAC2IamrLCyQMmgnoPJIRm1T74r
nzLEGAg2f7OLPYEESKsN8M4CjQ+LTLXV8oLzh/dg/UAlEgnTtt5AYXYjT+4f+pXX
adzYPoP4KALutw3Z4qBJXAbvRa9qxCUdYEZTb4PgMXTr0PJy413CBMjifqs80fz1
CjTz/WJ4cEXqF5F9TVEN8jGrbs9kPCdLqz+h5azPVxbB3UETIn2uVcrcErrNnQDy
WHui5tS/eLT77hlFkp75YZylrr13JzQxMCAtlJQ8qW9knjIrP1a76EdFoYck1LFQ
ViCqPMv5e6EPCBXb6RZTCd9kYp53O+U8JYb6l4nbminpjSu0mvsdoYdi5ebyCjqU
BjkDfcdMHCTN4bEjJIz6/3iIxaStVh15CXpL6412cw/k4V5u5dt+aeRk62wCL0Fv
dCPJo2X+wTj/ZQx7NuqYFAp0CdIQWLmfO526jyZK8FE6yQ3qJxEsvM8j8wjdR13f
SYETMOeLOdvh4PPlC0KQY4azveu3ITOvKLfEY7CkuS7hJ0gxkEevIkO4/FriBxJP
iIVf+18cc1WQEmoUJwHz9S9DB5XAHdHF2tvL0A9jYOb+fgLUSyNzmYxq9XDvtpRg
+KQJz4YL6zF30Db+2wBYpljebxHEpSgHuYoHGJhmDUJeYpBaGVeShScA2J67wBoB
bC6vDqUjE8aZW3ortM46cYX7P4W4el0RCmO1R7Jo5M+Cf9gYN90uR64w/2WtW/kO
Cc/hWUCKLTk+N2u3BbxZNGThZlwmoFThmYv9vGVlQwxgkXdWtchw//SJ7QaGcJoq
6ej50CEmAeCoHzFBqWMuKIn8zlCE5ynsUlSkKu3CRqwF4rXvl7595/ARb6ZWZs60
U3IuFf9WOlt1Xxbe+zwr/iuXtZia1PlPWpbEUCB90qVzqcDb4WeelR3e76yjIUL1
AhUwm9/0sbLo7RpR14X/ss4eLSdeaRhVobxn6RtPDG2N5KgPBL1c9g/ejs7wbkNT
2wJZBO/XyGpY0LGCfTvnbPdYLzir6H47b17vD9TAlQHDtHPeZrlVO5npWZNxN0Rf
pEReS1vlQKOFAket45sIWy2Jbje6kzsyw+KeEoe3tnLNoy+fbIqyWB+IsJBXqB+v
41rMtQ+ml6b0sc53Dbo/Wzhyc5JsftAB3yQGq2D1cjdO/G71yEk0LqVywTkZ6fqh
OGwXBlAYODQLysRb6GYlK96pZTYtk3CoUYInKiXGZoSTMUn/7gUGCd7r55qAQOFk
X9GFyStvV+89Jk9SoHOVEIZ8f43cEq5CTklBtepjnJideje+RIwZLcNTCQjw4K8T
AwJbbkLq/iM1lrDxl07ITLVxKHTcCy6K/LTBTRF2Enbb1Oa9KgCrFT52P9wv1Kzu
PPJcSWPVgoP2aqPVnVk6/i14ENDrjrKAi8USuoiUsB41Ey/m9gzQadWkundj3tIa
8YHRolnHZm2iquB3qVoo20JGR18qoWrSZM7ABBH0UpT8pyab8ehqK1fBbOyDXQDB
eS0ysqZM6vh22T8udJaVc1ykYs0T3l5Ga4ofT/cmeO0crktElptCa3s9WZ2gOVNj
2LPes/96tiQuNihmjwis73TT/0maE7CGIK8Q2XVDLginAqWDtzDfVv8vuCcyHIyx
aAbkymrNei2P9sHWWqduw87kr5HVDdsWZ0/Qs4xwqU60ck/1o7jwnMNaaqc6o5nw
rysveRfVnMG+JsAsj0xaYTw8tKpkZe23TEIjEVg7bpFwIQ5hZ1nhxSQMgSKnxWQr
/syb1CSMkOrdxJZ3PsobSqpS/JTvHm2bd+koFD43hWhAOEF+mTeOfg1Vzmxiz5/W
qKiXtQznPBwh6dYhkAbGgXnnsPU1VqJWOfSnA7+SOfKu6+7hE1BkMZVNtPgCwNHS
QaBunqrOoAwggJ4oZrcHcXcO9e8IvxMUo+GYNPg4K4Penk6Njotaz3FC721JpSvm
RB6agvI0HZq1bdoRI/TsdBYXN+sA4kSyh9DNqYN6+CAAhCDMS/lFpNn1zAT8rN3i
FKM7SqM1h9+Q/4u7IKklIxFB5oMgkzy0lbr7k0tlKC11RWJ9W/bTK6XIzcbyzfGC
nZDxkAZUi7FAxI5kaYE0k6PkI72YOXfTa9RTC8Q7EVNxSztWXtbb5p9+JBIDyHho
GKjvUUpwGqoTaJQNxLtuhqP9ZoQ0QcL7lYKV1cdrBBY+rEplxA7boKNjZrWKNsUV
BzdzgWJ2+h9Lkbi21432hIveGXwObIZhbxvMHix55y5wLk0egF6QT/H5JlBiWJuw
VS0y/lI9o/4rmkXT/brLoEL+JNaCUupsrQ1eaBq+0DLqWPJ1SB4BBzAs2yt7M6JS
D4Ukng05QSOjwSQC1K2ZxJ6S9RurU5nMPYTt1Rps7U5sW0rnguORtLKejg9s/Oxn
ftmypKyL0TG5U6GLdpvpngGqjO93nGEpWcCsKLxeI6htlJ1YVOvfh3KKVfU+4z5x
Nu82+8emvGRGBXGS/JCX3zwbwVKO1b9VATGMSf3OBLZO3O1qPjt/rtAba9eivOSb
/fstbFDIUPJNlA3rYmObHFxHfUrExZjokXxLJZYFexIgPGDYJTFZTZRV15BRwq+a
Y82rP47IT509/JXBxJjroAfbxB1r92x85pPWZpmM5Psx0s72tBQhfMeupuMbK0sm
9yZ6idJZ8cJQM41ZhxrojEpvEJlKxvHbyrF5hGCkEylOGS9+d7uXR/ZHJEcgZeKY
rP/otYATnTC5oBEQyFaqMrF+EdwHqUB4Eh43bL8a11K87fH6xUFljiNAMwXYCOrN
hr7nUsMJfHoh4N7lmQOFyV+/RMRGi+bkE/IIafVE9hQF+Eo04wrrWIcIoZgeIQ7U
l/OGHVNd7NBCtSHDFM2LpIokt1dS+4ggdtqo0gNIKoVCh6zOsPAsME36eTmAyz93
I+PClReEDGglGuiwTlSnc3DrUYLpsUD+AlFkxNySgzP0oGNAdd8fInPPuBVgJ1vd
sFCLSOSaLubl+mslBubJRJe3sXIfr69aRzD2fvUGHDXqFrvXayQEUwjiOsqzkIwO
gPFfd0c4PZevIX4wUu/fS8ADrHopwazik26T/9K5QrHZGhJ5OTPjbzhWVbQ9UJAv
BQrxPceJkNvv8PhH/UQ6oLNSIGrIZGFR84+sCh0fuZOmlQ9u9US/GLbsdsyXCXgc
fW9LL8byiFT8oMuRFHES/CZqSjzHyS8PiySf77YzChljm/fQEzPPzvyxbDNfC1SH
nLxnL/fG2yHTSaJur0ZmBH62ARc0BvLGBXxUcHBhJymXc3JEbyaXX5Uz0YQY4177
ZrnAkhAmspdHXz9qYNTBXjZ7NAZGri8pIZZnV755hpRewucxfMEkH52ShhvRyUsE
mzzEKoWXCDhEvIoJ2PcaTQgbVW7ZB1vrj521e5IC1i0jtPUkMURbml1AkGzc+FYX
k0vfj5QimvtSaAv7MCR9+ztNcB0hGYSjT/J6r60/rP5igp+hsD6klZy7areAU+dx
Mmn/k9yERzNXIjeoDnZpVFnk4lTH8tmP5bI2QAgVCYO8gTpgECj7klHDDXD0dRyt
RbSVOSk6Tbr3IvUPjPEXET0Yp+102XKkrlvcEn4rqlECoaGoFrYItj8Er/vAvo5n
LPzhUdqgaI8wDDklewc6ixsMlkcakCFSE0dO2y5R1z60SJhH44J+KkdnV4yxp2BX
t+IUlfT+Yi1GA358x/D2mEeXDVqMg/rvD6ePQXt8BjJko+SY3oHlGx4Kc/z2lk0o
7xSpcLZrFvxTOLCPDEk573o/kUUs7Dyy/k8+AUsvyHZWqSZRJs/kYE6PoUVI7x1W
oMLjnTupbbemg6H2ENOXewsEg8uomW5vJDAhhuRa0O2Pr0w8VoS0Wmi/iL8nMRk8
lcrUCUwhlXJinDpuQ+Yko0M2fLC0nCIelmbsEBv1xCW3Fj2lK5dvbqRf5QWZ/acS
cHgz/spCaABYJxLdhei2Ek+iOO9fE6YP2ixVnyrmg35tY/FrMrvnyX+7JwBcNNDl
/LJ5+TJBWm1St4yCfK3ReNFB5hIXv/3OigEmSupVNq4L5hoppD+QCIAAftjCLCCS
d34PdqnJ/MZAPxXm1zAhreXTIXUjwXyhp9DSyfMSNLIjrN7MBPJL3+Sm44TLgNn8
WnD+uuyw+s5cnog4bMiZCMCsZZot/sBTAm+BY7NZdO3lGIl+8keQHhH1av41njNI
4bS9HuPuKRYgJt6PBHfIvljHjkg+Rxd//8lIPo4CKsufe/AcxEB27ZvDyrkmOXam
cDlF6EkupQkEig8/6M0K1veSpUVBoS5SkmrbqjSUmln2+4UQmwnWApCkwys8WZIm
4kY61lCmNlMcnJeBv0/wdDEX8OG7gYBSmXgBQofjwFhXxgjESL+MMIEGjtCI3I1S
Lutxy5YXXN5L7XWrbacdteEeA0az0qx7pmxJTUSrznp3/IVN/ajNDFf1uSl33uin
SvaKOnxIv3OEn8uxJP5z0rdUwUTFU26GSohIwbTBrMNOC+le0GS4HBR7hh3FU+uN
QS6Wr8P7CIMKX+kJ8V4K+p8Z7Ri6xrXJpEs4gN5i2y76RbQlcag5pqXJSuTQ+SYl
neoQ49Ddj8sbRwdVQhstk3/e7w/VgLjsjCPGusb0ad+v5g/p3RznbOVCutRz3QEs
DyPPzldhEI4zjeS4c5Lm1rPze7gmluvbNcj2GIv3mEazjE8KRZfc8YOlbLb54BMp
P/jXn7D9kcHocG3MQT3FDluGSFW/8I8+QFkcBM7VDXQPHbjuR0/e4iVNwbMxe+/J
N0aNPaonKSNPd/PdmP9zonfY+YZ4bemO2JcfcpPVKXJTWVipJJ5YAGWi59XCz5rE
77litDa3mXESn5kK3fhSzQnXWHdZX1VDvTYFK87D8EJo8+pYT8eoWbgewFl1GDVl
aSyHXwUABUnyV1WHqHTYWHBe0YLT9Rh1gdhY8AL6KErIIL+llYgDHqnvLxzco0iD
8rzGkXCykjuD5t1EJxwK26OXCG9jZGyiBh2vp+9PCmBvIvOyqMk5tq+fg41oiyPl
uKnIrOrHJxsByR+ftDU9iIwJzj+Ot7BMsCJZ/1Fe0nBZ1EhAPR7RAvYqRLHC/c5g
zI0ufeBQvQvnnIQnOxf0ofWZ+iylrYkDdQTU1s8+toHY+P79m1Vor7EMZqp2BD9K
UOuuQIICJzYMIaJ3Z8/8OYVR7XLYekUuDbOPHQHXzfFbxGsWPb7KlfmWyeUjE2Dr
JxaXKmecPT0MwdlWG4UNt0CK3A+Zp6FzCtRm+Kt0HJdoHWxjE1fni/5fnhCJt+yM
mtvr4bjfCAtNyTMxWbmce8XVvVbaMahdD2J+6dH3C0wmd11So5et6GdhKvd9F/vO
Vm86C415ET2XOYzdTOhrhTdgdO4O+KWhZIXeFPV7j+vidR/BDa3GQ9fpqCQ4GeYa
Jje1hq5vaRzfgO/rMDzU1hAj8fMD5IQfzoFHTTSmMlVrFciAHTNzZhfF15Ckta95
DkBSBKoMYvu91fMKQRFKjhB3Q4DBhDBaavi1MTQWDuZYGvIMZhRSLwdFhvx7NLGj
fkgzAsGT0TgGd1eJMyP4CqrhNaMHeHkDaobzZTYfTElfrUZvO2WQHI2wbjvRolH/
2WdTjHZ6Bth/okVDnWokpPT11hQlZTIvFlOmhcH95cdqK50S/XpZopXA9I58OrF7
j6pmJpSfTrsicnGnRCwdAFk5/cGjLiRf5w1FcLiXzip6NhjnRtUK7B1r+OzxyOf8
qORKsdVTv8duJbs/VrrrdCd7TAhABYj4MWhTCI2Cg8aCPmU2+0TDW8/b0bDt6m8D
GVCVdrEYWXxl6dG06Em39HcpV0GKrM3JWTf7QvZAHReK/z/5Eaiz1HBap1f611Ry
/kk54/ZCEI7PJ6fWm9Bj0o0t1H3guG8KWUPrAS5Xv1RTq1brhe5evW1OmX/AR2/J
HLIzM+pI/ri0SL4o8F9NV0NX/qQpU84zeNOBs5ZD+hscBoHP0WMjVd33nAwW7Tbs
KU842Az9WtuDOftLQMszddEMfhKpglRTY3WNhWmdRYbivfl8S8JyUpuCoqCbjkNz
PsPJ/QAESzCt1l13MYKoJXoNKkr+x24VKgYLIeJDAnkeTLoz6sdU3KlBl37fHgrr
wKO5qLznRhiGn7albe1bgOgFnCD8EV6x84D+N2ywhu4/OjvEftHBvTobsAZU2Do1
fbqgB/tNXjLteH7UFS6t7aqAXs4bgcdLkVtg5cio8L6hFnrpjxBCZ0orvnuez0jQ
Jqr9Q3xMDGH+LK8sya1wtSkVyPvON1ohDJnP1+frPd6VioBOblyFqAtYU9miNyM4
X8aDJdh6czJBeTXmx6Ichnznp5usqzusUfGzga7lXNxnB4IBldlalE1TQqSP0NU8
VyFa7KmRP6VhMXFJVyEXdIW/wQNA7rOItdn02hlA6Q4SazhSQP5+t6/aMyzRdkgJ
mwISEsvEySAM8sjmzm7gqv2+OAzEjCFKLhc2xHjmSerXVWJWXr5ntIIz1iBs8WYP
VMGV0JhwdVQqkUow8ub/Pb56Q2CvqgDVyIh5IDQNPpGrofdGFfNBlCobH7XIRqtb
56OIyUpCHyoLRP4BVjWrgiN2dTt8hfPMOwFa0Q+cotvKghOXcgWhijJtcSlJY5aA
gsy2GRsx/XRk61bzBG04VXmBghHJXZAtE/QrHjzXgy6Zo8ZCE3UtmQ5SmRygSY4M
JVrSsZPh605x7q6FdNRHhos4DGMbhy9+KDyYzARo4y49Ok1uqfr13dADJJY0nEH+
GxfYVdNtIh/I2CFa4mgQaEFGXVBCZJ2cHOn+N1NmzqQgm5T7MClKBo5WMrCPHycC
djLuvVZTlewT/xMHis2p8dN/7amOrSbeyE/XHOZM0ScawekbhBa9Bs4F0e+qE6Vz
zHeKKdLgC49aMqsTrS8yJQ8Uy3pwWn0uIGiJlPGMhwJSH0A+8EYFfBCqW84O3F9Y
HfwTEWumJCqVvN4jbq4utu2S3/jN8yMQc6t7ZI8GkFOAuzoN+rNOtho0aH2XqFUY
u2WA2b9xcT2l3XDI2zQFrCHv7rSxye59Fw83oJcElYXJpb555+jwfsAz24qJZq/P
WwsP2wzEu6x2I96rm696v11v6yEw3KfwKfw10tWriV7YjI2MBMQ12iKv2Hzdsn2L
X9f2WoBE2/dAtbJQKfreIo5xOXo+o4x1qprK9h8IcqN6kiEqKI7db2WvL/89Ips/
sB+RVM9JLobDupSD+JhUUJ7XRkoRmSSPzkIzxcVTwrl8YD6ih38imZvBbjcOEFP2
UwrByFvCW4w1/PYZZnAH0tTTQFwyCCMj542nDTjLsSCbL3wYofhINGTAorxUQzOr
OSZwmT7nAhx4HD8NraPn02oqRm7HnVFuP8AYr6NjCDyXuMXiNq+HZYcfal4XpTGr
FPt68UMpModmPxPnSuqB25DC3WRIb4P5hRELMz3aozwG0CODtsFLvGB8aGGSyOfc
tEFCa3Qygk/wPE3qc4xTntCryNeHEbj0PHRqZoky50UQKrY1KNNcV+AxfgDyKmj2
owfHkiHjDyrnLH38tdSDszGAtBCP5/G0+WH14FNgkKRqQE2JAJ/S/4Fge01TcNvh
3Xie/hfhCSWkLIvv6j+cvxVJLTmzj3JVO0EuHq6uF9GjoiUiwB6I8zsmn0p1I38W
Oi55D+A8SISNJQ+wYY16RAy6E99a7SSHCAHAksqIeLfvLyHqSoIGpF3tSsHprJqu
WPEnpEL39QwXk4b9ZOXJiuDSTnU9cC8niSmVG6iNbkt3I1iBUXsTNEcDG8lf29Yd
lPrdVTaEfHXneUYq6owlKX3rchj7UhC5SUqL/Ndxd0pRjY5qhiLYzYEMMqz+u3S3
huzWealQVvC6dexNAkSiYFxQNd/nMUHLPpDcf5dFslz5infQ/vfSV41832ZD/7+G
xUOvJkMXIw752W9ufWVd4H4sWJ3A/byTSa8Rznbg3xBBNITsJbwjbvTqZrRjKzmD
BIJzHC+fx/n3e2+ch+Oe9pkCjcvngUHb19wJcO5uuml9v81RLFwgKgWwkAooo23O
9IkUj0bx8lAizsL0+LJaDJeXMFlKvbeOUbmejWmFdOh5SnnOpe2lgrysFUlk+vUx
T5MLdARHx0mqBJiqT8XjTigcQjShewFK+elo4zr5mT2zYud9RD63lVkaVMmc472W
PF/Mkn/W0Ms3RnIZGXWqe2arSmfdCOxaEFFWthKharL5xZTmY+PHAANDlZ+GWz2f
FWvX/ua9iaEbMj8kYkGzHEHrcXezklKBqSl07MTMpC23y2sc6tEEDAWrbb7/WT4Y
FbHxInRyr4eY3vmUyDqlgl1vp+AAOyDwouwICPlRpjQi5wGTZ7C/eblBBUvEea3U
LbdLfr69K5YF/kxow7pTfQ8539dDbq/YjQSodM+77z8rz/ZqedvVAlBzLd856B/b
dsvfDI+NV960IftTD/54EuGYhvKtNIi0wyx04KGIfWJ7vacUL6pWuZmJbgqG7wNA
LEwso8A3kGYVioKiw0zq7tKxpDWNH/6dvyKGflGM7lXxkIgprzOLubwYEp5O5X1E
Sry/favKvNZ9VOqzGOM43LK1QHEqc0EhjgwFTjc5Gd36qBg4szXpl6WUQVvwFlVt
Y6ADFINhykCH68n4ZUTe3l4QC+Ez49PomRa9dKU1mM1eGOBfMtSoXlpWNXDtieY+
RrbgNRzhy16B2K/aIfu8Od7OYrSNHi1Sml+8hXoZyAwvRGrV8NggBjNR2Kg65X45
SORjYh8q8l5Mhxg0oM2gcfCDHVk6pdP29XzGAd00YUdq0u3pJ2nsoIOfGtrTqcBC
FFaZd5Z52Z4AgPR+vhtJh2EldgyMaWhlUnYiHNeDDAmLKjI9FD05OSzzNy1yIEGw
fCSbMx/DJB9uwaSO8icEbhnY+IJjhS3UF0aABh9/cKZP2U8C2Kf44mG+iX/3pABD
A/lQV/34HAevC1Bl/sigOAgM2o38eCE+ibD/UAQZSwVllftuMCX9093NSkq5Al9g
abQCEGVIzHfIZYZQrAgzeSZDDiTIxZCMbKMAcwKXZjdlOd1aMV5c7QkkWQpj4bky
HS6FtmIm87DkzM4jaFrKGIoxgq4RPQ6z1UGb0u/jq0yQ7izmOJK4/qEClHsM+PiW
jLxGn92osVIpjE3IQ+PwAeWflUgC7ysG/aPSv4445fgXJZR9Q5lcDrwfAo3Nocbe
XlyCIF5owIKFYGHanzQLv2kfeIxfd2RYSKEecrmjAORwX6315bRbdHC5LOVd+g5H
JELxFHuSYcMBRJvnUv8HhCquQLPMOmRM9YUnW8zuq4VXwtBk7g+m/Z72ZL9se1re
6oehE42bwfZnvPBmFmpQeb4C/ggs0A53LbDzDWM/fHTVikqYyZ0P8RtKk4hyyN7U
J0i+iB4739GrTGgKl9vhIZIitGMI8jd146m6J8/3+mJtvXWzQxQqp9MzOPe1XE5h
ILAiHEpIIiSY57ZGWjNbg4gNHLX0b7EMamtAfvD6g5T9JA9nyoLZ/+1abDjLLGdk
fe1YRiVGcOVRqomMIaGGRtsa/yrLCO14iCUmeNE6SfK2CqHfLs3BcSJLu1XfYVWF
JTRAYz6HANaH9wKqGgaSFyfa9E3fM7rlJMTnu1o6qVUXtsosIP98na0j2iO1shWV
IIYw7IRkJVi13FK5bGV2kJiLz6km6AV5Ty4jgL6odPAP2tKLvFN+RVXiHiflZ+DJ
CStzOabzfv3lU9xe4ItbeT2aryI9jkzEszcjMay5Cp9GYKdm//E8IsuBqrOF6oQK
o23TWdpIf6LxOwrk4+HMRZ1wYWl7+Sd5VDL2l6R97Zns0CPnn/rxgWADXtgZeJMO
NwienVnEvUbXqw5I63ZCxp09vat++7b2KE+8pjTm+XgyAyzQevA0kNfdLFenQ/gN
kE5M0/rpflo6ULyS9ELpWzaIPQwjsFdKsQ0+EscCnDzFfVxKCEIMefs8rrlYnexk
2c/rzsFL+4mW7oOPEn7r1ts+yLWP3zCq8N6LapOFUuCMMPJMX9nc0Ltl1Oj4JA3W
rOdCf9N86ZgGBJh7PQsi+2mUV7qBMKlbqeqtrNCgBIAMRRfarSVa4IRj6S7tX2ai
knxrDBzDJHBuqwECKKNre0nx1TZUFHSP8AvMXpe05gmF43KjzBt6BUZEwOS/VOco
GNJrczSvrz4c0AyOAN6w0yruyK3JAlf3f2XQ/A9xUeRsXLCC3zHB0oNNU+u0xYMX
0B3NcVT0BKQTW5EZRXoIesYCS4VRrDTLPpCBqULQeJwtFlkmFl9ygMewuWQ5w4/c
wpLQMGoz/HAHiIF4Xl0t8hSYGWYVcXEsdSLwMxwJvvSPZk9WeIsg5qNYHhpLC8s4
aya/Z6MdYIUb9RmIXIBuPJH/wwQWVAk1Yh5bqzkEPgCjRPtEKYRVCwyWe2E5Y7Bg
Q/zoIt0uX9Z2MVZPI7mouaZMHy7gxGSiBMfdKT+gLMPqgd7AU35ARNUQdS6lMrJR
dclSvxLSnQoQHJJFZIWIzQ4PdLyg0FPCsGzWIBLZV2q4Bpsgwr6bTrw4LK5G4CXQ
VIP3jj/MTt9ZIJnJTqWopGhJP5bDCgEG7Ko/LNdgETt6+Q2Hs2Y5yUK5Q9d0QpMk
fg5T9tqVrXLWv1aWPkE720OCA/mEY+8PKB+FtLgr0ZZZKCuScFtJYN3ucZGQXu00
VttM+JbTLXw/Df0rK33a3q9q57FcIvS6piLn1RUPQs09j+Wb6WblFHh+7N9ejh7S
1BGVVBQLOqvpjtjrdJ7hCQCStDqIgNNMsKL0mbWQCNjWF1z6a27FnyGwcho+6rcQ
94ViSdEJCdhU9jnS0CV8pF5GCzDu0WA6cwtJ6wZ6CqBZMOmpuBat1j46VI04dJMy
Ju4A943lMnS41vsensonhZfOyxJfmzNikq7OuXVsE1o6MAfOLm+RddqeU1gtIzRY
ogzCXfPOKPryjRh4rodmXJ+Sghn3ydXnq4dKXxuWuhpMGYJMEuT6dLrNKDhTCDp5
6ma6lbfAD8P+pchQjDk3VKOouLPor05qZZhPRVFFjsHMoKlPs+iqX0sz9r4NjVjV
6xmUrO0IoXkgfAPxph3q6pOfcGzCexEbsFk0geD0jjMssyrX8WZBD7wFk2nLBCZR
WgqBA5io73PY+31MrI0wCZyOFDjrAgEKAnnrFfV6Y8pRIwghJhC/EFBzNkP2l/Wb
K7cW4G9o5VY7octTbTkR24CnsNRaaVGFhS58OfaHrAMq16ECH19OOpGZiF53C8wE
G57FJlKhrDyeNH2FEYbSUiaWd39wqokSa1GEqccVKvO/noj8L7DTjFd37B1C8BHK
CGFUQlF3bRABXxZZGPahg/DER3it2H1SFhmM56LPvJOyEj8IxgJeR9wVs6ol7tS+
W2vWt7Y5oQZ7u2BH7hQbJCo5qkTYV7nWbmyNVQ7+c0q3CsqWJoeEToXt4AuHNGaX
u/PFZyNMdoKM0O4hib3mXTGa7NKqmfANe1pZuHGVI9YQUr63GRZDgud6ACQYcBSw
OwSsx7ECd6gp+y7PLqHbKY44O9TjUXy4VcMawnX7dI4Z0xIoKaXPtOCJunZByN0f
5PuKrgASfw3HVhh71IIgrQWy1yXFMNXOlS6jsKtV8oAyzlsZVnkSzey546vFDw6K
6geONeAjY6cTi4egTFaKEMxBqtz7bN/TeCXIcjivd/RGnQYSyJR2Ins6WdQ9kI0F
YNlHoJI3gxaXZ24FpRZgx+P0aLW5vOEPm5f7vHXuhC7WcxNj254ucsiQxCN/mlI5
L/oodBkL7BOtQuourgSy7wFRG8RgcVdcSAtwswGAavfhigj2Lx1/mHWKwodOaGFp
tJcwAIgxflLLCmHOnNty2Q3V0+Z10tbgzHJr4ACW74Iany6IT85KSPsLJXUUjkGQ
wNYt4cjnU9dp6FGHrvvMbV5gr8MhDl/1cqVnZiuMmHF6qUZAUn7z621vVWNTvfma
U/sRZ7qytFLTms8JusTzajxcf/VC4PM+lD8F0n/yVXjmwBh08YYRhKkyXoNzVfTs
RXOCrcm+tdXb2bnoucVWU62j6Q0m/e60ecPLn9as+NVarsWbRUSWaGkUvbzTwUqs
H10lFSuPR2K+zyK9lzACGLTxANPhs2pBOBNIo4tv90d+w7mwzgNqrIKvOLSA+70n
QZXB178gt6QNFmnj7XGGSXLlJBfMgWz3m7qu9GIkhzMoN6pFH8klS38roUmTvFu5
4BFbL5LtOOqnw7rkdr42F8S81ZpL56FPdvYd70BhEJGPHOTAKdNI0q7NJ55rkvq4
ofwwRj2LMKDeJivlchgV4mnrOkWZg7lH6nykIdtd5j1/JN8hkRXubX+reUyM5qnh
SiYhwliZ1Ut4kw4aSXiAjhCSwFU2DiBzCwFjk/Or7ls/FrAqqFX2OVXvPI7hKJne
odj2RqJvDySlsSHOWx+mnKDtXVgYMqtdfQDo2pCdqUR+67xk7q8M0JrXnam3QrlF
Oswz+/vadgQVbXOVdhRtDinZN2P6u2FLiumYI7gbNvrgJmRWac4E1RwqVpitABE3
FOPGCGASwTrBD5LGTnIAP8LUu+zlEpEC+jASydoCzsEnYuds0LGeTf4LHNT8ngoM
FGs19LTnuENdzHKdD7f7iV04PCSxQG1f5utmgwFMOWV67qBW5UiYLyo3FClaYAxV
1uKjn8d0MSvMiM4XKK4R3ubEbzRIa8Qe4/LrE4QhxGCAFh8vN59csDGwcSMIreXj
jt3XxfQ8ysGci5omFrUMm4lfb7+D4HPVO9pLEeSlofTbt8Eu6PPr1aVxrN0bazFU
tNp2sBGuUkW6Gtl5csxriZj/kgtHDVZkokuuvW2Zv7jVMOKoWdxZtskez0og3lAX
3Qwt/MpBgCuDEG+06CdNJSjGUS15b1Ct3bcsS3fxAwZ8k/OFdvVaH92W3ATzTZbC
c98S3l3fD7C+yBOrk0/qzqJg80KqZjCQBhi2HRkteuzZ8+eYLZn6Ai5cPhir1E/M
CPuNSMkJthBlpgmLv3K58YfskQ1tCJZftRwwPm4dxqWMQyJk58EGi1QnztHVy9yf
Q+N6GpZ1aAqj3Bjt1VLA9pQWJPWe3Ip99V4zw2nmBZk0P/5ol26Vp8p5VxlnNsmJ
7BvXfElSaQxnbmsQKgBdzDamNLXaLhNMIhCGDEC556URkYDlQHg3ac9xWS2Y2D8b
hW0N7v+deVCWCPkpsmzrJU+Rjqag6NZsbt1xH1V5VBg/XX86COl7mzTySD76iF1y
qvEa3wSF5m5FkMdZGW5kiJd+698AFP4ZqZiDS5i1l6Mnh+cHc6cdkH92qanCyJaq
uA/MKOGWb4TC/nzs4lHsqzqQeW/xW25fEw9e8ylD1+zVL/xUmKrrmpbq/adnorLN
WXbaOOlifhBENpTyjr5+UruhZQlWalZNw6FPAgzSJHJIofev3PlM+wAIpPHoelRS
dwRW7yG5ppTbaeLJMcf96v/Vf9i4GV55gQ6TwMbcvpvDIOCBy8cLfoz7qHfEhYsB
h6alzoKE9DJWzq5lQLxFsivIrjDbdfefG/t6LkvtH5UGz/KETbfaYAHWW8qBx/Mb
0jBWY0UrXigYdNk5faBwQDNK6cnSuglJwPmaDfSr9Ib51MQpqmiOwtX+h9A24oO/
d+mMhgWYOLoXDhi95BSOdVRNMDdOuzCdAavzGCrfLRupYIHVTazT3ftO8RLAX+tc
VLLr9x1xsd4OPlOQ5Fo7YigUD7jQmGtmWP1+/PvmU3sAtMqtUTIVJn/r+FTXR3WN
FSaKcR/dZieIUaMv3eie+9D6vghGU2Zjwv+EKwppM0K9i/BMS9ILdjx1FI17JPZR
g3eI2UQHrKgl6WJ/b6mrVPi31eWER9y+OcMDgMz+rC4h11W5lvUBfF7Ip77jGG7j
ho89R0NttveMBTHk6OvaHd1zsG8yxO3gzyV3oB4eEnyxotEspuA0UzhSeOrkr3Y6
heitpcJnQWDjcVCxJGHSPSCCYY1/uxD8tNq0zCC/Ox8cyxIiQSBTdpDAXXwUZlcd
E25n457YgrsvYHqbeIPUm4Z11zzeTrah00SM3h/3mhMoYYC5zOi8sItMzYiukt3D
TbkRqvytaiYQxpc7SirIpbNNs7nYIyfGLuz6Ufztq1kyeXGcV4uxPKlTDY/o/ywh
HdB+vae3LbYkqUqTMBGPATqpNWPWq1kB433YA6sc4xMEnTVbP2sKFxfz1Vbv54u0
Xess3Xv1NgOJ0oZtVHjnQ6Rm3cUuu0rRtQoTRqmoKsZX6wkMQuFbzIeoZ0hvILVg
ItEULOvsS8Seuj2tzfpwiufkrkwTMWXxTlAKLQWDURcOlsbMJHRmzaGK/Pfp98yj
dwhF1SokppQDiw9v5lmZusBGc6q3f3FSyxxJzYs1oMzs2TtW1AzVf2CRWwLkQ6iJ
tNdzb413YvkSrQKKP13x/F0TDteAKsjb/dMxdxFW1e6SlSjUGHXdhZKlaNW8sfcl
ibN3wP5qJNpEAxcc2AwrQKKltP2fuggsE/00lMqQap3RgiMuJLCZ8dSB444GcrXb
+Ed1ZKG5AuJR6j9zKln8ucDHnYIioE9SGWr1yN8SHN0bldsSNHhFaXzVafeeG40i
PqM6CMBgkSgDZEBFxHNSoNafi24RMD34YG2lmPghgeonCIP5BAvnZEm8DKCBfhQN
BkqfukH3Gdu+czbwKpFJoH2cGsBngCik5fGtPe0HXQDbOalQetQVGXhBcEjLukSL
LzV2YmaW8I3TPRJjc7sQOKaTmoTTmeiQ6W2f2VhCY19/HDhuM3IwDVBVJbXeSact
GGM43LXIZpz5gfURGWtEzjKWUOYoBE8ff/z1J+qDYpP6kTG/Ahde66qlnIfE9R9V
2j9Y8tv71/ktmmM5sVF0fGh3GG6ovceuJlnARi98u7M1Nr2hv/KdLd5IzRedLdeD
VeNLqNa+R+YfM6z/upW0UTFGRPKdrHxf8gRsbeQJIr7GUnTXt7jOBe52ILjcKyDm
qDq7hbkDTqqoHvr8rJuJlsNj1HRE/kBvg25S5AVIYQ0q/8q1wRrZA+SkAtw2hMmY
SOeeYAcnQaHQ8BHv2vNVu1EW08FCCY6HslS2raKly7g2TUjIfJ0/FUmtXEjmHVC7
2r2JCFZGrv/GrFSEmNv0c/mKZfZP6JRerP3HnJSD0OFQpXrp9BACU/LYVkWDPpPL
pKP+7PMpa9cA6IV9/ghPaDZRchKAItrCr6x+j1azLfXxeq5FnRZaQ4BXkwTHLzyN
AO1xp/FgIojwJSrzzwU/kqNSWT/f7SYfPHTvAqv6pdsgBRcq9QDWUfxFSuW6d0Yj
m2Ue3LdBtwBu38cs1MckJhXxvUl6zz0ON/cl2IcB5rvw3GcDKl0JhtYfuxhQ7caA
4pwFh15yGWQ+XdJRFc0eF+Giw+8jj/PWtNneCobWA+PX8EIBE/lIIZfTK2sIPiRO
f/LzyA6LtvaWFOnbWN82H8tfN1QJuTmjuDsPG5MCJkjV0IolKn+MEYwmS1+NaXkn
VUdoTPqhSEs4c1gN2j9WAuezG4qxRJ+A+SKb5wxlstblooo8LuFyJefOIgIEjvfq
boy9U7HadUWOUGGh/QlhInZ3Kj7iORYjsRM6+9VV5YIvyMFw+3SO6ZCcqrfsTVDS
oHVy2Hhx5Ckf2attzDhW0vKT/thK6LpnHHY19eyd90e9vQgg2NF4aqyK+bZGAfoE
5XeWOk2rExYR6V976th+fytocOMAxUi2X8uNiV8JIOeOVDcbUO4AX/s4qBQu04AP
mgGMhEaX0h+ZetUIvNWLX7vqbKw9JWjiTa9bRziMUZlnf+eYmTfJGB9ZINIY1wpn
qaE7jA09uV9Td+WIlgOGrRjOzPhhtwbcKc3nJH1BeeiKD3R8cy6/Mi+qjdmMYC02
s40bWwIfcM2I2RPJnVdkC041K/R3tDePetV8tSDnpZ5lGG6wfps3dxQYT5flgori
NcKVBbSfvrGVGIEVerqNYf+CBE/abatqgbI3B4hjN4GSgWTRyDxaGYa8jFDeXCC0
/VcTf3f4I8fQm2VpvKvy8GnB4JRNAPVmwL+pOUoffxBqLQp9ljj27xlA8C360paY
bSOcZSw27wLcaaHy2MAAlSb71AvYBZtc4VRCGiWE5g70W4PGKxqxZ2AuPVRLsJSc
dzR6uKBEHK8kR1t+O1WFdnIYeNwzb3xrvlju+sO3bfOD5X9fNzBiJLqOLX8r+udR
2pRO+A9KOoUEDj+Bzzq7NXZVhlK9H0VHcBb/AtrE61jqr/xolTUa43Lxdihfgc/d
sYYAoIsOBIoFwTO74pc4SGtLNjU96Nl23i/p30ge3Ftc3VC25ifZKT1EoH0y8mHW
jzh3UpjoueavASp0mX3uW/RYiBHD6bxwkWT5WuAZ74B4yxjU0jCvPyyeclpxX6aV
BPqdVNjkEP65A2mXNchqIwwP1/pPH6vU9EzeIlzIVlyNbDqJRQBh8wyvfkvlfvP8
SurAII8N1QYE11XDp0QfLBNtCtfhK+KKBN4mUIZxbCs39IwYR4yD0ONwVG7MT1ao
0PC6wUkCSxnMORVzwHg2TsSd+5eljetKHRBVFr4Ri4/w+UgBw/ylHYFl9b46gS0D
skpzFp7Q7xLuZNllswYc392waay/Xb1VORVtWuCJdIpIgxduWGArW4aq0SoEytTM
ioKrESVZszv2Xo9nGt9+qnISKJem3qeAFLfZjHwpVjg5CqvLIGZM9Vd04Bscof+e
l1u2MH29tnTAC5upU/l5O0NgEKPfhjY7TiBXF/HfLw0kXrUFMifwOMjU5VP8Qsex
pJPwO3BUiv5zdiB1OlYAKhZG5jeZVqZhRvVm3SiWnFfjpESejyZn4QSAI5oxsy9L
YXEimJchG0iyVFt2zH+EFThLWWAeq8RQWZg/BVhC6ZtgpH+NglI65l7a/b+Y1agO
DVaR+FreNHK2B/NSR5AEVEWJHRsy8AS/hq5T2Gl2bUL9wCQxMX5yObrtjzZH08kb
9UZYeCsoQiqoan+F2M5lNF+E/LyTJMEuUJr2gYXc18sTx9aHjEeDTWUSIQbo1rTj
tPG4pR/N3O/1WPtHkrRgqgqyVu4bCXTqqWnHUZASyMsX8jzhCk+Gztxq4ouKUT/6
MXRK/xaWobDH+TVwdMhA/8C7dJRvvWNVK6SqRCNbYiW814kASlEBmb8gvhcEOKsZ
mpkCPoL3E2dRcDuaebs2dkm8xnfI94QYMeGbGOpVXGJGuAgZnPD4yRCEUcR1M7/Y
7LPGLTdcIlC4/RkVXf2ciUj+NS4Adl9CNQjtF370Zjgb6JjE/nPoYO9D7KGmgvGj
BMIIvSAhiuQsW2/59f29KSQAYxZCiocoEtkH53hDQz14HVQWOWptFZu23Eos5PRv
ywEAGPoReXbDhKB5wPpnqXT+KNLCp8ZTByproCuA45mtnDdfTutYYZgywEeDdKAQ
qBrHU8h8Foe+/QDBPD5FPyrq5mVKpWI/IHZpE2zC5KXTj08NwZHNzyRPPudg0Diy
uOEmbiKH6SUvlIPQcSV2z90A0cLoGMLrS2JHSkLKUr4xESwm3ukLjl7N2KDx6ule
wZi9K7btazuaHJarEmkUMWgJprcacNOZNiB0rrj/J7iRHPSjzAvjTtkvvwX/ODWV
nWmvVd5pMgcI5EFo/HsOKHdKXunMkilmR1PC48deI1sRT9hFDq0aGG0dRX2ADmYB
sJ5Nalcog8jS3l7IO+C1qJJ0AeWf/eXnB3rN15zslvNZGafRjvQFo0TdUk3gdtrR
47O+AXb0hmF/o2X73fnds2OCdKa1U3i+rVTRvgB7PqxYw4rYF2mYVIVQa7sn+tlq
drJpbOwV6o2xcCtLMN26+vCclxKWw++8xl76wuqLjc77+bcXH7OBBUrBb8j3GcBy
7n0iytr90TdL5rqRWB+qQsZQr4PNsYxCOHaUX3bmTucrZKdcnTmZVYn8QvaA/V5e
7TCmoYraVxr50LU3N1cK4nlIK5/GSQouaI+s4qKQxrhs/FuWiPTw1pwUz89ngOnm
56fVKkEwXeXGulMi+k643StdRC01hba2DFQYX/4sp48snvkvUiO9i/am6iir4xvq
l0E75S9CI94Tt+CcPuTofAEEym6UTiFsyNAz0JO0vCsXJt0LWXp2IoRg5TJUIRwZ
uXoDZyJeoyoSqmcdNjURN0r6dmJ80FRpEFJDAIJGM4eeXKir8hIFDl3T/kdNrNj/
1g8s2gI6E5Lu5LZXnPYOoKF6kDF8EHTNBP1ByzBUAaHGOsLj6+M3/lPqbi95Cwj1
v7norHN1QeQP3EZCtv9+zG+d1joUzPx2iYkN6gX+2AM3zqozv2B1mevRcAjYuVTs
etUT2xN6zsNIZQigCNxzNAT5NaJ0CWMYew4Dh6IwEYbd9jgRAE1pODZ8XBsjMNHD
A81cagd1awf8ZEVbngSZxUI4lVYy1XYDZMkyAmrP607WcLhpGWpHbxWIAmXc8OV5
y01Xvgur2TvdKAY3w82CBX/RNRLteIsj5ik0O6KbnsYNsTgp3f0tgTSCBC3LoRLx
kzl9gvfc8ZWXlhHf8tn2mzUSrHi+lfsUyTsQdy0vQf0yfReB9i9s3ZORlcgpKlla
uE5Li6QGJD9nr9cgbC2kb9rydk5QYbE1wmNKj5R4NAVeT793LrOAD0ycie1kNEU0
Xcxe2YVZ0uJQNvrU9m3/MOJccuUcC1H/KRllgR0UVD0UOZ157A+fKeWdQnmpecl5
Tm7NYw6WX2fZP4yYJ7y+7aUkdVuHeygrKAmy9eiYt0WDjXBjcxgSn/xcmXYoLIg7
Usnx6xLxw2MKb5Yc5Q/qUIMUz+nj4OiFIQp0kZP3+CoVEtguk+hgh7ASshC4XNNO
ZM/M4smmDV6IlvK2DJ+DXUeV4cEZCqKnnaG4vF2+QqC+V1HajJ33OeH7dBMq0lvx
TNIkpMjB0Bz6LzfkPQUJfkJv0PT7aK0a+lgCczNbVM3v3VUcvTgcQtpClVuCc9ad
Smw3RcOcwTOP/J2JDDwG85E/uyJOJAJTcT/r/u9gFS8bK6nOJPAcL4f7W8ismRkO
mgZreQSUCCHt1OSAz+JOKOBBDiVkeY2Uu/4ETIRK2jQQ+6OlumM3S0O7FCZ1+zKB
yg/eD7WRfxYY5IF9zTH6CDuevdJovKWP0Oon7bYNisdPc9cKHaAAMxprIWVfYBd/
FyTiM4QrEw+2T0RtKD5kEki/+eLcMI+xdhVQ9Kmq2/2PlF4L+NIgaX/pIhDXkdi2
EU+Fbx5xlWasef5cH6jQMQGgnHaNCfqdiropoKJ2UxslQwMkUihl+iL5vX/PnVfW
W5y1YM6VbjJmFdEAS8B0983ECqSsma6eFwDGyn6caj9x+QkES/n3LbQRu/d/7jnr
0VGEesHnAIHntTJQ4QBRQynqm/J80d6RWjhfH8NN9bwVv4l/ZltkWZFvsbKCt3n6
C6zYwb9h1s6Ybrx5UzgafUC2WnixJOa9Rp++KZsbxq37pe4PdJmC6yMTNqu0nmRP
WkWsnODMQ2jrYX5P/OO0suHzw3zyVDoJaubK98GS+hiygDFZDbbVIp4+yfCUGQ3i
n6fZe8sbYIUvFQQEKf2G/6emMg4D6DL3gbcV0mqk/HGl/zzo0MJ1HhiButfHBKJQ
mR4/Y5NnVLtKIzhEqCLGdjYp4EtM8wfvvIK3rl4fYkiJef1DcX3U09rtiNzuvKDa
2BlgulwS4orKzulKLbYyPE/omFKb0t6jx5zjnYdJUXYKDDqmOXLDtmCfNdH6Apj+
XUK3rfzpmKJwzs28GpfA52gPsGyHK8zxQrmQU05fHWBgfm0HLGRksJudBIDhFN3c
TOKeKM/ia2GmfZUcueKmkfs/UySg8F53qYiPBad9UkjUafLrfz2GGWJrXueLzd7F
DaFFI/Zdqa38STH9H+Q/wuyIxJjhQHCQvNEVQvBp3m9e9nmjKuMoC+rGYvUV2hku
wj4c7He/ICU/PcYfX5UA5xLKghXrLmb4kiRH9Oo9rzZbO1kNm4kt+a/IlB7vtz+9
BxcBjkvHpKOJI3CBAL3uCc2uDgruit8HUrQzoFCGHH98UHFc2xcal8w5Sflr9Uwn
+t63rupZ4haQVZsoQQCIGLKeoipvYQbrTeGUqCdmvxhlIfiBWkA/0P/oAtS8cO5Z
uSs4JUSVvnEt3kBEjPYzNxJohI4CT3HOjGrWpxVtU4K6CQbIKBpFRN0JjjXEh8sY
JINl9cfO+TVezdgZe7Z1R2wAGgQMuednY9+F/vvpSNSclg6JmWARYZVfjHYv9SVO
izSbYpHMLEjaUZFor6kqOseUyYn5OrHFT18MqhSomEPjNfqWaiT2jrHwNA6rFW4/
yOc+FK+sb3N1058LnSDfY3l4v9OVIBoix5Eeabr6i3pYHFkAiV1tJj06BEJFATfv
/enpTRo7DAJ8h6yf+5Q3qWfCy8ce5gFMUIRi2dwxESRZRCYdFoXg8vonfUpX+x1h
QgEDI75CcVLNfAGw4cTRJfvg08bYD6maoRJoq8IwNwNB6hNb1RXwt0fD9Bo2YLfF
9WNaUWuVEx32cpYM2/AzRdMIIQij0QAE5COPmNwTzH71jHrtAYEr/5956E0pTiEQ
ursJD2IUC8PvRCz5oTlaMnPGCikK2/CM5tGe4qmKWMHRPMhctDwk3T93DMdS80ek
A36Unq0EWbkDbQZCJnNLglwdFYCaFBvPKxMKat1sITf7z6r3DAWrEK/B2zuHuKRc
BaUW+RgsYoicb9hJJ5qtQtmvodmfL+HRSiBm9Ua9+a3W7l8LSOx/B+Wlp5ofd+F4
JXwAgqNvM9jOWt6orACuk3Sp8pad+ka/QCALWIOd9epfKAnmRH9Hq0cEl+qv5QrD
VLekQiPvwCTGy9d4MtHFEzIWY2zS3Jydit0PnEry0ta6B5hbURTiMv6uRmTW2JjB
NmqAx2GLsNPDltSUWIgfqHGMKLjG42pwWX8qmIn97M6bdbVkT/qgIdIKpeQqHdFB
XNscb1Z499dY2C/C5w9yARoQDCUjsvxHwwniI/2qTXgEzBHJ36gh08D2RdqzwthE
0SC/SsBuA7/KlxQ7sqfCJb9X+L1N5XH6OCDrSl2kzQvixl/p1oNakiIn/YI3nGVq
7r6YcaLwqVEcH1JpXOr3F/TOSDpOEcB05yz6qwYHjmiU+HK5Dpi5lrh5f0vzTqtl
ZtNtGQ21GC8VpyG4IannjHVRfzV5bHEKNem/QmTNXZYlHEmW93Af7pFm8M9Esecn
TNr5gXne3/+ojz+3gT6BXjc5bdybWYdcn7omonrDMxryzbLA+LYXPENNhOAI1F8c
r26dGcksKa7V/iYarskZqDbpkzS4R5JXKqQzUm06dACnOdGC4WkwSeLG/kip6bzu
fJT2cElij87epmT1W6m7MAd0BEjuxbNs8psLJIVgjOfNtjCWanzmBnfXtMevJfkZ
zQL0r3dEvd+v/fWncY91CugUHrwkVi4eEdEITAPSt5zVzuA32OS8ZDH0sCK44Byp
V82axsgnRTmbmzqt/3/OilWD6k5vQkPm0sg73U8UqNkfzWSxfg9fLV2TdrXuGhJU
LgH9ySIlkk3RB7MS4wg0DGW+HZrwn8dCmn0cAxdp9A0ykQD/PYxGKY+98anFRss6
eqvP4d5NM1a3/RcYZ1RqI99KdPTuW6KuONQAfOKiwJ/Th4whzkGU/TnSAB9o8zkx
C2XhKHWEKzZ0Gz42aCMSghvtAq+ieqTQuWuk6HVb0E4wAr5cXq06S3tqEMPcvuuk
VzVoOt80mLcu58j4fSjb/t5P2YNmxvh5dzVD2frqcmKvLht02tocDjPIGC/Jncfj
ePrybGJFvDSngMdLJt3V4e6IYHHyZTy/9HybZ76wbPLXYqTOs3nFBK2wP11fNh8V
lgctl+nbqMUCRG/2byveG9ewEK7QxgCFoKTLIRlKabYkaPh2stFi3fTgUcZbRlro
dMpxNpCim3AR1wXYJOWqvLdPKxtIUH/vkryF7fgqlqhpechOLzX2EK9bDbFId0mp
6nww3t9RAvEvDEfB19bfsT81y2ycJyzoWOGKLLqwnVUcVz4iIuZtnzof6DHWZV2o
QVw/HgF9+iN0vZZZjKrOwcO9gwJ8ovJs0YaPkn9vpuhCru8jTWZwXqeUJA5DJeMx
zUNmpy2GQjPit81NB8SQrnJXSo8lDomPBrjjkuwlQYnHX8N97lrN55RdXBOaPhZO
VPEfawnjU5IbnTjwvR8PrTwZzeEOv2ujwzA2a54JmjESIlTXaa39Ao4yj3xqmhPc
wJhnVc9r7sYyy9NDjiNMXi4oxgqEYWZtfkKKjN3eod99HOUM4fDqPOR+XbXTrqQO
hK1kFqfXf3/7i9Kpi9x2kFj0DoxDVivyazg9X9o8tXPvY4dzvkZg6DFxhRJPA73X
PWEQKElcEvc+73R9CDxsMXiIyu++DC7Av+XplAg+DJ+HjxhBFPBF5Jn2YiZzuvKy
D7y8+UjQvh+tb7eb0SkJ214tJ7x6fSDhWrICvHThlz3G+AlLkefChICL9M3W5q+K
3qyyXHRfKvzWbdRV/77OD+bVtcy39RPxVjlwznUFvWbzL5N5bmDf5gB+3Jyepnsk
3m2go9z21Br6NbDlwNSI7mYgEvyItw9oqYYIHWrHDKIMkMY1StZ4if0niJBoDJDu
xjVKhndTFpafIxHukoVSFS+OJpCLxnDzB8UpDcTHt59xCf2iNXqb7CzDZaINBFt6
5pbcTO8X7Dr70ZHV1ZHCsEJTa0h4jkNQSSH4qyOmfzKErXh4XfP7SfQDHWuCX/FU
cncrXjXNS2MnuJ6iUX9YdumyczazLmfyplHUxtJPuwvyR9cTPg1IUDd2UmAlwgNK
vXfkKq+5vlss2rCAm3Ja0UBMzyFa3nXnSywavtpCa7bbasPPjBkuEM834qTqGTE2
RLDeNCoVh7qT2JPYrMMrB0h4fze0zvFAC8EuXKvJ4ki6DcWYEb40FQJS76bsVkOA
/zs9w52ltxiWOX7NW2bM3JhHUbtAfl3NoTlD3cxumn9RD0E7Owc0rwZUEJscnACx
9M/GIV3B1zGDTZHHUQPBsRVn2TVwmN1o4ZjwvAjF4zwEHKdvQt9lvOIPVda6EC/4
h/5FBBfRt+Qe38K+6LKmqjZrnaFqmFhYtfN+t74zSswq1sMMvHrquh6j2xCywjcM
FVWu2SZ9WdVRIqkXP3w+k2Wnr81b6sWfhx1b02gvAfTC39QNzAvCe7C8bJH6RQ2y
hfCnRNfqbW2i9r2JdSs53cOoWP0YXYc2pqJEquIr7dksWUAt4yJ5E4575744hKPi
nSk8G7Li5zKMtRjud8HyM48Wu2atUtJyZ5RtOe75tEdH2h9f1ezBVpQPnhwtQkO+
zc4NZ/6pQiGo/DloIAhk7NJIxGW7X9dZpM2vR8lVDjn/9c2aeePLLaII/FdMzSQY
yF23YUV9nc240BNSFtACJZBxF8p2bsBWRIa9Ltps7cenXrxHcb39Z0aeHerptd1S
hVDKeot1Ng029Big/1nGBoI+qk391OAh9Hn+Ewj4/NCqBfli3wEy/rHJ9T9uL4zn
gXkF5hvweiFY4ViVPktgtp6qP508KOvy3qKIqsskDJGnFBXPJLPEXquIZvfs+Ltc
5ysUBp2BrxX1Z6wHoxHi5EEQXYw7BvvryBqeQQe1uR3HtNyW2xu2SvWY7PWMDuPK
DIyjh379BXbQwMjT8uqKdNjRmTOCYLNDEiowfV6rBatUF+CvXaXfkiG7xyHPzINU
3dAO97V7WRlWVofea8ymUV4Xj6+0CxI2n047OVvK3MQrjeD14nmid5vAUX00dSqy
zhrquxEY3SdHnn55BC5gz9aqyT2fGaCfKzrZ5O0f2Bu/0yeJrHfmHT4m+jQWNUQu
j5rG3F3fSOcvWBII9X7W14w40vTM+9T1twDl/BcMlgbMbWdZKO+utnG5jSl4Vsz/
pnlLP0Igf6UGea0Mf5uKSwJEkCy7rRfG/oiB8kOFuVQ4i5nmjhczI3fTz3V2oZjV
pYRNn9u12+7bYUvJfSDr3WacHOgE64pfiL982ZXkysJOaTyX7SP/orpgr3PSPm1r
50Gh5b4fR2apOJlFRayVLWwEB2pELzKEAQj7k2sfJXW0aF7SbPAJr5NWKvM1iDfL
SKU/Te9bL9VywXXUNlucmZnWA1aoSe12WRru/NYZ6xffOHeLdQafwfZcPQqSO8Gm
Q9Q3E6iAC+Q5eHennwn9Z13qKSdD7X6cSiRiqFZNr7yEVdilpYXBDxMLgq7o7GLQ
QIxsbXUWhW+F63zQ7oM9NtGq87pPIvqAqqs7jLBkDMJvU1KxriFjIjgTJ7VDL+3F
GrdYGe0GV99sORq1AjWIuwQ3qVoV49tCVv+Po9hO827Ya8E/LnRVUzC4otmr+ZGb
WuTOfaYY9azo8asQI5mDYiljelb82iZRjq5F+blY/zQOmhkkraINDbboM+v8PCmm
bGqYYwnr4xm6tIsyquWo0o0E4Ud1Wb0rTijpyaGR+MG4JECr28CGHsRNdel70jRC
kG6FQvzzeyGBeDuJGKS3fsQY5YvhLRW0sZDm1/YPh0BiDqgKKHHofEwFuTjs84zv
DCSkmKPQGARTqxOoXdv7/+VmGp0F+rT0FQkfqipzsOGont14lvQxAMya6EM5ZsQK
1XWGTDn7buAa83zO3kYt9xDYBmE0pCPsMSgfHHUni4cM6T3/EPNPWe7VwpP+X46Z
Irn+uukAKXLreCG12cIE0V8/Pp+Ihh2P7BDcRZF3BpABNBVv8woHqh7eLY617OYi
38UWJHHM9fJRCWWRQfXXPYKKhEtFivlse52RK7hUTKwxmiCrj60toa5eBuY8KQlL
4T0sxLlh84xxnTcYCv9nlhP4618qbrEyyGC8/ODXPGfxPf9BHCmKTM9yhiSdFkhr
SPw9xnDHHVI59xU0/cyk8lSjejS/kNy+5kS75qWrAhpupoAeUa5rgidZVLPP493b
63IwCHsgimJLGB66jWeG8uW12Y8q7wPEFT9uN//CjYzfXakc/2mZR0IlUR/Ds8pF
XFYONvtaNvqOazQ5KlB77/OkF+SYJqP2iZ99UwEJbylgknWdEpfDbTQ8xDIP4bvL
4StF34Fa1RJ/ie7fwDJdLnch5hNoM24fOlZQdvqMhNjhRTaFhFUA046/LJS9lDb9
qP6cQkNdT4LnB0+Yn+Rmlj8w2KOpb/Ummtzq39tQX5g1zpSTMcbXmBWOPf0jhiyo
SlqxniwPi2TdXT0yjwjrlya+/gYV4MP0FEomDIk9GgWkQaKJhUcwrfjoCdrgqqOj
9fU3Ye4elmlOebybrcZGaS1I99ZriCCwfzue5Y+VSEiSsf14ebckIafWElSoFDIl
iAuR52cLd1+kE86AE9X+99mHT8L3XDO6FLUIXzLemyZUmEAdXwO1N4+swZGDLl3r
RboR9EpJzjFcxg/yL2cj8qFZENCyuWRq1L6Hfj/8OHr28vMFLht3qBCwkGgdE46E
qtunWftmOmKbYs9x1rDGExuK3GrHZKdPHw9o6WChfedHn1QETd0Qkw/3klhv8g5G
KM26/ZKMBp6uEduuCj1HG0yHpLWT+MVXwn+5OPvw4bZ5RDDUmE20V4dWjpSZ12To
34dZlg8HPoarzKcELPlXe/NXtx8VzFXJUPM6lFb5IB1DuXiCJO7IB2KKi2wcfUKq
W8TywZQeobgYfUSt3PeU9Rt8Y/W/kLVid4u0i8g19qYp8R/h+no2W+nsigf8GQSF
sMTaj3FK3fGNftG0xHjNsDZETglBkZThmDlcpRe5rP5Qfe3RHOtSd8hqGrBGSLQg
7H/yP+Ky2lbCCJnuBGFVu1SqUF7Ut4ahqZgzGRKW+mYbn3bq41Bq373Enpg7sj7l
q9wQK/TMXcgJBkp5/vFP9jyOOHbKkqeOBvu9pTy8zqAd6QCXmaUxIajpN6lcTJq6
WT24bbBbq/0k0icyd+2FoUxcZrwxNmaZfSEfkD07LLw1eLgOqF8LNhOezresVjeV
HpFXRPZYStTBM5vY7ZaWlIx2akjepyzY5MLeMmTXh7RibhoinOl3fjtAODXXPyTY
Wpj1BwQm2cW4J5KtYZZtfDPmAb4vReKpPOERA2cuAe621N9PiuG6HLrSCAh/qDy8
ES1Sn0s/elt49LACsjus78x/ae+44ZiP6rWpKOKr4rSv6OM+MNcNrAo5bE4yREr9
kb8KvJ09D8fPkNMmpMRr2/+1x8EMel/gIXYfEf0nwUCemgLLyOhftaDWEuBlMEd+
fYHBx8h1fhjTymP4HuLrmTc4391HMDVChDm9i1kUV+8pnk4e5R03aeTp6MsPH1rR
0UAUT0Xa7HDpHSaahK19lKblgrr7+0DoEVFH3D27vn6GZQYPHr/krl+0KdUylniO
O3pfGUthA+vHggtbKqY1DYUJYHHYuskpdBDRuOz7miBYlswCHD5DvNxWP1j/CVC2
jMMl8/asfsFmK/5Z3cddgwJJUAcml77XZtjLBrfWHRbUM31IVomT7lhVFOOxQSAN
8pxU9YFXGh+zPWZpqAOwEFMfz/Z6tTae2AeCfqzKQA4Y6edjAHVTGeESQzNy0JHX
dA7iczkRHQzo8/PlB5Hrj2eOcyn1cH6OGxfFpoebVYNWoJf1rq5WmuwF6ocS01dj
kEQCciFdpKHAsQcnrgdibRLdnI6lL2/uOP/864d+uzN+hz9b0bZbSLLJawbAUO/u
zrBkt7y3F6cj7I8iScqanWnG3Lu0ZWVU7h9r7lsDSdCEhpADLL6J9+N/TgilRqMS
Od4HBC+sVKQ5VKtYydzom3Iww+9gRiMiB8HDd30QjK/Saif5LaX8fhoOYQHSTOmT
SpI7rd1ds5Y4mYwGV+7WHF8iboV5Hj2eHVNTACCI6NEYSrZIwWKHo3BKxjDaUJTT
QH5N/ZYP9XMvuKyRYNy9Y2hBu5tsYICe/CFz99zwbw4+QoPtg6p1Xy1J2M2ToVBt
x2vB31vNNY8DbmsXNdFcrc9+rAkYf255E9zO+NITazWk7IL4OnPxuNzixTQ2sZlp
ewxN/3ITr7oQedxf6tRbfHW3N51jtQGug4GUOjLvgUxbJ2kHdJgRuLFnVxPkCrNc
6owtSrRnYBYlTwHJJJ3QJdwkdX3vIIq++6K/7Wryp/5iP6xYE2pju/bZhJ44AFSc
jZvuPz0EoRu8P+rEQRmvJ2WGKHcAsSPSOSySYLpAavAeUzi6pXlfEbnumvCEKgqt
MimPWIrqIVh/367oL/ExYtRKYyWVCyvQPu8AiW3aIA/ubY7kFYyVINgnOz9vOJzr
TcaCokkp/xf2SoLPAPWp99C3JbWuqd9kTY+sNaddPmovai/LesfXV5wfZfRItSL9
uIeA9EAkT23hzCi3pcC+6wQ6NZz9CQ4/kGCftUKhF33Izxs2agyW0lbpateGUNIz
7E40/S1DWTCNTq5qoe6MirEgFbeMQApOuJz1GKs2N6Zb3WbM2iwjArzN391IL9tU
H8OF7lcU6q4/kRIsVbMMn2YCGdpDfiMZN7n84DvhIUUXomW+EKZquaX4eXSRwOsp
kfc+Pnhz3Ew98/+3BENsWKxwDakpte0wkFHoQvbyVtnlr4oQO3JN/90H8CWLNkUV
shiksf+RU4KZaK/VkZhvTsbAkN5BuBK28QPVdouHJ7jcTXOpTvluDOC4vjo9IIDo
bgs8GBdwKmlCtJpzMT479J3Am8O9/rMSKQgWe7/gVVUbNba8VZX31UBemM5OkS2k
PiLnACQCp9woEl6xLIY7Pzrw8VWdD4e6Q+/Upf+ZYD5GW3JcNyveKrcFi1i9iNJO
kNRCVH2Ih7SAjz/uo+0JJJHBHYovUeLI3Uii0lZtP1OJDjau5WKtIpiQqvBg2Sdn
j9iXdemedYLeaMDSbVUdBZ9cBq2zu9BpJPhutw6v7V46WGWuDh3NUBBKdHLsCOPi
243+Csw7dYWCeCrXPSzRMBag+4CwGWRdtyizcI4DBZxqnAXZkmVuEtBwMGmG3Bf7
I/Yy9T8//EFjHcmg4ToVRq1KGVfLIrmHhFWLG4yUIYnUXaoPTeW7kThACDJwkVrM
fTAiyDZQZYprdRD6icRQM4aJpxz3E9AttCiAfjX/NsD9Zql4m8a1utEPva9J7wGU
XWjxmh4NfRUoMyAPfsj4hSGbtOdaujJEt+IBRNauYrzv2jcXYvc9a9AE3dUZC+hf
ebQVP+ersOU+/h2YpKsJAUzD4Udy7Z1DOaBe/+LPXEDyQCux0pN6HTfH8uH6X4GW
fVvb+BEh0WKHNibfCJAakaTyolcY5+DY9xQctR3wkZIOStWn51v+5K0wps3ZrNk4
7A9wSBKMZjPzCLtAmopVTWmSeTWHUwe8RKLy0Ej/URgApmE/tFOSIcb13EqdUkle
jaSG6odsI8bfJVJupKbVLW8JtzB2zwKaxyKke5N/INA/yMti1Ua+Sh0Sky/w0NGy
B++lqIBvQ4fYzbRSaRG0R9ZDMxtHCJraIgpx4cVDA83KitclGBEusAlC9DF3Dsp3
6JDDBDpTnkh0q7Qui65qrlud/V0bM7eliGJPhhnvcEA84WBj3Zn8Ymn9p4LZcmu2
3sqhG/0Yx5+/ibYGkGqZKMu9Ofra8dNoOflJRUv+gp8qpGQTf2bGOx0Y0k8g9k+S
nGMhcymeWr8JMWWsHMS/TeWhZa+Z0NvJdgaODd/TTdkVskrlDFw1YsDYy4xeBs/C
pw1mhArMm0LGjjUm9YkZdHrpnPyxY+OFONZTecabc9eZjvzxseFrsuU2R6eqH1oN
TR/9OpXH81J+ttYTt+SY/XY146+T2nx8KEUlyju7a0CQZDkl2e4JuQc0LDbg8+dw
WNUGpQC5kJ1hPNY161xG5xmbUlz6ZYnID0KOKYNintQIDzJKK0n9Pl7hf3AM0QZW
PBhRa5gixOSG+ZqsHxceaR+imfNUl6HCqVoSmbMW2rfEkutUrhJT922t9rotTmNn
ar1UUwzv8SxEvd+5ytw3rgCQeoWL+H3D+SF12+cmU6BQfWjaZdGwDU6y8o8+nwQF
ybmJXCcVolvCInYFQLp6/RXBGLtKc7hH7E16frvq/v790frLFt3ne1ysEAwIw4ag
aCTGQlK1JLKPpv5YX7IXk1/6npGqc6RQKpRCNcEjLSOVyvGvcTZEGhhF/B/cNkMW
ddeiKXgW0+YRH+KnFuG2N2D4ZotWmZsR2lV7gd22rrdSls7LT8B9bPuqOHPb6Yh7
uJrphxMuIayecu7X9UWQb6DGCLET2VuVISmWOBnU3HUSFgAZbrJ0tNmeTqKiWoPK
UxFtSRc4F35Yu9XB6h6nqKstoAyFke4dgfiKyuMy3wd+J54xhb+/gTkJUkTmbHV4
kQcVKOahwWolaLcyoV7P7V3ngAcgs5b/o5UPaK5GGZeirjtGDDBJaWQ2tzPCotwq
mJBmdre90cdZrQXhp5tvXr1larVwnjnawKUcj/Cca5rE9zHBymJVmT+3mfbB7VlU
LmBZOf6hkkykSbcdwweBZYPVrZnURvOzdqkz5GsJ/pjXlOANHBsUt88OLaf26YW6
2C4qytCUNBpc1ktdftgBRK9JZBVovAX+9b6l6/AyGvLc99CQ6hhRDTuCQ28x9IYv
nc9/IDYVpU5hIeXrZW1Ydpm2P4XOoEOqqNV3ois/mDEGofu6nTpFCNyCNqQ3nnL7
6UjdecGf0Sjw+t/g207InRJToiCPM8lqbCn5PFAsPPx0G1B+AqGVF8TFwuA1odyE
lVsXClGnvMo4m7jvakZ+vVe2o6YoSwTs640GZzIOAQWslwB8qENutWv48ju6ifNN
koWHbzT6XGlmKvQkPMPKSvYvcM29rBYOaEibjhXvFWImQ43iTtpxrk0s7qmVhCZe
WbCuipLl8pgGcqtZcGCE69o68q8X6gift8VIqljEwYHK7Evu03fiYlzNcQ0V+c2o
VhuUOMF7B05ebOZB03DEI3+ZNY1aUJBr1CfSbXtyz+NYx0l9peFZMRUxj5hwFSCe
VGbN75lPmEjVITYESMcN05KUmZNHjW6K9OeVPW/xJyPSvF0BeAsWiMYE/0D91fUN
n56mCwNCxTPJfQnAGXgykMEKc1gkIWyCaQiUmU0a4IQrvFTwu72V438Couu+kCnV
XMC9CvVAmDa/BrtwNNrapN2SoA3VHykB78+MODr+wfREZZXdgOmFoYsBcU+0xyp7
LFxClD82KlB55n6rGlBlnKF8nnGuSfdO5/kCKfI5PEEcYXZ1g05eharTpwnbYGRy
n5S+7rKTu1MEELEEdX2Hd/h+UB2ec4LQaXoU2FX2IFf+dxVgO3B0eD6G22TCR0YT
WlQ3RWuJogO4M1eD0MS+5XWiTQN7SZIY8jzia9D6mp+IS6ArGauALS9df+9kKtGL
Wytm2kyKHbrWMC6VVW8rIPl1S0jtOZ/tmBJN4lkQvlZiAp0TjqgLrt3DujtJLUDg
y6B3bexF6naMEv+ix2nvgO3sQSsjS/4B+05lIsaR8Z+/GsfUVFFvmFdrqvpCU/u4
I+ICTfvs9pIMBrrwZ+QRixGW4Z9JsVzjR4FhuMfLd2dDZO6oSF6YvbcsWUDzr/ux
HLwnMSJ0gKEab8g6Ni2MJEnXLLv7LMZ1aFYsBCSMo6z0pIpByRMUzjQCRZDvzGAf
mXrsnTpD5vxcghnphu2cZF8aVeDzbVzTz7nnhheDRecZqy6QVpQNX6vxcvV7mBfS
BVjiS9VuUNID/H5PeXjPChQtYyDxF27eG+yi/fcJ90zAaC1sXTpcWZ9Qip2yr4j8
f437fjrnm6fEQ2Cdkx4vO6ClhcZBTR27il2eZHAlk+VXKDrxiKoGBjZ8rq8hC7oX
lQ946ZqNE30GlN/PPweXvCyHzJXNWeeF8eglzJELdMP7NXaTWuWwC8X5Wpc31sl2
oivSXgd9STa/VdvaaFhSWmJzH5jPuH4jcrF3o4SE62ziILIMfcdvBWR4fSOIpuhV
R5nyAiyLp1VrJOLkNfZbv9obQrxUH3a53BPCuXlJC0sZyj+pphkvOGtCblS1aXVw
BMG1raKjSnOTThWAe7TiYH/zX6UpnPu/0LS3UcKT0Zx3yI3X2Xz6xAgAXhEPR1ua
L5X+qVYFqmqEoK6Qsf+k4FEMP0xy8pWhKaJQO6lvS9T3DvXxbX0Er1qI4C5UuGGP
PuMeuut4fzbtdfjRmyQNGGAHx6fVXWdP9I1EmJ0PGxPT1o/gY/aL1Pp8+rDxCNA9
pLav7BTsOatOz8xK3E99cyEhOPiqhhjILQ7h7NjXVAUx9I/fT1ysoPkXXHZ4CmhB
NVPhtQHpLjqVNJSN8IEtqVV0OSS5P4ToFDGqAjMq9CbYf2DjV9Kwas7lQ4BEs4f9
laDwEX2lXg2OaHj/o/OZkS+AU86vxqA7rKvIKunD7eC1uRQUJxucpm9EO0XBxmVQ
QQjAvzkyi21NkVJGG8U1iWk/3LD5HIsD/scwL9mekbVFKLoRc+gGmY10piCtqTOz
KvbFBKj30Vj6gb9rTRgYogeWnyM3/FhlToKWS8vG18l3MWW7osBszDheXY6JRLHP
zyEC4m5NjBLESbPa+2uHLLfsoWR8OfLE6hjSQUVa2BTHkOHMEK4OOaquxDLZcvCx
Y4B0JlQB7AYSt/tPGrKLBYbFwafJlmM9Vd6HGkZcqHSS2Is4AdE6wO/6NnCt4PDd
YRHlz94DPBQ7ebQrPTdWQ+vb/caGcWgvx+xrC1fj5WIKeX3YM8SFKDNpwdttdyay
hLXg/XCY/lGqx/SD9OKFSEKX4Hvrl7YPXDc2GzoSWLrqS1gN46qwBSiZycYeBCdz
t1feGmJpa1IA8qbWFOxjI2Vvv7w/4pQYFzgJqq9XD6htS5e0z8uFyoBTsBrATZ/W
2EUFiaOuK9HCFbQ0jIVHlSvLyV7eSHNEnKRd+4GK3r+DZLH8hDuwDruRTF11T+Ry
iPPLPBwtikduDdQ/60P/7KAOhLR94aikF3h+fN124S/EtzL/oteFB7iLhw5aic/k
rB8fXM9702lwX8876BHiLXBATn8Ag0KG2Fl0eZc+Rj2vbLGYd5jNdVWJGO9gowVv
Z/StJdfvuFkcdaz3lgsbJ1Ic7EsBZVFbzu6OxJ5Os5mgTp0QCFw7lllz6aO7cJIh
LdJokXsdZuvpEGD2I0DaTbgYPu1qXf024cRqMhVV6GN6Wp337/b8KdkvQiWChVVT
gTkIUPnZrVK4DCqthThqb1Cl3SVUHKSEXCQTgsttt3KkL5kvb97ftB16siR/ae2g
xwY/ecvTgBQhyYtN8VKQ9DYIYbnMiBcGpwiUgme2AZkxiy7iEl+4Oum8BddbvrZi
So37NJZIFIFhkDbJDES7xFlWcEYSfnTQ+W/B65QEg4fDrMhs/7bez4LJlWLzjUD+
IzAUdXw5quOWu6YuNKp2XcFkJm5dnpeOYsrBtIICeQlb5Vl8BYLFDytRWgpGRiqU
CA1VzNK2z5usfzH9G+mW+kd1qtvyzdKmjl9IUrTj3Tdtttm4dsF62WMPDCd04M8y
xssQtyOHzx3WwbBz4N7IaaT2HvsxH2neBTp6r6by+JASFyfkfpJwxsFkJauVodbw
edbHLACHibBg2da/PPARM8fYI6Cg/RshY/WD0dX/GxTOjiQMXe68Nu+GB7cqzMMN
nlpKiR7QwfUE78tniQ9GjBNi4SQ/OpaFX0UL+yHfSVmSsVk9AWiQ9c+JuzlnhiEX
JDeaa/R9QjlTwcgHVkFVo0U6x2gx2Rq+kIgnoExuf76rZ5uRqh+AoqMMKiiUdO1Z
E8vt2vuBE3YEmX5EghEr+8Sfsb915gQ3BDkaxZXjSbmGqAVi0H76v+9jXTGaGFlW
Bsgmc1UeJShpvBqe3FkIo4Jt+XSRzze4frkGpc6acGJ7KAHSeZjCEGj9IOTE20ov
6OL8Mpg9izZ/6+s41g4kcrJ05QTiu9L1LlSKJ1owb4y3XzXXIvVZyV/2/GswtfgP
vxZgOTIjHYIisbc5WaZhnmJSo66Y0Ew1I5MDFPH75SvLHEYiBNuQmxQeFJm0a4d5
JHEoCMPiwXul/Uq8YrxQ456MlDHQHjXXYl9VFQPQKzXfBdPJpURoVnjhWolhUbcn
ChlCTSUeffMKl4vjSgAnzboZE5GERrcUPus7TkTh9Q16NMDFfUvpzCBrJ6cpqNn/
/PnOiL5QGFKctC7cbnudZvAcuEmNuwOYnkC3wskZi3vKWu8CMftSt1cy1nTyq+2R
qU6dZBKnG/W/KVe/VO/RuOXbnVT3Ub4SC/da8mmF6gWdNBh721pOtEwSL8/JxMUt
msN8q15NtA8h/+H+2qd9ffmGA/5plLs0TA4qg/4DFsUOc+0SnKKBHqPFR4NUs3hR
3bTzNguME3z72vt+7MtjcU14NyWT4J5oowbhFnOzStbXVmfoU/HkYOrCVRYb0R2B
vT9cezmIS0r1KKg02xo3QNiSIQ7ejYRTDoJiNTtil4rJlwl7kDZ6eWOOzxJI8X47
8kbfExDiUgaPjGTCmVmKG960F5dS5zksHQneF0CyYvwjvGMV0KCd2yojKq5fqtZk
XRx6vjus2skLCOnwhmm4cv90KrlPppEgzyOBIj5tWo1Qyn6MPDf7TsnLPSROx3MU
1BNQad9PKOYrC3XVHIU0mjpKa1ukpE6eryopsukuP0/flRee/yxzNKzExzi+XbVk
7/ZlnwhU2ww/PyINnaKSENRJkDgwfEg79GisgAWGKlvcwkI0abA7mgoFUyjX72iM
MWJy1etfDGQ23S29UcYHGMy+KYpGfitjv5B8Y8aFl6Pm2xEL73NTQX0YwXes09Rg
1laYvG95G6z0q5rRw6bxkR5W2xZOrixSm/ANPIMZfcgYwZCu42fqbZFG0glKsKe/
5VAaNyoiK1HZTm3AqQeJvKsMVdNaClEyRorpMiGRc204hArKCDDz+g1lBqk+d+6M
3g+Txt/QXw4CZf7oqutl2l6wuEKK1rftoBi+UdhAmfhblVXgvXDH979NZS/xzWn6
TiQAi2hZpFeFwAUMvjp5q5aeZI7KCXTP9uNYsmI9NgR8hTbHyh7jmmBQiZGzQg3+
3jed08RXkH8p9YvCXb1cjCmeWQYF6am/3waALR8QDkXHkjDTC6ZO1lm3m6bizdJI
PCbuBVr8T7/IaSHBx7b8JrnPWr1tJ+MqKMkmzfVv1BKBWAijeMSqG0sHLdFi51LG
lstc1Cf/5bV2rQ9hsvuM1lAw+zjUat5MCfhP9DtXizIRe7zFkDvPC3mVDaeJvlIX
HgHUl6CgyZl/LnmDTsRqACpaayQW4Eqp6+xPsqVhMYN11f7n5E07w5WY5OcuS24O
OZ9QYsr2crZIsg+/YjC1iB1nXY/AnaJt1atG1wv31LRqY362YOYvFMVZRV/Fc8VY
/Sucg11j2HozdEMT9AFJ0VX9PNO2mQLHE4jlyOO9QK8VNPR30MWbgBGb8PWXEkk0
8hrXevDvricDi6eHjydPTpLXSOZi5f7csyQuYBCUkMvxluzvRCRjvknvPm7DTbRZ
TPAHHize7y+9rQlno+JQELeD8lQTh8/aHjcAgBNPFcRxuZjIgVVHdb3C2XCsF8pj
9gFR2IGQz4H1Ec8+gFtG6/FrHnuchNGX+9rlQl+UpF2MNJEGfcoBGQr0adD9s8sP
gQnC8DPLkA7Y6VO6Yq+wGJsSW2w1V3KQM6I7r2Rc0yNoezgR7RwdeYfhy0YfDJxc
IoqXQJjJaRfsjM7966GXkqz+EgTZgo2aE1kYQlIKQm647K8hSOEjiOPVORVGVGRt
5W0JWtJnVpKlqAguvfq3GJhiFksETRU7PHKkWJEl0kOcuvKLEPWHSn3TC/xljAUh
go5GxcELz9dyHr2+/XXMhpozPnDhQPw5KBuPLsa+I3RsVjW4bDcKO9IxjbHopHeY
tarOgNFjEVUmbNRcnE2SJUJ8vHMjge2M7DurVI7/7vjC0mPPoOnKFwVQdYhu9fhi
WV0A2kU2UV8KZba7AEwDMA5dHRBMF7HBfrTZqVqd0hd8WPErhYeKoF3CUDRre/i5
eaikTMAUCmyITGf6F1ZM6ChAG9SHxCIW1hJsKJ0/J8xawLkfUexE7u+wAM3bGLSC
q3UcT9G/tb6B+7V78q89ox1xqYPnTKx37zqrNaAkhnGJdqo74JIDf2yqE6VX/AGS
bv0xp1kTD9AGaoSI+mYYJub3PbY6lk+gt9jjm1UvPH0GDil3uTCA2s5PcF6g4LrV
efFhSxzmM7XawgGTW0YdXZX+h27RSeKJr3mUTdaoYjSsZb00uWC9hHPRDKKdVNNJ
rVvhG+E2lWPeaJ37+WlXkZwLnpd1R5+7Bjy3sliWvP1NdmgmmQS3EdJm6fGfbEYU
F2OzAMoH0tm8Sg244PWfJbx5jRtw0M+FW3lKCoJSPBB9VwqzcYuwEwVhwfOsp72Y
IHTJvph1KHeNpUadRgRq05zMIu+LKQGWvIZYShODbWrZTh/9OAAHGAYcoDsJfEGB
GfYAEwsSZi2prdASGdV1GVo7uGLoD2vmTF6shMt01IgAJPUgTHFXxpSg94low8ac
VhBwP+F/xKx64c4nP8felnxRscWO+krPSGzB8KcmWyReehhNJ9qScpIFycpfi8rn
A0qz8YrpcFxiERzWzzxKf+horGjpRLDno59YyGuA72nLe9FhpGiU/feyHs7Jh3Py
l4rTlL8Y+5qMs4dg9g8lDl7FoScL+I6EUdXtXKPQLlioMP3z14614WF5PZRm0Sg6
rR0WkDtsFtKla8sdoCKOWLeORUpdLbgQ0uA/bsk+dSnGCRNz6GVQLBgCdEOu8g7D
6UmsPyl/13d1pkI6ZOuoueYJC10I4osI0YdTA7UC4rPKWeTkYOYc2OKelg6UWGx3
FBroB2WbEwZo+miQTbApvnUFY8hYRDvrAyzZoNMKZnQWnTEvKlUioRN0ggqSgmvx
omOBuGM0j7lj4ngyKBfiZUVGLJVN21P7Ptq4iRt+5Z8Tetbbcurns66pIjK3b+ty
/UXZ/JSMOSdDpHk2IWdQy6ez4ehVrKpBLRT6gnhuTAoYFr8+S8Mcx94nRtfaK+Gn
ked83yWU+Zbd9yGq4ftPdhA+yV+QJQu5bJV+51s2rSsBoPcf1G8NY2Y6+cj9L2Nw
BZbFyW7tGuDkcUvENKwyUAP/kYNqEi5kQliEj/ehFLi/51mcR+L0I/01SL5VbyQn
PnzPJ8rW/FlyzOtTtUgm3BHeRbDx1ITxBfMVR9bn2WykyX9Bprw4Q+C2Au970K2/
ita/2gJTExG7VFLr4Ia0o9oFhmRzSxS8SbWGrPjayxp+JU9cw5roI/MPrdrp8Moq
0om9PkZVMIgA08dUL8pQDltE9VK8iPCl3OtvSkFOYm7p+ttL+Ocohn3mqNT5zRr9
lf+HIzuHeKdBvlMZzyS3G+4qFVRhCnD930riZtnnxDjm1ikKdyqx+WUF4Emfv0tK
4kNdZSJcS3TVapldmiwwlZw+eWbUlXan91d5hW/BTtkTEIDGRs95rx9nTErMxt5n
t6ZCuvDKBXr6lHUMOmOzCpxwEmXLvLpDPulp09Ysk3qzJkjwVm++19QOyvoOsGw4
BUcq5alYYbTGTs+shaZvo2gE++KCyJo7fydYCFYjY+gohFbv4KXVtvWuGQv+HtW+
/WKs8rPC7riJY11REWyhm10lFGR1aYmdi3Hn4FIkZcAEO66MSthGDdmSN4KZijaE
WABAVEisDnR688a9TxYDFGQs013aa+1bYLB3VZPL+Q1govSmjpZXXuNg4/o4ONHR
rXDjBPO4pX4PfbtUbcOZEpLSbB8yF7J4E9bTe7qZsnH+GBc5Q3Rq5/75UcSK/2LU
M+1NWsA7jkW4/PeIjMJCkd4hpPIkEbnJrL3htBlI579XS8CkupON6w+uvpEDEmQh
s/68RfPe7twMScCqXV+q+rlio1ZQAwHolDXslms8d2/GxN+nwCL/yr2Pla0dY7xH
59TtEHLtzGCgbZdoUHILMJQcmEPmA6Cc9nm3f+Dr7M4vvuRPG+16Gb1Nlw+tckoU
4m1c+iyx5LB1OtMuBjemhrBZVsaRFpIDpMlnJBns12+UeCvSy+uGsPpeQnj7vP0d
CdwPpXcil+6AxNCfa/AVGsqIv3duujl3H6UDHhPwKcKHW7yYfRVsWEmH7INR7eGs
EVV7FP88NWi3XaMrRijaHKJ6r8HRXwB0U8eagtOtEupFWSnnkLtODNEl8O7ckzbG
7FH7vsOvKJ+6zXNxvkTMIkAjMXEr3EQBVFFVEcWqX4M248nSYOW095u+BXo2SwVa
Jn+sp4KYJfd4tvFlb+GlJieVZxLn1Gd79gpy+5HblOobrTXEBm1obxlF0xoWOKNg
TKnY++w5YmwFZEZ3QZbj+Xbqz7CWybHlCby8nmzj/L68UbkXbgDqFTnoVuTNopuN
t/CKnPU4zOCw42WNPjzg+xg/UygttvN1T6bDSFM0EUs+2ML/Bva4aauqR7UIscIa
c8rPfNFseJ2xTi70xXOYdSJw3A79I/dblTKQtQ0WL4lhQHNoBDd7FK1FBl6494E2
xsEFj2HzedC81NqjyK62IC1ZWrAGvMG+z9sTIc7AECUujGwnnqRNFY9mkajd3pCH
bTGVT/Ji4ERJiebthkwrPEg8/641lJ0voVsviE+kmwbs4dGytb3bqrVjxffNIZE7
b+YhMABLbWlQWnkoMVsg1prSYvS6nYKMdCKP+0ygN4hX2atwnxz5ZsTdVIot6Scc
D+FPhu9eiRCnmN7LCns0mEMdCkYmKF4JBSKfoKuslOjJo50xzLhISB403vfykzqW
8VJeVm6YEn5e9dhAMWvdQRyeQFmFXFShvoTI/EmOMlMr9Z7TwucpBF64ufenx/oC
Vv5KqxQq9pxjdbOq2E1nFXVs/g1fi6T6I9OFbDyyjXMJJvVVMVrwCkfIO0MEBve4
Q9MQa+WNjSzQ71qSSWO2eFctANp1jmtJemejga8BhV7S6cRPuTKaeqFgXswQ7tv/
FPmTeNJ43cie3g3aeP4hOvYEua0ezYuqk9HBvDXsIaHQQrm1fcxjsJ88dCt70926
tjhaDK5lkia47B5wpuIplvFSVj6aPBuL6up3iymQminVLnWfyJ21mDO92netjoTC
wmO7HZudVoGE+xIh+cn68CxX2HfMNyfazt+tBAPDBMB9Z+9l1Q4Tua8wk6hFqn2R
iG8a3ozheBuWBN9gTxM7UTTrMQ3hzG7zd7JwK+BBOfsG2hDrc4ZyqbM/JxHHC4b3
e3FmKighNvsYmpHX4Ms5xM4kNs5d+IRk6s9sd3UDC/3BBQ0YZkFk8vSuE/kYeznt
4fuOZVA0VTLDQdn7X7gi/L4XSuU5Rw54wqGqYHsN76JFf419xeKfI6BFhoOCos3U
bRZtPbFgDktYKGY9Cx5Wxk8QzyP4EYLdF7NmQ2xSNRe5wchuMLUzfTme3gOsNM6I
GWxCB8d7slWUSn1MxA3zm7fLD2ODZsi3tdoDFcniCmD0aqOOFiQfblhHPlqcLi60
hs+Y1LR1O8DDtqKv2HwtFa/LmuvVNrrOxzSJDPe6O8sgHidM1o4oYXthUnckB6WF
XHpFR3vN4WM6THhZBYG1EccuipI3rZ1Wc/IP0hF3IEobkNZ4cGWvWe3f7VTx6ef+
NZwWMUviDSEjxXmt7hflL8on4OnzJTzuUU2Lgh6QOnrKr/cxlq0+PTSGuzGDvIG2
QJf6176U7eVozha8GPMCW9tZBxBQDyA7nnRVxINaOdjKwnXjGl1685ougWdTcU8Y
B6k++3aMg90d9qgLA2eztzSgI2vdNj3sh90fRt2vcV+4K0Q5uRAkSmNNqtHqQTHy
0V1GDHXTpavKJcBWivhOOk/zOxb976rAP0/lH3u6WGlWTst8pdsnL4YvP0B4p2WQ
6XkmauUjCLg6LNphvBWf32PbLxxZNQiU2VorvBwdWzy0NvLZQeoBrSJ6kFENhg4F
KED9fXZJcuKlR/D5kanpqdqrXnicViDHlXPeLZNEZFPlxeViktyKG6m2PlPhGPNX
t5Gq100nT69yo2Qi+0A6QTkz/MaZEZNPo4qiBnS4GY1bqbN8f+w6CS/SX3tFfcmt
ouFF+wl2441GuyJ/k3H/HS/D5N/S/hQG/+EPC7GB1vTTJIVhWPKsWU1VnvtKTm9j
DRnKKXNfgyVhTjsUgu206Bk1K456DgD5BvIsf9ctp2AlInC4IoMQehQ9AYLjyOZo
TWhdeSp+6U2u6BZl2XVXI+eiL6o1NGEl9uvrM2Aut0JZBPtciviP+lg7fb2Lf/JX
whOlIjVmjOdQF5/zfavDumoZuMF6kbLls7mkaTlsA+BFnfLkrB4TTt2Ikgo2aki8
WkirKmh1vQqNnHLnWKRBFSLZ8jrfCI5YVFlm5mm+vPjYJ/yh1OddONr1jccczuzR
XSX6Q9JZZQ7/uVPPx0lRMHxhawbgEg4XUejK1nch8c2qim3tC0Ilw4apGhEO7C+u
oT7lY/D3HC/lJHKzUXyXTwhHdpOpN4sXvsbuD7ER5gQW2T92gnS6r/SGdOc3+Oa2
XqcGBuLqoi482T9DQ6+2EWQ6Ml1HYxWoZfG5NI5aw8GO7PJ66ihtbMFsMDyllhVx
CFOZJD71zgqFIHb+Yw95+mtSlTTw4O4HMngSIgI+nXhYAF5GvLOfAXvoMfQRsp6E
Bb9TzcT/+OfeuQBKt2mChg3npLDxhcgoUX0TFWwX/7UyZJTPBO15t3DVL1Bxxb5R
G++osi3RQiXIKXSWsinQBExxXZTQVcK1GqcI3CgTgLrZVNAsWy9WcX5nCa61UzB4
GVfILQEKUj9fAdWMJlwwIoowYT3ZxXJlx3OoRahvdjZSd8jtJtfWsybQIVk+NeFh
kPrt964nd9IDI2pWul5+mqwexRkMLRubH+PCJQkg/gatalBhpZWW15V0BhRuyTy+
6oW4s+9jaWFEGSHAKSQwhv/Chm/W9Cd+HYGXr3EJfCG4pwL/yPXW7NYRKRfsDoiC
z1V7eLKuLdcIHSx4TWFwBq59n510oQ3/8BcdZSAIcjX7aIXtRBDlBlv/pgoc+/fB
7dzCOpP0tAJdIKrkfVbwXJGyLrDfRnVDx/JBKb6IA30ldE/xv2DffAYnxlVvMwoS
jYysX3QlDfF41k5wKys5G2LPEsZwwv5Mzj07pynIKXG1vqypPYEa/i4rNxtthXKd
ERUNLtePUB3l4PZ03ygVu9t6ZaNeZM2anA1W6+ek07rINrVy2sLbk0EEk7JjFleF
CFtM5xGJSCqCcquh0r4jCoIRsAJ7TEMn2vLOcIw3zNawsb04AAoCVVPfr2g2gZHw
tRzeaG8IOsIHJ60zgcWKaWAkiKR7av6easVM2GQB4paj0J5AUSa9SSa1r7iYea8t
tN4ysy+EGF9GtsCBmYUNfDPWvW3vvlLMvmJqbNI8+HVmWH4JXGeNoxV8Gg5SuJiG
SuVTniredcxTGjN5/HRs6vT9n87qRsiJjrc1vRenCdL0M1d89070BthoosigplU9
Ttnvox5keaumtgJFb8fHJikTHlkS2llfF7hjI4O1Ro2Tnuk4KAhh5A76wf3ijuSa
rn62V0Aj4R3YgzhEnpTt9iKDmmiS/nTWbY/X8SKjpJ3nBwRFI7pJJNBQB2nDsfEp
XGqfxlUpOEmPNWliXrfdTCnE7j0rtatwLzLLg6XQ//T76YSuDokffLtVZwQ4Q0Er
Za3FuKLT8pauhb3fEtHhrY6d5n9Yf9rrZ4XWhxRZaiN660rSahsWW59FcT8r/wgx
4j96nFbieg3MjjqCCs1R1T30Ohos3Ep3RVgyae9kHUFiy41WcT5bDVDe2L8LSenm
J/zJ9maVE7wtR0a1wsYDKruQmi+yieFDj9KllAMiaFmWYcLNvB568knR61UlCe8X
rTls+louy4HMtf621v13wT/tvvQDcoYcwMj2F0hMEjq8nT55N0gb6xmRrpGk3q6i
ai2FtTmpCwRCun/1bqBptFqgLN0wJV4+sjz5da8pW37Exs+NXden3GfRBc/SBE7i
AcmQIMC45JSI7VQgEForcbd5zgUHAuM3PlY4VaShJHId08QGd0DWEDY+D1rhgFXq
NuCDol3TobrkrMBXeqXbBY8bEXFFPmq+skPmNonoEpBPtxOqxAlnaK55KKeX5M2y
DCkoER0wDhGOT1TQ37DQUy06d6aUJ263Z0zFHHKytdUdq7Kat4Q7Py6pVo8d1A5J
5X3T0S3t9DjHLYj2LQlq6WGbJ/9WXSv1uD8HoYMZ3vXrM0wCnjT9SXBzHpzxQlzC
3OnRIkB0ic01ePwgBdIvJ1HOOwbGVviOXT162GtSAyqw2uYIh+Pr0Q4KABtTHNuX
xEgm0EfSc3fatbRsYrZ1+gArB2TX2WcTvFdQtm75DGY9DwsDV5aGBHPQGnx8v0qt
ezLU4cSuGE6fRTnnFqNm94NxiKn9g40R8quthlawb8D+MriNreU4YaqKZBJUetMz
kPNUSl+BKDwekE5dV+b4QqnoAgD6wXulvu1/krYO8vk3g3MiOrsL+EKtMgsy99Kp
JA5Wlgwm2qId5x7RSc+bML9HbIPDo2Fa86B5OcTceXtI7juWywu7tBctsbWZTpFP
IKiULBkUCcwStnGdrxg2h2xInyYznsYjBxZqWi7YYOyNAlyCMw5zdJtgCny6+lrh
Iwcw8dDJFcgpYprZNZyBs2+ed5Egs2AuB2HA60HDrE98ECsK+7qJAISIJPl1lZ4Z
PeCoOpIocZzwpov5DWNLc59d9GQsg8ElsC+qqBrCSst8Qw8/FRidKBxRHq/rltK/
s9XEGgj7GW1UiI+AmB0IeLu/9Ud8/R0kxXcx4X8rh94iZvWoZcwv2mj0Nc7UucvM
etjF8ixiVIGpQ6h/F+DnDwiydZCZEtFTSIm40r8nrgbStvfs/R+LLk4A3bSfadv8
HN9TKxGH+5dcb0cW+WRp/F6KXIlwUQmYL3pSQLURtwJbrHAin0DulLR1KBnm4RFz
tzbJMBAVZ5RuWSTprcyxDSUYLC2KPz5bTOg188yVbkZw93Yrhw4o4q/no/Gkza0E
ErctR4mPf9apagN3CAWviF56TD1eBQSRAyemvaTIP7X2bw0k0mrLVyNTEzKFd7OU
tRNf6ulshkl+D7x3VTANON44n2IPPkYgXSnJCSkIes7TdEtcXORnxyssQaz5ZuEL
QqsXKWv8rygKsKzg3ZMGiQ4aKN5efbEGzed19Bjn9cyiiH8kwE3JPM9OIl9PHvw7
3HxxcN6l9jF8v1x3MeJqwat+AN3MbJ4nmylpwUpeKdd5RXvxQDO6oT8Hpun9GXNx
h/nHxjy499u5Ln4wylToh4a+icr+wAUZdnNFe8DGgdHW0Pio6OHDeOxpJpsjLrHd
0X7n+Q3OWqVlM0d+NWi8Twco+PjtudaH0WC77gqo1YyxmDMj8hIAj34a6EzHAK9E
Xfcqk78jNIKq2o0deVTn6fQNPhO+qiC9wIu1f4xjN1W2u+rCg8kMW5Ud0enoX8cB
exfQDCiTbnWKrksTh8F1Sfn9YGHOhyIdvIaMLUGbEq6v9rRlV1oRLaWP8kO51c47
ntmVQ8mhR+bJLnvzz5CB14SkJghHL2ghV6z3/wHIhFwv8VOBZTYikLa4ybm08lJ4
UbN5xPTTx6JcweDRBtG7rSngP3ldRkqk48Xb6RTqJdf9Tob6Klc71jdstGqlOnFu
uQWFsKnzUzUWX7AH5BZigYFrSj9CaE9wS1rCXMzvtsL2NKwZn/3yUD/eapcicrnG
YeAs6QF/rl5CooZEMF/367OrDUgvHsIm7kckZOcDJuRVpxkqLmmIjrLEKQoVWVOZ
nMTJYdZPrq7E9QpS9KFm7ZxbzU7TTFXg53Q5jCXlss+T2BwcR+mYpyPAG2watCu0
ljyNETwG1FLQ6GCJjUWuSSdbfJ2T/Eh2r8SSJy7LGArQBu8jmzUTYuJR7y6xL6Cj
XljruAbT004WEozmrZICVPRDc9YhotgDsrTae8ErVCpwl7P7HWqmQQsXq+Ut7L54
ylumBtt2qGnaCxT6YxF0WY6V27XF6YtgT85xeSnZGAlibiDirKY2IFcWhSDfm9ca
/zgTLol/7DMFso1TvQRHUIDGAL+yEk3I4qCrBw65Qs9ZK1Y9oVzXBYU8EAiOTveA
Wm5bGVKFOZbgHIpzD+nazRNzPW7nXIPXPYK8EkzmgyJYOS1+gnf9TqYI1v5sKorM
wVKUh67Fufk6HFg++nW49J35VEJanacbxQAX+EbyQ/QliX1wR+lwuV5Y4LENzqRK
PS7SDKqfixqtAQNQW2t0xKf+F1kG/3/idpRx5gaRRDLy15aFWFr+2WohPlHTmbRC
b396J+cSVx39UDr2SFwi/oPNV4tKvSy6C+tfEMC9CRqY5r4qmtgmVgF28v1+DZqp
TP6ENNn4c+5TTOqu69pitsaP3VKeDl+mlo38umnoGU/cYmqZfOb/niGFP66AoBDZ
TH+sALrmEI+w0wEQRDVGxGVeO7ZS7qANHFLzBfn+sjEkHcNeB4iBXJMCj5oeeL5u
VnAfD5scw1Etmf+fn7AtjRrdQtC6a/S2Vu7aTfmparnBMu7Pz130dWTWm05HNZau
WAwu1i4kAmXbxVdlu8EEOL/VzuJ4YM501hX8kvkedaMabsStn6Bl4YEjdYG6E7xj
MfVMcYCdq55r8uk8XoLLEaMoxcv+W/XkKCNPeHt91Fy6Gu+YlISSzayNsptGCXii
Qkhd3X03X3jtV7f5kAQ6hBDm/j1ldiEV8B+aCpu8qk/9pfulYW0gnO4PvoSu+mm9
yDSD+m6bbsEaj0mGpKQHIA7epmoq4Lx3cQlHZwUawijRmMTTA1SXEYUmkA1Iz/Ao
zxjPIkt0HJFpn/vTlxC4D8LiY1I2gvixKF1N45+JXiAw3AX+Fq1pqztzIWG5M+9z
h9UBhITVqb0Oq7is+0cfcCaesGcluAH0tr95fgGtbXmIpvcvUAX1+suptUy3Urkb
DN26CLwGt5BcGOR11RT4HzIGvYXs9jq5OTZy8F0WeS89f8AhgweqIboyfKqnoZ88
CWbny87gHFGVVFg/aT1/6dMIsR0vAOnmEKidT00pjDsWuBsf59NadIqi/eiY27uQ
x9nbV2kIZrMuTgqib52sduQiMVlTbeo+eJoK4TgF0WrWP0IVUSNZHjcd7zLm7Znw
5BkE37WsyQ2PXjAy8JYEwZwxRvjQ4eFmTB6dwvabBDH/+NGhPo/h6ZPsctoH+Nvm
0ifd3NWnrOz7xI4oDLOf6IrSe0NxUb6M3OKgZ3R7CECwKNThdzYcRrViTXhIEjim
si0l1mIaFBR3sL/ErmgBsXODhYcWq26ROXk+5CoygE/KsZvQJTr2BPwLjA2D8YgV
o9jsrqQwWnvXzTK+YK7u4118Xff1YWO0+dSUWI+yq6GGnysI3BqOpuRq/V4QfnZH
MXGs6TJQJFiP21yp0gx2wj6mlU3R2rb6Cd5ET9en8RXxuRhipRMXzyAcPR+P+1cu
CkKxhmwwjZn08e4e+aEKl/WvZj9N4yFC0IIWsChu5j8n/SjhFTgOQQ2BDdHcllMx
xhRjpv5NxXAVpRDFl6ewgvB+dNyAaeT2ddvmmj6oWrJ9YhdgqaOfvVTmCLJ8gMCR
7cRCY2ON8CYqQiofkHAeXo10NZQd7UtWITOQYKdzE2dM442ZO6dVSiCrOtHSUPxz
zDq8yQXwVl2ym7mhKC6MI9A3J0JePn4lck1JRqmtpNnY2xOAHfQi6pXIe0e7Fmvp
NMfEwWONz3i7RKsmwXYQffUgvZgyFQ7CDPqqm808CCMqbolwTdbRdQx6e2VtL8fn
3laoOf5YCODrimfB0XA0NsAEamQx4Fl5wJf64tCCshn460gpDLXNoG5NByQCwEF9
PtOeYdIpDvz5xybaFFHIwoXrpHOqKy8Tg3HwkKzhOVoYXWqpoaz3zE/ViOWCL7AS
Bh8gqVFalnWU5WCdmczq8YdSC35okwVSuRhwz5hhjFoi7FM4w7f+mh7nBCcEiReO
MRSs4zucO7TCoVZZ3dI8GD3wf5dJYK0b9PXN894SUApQImqk0DUig80Az66TrZA3
Qr9+eR/v7hIaiBp5OFws/Hsfu/Q7OvTdUI6CqG8h7nq0QTH46Lz4NCCyXzCA3EDj
r1aHMb3Dp1zLWgzfQij/ew4zLAU1I/JcoSe4sJwxmPqwzrCV/YPcf+4CeJOt23lg
LVebYBUZlrlJMLVY48ja1YJ6CrmbzQbZwXpXkykMeHAbXEYwWZdyovo2VIDq+SGl
ZqLtnH/3HGwuW8Nr0IIyFca2gsUQqxDmwOnel5d/xVLnTWdWPh/BMvqz/n0PI2Yw
ZbcTRjDPA8hn3mSreczUOUZ0OdToZGlEwVMHhZs3rrQHhZjj4nHchwsdLKY8JoFJ
p4k3RLrZnVZaUCanCHO9Lqee3wJ6TsnAnVogFX99LhB30c9tNff5Y7pEfmHnhmC0
4EuTm8lr1C3yMqYroSW0THuivDeNjYCEZn4FFg2R2KJxra0I26suNNrOfxJRYrDe
BQy1PRceYRL2wryLg22Yvxq1jfSdv+PeNCKkYy3P+MVchYFAMsyMhlzgtcQUoRx3
W478k9F8y5WnsFBMuMawg7yZ6295DwK4erHRzWkF6fhZ1uNb68FjufpOOQPJkgJT
qqmBeWXNYXphdg118T0B2KEGgqyo5SKBjgqDhaKQRFjwh7c/ueWgwPdwRHvIiBMR
TAiRHhdY4o5AwwMZFcYWTMnltx/GqmFbAO76NH98yROZRx/wyVsLvQ6f1WF7txb0
E175Mak0Nn/jubhlk3x3rMfOKVyjAJKsusB0NJpwsKpv/u16IQjoXdYVoPuIPB+y
MUp3WWBiKOLbJ9KNhVYaLyh7p9Sq1T4ioyUpABGvq02EfNY1cqzfNC5A6IgcUD/u
9lEMEPKfQkuAYXyEbuDnzT8gmpKFNOXVSWuEcD/Gfds6K2g5PF85h+B7NfQM6Zh3
wgBwIiy8HZH+UY0ex5TovGnvCCNV9DSCP3Q6gQUNRuMwE5mlh+diNhOIxrWpwxfF
KpS7A0S3czQDYIsAQqQ+RXmeNqhEjg4tp1jfLxSLYN85AuwkeAhf4TzhpveKSuRk
WXrqX5d0DFDyJahUUxpT2muddtCIzkBIdIenVeNFiUsckn/ICmE7BqMhN+1wwF+8
ku6pj4Xa/O2M0C8lp5F/c7WM4nYKWEnHunrf5EUOcATw50W3lrDRDZ4jDpVKREbv
/rcsyXgRGQ4LKcvyqVzCnJrIPA+t8uNqTRpkuzrpSbta/g6MelKsJxh2yORHI6J7
3h4DFnzzy2GwV6zFxy6Y+ButQo/45FQbt9F5wTz6/VECaQJFcnTroGxmpZTCBGyj
8iP1bvMycqwzofXSnDDYit+oqDnxNfN11z9r6ZvHNJso0tBAqICMMqiSfipIQMPi
Xqk6Z3+Y1HYHeyTjFIGqUSYCybwHcyB7h8VUw+uxuaiAi8Y2I6S/nuKRXNLvPNta
Gavhklns2pIzXbBzetX93OskWCttar1OFFkg3//t+WTQJ5TGxjDr7UTp6lqwOuGg
BO1RNTYK0MQB+NXD9tG859uqhbwFnH7clck81wcGHrcqosMogczI9U2Bda2BPUeE
kA0kEFBC041oL4mu1WAuZdCPhAIzHdzfY2cbu7l8jk/7H7EuYBDGWUgm84C7NV7e
Y1p/+fqLheJTz8wsEBGeS4zs6gTJ40CQ0PUxOsuT+d7Wo1vAhip9ij3D2lDhsERA
Yg2BnKpmDTnZauP2hj9DCXyEcKRs5iT8howCWKbJOPvCF0NFDPqe2Ye2w1VxaRjN
k5kKz2T5CcRV0xao0uePGW+bzohGFg5MTtM+2tSLkpHMXRoGzfUc7uLae/h2gQSh
SdMMNDK76Y/GutexaP7uwjCsGt3v2gxPAmrEx9jb8Q7HTuiIPa9MCOtxHhj6Wg+J
NUKghUoOlnlbO+QmnTwn3Cp3KZIyeu+Lu/gs2vbPeCVuEdOzM+/80hw9KZ+43+qs
I5gdHmQkqGIG/Fbt9PIhyMK2iUl91fRTJxHKoFz2lRLuRJYnZfcb7HThNPeVmAsb
w04ZfVduxOHT8L5uqd5mJpYncBvF/KsvNttpD0l6Di5/TEkdwQsHT1bt5eEFhkCt
+9Cg/sdqcV5NmAeAyC+1wTcD3U0VjT4tzj1PpkjQvjKgioQY0SxR9nXS+y6Y1iKI
R3vpfvDf++z2j53S9o1lKhOkHVxXbsVi9dvCdstS50VJcwUpGT5JdhuAoAdRqgsV
jA3cLITjHtuv5vYfsr6fntbATUnkuFMMnzYU3C7YltqgFeTZgxrarDXqWpfx975F
2R/2ULzN+zEFicwTxxpNpH2w08+Vctp50B2TDe8c6/qFuY7eESCdGDmt04JkrLlW
cu67nCRWsGXTzeeMVvNHSJw44U/tWlyDmCSXTzNMNxpq6BIz3Xu9sOu5ZT2xSFu7
XJC3oQyWS5RFumEEFqfAVkmWXw3DfxARDsaFkfmmk1KgM+uYMat8T7DfwkIHrs6A
FAEME911SCY8pD/6Nk6ivDwU/QU32+T8W3f0Z1PeWtv6s7vVc2CCqNoEMzFgM0VG
iuE5v8eOWJXJBVLrcFSP5hws2+CsHwKRlbutNvK9x+qRuQ66eXfM2pJckh0kBg9f
e1Pv80QAOJzfpZak6lQWzeFzBcptJ3ObUIux6YJr7XPRSCIprz+gZX0DMDyWTQbJ
xgMsq2mRYIM2JXZp31NtU4c3vLrXO0i8+2WsRKBBmMgfgjjJpTI2tKH3HhG/M6yc
rgQyPu9Bz0KaY31Gw4q2eDayXKSUbKiUpiensAHpZpsVkhCrqngLSdRromxM2ixI
GhEAyC01GPwBFiYmrNkiY5jmphpcWBst+EJcsVp76YLURS7UTExqeBfm/DRF0VuD
iiyvbinuFR9j2K/azAWJpbx4/RaL4cgb5Q7WQpinDFcaT+MffeJPSSqLpTNWoVd9
/we7AE2j4/cvUl/TIZE1GkkcmmLYEeOzGx5ExFIXI0hzkdx/KDHsuv3Rm/VapXQL
C1UEuX63aFFcQP1+LsFMhJWmyq22rLy59bclx17QJyJlryTmgiKRUUAXLicgN3Cw
95Q9GuWL38CMKlSAkQmJFjNVMofJ8yHnacgndquzgci8ef993VNqKAEPOTISwSsf
be0tfDtt5audCEM9DDTxvG0T7EexixgyCRDfTa9giyjpKaUU6P3AjK2POOctW9il
AdFJ4FhPw0b8n7r4YBwmEi2LAPEI5kOJj2l3BQIhCZwBy1bl4AOTZ3xqG8OX5frE
kt8LeFTT2OB4QCShb9OqShZqXkBhLZE6FjZH0XOOTeaEsWNn8Bt5KfKITtESgLAI
Jo7xAOFyso9wqreuqlgK2KRecq62t3GxyRmwnFVwWSb334eBMtzFRhsT0BxWm83o
3vZ8Y3JjfHs1k0xXFWf7Rb78r5eBna0SuDpC/emxnGJnRoSwZ5Cb5MQUe2tHSU3B
yNtvK9yummUFgn4q3vi/4iDfgyGbQptSn+V4YnHtYgnM2JaRuYF6iDW3a/ZAVVpf
FiAKIIhUDH1kMblhROJP0Zm7LO7Gl9PV7lgcu+KBH2QFS/QFBNJZqlcQlx1T867a
fD0smiYfDHAv8TD09ngzORrpvlQvj+uC1YP2Zla/bLxsjli/Wzi8KQsIu+/8OQMQ
lVfETVWgzsfMWT6PXkPdTPDjrrDCXiNjZpavR0mjhnD7GeTtYcPSQ4iqddGfFwOr
Jhe/Is2U4KV6yxnpDy+Fn+RLnPbdB5wc6RfESAa7Vj+uBSjE29UiOjj1GUvBvmov
ZMm/LAIEGuZBrnHF9CpOdOKgY5i13vNoIbz2zG/V9iGbxaAkUroaIxOrm1nF6hSA
Rnd7RdF2wcPC9aJPUkC+UfkC70MP7Ssn8PfV251gyH7iuQCxa44bfv3gaUk88HFo
h6rVzHcAAsFDuYXuzkEmoOj88hi/+JMBJibXiGuE+DM7Mio3ix4v8zobiB18Uo+6
vYBQpIQZw5J5lug0AqX9C/8MYaNpIfD9Dm4uJra982orsrXjV1WmgeMShnqNsOtr
cCO44pzMnKC5Gm7OmXywscuP0Yk1KZkrPHKDZbOLb8jyZE2ro3WPVrBmCxhQtULV
N5A7hBDVeEUHsgpFu2STKr9b3enyc0IhtnHbyh1h9EnzF4bRajJjW5dkeo07ESUC
oOJLcj4pvIQL7ZdPnmKdSHOJTxhcwO+MS4kWkj2PbUgqJdCR0KGxszl+nflYznqG
/LEwi+OVznz/BlncU9srk9TPrS8hPWBmwdoBeivOtpQihsfJnPY9YHoimrZx3aeT
mIyvwvPtBMnltPLQBEZdIndXNlmFEBsCmE8Cb4cShIskbv7sJVOthHa7Vf6s9qzo
IQcxQGUuZKCL7zcazkoFKD6uiQfcg234UgYd0jkE38ad4GqmUSty9z4oYS6jPk5J
BqWGHXtN0rGRasMELoAGJZcj3yLE3gVQT62J8hLYJjjg/ezG5ZTiPd4eO9cBNN4v
Wbr80uCwSwK53DniYcVEEusAd4ybDkx2GeQU7oUAHnWCo+eRQJQzaQz++1+8ocMX
WZf1VXM+gk+A7Vd9bPfsLd+wrSz+fIl1T/K1e/z6rttODRrDAyLV87mocI+nfcDN
I0tXM2oenSONc4WonN4yNChzw5ZUC7thzx82eEgy0QoLZ9qJQWlpteXi/HeQ/+nQ
PtoOhKR4of1HN7gLmCErO9xfA0ccG3g8ktrrh8cyUH7szggq3Eodlh65btnd+HFV
5C1TaI+ZUUATdedHA2J9iR2Yu/cwSqMGzdxg2Hi7A6MTxnvmZN6ZAt1fo3okt1KE
BrCEXyX4DFthAcmjyu9odX4OTOHwOnoHUFkrONzrkrVYNUPuupfoFQisdzV/5zXO
uDK4WAMLOeY32RARfJv9JMGQJUpT5dOtD2ihsU1g1Ymuck/QYbtxYDKJXIhzVymx
RtLEnLWegO/scLOlwSeZoXhSoMdq09/PWWiX4B/knTph2pttCt5z5St82EpUei0v
tMizzyLXzIotFgUQR7ijKYzBCo41FmFSTj8LO5N7Dsr0Qm9kLWFPRTJoWfwWCUUq
EYIP+Jjvl0cb6pvfAsylx9Xf+9yJTE4KUeIbCQL0paYV61ONmmYLPIFTZaUCWCJz
lCTlF0CxNeln/kCHz+iAqutnuuJTWb1wWkblWfE7vlKlWpM95uFRV0hIS9XGvD+g
RcoEJFhtiL4Zp6rfGlBh94x1Thy0ikVTh2fNNO1lyKP5DGA/Cvgt6jh1T1YaO7Uv
9bBB+k3OJzjumDRsca6TNCBYSXMDboX5D/CtYdZJ4jp7riwP4adTY3X8+bKlF36i
DdSC3HM/nzzl5TqVa277tqhD90juWO09aboeeiR68ZAD1mDcYq8rL1hYbcrUkEQ1
8/fC4mg4arBGPNyeO5xgjwwAgPNFDHfIP9JekDvjZM7yXKBP04ZzwyGci9/JXshG
OSilRk0PSrk1TnuGIE2p/8ucwQkY+mGoCtmzf+MpC6LySSK34JA8iTWdNcGvSoMc
c9krUwnGSJkYYxG/0g0xUbEgt1bdWGjEtEyKtWPx3NC2qAd1jNlb7FFLZWS3vhqb
xMNj1JXtfniIWiMFsHLKHG9mvgBO4bNfJifF6D0wbVKhbscbv+63JKrSzcE0/sJY
fct4UGxgFw1hXwk/hgAzJ3nC31ROmuqCLiSPSCCCnvSbWYp4TEIIqGC2ibevgC60
6HtS862mHGEzSmLm4nY3pMIEICaC8AwzCu2IukqvJmohoPRclN7jZPzc+8r/jaCg
KdJWRUkv47dIfHi8hkIh/ThbkLoRnH06CueI5wm2BZv24Bq+a6JCMVLVeeqR83lG
iCiwSpotz7P9GEcOFE34x6fetvfcUUtvMqpKBFkjGfcWiGT5YT6qyzAbh1JXAX1v
xfnNZ+UVwYFU1R+uGZ2h1P3Zd+cwBu+G9dhGmflkKLc1Gitu/WHgjFKHMHEkKqOf
f+EiGfUJiRqTZUV00GZedusOIkW0BOrnEx4R5IZrGvI5Bvk5MTTxkbqDvzLMkpAc
ExouykT386EVr+gRpXCIw8Q6WqFPyPmw1BMR/8g9unWp0SxzoHMZaNlP7TL/1UzD
uQ91hmZPmTuWxeSm1StANfDdLKEahMvs9x8bqc927/JMdPedc8yHWOMbyAsotJ+m
wM06tbReWBie9aB8k/ZWi+i5uc+A92BjaQmkSwkw6ENjkp0WBYJdbs5qfnKFdTm+
lBGMd8BwUAQeWahgfKSw9oNQNfk4Gll5tUEtyK7kmfsjG4e04sOz+5QsWdL2AK+I
vfXgHLsrIj5TOVNad8N66HLh61xpkGevTf7ZTabLt0yTHWr43nCe4RxviJhrfRVu
3gk4mJrC6L8Byg3PuLdHqcsCJ2LKxzb2/qxCa7Lpz0u8UWGUiXvlAtz82p2C4Z/c
kgru9jnECB9OgK6zu2BtmY4XiT+ssGKOlutIGwejA0BvDVC8NdF0ljLJ0NEEWE3M
Hd3hUapvbkXo2622g4IsXRnjrttH84WaP1CygD6zkLNEMm/0+akL08qRUkFPaOsM
6k1nq0LWNBM3Sx5/lsTpmjgaju8Nlft1FrPWyhBYcilnYZt+FSuIO5SViRWJN7Bx
NLrGhU6jo7YzwBoaB4yT0SEFsewnM37TKPaVOxaXxky7FEU7+wdWWmdSVeea/SSD
CwYCMvk2dlU+CVPK/0LMD/JpibtxH7wyjt6kKpd/nIpIDWeUzU6RQ6KywtomDRoD
jJT4z+x87p1LeRCVNVMFKNHnYJkJkH6TtOJV0ZlH26lKwBjem54d2pkeuTkmbXHf
0Lj6ImpPC4QrT56mcquFiHlMdmfeAg+J/Rp9Ng/c21fzYlRXLqRj/VccujgMq/li
svy9xsFbd54Iqu2AOHvxd/w3oommJdr099HOleybtx8oJClvxEt2/uIT+7awsvQl
lmIBNCvujyqyabTCZmOZFtlVVo11r1h69JR9x6GPkTd1+l1bVqX2/yHu0Xo1kmEc
soP2Ik6RH1lk/nGIuMhqiUdnXvwF3E6coM2Ib03ENMjMZZVL+zPcg64BJTXyyUvy
J9WvtYUPFyoZ1WMwRZWQmfwncpHJ1iTYGGKXAY2nvxfUGUlLcR2RPuY+j4L3JLUd
JD+2D2oAXM0E6NOdy/Rl+ctDIBOLcPxIXhcEsjesg9g0y3FHfhH9EylKQstcXE+V
Pz0wLsSUvFhbm/50owpV7LddJRo6p+BySyib3ZAyKavqsA9pvCuBCMC4RErdmTZF
31wsQl7QMWiQGsjDTHCr9oD3YHxnVeAaWEwiwH/XV4k6u7vpxCY1vxCzFhNslNO8
znVcF1Bl2PCtEb7Y9SwaZTYEJL/gS8CVVafgr+HiP4OLcKqmGhQFch+ZCnR2NiUD
Pk14VcHKV4B8511R8vIr1q0Eic6Dh1drN03YKU8TjOx2w+eQjQ+8fdHLZwcnZXzu
gQ6ok3X/AxjRiaMcpSWyEgAL2LRlpL6wRcuimJnTSWMqSHPGJcJ5srZ2pyslEaa+
vHSouxnztjzS/fSU09qtupTAgUnEzRObmFlOoSy3a1OB4cOon7Hc5MhiQgkl/xIi
0MtqpgBDF7A21G6wybbNJxMRtkU2T8FUJZPiAuSjD/25IBmUHcz0hZ7aWE5hZzAJ
GBd42mYPANDtLdmvB+p6eAdmX0fXv+kDc0QROqAK355zsHlLzJQez4g3zXyX3tJQ
LqBSXIvon2s5wrvV4OjltUg+KjdlH6L+BdSiV12UvSxGmg8rQkP38xVC8J1R3fjW
hvBtmYzSkD0gp3qmnbsLm7RTS8ktE4hPY2sqEmqxtV0k8nxf0wk8zcYd6slnqg48
DqRYpXcISZ84ZXwfDk/7okeOmhirwzuTyjsQDv7a8kxuJofd9/rM5VP8Qrje86ym
0iYCMk59dw+LoNBB8pF3URNvXW1nVBmWo3dBLRkN/NZSBgfWBk0dRdl3iAFOxttG
35YKKq0GwCsKS05/NLPVdM2qqpSh1EySqca0PvlyAI9N9U3IccIIJwWLmQxvfsJw
rcg8hfoJhYzsafs/NYNJqFNq/jTXSFeygA9Va1EE9tJGlBGAItof6l7qhA9pn0kN
lF7CVbWrFGYAP1GBwJ9Bu6EP4oQwqgQV0OniG7hBMTXLFG6HN8nHYF+J2zJkZbns
mOSDFbehpDvoZW07uBgbyWtzi2u1oIsBq3gica4kkw4etctpJrDBA34v1MxKSHmn
7FfXjmk/ksxJK28ukPPqNBu+Qlbq6dLkgZTCoqIEPL+d7y+n2aUJ78+ALPcFO+dr
M0yYIfOXhbg6enqY9mMsqj0M0d7XyG1gYC5oqyEcj4IUZHwOjlIiLlXbSYt5McRP
OjE+zXECfm/h1gr15gmyY3kWVL4kx19rPnoM/3WbVhfXLV2gtTIb44exkH4rR4k4
rdR+al5S1bPxPgyxdHq5+SVQPrDC0iIdIihgJq31wryxDaDl0cG30P2bYbFQ+IAq
108DbYpXS9QYmZXHvuBlSfFlY2B0NldU/k4coACxEMxoReKJcecPcuXcf6yVmF0f
F4CljL8TJeAQ5qW1ritzQJjAgaM1Oa7DfJ/pVYct1Blp9u2oxjGFAtcSWEbYXRr5
mWgYp31f5ZQ5NIiIlBtUM1PDa6RbKYtNBMHG6dO44hkQbOHeIwEQuTjxQXCwpLN1
6Yf26e33N7YvFsL+VQVcm8VhKhgnUTo4I5cFwBKO2BVpv6N/y1q3aiWhCZXqNqaN
fn5NQdL6WkbygXtB+aFCNB5V81VVZXpnU/H8jwtV3+zWWMqGm7KcxZ6isObBZSy5
x06B1fJzrCJPNsrFhI+5L/3wlIyeAjwtaU3MAmX3LsLQ0Eo56sXIVyLtvZXNAxgl
LrSxqoHvgANW4Oos8EVpZkvDz7Z6yBtt2aEcTB8AwpQ1z7Ae7mgukFpcy8EaPyvo
P0pwxRZdLmaDwTIYSH/SFbzfY8/89/vdblkF/x5uXj0pR3llJfMOoCS+R/d07i0B
zaRqaVV4Pn05COdCvUMSx9pmPtHyrYsEDvAjP5Zvp8aerH99tRch5wMKCWdkD5yG
hpgjPPyu8igYgsR3YbTwb5tv36o89EEE2LbsA/JBnJ1NrEy19iLz/jEv54f7sw+u
FSGXFGSEu1ZMq9YJU6dzbPjt6zhHx1dzDirUmGqZP5UI8LrtFTIlzWOOTuUb/tGK
2VJgq/3Srf6XmyQvZQifEdMKycaN6k3l9FFmSLLOFethhFUOCYWO3ct1NCGam0M2
BtBJg6kYjClk4wQxNKWLLirT+OxBvYQFZRecrcDJ1vA3axtFaANc35TlI5QK2+2r
3DPNDQpO/Q6NnHCfFYocVIIVgYi6xLiNfEFnoTAW54xjeas1QishGHrEwa7ZtdNq
oV14z6G1Udn/sRTMjhX9sCnTKU/wQMK2sU0IzFBdx8EivMPecROKuSwbSPtNuET2
0/sqGWCZ63xCH/XtZRLRXcnyMSHwKztaoG3SjvujY9JBbtGT1YyCQoCJzb3I1e+7
1D8+ssiruA8h4u4y8gcxloHXRHNp+/nOUtBOl2hLabsGxDxE9q/CR/c2eHUj9sbi
NrFR53yBxPpn2XzGB8Vw1EYKsFCv6OPUbu3pNG3M6IO/8S48Q+skvdOznDPQQ+4K
CaomX385rQIRfwuz7w4wMD4coKsLQrxzKv5jJM2aO+coPp9I6yp9pbZfSTyUR2+i
D+EUEEMrMbpLKHZsJKUq4vEUE/Akanfc7uuM10oFGAoSYSR/hV9JnoAnGeYnzmU8
7Vv4zR8DnCm+09JXZo4F5Goajua+ThFuLSmHaqeGO+MLBHrRv7K0i6kj/lCBUxu7
gu4/qHbUQZUwS3BHwiczcGbA0ww2Lzujy1ouNFLqjNUNlYGrNsz4tHxTZYn6a4xv
PE8WcHMtJqKuKScTKjv9alZmsH/5Pss4Ax3UiwzX0RPMbndCmKH8wPXsUpvkeweC
gV8roqTyrWVHmEBl636RmJFcS7a+77SywE5uxr2yAOj5oVAthT2IoehHcyx1N3VX
Vqcxy74/BbkNXTbQk0Hcfu/T1JEK7tTnMLvilEunbEkFVg0bXFilJLDHWyMlkIUF
gSBzYc+nOkR5qgZ9mKaqKa5CuPPEL/07RCnYx8oDMeMC38gvnndYJnObG1fBTo1H
7zVHfZIn5eMkRO453nGPXlzXH/5+JYMaNeUkv1TWEHV06YukPa4xkm/14m+S9qfM
YX7vN56s98LARS5PE2PwVAWrIPezYwr2fn5B74EUh7tyZ1m2vycCXBV4+dHaUOYe
NjLPuVk1YBd5Y3fnL1LrsiaPOj7t5Xm71+NcVctoUX99ILjtpGprEwRauEZHr2DA
+KO0t8TKxlSYWHpl64151YoNwBSaMDViPwgVtyCpUwst/OPWn7tuAfhoEBIPxF6w
JSJ4Obe/RIuCdquKA/h3WOncw37BsFFctDC3wYrf0oh4G/TVOER1XE5VOCJshawz
xub5iyKzX7Ss5eOFg5K1I48Rfb4J1irIEuHRxZxFbxCrZu/skahGueUVFwFOmGzY
+r+y5c8MU857NGb7f0VRYoEJkeehxx+JLoi9pujfHZKolUK9sF43PeHjGELDGvyD
jLqYPxgmD3P6bFYFN1O9HwojROg0f6pqxFEH0gflyRv2VSBn4wbh1aTE+gk12Qec
/zu61EvKsGt9Y7aJANv+nzOpQqEI0M+bzBJEnFXIIDwnqIYWOvXc8Y3KG/ROU88m
71A/7imt15tqUPiT9g2WM3ZdQbDyK/wgx4Y4fZVRgP4a6kGDGRBqKJMkJ+pGuXZv
kQCEqmeBUGpZbB+N6Mmvt8LBN0zdGCgyzXDmEHk2B3P8a3gcQ4w7qPsmJTShcI/S
U4Jflzl4Hhj/wuR0ERJjGbbgRxH1aq7JDueefN0OT9VHDY0eF0FqaHPXTp8ZNtrs
EUj1QaHfELYgKC2bAPfFLtdTDPnAzMgc+xNacuXHeCi8mTsedbuMpypmoKHWvMrn
aTHpQTlAKhokEpuiUWQ/cSsyIzpuig8m/RfaVBoqM4JmTFlP+rsSM6jEDGsK1oXO
npW1VMJ0lHhzJ77BJA9d/mCiHjLjlhYqVd4rXEEAutNicCYwnRKw+qugQ9I+R+S/
IxirJ1ljQsZhwJzxn0KV98oJNnSUX43DUkO6LkgoORx6MloU/hLzTM+xRc3HrWtj
S0h3PGYrOIWoWx66ckEC9eFiti+ac2F+RDwCq7tWyn7NnvxYiH+A9fjj/1CpbZ0h
sd1nfd/lr4CUiSVLEn1IKY0xbyCgf1J9RZ6OCejXzH+1u2++XQokZOLGZj/mXiX+
8AAhw2FHKdLq5Y5V4AEDkBksu28I6FC7SU2ytnIbH7Ns+5kX4adWr6M2E1gnHZSG
xX43o0ZFkqbbDG0gFAIyB8zfdC1Rwqsd5RMjWn02ToKslARpLl6j6mIPKBmGmME4
gBnNd01Nqqc9/05pkej3iN3jjFqo12Wf0dXI8+EymWD9EcapBMdT155Ro0ZOcryf
2KZ6tVCZHORs73uvodsEduq1dZfJvgB8f92rdPgdmlRaszE0PI5ZeyHzWxG1prPb
eIjS9UdEu9z0HNzRj/SFqUDY3ULjXTsTHSocQcvc1TcgsZOvDHagzSGrraqQrSQa
3udIHTM4eSeHKwIlLtTmhQDTtdaECX5gmzA25UgWuMYJ8OcU5N3ggv/Tdwn2k5TU
E15qThOa2gwwmFudUg9ySmW1/q10LG/ulocfIdwhCj/onKDthVaJLnnEmaYYqnUg
wkms/MOn62nYYvvaY1Jkt93B8SWUv3JpykxBqs0hrE/FRsa6Asgy+EiXpvYHiVoS
HxO6PdhJc3PY51MeBbVMbd9LTBEvXdp6EpsrO7xEEVLBJkqK3mYifnqBRQ3RT/pq
LNxYrAhd3dUgFr+6dqmfUkrjNwBcpyFvH+qdXRf0oknJ5A7m7yvd4CZrlbhVVPmG
69wKXABDWYAWa1inE/VZZL1EZHP7AIkajZxmtiQdDdBrAHqv3L932C82xmXwjw67
g6Wb6bvv5nC8f2Wi6a5dTOcmqp4HaRyz2lGkYVpfMOWHQ603sdFNbHqpO3b9HE4/
28RiSxABCBZDiNR301O/UC+bySUeiPSGt5obkEUlZwGdjXniVWmz51SJkMNU6Fqd
KVFZJ3tAQk0gv0ZkQNmRMZsEPlHJXUwx9oM70fG/4qShBFoeR68BBGcFZcIBhxp6
B6tUypsjKKCYYz0nQWoKm0EoYbcyEyppkFexf6MAbVQznbr9nBB2CAuJOf0u7GO2
c1CkaRplDl4KpIJJOgVT/8VG6dLo2RC8OAS4HUxAzrhLphxM3zFjo2a+sPQtQ035
2+zZV4qfPVNh/zuIFuE3YlY79Gp9pMUMwqPWh1UJ4nd+wNfTJeVPgKI1eisCBTHr
/x2PvRopUdCmL58GCacXEbYRpZiXW0YtuQ2/1mNMsysWQTLjkcCivr2LGSgPaKbB
scaqdMlKl1UYCaYbUhfXeuX+5A5d1MM4tlboI9Sj/8EOaBFMINad4jLz8jLNbVru
36LF6s+OphKvA04BfycGY041knc9OLRAqC5dDuCe5cNGCgVuupRwhKuPDBpiFwDV
vh9akLJTswXc8WSKY52Y192d+duEqxbUzHkZT9U8S1JvNJsyu3mwCa3Iw0wBLH+V
CYdbj0+OjA3rPWGCD/DEM35FakdrIrCoSUcQ23ofJns3dqB7sM51WuxgX4ODcsTs
90PW2Gi+lde45HP4AR1ok7aHj/fLlFGHwVmvMAUCPY2vgCsAMnV+M3Z3TyDH4mn2
e99cu7lxBq5gz19febmpY7VXqh/To3arBRX+FQgzzL0VENYnJ7paVqr0W681Lv8c
wAPKK88Q8rYFU7vt4OLC1Gkg7ll3CBmvpp8dwKi7IL3d1Uqj59LX1E9Fp6hMtpD0
a+raZ0Y79hdPoeVoxC5b1K3BfscPFIF+KdD1oNPCeUEP9ip4SEZevYWJDBdh2EoT
kYMgOsnzhFAXSXb2uZBowc2fmNQPk76S3ZMBxRy4dF8Z2relWFXxeDLaIvHRUw1M
ZGLZNx0mxEg25jXJcxSkT8zvehRvKmAGkhQZuDVhnl46r6/oc3P/8K4nJ2ggRo1P
KE8qyN8RlHJbxxzdndeFZvIwXeEMvy/7PFboj8+jyRqy6CZEsm2soR8clrd6WHDU
nPKz4xl/liZ+pLeA7vn0u0FJ463NS0JAkrn3I17nCkY2uI7OEWvSEbj5bP+Dk4Zy
06ONROxzntzLRz4K9HckrzP/HxBZ8fbXCWcqzv9gTNCHtzvQxKKuoHZ8f3NPkeTX
nwo7TDzFgwGhWSij8wuTL+kCsI6js87aZDMKpgmexfb90Uk59uS8Pe0m+k4jTzjI
IJFnJHjiCHaN3ayYs/kEmvyyG4AajRwRxlYa71mGjrAkG4+PvLMv6jBoEv/wts2v
PaZ8wXbvA4euLqrGRxmxAdDuiviZ7Qg7RdhPxauX1iX0qU2IkzAZYX4W1hb75pPi
5cdG2VQRf9i4VNLzPm0NCheChGyRZDXPFy9UCgTxoShNoLCyiGY/56SW8zAeCqO7
HuwXGSlvqeojL49wa/JKb+Cfe/UpBpXTx6GqCxXN0LfuGl28GQIQ0tCZw9R4PC8V
IwLWG1bB3QZyvf4LF3Ajqy3ncX842Vd1O7cjm8orsDS5x3V09WvoP81QC7duth/U
7VNKRr5fTUJTKpRGZNkNuUFofGsIIkXT9jofIjICDQYjKBRmuVvaGR3iDpcPfnML
n2BfBzQGpPelTxZbWrFF9GQCwaOa/f0CnsNF+hmKnmVh39VyR9YS3gp7RIvZ6gYa
tqZcl4UULHKt1qGxI3opuudtDg8Diijsq0KyMNBjiJcFMuoAdfN0RSDzCZ2sQ+1u
+Alehs/BZJRVdKnT3VGbsVs59TWMBpGX+xaQ8be23wVLQi0IqwYFfeQRRelvwgYI
cTceBb0ZfpbHyqKtRXC2stK/xtVD/rXUcRqHBwhUJdTM3cOeUDQLjEaKRzj4hTme
FM77AilEa2iADacMvk81/7CPIzG2NHYYre01rXe2I+g5XMMdcqRCpmtS4TAfBsiK
x+WTJWZmPPock3Yw5PdGUZdSUdMfa0YB/r3uoLS91Gaqr8MYStul2JZc4ZcwuW91
aA+Cad7qiUyXjWFDuM6U7PRjMake8aGl0N+VtiaYG7TPeu+0VB1RU82aDmyFoNDs
VEwM2Hoghuus+gqlO9Sz8qGgNhHgotFK4/llnq3GEK/JTouDeJD3I8WFDkJnam83
ruaY6Law48NHNZONmgYvfWExMMerPoL/zsz3UF5e80NSeOIlE/6Eirz1ZcCcPZeP
+sYP6yeEMDerLIhYRejCu2wsE0C47zBlcXMHt5jGxyIGyV6TAm5cklBeLMT/TyHu
olg8ICb9ux7UOnZaiBaJ51cgMQKVAQGWILk+cYy5JvD2ve6v3lemYhZIRmJRXzHa
lcr/hkBhZgwic4tKjjWmz4LFrFLpAB+9dQoGg0ZsUP6KMLyEDDitKLGCymWWFbvw
5/VofhfECTxd53swmAQzwhf+TAfF6D7v8hOaoTasLkX8suo6+JoowU3GYMatpobQ
OJU8ir1ZbIh7LEcxiQeAAV3wp7s1yaoxklTTnWBidFVxI6Ep5JyCOWRUfjr/QVds
QUhnNc1vVR9Pd1HEYW7C8rwSEUwYDMdv0OMOWjpGPxDEmhA2y3Q/Iju6nZaKoPVH
F5j/4iOa7WQQoUo5/HgAoCX8xqmbO2jmZWXcP4NRD/SCQB2C2fgoyR4VRFX7WgDk
OEymIzoWoqdxX7uo6+1TcpllBGzH3yi/yVT+VN1idhdDEBxRGzJXq8ZkvTgAs+Pb
WyblvciXcrQ6UZhFvhK+GyhDe0yrtGFutQsUCs5n4fxl0uPr8sB1Xmfba7+Sx8dZ
UxDimrmIjMX8EuRLy7HcIFaSWnlg3ijCM6vUVLUuueoexD+IqlFv6DjkJEWlx7tV
tFGy1MoVD1lucBeVRS/hjnr9+LKO7PdtxPfdxAqUzpZQYHIn1Xvb7yLf6v0KQZwK
McWtiOPglpKH5YjdtqALyuf/ydnwsicSjLw5rg+lUlgMNSNNvt5V2mGBUotWnuqO
ViZ+ZucQa6YE98mBBcWyGbMwMxTNDunxt1arXJBE27MC4HSr1r4WOTY3Ba8j50eL
JOTA6z3xRsvChO+f1YcQfmJdLoPWfZkWe/UDtjh0coyV29a6oqTM2af07zFoYPi9
CsuMM8OZ2LJGVoMA77ofqCEJB2X4ef7wuCaD1FVZm2T9mtfyr1QE6haIHoplvyak
Bfv54FjHX0cwbBfrjK01zVT3DFAxWO4bZojA+mvFvHcTQF4hFF5IsZz7iyTxztZX
GLEJ6GsjKfWxd/ZXALH0DNYZZNxB21Xr1k4OHXPx3TS80jS4sgA5s2Ym3cYq/50q
e3iyO2HOLWuB2YC5w1zalgueQsfqzTxmqPWFR/GEe/RIAKtixCtMJnZqJ+y7DKAk
kB7YDg+2UWHHAt2fK/7EtCbXk8pSnuIxrVXOk84WEUhzsY3aAqP+bp02KlNx05hL
3eKjFiFO6p6yLTU4jyLWXQR4vLJvN0oc7Wbc6pg+2+lMps2IsbHlhPLtfoknwLnv
6tOowSIQ54REXq+gmsXuSmfoEgLZ6pwGEXWSD9iFYx58kaMkA80qH/Rk740vRGQM
ITj7aKJFKKA3NpSXo5jI6znvVeo0wuM6KFTB0bRL1zmlv20aLW8o5gPhGVoS5vka
lH3X0rOeTejVLRP//muHvjj5m9z0BrCXyGYNFiyhZq/8rUxXc8YIJqOmh4af4OTr
D2clcaz/ctLvOGWzD+TdiIAOL1s57rnNAjROZXHibJB4Y2+iiJOMud4Wz6Me4aWs
vrUeFpjrETokobAV+S61n05xNCpn9v3Ji4uF8gLFaz8WDM4Mh/i32wMqqsKpMRAx
XoxgQc9lw13y6FvssblYOD4/0WIU3UwvTnQrGTXJoTc+rpxERoXN/SGAt5BfESNl
uDc1YcQkQ1zTcE/o1KRLZjcf1YhGvPXS2N+TE8ktd3Wsk6IfKNQ/aUvOfgzJnOku
D645Drm9GrQTHjug2sddQfF8H5M9jzonbrL5WWCNfDlPA5dBGG0Wcnl0NWsLZVD4
G2j/Pd0LLlXBEGrgf/eKjdyulKxqAx3YLR15D/Y6Eixf5bQLVqL3a/GLT5D8d33C
nX/BNHUWIO61P4eB22StpzQGTL8vYEimkRhZDkfbOEGgarUNTCUoKDM6+qBM4/RS
zuH+GRrjCXxVvPb7rlcd6JISgBhGI6E11Ta5H0DnCkceKtRsuHOeQZaPAwg0jnlm
VPbl3uofKAk+327mS/LoMvbgDiheABODUR6oV/potuHUHcnmRXyTv4/W76vhaOr1
tmd8qUL9qI+N1GnkT34IZToIoE6vrP93J4VYKIeDz0eWwVJEfAoNd4dZhjEJriIr
cz8wx1b8yeFbyGW9QsEF9SFtGkPP8eX/+w/RRoX3za3zMNXCd9dxRi/S1CnJ0xgm
7pBaYhTEi9zJWOERSoqR4FxsuC5vYQqyfib/I2zpVYaxfIaomswf6M2GTpNNzkF9
imUZBY5lkM3Mmf78/BSvjWQ8GhLpjJKg0Ga18I5+kpNZow4QFPjjUPOHbGU2qDTS
2EK4vA2xfVtybnh4f8dfBTk3S6geod4lH+WcovUTgHQ600PeXOfin8v1HD1VOVFr
iy4f7ejf62SadqGrGHH3ZNAr1c3aZCl5iYouGQoj0Kuiap+BtmdRI9j2wXesxCOA
TxvAgs5b/1ZV7gtymZQOqh3WsOOtutcEsuhan0k+ZpxwAcCGirYKPxfqgv9Lj+tO
ycjCE2LiDgx5sRmqherFcbdu+JzNGKgen5+oQlAme7IInkBFURSdVI7UaP0R35kz
QoKxubQuY/2fPYWF54iy8ERH3aJ+3mDQ4HWPhIKFxCLLDJTJk6IDReM9pysKSpRC
gqtsVHKqH95Jl59mhoonxSciqHRjiRqhaPnngBD1UEeA+2T8yef2nB9+ao+STke8
C8tRvETrG/lChitcpIICP8G6wYtWg64Dnt4JAm/ra1JyuwkaJvS/EgrACKD0axJp
1RQzvDCm/XKChK6/gbU9JaBuCkZitEyQrbFZo5qcizusam1llaG8cVQG6QzyKsvx
m7FxXxQ5wDXoNstOrcoFtTGWGsMPp+9dNykce0eGL+iMZWqkN6S/juSFd9rqrEb1
mHVg9RUAbgkgjcHHPs9oZCnUdZ5ZImDR8z7SyJQmHz0iQBI4XyD9OHW77GsOj9SN
rDJj7epc6UI8dtHguGV4IEbuhPWyAYRCvFL8NbGY4uvm4t4CVvmFoUecavmC4zKf
axVwSucP/IhbK/62YfktRTCCqPgqk1I/hOT3Ulwlq0UyD81EhA8y4MezuZaMpAyx
UWs6CKFKmFdPk4L0DPMbFU4liRqONMVscmROfbVDeWiAoa+rntafrWvenHPKWaNf
S6kLCg/zpZimkZiZmM8CrBP7bSxOaCe39O3NC38ZgYZKQHV01PDqJT5MBgXIyw59
u7ScYoPNtVmorOwP2xKeGMUw++wv+Ox/Aq56crsNCcZZ+KNmD8Vo+jS4W/U47O2c
v1xzAQ5MSx+ctxPg1Dj4Y+pUAYeyB1A3+z6aLYR0L2+IVPva9oa8xgxUwxLrQsuC
rwL1pX7Ip36KBsV8RTNvuiKuXxeAvs7xY353+T5MrOoKzpjoqrK89b1nVp/EDnrc
3IuNjvH7XETjptrQST7Plf8kXksymbPA0prrsgS8h6AyjrCuKz7PJkwVtjFSJ8bm
YBpW1LrZXmbrB/e/12wSuji/zHx5EcHzdDXkBHnSX7gg8YdNdJbAPd8dD4o3MuPv
BCgZyxmxZj3A7FLI2rHYM8XmibfYdcGBwnS6dPvYSxUvoam/cO4Va202vDInlihx
Rroyviq9obCECbL4l5XLCljmEsExvX+4cLvZntgZlHDdf1FlGvjBun5KrWiFUc+6
jFhG5ruUdhTJGuAlznibgBgzQ1JFtzJcitmdn6FTfTQGuI9DixopPUiBtz5BOHwd
0uYQRwO0iM8BBsrYo1W99cwIkwHvLa7QudjLgnT3vfGK2rDpKp1f+P4wlZ87GqdP
CRH9JiDm43zXO4oGlX7zQoK+LVetN8o1S0XUar+LfPewt8IryaP/Kq8/vqBgKStb
XCaVojRrCVNRl+PwkstjMhnYDd+yc0U1jerVVcnydGVcAfPJFkF3k8rw0f++Uyyj
/ps1QKqM2NS260TGnG9AFvQoVrbrEQKTuCFnQNSYC7TwTmGhIjFjk6w7LWNi51m+
TFyicOjMtHT+mkGwdeborBGE3vw+y1uVCY7/ORYDowgbPLer7kxNjNokECrtjaq3
VRHD7sNwz2Xk4+B9Y/iTStKt1XhIsODGYeoDqspM+KUp9okwE3iqWhUnBJOVQQ2M
6W7QygThHFTh4VGHQ8G3laxM8PYQgBuq5x6G7HFW9a9jKiazdqKu9SxnJ7D5oI74
sJT8rE5sKOHeGRSZM/V710VN5x9H5W0jplUuBHFJQwA0zpmA+p9VTt9n9ZVjgGIs
FAu91JET0JGP4KTf0MVVSeCIxE5YJXCSpDVtZBw51BEnW0zysy6+EKd4Dzr3hBcI
PrcXzjp1+lyFA0pRB3kbWpuXiXWANf6pVkmrmOyvqWa4aANNnAcWFy7ev9yS8hXt
ReB6OvUtyx/x5ELGRF29bpE6hZB7OtGYhFdObB5aas1V4hKGDamB0AUwGQpbIwgN
rmBVSoEAgsVYb1fOdz2gFYX+XxC0D9jWCvxkgBScrJIanYTZogfVK4Z9kcMRnGwk
Naf07vG6RlG7GePkJxPaLaaxmdDcMwNqSj3HNL+8dQI0wIe1HZZEw6s8LtLsv7Eg
EmNZ0mkDKn3I/lvU/Hkh7ajPKU47Xo3yIyGASBWrf8JK1prqWEdvMC7g5oy8aVVF
/7JlYPybafhI6HnnAwM3mHeKgB6zvsTjuNNyKFsHfdBgJBRI0nE7dcded8UkMvWd
SUIqZZY9bFIiUHvNi+I8xET8n1kSZ3dIOIwKD0EAXaefqdHF89I7nSvFLCozuMX6
fHPFrpOBRuwtyW1iaESkS1qKP5Jxxhqus/7QD+MQ44ip1oscIzlf4SSPDwGEP/PA
o9QyvJlwEWde1VErDro/3bC6gZM68ZZjJxPVgg3QS0gc0pDztzZfhOvZbxfhfIQA
sk4S2GLpU9QcSeqRKCj+E38cuvmyGKc4d0+OuPiySzzEIT8lQlx6RNxClWx0yo7O
ZJwQTYn60bSd8n/PTtBXzYaWPSn5wI740ucYIR62ymLAT9IQqDDYLuoVXdWq5fvM
1Qpo/I1d994PymGF4ZdBq/qDc0gsKdK5q9bIs5aQxtSLtHET72Q646sCLqqS9kYY
VIteb0CTHksXOnMYUND5O2eYuHrlnjzPv76TkVNHGUCsROlzTImgQo3jm62MfPM8
5RuKxCkSK2hbzSGlyYLoPBd4zi5AcOCkWL+/32twUBpJyX6YxSEV5P+0DnrMfY3H
mjRDpqldKStfTiDKFnax5bReXP+RcViAScqg2fR8SBAKuNwU7PCiE/sxMIPoKFIh
edK11d63HWuPvt0NbKM8hSEM1YlF/93H6pbVPszxCt6HNocxTuPOnMx4b+9CyGoZ
I9CL/vQn8Gk1lwKQulQMjO3e6SuIEc22SyPrdspxQPVOcIar+ytkJijFmHF/OYYP
a3AbD7u7ATfKuBA59p0V4X7lcrD9XXHd0eNXGx3G3LBlN0aYqYDPRiTz0+soubbp
FXHOqPAJ1+TToOu5V/jgGek6D0HVa03E1SK4GUg3qAkictW8JbxuED9+Otz/GQ6O
W2zjE9ZzRF/ZDCSgPQc+hlFBSNi7A2pzmE2bVZPQ8ti8qNESIMyo53BU9J0J3TDy
aJvHW07auT9cD9dxrASd3mz7cPbAlLIF+QF7Wt96a2u1pfnC7RZdxbMYti8o+wJv
FrLusHTwCDhoJO5olLYnLCx+L67dF4WzQPkwhVHvWGrSV74NNOmVT1qumsjgbQ4N
J8a9B/bESM7tS9rW3HdM59TEiHvPYFOO45Jt1O67jr5ORF8hGmnpf/qc9jCKBLRK
4vujT3nFg+Mpmoik7pegxpJq4tWFnt1OtSOsr1tu0uafZ88fs1wFQd6vDGYOzobY
emVGDwqYQ+qNontlV49EdUClXVO/0YDB81WktamtCihrXHjCv2nkAlehr5Nfx+TG
kYD4hh10+UWx750Ght42a65XsV7RKlH+Lb2uQfZsWI/HL2bvrLbjwTKUzNukaolq
J37ATbrYFZJ1bJqTF9hFreZLg7IwawuUgMcHMwzZ/zejXhy05HVihBxbOD211LFb
aOP3466CqrcoJ3rlXEN1hxYQa085d3Nj/TQ7DrXK/fLjAIdSiO1OQ+wOOX5SLzcB
7rPaajhlLGA/wzZ1yZdafQkNVWWtJ2k2WVEUr8TeDEVZn5xbtcaURVYMUE3csuE4
kFdmiYJBWkqkFMmQ5oiYziWTRhXbxY3+xvdpqWQHyHiabEe9p+tNh3HpIQQvGHak
c5K/Aet7BQrAw6CJ9jZKchrHQOMCRpoqbCbR2x4M6EfmMRvYipHkCgtf5iSkeg7y
vpBoHvCYsAQu4ifvAU+TS94TrjCpeXyvqETikJVsR3eVc/qPJguF2t/UQCzFs9eo
Waz7LghCol0eN1UcY34LJiA52cviYm0Z3uICrufMEhCSDtH29WzEvJ3qhg9UYFXi
OOdCnVzhbwf4Msm9z7fYXNtjAxgzgcyErj5hBNQzp4bsw6bCKHPrJNVwJ6+AxBjE
BCHKdCBfCm2STh8hT/yrVmfHR4o6are8BJTHp236unsDN+yRHXd9bipDhmDBDsHL
KAUSZpEa8oZF9xHfCHv36DR4vyca0sEW4kuL/g9Hpc+y6CnFE6Wg1iDXW2YqLfW5
EZ6t2Ka1TVyTlOsy83mqfVHTLiN/5UVua6QN8MYfCk9uPOaFoVr28jcUZNItMsXL
LyXM5cQCTIN+YWbv1Hs0YZhqpbcCe0SjhvceoAFQNt6fSJ8tfxiftqpufFRXSxWy
RedC/YzR/rMLhjTgTi72HYQqc9pecTbrgA4mGyHkxHNGJmJy96RxnDVCQIMLYkwP
vsFshQRamUlxSjqFEHHl6LI5yYQQMqOSMu6SNr1mrNYy7EgY1iX+NzQ5ABToJHCx
Ul5m3ZQuBwaKewnTsO1cT8wDmAA9yoFDbgfBNg728k6bjmQgkwoGH9gXBmDKozXy
hfXleUlJ20sCh/D83Gxb7Dw0Dufe0NlpVogGUOVkTgDdrs95UM2uzs5oLD03blY9
oAWjNXfZY5eesersXM0SBFkqitV7yESLn9geiU9U4RuKqqAribQ9S7UpauWm3/Cp
8Il//VsK7nooxCSMCisSZR5HuKHNObgRtFdyaBFX1BApq0YkC9BrvSgutWOJY/pF
LLfmPVdjst+lC6aSgXib9KzcfhvQc3QYqN+D4khXSmuRULsDPYm70poHMdHj7J8i
60h7RU8Dm3RdVV2IpPi80+sfT+2gUBs6Bf0V5HHD2AdTT/HoW9PBZonEhYlvmoCp
kSvalN3K/WfmjzfBrhYEhxgxrNyEIfsapuuc+vPmqJZZbhbwa8LSvNENel9I1FBZ
4ZB/FPTP5NyrrU9g0NS/reWyfLnPkNLlrGfrXYaa+Z+n1kfrB+3kXXChzxCRXq8M
xkYj1Vm65fVnwX/3tevskG++9iwEoQ9aTdit1XWXQ/hMT9zCvTJgrNNC3xTAhJIz
VmYpuZ0H63/tOz+pBoDDTObwmWXQ+1JxXAPiqR6JDW4ABNJQ8vrd4Kj5XlAgsK+e
QSZSmRZYIgpN86H7B1e5J7tJUGuA6ic76tOS0T2nlJfzifqIll2TH9cL7RlmZtrm
+/JW3urB0bTHb9t9Mr5x24v9qo7A8IXvt6q1JCpZ7E2hPx6WmhYgSrf1UY55RfC7
ccv+ofaH/Ox48MmvU8wk8agpKUEwGbXkAprduuWS26XLOWl74NN1d9EKzpb9JRzv
XgOUFq2kN5CGAFf+KEOX5jxo0P03lUKyo0SBpPFI2IH9uKP1yF3EeRQ2Y4Vzql5h
BwQRuOsl80WFfEMLJRLxMa81V9uhwwM2ChPwSshMMFgYP+vLxo1aRXIEbuZN3b9m
KkXRVFPoe75mcGWlvdvVW7yYxkbA/PppmE+/qDvUPnWnpUIGbKZuR69VfXfNjhkq
DH4yPoWITyEwh9R0RKwz6ihM/T9o7UmS6ym5uQY4tAT4p9gFhMKsXY79TYNsuOiW
EnozoU4qeNzjU3YSh3wxOz8C1m0xR0cuAhhvaYWipFV57y1vvK+VfRAjBQain/B4
Vlpp0GNXOUlQHd+dZd2lwMiu9HhJM5le9ev7wlOcEOwNg4E5YW+Ccm6RHzJ9jdQ3
FZ1Nl9zz3MglNUuSDiJEsMcX6okRd/nFgms8lXqW5lVGFox4Pj1a0OOMBG9KT+JK
vEx0+SBxXBXNjIDKRjtGGrinW7388pLKYycOxRXnGUsmlPE91TQz+DRgMQm0OQxe
l/L6qon6yK+A/qrDcx+qTDV6YYBZ2d459OqPG9hvUOQx/xa5+eUq2+w/JP1T6tJr
RaGoHmdCoURzoVntEM9/VxSP/y0NrigbP9EMwXlw0PRDHikoDeEgWpamFGdD0YJd
iyrrCAFfU1oVwvUSSpJSiqcdt/PxPQStg89ADWtHDr/gUPZcCaknOdnghbnVmtPv
hR0TNc4hz0APuIhYN1IpO0fPrTMY4rdUHgr0br/gvWLgORxGR+HkCU4bWFYqxxQY
NsINEp8+GbcI4g9QxzNN9oOiE6FyU8yDWjisCIT/eYYuhNz9l8tKavm2ZDdbqY6l
VmZgSCbKDbS+D3qhiRZKofFFKZDqARRDGetAjky4ePWZHytzunG9isPxs91oCF+8
EbE/u+A6bMFTv/+O3eFdHHcj4IzJBTxMAJspWg3SK4GtQGZYWUYke6eiwznDSLSi
1v270yG1w5gdVeD87RBNu70neK2o94PLTCyYPP/GFSsP9xZecp2/3xXQO6TRiglm
eFwgGWcZoL6qSTTmcTv20mUhRPjugEZFlJZTZBpwxTrJd2YhsOthdV9bdgOKKTnx
Ao35duSQbQ6DD3IlsxO4SdGJzwByLHWv4xlQhP7ckgyAkuPpiKJDJ5uw6eU4D8lG
fddIGniEg6FR9GvGBSnNPIj7+jFNsQworCwUSfQTNADO7oINzJ1dkPpk2VSM+vEp
LXWWyZvIXxK0zWK5zzAJ7bDx3P8Oj1/fAA47TUIKR9a3wU+KceBOH8KstPbi1xKG
NFuqNetIC1w882bQu4FtuYv+rrpaoNgAUEmChhLuGIGJHAB5MdpTbe21U3LqnlxN
EO3dCF5UYFS7YtDEu1WlQniA/pDSLVEFEispMTAw24mb9dlnSEoYjB/l2K6vowoJ
xtUa/8k1l98RDGzRjdQl58h2yMOqQw5IB8IzvtH61ZuoArAqf8UlU82gYxMn/Djo
WV2aPhAnAfgYfniKZ2yJ5c1cMVCC0LxPKeVNRJJJeQz/hRHvlF1F+/TyiBXqkSjT
dyvoP2Fjd1GWyVqKUSn0uaXhPpjl3qc++RmeatM4CMZ8c53ikyEzmCI5+t8lqId1
TyEewtGKksT73ImCZ88EPWFszm95h6S5Ba65cJpEWDK46WVifuQO6Gr+a8dTfQZ0
aPekRQaIoSMPzEpvoNh85WNfRveBigI+9zC+zDUE8QqtybgnwZRz9uGb+ddbJeny
qbGdT4hqXIZRNO9E/4ACEDqCgxPAMz4cu8cqlfTTgoWSyVYxMJ+TSA8Fgyoe/WO8
SwaFSvPZkvDfiqSSd9NGQy4PGclVmxPDo45Ono0ziJqfZHfZB+g7AZSCoW4g7REM
WS93AadzUnHIjXokmnCHHKbyelodRMHCfIGPDeshq+luUuX6twtwSoGC3bfvXwt1
G6DG9yeT7tk+9Y1fr5JidVqA94OKGa6ZWs+Zz8YGGDptE5WcGHxOPf7yg+JpBlNO
q3YrAiYv2urbkCiwSMwhzU0MptL23KHJnzTBj2C9aZOxeeqwvGwG+/85RjeOLfyk
ZRzCc8d2TWsjUgtsOTJQoh2fynYEpMVPS+0gaYv76ZH7/MUioPXCRCjAczPqKn2B
57uoBF2q+qRkB1b2WNg5aSHct1uiaHlLm1SPCQxerBPgLKdVUUvduP8e4/A6jpLg
qnYDuh2z6y/iW6wyZE3obJsCqRd4QX6lVZxo79ZVZVSmgfv8c84GPE0Oij0ObCIP
v4Ntaxk1akR8fGkBxzxeo+1jxxBJGErW3t5djNyHHAPRhl9MIHzsAOG0zmrrSC2t
mX+BSU3GpAVmu7s7XZP9BJ1iW3ZWikAAXJ+c6eXjJd9AP6t1JK10QkKKkfC0pSKI
xbyoW3SGN3TfMFiAZ1CuafS5k1Fv1hkFpcuJ/CaEYLnltnbPw/Aj1RrvrtOV2qcH
6pnC2DqTwkBnpLts7gzRQb3HuJW+YxHgi5km9yVhNWCCe5unjuvl4q/YHRAYGA2M
bcwwBtzh/80f01/6ZNlmvzB/JRy/Bs0W+ylGfY+DJzpRew0LG6bZ47FaWz3mOAGI
bC73Fn/wI2kXtDeWi6g8HWpdfniL6eyw50KFuItTKiKxDY/RB4qqZ3Udwg3Q5Y3q
CHq0tDpSC9uKJTUIOYYNmFDi42eFovlBs+8FW0MR+ljG5M6Bj0Gz8Id1Hy2tGaLH
CLxzAASWoBCc1UHoO6CFtrKylfxyUQZOtk8FsrtHY+4O9W5/Rk1G56838QKY8Reh
BGEUgtaw7xuph84Cn9O1k7EpDIC1UFo3hopfCghhxoEMTmIIHwqG7qHDcQY2sMfi
1GKpV9myHffzq92ksq4XVElghAekhOqHyLg3wMWoX1ckHF3IIHRXy7BE5ZTOiWX6
5UQpQbE85T3NmGqkRvkR9Ei1RYTFxxT4oTrz5pifeE3g9Zlh/rEw3vGmNtzkghpq
cYu6DxuDlZ/RRH7Ax6iO8kJnIlD8nFR2FvAbSZJbnTUmOE9+3cPFCyzFFAAONnuH
BQcVWv+YhMYNQgUALJytEHN+bhOqlNspd6grfFXJx2aSMYvb7nRF05UXqY05174X
BJRve3eXmC/wcoBL6XjMtPthRhwiy9WEUTYnDTDLnk8XNGIM/jpY4sNMUKu+5hss
DyzhtVY6hmXZQLKwkcl3ZTbt6rChCmqsUik0xfqusgsWf6i4Ah3JcGABULsADfoe
tAz/Q6BlFP3Ja18dy8V6SCXTwCQuc6B8TAvQb9zxQhr7ddUcZvg8kwVxSTINwgLe
XtBS1Uivy7et7POYCpOrIj98xNlxvX9rHi5ky05r3Y+eklqH/EJD4obEslUnxOeH
59099nXbCVsSg0aJvwgxjAU9fH52mvEsmLkdKxaFe96SG2qieii8QejljCHSg0wU
WLxUB6Ap7KnLSik24llq/DWr9Yh1YGemhesvO+pwWPC/a/l+E4iPnwHIT3TXJcyO
PBtIGPXQ0xbi1aLOjUzKwqFy6NarIrIAdbM7S/uVaU6zZ3LcxGHgimMNRye5DDxQ
S5qqsYv24BBucxFv5GR/yGcqq8RWYZ6//JaT7/qv83f/X6VzdZdEioJqRfEE3SyC
hJ9iHzTuSmWVH8sZBzwgYXfff4dvLhNGLoj2e+O0zJB/dsuvW1WnCQflEVxT6aXp
nhtYqlGyCsLRqvF5BbcRT4NDcc6Thbh7RPGEizwk6nsRePG5r2Nl1/GWThJ2hYFl
Y1K54ktZFH0T0oFDoTesK+lw4c3B/WOtqKmKW90Kcgbmu2yYiQP+3U9cZl8hy1+I
gpflg2fnMv6fOW4rPxuC1YbkxsY55Vcs2QXeQRr1EmdNGGR5FUKzi/U41n+5NDp4
J4H36XpcfJS0mk7kYqp0BT5juVXQjqN69LKdK90ddQYQ50wpmQfdUst/toiXziNI
0NGqhnKWIB+8fG7LUylFGa6/ft8bvWGbgzHsmxHJnjfcTyruUVSR0O6xOsapIzXO
Zv0iT6qc+qrRC3QB+9MsGmhTsPMcdI1OwLrjkr0FzIWl6YAPct0THWS3Hyp5wecC
iuSp7jdyRBOEQ5UsVWINUCE8fZVUpfOdSUQt6bKZA2AsaFzQ0vPv0h5ETU5gGPmf
kPF4qaaWvmwUMrLq5GVHLp66Q67gG8iYrEqWl32TB7HXuOz9jUjTVtCEHtNkIHB7
Gf3b0WDkza3DvKv3ns7M5R5pCVEf/28OJ3hdEHlp4UyiiJ//4Vi3QcUeDWlpravZ
3HDG1YGa5FzJlTBHQbIDjGh2O3iNmscKplAUBiUhbnyYZ52vM0ZJzHXn6cx5Ix5k
VyEqD/1BlNmpiVpCWZwvVLtuJiWKX2GiQzwY2lNUxCNhBKjFJvPNBkmnoaqR+aVv
yQw8fPCigBiUKSUrECQxTQvQ2oxTnH0AF/HEZwvP2t/ZmGJtb1WBdkI24CjgXngm
0sSgant0eI2PdA17laFQ/1hQIsvitLHbJivOu4cajZiD95WJARBdooN1OPZYZsva
0zJVw3A0NxvWFkYlRyxLZO8pG8xvjPJldLvmFBR/EQu59swmkKXgHwqTGTogacAv
krajFVgNiVOfWDDzQRfkVEkGBGAEApOLYqoHcQb7EmEbo0HwyUAlm1xvradoRGV6
aUr8WVUHOltZ12woR7ZU6O9CnxZnd/RrVIZw/vXVq+gzdX+eAnGV5YduTZn/4v04
EWUsqL5rt2XywYbtvQsQJBw2bx44o57c+HfoJs+Sp/Ywzjk2wDNdjiqz8HMu2n7x
t5PXyi8hYRlAoxDCU6ql/ksNPw27d0B8WWB6N7Ho/9U7TUNZgnGOucsDj0KVrNv7
GafKv7s1ojk+5AA/xMGhwMpJMz626nK37FM23ejtvcXZEqRzodVdDhaMAAa5DlRO
F5HFoG1Q7dB3r2usLEWZSqzFtH84xhyBTBoFRZHh+CONGJmzB8rABejmwkvp+STJ
KVihl8Jx+TWTN/UK0RPmTdBp74yfuJz0GT8SxpMvmjz6Jw7kasbxeowYXZYQhXdS
+9FW59FwhKE6xumbApo1MrB3qTv6duahk7jCP2GxwXi9c+xESsiE/15u9253QxRn
fensRUrLGfoyuNuQ0JR8/wYu28pvxTRpVPTVQsZr1xKLRBTUbi+01Dg1lFKTl3Iu
EWlFVyLPz39spxH9ca3WZhhcJZW2+Yg/UUa3PUbNQtpGETTIeo2PrAq+CaMZE/Ff
I/jRrE8ytCY9S4WG+eFqa2HrMjISGbXombjmp72HCWoNEyb/o+VRaFNjCMe/tJcM
7YzwLBfftR67JgZq9V1Z9me1ImAb0o/tzS0f4GgTYLYGMDEMfRrc/NjntschubVw
c8lyYCVJE3OCLq+7TDp6tahkxf1wp9MnE0JWKwE0U/2YmXwpqKTaptgE2Yk4HfCZ
j2GhcQXK6vlLp0X5MzjtUOV2SgQAL0Jkyst+mPRQEYcSvn/etOH0D7PwmDd53H96
Bz8IkNMBiVRXarLJaleU0U1eqWRFY7pketyRC7RPefWSqLr9i9FqHHW2tuDs50dH
EKguL03t6jlsAtDiyh/qcW9eCBDg3qrJCl+CZBnOHrS1PrYE0OlqQ4+eT00wIj90
HPv9305fPsyXL/rpWmD+6kR4a3RbuJc1EbJ90C4IXkLonIMivAu0eSe3+FitK9iW
EYurg4jdvJl+2eV55ZRXstKPaK8jkvk+ydCe2fKqqx8m3UQT4x4KgbVigc5eIVL3
DjSsbXkIitzvmHzpcCFEpTdEcmK/RJXWaI92q2AX0apq479QCP3g8easN2V3tpWh
bNLTX8Dgu3Sk3X2RCqe7r91BKIhZMwuyrlSWn7LyJr/hHUulkvDoaNboU+loJWXW
JCKaIH/3M/yRxeSs6g/g8DiBl5tvi78GgyRTO77vFBdqXmsSFPW6SoZ1+QbiLu4U
Dfgfz1fp53u+Qz43xVOCvS+J2ProeOmYo++szQvOVqclr3KVQ59yGzljJB2Aj5N+
QznkYQqydbk5+Dx1RvxRkF1YeM1GrNR4gCoxcpFOa6yPCgQgtZ+9MSO8SQ5zu5n1
n7+boUqXx4xsuZCi+oFLfYn5uhucKjv6LDsUsELBbLl8grZ82KJ+223ScU3AZRNC
ps1VrjrI+XgCgk8IF2hPsQ9/lG3gQzlpsKQv2fuZ1yLfrB+bIH7e50N2sz/ewJbz
qL6agysSKXrBaHEq0uWCS36WDjP59tfwINSc6H/hcBrXoDYDzr8yj09cvK254ey1
ObvXjaeSv6M9Pz2n3v3xlL/i7ELmTb1mfEZRf9wT77iTqmIJb4w1LmNbDWFA9QTZ
iYXwbzLYofHdoggXT8SBXf5FFUFkOs6zKAvu6HY+r5NUlXkaRvV3GPTsT9g2PUjg
oHNch2c3ifUB8KVBS7PiTXzPy+NU/Agdw7nYI7szek4S94tkRetB/M7qPL2xma4T
ZCnbI8OSVoZgln9t6lzGVRhSUUtu/kiPO5RHcuPMV7OKNcIDtIwt6Nw+onvZEJSP
kUNjnPKJB35lI1JJcdaqX2GWS1dDRMSBU6hQDlP3ABaEIVKGe2bx0xjRnJChoAo3
rYyRTEKkQpEJOZcmbBF6Y+/a94qATqm7tmWsECgf4EQdZCMvlsm79GHyxm30T8pj
9mu0OiB4pjvunZfMNe0FyQcVtRbNBvZapHh7uYcZDbVXb8fvac3cWytlnGcdeW3H
+T4QsEvC4ajKyNv6dRn2E/oIMPhhraGUJYHO6JPw8f/8mrq40i+nJyKsrzFUFD8u
x3hoa8GM0IPRnnhfzpguJQU6z7lXp9a+cL2ljkmqiZo+5f2/MKHESWdnFkuR4Qvk
rKxmIV+yiZrHZkCQKcKMbCV4t6vlFbLtkjCqNcp9oGJiO74PWehb33L9EcTLzisL
KH+lM6J4cjUQcEFxWoFDAzTGf15BsvhstjMi9TsaL5Uu8PDtxjBuYZYeaiLolu4t
f2JcpdWeDBN3UyJqbtzrU7CnzIfhPqCcXwrKQfIiBfGfnjgUhYUiM/Uuifebp6Rg
xTuDJ6zUg5A7trG+aGMTpS2vdtx7Pl9S9xLoYMFvICBH50OogSHM7iEX3pmh97UI
az0LD98uB0JG0pRHTHsimQSGOStdiQjZVwceoYVGR6h0PMlgFuKTiCwtow9dou6I
+/tgeM5BXKdbQ0VXYvZgia9cJ5j7Ql8XAOPUwpY68h+/3EP/2DT6QQIUa07yzeAZ
uXDqpIyANysa9Ja040LO4eP+kBrcBcKN0t0MQhiJTVWiHG2fM3bR4zpnVpO9z4dr
KL7Od6KHGM3drc3jiQlNCvq0H57dmlG69u7XMW0eHt4Qwbk8RSRUr4eL0YacINYn
0CGsWuFdM3bH2qE/U73fHolkm3p4h3ityQdh+oFRR5Bo0ag9MNaXGNMb/g7/XPF4
R7OZ3qEYIePfewNYr8j07s/BSbzKtTVgHK2+418HDzi2KOP/sVC2IlY5vZwlQfkm
g0BG79daM+xGpvnxptqLULrPsBTUV6MkLEsPkbkCe9jQx7SzZtwBnkfR6YLp4UkV
Njo/iF3RZu4f36ZNMkv/fcEW/NwYFsUqnNCeeOqWqEzp7QtZChN98GD1+au8lFIk
pNQl5PXm1zIxD724nETfiHFp2C3TqooC86Cms5r3FGOhj9q/1ODkZs0dijtkJorm
Et8ANUFFKue9lLfnQs4VD0Fe3i4Vm4hlyOiUdVN4cTQ6cF6YkXdlBN2az1Ws8G7P
vH1NjVz+JIsiMAyvysa0etJL9VRdSIEFBShG/0L15hbkZM1/SXEKRS0WdTpce5KC
VivOyA8pEHgjjkQ6VVDXqp++ndOw99HZL7dHr2oEGgiU9mVJp2eUDL9ahghpGtAp
Ya1AQdxiyDlXugCJq8We1uqyt3iLpQrlH/h9m7sRsQh5eUngiP/9OzF63EdBfvol
Vpke2CsGGW96cGBnfNNUXxuwa1JUg+2L8KD0ADzcRSiyxx97LMCFQBmpbmmcbBlq
hgEMGRERlIU/bq74x/OTiG1blL5kp0o7XKhPpD88bf5L17tG/RbxVl9S9Ho4US0/
1wxOkSmvFTA6hqDcU6FlLC3imAXdV6OZIGUXCWYb2hx/o5xBHJ4/9cIo5dJnaxY3
sTr6nWkv97Yk1JNrw8x0FXnMEVq4whjCRXcVmrnidrtTTW7adiUJawNUnAnfEMyd
0GHtnKXZyVZbH3fo/LzuxXzxiG06F5ItfZ2s1c2ZOTDK17CYXWOZXPiOhGXeacLO
HinH1IBqHUs1nHes0vRf0+zPyAKgGfG7yIjw+cnhELjjHIM1TVUzXXxkKXnF2vtR
bx5rbTN2rdj4RFlcC9RrSGNvBx0YeqRbGs3MCxlnxCteJ3FOnTiE8zbcFmc+vQ3k
4A+DYWXrkn1eCrxSfuMAJxADQ9WKYOhslCaLgZS3pggTEV0U5TOGwJRWt1kMdvYx
/S4NTuw0rsb7UOVCXDT6NHwmV4H5zj7kzvXCE5Prkgb9xru+T4CcF/j3QhtMLkSh
dw1+LtCKdmw45+C9fMeIibY6QEnAjw23947tWDkKTeqyDZY+HTeisaONMAqLyDfY
++FhH/UVp3O7Y6DuA0/ULefqMOE/ML9zXS2sfsCsJAIu+hcBUFTvErB5yA3JMExd
FVpINw9B/TMtnMBrVWCA5a61cuzAnAN/fsG1Cwb5e03fnfTg1RSngR67nB51o4v9
iNMktx/7pnQpK0lgvOi99VPNO3iqgYLMbwKlRV/WhXCl7NtXYRfbay4NvKKwxeGJ
ITvwn35vpW0WYrrWi0gTVlPgraEJeMeKqvDuDYS+OQATEO1NeVZcUIh71sis9TrS
D5p14ULALFrN14KCkCMm86qtCUpZOGHwa4X62TLlCuxYuk7tUHICgEk1/suG4Ucy
p0U8A52/yNkVHl3a98rQhng+a1XLF1fe71py+rV9Ae17R2qM8Q044VC+0vUqY0U1
Bszl5ZzrB0+Zd6eANQAtUmC6ft97wB2PyRFNc2ngeQ8OCLsdtpKhB7fQuZpc+Kgf
jqI+uzrbcrMWqGd9q+Xz2zon2dxYyXHh6JVu9R+qk8UaeOFxX8KygLCmSijAfURR
poE6lGidF/mOYIeZmQOd+23d7572tsLd1A3FVRhX4MUtUlJgODosTs9C/lX4noO8
0Y7Jq0dvdp8U+4Yx6A1uVjl8sVLRqJLmSz/4gLrMTyD3PI3XPlVR2filjAEZvDyy
XA6Jr3LWSNYI/0hG4uJpXt/6lV6Cqn6TJ5VU3NgGV2wL3CUlzuSOEDeICpoMSXxD
bOv5qz3Ok8JZqwtocD9R4zaIC9wA28GVO/vfJ5y3730TJFB3mwSxX1+Kivz3WGR7
FMSMQwlmHWO9b59FRKiA36Qzq0DKCf5E9xZ/Yx1298nscVQZvWa3NfXTAcA/8bwc
n4F/156U2g/iyb1MOwzkcXqPo9JfAg83gg0OLTzZSSrbymffHSMockU4ZduH3Oac
v+fWOyhHmCGvBb6yz3ztD8Gd3pjjcHoLYZZStHvHWMSx4SxZR4EPQmlfJYoHKEAs
0iflyFbT7QChNbPW89czTT+QLdBd61mBC4z0qw2r//PlJqbKEQNk9K6jWBPqpSEq
RswHN7hlUuuc9f+vqBWr1T6qm8XXVjjyS6tIgL9uyw3guTkMLd/UfL8+7D+SYlYQ
UmDbS4Ab0H/XNn53BX6XBGbbCBb7VWbqy6L9YIpCqDUekUt8SSEqYqs88PN4po4C
zPWLSDNTZNa9E+pkwuUjMngGmy4NFvRKAyVpw7/li2S5QtcBP1SaztwRh52m+pGs
y3Q23HGsnlYOwWYfH/EIVfYPthK/MZVbzSoPQghn7SksNfYJXvUNTaCQyGHad0fb
uDA1AAmIlEKaVvvwlRQnwIh3ff7mkVIJBASdR9cqFGpZwV2AMLnWfSTav9bhSQKQ
Fxuz2zMaHVmi/8iF4M/WsfpfS4R9clglqos3zIKklcmcwRjZRLTA5J6p+FV5G1OP
qRNea0cUVJ/MIPO7dUHmYnergvU3k0BIFUn4J3PjcaEppnlX61bdy6/gr6DfyZ+B
wG7SCEWRm/6LiXsQfvgfZF6OQYoAg8ixUCfI6lA9KdI9PGznIGuRPAwUIkoZgYNX
dKcIHss6UdojBhsJDHx5+rO335E7DJ+/LT9UILHo5D/fEgy2D636WS4Qa/Hz0kmG
kRc1jO6CtEKvS/qJdFsH0ijxCTS3UpzW08K6g5K14YWTOVlizvs0qKKoqJSHOJLq
WWZ2cIu+txZsP0EFT3ZQ3vx6WIXySwZW7FcRU/ZnNwKQ8uaNP1SQwLJ/6LnhKTjX
6PI32uMvJtz13QYo5vdpkKFGmREIOsz3xWL74I0kpeYcVRcx/Err2u8eep1dNq+W
chwAjuobFw1Q9oO1poRTxDp5nqJlDDLvyByMkjPwyQU8X1joDxWDrBivzARhtJWB
XYgDZPBWj2yxpR9jEogQUzV2HrVGj6oEuwqPJoNeuiveL/lmosMeb05Z00tHXHeN
wLvLwXTpc/lepC8Ca8E+SeDsn6jhys4K0tR6BRZX2csAr6/iOnP4hx746bPoXP24
qPh+086LsFNWJDoVLDaRW73dWgGW6PA48S4avrTnqi5odLpfy4shzLveWAHxEwVh
IXyIHLPewPICEecukPnnHakNcf2peQ9JJihaM7eWoFw9JjxdF4hFpIsLNmloYZt0
4RfHu2x6mSoIhGsEe8MnbBPYJZ3lvhUsb1+kk95dZbmzDfd7eEsA4JZKawtJequK
2DaTzwBjSXVklFdY2BUTOrB3cUqOq53Tfv+PElYcfzT67UqDnm5OPqchJ69cfZdj
JPqYOkVeJRCLYNC24v15+RCK2xuheAchc7dcG62TppwEO8ckybF7klpZSv1uFmQO
a5bj1cj90OCUME4PQpayTBgo2L2r/AY5Hpjn4F60tbJlutSO68wCFdJUHKZ6EdxQ
8BEqcU/ytQdOnkDT5BEbZegqwNtUURpTl9e7+OWcO0E7Tk5IeEnRmH0YMaBpa3uv
TjDW0X8xTI81d2+jIu2oLUVZmxQxxtCc4+2z8zMnPnE7bIu40TN+14jfiNDiwRp8
xOxQqT+Pl/vjHqbLEyaq3JhzAFo6k9fxPWrit50fdFqdz0dnbrlTxW+kwXGhPgro
avIj2HuywPK2U+A+35S2gIal7zggOFp78oPSQtTAZWyqNFRFNllEcWgxOESpd6bK
rgHzQNUEz9AE0WWzFSzFuv7YjDI2Y5JgnQfH8llOKpxR4nPYkzfVlZfYoNzkcajD
r2X3oOP4h58KgHgH2PBeh2Kh7+YUlGY9eKHmOJmhgT6Joa/ANKeWOxLUf316WinS
6hXuHjzMMZQ6+FR4U+gNYPt0AZF/0mJ7ln+StseGARb7CTaXSzWFRWoliGL4//x3
2aJlbYgyWuI+bXzxzvabAB4fupsoSI5qCgUIZVxWnWJDZT6XmbBeS479Vkg/glgj
ciCaz8EyTSNLjCy9Zgs3HDTyBtM3FODGkFh2FEQB03r5t+1cZ5IBmWr3wt7QOMIS
CZZFRo5PMU3Yf2S503U/2xVGtYoiWUE8lDREXCIuT9ZPCgCk3zX10XEerH6t3Btg
m8zc9nnDmloFCBrZpLN0ODk6EuOzbRTZVLEnWBBlF6BmqaiVj/9H9Ja8Hwhn3QL7
Xu025lJfj3OeB9q+X4qLDx2cHd1bkYPkyAN2DFtvgPa9SG0vvOb0Pzma+Jb0IeiI
Szo7GDWVDwWRzHRBvGsrqzhVpt2LT2saub93tTLZOcjfDsoBdLYWVCQVyLCXfwW0
Cd7MX3ca1dPsplE3tFGtCk9HLHN7rrLUrYB5MNTMvmVExOezwyl5vxY6+AL/XJKL
10oZaZqivDh0J/v9ulElKrrAaxUxtzfoQ+SbItN8KoSIkE70xBR++j50jLoZVlDx
j583Lh96gi+BTjOLuGZ6hIOmBIpMA6PKZ0iL0oIqnKCiFYYXcQ4/DxevvV1O1QJk
nH4bIApCBJBF8BAlG/8S31fx535ML/iyLOoKe3v+HqhmLeZyddiuhRC+DtEucp8t
9NrOfqTJ1OtuPXE2l4I/RxmfJBdl4HzwwJp7FBNTSgqOLWeN+XxJ9y5qwToHPV+r
Au1jQMqeootAbWOKOmch6FbZjlra61XXbszjYCAXRafjTPKAyFv5hGjaE4iWLgYH
Bu0u1Dh/8hrMUEphPKPkOX/gyF1MYofe3Kf1gEKkqmqasGPBb2qFMKFS7/EXLk8k
q9cDhqxjzl8gQWkjEg4LBsZv3l0s8Qehh6b6eohHYTdQpWGlJEoBrOtx6TRS6kjA
MryGivkCjAByCFh9vJ/XK4ndTgBdi2qCY15GNpUTL7PJMPJD5Nb/JLhCNNCHIMgn
lyNY/RGx+C5M46i+M+oQobzwX/eBaCDl4J+Cp9TzQ9dWygB9OhvWJeKw1HIwTIn7
BphLV3PeZcSd7hjwWxdHzK6pSThKzCdQ3lT6FOfeTwEFOQ9U2PpExz8pdR4Xgiz+
GJHWbNVnf/icFTDkHzRFWajNXgj+zoQrI0wDP9hdY1fGG7r5dwHi3Slq72AjNXHj
PVDD5bKfblanMrK2NOeMz0dU0rIML6TCwILCu/FoZoDnOBzi0QPLTIEB1iBpMxDv
5MhPPgVp+LzjlceJeWGcdUge3mY2EYEiiGzvjeodWxjcuIVc+iVAMwwP3kLnUsPM
oRLSIWfoiscQr3RPH8AwVoip9/NMGIYkLNiXTfSq4hNY3LSt/BUzASMP3LTygl6j
447oqxOrc/W/mI0Uu0EtWEnVrADP8llzntU5rLxNi3m9FMGemwtjITQxVL2Dm17S
f7DuX70JxDj6Ey7+aKu2odALgRGlFdM9pKXOeR/HQd6D1oUwl/9+e+FznGfvxg9M
f24eu04v+U8XpoBr1cci8A4YcQdDxwBqnNA7WUWC65r5+37Tv8LPz7p42TUr8JlE
xlGDIervMgW7LRR1URiy4h3sbXIzkN8OMh9LXGof2IBA5lXMGlgG6IIffYb2YzyG
9fGzDsUYQFLmObtRLPI9Pwjsja1+f6q+Z9nEi68O31ZAEB/IAyFSrs/UIp+iAa4l
az75+gXWTYGX5Xl7KU3EC73AuqdpwA7LZo3ip0BFRtz3gmsmwLlKaG9R97C8jH5G
+GtOAW54raZxWotR5iPYvQOzE9tw68cvrSgaGHgB47Hkhwo3D1t05P1tc9pD+p4i
k7GldpM+zkyhtKVpHsZG+aL1dXwnIp7fjtlxwewQdNWLHzBnPvkIg3CLxuFOZvUD
EnS9yGKaHSz7IJnWHKx7RxeVmZnS7yc8653u5jeNBdJm7aCeZwMOE4ebaH5Sjmcj
uojRZuUBE/yULTxQE8W4cpiKrVak+IFTUwn62dcLF4bIi3CHDKJbswwQdE+O9Jvv
/DEPqCi+HeX9i526VF2hG4gFeRNy1ow2hzu69wcrNkD+woQzeAb20akS9CAbMKBv
uo0Akqv/6RbNs7AZua28s8t4aLKGxDi/03mySQhf0rk9J3RLdxZcuxKpdgdWTEFv
LibvzQFWmBWma466rxRoh/GVIjqqcqmg2n4uHMACS/bicEGMLNeU/aHgZtdydgxl
5WGIiYtTg8ikZySacMrSiamWkDZmrdhFE7Raztp9jcp002MqWeR1Ot8+Nvlskc7y
F4QTzexSm26qVjzEQaAPFpJawF2OqXKiOvil7vnrFvJtY2EeklUjgO51lWzmhwL+
0TCb8xppmWM1tQvxm7Uygh/vEhjD2XuEUC7pQmjh+ylGf3IXRZF7+h++bd4hySFQ
mB/g4GCM8w6uyeQjG+kJeAxMAGXhrAUDJ64xxko24KfO6j9mW2fYHfR38IGkWM+7
9lUPo4vIHBF1v2cm/bqjFFI5V1/aNd72eLKlJpLyvsh1WTSfuFbDwN725gODQvI7
ySihre7SIcqIfqfomva+EG1nawoZr6tkxnuV/ujQ8r/7l7UnnEfz1VVOska0abBA
8QfJDVuSziHUJ7e0hXoGUyMy+yXV0dxvAWamAo/v1ohyRsVc/BXnGFBscnd5fBfk
3gZTRet2lDe5yZEJLfS+I1phkiBxdnsLaa//1k2Xmert3z6ZeZ0TFAmuii1yTPPh
V94cEsDh1/M4PZcRcpl8QHa3WI4vt8w8i8LBqPQbjZgYMEYQ7lRBoS3ejgk9DFk2
pZe7Q1IyRr+p7NGqK4qDudjDaJqSHxXKIfpXz2Q8zR2YKXAr9md4DdvJEH3CuUU6
shEBJ3/F1LVe0D5iW8NTZCNdyxU8O1h7ftP/9JKfk06h7it/7U6bal1xU5Fw3LkS
7iQRhvjrebHjXMvDCZZy7yL6w3k4ymGrdJQXtZbXatXrRvfFwgXNW9zE2az2aHXp
rVZQIp+vcnST3H6m3b209XQWHM6nhqAVWw2w0jSKJFJU0sYpUUM0T/S+8bJhtqf1
j0m74umZtyTR9zuD45cmkehRiu8Kw9yDL7oDm06nxk5gRMylNkqqRFDbEX/8H4bA
toc3Sa/UVUAnu2Lx++VbmV0hgHo7ZXGsT/w5PAEeMN+NucczOjgWOkx+WqKFqxOC
kiq5GcKVDWmZNvD1MejSNUR/39FZ13n65YbqXIAzlpb2afOnrRKolPr0SIcXae0A
fsk40ob8aW2g2bX09jHwOzq5CtNKISmwwbvIOPsKxIRCB8J0yz1ZzAOQSLBDd5VA
SbbbCDEiUKkQ7TgfFIBgSVs+4h49Bal8vouhGqNapPMjx0X1hR4kFLM8n9A106BW
Pcjv0mZvWwZKPxJdEo1RhZrfHlEeJNNi8hYt7N+Lx2h4BOSrGFM/hBIINGJYEPs7
biW6ZMKYvCU/j/rfRr7nfyNIOz/MziQbUANLOAwoBFqNSXPFfGgKy8JlNSGATOlz
juR9uNcOIbFEY2xJpPKnPQ/QSggzUs8Szg6acfYKAg1qHvSyLxYA++8WgOWcBhDK
CLcX/lN557UcNTS9aGqKnhUDBy/O+FwGbb1Px61Lg1HjSpqKtzCIeLMDIhKqsqSD
5kzjCPaQLkwJxuGnUiLuq53M7COh1tNlC/CCyiyJbpbMTclwWr7DkuGOloqx6YHZ
eWwWCzmftdU6lQ8NkFts7cHKbYMdklL1QQnSCRyi1UY/NsPEPozruplkmNa7M5nx
jTFZsuVlqLocvc4NdtAgYe3klkdErl1GAMPoV5ZCp+w0NReUWM9eAhQq1laY8lrq
beF2GZMQjq2uFK7tCHhb2y6bluHTP/UMjAPsThuclmL/T9VyqRpOAGXyBBXJmIOE
ky4ppAfURbsEcNx1Ezo7Qgtl5oCj26RJIaxZyWqPNuso0cVEUXmxu3NJPyiadof2
WXpxhTAyQUJsf+xgIqLAwDb0ibQMErAB+AxUfmovuEhT1BOW/VnSJhh5blowGZ9z
SHwFxl7pFVxLlx8K9AUB9jMwDsQsWMuiKuw4d9V1RwNCUsta5IW2oecjDspyc5I7
+jzI3yja+2DUynuRJ6/kmral4RXAkXmJGkCDuhe3GVMeiUDDfGrUdriUMmead+74
5FuJtsNtvTVwskO01t/NH9fgwDXxSRWKZ9bCLE0N0evuvU09yXZopJNZ5i1zcXiM
Fh/rCpKbq/mre7mweXlTZvhPIhZCiClvA223Phy5A+jO1Qzb+PN1lmFq3TuqllaL
ohWSQnyqkHmUblvR9mYeRMbCSbXByr9JFlS4e6eaUyKrI5UmQn8lIGt3wXWvsMDy
vVWMSA6Z+76t4ZhYTfC2bSnHPUJ8xGQbArbKhPYPp2XsDBmAckUsSK1ixty9QJKf
x14ZywQ9EPlriO4HuLSllrV7XXdDS6MteigZy5ajaIBLFwyXJN+MSfWeggiMjPW5
MWmKEKDXv/enps7gmBzhmzCGOKf85OlzPOJ6f8f+ljOoeqCSLKuSkfcsu4k5t68H
8bZyVupOI+W/R+rREq6/aGiLYDUqrwYDcFFN94XfAlaWkC5AhO4zmRr/Cd5H+wfY
RFZVg50/dR2WIggOWubvnYkQ4bWq+CaevAZWLqKiLlCy//oNcHcYVlkEdRySdJkH
NfpAZc9GYfEnSTdWHGE7sAhR4jk1FA+UwDhbmTPmf2iLwS6eNUcdDVC5w8Svq8Ab
50jBn9uAbV84HuXCUiRIMX7sHr4aCgDxuAjn0dQnbsShRxHQOExBNyGjUG8ybc+P
AaPL2WZ59GNKw3Qv+X1N4d5uy9rNuOhLpXHQYauamINVUgWacUZn3zG0+xv918iu
4homWy30ziPleYtrowsA5ShYrnF2/GFisWg18IuMLWEV2ute7rcxfcBoNR7xn8WF
0o01ZDg9K+U6V7z8rMndtteGLbQEKIsWa9hCDyVeKBPU4757oOJTKh2P8zuI8pba
CCaTLodbllB8DNZZB0HdW40dn+KbYe5RMZ73WntcY470ss3vJRrBYY1qELg5xrSr
2zKlQv8HQ9kKsHGGtbiMqQFSAjoTmvcDlwAk7ButSOmE21JgeFqt56JzQinnXKia
CObQ1fS01mT2OiP1kW6LxR6wQHtBuy7dD4z+8PUx4SUF0I07XnHCYXPiWKoyfoGt
TqX75WgI9FKvEu4ZrEi6OciyCW8//wiVL3Y1jdEaSWUGZmUYojHhJCRXn/6LKvGg
tEyesFUKxD3i0hEB90LeW/occ4AItg1w5vkUKGy4yeuThodcr/2JWmxsA6fF8uIy
ilWXQcs2a0glYtZ/EdQomNy25Z9GOv1y/FTYDkmAnjFmrNe0h+vqAJobvpBDDpRU
L8LKbcXpxnTauDmbBk6vQbizyu2V4MmJffIDA7/D3X9NJ2dsg1fMY+GJd/2+Kh7l
8e5otgyDh4vi10rksGsz0HB1a9l5jJ9VPTqyFge6ebeI78sCGLPzougkbbEgVKR0
iqFcASYOtoMKcN7AGZyRChAc3vXQSeXppg9lIAUIrA78GGUZYpnpjfK8/I+6FMVU
tlin47trzN47Ik6tfF+ReZMLYSeWr+SiRDGqWj6OCd03kY5OdGj7PgjGvGryz36Y
V5xD3FUHe0S0rNJywMJCdcRhuDSVpR30/ekwCjryKR7i7H8gzp+kDwxAPw2sYL3y
TUAfk+0lyfmASwJNUOpKS2JiXTJHDf1fRFd16tcHAiYrUrEILDG6A3wU2fvSZFgx
q6i9bdCsDZlL4iAx5BYCCTeWwPS1m74GHV3MZ0/t4e1F4o85Pbl5JaSTwOrDwZZq
qC3QQqlqkj1X7IsPAFHC3yGpQlxknYkwzmH8wyF3cLPsZZ/jluTeyTaUUxq9ZTw9
45d8SeGSKfwzqJKrbvxrl4VJbhMTFIxYOTc6CVFhWmQQUzl2MtvuOEj4+RLmGa9n
0FiRkvozuHQD/mYyd5dz7wKAkcr+/BTGMR9FK2VNIdKBWA1mBCAz1FZoHAohEmoH
Sdb+koW+HAZoOdUTyHCJ95/2ks1J6t46V6Pvd/2qGwgvQWsjnglVgTPVm+iujPWg
MdOSb0SQHK7+7uimFpWUZAwj2a34aMGedIuCiuVGL6n1M8LJc0xydAPL5lTorfzW
hFOnm0Fx5jKrNp7KwpEYYbeqUWQ0GpSO3tyijjgAx4JZZn33QfUjN90BzLWwP3Rb
bzYNIUnTr2aye4wAF7FNJia1fRvw0vNEK6eKrtW+Vk2dDV5zJ5WdkCxml6OM8xYS
cro0Vbavji6VOofXGoRN2/odIku2DcVMsUP9ScupYeiFiJ8WPVD5epxPaRVE3L0g
lHsu9W5FsBfU2AmYfdZYZERE2qHxU7LJAbbEnxKVnHcU5m8ilxya08oZsxMxwH2h
SWTGb0YFrxJ0Diqcfa15Jsi9jP43enm4P+5KRDAGWXjHsjq+ajjpQxSWc38ElcU7
/rgnNbzo49PZU4OGnhHFkpoAs86jlZsDdKSAe6nMgIyfk+WgqyoMhL7ZbJUp8JZu
YqjzdpKwRGfhfkx0Pm1+dEt2lOb2YNoYrTlE/dGvoXClhQOhParWzWnHPsX403Oj
7WQR7p60cXouxJCCwzocT64SLRjDR/oW0W0DNNX08o1ywvKGisfetAI6inxrXNGB
U7rRKG3iQXQAdNP6yQ4hXQHD8Tw31jE3YSOVVAe3YyGTYCynAZ399uHNs95lTj+v
vRa4+I231lXI4/XyPXMLkbITBKqni30PkjeFwitOVoUP8jqPOfYikFUEqHkpJVeT
GqT34pLoXVelOvA7Xt7CrmsDfCncmo5RZUOeMfOBF+/xB2dp8ck3o1rYUJuy3k2N
V0+r6m1zKKCVCAFJsC/1GalTqIreB6Z6sE6c985S3a9rbE/FXTS5jLlwrYMqn7eR
IHNoiIPnSCcDjJaz3pUFWLKq3abbDvrY11wTIdPtEPgiV/0ym3zMc25l5i+88BK0
ctIXmejy07A8GaiCzgEYwJ3nxzdfILf5zeN5D6ox9qEiLUwCwSmYmtW/OxRtyErx
WnO3fa7AgqsignP+0forYkKIe2jwDqYBEvSzETdMn9i0VpmkhXT1UC6CLoX9ZHTg
3oC2BVPWvOEjYhluORc+cENZY8FjLscixFef1sahnCuG/8e136bKRsTI1VOVv9DE
L+TkGEI0M1xJZ4k6wUpMlu2+6ErBaqKhIhqMmziMjWI5FOMKWvgnksJlruPZGRog
q1GoTsLa1Vp2kyzJ8vxVIf5OXWzXvMAUd403SUxziMPI97zQODEmzLgg3C3KAEnk
tU5iOoYjpqrSLFfsQS7brrAWyBwF14X2k0tBvo+x78EQ9uiz5A+WsvBOQjZMYMDT
L4j4nICguwQT8x1pMQY7dgRBWFPLv0mD8hZq1x+BPP1aXAz/2Me+ojAyaGRZwLQs
6LP0wW33JvNciONE4SbKxnPtmmGphAJAuZNHCaFeE0A5IWcZszU/zPJ/yAx74o0T
9rtCSAIAaccMc/1bWLTOOlfU5YOVe7jG73lBzgka/u2zsNlApDUDVuLndXazj8Xd
miryK/PXCLOLAs6pJ3DP7qmee9r54+cF/gGsG4tJz7qSSB6CJdIc2O8t80a/3zWU
qrAP5HRRmvWgNKJMlt6iN19f4lwkg/qbmOaf6Afe8/YloPGrmQhSW1OXTI4NeGKC
TH0dwPSrGI4yIJK7dnhQz+pZu8jv1zy1ncfp0feK4GmUAKtvPFqwBGJeyuYmNFrw
sTqX68pO4zeYUk2j3wDSMWhTGGXzOXJtHh+iFhxDFxhQKE7udPjkt018fiYmPNVo
kRnowUnbPkh8i7yLON64skVsgEaqnGrGcHnHwoBToAbvkMWtaOEVO55d2Ef94HUE
R770hmsSmqrGjG/yLc4ymFwhh6t3CDQczhN0Fiqb7TM8cz+NUUK2uG8VD1f1XRya
3CApHa1IYoOfqst2e8Z9vi4QDP5B9aSobhvmNUEE+Q36/mR2YjfCCvD6DxmQIu1q
/aTdAqg8EznMpcqKby2y9q63zUiUAbZAJKh9Yn2R9vTD9BP8vi7mONvm/elcSjpt
zbxlS55zPXDQN1blBdhUKImHw3twgVlTTVifl15yFOMB9QppVr8RLgz4eMaJSIna
fb/veoGv+s8gltxf17vjwpKrH+0jmYAhGdLgS8DesrXdHEAexSs4ats0ZsARlliY
lmLJHs8EGv4HvrmPi8i4HmJjy3gg1ZayKRCeR0sPFY8RLxk7mblgP5BPLRjaBqt9
QnOrxvpvl4glESS1vknhYj4d1biqJgXwy088CRB7h3v0TBtdV7aApLrbk1k80fhr
My91EKTNh/w9aXzV2MTyz8dyOdXHeIyNRq8EhwChaIyD/4H+bFA4ywkZBxto1e9I
l68G5xFX7rW3ZMDFisOfzWyG+ns6d7Ae+kws78vf6gx+jGcQV0xTBnQ6gLnk/YHX
OTMe/aGxY/20ep4sPbiBvoN14hqABR5j/cqeMfYgVK6cO+0mN3Exw/AqRSIKDL58
cUGVl3pIUFAJrGFSiUYeGcP3/iJFMiBLvNAx98zRVpWsddZqSfhGlCkPcIAx0/ZQ
n0AvgTpE634lA8B/oukSVy1Dwk/1DgT4bhCGjeuT0NtPXRLrwK9D1OFfPtXLTLxW
lx5+RQJcjcBujBKm0bwqse1mEYG5kvuC0SSMAd4O9IwQeFzYCciJfsZKBe7+fGSn
7HyQb9t7g3j2ct1UR16X793zj5UnFtYQeaMbH7sXDMtvMFTMgo956I+tMarnNMMH
BqqiZEQqhzYmfNAqhXuzSKbGPQDwIsLJ39h+SDTBtNTWBS+zDlNdRz1uLFz/JaRK
Y2fK0fTbttu/PUj9PkNU/jnxUrQYOclXZICDIosUqLT/P/8i06+GPwE+V3/kju1l
2/hQOmisGuQB2IXXnJ4ZAclXgQaKVAV+uGpeA3FJNT8bU+coc7bKGBQlTu9ha9jV
i7mF4nnOgvzYYLTjS/UEMu2K6jIwjCSWVA7GDvGavvVddaVGO0hsmftSUTvJHD+0
mDZJkTZob7QCIoNRwIzb535Pa/fH2PCURO/SJzRxpgbEGRxZtfQbOhaP2FupzpSd
6bMGJTfRf4mS85OSnAku3D4kuhnRyizEQZpFavF+cpwl2mkqD71lgP5dRexAGN4n
8leGyOyNXrZE237kViaasTXFzQUhCbvlsj50P9t/fgbi0bIlgTvZq6QvdUD1OMkH
NUOBGlHcqBs8gkw2nu+G1y5DWewjv5P2lXRUdnXpIrSRgrFTXfptDDeCvqdmeids
swlunp79yH22eG8DSbVhhMVDLrNTG52bA+0fgmajy/o3hwJdfdUnHapKu5DI6Anx
GMAwrtPdj8MAnzYktUFIIsIk7ubRVYFNU40bB3dNgIJtf3LI8NrOMt37nolsIA5t
a00KkEH5AdgNLzscVoLmGY6/EGMW/wAxSoVam0o37WafBWAvGKAZ1NTWpe1fF4cd
tWIsCSABKxaW2q5tFLnMtBhRU4YMxbyjtkgZKTXtcIYHc3sJTVS/VcFR/JmHS14n
d5SyHhrOMGYT9N4WNv5sL9Zwts20W4Nsfr9uj9kKNxdrN8NMwFzQWWuxwPx/mA+7
Xfw/6rTEweerNX7LC8WAHWuGbAOzkusmIptEAh4rztq4g4TsnE50KInH72qkOg22
IS80tpLaeHiMBbtmNXNZrQOq3oulVA7W24lEDMaROubWzsApG/295Df3kBkieLt3
biIelFORUS4o1llA2f/fxVrybuqZgt9hZy2hCwmaL2mCkJJDuGqRfoWUJsw0QtqM
2XhDAVOk8+ohvlWxKv+BdsvgDY+MBEOCqb/JdnOF4erjwDauCKyGuYJF+XDx63SF
rrbPta5S7HUrLQICDG5EvMglgjgbwku5PjKWt086t/vYq8L0Ozao62lB9MBBPRVB
f+Y4dr74s7sOBS3jvwIx50o+ZPhrw5mPjwkgUe+LITETc7Iqa82NfH/vXPk8LuaT
5srqT+dZhDvAFocYFl1DLLlhW7nKxFE/gQ4Qt0LHcbreIF12e0LsWDiHQYGIDOJN
dxqqIOYe0M5CBB2+hteX/OaLb+he9MvAaaNz1R52SCkh1hRQNRvYXzjvphy0eWgd
l1YV723MBaZ5OCvKMJwudZNWio9xMOyaWKKOn3mpxADEFTQVyyi6lAHiOg3Q4SHK
c9HGjk+f8wTk8lNgsFYThLVjK0XgIuBEEvsTxKVtc+md/Tz1clOCpoMwaxX1XJRn
maDbWLrNGgyjZhnCsYpzIR5vMcQetn75KIa18ymCjo4+mJv673zVuv1OWGW/TDQQ
/vHz29N7z2jftxo7wYptH5oCu16TTcEVZrWHZn1E6ZSL03rt2uR/gEjUapHSP39E
yglPqpjIJMjwpDaTKiiJqauxVcKobfPFhONaNHQ0ACp7o+/U6IlAF59s8IcpYG5k
8QHpM4U3uESWdBNr4comHa9LJpQx3B0gg64MG0sWpGOtwRb9HDB2yz/63YHCH6zH
EDZuzM6EkaJFVH+IsGg+tsZCUjQCP2xiF9lbx0VkE5y2o9iVpezll3QAjVVD7aXN
N05sNiDKBZW1i+mOrjeArnf7Ks3NYCo1+pZsOMa2AldR3GuYjwT1rDAktyBYChHS
BLikY1FLmWvRMseROAXj9S22VKgdsEHVlX6CuC0XXcxk2WhfqCqcIgDuxiX5GM+j
nGb9QEtUUgB5TU4y3ZTEhPg21u19Q3zbe7lxLewC2Bc64R4mez0sOeuUX7FNFpZ1
26tCNKqW9jesv2Ei755HNLl5fmZuP+qNXLb76Lg9znVm1QAE/FqzVRTEVuqrAAmS
DnDgol4HqcE4Wr054Z4QdDqJQkaPgs5pyh+8siU9zhiUiQaswcbGXgOQc0i6VJj1
EWuo98OFE8B7372e89eYAUCAINnK+nmvfaENqBlIyAQlRyGqTeQXdFjuAVAzNGj7
cD3diJu8e5oYcXacMPJDliM1TLDOvtqlxhxr+Gwth1HaUTU1lyxgTzblm2AQTZJT
+XCBTvg8EDcjDGvN718hr12uoie6Msy5g4/c2OyFiDUtniduudtBfc0VAJQBw1fh
pds1UV7T/P40QFKWv0ZNhJiBc/o9Z5qSronezhLDrq7RHiHagC8u8lKVdiaps7Yz
mPbFCD59IvuU9LnKlLAyJIZ3vfjQtpi27q72a/dw402zCJYk6y1PIj5jYScRKP4T
J5Lz70uW2HrDN0KdqTUJYxmH9uFu/KYgz9AEieJJ9x/ksarvQ0LLHZu+0so/zFBf
ED5IztV0PXv2WPYt75sYv1iZTL1FTLsBrC7RGZ194O+gYtGyNqPw2Xn4Xzbg8lUH
56EvwIjZAzlPnnTbnTZd6ci+Kcu29Ld0umjbcgG3K+69d0j2PQk6cjzAZwXVzCmY
/0LbxGlE5SuQxvy0o00m7n7Ptpu4RtUeUlHs9+JQb4r2TU8tBAOhchmeyviKpsV3
JlBX9P6/N8IoT6j3q2SIIx6pJkcnmuKYZl+oApCQIk5YQIzfUsUjcEHGtusZHkdm
ktFaEfXBz/r8CB7/gEokEYv9pPs5xzbmTS91pjFmn2zE4rBpC/mzTCpgl+j6DU/7
hy55gtGULiH2KLX0QIXFMD34V1uC1dzUzxDXn7aHOZIPY3jsmegaaa3mMj3y198H
F4i2kO3E8Ycf74AtSKaYf3VpU26/gageSb8QE044C+srJRl/B5bJfkDnjcVSrvkD
D/tCOCTY53XyFDXgWAhSh8jy3VTeHUMlHHhTrGHc/h1wiYgMmltavdl0Ej9MuXmi
CDqJNbLsW24kdWPvyHaCzm5v9CNEtKbmUYHjeaUUsmIZ5uuw1BF0c8bJRoe2BMl5
H9A03P5yneMKUuyEGUi33EQ4gLJ/5VCUIJrKV10UMPQ53233ZUM1sEEHfPLrIb5W
yti5P+oUpymoB/cVl72fNkBPC88sjeLsV56QexnkjHbgx2xEAr4L0bMP3yFNtzXE
ZDqMbAUQW0iEx4lrRPMUM0aA6gk0b+e+QcZyvXotMMuNioxcbBSWBIgMhABz6HH0
2KPMche3I9Lo0tSzt04qvHyMHJmm2FwKylY05BmgBNu19Cy96eAaOyAaSWKVLV3i
9jEuEMIm+Km0ICGclonA4/ATvoPt1D2C9/0KKNG95vFnb5Jmxy6KcxKnO2JlAO7c
DE73YOduWZvhzKsZSt3PETB0CfmeO7dt4TPEBNplZU4sQlJ1+BDUpD4PiqeHopEl
H9rKe4v5DrHV6xUyIk3szT5Zr2loci6e3kR9Bc8edDAz655T1bnVSxEwJGgDTHSY
4diGh/71sCOwI9Ns4pwOXe2hOvi2Tz6Pxp6IKEXGE1i5rxnyYV0i08MkXZaXTNsa
kASBtp9oGytzBP3fR/kf4Zmbi8G4b+RjpsW80kY+ZrQBvmFjhKvQ3O5JE6GJPMUX
pwNIc1zO/pNxWisw67qpxoXwTjeUjKoqsK3xy2APRQO7CYmLsXuMvdkl4SbPp8nV
S3vYXfjjIyl6pkax7GN5lrr3X1BkhuObtb+2nIROFmNkGMj2cAMPP2ifdHU8KdJl
WGU6qFBsPFCQq61bMMKymsLF1nD34u8n1HAHUJWGSg7gvSoKCXXZd0poV2pgLYwc
TceGCUOEXZw4CJsjU74XFXPHtCpIoKPKp3RiMQzQsEhqi1ZdKs6W2utzk47Z984a
Tt3gfHR12NYjWoDJJYVR4BCZUBtnO5yQzCNDZy5kLe2hK/rBYlj4rPtGCkYV8TNy
p0/q6SOqnr+vylWweUisWWT609yYB//8GuERamQni09dRf6YCMKpIwIstLdMNMVg
XoF3vT3RHMQWQp+CtO4Y89+VSCDpa75OFNdJE8Or3ux0vFNsx/qEPOnLZLKK2Iap
Oq/eXsinrR8ZzejGTIagT4oAI9ahthznBbpZcUxPnzl1v1VWYVUl55hwiBiivOcP
BhKz5e7tdEGI8If4dFcxMOXpzzOkBroB/1E0Fn5hgi1FKCFcebtIfxLQUgIJq4xg
VYt1I6I2Vb1WJho+6evmJPFwBjo2TqdGEHgdFq3lbjGGjgi5pmIr1FStz8OMObT4
gpapieXderMkmYdfs/j3h8U6wXw8CHm+PFb+b/108RpzDNcV6ei9LIOFZaSBoAlK
gW8C81uWjTC+8NBqe0dl/352s4jr53zT2DB4MgRl3KfA4mAuHa1RyqXeaGMZlD7S
Fdii4xEEPQYcjcSZzZZFiC3bqAJRIhoL6DygWIxfLutQcNfRJlGbMVV89h/pQXdH
iY6inGngxUKN7qNmU99NSNWFhpiSdXInCa61i3KD0rCUKZs2nGTHTNodgE0B4sQ3
+3vIz6SX530ro8O0mLgTVnwYXgZd+fejVewtl3Mh7enm3lh16qDTv4f1lZV6lzt2
tI08S/30gswXjNDCs5fEgPLxinTG+6dHYBV4g6DTS9sGMAp7csiARiHNrt9OMKiz
o/kfyYRM/oCHWDuhxn+D4quIvBMjrHfPlpGfQx73UgYIAUjuz0BabznKnsDHApB/
v3HPUwu/W6ojFtmVMt+XLTnVBFOBkcL+tq9ArO/jL7jO2LLLIyRatdpucn5ucYnW
djas3HmCoUYczV98KjSp1Tegp+8GMvSV/CPwwqDQsh7dvjg132FpygIu5gAj4CyH
vSdAo5RRHi+jmUbRpnlAPeCst8nqV8AIfMSi5cwtXIXKkMXQqx3F03z6/v7AROfG
ZLgGoqnOcOWSCgNPwlG0W/mfP8x7Yk8BHOWO0agtZX63hJaXMBvYlmktjGUr0RyR
CVY1CZDkoNP6/kTzI6GOi2YMEI1W0UCt7NnmCngV6hXaA7iEKR9Pzg0hOmfGSUob
zN5BgZ7LbtPfRa/lI3avXr4CBqa5+mLGg2Ty6pDnUkZLqumJ5ZjBA7lDVFUu+7oW
/cnJ970hNEFv1nYXjHzTYKF5Zj1RqAhE9K0ry6+YFKOHlnYG7H/8MbudrMDv+ZiX
zBqZnpWQdLQJLjHCjCUc4rngzjEQrgTaNOrpP1RfBB2iNnglMXsL58xZbCMGMVbl
ZcS3C2UAbTDGEQATl4nnujt4ePxADR9BpIVxQ3ijWOVsZtaStMrlxXN8syiC/DGR
CuTvxHsUxl++wEhrUq26eht701Jvagj106Sd2YjKIyhl1+uf57RZQuE0/IXCpGDf
0vl+n6yVXk7VV8cANUZrHdY/jicUDz47nI7nkbllbzvBlTV4BQ53Q2wbuFyy+fSG
Ihg2DmUEUFzvsT7V7Tp71PeFxt2ERca2FX2/wAz+egzFbGSmuQDhCFdoSSXp0dG3
6x0h2OkIDnvwuS+oM4UxoPQJD47H5TfnTL5rKSyG2I3jmLPJibwKXikpz2Y0LOY6
OqwNcFE2IvhxR2AFP3cT2xcKje2uf49i1keXilIg807P4q9zkzkdqC8IOtXgeJ/+
ZsnNnQNFzNv9ytXxq85MXAwUjBCxd99Y7N2u3DfJ9u7dD6ECWqSEegyiON3V1v0v
5h0ZXMrBk1IpvmIikpRhiy2XRdY4eB+J74+WWJ2GgKS0MFHKbLcKmEssHYI0EgP2
HmvbHLhB/1CAsE5KqyKKuWKdpJvEQFglOS9oiPbxGE9BdmCc4xfzKu7+ljwxIVhP
I3nHvBxTezWCk9tmYcK3izsiq4KfBieb7uZXkT+mEt6smryhNrK+C1BOZRmYXVsm
z7U2XgFYv+nyKpS/Ebq5U/52IZFPhKX/TyG+Fu5F60SgzCF0P6hmGiMEo8xYCWm5
u200vWxIVB56FGencexOnQBBEsJ02Dw2ZVLpp5MI1YnlWSbVyKoc2Jqx1pnW/sM3
4F0k766YmA7jAlMP7nlsy6UVyRfHV6KiE2qeOI81mXIUUsye0YYZLVhiyXyOmJba
Cu1BaJz7mXvjitLDOPvwqTx5cGAwWaoPLDvhdigJxg1G7zjeQu4luToByD6MbSiW
2l3FntISjJ5Nl9NFazWLjA2P8KAnxCv6kI2j/a99eFXvhhpY0S8UiIq/+3cyzHLE
ux06IwO/7rk6G9jpfDCxGhsNmNtnavcezKuEMyJBfwLliKyTueEjW8OvVS2Y2vE4
EFSaFF3WTzUO0VYySpFdObuQgK9Fgr0jDSKlpqzjWFzW9JpRv8KuVgr1M86ae2Sy
v09NID5Pk/+LbY1VXvjSlqO3jxJW+M42KLE/Qd2WfHpzBF5tn3wywq09HMWSlHg5
2C8TINSvixHnR0EwXGP9H7tXcmxVEyJSO9v1YGsQFZ938NLcdLoilTy1p3VRMO2G
OFzujYovrVCDEfzEU+bBiOGuH3v59vmSZnprMYZTC4k6+HFTjFt1oZfRp3a53tJn
7fmwTER6HSbSOJSpYm33G/NfK3Ke6ciQkNHEZmI/0wyVMftHXDebmibGMfKPE7x/
1AZxhlwzg0z5se+08VthW2P4fiNGFmeIy15J+r5hkmMo1wBlomai7l7pb6g4cvFw
a7pplUBS7HcTAyK9OOuiBkPJcjn23ShEY5S0P6G2wqHzzm833flAPbrzgHOQ7ANf
LE5uaJGMSpzo4fp08QDrXZhxix/0grbLKaaemJqc7el0KnSCDVxuQfrzdNzDCwJ2
pQDKpULjlCHtztXebL+Ar4KY7cMOMTEJLlaKdNSEqi3RdLXCIssNM9nw00hCdnaJ
8hBmtUYCP1HoPS9SAtckkm+gczeXWvdnjVamCz5RWVjst15PyAttzi03PEGLiGSc
RNzbULEmN4MzZvAFhPwPkNK1RkT3L3kqp+SJmG7Fbxaj5b6QOHUTZXMwAwIWoT08
+Dk2CTXuldq6327mzDwqzg7EzDpBSBmezn7uwlzX4JII5Qf3lv647CjOHMvICxvD
A9NKebabK1M/VoF3ekKf/R0Ybb20Pp8x0r+Wm7gTxAT7L8DzdH0ff/tsf68PKcQF
3YvmSr59T5pIOPNxjI+ZSP197Bg82jwFamxE202U0BYGig5Pe8dWfZaIYB249YhC
oofOrwGh6Yf4lNOq4moL6PkQwcyBOaSJ04p/YySCDNVY7ygO/pNCzM3YIxdZMgmj
3QSneGB+jMcVjV0CJoXtQhsE2JSvJCIVC/Ek+N3F9KxyX8QPjjm5ohC4CCZXM2mG
zrZdwak5kAKfo4Q4foFAeuM26jc8osV/BvL5hjmUtKqQ72tMXK07D11wqUzBaol+
fsQ9XKKEI6MkznONV1rAR9WvkKHeloYLcYEEYs1GdSwffPWQ+KZv3agORTGJ9fbu
JydZ+CbE9tDMz6iBq1IEPyxFyEu5N9E59rJIwaOglnLB41lLreA60Qf6Poo8qCAq
X2/Shm1iemhYio7vGgq5tYoEEKZyp5/EZ+x5rqSPF5mLzkCnBEJUVu1m5ueVjMxt
B3EcV7UhLlYjThEYtoYa8niNo5W3FcXgjakTheT+pKcEVBfGOI3IuU0iMsjHNLPh
H1XEGEIptfZxTavylXr92461sB49t8Jtk8yB37gOgSfDATkj2CC43v6DX+ZW3V1N
IsvwLSansnpPQNoH/vwmNfVJjdSzKkJlQJ1Hp+xiQLIGeH910lyzxaWTHiEOzsC6
nngPlITiWHvgJEQXZR2H5DOhdTbQLguxKIDku8vG+N7dFIEyxWmtGtrGjwzQGUbc
9qwMYM+rGvAjx0/IhFqGOWnzLuyAZwR5SfZywwjdwKSKsy88BWJtMhXp1DthK9La
0a6r64cFmAiWUtsXzwN4dC292kIEAN5zIXt6agsot5Xfl+g2IOdvYkIvgeZtaub6
BI+OUP8nRFa9luvxZegBu4ynMCBPrxh8LE84VoP2XWGjWb9jcLF9bVxiZ+qyYEvj
TLEXW+/FDju84cC7TqOplRSY0+LjyB3BZ8eSFpBSgGma2uzGNwErfBNaVTKhjLUu
P5V3/o8vzdYUzAksHtmUt5QYayUI5jF2jyYUPSLODuYnGa9nDq5vegRpiMR7nsIO
JVlKW2S61SAe6Dq6FujHAiyDgEUXYCBW9E+Jagngx8YImlxf7C3aQFU9ufF9PORG
CkrRuBMRu5sntmKj3S+WiBPtwhlopHT2QJKr5I2wRwVSRbDehTUC9701r8qvQjlj
iVE+S0zU9ZjFqnO1s3Fe9HE981tz1xDM/qDZDSzFTn9SeqYbAv/F4wxAMr8Iyr7W
2PrpvgcY/413MwhnmGS1zMgkzm5/uP951wOYlU1stkiDKwzKuHBBuoKnNMH+Fh8J
iYjqnMJPPuy7awDUWujot7asGISl1m9vNYrL+KeBZoo4IpcOFU7sYPgb5wN4HQF4
aoiglRiNmwoF/Z06Q9hdqXeXFFwj7zSryPke3D9E3dhDf/4Cai+voysoViNRps+8
jv//PKvUucioMBkY6uknQZ7XcC4VYjyXjR3Gaf5+FM9rBYB69OBisZpU2RUjLUky
uWQiMlx9yiVAgj2V3y3jd1eQKXmdTw5UXxy26YpUzrRhPkxSmWA6ozXDjQFRMH0x
M31I3GXOojXNbrbZD2/lhrn2eOLGdvnoFkdl7lP0JwFnzn7HOMG/lJDy4fKaLFPy
t2lB20dlf5fJMpTUDhacyJ76L85XHOUkIw3DZugFcEhaNnh5ptr42rHIivzp+J09
06nPDGiHPf9/mI+Pffsgq2xbEeLgEEkuVJbK6hbn1Bm9CWfgT57dPkZJEb2CWgbC
43flfLCwAhH+RVny8oO/nOfxsXItB7BbXOyiPKdhP0N1GmObVRHOyhewKG46eeVT
h6cOe3spR0sgTKyEtPrniIF7vWTbmZjgUKbHkEJ5ECWPzTTCTer5Ud8aIsuFPNkr
q5MaiQ2eN4oi0vCQ4eZ9pICc9lUcQiijO8NrqvuBp0kT7sUrkQc3WYITwwm+k+It
z9IcwvoAcJ0gaKh7sLxeYuEkVymxrCx/e020x3UwW1RQqgL4B3LWJtUI/dBM1xV6
2Pep4EUmZLuI8pFEGIoBx4cHGLdCYF9t5dUGmiAxLNMkz9HDYQYMdapzMy1GEPsl
UCaweKb3G44XYCE2iYYa40OWVXcYCn8YioVBTSiQfSuWr0DeraxusTbtGfqhQMRu
epEi2Z18f6Q3rnUpQivrnN9/mZs/t3sN5+SD5DVsdSC+wr8e2LMScTFm56WXcSNp
c5CC0xU7TO8W7sPgDw4blzTmUeV0rNuuyNOYtRrmd1vP8p58Fx2H4rhGUm4/8mMv
+kc/G8QqIiiFgrYDYe+c6wxELBsO/eN6Bhh3dXr+efVOBEnWR+UztU8ltRWAzUqK
z7xPiuy360+4zy7VO58WQ1oQBc9QegRLrSHlqh9OtGLTEiKCxR1azLobzDEBH6LJ
TprSypWSv9Sr6wYtJo+QXQbgy2fO3xGkG1pOlZKMOLDmxTZc9NmNqWXidPiiHmSC
WIgD2DDSmQiN3rSx5kTQi0SWR14ERfcPhXCAm3hp1Yg+ZLxec7Cl4NYhLodokkCW
XXm7lusqL89e+bfyV4KInqCCexKnqI427J6vn7u0hDo+g6KFKLppAmCugVGuEmWY
HAeaBP2puU0D8SpH2KeSET944G6oj96BNYQYwUGqMTdnmQOHTwLbfUsp1ivKPdzi
mIOio/5KEAj5RdkifsF6cgiJaknMTUUmWyABS2wDZigf1GzAbZu064/iqA3qxVc1
Nj02dJvJARUd0WdviIKD1lymF1drYsvPweZSnScdIcC7fsEqyp9oG5Mb1AWUVBij
tT+E6vTui0ARO4BFV/CRl6x7UX/Hl3e3hfRQwCeiObxr1GSwLrf/5uL3cM7k/lNf
nDu89xhYc17RKts0e8+ooQPkYv6qISSoEnvPigGbuKjGtfx3MFB+13XsTQspXiep
T3R/Kh0wlWHQA3/OF+0wX+xaXI1oD2e8I+We0Nj08jhAuh8ADAlNps+DSGE8qKyW
dBCVzsRMAla40kDK9ctjJwUk0Hbx9yUarH/trBl17K5hL7tys39LLSxEP+M9swMG
yQn5pszl/9bxD0YQX+QMnmEPG1g8T1byDE5PNMT3QYQyGVNlmP6UZ4tfa240PPKd
tr8SioKKrftQ8osa3mYoUf59LjsWocyiQHq1RAnKgF34hIAqH7qjcC7kAghJhwKg
1n1Bz+ihxoPoSmuC8mhFtsKCw48TDKzFrCiS6gjJCmeCqdV0/x3iSyzPTJbjCbR8
glNrN3G9QxologmeWZ3VaXpeneWpBMVh0JyOiuniVr4WPVhUXl2WEDkj5nGIbTbE
ab/lIBojcMDasm3SPR1wg2PClObnUCTiSjlotLHT1w4JDihu418z7JmhQ4CihbZK
oi9h/2ZTkWqqLp5ktljHr3MaU6Igll/XvhDIhnhVB/08I6kGWxO/7zVuYonP4ZE6
nm9ksdTrj/epicovNF2uv1G9vOfehy3WMzPE/SiwGy77sHtdPjq3tGhDkNB5TvKU
mVDEZ+beqvel7ViKCcWZNqaxExOdq/0wS5Oq1uiaq1BjpG+G/qbtjjEvdi8dWSv6
T0uwM9aM+lzjdOvSNn8tmUoIUw92TjEKvPuddnoi9QdUBzXKeLfvdCP3TnIuB4Sy
NnHw8VrPnaHDsAytcAcfiSQf73B0qEay4DfBGzAYqiZU/uv2VUg0LHd9Nt2YMScJ
/QlbLYDw8jVtlLXQqOhICNy54GjQIdt1yta4vS7uby0Y5KuL1DuShoOQFIz5U8XC
bUWLklmF6OhOkTFpsSFQzSs/2B0O/X8JmLgwWe7mCJhU/GnHWuy9od44V2w26U9X
s5KzwxASrAPd7cr5EXQHwJjz3eXiyVeoksOEjEyoc9tQtxbwqx08w98O38cjfspv
e+M8b/pNam6tT69c9lJv7xl52hI/eFu9jfpwLr647oLN1WFBk44ZI7oHLCWRa/bp
dKvaoNC/iF8yP0Rj+MHt7yjvBBxraF53PIqu9l8tuLBYYMhkuAWNaDibyevo20bh
P60JsXTzSe5DL+o7QD4uE7AyCtYkA5NGu8b3LB6puHhrYyHraJOBRzrlfWCOlJ5u
cLP/Hna0jPWS94ELeJCl5A4xKVz02IKiiB/1WIl6j8slj879Iwzcr6rG6IBVmh+S
wVZgN694MpRsxSEW8XBBVfcF8hCcYupo1PkNR5fEkigWOHkAaDDfBAQJl+jkRR14
CVV+Dz5nv6Jj07GY1lEKVhN/rqBRrx8Z37Y9IPEjqE4H5PmQ7e6IypaYKbqoYNT0
Dkss4Ns7apkRNeYqfV3UARPg1f7rF8cU0AwUNF2kg8y2hhrkgDfr2478Ag+ygrwq
BiseR1y4shvOIvsvvLC50226mT40Ku21ZGqC6nHnpC4n1iHKbbTg972ACgb0NmSK
3OL9LG+NvDOg05sZJY3VpxWTzUFamO8B1YguillEys5P82WAouu2my5IIUilRWBp
vQW3OwfAGVf7087cJPTs8H8V3locwymESNVHZ868RWXNx+tdbl/A6IPeDtQrT8AX
7kK9qw0FNj7KP96SPNfhUklnLqQfgQ5mx4IpkNAbGkJfaHJdeyctubdt9TnIQgIt
KtwzaD+tDtbndNtGHxlaJtaznaqo24K5IuxYp2hmSvxhE5m7JCZFv0KPfgPI0cAO
gJ1U+X/qXxu3MIDIWGagcVqDuBN/uBbyRXb6q7inMcdM0EzC3Uf3K+bSrQeo3vtt
sMrwgbyhI9ee3kiyH1l7anLi/LlDlnso2HQoLcL+bIf1xIAVzJtrtCu4Yb6aKfLr
EdH/JlEnFuKm0c4H3ptreA2vh/tV+rkOFntiqSPBfvgNxf0F6bJHST5pm9TiBNNM
7+/6ph49Lk5MAZKjye4auyqc6k/MeV86hZpdIfdPAsEnNE0ftXBgEUrW8d3K/BFd
/nepHr8P3xC8FhkWXwJcu94ySR5bAInv4neU2sXJH4YTjk8NwIGf9fmyEy690hvS
DsfVVd9S4khUmm/o3W47ZWiKmpQmi1EVmoJO8IEl3aw+wsmQmwnx1GD4282BlS7b
GUEYfxO1+C4EaJZ1ZuI1nBFer/MTQsiCUZrxHvRO+O863jOncD02zZ9Eg0ZFvNL6
okfb8b2qQC4y0USDZw4vg5gBiPGr4HY0sgkJUf/vnw9wzTD2m9iy38F/hLSL7x2S
0UJ7CSnC9r1w/pww0KK5zc0G4KlqnOHfB8F+mVdU5FNt7fTJKKJWr5lQJUH+y9Xo
SgbXZYG/ZkY1Dtz7960cPJm9ba6O8bRnRylrHDXLxiOIHkW2wRG+xU52QXXDvwrX
/t99rjaW6aJ0SJTXW9qCQgY6XIdPQ3sHhQy2wPtPj4rH0XEaAKhSGBhHz1B/Tt6S
kKM40zxkrsOm3LLdK0ikGnoaCDUW8i77m0X74kO6ZK+cfYA+ESITmzHmAz8rEFlj
ft2cHOiLNeqq2l8grXMbjaklv93eNybz6oHxaP4onmuGooMHQOvj3CygMHQz4O8q
5HOo9ZZaezeDuazTYcRshXMC5Ig0UzhzPslXh2u381EF5pyU47uGDwVYdqo65/QF
773LmPvX0f/4cwkaRi1/8dFnRZbmAaE0AFoIeMETko+av5ffoiYjmT8Bh4j2kkcW
2WhiWDCKPzjY/z0AMuQW20za33iazqRQV08oXOKEnmgR5l+imDvf0XhvmiAQ/Jsy
OcFaGevnxAdoWCwE1yYPHWKG7brkmSgzaj5jn6mUEg+ifKdO3/hGalR0iZEoUhr3
zGOA+updLsD0Xll2KjunYmo9Fm9Y9336eGHKh06VfTIVoOYOGjM5mcwvtbbEi0sP
HVRzc6GsBEKeAbEujEz4/nUg4iS+Eq/XmxhLyFwXXBDB8oxODRunYz1r6USiUUYY
zKJjawEeMVSdDMvWGGQy+BH0eSE2iftP13H0iI4cEDWH3u02G+tjbR5QZ7aj8X8p
QIjmL9L5GKcXnxc65pTd74JyyY/SXL3/Sh4qkIK3/ljgMd9LFUvnrP28AqiHcl4W
BTZ2PnVU97RTSyTTzRtkRR4xq9U2U04/e4Aw17D5bm7IU0p78747FS87DEHEgSYM
Fbgko7nO3OOS6klUr1RGWanY5jBEoEIbWRvjg6jOEypC5Z9df8pEwLAh9L5APOai
UUYbamJDBLotiHV3VP4/sh8Ex60H8/8wSE0hW3PYjUegmzv562ehdmWDQQ0z8ADP
deG6J+qVYTd8ClKkP4DiGtZk2a16FLIkuCbF77QvD8x3kQ9Uz34zixP3ykJnR5R3
VLRCN+l8hJ8rvKo0hn059S9GX37J7C0VaOlOuKZWYhqA5m6BsZPEEkr/OPMYgA/R
NDBkdZsYAGX6by7vkheEO3O14OwrENFBG0fkfzptM3z+f26VnQr/en6b2KX9x845
HTyvSLJtXnDaRy/UPvTFDTA903WcbLxKH68OpNM/QZaH8IBYI2p5CzvXpwCmWdRv
yRNRb59MJO7xLqul3r9T0HoFQmNrk0AnxgerpPtEiFF4z96BadyT+pJ8QirkiKGS
yweGt3dZnLgN8erFm0nqbcL5AU4SOzqqlE98jrRJvKgs1qWSKthmF5vL0ZP13Tpr
2iAWqLTekd4ZluExZ/jR0r6Doh+VQih1NMOIGBkrBAmMqqNzj+QyyOYUPytdSFiH
1ZuDxYzdCDk4/qFxSAfrSQdrrgzgTQzL4Qyhc+kSQpu/o9XpiuraW7Ek8X1eU9uk
IjWNSkMpzAaP7YJBEspcRn9WAYS9/pPbmDxow3JP1PlX4xYEVHeyNvXpPG8aMp51
fCc33gtu08XEiIQOJOrBKw3dw5MowNgp4ufDaNsxn38+BLWAeBdpuuLp0kw2CjB+
+DTPreaJPWlE4A/fJBXx0C+NSQ8qBFsu57xRApoHguw42OG1v7WYFr6Zt+viFJjs
SwaFWhBCOcY4BhB/RwECuROokOgMYEpl3AI4deZi+l2aVDpq2T1b5hR6I1RPKiUN
T5MQuhaWyYkUpAFjfl8LQTKtDW/U0t6ECCdA1T6SAdYLJOg1lHMZsumDssz/w98B
aNxYWRL51ONjiZtYrjL6ebD9WePChYqm8t/c9ToJJ9t/iE3Ye/TVtVcqH511FP4g
VAVr07oMNzdsT3aTyeNZtoH2Uhq7vJ/q6QAMpNpzoDsDKAhUHzxpvAowcIWg/px3
dGpY5/b+Xno0dawdMaMLm/RY5MgO7L/0WKMd68giXyovz6D5Co6GHqTRAMujYnUt
inzncFrhMzS8J6hh2Ly8eOpPOu39uAbvaAgFZrGUqc/eL4FZkrUOVnlGtM3zARXY
GKykiiIOugBO9FBJ7PHEld9CsgsMBxr+zyobOJQWgnfdOuK6u2iR/BHuTNKGajLo
VcaEdlhdAY/bbAciHlC+aeaj6OoT5ngYheLgw2t+SBRNu+BdPvniKrKGlD3GJQrm
QC2YEVOQB+eHAb/dQTcN68XhK3/QfurfBkPc3dkMBEz11pcQWC6HzW3G4wnRKI+C
C9fWETFqIS19XeQmbcT+rxTbnglFAhWzx+28h1Gsi0Hdvry9pRN1PESUp7qNLN+D
UeWX33W7J4M+THnTF2ivuMiaIlMUtJXrQ0/+3gMicCTNq0rQs+WUeVb/x7ZZiWjz
9Qsdk9ndfp5V6BTXR/0/JcsjzUsQafoPHkaZd1Fxkuz4R38dIRMxrbuID620Gp+5
aNRq3fgH8epDd7BMmNCs/95mrPpr6Jq5i2+7oXR6aqex57pRu2Ax04E3Rnh8nIXX
pJUstG/XW8no/TNi/eptyfYWTrFDi1KkFLxPjzdyAEhVZW666pWqRXwBbo7aaUVq
70SBo4w33/sr2BXyEpqCTyt/NAUr0kN16D+NknI4LRFAJM2po7vHbfNT2Jek8wYD
wD/gua6n38xOQUO1XjWirM0iPIyjBEZUEZ9i/m8Bqp6xLRazpvdW0gq8bR6WpPqj
/0XjJCq360xgvvR6cCjnbPFifrshOpOADkLdolvWgCJs/K+djD8/yjsDMSOfXP/x
FTY4UJ5vFLj8LmZ+mmGtaW/Avg+LLC8ZUlXPhbfjiJUf7nOM/yKYqYbZlEzQj5EL
qRJJ4Ai+mrLSNemzmw2LAQr/+LiKQMc3kXKUJdNOTPKjy1PLohwu3EvP+CZcbDO6
68LjI+q/p8RCuGOVwu4ddlZb7lAVbog8UTzl1/nK2Mg0H2Lx9s0lVYKUTUL9rU7f
I6Z2aS981JBS5sCKCujPnxgWziuhfmG9rKvcmBYlSp02CdLaddEM2NETS1pECs2/
zf+SAKBOmFurTXVrIkZb0QF1dhIuDEkz6U1bdsaFNfIrlTCaDE4Ra9NMHD4sFwHu
jg2qSTZxAhBYU04ehHwwAL31GpOBfX2n1z/q8bwAvOWIjdJEu4Isf1UOEeJrJC5x
XFYxwf0TBgKH3ioUmHgRKZSKXmdF1gzKRZsQkdf836lQOAQmECEUh5wiCLvaPHhM
FiVBp4Qo7vY20HHwLIpBnlAQm6acbRTFaKsnawbdSultJAdgL+BKeQNYvFgEvnyd
iYNWC2xXXMKLVVlZGXX7St/fFIwLF4nsmmVROMKd638FKt95tv/yecvjbEiEJqEz
1EfjhgSOsMZG+2b6+cpvYva21C+jeLCzcmQKNneQ9Hnp9fyVBlOsz1VUEGALkOuV
aRy9U27yjITGRIpb/ctUqjCC2HUyat4PIoEETbiS97ZQZTh+S5/I7DsgKpuFItEb
6ve8xUywPXVX1npIaw70OlJhv1YomZy1p1GBkFkf0KznwFFiZJhMUQr3K+01W90n
RSslF3KdxGJMouEj1KI8UAHoY2afbZrTyTWx+y6D6bQ+wS0qi0gl1GcWtVh0nKs6
aW8aAScHsLIiSazHFzoroOSavqVKPaBVHSYxLykf2ucNcJEsYa1sFKqd5DakF4Xh
tuKRkmPeOtGk5EABbWQQiVTRYzauY+vhEMfXE8bmiS+XChLAALnwzMwhqa7MUZhU
IIXkAlYxKtl811jza3+N6bWdfNGG9nBOO9OXS0Eeb1sbUuagqDgg57XFRBCMsK5h
vy0t4Bi6ATuG7ncP3wNg/Xa6tdl2DWfYh9Nc+ZRs3oNp5C5qbBh6sZdvlbuWLMLN
N5ouRIAo6eYw8CCza1+tMWpBnu/F1vqZHQzRG2VTlZ2mTSAUJMz/CbwU2xBJz2Ht
j9EOEy4w7INkbvR29cfp28hRZ4EK5E+J7/P8n/kJASbZbsduLsGB90OmXTT7J7LP
UnEIcLDPjiuWwTb4DCCswT/gAAPL5FDg360x03b+30j++x7k4Qoed7HgUvbqnLJ8
S/55PzggqmNyk5nyQAvSkQbnL6XJdNrWhAwvRQX1LXjEmi5NU0B+nrO8sfRDKgOS
/gfQxedktO5ypa0LlPkatnuU+0obzRXHBRf/8zPgbS2Ao1ubtqQfUz5qgADNrs+P
Y6z2UjdEHChKErZijX7eeDfVoj2out2ynkvMVyAUnSjkM44kwL/wTa3gXj7/cytc
Q/1ECnDCCv+sircmJo4x5zJLyq9WIq+57ESiBKL9JMKiGNSabkLgRYx5bpaFjyUd
2UEj0DVetifLKfupkJYVLkq5YTpXzZkB7d5VtUzOhNDYTO5254ImaMVoY1nDoeng
tAC62sLDk49miH8QWF9Uv+bP19AGx4HLxkwvFsOZUp1J72MB+Ai+Z3p6iXWNAcQb
7GTydxZF9UbJAxIUtN077ZzExdwSLfIcFYVjsrEXl4ElEIvCuL2b+NpV0EwLOa5s
TnsntXQbYh/us41bWcU+n9SxkxXHgZ9UP5SaDjtTgMHqwAUoU8PCV1u3w28rEEr8
+v7TtXF91df7NqfWCKvAy+MaWCUNu9Vp0gbeWDagdMVq0jnhymr5G+hwGbw0IOrY
+PzfUwyH6LjPGXEycFbLUNAzaJjOdSJZYoWvibW9hgmwvE5N8SuV9JStao6otNaf
17mdjSogC2wh+lRYqZ5uBapKLI9aUBCvEJMj4evUhbE9WDhZYtWyHVoaw2rA4V5V
CVRxqCrY6rMI/q5uG055IRznxFfJC33fiKG4ra7hOFVDHGNSsn45FcTBZS3vQaTO
+3MkocBPNnM2T1d1J1n8gzJP5oQqfF/qrEHmBURPqPIfJRH08CunGxI14XvyJy5W
/wBhwzBbZQAiJ0hhk+gk8qzcL/evwldhybfG8hCuPG3WnMVSpGp+tonQ8Y7gDonK
67PFBF0imV0oV7kcnlV/vtyFusjY3k4brLIG1fXdos/6NXMeTbCHzyzMUTIZildB
ArtVhwBPqIvafcb4puP2fCd7CBFKznrn8+BqfClM6gdgTtZBHilAzRZy+mCwyPeY
/CwAcVKXpWdfqTTZ6ixpq+2YEB42cLZdpMua7KwcJVPSl395TKu3BezV9k9I/+F1
xZr0vLKUmKUCVfi1Xk8j05h22Fsx6XPr7qKNWpJsjGkJhepuCeVjvIC8OTm/wK+1
SfknlQt1Mp6ZY9U1i0nazPFqe/+KAF7z6BjHCEVpAX4O55uRRIHOpXjwejH8BmRE
0HBvdenxkOeAk6CIzB2pSeiHd3tNqii0SmD1MSkgJrFzsHHJpZ5Eq45o7P7Gs1p1
FJas/nBaQqB5+8NVfIG7jeaCRNdqQd00I5vKz69CS3CzJ9RaJhWkEu5l7J/DUb9F
i2wQRAme59n/+C08odA2p4elBC2aJE0S5MJPe1XEeVQQ3M93tO4eBD5zDeUnaEY9
hBaBLxzpXVVTuKqKgCtSErmsGAHWO71211VuDaikVZGZsWS0NvrZ8734els05GFX
TrX7r4yYFK5bVNuzKPred8KQ8qRp9Cxbw/v6a21fq2hskK/p0H6YaTjkf30oefZp
zHi52m4NE47X7HuHbP73GQFl32yNE8dwph7PSJtIV8nxjOguJXELQk1bmNjr2a2r
MdFtvNGYUMuOiY/VIRFWy6+IiVcBVj26G2AdScyjfWchhAjqXLeB+wxdKnghLoqY
sHTjZWZnHZAoSundRGFZx/nTwEEUhnjhZxHbFxpjhCISVk5K0gikXvUK5cqTO+B8
BiVoBa5MEuhl4UpEcTSXMsIfqFRJn+2AHRYn76kE699eoyM3J7B3GVfYlT57ydOk
SWipY2Yn35DsAuSm8H1UO4ImFTItcuBCV9N54+TY/wzEu1Tr2lFgq+PKK2rcIpPx
wSIlZocpkyD7NjwQE67DTubDwLZf0vSmGNtx09NE3/B5K2vyr4BYeQ3/FIUKJQ9f
BST88Odjcn6nw3Gb+33tjyRXg1CoyJs6RYS4JuX3RG5anAZKy9khtcKyEWHirFsR
ixNvyc4oFIKriRpyuGitoyxSDuFvBMrCL9ESLfrOsi3rpUyTUKdXh8C0JTCewdJq
KVzMDCJAo0bZ3gsmQVn8NMde4lIeevowVQqBRWmAdLIDye2Mn8enIKOV3SRanh0N
DJ7Jg6UvRQVgLLdICr7H+5GC6D3Y2x92Gh7uVWp8DLGV/aRFnZysDyt6Na0UDvjH
165pfekyso6XMHjTIw71e5CzdI3KZyig+n2pX1gJTMnucY5OR0YMMuuxNSdhBKkZ
g2mUJtWAVinsU480FzLZFjj8raD2mDw3WA2JIKO8xXhe9ga6yyI2Bz06h8SEPgJ0
pn29xR0e7aA4bjrlD/78jMmeWiec6ZsKxypC54o3l8n/wiEDoZl87N+UZlkAfJnN
LH0LMacqUJHOKYZ7BznAAYracu7hDd3zx9sJ5jO+326f6TaBE9c3osx859SmX/7h
DkeV6qx1QiWbA1A5hyB24eCG1aIHEhSLSd95e0cmhPfLFQn8cn9V2wMf/dpjffDM
xrwmXz325F56AscwVz/1pqCF3o2tGSkGKCQ5rR8tGKUOtNKLkdd5P4/oum+LcKFD
hrM6QFjrDKyhJRgU+jlkGNy2WL8HCSmkrrZ/2OzHggR0cHF+x0y+CQHijtIcrgan
a5aTw6PqqLfA8DAaKRAiz/3z6tv1eOgaYQfSMBfbuB2DjXWojbaZa8TCbCwDKIV8
ptzp/tiLJwT6JhlzXGgHWn4iYqiJ9YaDVmG2mEgzd7h0VUOW1tQiIeUFaZdu2fDN
+65xbl7g8b6x7u6y5txafvkSktowvzXsfh4X6lTnsp64rLe/AiDZOh0iB51DHQpp
AZuB5EMoknnMcLE2uafIguuHfbYKTOAdMq7AWU3DGVZCTFFRHwgbuRhjPFKY3q64
Ab9FLSZTsGoyNkrnZ5BIpAhVmWZf3mOKXs9ZEEAlego1i/drSKsTTSOArytVHeh4
b0E7OeRmVUa7948/+mV911PCpUqHYG7KB/ONGPcIo9rH9wWKL6c2kMtgsJuWkMty
boBqhrM/CmnSG2GlpKFo3PxmYujBLnL98FaMP9bR6aPNqXXaHSV2Z2yqjKydqIYH
7YGWbwQ3KEpdczdDitTlXREyQ92AANiQGyYV0w4bkuiMJDpgvXopUI31gYtSb3GY
dIyWqQOWoUoxgcuOoYPI6CPJ+LNH6pc91PWPyJM+qEtMNDzNJgfU3oo3zlwLzEXd
pn91606XAP1MbVPgJcEUjGRKkGrrYcvHdDQE28sEEEi1QcyHcaPb2sHlh4zhHt86
IduFki62E6LUtpPgVV+RpQyMdatTBg6Vsc0/5wr+YRUbdjUs4AF13T5rR4l0QDp4
DS5d3LGk32Y5LO5tlbNOBmJ4EeL53PEjB3uZQPeeWAd34745yJUmAZ3PCMb9IY+a
GPMAq5a7kux4GzRXWVNLA2Jt6tEGcte70PcitsZwJlUsUZeeuunTvelBkf0q+snD
d2zm117ruZ6GvF4BtKUVIqJTp0AVRA8lNy4RRc3LRwJDK9tZM6Hgy83NH4xgqjQ5
io0TDA4EYcbuMXB0oT1f5iKCMRVden5z1yhsRqyXVP2Uc/jD2m8JFP6hLqcBcp30
V6X7BZgBpsbFKoBjCLQJes2yLUJFRtAAnBTKTs23kC/Qa0ZbTA14VZnSunGP430F
M9jZnVaJHmkunaPiHPLQanjNZ4I/AgJCELydlJv6C4eItCNf3LGgvS9+rHir5vnk
u1dO1YIulOfpVH2bdPt7yG8nmwRCRsm5p+LuOinBpCs61bgBJJkVnakz9LMMaEE4
UptqmUo8VSFA8RC81oJ64PaIEKotjBXpnXSHwB+du1TJJDTycV6Hp5SENKcoLxCD
wvXsTnhliH8B1sqArocbUemfy82Z6gpinw4svljUgk0tLFnWJxRzrPzIm0Pc0M6E
hNYITPZlH4FQxJxRSVhlP03RCoBF18uaFsGSQdff6oAmyWjh9cfRyEJ33gvuDOpz
oqGYui9hTQE4IcIF3X1TXU6Aw7yhqRLxi65voHXBvQZ2Xn3fObqxmb6vua0MN+yn
1+YPnZhuweVHT6yxWIRQqd6qTwIN3XQdzE4DP6PQd9iOI9ww3R1szE9vfZi+qyFl
5cnTQah1et2HrDs4dLH4vOiS4rPCASVsKmOr6qIQHSOCvkR3bKlDY/c3Bj9cMpa0
K/5Or4mQKRiUtJDmY2/PzxsdHBAT+96gPoiFjDWyHUetzsQz9pKu83jkTu2ILtO+
3Ts8KzdtrFPSwwBcku4G0/DBXcZdaN2J6+DrtLRW4zqa7X/YKWpLCp17aXqyPrse
OZf03iiPeLEIEm0f5sIRVS6zTithwgmwzwB6HO+TKLZNCPJQ9Klx6jTmqJ1x2+MU
mtBxArpYMl27+KA2wViXVX4GkiIE781idbp+xQLYK92eTJvD3+P2UbvH3aQGkQ48
tv6TL3NZwlvknM9Wo+C76x2zIPSeus5WIQKgD+xb7CkskbQqjiCYC+iM7lxpZr1l
5HdR2lee+G0LG0Ju2E7xEvn+cT5xrAkTtD7J11nP++NNRuyXM4QBZJUnIV/gICNQ
eYMZOx0gbPM5gGUUdJwtz4NKBdjbjMmfpp6vfcyVQ9Rf8vI3BEo5nKsYutp3qRLD
J8o+z93n7AlHKIIhWdAF7Fjbq4PiIq/A+ak9yBAcA2GhIOuWmLt0SfHt3OZXEQsD
2kPsQW/a8FThFR2xUljzkGciHzWWitXOlt7LLMM63aYowdK2dsGXf6HbHQD6wqDe
Nps+ky7lJ99EcjMQSQJSKzuVLVHf5WzbZ7XKW8hiOOygxY8OPhd3CKQ0XgzmgDmo
JUY+jF/zQAN5+tMl+C7vOlygVUj6RFMkw+J7VDKyhAbtcGiuLR9DNo2pAxxX1jrv
gIVdLl2YIxylP9h4+4k7kk/MlCu04Y7OSNtgctRpHBLmXF+LJBYsUElpzYBIgZiI
mWYeco/mPmzBl4u7yE+X1/m4/6c0YxuHNW1OJeBgSXvUSaesTyquyYk8xcHTiIrA
mrW5HEQi3TidukZ6caZ8B322InZ/zy4Vz19ELdI5JkXYj3b7UMC/5fxgiAyNEOAz
8tYQ3GE2vzmvvgOIwp6dGWSCO8aXzpFo6PZjlO8IjHe7S9iyJLbk2ccq1zuy0vtb
WNuh8LisRcWeHUkl1T/CMKBBKlTz6QDmev7JdVYoB4AZxYhWEkMp+1MxRT3Ez6fc
Uu7macWGKQpcmXTZsuagVNvowqlZK2glQ7sh79G6X2xHZB0BlofwbD92IlYe0WbV
5h4+VZAKFhPm49BZwuCoipYVmyENTcfa/d0VTmyZVnss1FsjgcP3I7q5IfWNXwr2
v2QKwSJ4zVD8N763r0W9oMLzCoCF13X9tZiGY8OIrVF1QLo1n9QWQNGBtl3zIpfk
h1+oa4O14ekZCdTbmIKK1Ns9mmxKJe5VP0+5UKFtEVip75dSvNr52i5cSDyfUJBO
Dmjyc5vnXHP4+WbsVPtHcE6RN4wYzUwlOhtQP9235R7YJqe+hQLlvKlxCcpvjyvH
pgNJmFrxWIfeaKjhPRxrBKm/VVmTgmdMYT85DQIqqlP51d9tBTxgoNG4WyA3UJlI
72jI4chdjD0+7mrlDT2v5qIzAYyMjqc7Ky2waARTnHYlGBejabupl3r74PK3Tve+
9jFtK1VeprGp6Nitb9T5gD2kWoqOUe5rzjlM8HoclgKRtyPg8kAC+ljxM4AeMbn3
50Q72rPwhz9aWRQU87gAVzKGERjjX5tK7SZRCO3dQhD+nfu4GcyRTM98rB5kGlSy
SroynjmKFCVlUNtnUK4S+L5a/dR6UXwiniwuzMMjY8DcYpnHMaUSpftKezbgx4cz
6uNgCnXlOvfwd2VOfcGLDXKlOENjlmGv+aYoHwUkoX6REI4jJ9PpNtpYA6S/0JtL
z+cUH7fvnd9ddrQPJQwmuCw23HLTpaAHHx0AqfSzVpLqsU3p/CyB/qRajJ06VDg7
dkv+J7R4NyNK0fHVksGhK5XYK7oHdEwJC7iWhohJkeHjej1HpJHG6lZ2EzGTZB+J
Hbis7m6FzQxQ1WQh8/z2H5qiWULgxKchMtx9xMYBNxvvjqsQgAFT8jY6MNvxUlXQ
nzMlIbSHALrN/u25vj9zDF234p8R12tpc1G3pGGTOVEn/3qHqJVLE+9QCVHUlJA3
ZaeztNk2OwuSuPuC17L9pYyrgJk+hFdHjHaTc8+VERAhsJpjsMgSHfPsfq6KwFKX
RNvzhKSkTH5N5CulbagaK9SXaJGQAaW8x5dRzVRHk9P0GTB0gH/p/pBkJoDcpN4F
R1u5fjxAMV0eg01PJ0DbgHWGnvYvX8GfUhAM/zBNhPuTqnwBNoZC8G5A6ofgeYvC
J5DUT4DJnJp4EiuBADlUNspyVaXdzu7iSWpElh7HKCLqeWdXH9EC4V8Gkri//mU2
q7YAu/KmCMqKKpUGcBMsnRewopihOg1eUzJGgvoQ5xluRIxjp0FiqV2N6G0kW2Mt
Er37NVWtW4hVYeQqIdx8Y0am42OURENkPxYnYEfRtvtC2b9UBncxopSsK08hgl7S
/Fhf06NbwJPzt95VX1r0Rwrfv2sYwaCzZeoOzK0hbu3NShyLvzl87Mif4pFg1B/e
pSI3nEKzN4PenYPuh9O+66M5FT+HKtnOSvZLprlMdMKE5j7Eq/AdCxxOfDSC11gE
lI5Uuy7UBF+DxYfZFTA30mSqmhHX+sgF40+TTbcEcV9RKzBTedufzqtIgjOiZmMv
NVMSvsVFlnbpy1/0L/T86fGmBAmEWTvn6ykiTtdEM0CbPdzbr1f54+PSmchNF8H2
cYhpcQrDfpfOcdKcOLwgoh7JxQQqzqwk8iWj1dl+1uaMr3/xJeKGOfWNJPq/sDMQ
LDPMZY9XVJXHIHdg4K0p2Y/kMqERYQB2ZA+e34Zw/7VZkBy/Oto4mOLllh98ugiW
dyurh6qaVlTCEdubUrSrWk0xT+J0MbuaU3mI34Btt+HamlTah1J8ID9DOKkyLZAs
QqVYQlmjKu7uHr+G+gWvR1SLEH+9pfbmcqOWWBl/p/Nu6OS3kNZPwdBmeoJUsRsq
suFTfGEoVIRLnauM+DEdQHZePTRMR2ylaQyd4aQGbO2DGBcpweDX1E7S2ssurbst
RD5aGJOQ2mRt91VHbiJ92d108sZzT8b0SejJYVaQc/YmhmMouJ0YhxOh+Tjw8JaF
Hm+UqfkITXSmCBaXZIvgzZ1Lkzx4ZThLy7PMDZCWwMGdXXDWWKwlMjNmo/di4dgY
HSVvqj1z0DTd+7ynLBYzcPhCfK6Wz0F34XHNgiVqrUotQTVJ/SKTag6hZNnN8+0h
KWYO+addEaFqTZ7iDH5y7mhbybPq9qzgMDcnkMVaZ/LmaGmfBeB4qzO8MXjnODiE
ezzf+0rMDhvPgsC5+xtwWOeWcHoNddfmTUCPeg6jfRJbd+fod/REaZQ1QAvpumqA
YswYc9C8Fp3hZkm/XqaoWwO4sg4fYPO00OSKPaj8tZKGJlu+IfAXqIGgz+QhwFEF
5iDjVnQLBPXRJteUzoV3kbgHs6w5Igy+JLQY2Oqya5E6lL7Gja1/EpGXhp/6OaVM
GOoBYAWx+hQprfBs3JXjHyqpEaJt218bl8erlkBhj4Jo/shTbrxfJiZQQdRiIqQx
0RKyQWQU+l5sA01gXmHONKfguWyZlVqVjkAPnHoVyJXmQWgaRP/xRt91fy29Lmc6
vOFyJ9DQUswvug3bpyrmab+d+hNHxJZCXqq/hqkrH8H3CBxEMjTEp2Jg9LOySw9p
YC37pM5DEiuGtvfE235+nFlK1YOE4bg481hW85SEz+kf7zVopprzC1HQ6muvbMLK
a2graaEmDLsBIi9NvSwBxT8MVfBF+gwcfaxcHg12HKiL9ir95jNklrUGwRKizHN+
I8P2X2dMrnwI28XP4XMeXyFslbl3Qm46dQBLApjTfEgE7hqAkn7h9o5jd26sFVeE
YhB7FEqPSMVNT0X7oxW35Dke+9MFjg0gnJoBD8jkmN6UMSA7Yni1UPCRp4qm9WAm
JZtHbTi8mSk9Utbt00EIq4pG2MVUhVeomo+kp20Mi5YsRye2BWwEIuwSQW9NjJIp
1ITILkO0h52/Ge402TnP0MRzTpxVSxs8C46qNGtm2+1rYs9pVpESpnhXKhi/kfpY
3zgjdPAJk7jx/dJpUQAszSrNWQMfP0WbF3Eki9rNyqcIFVesVT9Jnopma9wXCuuV
ZDsyTwRGZ1YlAhQ4B85Kyh3FyK2fbHDSIQEVYVR2gj/jQYl3p68gSXamuRrz4fjU
Klzj09gt/xeKOufqELoSUb9wxy+YXBJlVWKEDFfmfYOEx9AStH5PEnjAeMRHRS3A
PVZyMC2ILaO1R+snF+FeFPdAP4xUltUQ3RDcIEXexFs8aCB6YIv3TeCwHu2JTf86
+7CDkvfc7e5o463VF9Lo+Mhc+9YJEtLd+OdNRt5hazaWsf50JQSSWr7kFh1hRaq1
fnff9C5drgWMK1sx8nSvCZoojxKg8yM83jhTcl7G4cs58GWlfumgx6srElTlJv3E
yshHTLULpmfPx3xhYbKGvkS501aypyVWfbxx8FEa8Yf+kqRBbAOa0v05TPtZoja0
cLFo9p0CNlOCghaitUXXXfTuBa4u8vlGq1D/YNNiURNrB6eFtuFSXVs76Uv9WvAh
1f2sQ+vgFVlZdLxOdklY1AGzdiflGWedNXI7fiiB+8jHkc37HvjxOLg7RwnokqlM
Vrr0tR8j+3aO/GPXpHhHcqowvI0NfVA+EVaD6llhxMr3+fMsEQpwTLEQ57dnB4qS
uYkkeHNe2+LVQEwBhz/GOrQ+8Vwpvr37clXRq5XUAn8uEZYZ/NooPxdaz6JZqyYg
V4Pbl46WkQmtAn1RoRXQo8R0ejEplM+u6QQM6xC4dJMg4MrkA5C7HLwAdauUzFge
FXA3CRXYG3i6riZVYK37kIfSHQUv/D+hGcfn1yBd5TsChs3A2yXysAx0NSJtXRos
Ra8YM2pQgAiFFRItbfb5lFg8CHE0hNSuA06YpXS5MpmYzHiHl1Z7cCjyzXt274Sm
v3xpX1MPfJwnz6ZgNmdPhGhCvGWe7VhbROz7YwFtDGAUaALkuzO1k8o+bpKKRMV9
9ajWWZg87fvX7M11h08Rm9vwSbwjm2AtEK2PiASAlBbUnYWyY0eZFkIxN0xvR6gE
UcPm/Ewp5SLn82LQf7LxC/RuCMu7Qz6kxTGot8lAXIvWpMjchitvyojFzXTngjPy
7GOP8gwkvI/asxiyD8waT0DEY4HUiAf/qzOY0eWUJF8O0ZTcVJh4ugSeEYzZgo8C
Fk9FVVIeFvB4pmdNg9tmRHc9MlqNnD1XkRTp0scJz0qpc9uShN4wye9nw1uAF9pV
2Ta/sU9hcEgZzNeaIXmskadthYUn7LwWldqJ5oqDms9oS69J4FZVHfo3+wHp6ni3
X+M7KmXlz9wun5ETsfbrUfOyofHTobIme74Do4SADPiTJlFXkXF24Zx+XCqGIl3M
b1/W2wdRoE1gpXeJ+SaEjJIdGHP3jwJMJiwEVbhUAPRtlyT1i8HKs5kq+ire4QqE
4YAff8JgiNJ/5AswtGWImVvgC/6bIsNO7eaGaGuF7zUgkQdSbSTejxr0rMicnf0V
+bFodzl+OMme71EVSUgqWcXkjiy5mYPCDCr9PdwiYeWbwq+E0VlODsQ1uwemzemU
o/C2hO4natHTaIjxarihs4GkiHWzrobGsA0XQPUvCmHlsqvGo2LNDZd8FZjdf2ZP
5IA/RNLe8FYrqAXR1F3H2FGBIijxeNdzrEyfxEBHJsyB3C5uprMbVRSoi4De0PhS
jt/udd9Tl0iizDyhSmX4uu6kReQaLEMKlBnpUyMqpW29rv6hYqzSfXqLzDX/dapE
hLNu15FWHqgmodtp3dk4ZlwxHuF0jAunpMbjs2wKyiAIRaJg5TSDGLTBytDOyOCJ
XnYQDkCa1h0TduKimr3023bqk2obXqzjizTRtGQS3N5Dw0h/+oL1F6kQGLBEQNaz
C+sOOZvXRpydpc19UNLCqg58L49sdakWFyOj70TJ90VDjVMeRe+aUiqXuP9cCUon
0M83npKf97zNlvapri+ajQeMpso4CbOqU0Wuvsk1Y7csH8McuSyWDezcR+y8xuhI
SYHlVMsO8gIYj6K9y3Pf6iuoFHnTHe2oJm9jucXkbtrADF6k+h0bg9spiWBip0FH
4hr7og8UlS/rYQdvmsgRbKyKe0DSsHGb21uikMszwY/CE3NadRxC/K4sfX1uE2wz
soQ/4pCBEtcmIEiXQkTJblh8F3qpxgSfHfjjus+OTPoLDY37RjxpIz2E2iFwelD0
NXTX22HQ4mdczh0uWBdi+eksiO3GSLNRomxtKIE1kBcX9p1RCX8r3khGj2hrMe0/
vhstXYAdshw8yLxQx2rKeNbP8IvwAQSe5LnnW0T8pcZvoJ9X67Zg7mRoYHZb/rG7
EoM9OHSreDzx+yPoytzrBN5Z1JOhqoUnc1JRWPwh4Vl1rhLcoj0c6NAwbxGl6GBx
ieR64TD84wIxLt29jhnityOtbTVYWaVXDsXTG++fB2iUynVMIPBn0NUYOWxXUGtS
BSfy4MXN/NBxZcCdcwqf18WAUvkKSsmxaTxdJH88campob3IaYOBHFoIVyDMdyO8
rt8jOyLxyeYKjX8e+rrCxWPYCCcOr6ZDCIfnhFeBHD6aJLCsyIN0JghWn6OklELG
OTSpPUb4vqOHcpNajomW1ZbpusJCoUTdCQmng817VmYXvKneCgELdhcnmoTnB6kC
eCY0bRHXna0hZ3CaEmxZpvVRl9mDQ8XXbQSt5BZ9aZhbT6UC5EIt5gfcFsrK73FZ
5mz/dPYd9ZQnnQz8q2MuqxyjX0In0tjkwwD8I4os2HUCy/gBwn6d7VZbzjhwK3rR
9SaLLRDJoBqBc73YhdRoH5Hj5uxeYR0qfWrMCNL8ev5NMrps3FMLh2sw6wg/bo0U
5fq1WEj8tqK8R+wOyBlquEQR3RzmzmOhetPr9y0kgUpUEJtBYpUJakYDZ9p00EYG
a5NLIz1ruFfYjeDhj/5xELWyP6GOxvER5yV7Kfre4ojFx+QJs3oLVeq1oLIj3UMC
pu8/HIyy21HPkG9T87+B9cjKSkh4hK918mKpD5aoT3m9zgKCaV9K25GPnGUlWmxe
9h1tMiY4wtfBGXdKYdbdN2LgI5NsYlK7pcPO+4zajyOIxqUvnDErIAXfwht9Y44Y
ImF//5O88azXWIzfD2xiCqie+BxVk9FyCYrmRxKy8REZa3U3Ff0mcyixX3Pov0+o
72o3TESb5Xcm2/C1iwo07lQS/k768YfAW26fn8VuqtGlWl08l+bG7Qsj2tM5Vu/u
25YZbSEyesp/aYmrXrK2U36C9FFWOWS7jnOoy1z8KQo6EiXGWUmFOpAwBgFwTbeQ
k9zuTJeDdCTGei3qq+LCf4fpcUFrJmvdvelodEQgg8H0mhD20xvcPTMaF0Y0xIX9
AJU94IrBSGRAZsDCVTIUvz6R/s93qJjnl4+l5GbuXoq1dwpBnbM8s7ojx7+Qf/yp
StKPFJhF/X5qM02XHgQzIrDq2mozWUmhWyXqdw1yZ2nIkknSrBpEHHNXMVvQrP25
vIw5UUtHvIX4Ac4L9gqwcxYAm3sllA5NheFXMZj7Yjo6eV5caJv7R2vDaUNTrrqb
Bp3FalAcNm/2fQ7NOMMXVcsPMddImTL7P755g5Xv4/88sHAUVYX651GtenFP11tf
FyHbeFelcufU8DYPG3upGaKCJEMwyjaUYSRtCirY0BrzCVafCZqsIrGVljA61fgp
/r/+SCcIH4YwUyDz2Y81hKb4sOFlrqwp4k0Z3NI6t2iMIWUVo3RMIk4xoI3kztbS
OVyh+CWEn3s7eyE43tDcrlDz+8BTfPkwpWYLUrf5Vg0RIbiS75dLlNqT6M3v3k/k
lyTtZBOLrkW/ukTJamLSdlVip3xxeSebQ+6+CJTT18pACVaraykAlsn85w6/GZWi
tWWb0ZlL+zd5G05UkN/IKnYjvJ5qXackQbB4nnq8QtJTiUiGY/BMJqDF6oJGXf3I
QR2b1t3w7+bbEVVLL4SDD7CjDSaekL5MO6uwYi4PTIUJ/pgeMBsITVDKwaEnem1Z
RaLqgjfqCuCPfTG/NNDHrIXFa/LbPsOM7TO3ngY8I56piKwU3PdiZw1vnCVdo+Sc
WhDM2oWI34v9mn6Jm/PMNJIu3FrT1s3aVHZOvrrCXsJPK0Hs+/qwI5PI6e5Xob8i
/mdWJ3qr+cYJixo3PKvb8sh04Xs02cF36BOQcEsCNszrVH/spJNM7rWYvUo3naq/
BM2EOroYJOIjXqXVQBHvUhU/Z3NXgL72nMGW31A6acDjgERPptb9rF7xRN20B1Wb
J6xI2c9NklPTjbvWpR+fycinUWpsXOpqEIvHHr3YmDV6SnhDK3IvXsO7CLHy/CwK
Pspdq2yj5ZEzVCCsSqOMwFG0XqEyv2WxoKIMBhWTDK8ULYvlJ1wQt8tn0yHdC0zA
d9GSkmqA2duzaRINBAC7hwWn2rw8crnAsA9FZvsNz7wUyxiY5geN3Yv1gw08cAxp
uwMdS7/u/MRkcl7UanG4lCPZ+0cal3OBr/LUmsSY0lL0fRQVwOoTmCPYBeCYt4IT
3677txtgq5asLq3cH35Ya/oCi+pgqlU57tsDGG2pJza9sVU5j39xZxk2yscrjyRB
NG7CWkn6Rehd4NRYt1MIY38VyaC6g269foPKqL6yVV0J3a2SD/HO/xLUiYS4Lw8O
liPRw3Bq7MhTbE/pDZvwAsQ9SAtmlVRx0cWNvD5qZHknajxZhJ79jeVpLL6H7MsP
E2HtM9iz49UnBCpBLarF1vEqCPobsKKsRCtn5vUx/wJ3vhO1xpP8L495A+zFgcya
n3eRYTR+QLsqaCziPjDzuvq9q0S5vVCzfND/iOv54awNaB9YLrC1AOWm7sdHyGl6
WXQPQNe242QGBwvQk1+TSzpTZx0mrR2YwX65hEvVZVpq5x63ka4IhmcSYh36F2c/
sxZ2RQKkyr7G5u1jQkt/BvFee/d1JB8vq1nVye3l3vHbVNVGipIcnngyKzwRJIDL
mWeUFH5kXapybLufa6zyUzcSXuwbsoAs6aADyCPQ0RQ1A10yBpxIeaQrrhYDEoyh
WkL4ZrwxC+/KasHzL9TNi0mC5NlpONfMFA1lw8okaCjrrcX77GtJrjYxIX4AqyKY
uPMtIZXnjB7Khc6yXWMYJsPScFBoxwig0nbCqcY64iwOSdxfuJnH44Ct/fKuuiyY
/Gn2FXmG/Xd6mw6DlZU5smKqOv3MvX2nb0FDRZwtx7O/69tN6vJJa0djURDJdtEE
0JNeE0BQQPZBoae0mxzb0mWEIKQmxjUTG6opWCLH6hBisruNqoWvGa97gkTIETSX
TlLAl0HKS2brE/bf5OBr5Y+73xP0VjVjckOmU1LWM4RwU9B9dXDYEdzX5OrGkDv8
hHjCn1auxYLs+ZQI419XRlSmckSfZ4wwLQWjYUGVA80h9rr6QGw157+XEc9klQqm
U2VIYM2iMOgl96KU5gK5YIjJMMwPENo6GXKDdVwUkiT+MGst3RsuGFNlHqmSNOLt
eonjgOkO2EqDWZSXif2KJW0soUXhsrlg/suOOVa1Qctzyo7cKossnnpnCQVT68R/
QnSBK4g0pDKj7o6irP4gJ86vNWzKzM9TRgDlCVKPFP92xQweQ3zeUSAraKaPEItz
ZRKc0EnFfp0Bu80+EpxFi4O+r9VteWzIUyvjdfOXYKxm/fI8Tn+w44CCnmBm0HPU
8KTFFbGjKdNuJ9U1/Ao3Vb2vfv0WbTpuw42IU/N7y2G5WeB+aggH+HdcaHm8n5zT
rZae6Z4w5HhKifz5kmrChoI1AHJVAkIg10QBtAfWYyTK02WHCLjyunELHkiolRBS
WSWZYqbhTTHYrM1IxJhFPOUXPnHTPKC3v7Xnco3PKy43WY1L9LlkfUj7VX/rPUvd
mf+Qf554kDSMccvF5lw/QeSUhgKhp40uLvujImbT9aJ7CBO6PbtxBWatEYwewyp3
F8TomHXdxrSoH1qu6E7/O90b+NE2i3jpksr5Q10kFN7KsoTCrJfDbIhaWzgJ8+Td
iyQopTl8QjHIw1VuKwwI/fJ6JhZq6r7IPd+I/lXoRkUYNPfmwUqgkhCDf8QPUOIU
iH0Ud1R6idg0iZ5p4IETUPTSOAh3UINWcsq+wsqLnzOY/p9NwVRx1EGMAnNyC+f1
qR945HqJAWJWAlTHFt18FIW1kWRGc/DlgGvZdlP6r1SWBbc3wc4bi78hdf5qukQl
/j1NzUXB+Xrw8DBgP59ynoJ0Qc9Ux7T+vqDHEB5AYSclNxTZkltmfPFD2Rnd4ni4
CtpF+EJRDM1VR47VxLbln+axSLLOGsDSsgLjsffXizUKD5Calsod4qAB2FnXymGk
SmTPNrnW+6iyTCukZkAUyP+UEUrp7BkfNUgzOL9IaEm37IDhMfyTqyxqs4y0HUxc
g682tlztrFAGIk5Ugj4mhmKZSX51p6bugrgIiak3R0mPJhkLCQ2TyaPxi2Q0O+Ey
tAAiH5oZ+zLyovr2wxeLnKQaahHj1xLp3mhjK/hDS1gGvUkXRADL4/gVKGTnlSMY
+2hAeiwV5rTeJ8JBMuM1pH5ojP/dpYo5Of2GB3YAYo0PsBLQlHrwLpPrpeiXFXLh
cLtkUPkagbwLbZy1VkKN4oopnIHQopF7NcN7O/elTyI2g4Womuyz+IHxCYGT+piw
6WJnbrM6jldT7+OfT+A6t35xlIOW6rPx13yuRDQGgZh+SpPLUb8LVJVACVuzQjfx
LdHrcEHh1clbpXMx9QH3ImFE68j2e5VJp3CPHnqAiH69UVyJ7G7kVFMd5xy8Uw5X
GmskbImc960EQaiYBAngjsIHcvtZn60kFDclp9PNgtXy+nAjHUocu6GmyWXg1lT1
CHlqWxKgbXXZq+ReKcPHeLYThW10wz0bEfvxIk5V/a9oQ5cnoqydU0BDKbKIsVe9
6mUZPQ2SGxvxAgph0lgFLaTl8uHiJiVknYqIpT3N4dLK/U0PLOG3Qs/UWUXuUQBK
fUlO8FW+qWnBci9UOyMO3Q9E3icD+vXaXcAlKHmG3qzsZZ7cvQOxVLhN8zvULVRm
p30oBua3YL6Ydx3q7QE0UoxKy5AQbNTs9KXUSrfAZAvzlU3QD/2kZadCkzIwigNI
fOwLFVVNr/1t9d7BQnujt+DXL9NKbBF1lmywM/oXV8Vsg/jKAhRJTm4fLFGvp/wz
SyhGDPov/j1d9IOFf1XgCEnehVrIeY5RByODfKSfnuVwnfjxkJ3kGg83FzcnfGCB
rbHI82yqwfQhVBWUF6b5XEWFYuVSayEhvUNmM6OalpZuOhQT0ryfHcVUZMp1q7uc
7HpfltFZ9OLqra2xTU/Otw8EoYlF8N4zlwH5OgQf5Sh3mwgfWxOio8C+1zxtGYka
ywLXP4byuKGy73XrYoJ/eQxfC7btCO77l3+0CvQLfGCnyu+nEfaKph8LkAa+NsbH
UkeZMgTpOdPCgFzGamJml9kxZCQdRNzn0Mw4IOlRkrdz1QH+0L9huFNoPy9Nn2sW
vjZq+UpJgroFf9m3BY636CcP435LvoyZHoYLyyYfWz5Z8XrA4q6lghJdLwWq7KZn
GpD5AnWqeuA6ubx26YKjxiO3+gs36aQ7dkTZNnrCb8ezMCX6EBgadD7r/Hk6o9jY
kzNh7kHZPOfb9gx4cyYOheK2B7UH3VNvnstkHw37Of6YSHBMiB1lCl2Rp9l728l7
6k1cd35Zbp124aEC3BQmfKLPPxW9ruCeEU1MpmSKMoFQMnqIfuSR8LnO7aa69Som
Iblj3ZQ5AZ25MoukMeXe7eZZut1kC7ad/qWIdXmlQdxnyfE3XVngMURMx1DPRW9d
8Y2D+jyaQRNPgy2MVia2Yp/pp3H3FHEanU7mebLpfVfl/Rh8u/6WBQGCvS9AsFaw
+OWq4iegzXrKTUIPVrzuMo/1s6Op7Cf8mUVrVb4sZ2OMnl74xMuWrGGT3wwePxiE
DBKbYQXLtdpvPra6lBSm4n3Q5FW863J+EFSqG5iq2K0NWtSe8IK0u6l1aiLZKNs1
344qSwUSq0ptWeWcsJnCk+QWNOwtl3oD21fkMT+iZOpcRLkheGseJ5QtRI+0/ad+
AshhA1vlTQEQdVB2o/+dssET5W1gMcNgUXHCQb0vY2cz1Mq4uKFPxiwIyz8vet5/
zIr6zS0n5N2aNXt1h4rmVfiJMYGvoiW+6bfQyHoiD6Olo1sTs5HaAlv2nQyUiP29
H3CgSwEXWL4uslWYbjZlAZKpNvBWlnI7BTusl32JDIywemFEw5YO4sXYUJqXDmVb
XyVeuKWRkKSMhtUppa8ITeiZn0zJeiqV/FS+7U+ealwyN6DxoEK/B2F1Iv5ZHNGX
odLzGs5c+cteSjXoNoSbwZwvxbKqSjo/vuZ4brcYiwCRuC/WbvojHnVW0FAQG5ud
Uxro2nxkz6HfcJGwIW1GF8NROmKsoP8Y9o/z+/c4ocVvm2yWGLE6z88H0P7jErZP
ruLE5Mc6rvDqIPFvJ+A18qG7R2fXad2HIryhar/YYaN2XHQZ7vLEcctfHf5QtBQZ
lZzQDObcmU+YAxhfwBAp2ixsIwzOYySI/aaUMFbvuST7RUWL1V7vSutMwTZCnQMo
laA7P9oDIwAoLlhSNMNdrqXHIS9DoLMlNOs3FqQRGix3VjxY82tYlfO+N9H1VbSh
2lBS5qE/FDDruhABu4PeRgHMjK4ToKH5NcL66q/8UIpv+YoIqxfxDKUSc8PHOUOf
K5j28Mm7q+yAqy+IJq5GwKbFlpbu0uGTk4FzuC5be1MLr4rb9uDLBJRc0y3EYGTg
DZp1Zp2O3/4SgnZbUegQ6IOkhJUGC39gCqMdGcG2KqYoINtM0uYOEQOGbK+jdVkb
PI2t4Amym+EIeJ4D8KFfgRJTYQ2EB4AiN3aWVCicvW1aks3vSM18GpKN45pWHlV7
VWxCCAJKK/3N5blhX5pGaUL/htkaaRpdi/a8lP6C5yXXV+bBjhinwNE1cKC+moTl
JrS6Tep8KhPUwnlP98Uv++J/E0j6uuu/4xjZbDVklnI14723WOxbmJu+QBma/JBd
KGTvwykQiAnho70+2FIUwu7uLqECkZCT0l2bZgHr96/WZC69HjulwIVgwBY9ZENV
hylFmzeU35AYd7CN2Wp9mlrp8HM/XQ66DFb2oxDwd0YztKVK4ImRqYiYNc8QG2UU
9BKBKg8no6c9qCVcLhX+wYuDlPcdz5SJZ04x9taRv0NuddzhI/v0oQ7NXvaKDPou
x8cQHKKWsL8QUYhwd7olYT9aoxS3I4OkFTawOd3W3GT8926OjU88aVQykx2QibIJ
Vh8gmkNTtensW/aeeaN7Mptn51w+s/oPiYkL7kTsPqvvNv3c7Csg8/EZlbkWNIq/
pDqssEbfHBfNhPv2UMvUesewzGvQQsOg6lLIvaHvVwZvF380pjq7xYv66qcAhVTa
dYC0cplEpUzYwU3xoThhS8RCEHcRZNxOHnQqv0OM5SO932RGWYwCi4aPvDy1KWjD
dpJPm6D0mDcsdpoFas+ulKJt8OGM/9roIP0qG8H6W3v37i+ryqtaF0agIJL0Lakd
d736ppUM+pexdseCpzpsJOEUcgbO2VrdMv7nwGewa7zIq9jHqEnMjMy2klU1R6ad
/103Cb26GA085glKuCnjIuG0Dkk1DajQdM1nJLwgIPiK/xGCtjX3Rvzka3bhhot7
lG+3Tequ2OF4BDJCnr+Cq2S0GP33aFlAMYqfKBDnMm+qCeQyMCXKj/jawTjra4IF
76HqNg6wjGwE8oBkUvCDU/Q+1zbWJFin5m1PLpfPianMJpqHUn7vkIupzYJCSa8Z
zqQzjrplL1gy/q9XBaha23YZ8HeljbJv5x4W/r+smNEU4X8MwZ1Ht7TNmKhHYsGk
R9pUHkNKWHbW8N+riPD/SS6iOxviGhiScFzTSRamsOvJWWEOiIpMgliXkJsTAmLs
S7JvwjO2wtkTgMmgvoCNB8gnBaTBzLFwtZJB9RQ5wGmSc3ihoK93G42nmdzh0ADp
huTDdntyVf919u/oMk1Io0me7TU1Gi51VMVQG7NkLp9KCDaNsXtg/8DJ9MRtJ2GM
rADEh8NJh7ymPjkefXh+07AROiqrW/jSIITEFYdaLWFMHOabObs+cnwZAAgOkW21
y+6wHDjZbe/tXGbfxLJR9oTnbjfyRCnOs30lMkscfvubDqqGCol+r1hxmifRTx1L
jMNzxMP/LgaR8ea5ZiggSOIZNQb6vTxvDDcM6dcqKR1pOFEGegHuBJf+WSsoeCVM
TNga8lpEswOyXxBMTCFv55HHwYVQZ5oPZO2wIvuv8gam4gQVoL9j/KdumjhYs71Y
lcJLC/IUqTg0czIKs0aQLT51jHLHLqK7SI8e18zMYDpghGSAjoh8BCo5iRuih4bN
wP0Bkbs5eBrnlLxVl9aRw1KB/hDt1Js8CEOWFQuBlHqzx7JYIID5UHb1Q9DHZTpt
1ySkdFptSAoqZI0W3gkaVvDuLIDryrybB2pXaY5g1CiLy9MaRrcRp5VMHaaoFvnN
ZsrBGJ6ntao4mH2Gqy/QCzIFbCTRTvrSyoLC74biLW0Nuj6ZUagBdNvHbPpTfPCQ
1ve47wp+O2tcfff3ox6Qm/0scZRaGbgpYlRABibzZBWzFcYla9EOGgRjtttQjosf
tLulkD8tDOJuPdGfUKyeIyJXZZySDaCyubdMXv5DuWwLFkr30Qh8gFbhiRZFIDfx
qVDSbJOC7Vh4vEwyihZpxzFWW08DQVP/PyOFTmwpzGn0mxonmC0ghR2SUdqOXnrz
aDxinDOrxQjubPG8zQHLk0mEPkxqOunSVLjgGoLOnIVXpPFs3xt1LDKKplWGzbpW
btPZkGHqXJJKnaGd6xXhfILRoN3uOcmtmVL3dL29io81HOPzcmCpdMbyAFMP1XIx
b94Wg3Ga/+7uE/vWaYSMS5MUwNPFg/XS4gX/27Ai0VGOriOluE7yEy2XkmtzpcVB
EXRXAONlDlBhN/aULiTE8T0uIHuqxWuHax6GiWqHU+qslOugeoWim2Kqud1knUhw
zREoijDp+Lg1i7bhA0htjxVJMoR7YRbbykm/Fm1P9XnjR2gDP8ch0Jrtt6jrKiMw
8wwctQsMabVuaukr3jGnePPDYxxK6C5vKyB+fxyr6QQSXjNVoKrxviBcISn+g/OP
JdXoGNdTIeDSS6auNy0BGOPFuiaIT04+lKXK7nPYtqQJDEj2iQR2JuthqrKFjliK
cJx2RAU/W7KovwNIV0ubS9RvicHdIk5joM+ahRg6zkmBTv2O5KX8b7FD1nddnKfG
0urhSLuUvPxaIl5Naigr2Qm3B4r/+aoClS9NFuO72P5R8GUFxDbKXOYFHiVG6iqw
kGroZsDYHgr1OgbE8ZDja+2xd4/tVjPSjBZUkcTl8xZk91bTDtVOZihUSIoh8Uuq
7Oi7DcbyB9lqlchEXxJy0Lamck4mAMMUK/BnlV+BSiVHUmrOkL2uT59wo0hVrCh5
/3KgbfZ/Xne4a0KUGYo6K2x0z4/rnxoxbNI6nm5Na7sA7hc2K6SQL68SfQRh2Cua
sQOPw/njuwpQCJVnrEf5hvVBDSpaA0ZuL+Nt2cVcWij8DaxDbcwcP+PO4AzyscoL
ODP8sxxp/r0JAv4FGzaVINnli/ecB7UXqXat3W5hPFgNwSo+QjqVIF9mPNcRb64K
eCuPhPl9oeTTc01+K5fgLTEVEZPcwLRPzP7/nep6rdKcCccxeZ5yHva9imT40oNJ
TTbOKi1DFPQFFxmpFtVqPINKtx91DuM2WXyxb7BXTRO8/47GU/53sCeH7aSZ0R/S
ZiVoQZcbtjuB9Vkn5vEfCJzBoQIpAJrazZoH+dcvwa8Fz5QgOKpUVs2epd79fzJA
3Zrpf/pdaN67c29M8yptWHO3IZIfcmLGM7385umAP68fhF4wooyBVn7s3BkaDJU8
lKtDEiXVEQElqRtFuEcbcaMCcxB7FBxOeGK5zm0RQd9JPBTQ+vpn4PekwlGgfImJ
XsTnWjjpayywUDF4uI+q2TkK7GZXHfZ7DKk8wwnU/UTZLw8oisvFnzFNDnQcTpn0
xp0jp3lRNHgel/ssqXJxCI/VsjoRxR0L7F/Bvkw+B4bLCWH3+upTqYuFsRfmTV7l
oyJ0ZOohlTcyHOL5AeIdUkTTt4pntn4nsQ885ANj8lICCe5yT2IRaKIdodUrUzf8
LsfF4J9kRKQEwbYnOTTRK3MkM5auoNWfymN3jn0CYGsG7BZUOH7eBkv8GNkNQZb+
OCo9Pno0/LVNaKpn7JBZtGbK/mlaL76HRjOnIYG/jTuDX/0dZFVntyisyjWhI6Qn
i6u6BuFZaNFPQnz2lyugyBT0kQu7GaV3NuXgqSs92RtqkKFBoQEBAO5yxFQjp7Q+
/GNJYC8e8pwbahTbHPYYIP3ksTmlz5efIRYFXYS9R4bL7SOrk3/9vb9B+osMfhvL
mfapJAGGR594Wh8CQ5mvLprpGAG3NBwaZ1E8r8FjkglKojJtFbSh7C8czQEUfTvF
sY0UVeNdQBPUopsOumy2yUw5bcM9n2ZfecTx3XMpmGiiwaFcPgXZTJr+IEkackgK
vsvVTInIte2uLMr1XiVodI3hk0StrgqRdT/TRZylFUoomEUsVQSb3eunitKq/kz9
hg6umoxRZsaII2PKyiOCh+YpHu3GLi3iS6WrdJMpc+lmdGgTQU4/dXpEb7bV1dJ8
BLLdcosT+Xkw78/U+cWDbcyD+xI+CwkpqbBfz6wLJa0S5Azxym5OUHrW7uIlpTTh
0+/nPsInurdAlbvae2/jUvJw52MJ2bfD0PhaS/hLwKRqy2+Rr06kfUMexp2Vmw/w
MhmgTyCOZFzZgx/T3DpOOU72KPoa8DpECmv2/+wSOJnJjpDKSwXFfA/2Ar5qSK2i
vSgs4U6u9EavucqcpCwGG1A9ddaFFZ8SwNZzjOC/L8s/SnyqMd3bXs5xXo7rfD6y
nRl97mrzoFShFzpB0pCJj5sxO0BEs8k+coTxS/xbOCOu9MpHqYtgV0VSvdX0ANPc
LneeJzmMYqSBPPVP8yxtuLxgEqH+B6b6X2HGAghkKIehIuYj+TYUe99hPMzyvbqD
JOqk815n9WHdNzA2KSG/HM+OLF8bPYLawxy2pnbxGG1YuLjFd1MNKn4ueS1EoLhO
evQnKuUBdjC2w2pCPpAoAQCs4slGT9BJA9toHUU7O4Z1xUw9pLgQRGdRKYSjioPF
3C868cZW6g6OYE+S1+sj5DDW+HeKJFwgq4BSQ1zRs6J/hE8u4SetBPQd3HNxpz3c
hBeETqFv5MqepcFI0hTKm0b0QyIm16DuibsSJH6uqNz0y9VCQqscYxf2LDRkxdHX
O4bxvk87Y2hWHvlay+lWzQF8LnsyH3GetQ7oEZe5hY4ora+T5J9Zaexhh9Rm2LO1
7ER8niCMrqxsCzxUu6R43NbRx6oSTgBnRU+bHcSUI9zhVko13nTqM1KqTsZ3WXed
xGBhRbb8qCxFiYl1E+q5BrkV82MjB+/sADj1VC0+Y7/ZtsmLX1eWbZCiZH8llfY+
oZI2/VGPQhSsS2sipcTqL+4X7OUxAtopPIzz0YhGjc42FmHamC/5vi6+gDmk6pEe
2IIhFFfS0oYhb2np6URgxWKbrgh3jvdJVAj4IHmts0+tEE7VPQmpbQym/VFbUQR0
Q8hFHYBATqt9ZLqpk2t2zV5yNUuHjti7IaWKc27B+qUW5fd442OFe6uuA5O9ALvp
k/Yt9LFOnGWEt1KnZItHYnH7ZDoxRtU7KKJbj7lx4+NtfYNLsBeFIPtFn4BqTWH9
YRpU9pqDGF0A7SsST8bPPvKsTX1opYGt4IlGDnyDg1b/vsSdGMetVgheq8Yg7nYl
Wm+jD+7AS/TO2nqK1mO+MS04BOnSaq7U1yYLcHM81Sil+nNDR5IPEB8omAt676Io
h2AZz6rM81MNGAmiKhkVQBgOv5BC2X3je7eDIqGhy1krAdEffb0HJqwcWdOR9Yi9
mbD9MShB+PGfBBlqtWCrD707kzsic26PXKjI7xVfTCdZIlczMXHiVVmDES5iVf8Y
cTn6dV3/ccNnzxQiniY7jeOhICPIsJus+4xsKOroY4jVenjxtkDU/xsnwTgRWqgB
jeyC7T2lXEZXSjqD586EeEMGw1xtMUU0vM2kyUWTIiesBAzemcFzrhm+gID19DgL
d78EopL2zH01LSlJpqs5qJlcukNfc69OyGqytBPbHClUrmEDIoMpumvu9ivJIRko
LyTHyNzBheYIu4TVXkyugmP/R0VIi0vdlPlvXe1cwR3YgK/SshH6FJbFLmwROJvc
CEAtIcedN9hu8ZHuCfSs/ZAdIN1s/M8x42l9PR6Nbs2hfmbcyMq6tXeeZFY8PAyV
4YsEmu4VBFOHyTsJ8zjvrzu2tqphL+uTjeWCxsTrEVOmgweaowpMMcOcNJswSqMe
yhVKOVSbuzXjO29/cqf5MC4Z6fUFtQEYHcUyGlSve2Kx8JPMSBC/UEXQfuxHppRc
p4o9MWDKj/IWTz/IFgsG+03Y8BrfgipImJu6VoA472YlMa8UBrpW0cVo7V88S8hS
k++STt9tZPRPzIkNXs2rnJguiknEU1QVAWQhnWVhEChpUet+RkGgh2GbQtd/Sdf2
bl0JjqphSSX1BRbeNbCmB1cAmKUikUj/alE1hizlvqIYYHHq2O3ZwLNILRp1D/b9
GWY6deSkwrpolXLDtQUG7X4GGDlqi0wtmSUoISWw06TX3fKbAGBF8WXNCG8GtDzU
utQP7YeBycqkAk+fof9Rmdj4rkxES/iaGWwVjsrLVzrupdjHT6fsL11ptoFaNNtU
U1hD48B6AgcD2sS9JRfe73c0I6Wm/Fjnri3S3z1iQKUWBW2qcIhJzNYrD+elv5gy
zm+ot953ZXdvbBjYz2gbt2qQMmtA0i0ti7BIT90ja9k6aWNkqogeujECY+jUIJH+
3JOLDVZoweOLRMD8jXY3lJxCpypADCL2V1klDKtmfDIrwbnO66m+2WpiAw6GpCAj
A21auF6PmFZVEqeVIoU+6Mez2W1UXtqKp9S1OVhfjVDXK5K/FuVn8lHJRvYq2iUF
oGMFWjTLRBH+84/GDgxzS81OWmMrwFf5+vB/kOjEX8aEs2WIXr/28vuv1x6HjQ6+
MqQfViouBbIzjr/Iqn3tB052YflassIOJ2Z0UYz8YZTrGle5U0zKJeAeoYb/+NAq
CKVFERtue0N1AagvAtajGEPeRBVeUFWbiAIv+PWaajVkG4vMI7dPL9+ABRfqPm6Y
yBtcP9VfKjmzNFCFA9S8cNZIiRoacqpXDQyqoNyziTh3mUv05g4B6njTY5BlfidN
eL7ugSFw7px/BMlXH4yu/ZAIlQehDUVEdy/33k7KV3AUNCkUfJMPYZknZd48nYn9
yCuoFFJUvSHlH/j68XRzwlqi4KgSU/Zinxc8OupOUh+E42fAQYLskbnyRqBzqgZ0
VCNmYqsAcQA3mS8t4OoR7M4ew9u35hYMcfnFjJNZJUD1pEuR3VXM1XBEOJPXDzpk
AWVyBxaUv2UNAjgFM7Rh8G3y+h0iKS5DAKuu9DE6WNnykEK5FrM5IgrG39jCQRhx
EatcjUkKJklER8fjFoivb/Kdtft72yg8CTBXOgXt/QhftAaxUzUp7Fqyv9pU4Rld
/ToA5oFETmMGmC2UngfHK3J2Pjp5d5hi8CmBRolieBtGbz3o1QYFR1jZ2p7Ht2gh
IG2Zu8TuD7Jf1OjTodaPxzwbMRIOr07E7lxG1XfeXNeZvo+c42f/vfz0OYNGqjC4
Rhiwi20cFrDbXanNu3Tj9xhMX2DywdtM2E4XRpNYvMhesliMheYDSyKl6cxbnyXv
J8Ny8GMyLFk/KrAPCUdrEYjjXvM6e6JujTwqSkD6hEYvA3ozsPc3M1vONw8qHjuA
LzEfIlgazJRasRvFcA9KZc2/+lr4UoDXfKtapNBewwX5ohj7CjnSVXFUTN7H3a9y
IvSU/GPHIpnsnyMiNwFFgXkiuQ1w9Hwe8+IM26dNGxkYKei0et2jIz4xhJrQESnM
1Gudw1rKXrMAUavhAk7ZeM3kv25wERiXKvmUhXolWA31wLRDfrnR8433kGmmCYDz
rIf1gXpZclJYkPUSq0fcsXxuXNASgd/7jN71n6W++jhGVcWQfeZqcsrxz+xqTJGD
vJWOyggmk85gS3rcsTTg746IeI9jAYFrOmdVio9XrGkbknHcFQAt9IHZTide3DDg
CO7we4faj0zuKeVL1+ck3twLst7h4hmUKd6lsRg/GHfHa1Fmyi5VKTaL4eZoTSJz
XA8N1jFRapXJFOSFhnfoQSNaUwy5D8HQteljbNrT+exdduR5bwxAkV1M0zV2olUu
O5QGIjm9+J5E6LwoGixc5q1jKLN06ndTtwOEjJemr0oBF20ysr03t/slC5f3c1w5
w1/f+4yy5w8ytSZwh+oX+J4mdnZFHIODqRaqv6THIuOq6PuPxRmprn/gpf5p0I74
SgvkMMLKVDNkW2wwwTkyR3LbwlmTYpZoyk/u0/Le5m+VqZo/pDDq5XKUcTE0qD26
vOpECiZ606/KBHUalNv+SJu8rNqHXIYAbcxCLBKr44B37jUlElrvyhlWJxC38ZWh
x8NHkM5VIuw6PYyzrBjemiMFxh9w0dONMNty+W39WgjXI+eAD973DdDt5Q2gwK7/
WMjXVackLjlCzRoh5Iq2cicmmLOnyA5mXEuQXLHkfrRomk9BsWF+KL2bxQxeV4+a
ekbLVvBfjwFZ6BHtxd6kTQ8PNAf6k2ObDyJtQY3ttWScQdGAcJXP2k2I8OVRM7oO
pu1nlLb+Hmtgfgsva7+yMXYB8hdj+/cF4hhzAyh7HcievMhVZeIG+JpTu+Krxfi3
WwpCrHze5RZ9i2rqRdixJfwaEBYVSejBC53loMmQVL8DW77th1oIQHWZA20yu+y5
GeVUT8BRnBxAzuKOfNEBVaZr9G3yQEE5pLracQp/o+HvX9lyWKDKs/AwwkFeIv5g
k7JncDlSfZ8i3AmuZvnDMBirsyEX0Gtw2NqaI/WzMgGdYRf5qIw2EcyeWBvgsQlE
IuE8glzzJPh7e8O9nilvQg76SMTS/NUyoUzbYvX8yr3IzxlqJcYVl/SVGlyW2vPt
4gY3maBomT7aSxhYJD9nJbPv85vvthYzDvQ50n1y0heglU5a7uL/arSGF+ytElAr
A6d5jWGGpe/+BEwtCQUUuuXNX6YqNsM1jgmbGDFs659kR0E7+5ZpwXr74aAr0w0l
SOwPMU2E+5W1y40tu7gSvDWfpR8fNdNNbhw/2TmyBCGi6wxT2DT7MP5jBasyKLoK
jxkunPipxYHHQC6qoUSQL21fgSXqwdtdINnq/MNTSynLWfwW9M2tsfWec8y3jVpm
iSdYtnURdwfQCEL/Nt1tYnLcKPu6d2p7+YS3e7KhUdDfwvx95gk+9I5oWp8iyzJA
7RsnTPgTzYPBXS44AwF23R+m9KYeaFsKbO4HcC79N4ErCwnRvv1rRrfRRSFijOfs
wle5mlj+EBAP3Bn2VLg24NlWqKx5Kr+V5awtKv1NKvzVL7RjjpBFmB/ZGUbOA07X
V0uGsYUaXuPT/92BXiBgrZ8ZJv1v1krzQ0dqqsDYQ2sywpy6O85nGPPRHKuv5Vy0
LCzWCznn8dAL4olF/qdJAYmg/uaDjA85FjPZwgPjGI+yhoAu46E5R6HMPM7t35ak
phYsMYaDbotfrjpDbYaaOum01DGMZ8e59KPHGLw1HEwILDdmJ0u2TuPMoNHFA/JJ
uI9Zzir6yOP7u2eZjbmWPaTUIehdFByRmFdhxexysuVp2jTMTW6sbNtmBSACLLgO
Xacq5pwctXg+td2NIFBdsMg8yYmI5AdHJdD3jVB0AMKZEKkUj9B70K+DXwKW11vA
X3KShvyjTcT20urXLoySC6kull6SQaxySyiuw9k1KgPzW83qEAZy1yCerwiijSgt
lAcvf8HtZsUCxqPCthuHytQedpm1DQMsRNemVYOnqGEy/1uJHnlXPWgvjEQXtliW
9hVWRh4WbobEpBa9ugL0eHOfWC+6ga/GsMCTHcUltlajeUry1qsX3FWZ3fbBKO9T
3Dj+sFWyZzob84QhR0OKIImK9MWI2Xb4NfoPymUV12U4b1lxYL4Um8cGw3jliPuK
wfepy9nzuZVWVV0/WHe/yu+pB2UYxgZWk78TsPGYlsxHC9T+/TJdGq5XarDQ7bCz
Jd7m0f2PjVCpCc1naStQQQt+eM3iKNVt0iQF2SlhdvqQG5xeOSviMw87c6dQXwCp
mRx+DMrbrvDgsO0DrBeZxFi/iwaU15MkRvbc44C6VINYnqEHWMGZmt3M8Uscc4nC
qvdtDlTstwcbt3cO6AmHbLIqPsHf7wZ+o0lx39J0xKoxn5P0WvGqa50DnAIvNX5d
GKuALvqWoiPg1LMb5GcIN1EpIbW/4UULH7K/oZOHyH9zAachkByFrEaf/6ZNUUXq
fepk+/AdTLZs0Pad2Dm5PgH512hngAdfxPCQaHPODABdFqWG5hO8+LX97O2+YkGQ
vBlM4+2gi7HiEtmCb8fHlOqU70+Lvvrv60YINaqTWsC990UphNSlm/IfKlWk6N7F
Q2Z2EnIw06w0CU6wmYkXEfOSK/3m47+G5iZoLL8xq/i7Fec0BWqO5ETqxQUWMA3Q
WztbxtqghjEn4zxFTvyfcQgJKc/gnirn75wr2KjU6hPDNvN0d8JX7ZjcFtSExf8X
jCE9Wp0AjogF2h+1db/G/fFl3JqIOZJpnMnN/hsTBX9lYB6KKhCfhS4zLLwWO8wS
jsr7BtrTdhT7KbLH7mQTPtXeEiB3uPppPDa1jn6L5i3Q2hyYzVOrH6CmNRcLob9k
HWTxQ9sLrhaRifT/0E+O3FX5ESfpAgqqKaYzNsu/DDj5y+L3htFGnlSg9L3aAgeu
8R/wu+Qfhu/aqwSeI5fA6T4sbpNKguMOvRAwBxQHTj3FIv9c0tGDhu/VEY2rxxp6
F3nqcEosstYZL0dLacQ6WtuY3cSdmJ2B1exAZYmYouHDt3x+EtaHKz/w8B1ndr7o
8XSzU3+te7+bj19S4d+Yb4YV8TzGAmMy1kfHuXr/10lD8hflrEkwngYGi6uY5DyE
WFZP84diUa8R19mdk5I73wHO9jVR4ZPX9rCkRLHqEM5JverGcF1gWGaRRErIR424
IM9hnuE8GLJAwmVVAledVJ2/xMp7N3OYrOiUUu35ar/Qp59WjietRNV6jDSQ2eM3
mumj724wjtxkVSPKGn0c63s72ShTJLLtAQ72vZHaHg/Cj7DqONbbSTcexozMS1FV
DSdYzND0oeCU1tPtjge9jNHmy9qdrRMi01NQ1ScQS0r/v1uD7tb8xsvdMtPtM/ZC
39BhpwiMVUaBAdCnLDoHF+7IfTilu6TMoTyrpm6CPNiD9sE20zeDKKxIAZkrQM7Y
eJz+O1T4HdqlK3uaF3ouL6AslpYPSqKAfvd00IJRWUypn+dU9FxiQq3NUJjkD9WY
YuFKH8Jn/1tGu9xwMz6I/4hz8il3R07Hn5WVjnuY1HqfqI7ZvItRgLBLy1HQliuG
By7zq7jgsYOJFCekCQf/nbJp/6+ey/WqXw0AFaZ2TLloHvIZiQrophIAZE+l6iIX
LAYw+6O9FH/NwDP8PLCEN3BWiUMpx17MzyukgwaWalgRtyvKInx89R0TDoVWfJLh
QiJB9X+AYVZwtZOIkxxRTFEfqEPiCyzDxcbgohNd/N4WCCJLm1FHTgGz4PNaa1R0
OIJwUkjpHuizxRgAzm6ISkllGIL8ZwjPTZNpcWAvUQuenIbtcwqXe1iNsW+cjGau
H/GswEv9NSTGjH+tLxsb7+EqNwuV5fAXozYLt7sztp0EqnenMsRWAhg2UudZPqYp
ptrWSArIXpk3dGealrz4ckrTXWs9PumabUWHNtk5bKqRvRSkxLGufYui2M5/ihjd
qZH6vmS6JMBDX1OF+SGKQFmfL9rLm1ssTqqnfgvwKeIHSiRbQWh2BuE50TJ4TVyh
/vwLCrijOodYa/O6gTtYarpnp3i5cbT4Fdy/uKdQATKqVL2Zzy0QPpJwbgPjYDN9
thtniu47W4/p5uqP21IS4VaBgO6wZNYLG25oaITpee8fkDhEgKCoWSyV5ho42Q41
P956m1md8FNSXc1KI6QnbylDD18gk6WG60znKWJXc7WEJxn/HrMhsBJ3dY5msFU5
FtJJFG72/ICCDRTTrAgnOlZfd4y9NcKO9NQ6cNiiK/Oo9fjPYP+9PYLjt2hK6Z0o
o1fWU+dA/liCMBh6BOFckr9WKPB0RtTzDVHgpKLny5TMXpxDkrB0zIXfa8hLp5H9
2bItfltu/8/0rTri70mSV64+ZKoQ+6v3zJxRmVjMQzkw2XL7FZ3GPGijKH4f9Hrq
VoRyFnqDMcyOTPD1BRXVTCTqOwHR2exOmv3mNey5tf9Tz2if8qfXlFj2RbayD6pf
44BbIidB7tB7RFNOzUgw6ZJJv/Pd9NMbpKm2aRWqv8HNAi13Gmt9pke2LCWmzbyT
riWzhkhUHBKQYIFq/jYN+TokKVOF/XMWfD74roYWCl9S7Q/3PkX1VeUmI54PDHmQ
a5rcqRgzKsFKTC/3nOVMVH9+sLS3F1dcWCft0Ajk/RcNugzB1YjkX44IOMfpMU/j
UMaw0gXa7dRWsaSiN8si73kRAE2MK/Hgxrlpyt9KjhApywNB/ZWhpNLcCrjaAh0W
JwfkG/uEyr9X8GIx5sh5+kpFCmS3cgclo7VtjWQZ8010cjkL3C7FYjmsjE/SlDkP
JhmMm+BuDRLlkSWw+5sv5dg3/ufbu4fYAavNdwjIhTi+caLEPsXomfJsBvtyapZA
RYspgb5CU/QrRCk5UMWpDze30QiOGDxHDOatWWHQhxSN9Ia+KsIBCSZiDbZ2EDER
dLr+bzsj2NzoQzc11yvXBfGGbJB8rtnKjv4YK/2od0aqDhbXOWKUsg5YoEq56luu
DFXnSm+EeGgKHKsUeeHa/Pjaoc3TwE2TLFzqDRyJcjhHSdv1le+/ZyBjT/JzYUp4
PF94TQjpgDPEEKmPU0mL5JzBbmnDMnMzdAl8boC5+RSRGbFAzh9LvTLuGYd1h7B2
HprkvxomzdevnZs9EewAUxgcnOOXGvMzpPONKV+am0/KHhFRAEIkr4JHUzh6Taqi
pziLAnooXF3getfpQF1F0ljFF+UICASfA8a2BYWoHwIlftts0WNXRk0t72eAXPdW
HffIYz3vzpvCpu+wk5Abpd39QnSd1DcUZrv08Lyh5dahzwoCjg2Vch9nPEs2cDEx
e+zRQV0PtuVBNjI1DWGrKPpdiqqQd3Mi9w7c+4xESIOiF8U9sjQRH0L13tke1VDV
LHzGqQqNm4jAMg79ildtAdnlzZv2PNXUD7yDpi3PsFIjzZ99SvCC0RJ8Yc2glyeF
iqo8kl++Bow4uEjKt2vDNCNRpEYRw4OqQEn1JQ5fLYFKLObdzkStMwY9l1STQFLQ
h7yD7jm209uJbMMhHKouGygqSXrndgaoJJj7CxGhEqmMZNI8538JBOFo3EhP0cvB
xJSzHzF5iYWDnIz3nIPKf6CmU1OVBF6ubvyrMNf9Z5ywicOwPM/PQKG2zTrlbGJC
XTm8lQA6dPa75KDE52ArhIaUG3065S969jl9GGiFqWEVqTgJOK29kTiPSLL2fNo4
+FgTAqw1WvsnozkKFEmUA7dt08zFYy1eTl2nCyI1+UdvqtKFhrLcK8urAr7Rzg8Q
tI37njXbvcSFNF68jN/Tbl28wEPGMWFIqINSckx+zsdPlahpnBA9ZB1wx65y6kVW
JwsrlwB9RsSl9bQS0rrYksQPj08+xhqihqJMCO3zq7K/Du68ddgGL81dDATCQrha
fu6D2fihOqvZPtNArr+ZmMIgwqWbfWPBgLeuJ+mvnNSFdYO3mdPnDfU7SK9nMLTc
aJdJJ/juNdQiNgsW/DNibi93vaxsElNOkoVyNKtYa9pC5lPNEH5LZxZZk4cP2BRK
EAPZV1q8DYhY/IE+lC2cIOq0baqUkVwnDSiNSsZb3n/FRMP1ab7nEdcaDdgt5i/L
e8OJ6H7Z39TKU3kB2PTWCtQvxUFXAus8Mn04Fru58aiALPjcYAurcCbsfBYd6Tng
wuolws1sOPQV16WUdO9zRTVG+qumhPFMvF4LuoGacgO9eJcWHV+8/OkVTdNwYf3E
V0F0AnuZO4Dc+Elisu0X2+9bgMox66Vu784iYtpQXiI8OOWZHQqfAlJt9S0QWJIr
zGb8DE3iV6rXDI3KQ451WdGaQg2aUSGReWWrcIqY/jUKOiel8KmJt3hzo8GbHSgf
Ad0DoF7Dt5MPmx7B0iuQTkXx9h94pVputtsoSbbdH/T5s02AgXc5kYMKivwLityC
YqYeqdaFG//gIkPsiL5UOeebbkwXFjtccLCGkPGslgMMcsR+9wnoBo2kAMeI6HY2
zpByh510MbGxUqjTWO5Mn1BwwcN1fXYCdi98g9VfMF1SUpjTAxx8iJbDWlZJH1yg
TjTq90uuyQlh64+cLNMGogU/WhuEMMb0D8VdEEjDsFE4Gq3QZkKiEfn0yZDy7AKt
NWk9KBEXk0t0W8ilxbuNne8BV6CEYumn7zLAe6O9eCodeQq8yKsB3qGVU8MNJJyK
4kKh5oNQ9UTyHwG6LnnOZ/LNET8V6H6M+3jzC68NQrBo0aiRGADgJ/NiCq6v/oUr
2Y0q844Q1N1mcuYnbsmJ92I5H8qMREf1RcujBSk2mcYTapfoLgRvdLtYPNwaNnoJ
w3GFJw0TutCNsqkYpO7Fqw7EE/cpZW2a44/aiXpHppoUJb9NbukmJtn9Yrz1jRIW
ykjmQBmY4CG9ADdCzqPoeieYYkkpTSVBSUusXHGEJHhlOK45aAsqk/drNWcwjvMq
34Pkafboqz2pCqBOKDV8H4jzX/+MRKafemYTaSco+QM71PN1Sb4in6sASl+It684
rHJzL+ZUApWA6udChFNfwnzfDPhWwngeKxFnb/TX8jtyaHdW5tH40/Nxknbrhcnk
gMUAjjviGdPcnW3n5bRyx2d6p1G6V3Pk6f5rgYHMDqMmR7AVDex/3/CsgUPd30pk
XE7e/ImGDWZsbgJnZ9dMecG1ePSI3Q274j6rktxhuRyENUZMniz1JY8maNzIY4AO
4LFNhvcCjpR7pzK8Cr9wWpOAenLys/CEHxd7vW4kGLYnw+c6goX6dFWVO+xRV5k8
DjEsysC+56KOiAiv33F4OimBP1Ss7NdhSGXsTuqHRNwfdybGFzlICr13nU1kawGc
moVU7Y22o/0xeHTTbv9SlAZDgPTEypU9pPOlL2MIi6E4Zd5oE4aget4E/Kdk7+nG
IHuNOclapcAgfQgjrkj20jITyNQX18+7OIQDBDLnyHcPZCmh6m6OaSLPl1S1aMnD
IfnKwDBxUcH08OoaQrXdov0KfygSvY2ceC7vKWKu1j0WAC27daDkF8lnzFw53M0u
b5aQC+KELVFPHsC13Lxfy9qDuIBukt2ZY6bMXSf1tF3Qtro2IXgnw4TC3+8m6+LC
mt4Amd5fT4elRB4e3yz01Bfm3teFPk6sMU3LJvAKbq3w8qWFWVCR9SSts2AO6ny9
N0Lv7g/r9wpRsg+1ons6aqfNONLbEUxx2M/yZVnKySnJhpohizw64OGwcWEiX1+Y
OxLXXHWErGOGLf19k74nHY83QtIAGb2Y7ghHSMZ3zeFcDlpGGV2ptEmeT0d78+p0
yswnhYp50bUKB4FORI/HUCQukpxFsjUglIrPyFIViIHSqWNwWe4xGWP3wdEHa4l3
iqPje0jkXLoXAEdedIQFEz6eKvnTUbFpicHFNn0Dh0vBORI/WnRx8cVWwxEM5iQT
JzOMRqq1DqZy7C4XJPC7mTffjnsDkPu5hfrUfIMDs99xnsIXIm0ruzN9Y8Ft1GcU
jCE+uwUkgpNKH4JFXsEvEWQP3TZOpeQOLHllIex5Pc5z5jDuhOQb7Z6EOEEvxCZT
b3Zfs60QK0lVcSNkYIIjEtq7nfUwfoTnpCb9EqcZiWBkYF6QbLQeNwxk9Th56i+E
bu9fGf8KHh+YvWgBuYVdxLp1ETPJ29R1PZK6RbliyWEh+BSa/bmqBZj7NvLAuiiR
lsqsnwtkkoQ1YVDxtGsfByMFjABa1wZUKH7sx7oo9uimJkYhSVcvydRrmgYA+RGG
/Bt1Um12iIbLnYOSLbz6naT1MD4hwaY4wldKK/6CcRtHpUy2BsD5coFjPA+bhk1V
JsP1FNMgbEM9vrj4372MRst+zMlDr5/zwD/OkFSdQY9u/pbf5sko2Pgw5uDnOWiT
EFSvXjR3zSidAckzGr6qPXdEZkPn6eX397C4UHdOBCgzpGJq/wMKp7sQzn6ZUWKE
7Hjrr841sLIv8pnavJ5nNieVlAauu0ol7Khq9p/YVK55YUcN1AHpmwUhXhnOyntW
JTIBJx7SgM890dKpinqbAvz1svT1wSyTe1x79Z2L7OhnzWQI4kM8YK6wN7MfPzBj
D3UjORFJz23w30UnqvFOsIONdePH7t2DdDWbX3howXnX39JNjw4COyPAksOVldK5
rPH7Y6DencZ5QM5Djyhvz0dqxIcagxHPIbG4tZrJHpmA56VaX9ee4h/l+cqayRY+
upACXBBpFaqkQUyHRs6JrJd0mKZG8QsiRbPIfQpbskXEb2cvYcfvLrUU1kmjiCyF
Bb6QRxAKcLLcwagoYab3Nhiih4N6vBGL7vMPCZbRBMhkGF8Otbn5jJ8ebqOyzlJK
psATM3behfusgyKF0pCkokTa1i10gLlXSAHuqqC0SGQYZSkv41h+pb/Wa+5bNeBe
Mb7Wj5xgN+xd2uSsAHOy+yQvuXZPf7OJ6LQ2lLyae9pbyY5uvhdhkI9xN65kK3Hy
cjHmQIm8nlsmmt5dH7mxJnDI6bRfrkMHp5CP/ZLoqV2TZ9GT08OBQ2yQe5QerQC+
dXSRp1oymwoI2ND6cNlqNPp65fRu+M+WN1qHCw4irhrr7BetQEfo1iIUI7DLz7Q0
G3fUbWDEz7aK3KUu/ijgkAe/3ltP1fx8ZqJAOvUAlfcsWdZBs8KryE1Pnbclx32n
pcEtpEgRZQJR0GjUmz7I7fja8Lx4QvyPeCq8XU3xkNXALJRGUynD4RYLjvcs4JN6
9Pw6IgJFRstnRcDfnyKGctHOhZuaLASP7hQ1DmNZbAs5V+wRrVgv3A81mHyeBwJ9
GBmMICFUdmWv4iSfnbIWt0ULOB7EBsSrRZ7gX+9ttAqZy7Bt+wVNMhfUAwj/omc9
ijzGseAPPprbQ/Yuds7Ae7xmDf1c/Eta7UAqBebNTnUkX3axJpTBdJO0eqiMTJ+6
yXqHnePAxXmg1DqjIWwOcK9J39a+X5/1Z3/UMQQ8P8d1To7AbvgjNt53tzR2zwFu
vStVaLYaa2T2rz4LbANysAAKyUyVLagcNFfa1XajwGxEZ8WvTjetlt4jN3b5SzpH
JiREhGQUYR5kxDQzhOd61u12mDdJT/NEolSly6rCKUNcpC812776qXif3SudI/wj
ee9w14Svvj9ng0MW6U6Kz9Kzf6m7ttkHjeqNRz8SPAuOsxW3cnxzcCeIoXW4Ln4v
YWBVqQSz5YkOVQ8M9qUAjeptqwAQ0Z7HCk5UXu/CJTIG2dlMUglLbZ/h0zRGI71P
RiZ46BDBCNXceDt16GK4GhYSHlI/pqwlozyJ+7gyyajCKnGXAgaifnB+z3Ctcwyl
JaTg5LLW7rRxkQ7yfBUqy/lT23KDGVvI3IN56f1s9dAup3XVA8PnZW3G97fHhAGy
jiJgDrVJZCNerJVedlatTTQGY4Te2HroqnxkwBwJP5cMkRmTbnXDRtIjOjND+lWo
52Po/slLx2xPstlDhjT8Oh5+nWuluptzN7FUBvVJyxAB1/vqb38m03+BFatRC19f
tsVWycgP6NCsvRVfhKzzutbNTmNdcLWm1ykwftxExq2UAFMBg2/cf7q75P1D5133
ESu0uSOZmbCqUwTzNnSMUmQbZCPZgRgBprJyTLmTGJDRE0PqIhReNbjyM6Qdl+hE
NX8jtkxuiGTssUyxW2Rz/PJX8kpG5AcbNnYOmusZCrX4L8VUQ/gyzUY8qB6Uy6EX
UfEDwFM8875rhiCp/oM0Adg3RxgWuQoR7OIS8VoD8q1ZryrxbAA4XLyRjeGYkjv9
14vlzc7epkvOz5kWHtDrUaUvosEgdQNikiI76JzQkXspIQzvPCZ6mlr//sJ4KXiD
QTngZKCzUo+KOHMQbZHZ1VX5Y/WOsxiw38v7rPRo126/8h5peaiePgmln38JGS5Q
Zw0V56hZ2w5dSl6F51eEgjzKdyZJNC0JjBCCtbOE23Lc7pNzNJakWwxsiNpL9WxB
yXDNXe3ZbAZ4K82gPXX7ymF3JbPYBoGJkPL40ioRxXE0tLnL58JxHcOcE0QOqfeH
jUGvpA4ncbSquwGA5a6Ur5n9jU/3MctDdv6uFyG/KawV8xKkk38/CjOFSn8jM0yZ
06T6+4ceKmeZPx8YbtLITYgSxUyvQn+0ZHEHFEXMQ3CDb8nonuH06Lh1H7ftWlE8
b+qtyHHE8stGkxvFE39TSbtLjKxg+FdWQQBfRq1xeg/gcssmISNINgo85fGdpvD8
yk5kxdJoCZJmmmx0AgjwnBNW7ykdY+q+GXpziB0mp7wBSl8K/Y8vrkPauOpP68oG
IXCk3msblJS7fqGOVZWqfGFMG9L9K+7kiwuQ6UFYazKo76tX4fm+Llo0mZ1eWKXL
LiYEB9sxH1pldM4J3Lm/5eRP2mG4MhqVJczl8HWlZTaATgvmex1rgp3FO/C5S/fR
j6U7V1fiRatJUr/USGpDEg4lZN6C0Wz3r9ijaveOxR0mXuFEubriGmH5h3mP4BFU
0weIIWqmT9orG2WUw39GwKwqt5uP7F805EHg9xe6fOavYmgAnwroTj1XQbiGoo0A
TyOR/rW0sie5QMp1fNlDRSpy07THf73O5B6lXOgfCjZrUwShwm6fZ6eDgUqGcp0y
CTeu68psq0ZblICylW+SA1NCPqxR3AHRLQVCEGffRRq7BOeH1imwFJ0eqgOv5oRR
0nfnii9vnqaIYjFkEPCK1AsRJY5Bu0qHOwjUcK90vTAp8hh81W2q5zaSu5vfHsL2
lY4pFcH/M5vcOHqPAOwx8hYTLvOTcyHzS6pXDr1PzSd2chrmMD/7KBdbqD02LRyt
3P4vHwwjzJLVkc4TttZvcxch6WI1QhgiVs/ri/23EPWfE0RYYrBWh1AD+Gs+i6ho
FXPYYqMQh0/6GR5+bH3AHgABqkW88zdCGBhzTGXun6HNst7f26cnxKAr6xxI0gPu
1KOqV3BkBh89648rgMUM/V5Ao5tptRNWirYY/cdflkMQDnwcL1KKpKZfP8GHY9yc
9OSofFefeWUBtoGaz56sE4DmPYLG5qmY+WzVtndK0tTD4u+nrWj2K0psHcvk1DJM
MZ+/7SxmgJUXwfKLJfKZT2Y0Yx72KaNYFs7+CPJcHfSv2bkWUsAq0cvLptrQze8o
GG6KaFWHff6cSDOtL8miQwxfpsdQADYJeKkSLIEbWLRjK/lPCHk7TsSdZStSdBnW
Nj/tJRUIsxY5tzvex4LStgWcG2tOH1qX3c+GSk2KehXkAejdL1Ybm4bk29riZ8r6
6hraZhbvvmMD74Qjdw5tAvbYHId6jvb8N7wDcJhXD9kXp5t0NRPhwRgcOc8zjggi
BFN7wKeqf5heSTgkIj6VlphuUBE6ll4yx/95/i+UsktMAP3fO5FG1Xg4BQl6OhoB
+vgK7PpmMosEgqQLBkEiE27oNnHZmUMrXXHlw16RZx5EcC/vHInNM+Xr6fGlpXC1
69QwCq24loRMw38i7z1R239ryJmvXpD+DuZeqYn65q1l/lB0wavuMUMHNyOsvWIQ
tN/4QWvBmll+tWeJJ40qCkb4yl1qN6pfLkBueMJfPClbB2GYW+zIvKOF2Nd0Ihlz
5ApFiE/bB1A02gKFQ84pItjJ3wdGEft0LOsTMskYlIZPNyF3DnYB5caDCzkObdXB
2irTbCzvtseaeMeiHMSkEW+FzzpPiXs7Oaw1WSyumn62xhbs0ty1726nk50clJve
KXPWEFuQM4APnpPGUJKW5Y3Z/ruu172YG9mHjKiEB0YAwgx7H/Wtto2iQ37ZmSKO
f2RKjMMJJ7hzXIIDeeMEucHFv7ngNgfmTG91ZmfuVnWJ/jNcH/lP+afM3BTHMccu
jV8jl+Nxj65DCpZ0wTQCW+9zrLCw1dpaq54vowszEYH9qDoiAxXG3YfXontmYO+3
AAS/qM0HZSJg2KFo9aLjtYmhxUdYyl9aKTqAJRJjr2JqtwAPwAAgYGDlmMGe3Dji
r8iJw6kD2wI/GYcqJEPHIE0HcsxKmmjJ+KvtHMb+dGZhG3CSWEIZ27ZsfAaXp2JN
dMjY1UCoaXtkdiwQre1bik5H32hSl7LL6PCDEskcx7JEuUZNawkoLiBrlvkqKd3T
+VejVE6aibhJsnJXaWxYhkEIcSf8Wa/+WefpLygYKtELxeeS+SVTQgHyiPd8itoa
W64U8p2Q9M1jsuc5+kJHQkuhghKkUxb3OqYpWOQohE1ytFPJ0dOqFFCh+0sT0Wul
eHpr9OAIBI1IKIIaM5fj/FsBYaPxvz/U/Ppad/+WOQMV8rO/uwp7/V0R9Z0GltLB
CUFRUD4GFgLd9EJZK2i6YkL2Pe3IKbo3T/DbJzBxQOEDxcDw7+Y0Hp8QZ+xoLw1R
D9D4SCNT1K7hu4ELS2mZfQE0+05pZGmGH1ttadSN7GH702YvKYLUuXkqSypRhTOT
iyTywQPKxRKa5ymt/AxBnD4D8qV1clG+WyZYB6Mtu0npIBTwzztRsEIJyvxw14Yo
9vVCO2f+rUo04bhr+sW/jyvDtPFiBu87XFovK2xI1qiLE0QIuSsEOoPXvOV2Ht0r
ZDqvACctjgdiJD8+x27aSiUF/fVJDNaVXa9IyuSq1it1Q+IBeHQ4tINzRMVHqwJD
b7pahLKcxhipkiLkY+TyBBYVgaTZrRXQJ+JUdW3ZJApdSjPvJnVlMFGhiXbo8KNc
Zjfw9VPDy4P1XrHhyBsQPkVDf5M/uyxaQfQ4w6ZtlfQKV9GYbe6vzaHNaDV/OYZS
7lv/cpp0qbTSgBiFOW5bZhMUOGPVAuJ8HR/P2CLp00miFrNO3+3CSYmMWBJ+M7sX
x4ndo4OBPFGClkVfjas0t14lFrPsEMpLOVvbsaPEfD9hXwWoYRSMCP3UALj202D/
HokZQFAwYaGuK9sDDMdTUHvWzo8XKf+PHwCT7pVj7YPdoPQZthQtOEom1n4QtUA7
tisSEhxsqdviE+DzIUd4J59OH5gOIyiLI+v7DQizcHfgW2boUp70bLtxvKpyQFUL
V3+ygc72VEfOd3TPsl1XUAP9kY/sdAEOdBylJa8+DPQyQIs47aI/gvgakeSdLnHN
F95iaqvglZwrFFy8rDr/nZPQ4tHSujAzJCyFxAR0nRWxhO+jl/ElcpbfW9skJJvn
TwNa5vJ3bBQ5PGpRrlC4gIvxVZc9N9vPodxlwzwYf4Bong0ynVOEISGp2cuLj0AW
ogaWOd5riJK55gAUJny03wU/kpUzg5sWxbZ9O71JarxHit/Ha2Ms8YsP1stz3LnF
5piBYGxGk5qFfANo75WIDBUScS8ZxTJk2yWQZ0qmgxTWIHYL7BS6+IOvS7MPdKKq
TNl4u2sk/XYMs5v1klosMn1yffZHyU5g7517uDW7SzhnvMVXj4hX9GzejVT8vo5t
jYH0r9ojf8y9vvKkK90Psqx2GcB8wVG20Kx24mIymMdDadPk/x/nJ/e7ttl/b17T
0nWRX3oGSj7OUBa33hUE2d7gmsGsYVy90aM42C2IQVZFNjO4jOSbDpYHHtR0kggn
MZBz0h+btQ2EjA+WNOB6Sk7AUfpx+xY3ZYPOMr3hllD3xnqTN+SZGpCtJfkGMJGE
GxHdlrT5fqwC1ZPEK60y2f2h57RpbRw2M57XiL5teeqFj27X1+5HgReSNnAl8yzi
XP+1tcGWiZTva1V5o4MePLZ63Mx8YE8w9zhWJI9IST2Y/Q6oY8ebZ8NXfSJbqR57
DXcKDrIxqjPJmkmVZEDMTL1w9HDux8fPoLi1tS+LlWUYM6wuXVXUi2fFou9LOyKK
favRBifTow6S4M9O87Q89ZkGj9Oq4T6HmoqingdFh8oxG0CLtWKrJoErzzA37jqa
nPOzn1WRphI+2Z5OnSiuIxeTW4/V7JXG2YMqfSpeQ4l4oMTlMjo+8qNE4vq4d33v
4aDXNLfqN//t1X3r4mkb5zi8XNc0NvLXs97og1b2cCVtOoa8MtqjfIY+InSSwFuI
zpXXe4A0vNK1is6GKjUrNiEfmJbrQjpYrNZ9CSl2uXQv8dcnFs7vnaQBIWMSh06x
LmvmBq2kWilAEDFoxSLwg1+ZNyL0MhAOO7blgq2r2Aw528HWQsoD46TafhwlX0f2
qbh08NQWL18/6EE9P8VHphiT+nbiyl04vyD+ZCBeGtp+W8JoPzEaeyRvU7XEN3ye
flcIelSHTlOlxs4ouYSK9OcP2kVSYejlD9RWkR/YhBJIKzDd75NlJ2tKNN3W0O6/
ct8F91Nkht2neUh0b7L7Tid2cE02rtsDh6NnZyTRHGwNm12tnceRfJONSqsOdS9T
uBH1wbTXlQJIbeCF5drQJxW5jdCcyUMpy1jBZvrrIpgXJ4idvsXM7Afe8Uozp9l/
PGZ/OzEzt7uwPH4o2wHV4BQUWRsHfhpWthELgQeyp1M+w2wWfoAt/dmQ4RvE7D0O
KRBEo0wFzdw+0QxZ4cpxhPWpbTy89WdUiDlzL3Jhgt+YOooWtZs1TZ7op2diqxrf
27jFVBx1yXkp6pbOpg1H4aCI1olxg9uyi5X2aTz1zJcS4nmkeJHXTFDDhSRuxL/D
vvdGmfJM0GPpU2YLNiCOy+L352zafSGYUGgS2xu1y6xtfVEkIM7+OzPmqzdkBXNf
Pm/olX3CGVVt6FPKM+8MR3WZajy6kF0cqTZtxeW1KyQcZhrqroTOY6GJ0WkHxf8F
0ydab7FfymQOciqnJ7d5AM4jRMrMcaYpkd/N1luF5TYZ+5kVUeKMXyq9LkJs/keE
3eTXOxNfFQPoGnx5vb9IhLL39jG5VAmFUswJN5Mwq9gxeA61GNFOU8FybBFMbpC6
LQwuy/rMudnt7qixVpLt97hY/tKRe9cO/bXyCNpWJIChE2qYI5TqS/G10j58hGRh
Mxzv7OkFHWbxI6ucBVb4aIVofJDIGQhUchf/cJSd0K1GRquPiqmAV5FqZSXd/vJo
xeyJZQq92uF2XKwnGyWBPkCNt7uohEtnngQmUAFZ3hmAGhm24psj8mXpETCQxxrR
oVEl6OdLC6JcL1idmsCUNqloGpw5qI7D5zp1PIBw8RFHGfsCmmV+haEU09hr7tGd
N1fhya9aBj0698n+GP4r6+ISpJw8TXyLpewym1tcJe8IY9hteydsrIwie4rV3YUw
TgtgBC3vOuv4ad1zPEVaPDV82cDguLHGGIyOFSllC4NroN6Xx672a4ScByCr9tZu
vnoWy6Jn4cj5vrXgepeQskgr+57Jzy6ywN/TfsLGB2m+R7KuufRyfXXc/BbfX8kW
16dU/GkS49fhJsel7eNMZKzb/l6sFBByCE6IdZEg1QDSvHj+qUEEBKn0BX3K/vtd
UF++byjsjBvMH6A6mMe8BimdD4FN3htKRjKNKgj05GDC6tQfYlcLWijzk38rY4SC
qet0NXq3HObS7TK+H+REW2DHevyQcKxFjvURgb2QpnkBcUZ3oX0KA/zlD/8ei8C3
q81E8KxzsnuU00vm0bL9qubnYsds//ylqf/0fzFXYEPCDD3rLQeaw8tk/eqcnDbq
MLpJnMXSJnajmqFGf5nfonRgbBc8twqlQtcbTxRrGP14OAiCQvv6z/r0AQHtzpWt
8xW2wjq6z86/gq/N4KfsW0eEzxKIfA+t7jTZ15qrJi/+T4Rv+NX+WWw/raUBk5Y+
Z9fJmkE9K55ju7mSHpfsioeQDNC9wqYX5rjRah6TnK1ycnydFvTGONGJXlat0zqC
h9jDrxsshalIkUoufEjafXp8jm/IhidJI3DPdqjektCbhXbyfrSx8zLePb83JtJv
2PG9s6FP8NouZ6y8lxtikbWB9CdT1ob0dhkXW9s4bGCEdD20iRvmwcHvBlyXlq6C
U4X1MrgCsZkej5KnqeY78W99CgTmKNfVf54fNukNjsmHDqSwwJ/vp7HR1dk086WZ
DvoQwpGtPkVTVRTV7vk7tuFPpxc79xBr7v3TbcWIk2TcIiD8YXkx4zBNceMD15S2
rcayt0bpLUsHm8Nx3zYmGKTojSTKA4VMubMMx4m19d2ZKTOUdUBTM9kYHDzZfQsB
mzdNkVuKPnv15qN2TEAu11wvbMAAVQtMiX8I+LSItLFqhYdHycRhGAma/WxOm4wH
FlZ+T8O+Jc1U7ZOLm2YzvrNWhAxSTR0KHPrLEX/1WA9O58f1OPt/Qjk8/ucwnVLW
+n3mO3FsC8D79XVGQUiIEIILmdhuVzJpZL567jonCwJdsGsGe7FvhxxSrc4B6WGv
xydmjzmbfbrmd6ktva9tI8aRx5sk4Q4b1ZSP4FIk/UnLQh+hqwd6lM+RTJfkJjl4
FIzU83rqK0sLOS0NCDGEJC2DKWta/HcD7HRBM4Oq9KX62YoCiWKAmfbIYWuo7Tvf
RF3jx7bwYiD8eQpauEJYD6w9h0RgPwl+DrCrZlVPF+GI66Wg+XcwjYFSyyE+Y1F/
NqlC6BpSt3hFleCA7+xHtaLc3rZqZomMZiuP87ag1hddc1cZhAMPKT8kZ0ysDxwa
ku1IPBdzam62aDUH2neNi7+nOhTiXoFf5fWBStOqKTaCtJj1R8EeJbS5rxnBeICF
dqhuPTHS+Sw2gx9Wq9zEp5T5hkQpSaa8i/CfO5rO/nQ56DvohPHqyYuYRdAWv+Ty
HFZa1lF1stnaz8pmtgvPkdc26gEJ6IcpnD1liL8rWGGbd0e/J6oPNyGRqliB11bH
OQxfnHkXnwHjxAklpA8B5wE6FSXD4/XY1WXlfQX55rI8YBT7yD9iu1x9snu55FG3
a7InESdVf/ThKLneQcfR4wg0nkSoLSGrPufcpBp8DHOMiLBnQb075luZ+TIWd0Vo
S/x/s2OGbuJq4sW23PFVayGgjMTvnTHP7cf5RrtX4a6QuGz+CyWoigsxnZK/W9og
+jcUKvNTnVs10Xx5CkhYNZxLfsUqAYAEa/oOijj7aX6yUO5MOrhizcglJzSxOXrH
jPQE7ILfGYWlSsw/j+LDFI4sqA9CoZObskL3Hp3/f4wXizeOIbzu+lkxIDZJlSkU
XKNtxkSbf+yOQIX+gcdq5Nwpqj/wT4PS647Gl5S1Hps4nbsZR5JDWMx03MciKu3A
0X65tE96EH1izW7CSYuop4+njkIGdLOCi3Tpw8vDV7ROOrhvqMkzgeDGmRVI72zE
phvsiEhvgf5Nj8LXEywlM/CPHN1pEnUjxnkHOol+dfW9QkyQ2p0SSA4pd/+k7g2O
LWXDa7vwd7T93wh3ZN6LxQKrhtx+yBbIbbIlzYRZhQen8XrhXEJ8B/aUKJJTowc/
os3MN+TSkOuOA+vERg+RWmlo6xQBn5/RcyCbvbBjYx5hqz87oxyTJHZAD/nKqqBj
PAYqibWYf8zkdCsTJCKloDIXeCD4vKWHVPoqF45MzJwHqCJ1vXsaTol/dT1D7BbZ
//IxHjhPVw4snrldIsmvIkFYUzG1q4ZPT76uJmao6xKwnw0CWNMX70bQVJPtqMyH
jupMXqenSVYvBnf6RJfFwLV4OQdKzo6znfZkZdc7eZqBbUmDXDRLLy/DEjwoGrFH
Dg8shEdx92XYG0YrZq5TlttoJwjHY6vY+tW7taNfSModZIGAOLmQgKep5sFx0jBK
xD9xzrCHH3mgMjSWD9Ixdc/5T5as8lTcVvrBKYlvip5AjH5vhE+GUangz2Pw/fJX
YTRTfPBJ0WDZmNj4Jd8Ziuh/g8Nlkd+bJX9oRKJYDV3Y3tOBWBOUFN7nMVKXnYlV
Y7cllDZr5e3HGiXLkPuNS+UVN6CvRAygYYtrf7NBSIsZV4KWm7GIj9Nb1+om/mGA
ITB2N5yOonXM/VrdXgwbR0Z66x+osZbxD6l0V7oFW6m4LRgbJDDOi9SBLrPcLiSs
XoDZMYxalwj1EfqpyliA67IevPW99e6E16HTVe2rj3YS5Mrf19bU1PR9V/rzwZlT
mSnFwKo6OH8EgMTKuZW0iVqV7nNQggSG7TK4uvjWCjwq9YAH9TybsHUxoATn1zn0
wlLSHDZNJurmCXKO2+pXaTfbB1jTIoR4S8glj/rc673grgpxQK9p+A5nYJY1MCiw
b3H6E6VNiJFGFEZIit+MnPK+KU64xxKVdUyg7eby/i8use+GaSj24Kz6LBBxLEXU
vxBNXGypdCnO7dXyQ/r/o+BLfY9kLMrA3iuOFG6p0aBbSYNJNWN3Qo2VTeaGQL+J
XzuHwJK+5UxeTSuS69b0M8nHP+TBmJuDOMWBX8YNCNyLM0D/OZvmVnFb3Gf3ZyLs
KsTsgRi/b5O8qUDJq8sg7pSFHtMzICFE8naNFN/HRsDvI0mtf+WAh5oPmjwJcIt+
x7ZLxVa8XgIRpSiHgTM/zk0cZaSzG4xcOqk/fHkNR1KFNzoApjy+wbcmqbtfxIjj
XnWh1Tc5/bH8TcnT1JPXFU/a7jQOCqRD1JkrthdFP/1qI7NQ41Mzi9SGgWM1fb55
dICgXS9ujjTXtW/AKIXENN7J8+Cp2x28Mnwq6+092wbI5hAQQGnQrnClpS8cCZZ6
y73lUdIrfLrqi8VV10ftsG0piCIiRo5FaxhMOiLlIp0lrfjbChKfyOrJ9Pww6l8B
IEVD1LGTRSKHuEmiE7evBoA8c6GAMxuftz2Sf1i8vtWh9Zsqqlhga2RYYzAg6aKg
+lNB2tVi84kUUSG0pFYu/X6Uncw1chSim6cK4n7s4RoH2pfWeM7EwTFoEX+q0aGc
QX5KpnPnf+XnmC3j1Hrx+auzi2vNDXjNPGmPTFrlIhQsAIgx2QF1BMfZHzemjtrl
Y2FyijFJif/YDSO5N2A+Fr5KpILzQIAKsLFhVHpbZH+E7mJ9keFt/Wn9drlHCUmw
F9GbGo211x/VTGI44RkTDsTEbmvIdsOjFNoKKu22fwftmOBZUaV5KnB+HGJyUfqq
G1idHVVn8Cs74vEMNvwo35wtIx6H8OxiCKg6s1Yt4TqmI7LRhrM8TEUD2dHVubvL
huLM3ssLtLTeSJOnaiTQcQ9vmDebajecwfbS1qYxSwglBIK/yjGiHljikb486okg
iI3iGPCB+lPMbW+4B4xPHAIHW32Yep6BMynnvfFJ2pYEhAMH43E/bjCxkwXKMvz2
KTVF5VLAIVSolN29cU6BzS+F6umhALRQhXTt8x1PewTt9UsqNggVAjHQtMmO4UnU
gjo2/4esYJhgyOoSu1dq7ONJ1BoXTlsIsABij7dGFxucyoYhj9ek5ql/wWmaktJs
smoR36KZ6gIGGSofCSPNHWVajVSUTCURLZH6m3WaYFXFU7ieTWaCOf8agkXOH5JS
g7xOl6aYb0BAeRKoI8rTggZ8JO/enLoNzfLtI+QLjUQQFq4SSU0k/Uf4Je0jHirx
eSrRpF3xIXf25yargxYup6S7gu1h0bNt5dkcN7GDAeUNM9jR7sGI7RhhqtwGY7T/
he/6OFVQn1ydYkkFYI0x7Ct8qzmvAMDUd+iVEStXm9yLrqmLEw80TrHyUUHYq6IB
J0nnTmbtO1Y6FQ1tYpuUJqsc1OTAlfKTG/MRh+eiw94B8BVID21AvZvkDjDyiPYH
NbahwBt+uixs++9+OmiaSNwDukmP2rK/uIxjM+FEkMZxMHs9LFL9eIBGaUMJSdB8
jr/5trNivBTEIHeIR63rWNB2tzQbrEycxIDT4imCWSYqUafQNkJyWUVUcTgDYbJH
FkECUTrQklz1Bxt7IhT+diLw7+eC6g7+zbgdyxig6AQBQ+3qPreH11uR0Ch+t+U3
v0QmSIC4Yhg5536GoSSB437J92jsc3aFCkQK/n6vtaqxIPAsO/BNOoBFeTTP7H73
RelXguHyNJ+97XinCialkEAwTnmgGIP+slB6V0WXF8UG1dRCB6DGhDh5FpAG8XO3
fy7KWl8Ww1UYUyyuPddK4dsYgeAuA0ObEA1zItEOf+qb+//+ToxvVaMRM+NvhNki
9UMTmmpoKATOm2zBNsd7TGgFyHTMo11fgtPzmjCS8BHr1hisbCih0QYV/sWg8XXi
k4rXZ2cm461hn4jyH6pP2HLQ6QXoMpZgfP7AV8i6AM1iiR8B4vwShuJNby45TLQz
otxOwQejkt5B8lUeGSI4oplkKUTWMonyDyNESUD2M5SRr3ZBPmDbPOaftl//Nw3S
gPXWOn1kquj1o6E2bV28QwZdAQvS/ES8mzbhZujAiXk6R/b+AqhRXfBwlsurr5js
P/BtLdQ/1ipRuPoIMU0vL4mcwOqF9vItSvtARF8HDbODr+z4Fw4OGiIbX0pP0Esx
atqViEQLF1uJqR6aRztHXSJ92Mn0UhN0JcJ4aSGOZ05R2xouU1O6L8HeRzznOqnG
6hknYQ0rf0dxfT9moAZx9O6zVb8Do6JI93T1kGrzkNPpSCKY8mrsIOMOHXo8or63
aw6bmVlkGOFfk75ZFQWNhPFii+qTl+LyPnINHGCDaKSOFoe4wrtS4SL+jzT6FOvl
2q8Mo0QsCtcHxks2AO3c0yi0hMea3nhQ5HjjTPPs6dK/yX6M8UQzwX4/SAvLzzvv
uCW/8g3e/24FfBQ3N8Su/L7zL98yv6sVRuE4dlXgagSU+VgNYYKJyfQRLvIHaSrD
jMSo5W3KMwUXbFnG5KIJgC9sQMatzhskOobhxc/BO5yILOaofYA5zXPeTeObJmxz
zPdVUaXbyfTBMpK2nDHuMZRQ/Ng63J/KHqqVBe5AwnWlPsVpL+HiKRm4KsjJOeHg
yPZt9HAvv5ANniq8FHjuIsHBFGvlMhdwLaFaoCvNa+IN4bW2318KhjpI55tqcQ1t
SFzsKd2xVNAUTuFLaYejg2rDNFuUMtGRvOpdaQPDQNllnv1VMrCll9Omiy/8PohA
hBxhb5cx3SIteHnqx1L6dzse0/nHt1dSIUuAEp1z3bgJ3IyA5JLgG1ndPc3gYJ3l
vHaTbDpUK4jcXpfGuo1OabKLTpQptdvg4sRJnPR33KehUJcUL7NNqTVWwKrHeLlC
jDsG7/7aFhQQtUOzO9K+iUxIjlV1jp4tE79tNBVKLwx4UCHZfIDa9Ma68gxX+SAb
QTc26/pG+KKJrh0EqLpQ+Jz9XbRXi3ySzlXSwOg05cAXul9Dm9RolyvwhQ3pubhb
J7xzjP8OKNLYi7olUJ+5h2apxLyE8IatjbfImbBRUrDQWYcxwQdk4EbyaDwnyhTE
Z8Z81E3p/2JnokOqA1AfCJQvapYUQPE9dVJF7IY8PrALJfNoMrVLHPBKq2C6GZRt
+nG1hiULQubtcMq0kSDYRzxybyZq+UC3rR+o1WmNgYgw+v93U1HzQsOO1kLVXH+m
jiUWXWXbOe2V7nK5ix3peoxURRP71QwJlGXR5f3DNm2lBs/S72GSyvB/YjK7egcm
jfbUHUSPcwUHaWEpXLAqjMP9F8/+QtX6lsbNAfFo9OU5cIRXMoykg6faFz2kKyEl
9/GK3oywgGZQSn3+epNT3xBA0OmpittOCmLpiDXya6H+V3iyb2IzgojWN2l821I9
76+buRxSLWCfg8zXp3YGCAsG8fChhic0UuOUVdAlTNOHvo4xyWe3IvJqta/2/zK5
4lJlGEiFW4sn+9ZRsmalQBP4eqwhOSByOZci+RaTosYPsHlbBq0gLdlSxfoeTtZK
NO+Q63ytS2Fzee2CTj3n4j2IgrwYjUYnQcLjoz65sW0DsuPHCnPBP6p+tmlRrEOx
gOJHksaKtBRSlOrYkDq3ln/qxEuE0lFmkDsh60MclOOwTXgC6N+o8oB8+kubgl58
T6ee6Jr5uVv2kRyoQdBMpxLutFwvrukBNZ6KOSfpfWxw18aMdeq2rJi227qJTGIZ
aDbBPOopp/kLwnXytzySN6VBqPkUg0YyH2f4HnjHGF0b09ObZpXzkNLImwdovrM5
RkYDGch6ZMhDrA2afQONPAAOfnE0bpeDnVacebibRELzGgEaQiHS+A+uUTbFpDYp
6xv96Zej6A07y/aVPTAkLuaxgw2TfbgO82W7MaATE61qjijIVj75tXheY4yteR75
Orgl3PXyhm+mRB47divI4j5HajqFnwOAdIg1VXg3ulLbj+Befbs6RySG/ELtXto6
LZcTv/nJaUUbxtrc2VOnhrICtYQRXCkflEbsGgsU70B+XltflCstAhPtL3cXPHJu
zN0aMHK2m/XCIr/+aAr/ktoKYAZZ8gVpHXhmpHl/DAeblpp41euB144rrhm4MD8p
gnI6bxnsy+Cwcs0FPVSHFm6/02n5fv8wvj48M3ORQJOIJJx+wCyGvWiAQIkDt3Ci
yIUrzGX9G2rm0D1z5HNOlY9eKzsEtdwdkZCNycWsWIuhIZpPvvgOVmTqCQ2TzMx1
VmFGwPKlPLC2/PCBPgOEypWRYcOpBCKXlPFk25jMQV0i0fpad+79xPs6iUHktAqw
zggz/HB/Xoajf9YssQVfGU7hVzcqudLvmzr9J7/tZhgnzFsEllOUYHPeLmWrSoQF
mzH64wLVarp25VJNSuT3HCsxYn1KR6nnNxKZUbWh21GNTxByCr2760jN6oQEA3MV
Bo83JKobFVAvBuD3GTUV2zGo69wNSihBGoq4ZvJlBI1e516oJFA2O0vJformWOPV
g0WLBy3Z2fYfCGvzQK1NXB4ihS3Vwot8JRAGzMxXGhkmVAwzh4ZkrmqTIvCM3Wdy
0tPMrTnSm28nZoXfG+4AwEbyTlh2+eeJy9S21BsW55OnYJNEy3A7u0ukKd46tiSm
lmn6woEG2z7+lq6HxKUHpCO+Kfb8pY/d6NQ74zTeluCsvXmj70Uwv7XIASS+Ln/o
av3wKkfPicg6IqgHP1/iM9DFkPIMvByfWHZcd7yNH9xws2yj841Rd7CezImUZBB+
7MYjeDuXcFb0DxpvP74C8TxQ4ysHB00WyCezuzmsVCCtrKn8q3+Dh09MV0B+tW4F
sN1LPOUPdxSqHI128bP9lLT4BIvlepBNCJJvQoZiiliUV6A+BimgcEdN3X0g0/0I
3k/gM3wP+utBLbrdzCiw9WRKHsdCAal/IX8wwDK9M6iClIA5n9UN3EASaLwAONxC
fI16gUGTmyAe1fxzYbsspgAZ854oDOcSSX0DNK9jD51OdcZCWfJi8eTUb/jH0L9Y
xlgQehelCkZfpoPESlkK9KMNcL+TGjrRCwAy4pk4ZhIw06XaAZyFJ6zWeS/vmgsN
TD6dWWRbEuTKzWlJ5uZgWeMFJNpPNyHXqYRNYTiRgJWB9l9TifM262wqI/pV+Rzl
jh49Wj2XfLjIwdfCKLrC+qRaaXDk83ELBjlaGpJCkmZuGdzEMdEVLiW6ks9+tpPW
T+AGy/XMKPdXfVUs4IZ4SZsEtSOggbyGLh5GspjXLfdL+9ZzUl73A1hiMXPgvyTA
eI/tzahFd/DQlSYe/C50kiABZ2xrAIhWnNpplTAxMMklxkgdO13TTE+llk623bgN
hC/iEXznSXH+xFDJWvr04R4AAmtBCt+6RrBOWCmZOIyhXw7YLWncDXJAN8gAF6CS
womkEuvmLGKzpcmaq6nClXXpKy5oviislt4Ga+OMDXe8XGhIZZ29S16fqN5WpvgB
7A055EA+RnbTNt4Nb0RhC+vy1YNcUOvXVsUqfaLTF8urn63EzB/CpC39tx6900sU
ZsXou1gSLoNdmfJRdGmVUCyjbZz8GZ+2Gy7mk0gJJbE9o6KmWCRUZMwGzOGjU7H2
trkgs8amMwdBsB4oxDmxgGvqKKwMhku1KrKxZOkASnBHjLPVFYjvaPePrFBDeIAe
/BgHDygajpdpPbdtC8Bon3f51pgRRGdH13wGBjUFREdbWuP7n9165DgWRq/4nTyb
SzYJrBvav6WCcIw8emAcXsyD3gG+x/4QJKqQRm96v09TPctArvXi1zFD15bzuEDO
LypEeNKRDxH0iVvb+9Xj9Y9OollpEmOv894MzC7xelQni/MDYo0GATRZRiyteriu
svNj5DFerutpatleNaaD/cg6FTn9rCQykd+L8AshFFeaK5JodeD9p2/1cyV8qAgt
awLa3XTEbNafoGFLtriDRscbXZT3ICGRpL3Ri1yM19bvje0UEvmPH4eqdhWADNi8
rVb4A0vNjVS/byBl1aASXzp1eNwzupAXKTHQWePmqwsvibPnZHffuq/mmeohQKcQ
o/F500k0IIxa0nwGN7G/cWFeXZ391j/0hiLusLSqK4+vCCPxxXg1lMtQFuS8dnu7
NRvVZWllpOWKbF15MgbFZfI/T/U4SsimxBqBP6iO8OqY3M+oKdmXEliXqphL6+U5
9MRf8f38XAtZvWyNugJKIfiZfhTrsi4SLIF0LUQMMqERttVVLMnWs0y/rRYIY8RN
9IwEXi9UrxOU4hWWyz47vOFacGWXEVXaXRz7Y2ohe59rA3S2rPR8vNcikg6fUcNs
wUeDNTb/VLfpG+3V/BJAVbiC776+4n28wWl6iyBABbNdoR3Dw/UsO9KDaS3a1b1T
0fLSDAiDGA7VnV2fKhnNgX4oqpYUIxsdH2YyBB+V026KlFUppV03K1ixDr4cIRFc
s1PpB5MWPD2c7fLq1MTrSYDdNQmYgEEiGPvC0cC70xPC9z8+B24x/S6q5Vzs6sl3
IMKXrWOTU0IFTkKNrgK6ghtcBKXKxNaB7LLsqbsOrAzabgDMPc/BqPNhY/hLclPI
nHygIhW3YeXCxA6gLarzASn4lwB5yTlAivne0TClVIw3fPKvPJy8gWSYxATehguF
QzsQCzV1oL0onHJ0+iMgKiUv492kFQiz42rdckfCF9A41zBRk/29x7zTbF5NP63c
D4BO8TPyGBr8phWU94hwbAkr5i/NDTrZJxKF36ADcqZPZgqb+Er/0iBFhRbuIjha
Ev851NJftxNjLELe3QxmYAQpgiinD5Ulii2XsqhoQBOKUxz5m3o6J9KlBoCKiNCL
id5ZOhvkDmrwYCVMsT8sjeviOZf3acxm5zeb1ztlaVOaI+RknArCEHtk1SZ/1es4
AKIOXK6AEuMu40Mx7wn1oa4/Elki2OuXk7xAaQAD/UesJ+sRC/AJYbSzWp7zQeSz
I+8Saio03cRTcUx43bRWgamDAuhOPujVsOMK3gaCHfJfh1U4K2+RCMMrmTorzp7T
85Aznr9ypDJQYB8Ge1psNnwigROx6wEYMUPEIzGjyqqiqt7kYKcKdvQ12KyENv+z
bUT7wXBy4QWtWUv3SD0u94A9oVHZx3p7nDUhsmlQz84l2qjVGfm8/FVsTRjO+Yyu
dxXX25aOlwiRie/v69RoJzmDABT2hX8bIMoAhr9jv4Yc5tIDFoDf+ioNvTEKWz90
PEEgqeS2kgjn3V8Aq/1I4jsH9O6uLg607uWkkJDW59Obe4ZvZbH4I22X2c45o5Ob
U25Mm1yaLycSEtBSJ09fjy6qPeGUa8+0MANQd6BG3EfDtVOzyWa2SBBZE9vgGAzS
gGGuALxiXXEzDcMI25ijMQXGiDsl+vgiNsYboy3OsyY/kT1Z5uscHaX8/IZZgBR4
I4I6tPfcgIoXugLfZDArT1qVy0HmAyxae+eJTtE8OVRtOWZsiEWdTgHBi3rXiDa8
h1ijYfF282X+AC6dwSRb/LwiFJf7hpbLug3nIQNSGr1l8DVWDlzPAQ5PE5KBndot
j90efyDuxE2ueIBLDUIXBRI/PPJksIacRFdkqlAbnrzcw0QWfqVPx4DKxfcC1KN6
tAPjPV76WUJywyC3AvixoIpKA93AVGfAq56/7LhueoocrXQDgG6tQdOti899EODl
YyZVBzLQ++6oR421EdYw0FfaBz9XglrhPw6WsmCqk4QUeSH69NSga0FS097ZV7QW
yc9D+7WE7h7Gg39HDR+Ruax35qASXhu1wyoSrsvs4+BLucTw5jgwWS8Ld4+s/mDb
LtY3Iw7SCyGqaFkTzOQKxVLM7AYpcTbz6RUwJW8LAccZGeRGtWoWIyJJVLfoI+s3
Qw0sp9pNfUHqE0Wa12nE5CY6VqOjFp/CRHOx1BuZo9nxVX2oSFy6uXszL92TiSLQ
OsrFoJFMyEo/eeSIKySe2Or4Cr4ydyU180JXGiwbrDB4UhRIdEOac25luqlllOgR
vbYph8jBzYRQZqiiNfBmNOdRh9r5L8f7AXWKJs9Ww6N6sa1qgAjDo42WxTvFrDw0
xJfrYyGPGwWOzf7MtXYMjd0gfzjla58ZWd6uSb8Vg1lrQ4UUDH1EIz4uSAa5/HAe
XWu6b5C4TirEliIL5Noj4RUOT9DgApIKKPcRz2CZhofv2cuzWtpdHQp1GPm81d/2
9/kKkflVdX0maIBSu8GvnCCRv2UBtDcwDnsFakUxvzcL2lxBDrM3r3IZDwfYq6MJ
Yq4bEf1eULMAmG7npXxy/mE63zMUKZorj5lDyPxMQb6e6YnGEA4Ps/15rLqvdJE6
NcXBakPhiHpeS7Ko4uX1EuKdy+hl6ZnNXK7vDKAabajakFsWGAZAT6DK/SRn3Q93
WiTQiqlobVmDjji81FQcl22e/gaVxZ/gkxLYaYt0H2JnTPeJLjNAxTW2Lnfho6hx
JbqGBtpi2VQZ3qg3DWD4TIx+Wyz3l78Ux1JCUg7frSMkVStCyboPFeOUXZGFfewg
0MSDpD16TxM4Z4rmvaaotS5bR32OfwwhDp19Hm65AENJCnQXAwwKAMnjA4UGOEyo
cH9xrRP6vtkc+PvkCOA8tKBCngeimRV6Q+ilTyDpl6Dr3losVFti0mqy1hVahydN
Nso0uAKHRhCgE56RJAk+wbH0UUsr96Ht2BkKrUVYNDv2a35wghoLuGUI9R4LqL9B
dLrvPFt4DVp0A2vxC/i5TSkLq/FRojiDGSoDkuhDX94AKJuHWcLRvdSL0cNuwqhC
/qp0t1jAeg+bSYoWzBk8gT5QKEaCmeGWIFQKF/SBj9eYvW35kiHbvsHsPsaa8XIR
nQhSYL4380mHzNmli218CLQnW39WduW5HYVjX0INkD7L4Si58W7i1aeHbywSkubf
0pi9QCPF/Rh558hn/UkwSYtH/GZ2aRw/KHFMrOPpN55rHlnf/ioxnoYNQYRDgkM8
Kqfs6Ul/R5+LdQyTFZM5TYIOx5oqracQ0vmNjg7n4LOLQu/FscQ9lXjdjTew1Ume
xhBmYOPAln8/To9MFeeXc269mryBdHxpXpARt6np8fHya0c6VPfoj4+/18rdPert
yHBJr0C4me1daZ5OQYbHfK7ckwjn7RHQXtZ+amuf1kzz0CqrkBC73zmW8PkzDfM/
EDrfHGiuTnXlds2Y3KBaFkdRdJXPpOFGHY3l+9RXLQEJ58qzEAMM+mOL687ZinuW
tYV8TIlyegDDNNOel0BleusU3fZq8BLWpuwQLoOahlbGqa7rJTe05ai8DWyzcQUn
PrmvDt5Mj5qexHQN81WzrbTeiqtnlosP58baXyQ7QF2IsaUScu+OaIZeku+Ih8Eo
1FU9KISVyhozflPU7mIU5klTnkk4vlwIYX33059AsCDzJFKJcWHmE6W00eVXh9yd
3ie9KWfp8dthGRySiayYQU87OPHnmv/iLDfYm36NMYg21V7+0OyNDdPc8o6xFR+Z
1meSI7jzvpsslrmQRPXTx2isPSL/ELgNEbP/8YYCAQZUKHQx0+Q1x4QhOT3/bGlM
b6+RZQKoAMDJUoeID5BPg/mN1TdyT5NdrwR9T2M9vT17VCM7tAu2jVSMBjMH6Gv5
QGqdA23Z5tPMpMBXm1E/cEAMOiQSOctzdaW1ShSHrMQ5lJwm/g2Ca2Wfmgm4Dg/u
Lg2j1uaW7JrUn3diKc3tsA0jhGqdesjZaNPkZgZqu1Vbwy+vQtZsKut2N+EvKzVA
HKly2Uy7qgcHLCNvk4d9YTky+7crYrZVANmIuG8x7GBd93Og3A9nXibqstzwYUaE
l6ne0UyvK0k40j9Yysw5HhftpYDhj8C9lzwiuixTixfRB/eqgzTU7SDx8Dik+LW4
AqizrKSh3yC0f/pBzCP4qpfSrx/K0TO//QByGnhUOptyCvFrt3Eyijs2XVq0nQaV
bmcrvXJvvqOhTmuKC4HjALojGaRTog56FtJbsPHbl+a+i184eykVRkIty2beD951
7t065780ijQD67B34sxjCZ+KjLHfF/FtBlzPixvgDjG9q10JLlkXU7l2pqBX19ch
/kuW2y2lJPUTgxXeTzXXR5BrS4BGzRfAsEjYtHzlmKJiuAHvkLb8I91cLKeT/sLt
u7lfZmi/Yid0OtQ+DD6CbPcMLLEJ93OqmEUjvt+tC5dtjCi4vd4gGsywUqGM4zic
zcKVJSLVPySJvmrV+ncEqJC50pEJFcJgBFGwfWSr+FgSOANdh/1IlsHnwlFQGX15
zZtz5jZy9J9/5tUjC/WUSR3VqaLZbJUscqr5WiWuQTWzE4OxTQgVqxqyqdKxsbzI
ov7R4NizsxorhDRgym60opcwKSk/wPYlNDSQHE7jVO5LjEuV5m6MAXU2kzGUD3tF
syaCvk1iyKwv20NJrOTyp545hkzZJnfPYz3UmzpSY3sV8lwZwduaBmoGiTw1UxkB
4e9CchCKqt/xi6hHvv5DhvxSXiDD46M6n9W8JOilose8FcU0u+0mv8vhkma+oVxm
yzy+gJhIqZh1VjDnhealw3NX8tmA/e8Me7JHlb7AvPDdYWWylOFUjffM+qcPQm9r
SkUjqL65s/9COLzstsfe1ZDPJ3JylE68Eqj6J/zUouAovbr+LFzlpImBhsYyweGz
1jpAfHGqRx2IpuEOcs1Y4KT6WiQ4Jyl9wTu7fZd8jYSX1EH7U7skccm2agV2uojp
XwPQpV4x9kj5cpsCdg3+crxHtbP648QFNH3ZnG7Vssmu0niE/BSIH2pVkkxQYWZw
FLzampnC6pjyD97S/o0rFGJ9GiojJHoufj/wFI0PO/jZbr6kiArdOLVB/Xz/sRC2
bLEkT3nopJOys8P9iQfk5mjniRHJKC3Qvb8SIJ0JQNR2KM2tF7FLGEbPghY4TOzw
aIqiJmcFLLpc2SpbsqyfcuBCYD/tQBs4VBnmzYVE94wKIwj/WTWh3lDEnlVjVLkE
TixkEpMi84ROVYXPk5bMUoJ21ccBCSsO2zvXVoOWL73A+Sj8HbaNHwZs2uoqOC3O
XEcSCYS9+4bC80kPHhK5TZgOuznQpi+AtQibNEBZyClqs2d/m1O+Gq7HEI6Y16Qo
hArH4Edrhff5eX5wIk8GGumTZErGa7/hQd4LKAI8pi/pexDs+/GvNq3YiWDyX/WW
NaaTdzLPg5wW6CSDeaPLHHlCbgcs9una6jW0LrzJatlxVjv1UZN02m8+z9+crPyn
XPRvgRRsggGB7K27OIhxe4eKFr+Maxzm3mDuy75EIeJ+EA427QtpX6trKwIudcBF
6pOVektmP7R/jXIBQUbru8Q4UDhZiRd9lfCSP6Jj3pwlp451UQQ0SOJrC94qYYoZ
of4Tz1pKehNORa8bT1EIxXvGZBrJXanTJ1lyEI2q7RRCriLiYvB8icoWMo2e0Nlf
VYMXJfyJNDp3LhIDErT7YIsdmtklcCOSZoqwPDDdvXMyfj+jxKRlxaiRzXLW1lWN
aEuDaUFWy6v9UyuHIVBeIZzo3lLeAvGPz9abIigusoBvZ4vJC8HZwaLXgM+Yk42G
hOBAEXG2n7Gbni4qSj0+2Y3DaMu7Anem8Dc36j3jGTailHltSojhWhTHk/HNApg6
6nzGLvI62QYySTxtp7YfBUb90GG7frI12irpClsksDZV4sS1AqmG6mfxH/eIu4us
pxLSUu6A5tvF5Lm6JvpajAaiPIlK04hTgOHfOaKfJYwbS6WctEqXxoSIYFsTCKW7
kUysD+iV2n4Ue3/FE/Ku8TdPmmILSi7a6pdRP0Q7ACpRnci+dyH38HEfO+dwB2n8
kKGy5VHulQEL9jTk1XAZ5ytxnwJlHaYP/FFrcRB+aiWIFzMj8Mrm/wSLdrua/4Ly
gAMHR58pQh+oXXyE3sDoZ9eIjZZJotb0mt3mtb5nkPv2R0x/LTkYF8fdXTekv2G4
p5J7dtpgs3yn9A1WWQH780H7nd6zcUehNnJOuaBIe6HyIPZF46P3g0TTm5oA/lxg
KhFutu3FBrvV9/d2z00xVK/ECZXcGChq0mkSUNns3iAui5XwxcdcJVHcwK1RX4tI
ZaEJ7jiXfe1GzXu+7cwbyl+JHrZ60pgdkdlsmx/oaFPYTUzCalMkz0daVrIRl8dO
o6gBwzuWak/0qlyP9fAdeT2+Ubt0j3wynmcppK0XPxRki2swE02Rn5TBt7jY2Qbb
aO+W9AV304Od0GlBPyLiGkeXTeTkczzvV+DB+q/lV9krwGIvw9HDWQSb/2eTw6mF
bx3RibU5WYHvs+nt4C3Zb1QgF496kQVXYPQyXY6Ii+mBnPVHkegOMxaXzSueUOoo
KzR9wUkg//ek41RidDqHGlua5Xi92R5UAh56dRh7PwWYrDhmICncOkeJojUUVVq9
tOrGzbgm20i+Je/iXJrgVPBOtL2YqqwV0LZPv7FtZWXy6P2mhhIsNQyTjmwwlJk6
DypCdjPC1exWkVbuBPLm2yb1jBkgN7UcYW5X+mvZA8zd3B/vvEXQJbSV9DVqsNkx
YKSM+syssHFdq2qC3jR/odeedZ1/FcqdcyhMYPTelwE3bKlI/K251wXIMAmLFm5a
XZUXR4P+HU/b/GxqJ4H3EhERmssEMXwUJHU3WWs/wV1cswwGONDBjONhqrkqtcmW
THPNIJ7+8STy4V2XBhjCsfPCA0jgCEUjUadwwCrXAzIApV4oi5itJYaIbl2iCdIh
ur3mE+ZZoCeknZ8bn1FDMR2DMgZo91T+jI0//ZNkj4bb8WIrUmRB6ZgQ2HBM2WVo
amOlavUGx9TdV31iNZ8cFasieSu/Zo5hsNc/Ot5WLThGHMJ8a8Swv3o+941vfjmr
RLnOpHox0/8YfYKg4FDsbSBpeu0ctQ1zFVZ86FXUp/yqQb4kM7iXM+CEim8vdRHZ
sCnLB788OBHKt/bnlTi1uPAvbcFy0RUosNAfSDRQasBjm0pR+1HclhB6Rz4WsqMw
rSuq593OzQ/K/luJ+fZmkXthrqfkeXFZbMbQO1B1UtisJN37sfIHiN4NCg/jVnij
lLLUT1BpfJYmDAoOXQl9yPJ4tf+po6tF2j2DjnaKuR09cz/O/dYDH7udgov/+OGU
ihDdJvD8nTxnFWTfvRwbxH05ZMwDPykO1YMJSqC8h7bYwT7ld/CaFP8LlUhCUwhU
fvhmE3T/9WkvdwFozmkeHvKFCM7GGwsNf2bIEQOlv31Xj4cyVjvCKwH3s8f5pprP
Fy2RSfstZMtvqhg4E+CZA0ypj1w5MaDGu3P0Stfgg3bFx3L/VrOAYanrMZHK4D2J
3ONiS4hTteSjSBgVk7MK685Ts0Fj3pWaDt57PQWgMqZgVtEptNexwvLKxcYrCtNB
L2u2grmqLtNhWTitHlNdqiE1D9wdnwCMhbPCg9q2TLaKWTrvt7ZsnGpVnZRuAhQd
kFMosYx5hZgE2BVHvYDv7tCMq+rYISd/o3eLcZd4J8uJRI2t5ldP3YpsfUycLi4A
Zrd2dcavhFQoBPgAcfBF/C9MZEWzoDQzzmHP2HShBbNzKagPS3HQlXJpq5m6TEGl
oiqrFxxu53IdWl+6ztS5kWu69w+/+Je6vmwj61CayI32MO2JdtfbpPMzdEyDtmFj
pa9/9dDSCF14WW/fnx5jPw4bOH8KgSSR/xKaXyQpeQ4NfOiVVtzLWGOhyVPYjQbT
pRmr6DE9ulp9gVT2zvAdn99mjXEUf8gli+dvFfxaiUYLsk1MXjJYc+eURFN37+W8
Snv/kDqM4pheT6M63+XZrB67+icBjCj9RwB/A6NhccTlD4w3A2eXmr0fE1IhaEUC
M4Zy4pVMZlvAHz2LmB/KHi7wBox0/PQKoiB9J+aAuaMXvfEsB1VJR+GJtoG8J5Em
jRqymYCeNaUq2vrnBW7tsPsi641Hfe0qL8xv+wrNMqeiA/aFQH69JmFlox+8xsvf
678BzcfITq7yNyBmi8oIFrkFKluUXpnHa+oOx9mwkBjN7hNVn7z0bwZnMw4sRZkj
JLGqvhgNQEizWUozDnNIFmnaZo4cjCT5TNLjApja5RAyr8QuYYRdPeXQyXuzPmhO
wJ/YRZg4uQ+EBhcHQTISUjgv+RmyAIdh1v3MjYEDHmIaFviLr0Bu/ZRnMozBVy73
NunFPhRwNilR5Gw//8u9gj5x6y4LhPHqKnDdp4aThlF5NBZ6Oxsfdw0LSLGufV4Z
/mIYULttEorAfjD+evjGyPzfPcoAvO+ft7tBVb5oL4OuQdXaCAtNIEn/vX2WKMtk
SlcxExWhQRXdmanQ46SbAUX5Po/Vr7ZoxuaBlCKFaECgg2DZbP8dH9ZH9ModKN5p
Chb+QBqmNiK0q32K+Y6aSe59ekOT8AuXbKe6LdAvHwJl0UotlVTStGEgDpRf+vpX
xUZ8qZhfRIxpI11DvDtn1WRuaSOyT5CGEeHE0V4aTpWlEtRctTnq4Ka7K90/D++K
eK/Cmy/VQbpVMV3IgdkT8EY5fXFt6AZsxLXqpd53Ub352g5GrS/fvsRlJyjxkW+M
A3j82iNwj2nm4s9Sz8XHUIi/ILjLfAuj94HywZnkUNGDNfVY6ZSF85gaZk+L0CZb
4039lyXZOFRjpVz3O03KyS7g1idWLwX5Ug2Nz79iR17kgbRoVcRh+cIw2EtQ34Gy
dNb8pOwTr47O6xrqGEorGSH1xay3VLFWlsbwL9BhzSGcndyhOo7KG3CfjmVKHiYq
TZKDlW0vkP/n5XLS5VExPfbkGGubUMZLsey9VEFlu8jXXS9d6zTKnWMbLzNrBT2Z
0XAeJkSBZPcxowmNje4KtX0E/KapXne4L9n4bmbw2B4GeyNWKOeTFAR9aLAnXYh6
UiMLq94vmHmAEaj6QU/ZxH0B1XEDvIwY36l3jjev4GLkFf4YhC0EsvR6PCkRwX/s
QsT3iXkDmZD+Fuy1K3lUbFimrz0Q8YYPl0eSdCjLPuDqPOajc4LGl1VM4iDkNu1u
j+sQO9mbSf51fZ5+hJLdenZK/jvqM7uWG2hSYV15OFlZiaC9pj9KEPqRpqx2knBq
eFoVzpSVICI6rib62BehOctwWAuuiM3ME/kKVMgqv/f12P16FMuP4P+k9JIwvQA/
Lzc3eMEAs6kspIFXT42/3ZWespP3JlAnmmH/jIQeVZgOi/+TpLEKiRoALOmCcaUa
GgEPy5+/JU6qwpIIRYE2pGrKmUaVvD5Szs/TCNWxn23gC2zvzc3PzZJNB/nh/k59
GgRB8ARI4P09J97qnEMQS7HJiGITvx1uuD4dlO5teH9DnkB4QlDzqNIhYYVfPlXb
ND60VHLGzwe6rVoYced8T5SvNA4fXMj9vmX7benC6gY6SMHl/mFGYpnRSuM2C4Ik
o+ikDvkyTLWUlUYCUI6F5qIvFY8lbjkTAESTmoZQzT4gxEP9ul3bWd072+kmyrTS
rBbFofExI7NCHzpNNkiokGqZpNlL4MG6yp7RxUXRslTo5ToGSHKLhzGbLnOQLqn+
GT0FGUcOkApQHh+1zofX0ssWbgU0gNBj7AdGLYwrEsxNvbtudNbu6nIiAjqCqWRX
8w00XroU2kEtBxPQzc2T4sBxIU1oufZ0iXDmZkB9kTdNKx5CkNOXQl5VpNetqD4h
wnnOLookDC9Rr1PDKEumS9BOqDw1YadUp/9CcOHt/e7vWqissTzmRDEs/FcrTUQP
QcPwg/JRfQwuU2jQKD4hHexY6GlyN1K27sun8+NP6yzgX6CbBd62Jg1VOAfdqEJ2
p+9WenQGUbGK2/rntkVRSTlsT9L1zmz2D0PDRKH9OIyBfljVFMmWja/DrWgjB53k
bEh3cyWrayis9u5FTQARp/mRLagp5I3+DJ+pj47dnqRmzIc7iCRvPZZb/huFROtI
0+mPE7VSw2DXZkQw8YrRmQOTfMHYv7amVhiYFZVpUNaTQfxQ7fA9+/RKAThNu+NU
18XOxsPqdPKYlV621whBXHVPWEAxBOPvfcWt47/Gzj25geel+L46ybSygHgUC2s9
9mOFbKwBwOvLO5Njb8bSQiCt+3cHSQKhxlPofqs4h7hlzP/duWY8AtRQr9kLyvdv
p+fpWQKuP+Xz8+3gFzZv3cHhXS7XNfnG8n3eB8TGL76eRNSg41DOK9vyb8J86TvY
6PUon92BXP6RNcLNM6bDpK0ePxxPGo+F+vaG4U3iH4vU38uktg1tqNN64pU/Tm1t
bUuWGQ6ofAMvjyBNcapbzufuSy94CHykS7d3kTxbP9EiU1ub+CjK3w6NHVagWqA+
rJ0f9nOaiol/1ja+ZO4KSdXQzDKu32GvBzgAYyZCHzJB+wLqofaRG79cEjVoYZ+D
fmvw7MOxg6LLyCkZVtD4FkTdFo8axT0nRw53lu2bYah+4+q3bseO6hk35IJn4/A4
kxzzgQvqPKEL5CAuXW0i4XTXAAvrlLVguRPmo+qmQLxVhT77OrcEcgJqWAbhF7SV
skMvItnyAra/+5N6AwY6WxltiAszjeEC7WEIMkKVLswupTZvZNQ7QXsO4lm/OItO
xwDajCxbsZbFYxhbXAcBvLPqqA9kwmT9ZWajAlUEL0oX6FH+VPv9+1JXHhquOMdY
vlUPbaGsfXOwmEzmeZEbxIM/RkkxjY5e/6Ck/gXfbRa6C/GbZ03TPlzL+8ajEspT
W3elWHgulaGXrx/5hyyWUlaEUHWqDVhUoGxih1yiDbKDMDjkRbrKPjY5EEfovRzg
rHEMjdS0s+ClAv+bj+nwb0LjwCRKgG4dOzRbrgqLgF7LkfhNZZksLe2WptZ3Tr4I
r69k8yjLJQbryCSEpewhsgeRXmPA9nahG6ZDFfTVc3cUdJPuaJhRdiJdbFPIVaCa
nZgJgCUMrm8l+OnKcxxk5VtACCbgxq0PBoC5vhdJjgHSFvviM+DYbz6HxfEqaosq
uAIbw2SnJg18FftRoKuuQFx9mYL2qQGRWCp4aYIQUN0tCu0wkz8k04tR19HZd0IJ
nPPSKNijl4KAiYuyCR/JRif1c/W4nRAdcgDS43vWyBVP+mldd8I9ezEoM+67ZgHb
ieyV7UM3pxXwjn8yWgBi4NW87/veSDSPqoKZ5XJSNm7Rl/YKMKFxWWpgoRsCFllE
V8KLVgX+MwKCNno2LDagvsKFaBStRzNHoijeS6jftqATnbr1js5HDOtn6acc4mU5
9ziAtTCFnyg0UXpjIR0FjJYkthTSIvKdDEgFbUZ9BKDEymq455R5liAzH5j6l5Vk
Y3X8pY+uZh5pBMsQixLgvEjcaXw34fJb7MAGah6dmlAaj8qjsn4emjsXwEMJUcXC
/W30okwyPsUmd4va3djwGEIZjhQ9MdMBUcTzHsU+lB96JV2Xo0Fdr5Atf1P5jSC3
sI9Y6i3iu1DjrKR3Oys8Vf5S62O8VMups4IlmsTkvpJEdP9qPHVJff+U6J6x6v0A
IA8VSGkjYzpW8GKyWQwI1NjXI/xOrnIfE1ZMoI2LYQh3Vr69qJMwZz4rIbUzZPFx
Z17bL03rsQ8yzKg2/ttE1mAXSRHLaMVhb8l3STb8qzR7U1ywC7FMTVyr0l0i5rF1
ZmCl6l6bpWkkK2Rgb9NYeH2gPTxa3xxL/4ZxwQFXXlInCzCUf0rCAcQ2Gy5ot448
MxrWsRUYlpaJYo6Qm/IWFgU4i6iskGCChqK+5la60T8pil12RfcWOci+cSxmfDvK
oz1x7TI65YLU9zm9pwnqqk7VoskdQxA49699/eRumRGplT9dVVEvQte3hWkWOV7D
70k5trKgVzMxtZ3d7gxIhAu3opqQ4x3Dzm5FQsf85x8Sqkbr7i9ziBg7hU8TfmSC
gj+zuv5q5BDrePkX/jFhioHp4DjaUKffU014bJkChVSSkWhD6tlYkNKwKxr90uIb
aUmCPOraQvaNPORei0tVk3syUztgFny3ypnxcVuFTXnncDTfn4vlnAkunuUPnCNQ
768Z1+0VUk/vcItP/lAmmy9zr9JXLeLx9Zoir7Ah/B0SaHyNYaygKX6lsH1sPykv
aCIDmwvYohJLo/eWXuzi1zD6CixoW6M+DMZgvRofPhjhWUzPo+0db0bYEodTbQdI
KAtKv1Wx61DRf6FNVDC7KpRCOwKnO1wnZ3Axm3CexNU5ibvJez9rYb6jFwzfr1ZA
0Tv21zi/kJ1WWexwFB+m0K0g/qQRPTuwY661PK/V7Yx3h353fNVgQ17FbdqtwY1V
i55uSYZ1ZyqNJ9Xr3q/x2gru3buT9cRbP0dN1+5LO4rbI9aqIpbzut7XH0A5Yp5C
WcN3H8UlQuZx6rd0cUsRUjiUimEajCDsCRqZZqnb6MT0C2fZhvImhqLZKeUa/WzU
dn9I5b8eVH7iTl5KbfGmLn0nINC1D7j3eGyGfoYKc4POPQRPm5dQcihgKzXbdRN/
wjHgUid4EVWDQuS7nJCW+CYtXVxweML5pWWA7Dactg2KEP9T0e1EGza6PC8a4OhS
0Tapo7mgamjK4aUcAL1MmhbOtEZ3975UyggJrgiR28VTH1KSFMPJg59ytXq9vQHg
uNpdvBJjok8DbK72DTu1tEad3MiBOsO4vuf/uQ0cpFBE5CGa1VKpggfcpbxroaZU
1nhpCZB6vLfZbSc7rf+3g2883rsC5lddbTk6ZkEaXh8U5sXfICobYKhnQAVyiYkH
/UyxiViWjDw8Es7awfvPHCj/OBw1Rq/V8jKibS1csb/pszHLR9uwXPkQuMXeirVX
wYpSIpKAaZKN9dbewrCOrTjc4ap1Ib6PKXvpfvtIiHQ1DI9EOS5q1vNNplDCBQlb
KFxbVXq+3+MkT4IH37VkiMGiX88kXRwrFbr/KVaiWgS7aDj0w4BkxMg+hLIbUvcl
khqO9b3YRrDAtsBB2OhbYBsnfXdlaqNJAb17ljKEt9FqDheaQ7xaCZ5NUeD935X6
sMQbjFEIcU8DohzLZSkprmUPHwHHGvkO2TZNvhZdGTnlyyx4g/74BpPT3KeRwaG2
wPJWAsu3zbKmFLx0in8PxpIpa3ETm13lZhxJ6qA9et7qcR+1jMu0Z3ax7gw/COIk
QnB99+uF7cYFUX2hV0t4rh5GixH7ta04YndEq4W/7yiVqLSz9xXLUAz9kf//oisr
OOoQ2kL1Uz/zeefiKTSsBsnmy+7WQ46iLaktGT/myA0tRFW5L1yPg3gSBOyLhn6d
OEBD4uedF80C3HD7dkmP7JrtxzFl5raswbsxebS/bF4+EzLgG8OSkDgZOVIfM7Mj
yeA9qeyBOwcFJ1whyhcKJbNHhIv0Ox6k2YVYs8QTaXPrr/5gjzEG7iNCLFPtyAfg
HBZLoElsOEnGCpxj5AywGDaGQfLyWC1j6xKRggjzuXWY0hUUMwfN026vNUjY/VZl
Q6SURlUCUci96iW1gi1/0xz7EWbp5St/K3ofie0ieFJM28ex0ppKAx3NAN6ssFsB
EMbOPcB7+Flt4No58BH06Zo+M5ycLSaOsI8dLkNn39e4BigrwEOSIR/EmUdqum//
Orzx52NC35fCoiUo1FfmdLHV7X6JfYA2AUKP6lOCyDmmdxYBmSaQucdcJW589n1h
YMArLmmy8kttnNTQ5mM+iW8KoRHW5QZo7n79SjWZvZmhQEpRiVt/cSzlbtxB1NBh
rd+60VJUWxl4CNVbegfw6ziruq9l0Rc34zbmWisc2ZX+LlUre48ywVKyiCbCf768
bUn0en3PBF7FDo3WG7bxTvbtgOuenGohADxLbU2v26gQbxqlzkyFSexBjE4thXUh
WZbynMDmArmNcE7fvtg4CoHB6UfN081tHUE4YovtrJvp9bFjv08wmPp/PbfQQ17c
cMpL7ovjmx9KuETZolFUEkL7TqfxWe33V791KGSQXg/P+OHJu8pi4/RSqTYuDWUD
vr5ujLVYH7nSTdS2sQ8W/J6L6JVQ6wkan1J7EAOiSdKdd5w31pqoHVZBpnGFMIrh
+wxLvGO5oiORvWWfIgQvS5pdX8npG0DLHyUWvTDnUvPxUk9N6vXcDjpdAZqscHkV
YKyvqjinjOX4llxbbQ8e9FTShrVE6HKNZqL6a4ZBgOgXGMI60lOIIRXlmfa9pLLD
UrPrfQqmht0cBng1/Vj84tM6yLE/WtS4LggfJEb+FLPHBS9GTcCkF8vaLpaLve+6
OHRaagjsaUeEhByqx7Di3qYQ68qdYcYLJyrTw27Rr5rUHJP6nQR02h8gDx48Tdh0
GItTkCcWJ3eE8cDt+pT1Nmr9QPz3iq53z2ut2eDOauUJB4ZF+jIhZ0XtvriIL/xA
bzDQkSGmhlLYQ6xmu6M508dgsrEw4IbG8V3UnIxREaHH9upK2lXNH96h9anEnzvo
X0MCSNCehdaqv2vaE30lx8An/bzr9grJUhvXjwttL11jorClrI8799xCyFmaE+SQ
OYEFgcGxkJADxpz8T8Z85y0DG+AnKUMOkmhVmVgIl7ghUJ6obuSgTLOth5d/Heok
HAV2xs1fKuz18SEIxVImuThDWpj0va30V6M+W6CYvpPIbBS3QKVKkFRTQMZVqmbk
AU657GQi+5AYoJG1/+pCrI95cd5XGyVd0D9tmFyiSCjWmABjLZzxTat+87pOf7cv
2qN8J855rzPW74SsFzgfBKdaf6ipO+7XRMSyPQOVuzsYWs3xPuoDzNkzQ0PBMRlP
g8t2XAKXpAl8ot97ol87ZB5Nd22rjLzkPgjoII+PzWNcc/00CkFedN6CXbWtr68w
bqZohi5b+dGbpv+8BThBP/Q4EMzbTOgmOeA4DbskeRwoZ8DGBnJrB4HtZ38G3zTe
MsXKxsEsYgbZIJDpf4otnJj8O705j7ZmJnwqnwWsrqOgSXj1z8ceshgQqXJo6VNb
mngt+Ldrvmt8X3c1sSrsRsQbqy8vHJuxXwpvMWf0Yp0pFFoABShGnhkvOdb4oMoG
ofdYZHm+l9G/Aic0/9IxCZR51YONxWg1uGwq0R0dqhWYuSliqZ0MWRIixrDc+6uw
xK1M/+9gLegzNg97oWR5bv2GijIoH3pRkx5UNIP/RLLuRxFQiCsY4DXdAq4l2iem
+Y+Tngu/2YN+Az7NzQkwDt4rl4AXAZqNAtsyZXtDXEjL5Z3rx4GKQgmR0O8U1V5K
lKw+J127O51IOhY6LZ7sWhel0OWsGM7FagWk8LsvL/FxsuQf0w7fpOHblSV/YL1A
TnkSIPnEPYiIT26m/JP2Co+fV9dkGGAcWgsGQLS03cA91pCq13M5jx5baWnH/I5g
/69/XRkMyrzuiMXcyzdciHBGlSbMM35vwr8OUl8hOh3DOnbFZyLfvFiRIOn8MhQT
ZlQpA3WvkHi+ODLmzwjWkb6RAmwXyOZ3DCxkoN/HEyKOu/dZwby7KaTcPe/gegut
1Ir1HPnKsBrGmbbcWu+w2Y/ZyXOnB5JpWwzWAhlw6eRyU/zZPCCbhZO4u2Dcy0l4
FnokxThciT2j9Iz1BUqksWlQMWUNGVJSt6hC5rMvi2MuhEZGolxHVo2AUdMzvwx5
6+iAX14nnL01qUz8uCq3DuM7MApaCGRV3+pNasCXP6bmI64mQxR3GaaAbKv65gkL
/U+qe2r+LA7tPhDAGdaUtW33RHAKz7W8ihNw+vHyfACbqpXspLLjGyQmwzSyWBz4
T3YHpK3EwelF0r46WsMnCQPXN1WE+U5Y7bflzvO6Opjjw1URylpCt06qHyQINLHC
OzIFosW36gO5Ko3yGDzALCMgs6tDAZ4wev76aBVW+KC0tuR4A1Xtta2dVI/LzKVT
4T2IHLtCGAi43UA0yZb0XBZdhAwV9CaZA9BC4yzMvNOQY7uHgO+ctEGywTH1PO6l
aOzBCVzqdecomWD59+8FkRm1cM/jPmzbOhr+mpwfkl7lNRGuvOrKvw3OzPo7C5Ko
LfdZrESFJoJ4POPMNYMGvt3wDLXvllXk/6dSAoHB3hOJT3Krugt8AF70EPCkWPXt
XfOnNFojU36o0aNRCLjCwuVj4jiH31pEJyMV9NLbfAKX5/ogZK9HOzTXXTPSm0s1
00d8B8k66EMzI8MPfGavXM+1HUFRKlFK+7y7WMnIhpYYD0bFSKsTl8ybnCWwTtTj
h3R3D9vphfARgx2aZ02QY6c4lt4wAUp5WdDuMsKcQUQCxoD9cwjM/3LIjfCUK6ap
2qFeub45FXYPWHksGfGJkQaz2uYNbc0eu3fJkHKIoNSxyFW+/58PdpBaX/j2x+nh
Lm1MC0IkjAkkVYMQCM/q0nwJEMi8jkP55pABAbAtj6uxU9xkivE67WunG0zEfYPC
S5zSRnd6iA73vmXKL8fFDk9+Jol4GzUTGxxFWhfY04z7Cnpcnd9tqdddC++4Zw+E
0a25cjt/DF7C57M8zicIuXLtxc0E3KEy1jVR/m96SqjTVghuLevFzfpO2lB/zm4e
ZBKZyy+cCmSU1WbsjlXT8VqS8X3g4xiXTPl74oVI2YMBA7v1v5aWtnYScQ1WTlnx
BdtZkdLK0t3YhCi8Ks/lq2FpsRjo1XVymUHQ+d8zxRzUhbV6IgT7Cp2ZvmVDZQfv
hADq1s3UTZj56/T/+qreHiwVW7BOB4dtlwfBv770ooCTz6xC0zwUC964GMIQzexp
vx+mFgmQHcb+FEdtS56aZHE+LqDGlaOQZYoFp5VAwZmGDPyjDUycqZkVoEENVykQ
I1p1DbXUDdPRI1uscfokCX0eKcSVt6PBMej3/LIVJE89JYfhqqm6XxY/U5jG50Qx
A+mw2Fs24DS9/n4LowWYcDAKKyWbTcRE+n850vV8EmdZAgDhUOdGIEUNxPhQTQXI
+8NRhthvqW8wRCAxmrEruJGlhZ0v2IeRnaoiXUMDVdicZ/MOJ3HebR4vEknY9frk
T64LoKGCBF5KBfWZaRYix+1UuBOmSMLcAJjmDxjJDJpnEnqQ2C73PpwagwwSbQI4
q+7xwCGI6oTIpTFtapAOwMSRZP7WVfGWkE6JAvttQHCLCV/XZLTreIKHepq9avc6
wnE8e5/6V35BVh+XY9XC00JRUr/I9M0ZNwSGnEmwa0Bc+j7824OZmcLU6/yXkZts
bBZ5Q/n13i6TZQ3WnC5LztepAd3YF1ZVU3wXUwdLYtuJoqbZMjmyEwOKpMa6aEDI
htc69OATCcrQaQW2PNeD9aDGv1v9LVKXFvNk/CKXWEtLLHKSXTm7Wu0rhm/ZNXL1
hT9K5HdqQ4QgCGfFl0VU4kkpAyo+KgouYjOvkD3H4cLCknfRGrgrLsfzjovC5xYK
yuW0pzBpk7iDXcFaVpzfUOxHP2/lyiKTZr2d+UssCo5HndRIpzH5/UpVeP7ne1se
BFoTyWb4iAMJmMfR98dJLKzZN4Y9AslOEPcHNWE9TPlEdMlFScwOMpy+Sb7W5yri
49Dbq9dAnpBtKZAVsZTd6OvxNIch2Zu6P19aKYFaKQB43wbb1DaEg48Wpp9Arvwu
XeF1YChx3+ntopwBUh4oEb05F4XyJ3jrDp4uO898GtLAg45dd4NsIIy9pa4s33+j
epQxn4tPUxasYDMLZcW+GSLawj8Fz4gcST4MS4j3v3kGOH/IxNxqWsTJrLFJp5Ci
eTskSBsVyPLGmuOq/d8hYBeyh9H4a47dmsShR37Ey2mHSIOI4io80g2opB68g3S+
33Zl2lpgdFTnQjJcDab8HNSt9unz1Fqv9Iw383fzWWZdV3Pdfc9pZj0ANHSW6QBL
fU1AB5pl1AhxGYpNgL9DPcO7rZ9UHHz1bfpEs5QBT9fKb16jkfnUzGjkS+YguTAH
3pkQsQlcwCAMrq5y5KhVt3Y4VDMZZz7hP6Bsv1DZuCnaIxpcl07Z9Yw/E2APrXsA
8bRS5a1pOl9yuDiH+Mi7yB+61VGJrNlJ/3TGDvioIgrSQNKb1Gm3mbiXk60Rgt6b
In7kF3S85npY6NZcrNmAY4Ky/K/a9jWiP0qZSrKJl7cFvNfuUaWP/YnnWCyqlhPk
5LPxkU50LZUt0IXtZAmpWgMV6EANG5fbubUsHvImcu4MJsDOccKQmf6KjK5CdNp0
pbH15AWxo68MX+N3lqM8i67w8/NRfAjuJw1kdeRaEN79Uq3iO7F5fyEn7RhDdWbg
Ver8OsWqAjkECNP4ph7+oPHlRFvR0iAiyHgkBTs7Nbo/HBD0skruEGOAGuUKuR51
XxGNWENOpN5CwRljyZNyWMG6mEWZWL3+IzUKuGAZF72ZgQyDfERf40lIRX3fPLxh
FMP7rZqv8kqbIyQ3iKDBdyqmu+E2ta+2M7z2q19D/qmNuuWAxGlkrXb5l/W26XFb
38jdH3FSSoXe20sEGzTWiGLng3WAx9M1GzEjXbhChdH9B2RcM6mzwcxKTGBMTgN4
bAikXTp/dfg69GVALfUpwBW2TDyu4qynFWEdt7iLq4LCKgyXwwt8TQC7xCvE7plg
BHfA3H2o4AGE/GTb/InF+7QScUoevBYBy5wIZcOPfRLAt14l7YJrj4d/xKZV2N+/
0KJEMBa8n3esozGOMyBgg9oNBg0IkbgztmGReXeAhFjx3U+1Dsa2xu0Ds6KkyGk/
EgpOafsH18zehpmXsaktH8QXMGov+5yQfnL1HRy6ZCh1Y/xLKF2kdVF0A8gz8G2+
D1JAnn+rWPq2+LZhO/Q1+gQieanZdGGRjjsZTtGW+x/jWv2fwa4lZAX3BS/rWzO8
u0MmfM0vKQ27mdNCukVXq/mG4YdNmJs0qWFrmh+jzbbeNxSMaZQ61klsSQZA3TTe
VL7drcDG8+JRr51CpHO6cLn+UXP/A5TWU2L4NThCxiajECw5ke5lGgTYmwM6sWx3
WWMFTkOMO9YveSWMZdiLbVXYfvIv3SWojqFN3lIP3ZWh/R8Naau/ZxAEX3cwFSgY
0sz4HlIpJ+y9tW/LQ1L0MgbJFmvUV6p6YvqRoixxTI1PKK4CJdvUvKQ7Y8sV93FI
W+0/Rg1zzLu6IFSp/TAzw6TXhaifJBChOh08+8YSOw3/BVje7N5bTFz8WK5p5l09
x7kMmoyp3SLnqX82Svw6ofhATidNweQmewaSxXQBHJGc+FnDYjUCVCSsvSg6zHoP
2EyQkjoga4qyW2wdzFVR+R1sxQ1IKj4vmDgXe1pkWOODb9bvCEcTuIVCaJbSsWIk
DPMVm72zmZ3D9WAdYOWMCrlugesR+HwX+Px/TZ8c7zGp2wQ7zwJmPjFcYSvN2ZC1
GmoLgLs935U3w3HGZIRr4Qr/fPuVk8iAr/axZlGU1Mvr1QRcVGKrTBgy7yn3NEBI
ITweymOJ9GXMwKehs3voXXQSvyxcEypOga8t3Tn09Jpm1FWvqqXnxHZ0o0d+n/1I
DcoLZ7VzYjikxIJSuHetFUx27pkJUbwwl053SQfUymHzT4A6676qbwrMolriORSe
7NwH7xUjpbUQLrplhhoyHKDnVE9uwmCno2n2nMEtnerSB7LmkVdBfARqu5KIXykJ
4rz9jNjFPLQAoG55XK+2AhHdVZ5W4COqBmKIDfjL6919nzJgIWKHwk/JdG5yfxJE
bTCAlsK+aDtHZsHgn8hpZAk1P007scy88/VTVgseNl6fn/23ADKTo8oPSh6sAk7I
bs+0FVtURxPcLsY8e5ylDo1V8rETcHJue1Fyj0epHj8mmO+OqH64Ui4QQu7D1D54
48cna2AXvVPe17aYOWVG72ikcXTg9M21E4rYvMyGycoJG5F1j+aqFE5Cdz5+Emim
jIj4Ysu9EUTl7OLUGiPOZbp+hMxueud9MhgShaGr9kI326u/FY3dBmOGTLM4CRuj
VV6h64Dcy/duj8QTyWXU9XL6qZSsFGJdzZ7aaNvz5B+ZUd8xjJ6G4Fx4RGczs6Ct
25gYbAq4GLh9c2iJjcqCRGnSsk/x01DBU2K4sCP+h3BrF5Sid7NfzsE7Kjza/qkX
8fUVsomvaux74nXheujOIQT0hnGlXRX3rJoYlfaIMLslHc6SwgPlFE11sJyqCigI
Xzjr+REGJpE8VPRwps/d48Q0NHy6jWm4Fmu3LuLncdeDqphgjytm1fNKXrDRHVmZ
OqLkjrXJDLnTXY6+EPx66tMwkSdPS8Wiit2vOuIqcH+mIymGbUEJ3/gq0RirAW8z
hmQoIMsT7rMUnM4wl6XX7NRYqIiHl6HGZNAQEYiFmxnF32pYP36kUqyq9QZkxlGA
olgVJ5wSCpqmkg6BTmUabsubAG/GwfYQ1yCQfMOujHhKYsq7DOCGmZg3tyOT3jQD
z6nzxQVOtb754sGLy2ub6htUVenscrfhVVwSvkYKDAuistUju9HWZ6j9XSnrGBeP
cT8Mj5rm0xELSLy9f9Rv7wHV4jpCD+bkQqerGEBaH+noy48vA1CZYVjzghVHUG2l
Qmi1T+zX8ygirtVmk4MhiIZTrvlt2Yw6f0BUJthHBDS8Tgm+wiE0pqQ684Qeo+nw
hm7sSOtU5hKGOqUl/7E+G/AJbPPYajpRxZ3jFu2lb2RKd56g+HYXyzMbLD+IHz+s
qasXCA92X5xsDKpJY8VphoMSWG05ReIOWB9zWlgdnJ51tqitxB0TLN+X+7ZZ3GN3
TpkNMYjgqEHdftrm6yJ7O8tVsLnyuho6u/HSS5TZTcnDO3zphME9lTsmzH6Yg2Rl
kJ6gcsz0LzQ0Cwc/sdwqi5TnIBgF7JGe8q7OuLZ5AtsefWspMcpoA8x9skmFnMNQ
SK8s37HTb3j/JvsCII7NqR1SmOYZJos3ineh/a/RQ1x6sL2rFmCbPyDdiHw1KBJy
rklMI9DVTSoCdW2CX8CoCPSwsiO8j1u6Zs+/BLFWmUigxXAygDxYkJS/lkGQOHUA
DjfWi8tM/MMX0+iBXF4bwf3aNPXSid2nVBIWeQ+90IhT8QlhfhCzM4KRdPD6hv8Z
SA0kSgv7ibRghse7h/dOqlMQi2tFVRsnUDqIorsU5fSIzy8uuvUn9fCoDx6vF6zv
ImcbWNF3bgOEFqIfV8vS3xxPGpYtPOgiPHTPHPXTvkZJKgjthYnDuv1pV2sgM+fG
Kd7QBl9HqsPW5i3PFQtNX6Qh/MA6jR3MRmXH04tt05nZsQBEq6BRlTdLn4N/X3X7
/QOlp8DrB2iwfSM2L9px0n7f/ew7zHb6kpA9LFvGDfQmEZNmMmKZCmrNHd+Eh1aa
XPoimYXsXltlPG5TduiDgUWicA05R1h7c5YkCaBcnR3sOC1BGdgXJ4SvQUUG+BVZ
rzxzI4FVwCd8JF0tAWrnrBPGVCZIXbLj7VScD06Rs6ShvAQPtZKXJxcwv6BvnbOB
f5ZA49tP7QNnevWY8zq3Md5RJ9ctNtPmB0bjvYeW6YtMhYND7nblS71ZrGCQFNyp
Kx0f2oWs7QXut478aB43PfDTmHWCdfKObjCBuaFm/LIR6odMOzUGA735CzUH5Yf3
B0Nq8Gi54tc29EjdnJ7uJhoKCezWkNuANjzsNVjeirg4VWmk/NHX029z1SGsEzmu
AG9KhEw7GzrjlaZ/WxTKOpDVRG0TJNpC615hmuyZ3FfyAN0eT7SaepziLVWzRgSg
xxVfS+m0/Wy403lkw4MOhjF6Ac+1HOz7LEpi+itHRjHt6ujy5lW8vJtr/QHabBGm
dOcGGZgPSzRiWZuWp6kCM8yaIO0cwuTPaM44Rj5SeihPU73iL+enpw0WOXN2yAqX
PhlKVjhkRVldnLrn7PVnlDVn1bMzwA5P7HwolPt+WHDoWe6mAdFXhq5TeUuSxkw1
NJ9PB2TmnD2A395E6znLFswcCBdM1eiP4Kl53zxhys/6fbcK4FZeO8Lk6mTkKvRX
zHaPb3EnuT2NT3p7dqxZzCe4tjrNJK6jsXkIgsKl0ZwKhMAfm0hN929OHNDpXTMK
5CxiaTd1U0/K7oGZeOkOYQNyDHaYOQl09hCfvtb4BPbaPOvGt49kga2kv6gAbzmo
JEPeWo2gHzCZ6ipzRecUAQfFWaAy6zzrBt4/z/DtbX2IXyo5+hzjTuZLzFmPJ7s1
0+KxgOKWZwO705fMs1etxPwEHrg0MlPnfgdEDhOksys6ioTAPunXSfFTMXEnF/1p
2PGXcPDgjtqwX2tBoegnTvKuSfGyMIOwlyKoqmOUF2MStChT5OdDh+2ITET/82oo
zrorHJDPfu7JGXeBm8XfFziLg0vdC/PTar4I/LgDI7h/Ho7xVAMsBOpD24aZL3au
UeeFtgro9H85a2v7DyXP+SImUhxLfHKZIsO2g5HpvJkHxAk+dYAto9N62HQbKGHJ
A090lDN+p7tNToRfXqAW8IzHmDSFhDbzp81kdfEJaN6sKIJENE4PJ7CCF7KSqyMZ
HLlUIlGcFxz/hQGmZ6+5crUsjDMiKE4zeUwP3GbJXEZCsrzj7kmGAlmAMEP5/+Uf
QNgo4XdE8nnURH6bh0wv61tj+YCjNqmhIIOfYb7hQwGR4MV5HqCK4ts/KLQh5Fx2
f3MuWDp7W17knrMJGO0YV+H0F/OKCmuzTk6x40iRALyxSgYTsx4LXfYmPV2F/0qE
8EAoTut2cNLyBl2nTHcVvQbOilFA3Fss9EE2/mUw4tOW+Xh92L0IpAdPGItZhi7X
+cLMgAmIamNmv1rXd4L5FOBZ+UO9K5QMeBoRxW7QHh21r8Yw1X6JidLZPluZTWz1
QDh4KUUomI6UMK8FiJuCRTQ74FUGwSBC9MJKw7VlUVmNPIlUHU5zyWBmevQ0UVia
ecFQuEY4xVBqvBg6SIErc5FBF6hHc3AhwFOJ9NPnl82iPyEGEwwWecx2pGc/oQDh
MAnlqjMkpQWAsYx2rOdCDq/wrZhqME2xxA3i8Gp+S0uphAYnoRCZ5T/zNpRKH4ao
okb4iFDASaiS21P/lOXNZBoyyjM+FBYy0bkvZHu0WGZV8TquhFU2+lK6B57uRJqr
7o6iDwj5BcXCRpesg4C+KckJuo+mLpP0tZCmUFjr9Lxivnz4JS4O4lyepuEtRXg6
mr0yxsuHe71jhlFJ1Z6zuMyjfA3ALAyvS5xPcOe2McIh2msghKi2a9ovCcJRWBrh
GbS7l/KIFEMq5G9n4JIFYtAlkN6SrUjRqEmeR1kseFiogpQZ0gj56vUC6upv7GbQ
zKD7POgwKzP6uYRLtZYAPol84cKcngZDSuPg9ZVH3FoPZWJTQ1JDTMG5VITH6zdG
TFDb7Xe7eyTqekfVCDFaKjjVCoW90Yx9XL/zkG4fuaFvwPugjW8JavzZle0WCow2
Gpsgi2bRnY0KzUq2EM8FvqVzTGo+m/uuxfEbeq38zBKA+T786TtGurf46XTkW7jV
jlgkjoxKj9Eh7PJw83QXgi4NylW21Zwxcac6Z7seoDl/G3unzb9Lvl4teLooZWGp
4fIZ2zpADe+XWFtXTYLYu8KHqr9hst9D+g5n7lTO3du192h5HQMKTpU9uXR08rKr
CfDpKpOrXJRW+WZGdzz+Oij+xsIvJfOq0iohcHJUTJdADXiroWshWqorBBs2fGa1
eLyh0+kvHpiqgZ69lYSOnTabByrwh30LF60aYrD6NNPsfBJ7Ig91wMRe/CdDtXv2
pUKdSu7fDwEy9qOwdegb6OZ0WsaPBdWKf2eK244Ydz3w88MVgOvfNmaUTlEb6ySG
ZEoZahNO0cV54IpfnZrBdzGmbGAN8rYkZgWSl/gj1RObfaKeW4JaY3KmHsOJCVVA
adlMzutsX65S2sXOPIQQLJYLmnXV7FzjyEBi+gzzA9PuDolkeDPB1jvpuSR6M8CQ
7Uqif5xwanOx/8pPHXjvZlkvVdvIALZen9ASh9pT7DV17A2idgRlPC7wgQ5sNYBs
AE1ezLOr4qO9mM+tlisk94uX0MEEjbMjxEmTiEfSYKcvcsUwl6z8JR08tpH891G8
NZUcE77v8pUIfJxgCGLQPKTDF9RJEIjOUvNIBvhaV9efymXsK/+6Ax0dFub5B2At
5gISepZd+Qyw63sVirVd6Lz+FLBKSM68AQEsRDThLMveVVjHNmEeqJBMs8I0C0qn
fNr9NeJRQg5i88TC4CFN8451ZpW7I4zRLw9FKlOOYbIJzd7njjmj4dMhfWQEQl1d
duUtYxj/FW8L+lrfr8lFxWBoYd9C19sL92St4GpwH03J8FEHWQhyW7PPo77AMaXz
nHrILPzpHun5EamaPVqYLnRIZlh6NTzcDr2L4V7hpzuGePYQRmKjZBriYMf43T+0
2SE0U86R1L+MDyf5w4HYHGD8bt7v6YEcsaD6KxcljegCuOTgkepMZKlF80dKTH8b
PoMLObJO+U73L1nNfpcwMZs7rU2AcgWH1givoSYPT3YtWeUaL4VO6Yw0FcPS2diJ
eyfQgFXhZ9aMNk16sAvIPBhKP/qlf/XXfrOF4dGFoUa8V1J5tcuh1+FyemTYr36k
j6FO0E8fw1s+XyVqsq3/seFKIEGauvO+rE2Sx+ngmVsXkTXOd/4JO9WSOhFBocsM
AJZoJoRoIUf4M/CLybVu2IrzmhBeKquQwhYEdxWPSoilZ0sSGjKllNGkSjrnB4r/
QerEpBqWIrBclVgVhNqK2J1LaQQ2WTf7KmDMpiYbNRQCsr3P59tuivAH+MWqydwO
mCeH2rBlEOT+Svp0tpt2wuTDm+LzoNUzv0uGbIhO7KoAW2B16UNw+ZgBg78MKUzh
E2DAzhN9TqqfhbrXeTwbQ3YBidFKr+LpkgD7JLYLvouyChf0B/ZhgcceMOtqkLF5
eeMQ0GhHSsaCZAUlXD40pR7Ylends2nBCb+3XDFIDliR9ybPNLALYr2nlc392u7Y
9CV45ewkgzU8bc8gcs6pYkiWra2VFwWfo1lcYIqEWzy3pvOeY91Fxo/3m/W+D3V7
/Qil3Ng4YxFRwEdD8iowLEd2X+dV84EHh1SL776cEsns1Ta6GSoCJi5hMDSv5F3S
grFgZ7s6IXvM4SRXA5OFz3Bk0TUvJnRQU6+JLYoV3HSyKhZAFqBM2YvGaPClc8kZ
8O+pQ03Jx2UYuuwRPKcXj3JwpF+lF1o94nuEIqbTVsshTQqg5g15vJc1UwqI0keL
8QuG52ZnkJNTmNgwpxxA7cThx1+yrhrmvXtMOBuzgLeIygeedLNcAAJbf25t1VPE
ypHwDN/ozsKAJBJg4iHcKhVnqqG0yaEEfLB5k2L6g83XurbP4js2/qToNeriLQOY
E0h1K1dbdGY4JeXH5Zz5SHOmBfgElyCm/gEzytWhj5JMrpvSP8IOUYrDPSsvMVn3
i7t3zhRBQDKqoCkDnQM29XrA1VtNofupIjb5USYHHNlmSZmh3FFTT1WPcdElzSa4
1HmRWtY1/d7/UsGu9TztB+iecGZZqL751GAaEtPUz/MFdbe6xlRb6G66jCnBjhe5
JcMeedwZ8EscX/igDslaSM6Xp6hiPBnXY1eqpbOBFuP6oWY6xc8R6U2ZH1qUHTZV
72PBpxslFwJ67QHui0q2ZnAYoG/DPApSTJjVKpPOolLDyQediEliqN4CkCFmFHy3
HFoS71jsWTfRUFTr0OgBAqoU0KQAIhilCh2th3GvG856r6qEN3ylnkwF5tX9iAsS
cAg0Qunc4YuwXnkRVgGEu/gnMA1g7rA07OWrTo1rZmLZW0gvD6Ea532qkXXS4xmx
kTS87+e8Sp9Mx4YjxoHLSL0t+4MRc5e//Y0OM+A0E1CUeq3MhjRC6ZgipOxtLtwU
mrrou/PxAIbKw0aK3D5x7oE9vWXBT905jLEwfrgmQtdAcAxzGyekjXi3DlinSKcR
4MQB1jTkVGXLqPVp9XjB5OE1dEQHLHhUFW5ep+OJ3XeEcH0756/uWdfKpm8whB2p
WbazBkaY4zrWPuKzb0eN4Kt8XU3qRCOTUHC+Po7NULEpGAypuM9xxlV0HJ3bjW0V
2qvcMPgMzFl0IwYQ3BbvuraCi6IKysm+dZQ2uGcDAGkpstdJ5ahI+/QmRSSCQcJH
TdsaRiEoTcN9ehF07rdV/oy4oZAWUKAhOA8D95WjKG6gCqg/udZMTIJmy0bAjQwT
J4hspSy3bJ7JEZ2TKWw9G3A8U5bIpDC5Awom4H9iDE75Y3dfkz6j7mee2Uu78BGS
wkVuJStTLoBvhe9Zyk5t0M2wkDTb/9+cVhyd3Wn6WHyWmXCyRCU4IPrp1CB/abDJ
dFfGJVLjwOvv8NX4Rr6Frf81ZwmBWMFOnSFjepvxJ27V25yZJaz51h7SBBe/87Wr
TIX/wXg/gzdipNiLgVMIxWKc6dMfzrZJFi2Q8yvPpR1BP3IElN6UB1g1zU0JeYp4
tzg2l4eH7spuqjesNpxhpgO7ODrmlI3cses9D6ryMSDGzi6fa6yt0rqf5mzvt0x9
4nVLW6NRm4Vv+dVWezDDFO9k6nzdLmSOTbnCiF4MVdtMr3ccRTNR7cTt2oHu/ysu
YXwd372V+7PXbfRRPhnPe88b5nMgBg3HsQzRYaomvlcNORj5WiqGNc18m9/DminX
sYS+addDo1QOqTniaICVjywP73DW+9T7SeijyQ/RcBJ2x3crx7ux0K4S+Ms7ekeP
BPiqfxn9ZcJzQItYgBRthOhTKemPZeGec1cShwK+eKuT2SLi7PzPG6FCValZnDjm
71J4177wM3hw5oncX4TC1pwrJx0yXkQXqzP2XB3lc0GOhCBrsa/nYDN1BoZcesAj
zXzBm56yydDSit3dpyPGv414mTYx9FjKf8XkG+Nhz0JT8BLOAzS5uCoWtdii8up6
V5H31DVUrlmVrZqX+1TFrc34x4Z2y7vxTRh+osisby3Ifvu47ra7Qyq3h5GL7Ikq
Ac3Se9bFZsPu6FuALVFVzD/TQKo55PlgP9eIc+rNUBSylgJEsmvFdTrnIfLAKzDh
M+JaKIEzLDdA9PolEkeA4Dn81h4NhRbc94F0EpPTKOK2bx1wGjBIC56IaUp9J4d5
cx1ut+jkhQ1LxotVDX8oKn2oQbP3NT+FNqyWZ5A9p79zs7hznaaQ7qfOK3E4pcMP
ENjFgJGA1st38Z3MNlTkDcZLH8fNdlIKwT5dKZIrdbC+hQo6GlDTgayR4f3DOCeE
CQJIaoH4OqIRhQNSq+T65dUKFaeisixqkJtO+HJpL6ZdUD4D0D3WEkLmUtbuS4BS
CT+JWQ3Akx4q7NUWlJ8aTnO8R54BSWpvNBMM7CspmSMtLLU/fo2wF1Xvr/lObg8/
rlabtzHZTpovr/NEQt3mZlWHaAttwzO1Xrbi/XWMlv7mZDPdENlp0INlKLWbenxe
GHSmnzX8Qu3dj+vv6ofp/0TryZ7pynfPQ15ue2m9FyulqLeJG5kP39c8VsdO5z/S
2OEvAT22HFJRpJ6+DLAN+vo+xmWBZSjJsEXfzHRdjktCVPtblHSZKuf6SnKuJ7Xo
+oCseR0k/fgsbZ2gU0wfdY+1AF6DhA5mRtGq+YSbmhhDpurPDRNROkROCkK69flc
ZBuoO1rf9Berp5zo2FvYFGgHRW+AP8GVdmrJDxmvM2e986C5iGMycWLXVo2zZ1r0
RwdCeeQUOiKmr+Lgyxy3elzGut6LGC3qvcnG6CxBCY1xNKgfjAi0KNyAoQRKEJat
QqjYrLku7ncx+I5FO0ET1tx3z+8hZmgakFZs0COrfET0LofCgbICSbiGikeilW13
NDzVb0shtVn19y1uVxsHsRxEEr9ZuqE7xFK7AFxOV4axiTI48CFQfCC6vWH/o8m1
YbyuflZikxvEZuk6Xg3ZaZo6egvpCYzW0vd+LA+BStP+xfTvJTJuAVwYQaP5PJHl
BaV/AuhUNpUajsZwif/TPIT+h+8twSdlwAoTO7tEZuIDCH/DuIlxtVVJY7flFNTV
Ryefp8hfC11uI7CxOQSDOvlV9NkJdHzucOLZdn8mOQ2o6MYhQeFcFDsO15e9M46v
hwzHhoSMILl2Y9IoJV4L5NYxYOpLdb+2bIUlMmSjsMaV6FjuCQq24gjtIT0vUQlC
lzi4mzH9xquLIHWfMsndzGdOjHRofXwMzs9oJQSxSdC+dEZzJopT/8E3KtHtNQ1d
boqFC7NWGsflxaCXWm0jnZoQoziz41ZR9+vXpCHV1OEPGdOQ6N9GsKLAJoBxMLNO
UYm8YO5W57oaYxYyTei6QeJcmw1J6by13XAaph49Bj9GvhLp2EkzkaxLrZoouxzZ
qhA7GYNCfl1yZ4CuBrh0G4lKOjThU9+iTCYDdUoDuj7LeJONtT6BdNgmLDh71Guo
DR/wG8S1agKc6/wu7WuVtD6c2Ga4JwDH7aFJbOLUW70RH8iAuJK6ibh6XZqrhKK+
ridnTTS5rkjApjGOPGABooQLmCN2dxupCMnTjK8fThuRgL7+ycMJau0rPimLHZHq
pWcO0GrF62PRfLOag6mrWm7O6I0UFOIofC7iPUzTl4x6bGtLlkkq1ddpKwHhIbIU
FV9tVqIOM5F0BemAKShVWy3VshTzXIJF/P2bQZf9CA3inDHEfUG0CtU3lzUpEcae
mgbKOFdye5xqZChDAQdRM4qkDBibI+UQOg3I7EerRRPqmqEWDCSqvHLsBdoTKajF
uIRq1dIoIcGoN7quXjz41SO2X490bMaS+a/+8yWUBy5I8k4hjvEcXU/FX8yDaE1C
My9cgeng3mTWn70ICbywR6P865hTwa9HEK0I+hlJAIXSIGgf9SuhyUAOMv347M1T
e7EUZZ0DhvQODU8+Dk7u406j5QgMER9QC07EfYRGqcB2sR4qzt+raqZsRepvjLmd
WRvopYVkxN0D1dm2xpPbf9vuZQRR1nyP3HZo8/PmMtS4FTfe4Nr0991bdaikWJ9d
ttQMOebh3VRqqJyMXy9hRIIKPgV52QudB1Z85KAlWxnmv2oBcH+5R0Kr94Z2QWCd
4w7pkpQ2RQO4BOGv+/eUk8BJtRnOQniJnIXtinmUODCmmP05ZoWKsgUitEILUrpI
GIXS7HnkriVknb5BcZQUc7JwY7sFcjdu+iJQ2bBEy8TnP1A79UTUydTpQhZmXrAc
XcQV72B3flUXU3GBIRglEgAdD82BsshJKOvmIdzYY5RJvzIkYIt+JR2qjxAnpq6A
RFDJ50HC0NUxzzZtSLW8jW2stqK1ZpnFbEKb+SI8fW4OQKG3onSyxgqWcj4wnhCR
9oq9kipdvCuS06qmNRzgGe8C/o3lnRZoqnnjcD2bCm2fWFjvQAUXV/SwgDtk604Y
eXHTTFEczyVJrxOKrmMRVbCtAQ4J9F/0AgVH77Qx3xeLVFOYJQjk0bx99p9diM7O
WZ6atM+Jk1y5qqufRRDj+SXbpFKncpMLqGfydEnse647hcp9ObhkxG5ELaN+4tG7
jOy3fu93034PLw0FfyZ9v1h0aT0ZGx+2+3GJ4/Nb6JpPwO8LnkrLeK1cw9QTzeGx
kTGl2VjzNU5RLJNoIljLjIc0mDrWN7g2jDrRYh1EkWYOmzI4Zoq+cbU7Zr+gVg4f
UNqqoGN5UATxhl3rqKik0NC6Sn+s9ksVX96Zm7PUzWiQkcylnVK08gWMyWITOWlH
GJbzFwiY7p7XUWxj9EcDwJiCSTD8+UDJ6d9DNqLMPgF4m9+tk9aBXgQsZcRbfJ9C
h3HGM7ySStz/hDSMcArvKl7m87qtspOwkVNwKSmNGJ7U8ZCRT9vaqTmbfktXIIZH
66dGcczYQAyMWThzt30smRKGF+FRF5l+IQi3rPeGMzqxsBv7vKikRHi5psiDOCUu
xVRQoIPZcLg2Vu/B9P1hyU5/2iKyxrrE0aANxk7+F/t4xiIpr2cplt9Qv6EBVBfp
ggKcNWPpubzK2EzC38oqNPdORFiTjpgpAEsj53pm80CKHXMgzXcZsFP4k/g0iZCM
TbHRPSbFe/yu3I+rc6RCDG4zRsuPJGaOdIeL4w1PSjsYNBIisC0jLW81EhETs1qC
q2sRX2ehCIej/cbyG2PLxhSGMK0dKlg1WSNu8DIyitLWnDbZ6J05V1xXmjnZuj2h
lIymCv0XelqJfBs8za0EgPtW/PBqGykoDLQCG+v4ODDW3f2hlJcLiOv1Cv5J7d6w
loaYGQDHUHEzGHIwv4lvfncNUnUOnjD6CzEN6KZZdLQ/BSFfZbd2A/R7Ods0STaK
/AVHOnZvizjsJtnerVaHYkCubgHLP/GxXYInp1FBSafhUo74XMyE+jMoRoELheRS
yHtgl+Xj8XGYkAcpGw9EVBUyuDWdRV4tJo+ZDHNCjb1cOER38oM0QFVicNC54bRT
3qny5EIWUGDsUwsbDPSnr5dWsWa9xWR9Jhxwb5FLskHGOGgnRKPsSrpxHC/KPN0d
O/YBVPGR2qpLrNcQolPchy0ijM5XHdGdZC5XDAd59ibgTFrAoWf+BQSmo+6GOVvX
GktdIPN9wSEyWeOl08wegqkIRna1zG3HTWDiC6B+t38AGMQTYEv6nuZ8jaFv95e2
mxmWHeTm2vLjwbb5Bc1CGrEQ5+Xtpq/MTY8n3XYKhPn0ouDh7B6t6z3S7f+Q6SSC
hb5SHBOMl4pXDBUHOHfK9nvR4ZNx0ke1rwVGLlt0XDgq6fxHQU11gaP2fElq0NQJ
FdC+8FORJvnPDSSqOGVtLTrchK7xi5pdbpUHPhwopeFBXJ13B8BSPCbz1kzdYlLd
c/tPU3QMlY2bEjuRtdEHB34yzV6/KFG5hWnnT8evLgUgcVTVWiDU3qk5wx9v+WPc
pyW5hrRXPzfQByDjb6/23zpX5LGfWL+tFLWFoGJB9yXRjlQqHzudH9mnahHf2tC0
4fS5NSJkf/A0r5Wl86AEQKLtGKxFIQ4+LvRJc3iB0x7r8qLEuMMyf/s1u3UA9Yeb
N0ZYxJ7YWyRrdOYsgkoBI6IAlg6pVXKqH4ZqOInERvtnLz7SlfisiKTSx+st14vQ
EEp1ER157EbybK7b/YnvsxRbBU7YsZZ9orddoZ7Zv3SvTQrwDzxLmFI4WPzYL401
3F8b37IUkA8uauIeVlfz8PDFEhE85xQrbgeoxm5tqF+74W97TNTBtB5d3sYRxxl4
kesiNDURFeZzk5VNcDkg9EgbvOKfFGJJc3wlqe7hxgIswBytGtWi+eIk3mu/rfRx
nnr/S0LeYuZ3XwqAw5TT4epAREwB10XbKbuPUwctJQL78qkKRw0vTMPX3dCfahoW
shiwz/Qm7NqzCnZz9x+aLOBKvOs51GV4oA373mVIprgDcnxkiImrNdNU4O919L5+
xd+mKEXPTAJa9ojAoseAZNDpQ1OFzYbPWFTvlGvdyBiQhJoyz97To8hHtWHA+J4b
C0A2bUiree0X0QDa9hkqaxoGwaaWa/+X/uMMN+e5SSfkXIdRpYqsAp2fR5+Kl+CC
af2urcR+1rJdt8TURvdL91GnRADHGdnNObBiYmEcKQpmLGqULZEhRyx8tru9U1r5
TyPHMpj5e9epDxDN/eaxiOhOL0qXcWeqh1YalHvWl9ecOCFDdm+JMZDLFasxh986
mlbvabRHCR8y8Aewyn9gKcqct+kRi5dVWanMjkxVzxw4VpnqTvZ3GkVxX263Xpxl
sbAGTFKNXjjci0y12EE2rBIXzZtMCynMR2VJ2ws5vt/cZ5Npd+SbwWLXR+E9IR2R
aKFgttVGoHoGg/csQdPKns00iDsYyQH6j/5GjS3mkcPtM0Q2DnIsAb5S6jT7K0Ls
X54HwvxQSqF+0S/rkg++CU8Fz0iAvTMJbMxly83dcnCoJFl14fgmKwZtf/YAqqvx
M7FHYiPIXgWmE3Xta9BDihVNtltFQWu6YuZDi8kvqWQpwK/Rs4vZ2CbTDlBvb4RO
Rfp3oHzQvKTh7qB/7dYMMvX2HACu+gkkvz37aruZrqL6r0UG6ADIvltft59KqxU4
o+Bl8PcoDM4sLtglQRB5ISiSRlsqgLKsm4nDZZsu/jIdYrpq8NdJWI8NnUG8e9uM
VyQ87td/bVrMZiiDeQoe8mxL1NmVnsWxOhWrav14FaP0SPAknfyjYV/jXqFSxQzt
VuuakkdPNeiUepZWEK0UF9hLZaCaQm1MmBtXPRtLUMj8jYpy87pyJbeB8hp7AT86
JW8bJgvuRqipCX91xm6bM5SxHCH0gO3pDpmbc4I9sz9S0NuiIQyicUnI5yPdyUy8
HiQL1ODF1iPwVFq54oPkVNWb/i6rxlkrljGn7tQz/wT8cqnLjRHGe2kR+DS2Q2rU
hgyZFrCDKS7z52NpL5rFRsObeLSiYeHiBvkL4TTVx32WER5CYsPCxDZUyCLlhCMy
DjT9oUenLixTvzfx2/0w6ysAyxYTEsd4+/7ygy/zj3yzj6NFFOlk31rBsedClKvY
8vhQ8Vr3QkHKhB6NWEUnC0tBrExNjdmFK/I0FbYV/4h3o8oxPTvNSap0bgyfXcAZ
l0rdCOHXOEkCr9cysJowkEUbu2gDot1yo+vx2Dx7HJLXRPtbpJKtL6hgLuu7MWaf
QtiD1WJberwUeEfthHCJgEFATUR4tzqwPLiRigFZ/8w4RWM4dPy76DjTfdhh/aPN
v6HrYD/pXNnWfftti5tct3UE3JbfFK6DvQsvF8VL8Xsa6s1sfahMRu//pYTrPfyl
w1pXR8aKvxG5iFZSExAmAm5IQuS/GZ8FX57TfL+hBbLxMglzqHWeCeZxVOlwuCZf
0uwI1C4O9RyU5HA0IbemORvMaQRXkS/Qh7TUKebN8nKe4MobGTasCvwiGBDedyX2
AsuZyddxf22P4+crDNtavl0lwSMpEueerdxs8ES/5K64h8p518u0AbTEj+UgYnKI
CMdiisZVwxuNFEzai+1pjIhZXZLkLuWkN/UKdiQczG2I7egksZ7Hqkr3+NuaxvSQ
7tlqi7P/YzfPqmVqIVcx6yuOJV2404gvqgbfhbpnksH7gPmgynkaq7k69aNxf1Nk
9QNtOtHya4G32m8ghdp4mPFhLgzAfeRNrlD4+aEOZP7Q3igwBNq/1IupttwwrPyK
dmxSPOe4VERqNsyLQj0+gmcKK8O4EXuWiqUa2HkoD9qtRwVYxFR/MSpFz32USjjj
YqVtN/4Lc+dVAk41SuP9HjCdLfoIy8MpV8boLWKWUxHqrx2d4tbz4ZPiNRNjBZwk
/RVeQjvA76VfCO8FrmeZgenYdTXsXFJIRvi7G/03JvwS9z4wEBNxEC99HbMBgWOH
SnGLCJK+BBB0LRJOAsZgaJ/+fsVTxdXBFhDgj4i9SuyD+GOVESPsYa7ZDpGaTRLN
Om8eAi2FXbEluYOXCZdi17tdVNfZfG4mZ2zgPpMxbmWtNArMi+WlSOCOiWrfa/8J
anZ6fwL4vShSGlHPHqyi8xVG8nyl4Ty8/pW9dkHFBbTeAWRG4QdPFG2uhV7g6E9X
h546fIX31OAuhRUh1tG4hzQjbQb1hcfCDmm2pRjHtlzCZcvOm+zhaCw+5BKWOs1P
Unlv8iQwqy/X9clRG6X93PmflcQW/qBqbCG41sjiK3MMZavOlYdL0tbbvhFILpil
0qyTkKqM+fHcsCMjIIM533l1uzpYfzwEhpEf26zQGJ+eGO1vofsKJ+wJ5VX/d7Q7
Y8kJmo52BNJXOEwbxjoeKz7K0aJQbNxKQkobNgEywuj4yRrfWGUABZCnx8QXsz11
GRzXwtgSy74ncORROs7T3ylNR9aEGjs7A96XlczZgomwqu37MKLa9gv8LZKZI+nK
yKLtgVbhXYRrSe+MgDuKgRckftgPEQX+4xV27Esr0CjGdYz2wi6FFjXYV+E4q6Zf
lX+/nd41k3YW3nRnwm395LQJdqNSulY3CHpvIP9MeIFXWlIiKpll2Zb2sOFxF30u
/t9ONHJO6bZF4fbxc8//zfE2hl14UEdFd3cpaX/TOBYpKILXTAPpXpnOkKd+9FRZ
/W7EDKlkYD7HhQQIwlWVH8/nkmKJT3/sOvKtwDw3+df1sXWIOOvUSBh2e9QzJqS7
U75xYiUZen9LgUkOLuUHCI8lKKMeb+8LuUioy9MBlFJelMcmFHZWJgXHoT9X13vn
ZGDiA91GkESMT0/KOeoVZaUTk1TCxe4HCY19Zvj7UzLgkRFE0SL8QD20rGIyeEhW
pQpau0yeS5JXvNyBt/pXPoIfqerY5qMgoL6WI5KqdjYPD0tTeTj7t+v71M9bWqz9
m2r/txWf5KA98alPzxSUmP89IFhpvcfytkwnTdmMTFfvs8TKDRKfa0k78ke3M88J
CTTBuLTydskCIBlGAZfxWPg2tHAyULN2A79Tkpz+VTCw9TLTSqYjGGDC8BVPTAVp
eqf8uh3G8XLZzPnI+JV8aw4bUXRDhYPu8jvaVn7oiHazldQEaYojSWF8VcQ8Z/Yb
ObyySKwxC8rrziHQlXVeOqqQHYXW2idHIcY43k79IN5QhYit72j1xgjpn3j58aIt
fEhA1TqhxxwTTimx7o/fF1jc166IF7Mvd75SYsMQ0idl4rhyNuQaMCLs2OE55v7E
bsmbeu6C2H06e/jRXbX1II2to3M+wp3bhneZVcw1PPeyOWVvOakEp4VJ7J2UotdR
xey0LrWOVeNHSx4iMyBepmf8MWzsW26JF8y0mjepIDOiEjafTQVIOnndob1ebcnt
b2UaKtXzjBjdMx5gt1bs141QbXkcY8BwZyb1uHjl7A7egN3JzW+ANRViyu7K1wb5
HniqjsDi9ebCzLbLJm4ALZeLT2UUWNwY/TcYAJnat/UJy3SZ6wjIRmSqF8KoEKDv
rIaXhiAM6akLIjPp7uatZARcdw4FfTlk1N5zKboCaE5WqLfyCRQU3rcyijAB1q8p
rxWDyVEqkBVmFMD0nA7TMJFuATRT7ZSyn48TJ3IudhWZ5toNk761TCcixj9rcp0s
G7MUsFNL7nnWzW9fDc5umvJGIeRr0Ztw0Fn8Hkbj7gkVrjro8votAZaDIGiUsk8q
ebB18e9FIEUb6xLI103RVdWfYIH1VTfqaaPyrIOokGm7WHBzVQOUhS2Ug0kDcbdd
tEe062ODxet+RnAPazx2i4oOKs5J9pNtqtWh0ox/aXlLgAKJB/d3W1v455pgRmnw
t0pnU6N1KYGjPX174V8trfccwypdnjFvYKooZTeokLxSBzIrCke2q+46yl8NU/wJ
HnmuX/HPKEqbdi1v4nib7geLZpC7uUyLtuysofRZEXbYUtya1Niyzob7W5YJusEp
yzKkoVNtxxUclfXPvORQ3sVEaWJk13CoROdRZtUcSyTZ08onwHYwNSKKP+5MIuz/
AvoP6XOYrSE40fEN4tUEGR2Kv0PC55jS7B5GrRkkNPVDeJmYCukmY0nLfpLOHE3x
nLhGTecN5xgi+oXfOcCbECQtsS3A000IJAaappYSTz5W32Fz7TK28/GoqOTLpwX0
XjfOAMK5QeBut9JeuboyGHR/oF7ylcZ0QnKqju1bMaxkuXxF9MJa3F11+1jU/DeA
uBJdT874s40AFBKu/5cVWXPz+SS9t2C5YS1dPvc4Z8fdm2lG4RwCNM/gorrbau0A
7y7sp5lNWGNOSlNEa5Yiql4jquc5F82Vl3f/I9ieEOjuupADKFXYV48wn5ygTBzA
VOlit9qLcVdEytbYBBLlT7o7rcLmqy5+nrXRmaNyiqcE87n0IOp/TGSksk2eKom0
GyFwEK6Llzajbjyw3ivvvpQVcfne9+Tnk/v65m5wbZ46YZDa4HScnvV0A2cSHcGc
jbly5vlDJbkv7IIM/IZcYUip4vVn7x1wkPziaAYlWKFK7mZAzS2EoA2Jp+/NxC9G
r92KI84TKBuW75t0iToD+9qnR1knMG3MFv5qsVZ2dBuXgmIPCKCL2F2OTwbHPsk9
3d7vPU60cFvkl1yUYWSPPZjDcmoGEdjgEwTBhdst49gGeZ9VMqGJ+3MM90bVaAzX
6VyPa2AXcmEZigFLRbp0cwbo8ZHusP8ZyqNd5AkVshL7xhJcqPArP4Wo4Zjh7qfX
3m5ezUYaMCflYV+93V1um40M0hgx+vcs3nFNTMhqDeuryRvSZ/gzJjCnQyO/ebgw
I1O2/+0LeGUVrs13OxWvX81M7tQX5L/8oAHAUcNOvjpJScrqgubvvuBMiRE7rXPQ
K85Io9U4NdKDnRUD6XmArqAgwSWah58NXdY2rhtg6KMvs5AfbaPbRxRaPcUm6mW2
VXyGRyV3WEvergLrWtwqwBJ5QIFskdhUo3RDFwSijOcEuwFqVqWtNssyJfnP/UWK
fYLqD05U0eKA8ve87/iBcrF6bWcooRyfN+t5odTpxWIFNyA1W9A/5W8lp5mpWQgv
jPuSuzDvfMD1udyu+lEjWBI8/1aEBwGqBBxMoHvJR1l/M+Mq9YbCM7NwEN2XC6V/
D/z/zWJKE698nfX9MbklFUXqhPO7U0nQSLyfMpuPGP2r9x7Ar+NCY1XO7JpZMQ0p
jmeheYMMUDP/AWEV1MqkSdCTJroH8T3kABR/IbAngCZYU6d13FrmA5i7tnCveVDY
DVC4IGI1Bl6xJWnLKRZFC/dnJ2IXhED+TZFB1WAxHFDkl7svMojlcqy+5Mfx5QYx
q4yw44dQIh08yRkAU1GPiGrNT3zhMssgF5FGgx57aYmqb7npl9E1JjKpJoFUPavR
0tv1/D9Lc1FoeiUvgeinJMr1ZYv24ku1+NYFrf1/V1cMzAkJT4lPgfNVhqMLeF5D
gSVJ1RWX0FMdoeRWW5h0LuMP8vVcy5qvKFYtBtZN45tubB2rzfxRvrDnAEoZw8HI
XkFI20tqp5lhaDBMvjS2GOMs72J3BB/kH0NstMh6mPSM8qICc6hdUysnsz9dsN6W
Wa9+KYXpdB2pTi4BY4RGQRXOuFqqJKYTLiRUAdtev2DU7/h3+X7CYacJSCDIRnAo
5eCbzm7sFXuI28Pltjc3nAEKBLJoHbjLjbl/SlLrZh6S1J9cmU2tTSdTBRmDZOYO
ZQ3r0KkomQsyjT3kc2oPiVkWsU+yAGFR40cva3p8AvLNd/0JPnOpRTAgDZvsLRnv
GwlAj4/eV75HEQMDMxLiIQf/qNxqt1qizm6xNNfnnKGZOiOEvCG6QUP0yQuZN4UC
X+uv1tW+TMuY22N9C0ljXSt2QKpw/TgVAC3YBDjAF28D+NilD/dnuDNVZClGEKha
k1J7uNBxtOsNaYpLiFzH4G/Mp2K4yShu9z33Q/QMZAoRcWKTO+cdbhpbemW0HY1S
9RtV5AFj+93ksWNMFX7f+38Jt102JAhQ2A+W+G+HYmbP58YQdrMWu8Du4UuI4jt6
v7xyGY5CcMPaywz2pqAVf5CF7Q+KfXxHIYs2zeV8nZQ7Pel9Ndqqg0aXwavFzYOK
IAStX0rNYppmwmsXarYs2M39WZhHzOk1Ck14cPv2YQOBXFDQa1t4L1R/mA9cphxn
76TWgLABbhZKZiJKDy8Ba/71xmKvfJMfqt3/9vX3Q36e2BLmGeNFODQYK2alPVaL
Ku1LyqvaRoGMCC81LV0mMuMUNLgKdKMIybbZjA1Ox62B/qANB4l+qpGjKreR6dBY
MCew/b4VJjxpFVK1F/ZGnaJN/M6/DNnAX674qkSNPjy4l7Hi9D3IJidXUtZQl+sb
KXTQtnECYPWDGrSjfUTec7FxzUQgu259WR7dYmTaP2ZPRByXOPl5h0w1VkJzsEH5
TVRc88BQT1BVMqV8dtw1KO+vjgrdWo9Y3GRxrg2RFL/y4h8bOEzF7D4/SgLMuxpp
ARFwFfjJ4OA/fdfqOWaB+itGkU5GzprtxhIHkxC7VZw/JeSnHwVqdCV2llI9/otM
ipGEVaaqoBEHwU6Fd/TrvM1Cx2buZmckKOGLxmqAS0GvyJIiKSinooRBR5ScE70m
0sV/N6G3xUWm1T8q/J8pnvzn1IFZqntlZ/dQTgGVtI7+p+Z/fQ1h05lc5fL8lRs3
QUM1xOj8vv807qcVurrB9W0t7Gr73JnLTEQUMm/w2vyvom7snOeyL1CJwZNAlNsp
L9YY2A8Qor9DK/wwRcQHQQcJ2GM0Y+72Oxf2ezl8QYw+71ZrDuqTHLRygIS5RvkM
A+wTqRgNLbm0VR2Q1e7hVTYPyo51h1+nKbqFbNXvwBm/a2vQ9ubSOdGJWOhdJZdx
A2ugKeDPitTS4fCpNhJa1KtjKTHjh8abgg5mCSsi+0PfftCq0BiXgkeYMa7LVULq
jJu9A7rvc/fEErI2Dk8fsB30RDINkPodX0v9yCiJcnOgUrGzhapaT+CbhbFwlIh6
U5puKn3TrPUurvWSEEnU3i/jqQdCL7d0S/kSGd+/0ESANNOb6+MpuSsc6beS+oav
dKVQSOgs+AJnMZosgZyu+3EF/fT4kFIrFmk2JC3LtwO38i9iZViSbqcNJCIemY7+
nveILNp6wjKNh34nUI7y2Fc2CZ5ItvHh8Hb8CTdJ/kQ1jeLjcv7DbPbT7MHuB6cX
X7Gxq3PipU5GQfXqdM18/ayFET4cLy2hf47Q0oZ7PE49Wg2dKoUImhf1722UVJXw
gIUyZYJM19MFQ97YBnTOyRkmdi0vqIJAjJVQ0cNl8QCgOhxgyM60mN6BR6wO8g4A
VNVai3JbZPU6INKY3ot5HD/WcplHsDG0v8KWoQ+o+FgEwy+lxdglvM1UqGGkDqII
jlWuG+Izs4ar7dU9OtR3/6NeIj9avthRLXb5gAmTth6CIkd/CXfrG+zbN9X5lgpm
XbqgFjCYKz/o9RV7e+okRPanJVdtw/COQ5iwDNAOW+C/ec1ezVDO+We1u0jt8/N8
/19NOVHdeMyocP6g1KvZhUTbXO0MV+83AU8v/slsntAmv9oesGpO/JDrxObnXuHN
kuKbs35Qg+BFM4T7kY4FzNmY901L8LJZ3ZQo4U4JX0Tqo+vUXtIAjxMLNyInnGB3
izYmdAoO7IlKZVen2WlCJPGiTAUTZRV4Bvo0gFIyO88jha4X5uI+IxmRAjeDmI/b
w0hDw+oexxLavJCMJ5BOeeuFjY6B0JBwQU8quVGLDcaK9jWgUs/l6Ys3T/VQLDFS
wjeioO0tik3NbevvsQrSWPsOS/k0KzaZ+mHBr1qm0irUMlVHD3apVd12uD5++2m4
u74JFdkCABuaSnD86cgge2mws0fIO2+r6O2KFc4P9mVKbyX6Mio4F/ExjgUO3JkF
yeEV9U3MnXavLs64RAWxJrFR3+afAYDRM5+osolqedZpf+ytfNlj3ApQ3CLobNMh
Mdle5IulGejT8lixS98sYRgGYqCz4oI3CjBHoahyOlh3RGB1bWNkewS6vcRVCgco
+Nj4sZFqn91nBZllVBRLu9wdZjV7eSucKkpdD9yyvzNlD/Vklx1bYQnNH0/JlpPC
QpXsB/Gha4GDyItMGzUUykJFNq9u+uOZ3XgIfbd2gUI1qSdM0h9Tpobdn1c6kX22
CmmcUIu4jw/gIxk7Fe2eYfWN0T5Trc1Vx7MY7BTT3v6y4DRyzEOUBpIPRGW5GxjG
npNbbjdffSnIUzoiVBqkQOLm49iPq5nWhtTlar0NYsoVE+3jOPfoZXhQUsFw5XIe
11IfzTrtrZh1Mq4s2ZMTcdq4PUeqqKrraSydOGDl6VN4XIxjLj1hLni1ef8AzuMW
LXB538srCx+DdrDaadNsqwcoSfKUC7pQ4mMp0hnoZyVy5c5BIYYhw9vQP8gHma4y
Eyf69Mg4QJp7OXdL8hxPJVkDcAcGrhSITNKCKOcjfcyv/tE+/LmgC8U5njyoZ5B5
W/HSkgyKX8qIRZEzZXT7HVVvkHrjuF9RHery6o6ro2qi+Ng2yKFDVqCdI4Mo5hcn
9SX0mYyYYX9bvE7qc9FYsyeM9pwtSevYM5vsROZZLrueXqPH6AO75n77p4A06BkE
s15htH75mUre0woxgMTTKA8m6NxpIRRcxiSHEmmRlCY5mLQ60ggdfIMt1sDY6EiZ
SWu6xRP7Est7o/kboh7ARK+1K26YY15VvkPzvJo8G64vTfWMDuoeU9QKMEkjdEeg
DsY71frg9zKcdisYuiqZyhb5PidDKSiDmNNEQc4+o5tHP1hluEJLLGQYUsgjsK7Z
kOcNbY64SECXACTySWe9AnMVpluTdpNn0UKv7GROyBLXS8ZW+MDQJ3pwFKfOLcmp
frG34U7PMQHdsC7TfnvulQGegXN9wPCHTd2vae9ZobbiVzRrxMLvN/S2pjC/zzrm
pWzil+7TJxuOIzaA87Nd0AiwUTyyHkHFEBdkoT/De3fEdhl+KDBOEpjwntzruoif
zaqkr4+oO17qlSad748TG+oXSoOmnXJD4Emgu92pmxorJ+Pbq08SsrVEumQl1/v4
+KEGXWN23VjcKNPQseyhqSQ/HVazIW+4TqyKHHFbf16Nu3e6tJmyl0vy+rwUc1h2
BJ25n2H2Zrfw+KrPPQnrNujhsPsHhYkWyzFIJsmZ1TdDKmjBDDUKMN5on0XB9SoP
DsEaTTqQvI37AD4mEKILKQ4ct8DJONbgh0soUKS0kiUNbgTWR0qJc0iweEZ0OR3p
4UDGfL5Y8P8SqATi2WjxEQp55ez04C7maxYo6re3qycFHgZj89LbiciU/WWl+lGC
deI2t5YU8Ao3ewm5dd0xaFG+qr4m1NBwvsYr3YpaQnRvnVygsUKYrdPYd7FZwP7X
HuXgcTmkspxGiYWuJhkS42V52NT6HgKZI7JF+X+BsaAT39PU54ECKI12BEt5rA6t
kIAIQImhc5gvYurBCeybw2fCB54OCUm5A4ALpMCo4Cyr41MwGJxdolLWP0rUX0C1
jGro/SO4QDuyF4+B5gXhL72G3B7mAp1lv0qkeMYb/LenQK8rbo5zaELlYhAD6sZ5
5lHsQMhOt4HOAroLVSDN18M/7Y2mELXpwmkRDqiMbqz9xE1jbB0g2lOeX0GzcpTB
tcxjQP7JmQMIZS1YLq1JhivchrZY7HVto8z1VKOtktM9lhAzFc7fZZJD5/gSNznF
eJQoSowcz9PJISSYHW1FGEGuzAttblv0z3pL3u4zz+Jw4g9w/nW8WZzmKTbeDGei
TFDyz0XqtX9Ck+a/p3smkUGlmpEYYXeNVyq1jyECVoCOUzrhhCl2DDDIxZrNZqnf
wcBhaquLxQLO63WtVxR4wnCeLLLynoEFWgT38P3cNQbgdNvuOUC3gTZQa8vNJRpx
O8TEjkXczdmtZu3A/lJ5rYgyKrcZkr+ClNT8Rw9JjfhvYP21vvPkYGplPsXaExiY
MM0zSqGUP5oNlwxoelNTD9YMNYMbvBJAhBNxFa6am+XFg418MyGpms2As14dh+MI
QTxP5tExDwI9VCusxKQtV5grld1ifkW/wDbU3WPt9sBAm+10Cq9RoztR+9s4V+Mq
mjhuR+2QctBY7aBkicHYR+0md2olNlQa78CBjP/mKz+n2KOHAWh++5PtUBJHnaVv
xw9Z0Us/WBGmdNrsQTjDxUz5X2vzaBRjw4981OOcq47k60IVc9kXR51uwzzhQAwY
eJT8YVIanEFQpW5x4BRbuiq/5HHiugJ7V9OddCq90N1P68xd4LvZEoE25ouKqLW2
RODYoljh1pNHqY9w/0lFfOgYbZNr9b/4JbvJ2WSHf4+heM2g6TnOYmRi4lHls+T6
VtaukQ/1u+zquOo0S7vTi203Tf41mvUqguN2WjfARj7zuCDCdZTJwZbeV/RGv4kK
GmDyONE1ltlAKC9Z1gANftAICwrhXStj/KluBg7vsWyN8LxYbFJ94w3+J81EcPVV
fDzm2aTaYlPAMsxc4QNuPw/8FYEsvuM/kLivTs7QblZEsr1aNu8nSCqnxOXFqoOb
wrIgaZvS5XfOmAHVGduuvkdqgM3rPV1Q1MCpbDOhP495k8Fnk/vELj9I2Z4ykNfS
0f27tSvSfh8OUfv/ynJutpamHGy9GuvLVbv8+VrKCxCLy6Ju4kFRKpYf5reIJEy8
yfQAieSoAw82kZcdsGqJh8wAv1LA1Rm/hQeUMkrJdJqWCbS7A7tloMWxrLFhWJui
mPuakNN5FR3RvALR/UjtWPZPp16b8nw2qQYIFfTCrdOWe1sNG0aygRfWzvzZciGM
AqLVybbplxrPlmkXXnq6ijHo9lNzUSu8R+2JFb3WVPHGfCPj5roN/ywKECdvDop5
GEcvMGS11n5Bcg03nuKyRBYYdfKlG9dRf2r35xVoXhh6wO9UjxwwoZwtJa5Cf9+G
TspfezqqEiyxKexvVpNeac0YXYBJBI+hJZ1yDj5jW6d82w8Kmtc6eB78+gi/6O3G
x6IOUhRL+CS4u5iW77VhxYK2KZOf/3V3DsTvT4UveYFn9xIMSGUILPCYLQcM58PH
FCqGPBIp71iOwujIY+kfrKLm95skv31+mXdvx7CbFyYOHs1uTHCNe3/dddk/kXHP
GzMhZQyGveO8IWa5aXpm6h5C3O2QlUD5H/0JJnRZ+KwdClNL4afyq0ZraNEypXeJ
IcNW7249mnMga8r8KFb9WUoCDC5bvPk6t212BqGQns7tYQ7Od0zgSzj9MKJXsX9k
Izk8djV3Ot3FHhsYnpMJxXuDGpYImJiBOye2D/+TlXwQhhfphePSOYxZOGHqySGq
eTrpG/mNheAwpzFZwEUV1+yzFqe+XnNzyOP9sD1d/8AMswCoucTAPT9Yn/ZiVmd9
lLwZsnCWadBZzHTVjRI0/i6FUdMDSwxUp8TJSeyFLgQVNAaEgD4TlLIMkIxcJIU2
p7bV1JnjLLOEB46k3SZujYI3a2xiYmL+g54/qdTvHLcAARtmtCOysnjgT2MNhZR6
wWm7X6wj13fphY7sPG/bVTcd4J90jeNfSU9WPsUn3v3rTByRuu/Rp/UJ5L+I/EgZ
zOZJxlgFMg0jUIqES1FneHaS1muzTO0Y7Qfh/uP9wbj0Al6Rbuhmw3kKugFlvxH+
5iYyf8MXXOrX38uWaeqJDCfXirBpDSXCC7IlmlyZVXaHoMMtR8hEK7oV3aELN4BS
pLxfEchsHI3wihN8GSWx+IR69j4WH4QDb2wC+il+mReXdgRORgjDROG0ZNdr9db3
1QcAoJ2LXrS3gBKnTzpbqs/MG25eMP2jINRPhuTdu3HZVUZhn9NJKwNCzvhFlKgh
4GNhOos0nJcmd6loFY0cSCEq/1NUusZGTiSO/hiYyJM7NxZCiq7UsGS3iLcgB49O
gRJUob/yVMblWXBgdRa58IAYCIKg6mYnVtenzdaw5qtxW6XZJGzrmsnXRfJLp5r7
ZCPvWadK3y0PNFUWvQyHcfHgYCYzDd86xUQsG3520FO0iBzuQ9adxhEbqzKDl0uq
X/c87UnYquOQJBlGg02KM73ndnE/5qqsXXSg5sSzVwpyaDZSnqujs1morduPVlH2
cT0hjhA8RhRK5kLRFtDLeLg+iMRoGdzrWmFh0eWD+5skRjJbcyQhVKd5QwUy383K
b33Xz3guLqEgg3SstnElTk/ArtcQ7HllD7WfU8gI/jL3xgHffHT6oU8Wq9Iq9Krd
agCP4cesBOBEDqQFpJxwsajzCe3OMKHwTCnbsrLqJ1JxQ7so+qvrPGCx4Yz2u9A5
rg9tKcjZFLMePIdze9n4jO+W9wGanBJL9B5XUPN7XPHzjeEzHAsjUZi3h7D1FqVF
Nm8uz72O7VoUo6jT2H9s9vsYgjGhp/8/5mhjEBK6ReQkj56rr88wXFihkBFiRRx5
eTm7sV2AB+ma0kNH11pvqWxJKFhmdKEN3acFYPhw2ZqHBtPkv6475j9k/SkdpqCJ
ieHPe9CDyKA1fG5ipFF/kglhrrqTFuJxb8iSARfma8TBeIA4TGuSYsmKj9Dr/MWk
3nH4a4xJbSiSc3HUMoI3CfjYc7ctktAOdIt4g4JdDkxXQCq2l61pg+CBvUtMURra
HtFyfTI0zOl1iVBbB4e6GWYLMDDfbAjhE/a2VBSAml5lfkyeV9iBdkVS5JtdLvc5
QCE8zph50TaRp2yUStGmKxk0DyjgTQr/hgoJiqN+MHDWEwHlHgSI6qv20CAimX/Q
PjODyPtw6naHGZQo/KF4KScefbfMnE8yfF6RuQpUQbi4vBHqSqfdCpfp2dcMmoQI
yQaxKsRbCp74s8YNPvKJyYi20FdJkf+0M13o0GLoO8wT/Htj7l0PGn1N6dd4UQq3
YwEpHtQZOnrrW6yn7F/Th/hZ18I2W5+f5hPh9n/9QT3kp2W3w2ITCbFKUfv0Bki/
usGnxqWQRYmgtzYUxBRD1wegVepa8o0ElDhzChHBp8JoQS3M5V1m8tiNWlSYBHff
t6nojHZX3ktDRK68TXwUFwQUt1+/SWfFVfLLo0OVZlxYZzRAOn/XaTYW0xcKCq0p
NYnwRzHcN6p+g7625VrTtXvjzQ1NuxJyRy/hJUikKPKxzm4+E8iVF5vaQ7PeOHaU
xB06a9pluLsdX9GFZ8GFGsT94neiClE5FhoSOgILhw2UWPFiJlphTBQ/+Mmmi8sc
Rh5w5XYCG7ApHVw+OyA2yIrAnDZAJiJuyg4WYi2eMCdLuP5/Q2RyjvHYqZIabmhz
MkKIRCsh8UKxYcQbkzWJkR/SY+pVlVdYK+9zfRRAGIEnspVYoevL2tantRCsEDXo
iYM06IK+Y71nhCqsvwXgr48WujgzWU1WIHookF7zoAqOOgZbuzwF3BCUelKIxQ17
WinVybZSDY1tTVjWY1QyfL9uEltCdn+ulQ+52rM6dvBaQqalbeuiEu30UIuweZAP
/GaAMjMTzmD/h+JPKzAUYZMufuBlgo4MuT9tkfiJSIv3/M3BHa4NFUKh1u4wJqmH
j+PrlMMJ3C2N+KP7451I7HJm4SySnE/jpYqyjeehfyEfNQQPNUoOK19lonfhrqZ9
TSArAHBiJRDMgQB7vMD/Uf+VUuFv1MzsduGiea03VSchvuYgNcJdMnFQRQJ3NnAN
3tStK5fMSs2ozrxygVa+KBtkB4WAz+3ekztMb1Yagrh8KHwu9/8sUykGGFEYyi6Q
Udd2MCscftGHIvPCOU2O0O+5ycY0MoqcepvuSTeTC5RuLvJSp5+OH7Uxly+Qj2WL
mEuYO7Ud1uF1nsnsTjaOnVcLVUZlzWDOpIVHNNB6Uy/BFsbqWmwHehANFBE1sFlA
5YHXBv37F4gy4ONFujrKVcm7Ocob1E1k2keXhbxEz6hRv34yVm0NBEbxmS3ARV/y
WnH5T0Arzh87/j/cCJSABCN6BKtFVXLS/JMZPt0Q6R3v+N4t2WorE2l/20tqZkwb
v/aXop2+2w5fKNbPvX7NAb3ZQ2JPyZMc9QN/cPcNQAe4oK+oYkqJ1qoNJrTPNrUR
x5afkXodUMypHhyer19rb0dOjvaxqpIaB/787uljc6QfObB43N2pVfgxIxxD/6WK
2tTUj1yhf25qWoRjXSQi4C3ER606dvz+Yk1txTeXuKsMDXpFwlAbdwZHAHBCAEuu
714GJpSz3b7N8Rniprbkehz9YEd3qdF93yCpoOiXoJMLATxeLyGAV8m0i4EZwQIR
gHFukpYlLoFiPLrlWMhNoHqcGyRolJCOBpHlKha2I9CLzIUTf3L6kylYdCXPGAYW
AOR4vNpYrhSBpgkIDDxP0/yw/rdCIytaqbz/VW5PuDIa5ojv0kIhHBM6xCfMWiND
8H9Ckgw1UXC+6gFrEJ/g8U8zpl7begsu7lYDagM8+tpo+tUCwG3ZPADKj13ATiDA
zQ5LyhHcsRA695QqAHuG73TDj/VctPqPVQMZishr87dZUgmdQe5Rul4u8RRgRukl
fgKYNiLTeMPyR42a78ODqN8C+NhkdU5OM53xpelGGI5+Bdj+jpio1ZyitwfYdwR9
wORqUQ5cVHw1Z+So1dBY9UvPXHYJOM5dLPBtYTV2AWQVsHbPZiVZpbBhukAAL2gg
tnDepLimbG7Tu5UPE8qsgAVk2NJsMEin578ZDf3kd6pXHmSd9hx9NfYh5KCXWPqz
vI0wVtVOlEnm8YlA4HScbtxJTU5YGBdTUhA1RZXoxvtHt64F9MNJBmGS+NlzX+J3
p12pkpt5taGlJGJcQkPoV2HVAPaioJIJF5cVQ7CaEkJmWPl9BC+lmmd8ZEX20+rL
hIPcZ1K8FA4i/JtTHEEfWUWApv3ANIeX8h1BSYQRF1gz2hZghFD7FRsFEHw+0awC
4Shosnqb/2FsaDZYzatzqqtN/xoOqe9nmjtydlgs+AU6kJWOFR1dJW9lP8BU0eZW
0SvrRFwEfbOt3tsORW97nwBXaW+Sm4cRAfnn9hvD2llYTIYOdsU8Ib3enCD5OTJm
mhxhAJsgYXmRkOdtxwuQxTPi23/l4LEKvF6/ONJJa98CXkHR6gOJjfXfzHETCLLz
cYft5Xpq0irLUAC/eXA+Eq3I9VpEflvB5Pv/ViZuy3OmmAm2mhqu39A83rvUPSxx
wSg3//Q0/AigR3VRbx7uiDqXwSKa5HcSnhN9FkQs8nDkCxPZO/7b/jmHZMLnbN4t
xJyQu6oJf1zqfXI3eax8vtMgp7m+Ugtwfso1a988Ve+F2mcIEN9XuiDSKEd8d7LR
/856n2R+FhczU8MspzgoBA/lw2wPk3g7YB70WF0/BpNlJL2I/8J5BESUnYbjfpYl
gchYscwUtpBRU+XP7D5jKxvappI07em9e/uHzCvXMN1PRsWI/2TJaacjYyBPWFdF
SY+I7KzMQMDejBOTuzP7VPU3yNSK2/GEDS4CIgzFSsOuA4/tXcbT1qZ2HKsJ/m1d
rAhU0BzAKJGPKk6VKjc7AswX/DsovpJDsW7bDsw78K/ZfTqA8wapAvhorWlR5B86
eWfwAhwt+otKUIXknTOX4M9/6WN9BDITMt8oPZqiwYfm5+mGx0AMIj7thTxXT8mE
O8hgSbroSse3A5Cx+sndEEdCMgigvVhh1EE8keTpZAHeOvFZ/5M8zrOqvLbl+9Tq
NRx77I5hXgSNRBjRJ8NR3VYsgtAgDgyhz2CzLQig6Rz9YMlqM2keqGVsjMngUjuQ
blstq0J0DxNjv+1iHxBZWZR8dyZQMei8BOQSgMggEmawjM6yYLNA6XXTlDft7TVH
011BThv9rT/XZ7q4p/qHFqjx06AwIeOWFzgOOjxYLUsKTdsd+0uwMZQZoRWFmUce
XztcQz1kfoMMiP+K9sooo9iVV/5LXq6RZD5tn2VwIMwuQa3jQIy8Y4S8ouIE4DLm
IbQG8OsCiqdwD2qMYBmEXgmKFN6aS22pkTnhxiUXvARhpJP0K7z4Dt9JwUzL2KXt
bH44edtHxZAByikyscvFl1WNQxgGmBRIg2TKGBd2hvFtQNAXO9hquTg+ofAGeFZo
LE2zYmUOb58yesMvE7Qy1tl7//BoyvgND47YMKBWVSX0dH7EtP97JJ/LNGTwGKbt
emDtLiN1aHVYZFr28G84CDzQqiSVrwsNDrKX9wKH6BcvxQNe0Eu+p3nPi+7iP2BD
7wL6mDbDIG0N2FZMGYJ47Wgiu00/7BeDvMH80PyPkZAb4KXzHi7g0QMXgSQGD+et
C3GT8v18vSVyrA29kcLUIPXRUt5jd1wF6k+J3bKmBxwBdnLwIQS5+NuIYAJ181YZ
ydSfiqZBU7f+yHj3r35Crpfy+h0Q4ozMhDk7R39cqmvifvNU7W3zclQlLVwXFhnk
Y41DImBPHRz88Fp6WO4M/5pxu0pM5QmsImxjB5/ECcQsIL4+0iZou6kja0qlVML+
L67vysxtkUNi4aQiyVJLmfNVW6eJMdxvxy0AhmGRMGM0/3s86Yn8AqZGQ67t4l00
Z7+31dBkKo9WZ3CfXQ9jWAOtVl6fBNp5JnAvuBSxkai8O2uV5t91XnvYEV58s1Av
nosMEE8tWaEANB3kEbuVY8sKghzsDKTU/ekgK+xwfl2KauALzOb4QO28po4F9LEe
Jg2S+GwTherbSU3NDWO2XMqKOoOOevwmj45ltgyM3cgym1GcBeczTMFXVoIREuWe
WqG/9sJHltOz89FikCPAsEJdGA6WNQYG6XakOL2vJB6BDR+w5ltp755tJZjtjm6+
FPzUY9NI6Sp0G8HIeNWGjw5MEu4qV5GT8LoZN9f5pnjcjDbp4iErghUmgDKHqc+A
erWr3HQGb3736BaUkLLvznYOe84dby30b3XmRsVcCajZgHd+yphcJwtsoibkdRws
nNnpFI7nmlVnYWrTB0LvYl+UmKSm5iBR7k/A92l5Xv3ogi4nSkI1NQtN9KAQnJb+
ykLkLL4pJPEn80KQ5XxNfV7nH9c5alYVC/PidFG8xAw5FlPZljusS5jP9PTWy/TD
u2SQzztiWkQGxcAgm1r+foySyTYlLSTXDRUPm/pCVjAM0UfVu0Dh0XN+Kbji/LcO
F+vOA0tqay9ERNtoKj14kzkkxZ+OxCzMh+B/9zw6bYDJfYN9qNyCsYyT5p93PBFS
8MpW/PEKq4iuPZLtbcfb/MxTiJBcDddg8a3Gmgfj5pa424iJoQzzv9pui8xcuO/t
IVvWUZGaPj7MYzI+23tg1qfEt9vlrmsJIrxYtZvQxyJ9JIHoTgv/DcnTClkkCost
5jo6G/Zo4azQUiY8NBIYN8QXFoJu1NxCxJfC8L72sscD9H9igFXmZbgvYkEAKRRY
g2yGhHLYHfCuj7FdP4zmPoc7CyRG8oZB4IuBDDd8s2C60WOG3MKpwhiEFKXEgY+p
Av/7ixVi07MIwv/SYOihTa/xitU3WtGDi5/LF9Drt45d7+/AFB81ydugkZDQBWzl
EnJ9M6m1zL6MjgtbnEs0Wo/RNCNAeb9OVzPVnMHmNUeiWENzCI+kKhJhO/imQbcF
WEURy40Om3gr0ljAilwKyFxrxnIG5xfhANoCpZv9uyvAsf90d5IoQXBlmpZ9rAQy
cwRMDgEg6CCgPgYsSN4yyIUT4ZpDu48YOmUE/RB/ruN5yfMFxn1l31uk9Pbydt/s
2+fcuHAy7MgIVpvn49srraE8z9m/TaBnNprBl6HFzVuJyfoAPfeiWMICCzy0oi3B
UceukK+RBo4Rb867JvR637wbhejMtx7aweN7prAKop2xea4an24renK0HlbnurII
OU7PXzAjHJHWHYeFX4ZJs5P3X53H2oIYSN+DpRs1f9FYu50TStLAEdrf8P7Kv6O1
gm+EaYL9eBP1ftf1Dp3dtbu4aaCedZyE8nEyPxIg8Pn4f5id7FJY76OpJPjdYFvn
tw5sjEGLanWe1VcSzj1jSwhHwwQNnWVWy9iSz/OV0fyIdT68q4qQljn6/KVY2tpb
G3ffyL23eqcYqaVCWOTw+cp3rdhxZOsPV/R5jLbMxMsHG2c+cYO9DkKKuLsWaNFG
sXNSzwFlg/Vcllm/jiJEyk2UR8wkFAO+4Swe8n1pFXk96FAm8Yh2k6Jp43hMiPku
pnDnbNgsVLXnq1uknUoxT2tnlOt0Je1YVH9zni1racd5UdnHQAJEfpS/BSARKRq0
TucGuF03Q35R9tb2f4r/GfbrEizRIqVQUls+LU3wednUM1MoDC6LcbwLkJgaJv5w
1xMQ47AlClxRgdhRFxkBhUWo2ti+OTKGZy2p1B4Mt3+0ri/fQwaWajtQfBFRkGql
Mk9avh3kA/R5AiaHeix7pTxcTLQ/rnba6hfr/i5R4BF64sjJqjCq2dh+leKcL42T
F/33Z/8O4yWd5gah6/hymzHkDUYxPUaZtxNrK6Om6R+JYKpajrECfvnkkd6vl4Ny
3ZwG3WVgSYP8U9IhtRZJiGzGnIj3WLEiQVGQqTWgyTniPBYmDV8SN4/xQZMeXEZU
Rlg7iUvuZnBYVLlBHGc9+aGUER7Z/ytj1UXEIIC3tbmiXVP9hDuZq/88jbIK21JR
UZq5XDxzhfsVYEqXRS9Owc2W/oiAAmS+kTZ4xPfzIQSgCOyMzFaqqMgbVNZ0wepd
CjCfXIZOVR8D7rZXRwotUT4DMzDyEti4O2VoyyXQVxj2EePTqVDrtcS21VG2JyAi
OV8sQoFonfbQHh6mUYowOKX9RF+eqUo/F9dFXLH/CKz3IhrxeW5EUujI9aTQ8ebJ
bd4oinMAYMm9M/8S+iUO1wqgRjyDzeW+OIQQsAe1nUSv2du6O04VXBs1Yi1+tWvs
g5ak2h5X3XA5fpwtEoKv+pkmgrKr4+Jzrx7uo9drvgT+35oU9mcG4EPpmX7VE9ho
OmjLEwT9IxkT5UieSQ7m4U4l7WPfaB4texeXxms8aBEAM1r03YpNOMCCQn4H0ahB
qhfWaSBGKiz33OaYpkgmFQqhN3RD30jighbD1RKSWFqwzqZLEL0w8IgaIFiS3QDV
T8JHdtXDPNfJpf3neiEBj3WP3PPyARBsmNnXLWZL6FHbA+uoEFMkOCGuwKIouZ8Z
9igmqgM93bBhWr4WlME3zwygBGi9goGgDUYqlNvMPGvO3G/cJBZ7hLSH9wGPW/iO
M0D53K1n+ZmcSHeFAXMHCxZFqkfB64q0f2/FwkzNoDgvRuH3RTemOiE+VRfTqmDq
XA180PxOiH2YXb3f0+KN5ESIEbEXoKN6T36BP+l/KqPOQnnP204q4A9tXuSWqBTo
YGGnSZ1RMppjHl7S55Yatd90Z3KWaKk6pqL+dTQn+mwdrchtoJR3+LU/JpYez4lC
PXCY/M0EMV7Gt21KEEcH/ZW80XAOSLCP4YfIDHwGir/3gPuO5FhLPPPFI+saEQrg
fFqCkiD+1M6yLLYIz7SdrkrbqqdXofVEx3CXoY4kKRBwsXgMre7zQEtpYF0inrkb
dvaxw8OEDmP9D/mfjXy/MZFwlQEjR7xrq7jBrkxYmjbxtTONlCstGlVpCzSmWFar
tPccOZ4q2RdqjewACl7pW217XQ+e8eIgfHqY1znzY7BYyTIBgEQMRmbv6cvqyLHK
OkJ2j0/Y1x7gjRd56U7KxHEovg5XwrNzj9BqZhhJEnQvn7K4vIkrqivnspBX9u0P
JW+vCrrGkdnuwF+zrBnnoUX3v7hfb9qS+dh6xUH241rR064BFqBOuFh/eX9f5ZqA
D2sA+SIEgIRAOsNrR2n0lzGPQae0WdhFOcV23vXrN1XuAjhoBqSBMZK+yBML/gLg
jMLKs91VMp8ftd2aFc0fTCt6EcCRmtbHqtjjCkO22d8i8d7hbKwuqCJMxjgopYvj
I+qWkRn3a+Nu+/GDXCsVTYR7PV2G6mre/3HT2bfP8T11NFx2g4aEoFIuVOgxU49x
+EwtyqFZsOCr7b2V4kIxx6lpv/hytbGAnRmUnwICYnM+FyddNWaa1TFHrI4V97hX
KrWzFekSN7cbv1k11JhJHigNMBT0J8C+pvb28Z/IgohGM41yi4nyC4F1zTo1XnS2
veB9vulNE9LwWkjD5Z9XWHQkKW999La5RZOT5QpnPNuyvFbtTvarOVjl7XIWmFSS
QFeZvHLgjwu/mSJaufSz+RE/Ws2l1HJPJzQpPDyqP3F5iFCZYGs0ZyQtHWBDCDrk
ppr/V501WAX2YCdY80bS4E8edE73d49GhFiWamhbGjCF8gtK2WT5lCDyeAFDx8Ff
t4Mqfy7DcOZEIxF0y6D1hEs6NDlNS+G+MTNmmWlj74HdF7lC59LJfB/ICawN0oKj
dRtNFsdTi2I9mqUzF0lzlPkJ8KHVplZkuVkh2yWTXXTXLKTP3c45h55630in9MNP
LAJqXVaVTWtEjcD15QmHEMggcwc2tLDCQxcd3Vuq46HMiehZLtabl5nzxGdtR5/m
iwHJXo55FUWU98u1VEHsdeSSH5vFKUtLb1hg8nu5zsY8W1rSKCGYpxFhg1qIoz5r
VGIs/LmR+xiIzEhc2mJSVgBO5foxAnk4rl+ow26EbFR7I6PzE1X8rJA707mwRB45
oYlQ0EjoSAvL8CJ10ud8GXAcGp6VnthcxpSB6Ko/Z1+zxWRN+43Yzrhy5o9SahSd
xP3KuShheXv5mpHCsVX3PjreZ1rGbvBpxRVsyeomIcB9gBisiKtpqfnzdOo7xWjw
aJmk6daT0PFpDLGoEfv9f8VZxSSZV9A8i5uboGrT7b6i0dnJTdIvfI9GtL+t/OKw
GpbTrjHLSajw5SVzTJW3GPWEOwZYKy8fpNRFx64bYz3pjvJOaoNMxOgt5NtKeeph
UL9LWULzxd9ppkTsb8vlUQc2VzIkgnGMFLuDIylOvDFIDOJlttiQ1crtB4CksKaa
zIandHOYQknyzSyC4lVQSTiur6CY9jeJ5gXfO38AsUe9R30U/uzej8lUdUXQG5tB
Q5xXPLlXlASthORQuTrPnRsWhezkIHD0YvpjGlcdbyYWstcs/Enh/HixxM3G75DX
TyaRjgOic5iATMoe0uV2M8lFtSGPM3LVhhw9+aqtlidtMfuTcptmg/tg7G3kZ5jX
jmSv6EW9JPhy+wG+pGrBNhbIoDg1zkSWfkwo5FAzmSe/8LAwZOhrqzSXhzcrDcyZ
3/XqJOuyQNLf/4fYFV9HyeMAk3ebHmMQYtqVK07RJP1A/Y5d+asL/JldsewlNf+z
sQW1ZDBx86A8Swkm6pDeC1s/M61A2z2Hplp+gEy8rpOE5sHugPaGtyNi1CQtiSr/
ZHruO6CXHWaClb7E5c6I7ejlI0V+wEFQbrs3B96Ztt3aBcTCbn4AhOE0o4TZkzlf
GHmiZBkpc3fCU8mzRbyCdO7z5vyHFqDRZyQpziJXJfQdH2nfCeObQBCLKgSgi0Or
xzU4X1CQKj9Y3tYU5OD4VoiTxfOLyiOv2nASoFVUoMIzEw81ouyHpUkPnOWSINMQ
IudHLTIElfmz7wVYSbC5TDt2DH8QJUfHhY9Txk7ZY6xgptwmUSkkrkRG7hr3ES58
Z5CNDQHGZWLWeZ9pNTZ29U3P7HR9rlHrEmJNIBd5Wz/nuSZm6Cb5U+eEDlXkklew
hbGbOD5cIByDMgM6M7Y1JIFN0s6Txmi/byPJdxRrxEwUdzABNpy2u/2wxxdjn6bw
mtZSbYCjFgQ9cNIAAyFOu2lxynkhmLdtD2MisHJJpgA+pErwmnu9I2JsgZwo86Vu
3UQkzysaEOb1w1ULGQ+UL9gNmHLTER2C1hA3VeVA89svvN7ysWy6J4mQE2s6K1Ol
tkjVgg1L05j4Qohi823lYZfK3uEXGaFqGFHrARsvpmu9XaZIrSu84ICI1AXAfCSE
g5MayghV1s8gtyCkqudTRRPIKYVoGzXu74DU/Q4mIoc1upqRtGmicO6g45YVcwo/
0cYiJRCE0Ry9CMjSrLvg7d9uTf08KT7V1LcpTlyl/z7nUrYcDPhRt8Dz8J5IIkgt
QU4NpfweKJ1ilDlNSHnaV5B8JBhUbNwGt2/o1QAXZBY51W+135mMpyUD3kpaiAgZ
m3D6GMtBGI5lZLOx/JwyP+opamO2MBUAb42NDsy/+fZCj74wM3uWWMFdEe4R+yJu
OIsJOy/1yr6FffcGcQ9ZNzLw32XFSFjay5HrxL7sINEb2zE7r3A4owtOr5eC4n/S
/id+0IFGkrcrnZAuIn0NThGZOEQTV/rEPhHcBIg1sf9+qg5nfQ3N7a40dM0LfymU
7MneQgAqpAoXz5CvnjRuCjY04m5q4kydHhWRHoZ160wKXe/mkygNoLlH+5Jc/tvD
K0Ns5SlE743Vfgvx230MPBb854/f7ScTN/AqCx6Rh2W+5EDrmjTYZR19HGw1Tv6G
j3Y7CcFym/ImEcpR5AiKGNvgCmwGn+cJ0ooIt2KqXX0OS9reqw7lk7wW8ulrUfHe
jQLFUed2w9QXSr4oA7afwja3F5hfupsIccSuayK+6RG4wJs8Mp2hcmY/4lxFPHdY
zeFYQOdYFVqnL/4kriRMnrpfGhF6Jc0D/UwvJQjWWui3/CAp9UtmY1zwuLI2Rz9+
Ep/lDDrMXvMVWupsmUclvk+HUBo/YLSvdLbi1VbTg8E7VXlqPUhE48a52euaf0Ka
xKQxvAhAifZFHPXFo4OXdUp16uOSd0EVSLRuQnDSCzwT2QCPAbWG1bKMQjcuHx9L
PY1YWfjCl//YgaUnf5l9sS9UbfqtCuZsM/PJnqTUOZMLNm4LBXDVBgRZ6UVNuGLd
9DgYZctM39/sPYJwNaadBB4ygwZUlXEaCZI6mTEGnZvG3nsbl3vc4NRIOVtCX4bU
12J71eP/fET3gBi3SQ8SH66ypoLsXtBppwdTS+/hoL+T+g+1k667FqTgPGFeUGIx
EkmiKWWEFuTFZWmC7LYwQ6MoYmfNf5TTh/4hP6cVNzrJF8QxkBEXN0SCzRBCy3lk
FA6Ntevv9pzkPxcRYA103B31Zd0kSJNAo5i6HwpTWTCtHS0u1yb/SuCzO/SWZ+5U
dFNft48REVTlQ5nOccsGv0H++5nCZ08RPt0878K4Nt8R5VYYLgi7YuXeOwGYw4UY
QHP3gkoT4si+AIcx4H16uY3LcPcu7Rnf8vtoYgneO4MC9Lrng97b+PdSss3erxkF
LYkdIMREGUijVd8Ph5RZooZt3a9Tcp+CwZ0Hm4yrH9LO/674ubCujkw3ur+6QikQ
UTnq3vpeH55OIOVz9HytKsF+1WkZ52SzEM7OhtOILA54OdTSCt3RKZ942vrd/dDN
k358HxKTXWSx8f90EHwo9i19SUfl4hhABnanb1mI43z8L6FH/R3OBUnn8cpN2X7Q
+WMXo7oNaMpvWsgxbKtGV7rttQPiXXxTxcfgPNSm2o82TJ23b6Qb8FqwRhQH/r87
y9qFQqfbMT/2nqXt7UqH4SHSmQdQvEuOjpGUglokzsERNxcCeoWKhnSHEsuH/1XT
A0TH6yFfXJsEbJMFTvVIqhmNsqQuWVsEtjrQxaxhbHn++8pwjljMQhaSh03HogNj
2D71Mvzafw0xL9lkQrjf5+hf9hENoBcO9VIh8vJLkX+LmIsxZwz2JSv3LDRU65fv
3yWhEnAJWdiHsrPf4tonAhJQHJDsDXicSJdBT5krAJLegCn+QqtT7SRvq/8VhLBB
WTgktKOJBSazpjrGMfxhxFYokJngnSIzVF+Wt+WHkXIOH1TlZTHnVUWCgHXxuoip
8vDO01BxuSVCZdh/mVNe+uDLYb776csZp8pizw9pc7Zjt05C9FmLQyN2wCnJ/IpG
oyZ3UtmgE8vFN12ZyOuLLO81uVlu8N1kqRUkZRPVNXcd8A2ykeVHTczAjG9xUtm+
l/i3Wo5VHYW3EbhLkWcJ3W2lcc85uxFKgHaV4IO/N34P6Vq05fgqkrdxGSz6Reyh
rj4GeYCQe2Iakkm4r6yaSMbpXFgot6DiTG9Z2d1NIFJ8eTHapnd5UhmMYSeOvgOt
c6P/U736LJP69j1RXuymvoYHb8YIa97oY4/dUW9FZJxdV7jk/kDvXet0a1FpqJan
2bZ4eN9ADtQiRG28GnHgW+uwy5uXSeocw7Afgn28UxooBmAYckEdtIoJGoAUrgMX
j4Pf1IG1ptMkXk7q4kt6ie0Etoi52Ne78iGA2TDX/60Sntp8XUYxzKf1X5F6i2MF
1kf0XUqYi74luyuenmutNeb+g4yGF1KMjGUF/RtJ5Kz1Wa4J060uGzE40MMLHPzp
yuZa2DICr7CwnDXB5E7tiFvCcNRzr8v740VXkBzx0MdnhQDoYi2mgkHritci9cKy
Ccpt3+z6CY1dUVcABzz9QwZx8rfE00WLjpm/WfhQ/G+N0RXWgLEeXx3KHCGdQSup
4puw3ME1MOstLa2V92BYMkEOXsXlQ9MT65OI5j3qOUn4Mow1wu1Szd0X7vG+PYtx
5gKGBG766ilXuwZSzTEH2luRvEttcHZBgydQ10XeuHNXa/+RAmjK0rj+b6e3JHvD
f1edAXFYvVu0NDjOJkMoM6rq6t8GgB6iJ1MiljNmLA42dr+Q7RVcAoT3meuV5V6A
7J+Xzdm0zPsFAhW617GjxUWdPnW17+62Dx99c3tf5ul0bCKJbPbPBZOHlEocEW4u
M7gZB3B4/UfLT0F9O+PKRuf+pkvmr468cZFhg4TyLwYMGIY9iT29egT63muT+QXD
ljJiV5B8HtJpvW9KoQfrmNqWyIHd8S89Hbz2IKORfr1I9DezKQP23GluFuG3BwwT
tThX57+p0qsC9ZTwoO2Ivn3hBA0ERVgbRJygfB7qK66yA+DVEUluSP4WifB/BVhV
aCI0NcYwwR7hHT6OrzP6meAtOQAGIyAKkvcdcjhHfaL88FTiLKZWMF2OeYNp05YG
S2H+gijPVRkSd9Wck5V/QsYjoGC4sd4DuvjcxpgAmJiqUMO9N3G8sC3/9qkUk232
BeqQ6ci55X7pgLcOOWglZtTAeSW4UwWQiSPxQqAduiwzXqhgxmvJd649zZR+/VdP
8G1g/j55AC3TUSZqpORQ5cpYs349Fbga8po9E3X4mxyfZZCttX4N9A5AdfcQ8HVj
xBaDzMyLt/+Egk2GhvS2C1NznqQNIjy6PUNkGe8fvkA3e3E9qx1/mRsD0LtnOEKg
sN8uQwuBv48bKw+LtAZHUjjMZb5cd4ctNSnE5xYhNyueed6TSsQ6K5w3pwMqFvSj
2JRyIeGN830eXD/nnw0Yq9qrSv/WAsYobpk2u5XAV2CezQVNbtpOQ2ZkANlKPKID
Ngh82RjJUKTCY+eEkmEn9e6Wv06H72sQYo7P7fYK/T/7VRyL3z0BWhgtaGf7j2+G
F6baIOytZBWlRFpEkQLCOPxvCR1clFSyp3kx+lVgTUL5lVXqPPalrRdiNR8vbPKo
b9JN5BPy8Jxec5WPGRahaWA6kyiqoZEfUFLWNOJmpWngmBm3d9dtfTwLVKUls3jw
tHqehaQsPpo9jJv8OALzxwDdiKq9AmGeCe5N7URAEcILYlvKkl4nM5EtigDvUPDO
RQg4bn1vDfP6/LE2TEsi2/LeWFiJyyIVKfzKxp+7LTkxIo4vV7wpXYXbTyMjdM/+
p3X2mWK5vGBqLguu55utpQiJ8D3Dm9BVWAPTgOB8LOcl4PrHv3PYl41nKaw2JF73
lfo1/kSWftZUH5gnFmCpXDUkSGPKHV4wxNLF3zD5lg93XGTrqZNj89bY05ckKujg
oZ9o8/b2S87ZflZRneIwAVOohzFwMlXk2wQOal6vCLZSwKnUUcYCiJDYAJVwRxCB
XPKoM3H298O3RA5YLRcxwxGLfg/FQ7EAOYFPcYFbScaQlxQPIuSxDymkhI3ihSIr
4XffOrZuX+8T1ee9/+M7wD75uY3MuvDkngA/3EP5rdRoDIwExp2uRxxFLnym/G5P
clSaAgNWq+V5+g2R5UHq1+St/xgrD5z2EvvX0yJF93HVaSEYN5wxEQOVI4VRxRO6
mPoHcthljdrz3phugC03vl1fLB5lDv+8YX/3mMRDvVuOvWnq/CgcO/eQJFpFc/oj
S1Cf0xsH0k7lg1vjPyr53fNULrdyRfndyyx57Lq9RadLBMOtTCfKeuZQBkeeiiUH
4RcUdU00q7y/Zm/LjsHIfEOXSYVMCQA/2t7hUimbuF5+sLfAVTWvOREVnzGPkWWJ
0sZ8IKJrAfSlUfgB1CDhlyGL7HCFK7GKk61NL3zKNh0TmkOK0DHoJphwpT/KEInX
ss/PY764TXR2pgzxoGZXBc740TogvDa96OA9YG/RQK4n8/bD++o7UDMS1CfNwZaW
UKyE6HYNqaedXxrVMiXc6SbDPNhZRIBsZyFxqGJpAW/PMyT7NMwYuZFJnNzsQg4C
6kKPaLffEjC1BwGbVVIjRKwi9Tb+L3K/aUqpK7icrBonEb2XgXSEYGHxqhq2AvAf
cYzoI+x3Bc6av4xcsKM9cEQpi5GTp4+f8cTAh8N9s0bKhdT1ijYiRGPcXVFBdIKh
QbWFYpAdtMZRR2w5jMKbc/sMDNFU+kC31JcRNEpNFJIx4cJvm6kYxoWzqZvBSbdE
pOPa4pbIddhJOtbh8D3WNz54PgGMDVaVy/bvBAp96ZgGoWQAWF7qXrg4IsR6H+NN
e7e3MdLllOSW1xb4+xCfy3VUsYaVQ3Ux6ppXhEQXUTO4i1vpHvpBlLRECmNE3OJa
LFy1+nu9PakTCwjj7EM0ti/9KxKSP4P/rhDs0LDyMDY2hbxj0654Hqj1g2SNsGy9
qu01zlCR8zKdIvMLh84BjRhc8ZOnuycuZrZycByoEz8RyYg6QGjjiC7334NFse0I
IuQtxzmxGDt22iJ9CLO8HHEq3Q7Y1u/RrDRE9na1nZOmb5WwNaPrKuCfoLKC1tWq
smKG7u+zlUj88FItR1tCRWuxg7bvaITzJSmL1SX5OHpBJa2SE40QSLITsMRXSgOb
JtOF8JdpDrS1lum3atQgjNYO3NjHg84m1zGVDhKlDVUsCqc0tOBVdZ+xZtBpaU99
BjL16LA/vlo0CQA/u1Rdw0FHWHYu2nNqfkdr4dTuSDsng2GUwWgoMFeudtcyAH/R
5oTlFYL6nbI+hAaVZRj5YCxzSC3hWAhlDwtfanetkpkDxxWlJy7oQbi3eTPGNdZd
nD/WYuFuJ38NIXwx4ndao2/uZuapTsySvraML3FqMTQL/SRHZb2VEey/KFo9J1rd
Fa1exN+v6BgkLcqiK5GhamJ56ZqJ+pvJrApjqYwhi3qknsgbSdQrmKc6EFW+uoMr
wNJ0tSWPbw3hb5d4Cas7tDxTJngs5FAgeMNBvsAvzt6F/jJ8uDJ3sXChdvjYwpUK
z0Pq0r+/+NDfx2kxJBpmdNdjZ7doKwGas9+K4Fz82M5vSTSn98wIAwov2KSJfAYL
gmyOyuX88D4f8Aml3vnO8BiUSj3LDJ+VDvM9xe08TIW6UCgbI0zaYbGAFGOY+Cuw
zGI0HVYb2vszRquZRS5+uS2MAC1MVmxB+NnVP5A3YRcZtKNUPilmf6Ua/nsNUpbI
0Hy9srEqRsI0Xwg0PNBlrnYaBeucI4qVCSTWE3AFZFCDt8mQjXsnGyNICW1jFM+y
xYSLHJtyL5trETAlB+n0IvSnNQf19O79NceEvQIj7iZPQutCdURX0VscMnuPMH9v
uaVkyzMShbeZnEuq5zWVHzW1C/AkFp+xi8pKmCcSAEvvqn0g0PMWZ7I3MeoSIAlw
6KEMzxOay7K9zQiz0XWATCRmIMHl3GY+ydji+Nh3+fyu0gO/biSCWrNXsRhXXFSu
hUzenIMnlzJ1lf0ICYjez9l19FMwriO4J6dyo/jBmKfnuDww62StUF8gXN1rZbeD
WLoWmHOx7ATFC3OKeeSQF4J3AhYd8jWCioOaLXv5v0X47FyUgKNJKQ22IpUhh7bk
MxKOubSlT4HB9PPPCTls43Hf/WSCo6mnOngE6sHHEPZRAPG1X2yFHrWRA+STZEsM
K+LSUwFHmkfJVMU1K/LfTF2WoWwpdHFgPtN2au/yqhd4c+0G8nboabagh+0s0iFN
QuErc7rF+lkRmm9b1uRhlvbTyLa646HKp0R9jmJJ6F3hqowPFmip1wq+4AN7cb0s
SY+gxZjG8xKgqEXZ5bWA4vhjPy5pP82OgdL/OrPIgbxQeo7F7Run4dNz5trZCPI8
HLZx+L2cw5ABtbw16rWtSczIv/0zJ8kGuLVGa4w02iiDgM4jRBV/fkuNYKQhbLRk
tSua+w63hTZi17RpgMnrKi3GahlMTdzGZHQkYJeQWWoiJCtc/i0Jj/TUxrXaR9Rk
ttOR3Z6Wr86mbM1YQPNmMn7mpsBDz258rCUoQmtt02cWzwYzRz0cKQEYm8mPMay7
XIUZF7W/dI5XZQ+FVMfM3sUBjtHwl9gta/5dkaUi4SvKSSY3CrR3zI8nnZB8qeYo
3E3/PzyDycqTr9CQ9oqSFKaB0NfFz2rjD5Eu7j43732DwjauGrYBaakwrDWhbymo
cIPuEEmYXKLSiN/xrlz44/X1AYYKxxYBLyn0wBI+YG56ExykAiIACR6xISpVD1Aw
mBa+zFU0LtM+t9rOmS7NbJtkOLqtATSCtj7urMcB8BQ8HPft8git3OaH2nGvnjtX
HlhWvyYmDLtsB+nX/fc3VadI9PFWlrIy8Y/Pw7scgbI2y0O/PaS3zSCtzGuUPw/J
/hisIe5TRgrMF7yUxA3vnaKAxDou5LIXoVx4g6B4N60yFXDeUVVClYxWdPXh7+c2
RlFfUXXUu+63PIfwsr0PD+lw99NCivmy8jLckkbZVpX3iENeuwZbG4Sjy5RH6r2N
kVEfxpvSwa2pj5j4ze0Yt9ZzCVhQSpJdpm5pCVbRKOa7OVHlqebaxvB8iEzNOXC4
/OVu9V7Lnvb8JvLXFp41qtTAhFwYgK8Tw7SjxJI/T9QaftNuuyCY++GfnaCC0tzs
FeWZrXMFPJ6byccYucY/pFSpQ3SSWMG7YBrqtOF2a7YoM8LZMpUf5HRYVr+RVkp9
3gQ0QDWKz8SMGrcovuOb/THsl2x4SKQ1Sk3HDrM+UywH3FQIQX+Gij6UP05o/GOF
/CA771iM3svw4ELmPGJPyNvavETMGjeLLnVnKwXtQ9jEx+s5gwmu/6cUxeigY84I
cBqlGCsN20VmBG6TjqTnw31kXFCFBFAGSe+UYrgYSRGW0RGwgnM8ACW4t+EHD2vt
P5mQKig4G0ejNFeWJ7Ddg4dxDdH7uxKMbzjXumbcRTh5DDzoAFbnXW6wiw3SnsW3
7Hb4tYzUt6s/JNf96LWlKcHNHes9+e1RdAlH7P3HffoCwjhGqozTNT+Ji6oDC9Q9
UATgY7U423mFBc6bCg9NQsZ/hxCPy2gd8TWdMyxRKvbNk2Go3hZOvLErh2u/flzH
G8oNaiRA9wDvTI5juqd/uMRBsI+YqomS38mkYpxwGoLj9jF4pu0Dpbc6RUxe9Lv+
yOkP5y5L4N3pWo76djLEw+gpceZi4+WbnyL1VqLU1bdAlwlWsY6f1ZhX6FuJvU0m
uoWYvnE1nZ6Pahk/doFKblAJT7m6TigGCjsPBy2afcT3dK+zK0/4xpqCvovKmUlP
obDwTK63ymlR++3YOXp6lUXrWja6DlsfPhbHd8D/8437Uf6VVRb2Xf+LYQQ3r1w5
I8ycxuOmqBefJWIp+40FOQ7CEKE1uJbarhd6eAIakxxm+xRHyle696Vu3b94aURg
N87J/XI/YqaOywL3CWdyawCwZQ5i51KQ7SKeyuiu/ZC/XvshQ6K0kNUgxt+zf9ff
NRwkShEkXPV4H0VVXcmttgPKWIpsRxhAYLFM3fck9r9AtcId+Vu3Q+FA7Lun4Zew
QmRoQs4tL3kd3FaytebpiUo2eM58Rb1Y6dmX5Y8tEWy66/YpV0Ft4M0VYlxz1xSL
8J2eRWAkK8ncJfcdR5M8MOqOYE0GG7EQ4wV3YwjzlyLtrTVVMGcmwSE58a2zLHdV
kEZU9EBfjhTQIzWOlPgMV6T2LZvdltBzH/YaeJzIDEZpD1S7FzbaE59YhUFhMeYd
XG7zYkymeP+GKsXakfL7K2VOc+1/CwJb9xnJ0wTuohKJ03Vxv1hwJo5YtWQ8RCFS
yFBdYs5qrVlWrZQBOmDcimw1cQYiRu18X3AH2GyyegeZTr6+Z7tWQHuFq/b4WxQL
Dz87j370voEe0dx8Iy7INMrG5GiqNaT63eWn09sG4nrPbP3BcPXbCtjrxcYvgXxH
nNmmuDc399VsTAL8ULyjKtO8nE9GRnumFLT3J/SpGEo+qW4aG9uKmEEyerHB5nCn
1+swoe0g6KHtDsSGKYOfyIRLqHHF/Jd3zTtp9hId10/kxVMPzL2FJ0qDnPjFK01w
2I4378ZYzyM3ifSSfIdIFQX7QVgm3evTGm2lsk8e/ubJNmrfKG/WV8BjdY6sB843
7+GoDcY53vGqBzO014434M8v41Zv8yAiGt0bVAnQ/vm4xcimjFBa8j3LnFDp6XDr
4uyPFqGN3g9CGPve0r8tGuYYhEBG9lT9n+6ysOdYW2qjsVxhwgEdTBxHu1PeDcAX
xUL/M1VkyTC4TFaM2Pvpx9aC9SWLmpd/SoAE2gB46p3+Gf3knDpArFjrYMnOFNyc
2iGYzxq1XYtj0tXUGodlupkN9bkidGE4TT1xYUvsNBLwZ6cCdUKXxIJn4Brk87lH
FGyxIdL9syr7dGt/LZ5ozkYyyxPcwIJObz4/DmnUNynUQtIxrau9v2TgxFNiFV0p
GIVgmI/LoFXtcCiiAkz+sNycqH8HqwTCt1tdWpocETNgIcfigEdQ3WKawXDASM9s
B+xA3nHOIpaRg4IYFRF4lPRjv4xT+FHbnzw8xy1qUXjW3P2iyeKAPI+fqgOYhOVS
J5vW84B5pKiMiYNdvIBkLpKNgnuMwmXfX1I5jrDSl7nnWzBi++FCvJJwusOej4ev
Si4viDu+57jkaxfX2Nmc2augwR0WU62xh/a3T7qJ1fT4nE8Y3QQ8n7b8uDYnYgKd
uTPYguvBBuMDBWhpXHE4tRxSpLzfL/afR3SHPgbyuunziQfJD8y16Go6KWjdmuKq
to7MdEYTtEk8MyR3NKPJfWUsV54O0gvdU8d9Q7thzVmEDVVnZMQK89uNesej3AyS
WwPgO3AVc5o4icshkIxDTbcZSWXqf6inV+WBTnWPZ70J5TtGU6CYYsTSVjXv9qGx
E3K9HlL/uTdamDnCp5jseOiemEbNBtHhNNc3/AvnaMCnyxGa3Fdn0MkCHglx2eLh
oDxh5iS69j/J5HK0spwoyFaMx4BR9HRWiOPMT0R1zS9mTl4kS4WX1ExDCjhnMpsb
rlJVD0plIOAsJoJcZ5yMnEmUIcbl+Q5poF+lvdA5FajsRBBLQkWCtT3gsMSzEk4A
NbSVSz/YXXepvAX5tbSQLnFofR6Tgc/Kjp1mpPXio7BGVbi3f9ov1+0mWY2eGfn6
7UHdvQSTHrdJzWvMjGQIp0oFeykxMDrMPPjNts4Xkhxu2tNAwXAMiP47TY74M/ej
oGTQa0w3Th16wAdfXCSYB/mchCQ3K/puRVgXVWJYptIdOWx57TyPuzIJlpudmqo5
gvGXt7s/+FhjGAWc5/Dgd273wNysVJyXtLFO8zrr2JCakBmxyLhG2AgGHqybJg/Q
G9CfZZ0tC+QIy+cMW7lbgkeUZAFE/T0FzTwlYlqoBg7bW6ITPF/7rpuYphxVBftb
lZaE8jhfYSt2wNALTga8xVXsvWPajlKIVcXNBM1mKaFMCIoKUw2V6WoT7y+NOpbB
TvKrTAwUlBrMAyErpJdlkcm+zB7uQ6io1k+XIcXEROnh4IquwosflZd+F+Szm5MY
abL2vAHcIq2h1Rz+aXBt4hdpzpKXUa1AUum/o0RwNBE3v3PssQwI4ecTIdxVYWmn
BqFQBk9gpzq5aXH8dtLyAox3phtFNJeZc9jj7jOZCaFDOqeAzPby0amzPxllXurc
ixYbXWaHzObO1FH+CBIAXRBN25GNS7UpFsQ2wtYcVrT5YH1RsUcPGLCsuKvYwHiE
cQMMlZ00YKXsjZ/C7L1+2rPD37v8H0jThfpgdu56bQqUwRh8t6XjO0kiIFRjCMan
9xyXHOiLhCOTDKoHPpBozgIJLqe5Er9nbqFKaVTjR73QlbKRzX1RjGGZzurPDgsO
8rLtnI/qpjPRqlcJBJKr9LXBUNFxfK1e2/HC897ed+RVFVz5VSmwaGICf5ZZTrHc
eVYMHR0eMGqsGQd3KUFaSZzn8yAW1aOiR6j8qvuklWMMRuQ6eTwC9gt+m4DVXJFL
TMFHGkFQgqBDE0TsvpPMRlhOARULM/+3X/6801Hn6LM4RmnMPB08cCRxvEXntXY7
0ESeB+fkWL73+50S5N8OACKtGoBqCoWppvg24N4BJl2jJRORVvuDw0dTg0bz2/m8
lhzGzclB32RwkLYAnVNViwtJkMlXOZWjt91lAGu8tiJ7nHGbt4oFxssjAzVraEv7
H0KP7gJg+dpOKUJq4+iMHGdlT0JYZyQq7nzrYEHlS8eX7nVu9b8DoCCteabAeJH9
VHo8G/UjiOU4xaATA0+VGQvWfM8NjB1jahkPGwhByPd6XMkRRgfWEFB97bBz8ehv
iZutQFg2U0nQI+Vr8+WSEaKji29uiFXxXl9QNLZH4xBiaoBWu9B1UyHpaUeubG7w
LfP2lumhUPZZHnnoWkRXWrhNkqm0TnlddM+6iM5HdJD76NOHDfDeBUsOq9Dhp8pE
y1ikCYlzUFjWMGle0di4tYMqzewjF1UDB0YxPfbMCI6jQlAbw2q8ULSS3OaQPKCC
OgO7wwDxoGQl41IMfKngiiy9PRazJlXtWmQlnYL3i1ntYNDZxhBT7sDWSKvv+cqi
DCCWw3iGJLg8OK7o5HNgSkgq1iEpsAh/9mVwv2sA7Ai8M5IeMn6BMBVDIj1z5zi6
qlKyKCEi1fSDC3OZzcWwVsVRLUjdy6AuNAfeSLilpakdOm1RvuckiDNa4F9YFZ9Q
asIYSr4EVLlTnRM+YcrDdnKwzomt+VsDpdwMQY8ngxl9YvOD+BsKLr27r4o7EwTP
bfM/uO4AZto88oq20AXuUtYKDHVS422CUWmAm7/WWSxec3/jsfkTCqr/7CcGTr8z
6zMJW8z1Vot5UJAks8DSyd2dmyNzwp3vRgE7EBli+jMT92HXDmq43j0bho9sc3sg
jS1ZsP2U3NzswNkPIdrfCycM4iEsqpk3IPrMYa8I3YualLPnUSgdu6Tdi076rn/J
MMWUo0hAaql390Yqesy3VLxCSrpHmsylxV+A9RNzZdnn7OmvTskukQjMQVlQzRTH
A1e70oRzEqVh+7+HiHus0n+Ychnp7xoSDFm07c6JeyeDl6ihsxNYDmsdOeGwzkgw
YFyJ3jEOBAx55i+gOmtnESMWFy5kGYUzSYIcwAx/y15VILsUo1CUVwHytxIja5bI
X1u9RSRJ0/8gcNRoYWgVWscvtmGkUhEuOHAwe1ed9dxhhjb/9ZiL1+gWrqtlsyd2
AmEc6a6AKRdpWBnwZYr465ereFgiVmyzkkGI+33K+G+IRVitwnBejE4HZBgMXT8K
uAzytv9DsH9DP+rC9GRnBVP7ZTph7YI8yg0tW+C5t4OAODk9JZUh3NwE3heGWtm+
jgyikrTD/LORVanBZk5WVkO9khqE0e110f5pe4SP2qFoVMOHmLW/8zHWgikSa1HB
VlRXTfyXFdZPr7qi6RX/0mYMbvOqEuetAp/5VFgS4IFHQwKnSqv/6HVrZsMy8+Sq
PVKLb8kf9QP7eh6jwqMYnuT8L4ncNa1Z6ATLUaag2PzKbKjJ90IXrtvCVVN9XUJE
41kYzTUePAHfmZX2BGyyhuWLP0OLga+oisTJDGoNJmJ5QxmLgKfAgikt6Vi9uEzL
4kw3C34LcossNGvSCt/hIU4P4w6q3nXHBgjfLKJrtF1D9NCb+uJJv0jcu92aV5/G
AKwPfdNGyCJtcICWsagOCBMNNiCApW+rsxcwuV0AG9lOrzMNhuFTO+G0S3lBSFI8
J1P35Xfp5oxfbfQ0IdhyUgpuQa/M1AQXDPhxnLTX6WKJEGTKOssW6nJZVLmHBEJN
uWkOjllQf3F7Y16B/gNmRQxP/5PpUtDThSYACWNsBFTCT3fsxxQWl3hPdEWN4Jf+
GlX+xC7+VU9V+cC9yNUpIww8CwY72trqfi+cVAh1hmAVA7hB/o+CGiJa9QJBs/yV
Ld9g2IAEpnpu72Hm7SV33E/XtOahiEbKtAbUZJ2rkcuZz8z9hZdJB49qwSYKlIeJ
/Tf0r22oAON0K4h74Iw+u+HsMGq4SovsnQYDiJdoICQpLX1LAF8DM80ZTNJ+tNHu
wJn2Fq6sqoXDOI7HkxhVGCrYPD+H4Sl8yyQPL6eYYkK2QExKiX6JZ8aSaOMTfooN
K8eBdA3FIgglQFAps+gQm4SwFfC/+h4MUbECy+a9ZY7PPiZwF+cDmgmdLqpRFTQ8
WxBTXkv1l1FzJLyVje9jU99BxPCHY2yERfum5leO34yUzS6MI7iq8awOoRU0vSB/
pD0tGbsUjG3X+V0b9tNXRy0xxq0dsQiQ9Psrr7D8zpIDik47APSUjFM/N1IZHicS
gs/7dnNGqtLlz/stiFWtES0NMpToZdklUycGsFObIQB3I8XMm1+cbRZHx0hhvKn7
LZbZsJ7gNEUkaq+VgjYYW49gATDuVpk52JHB791bkpaa5u8TsP1KlID+gM8FdTqJ
D2I/U2l32/iqmwmZ0oFknJcOv9Qy7ceQRae2x93QDg3gQFkfVkL9UspEIXNReqcW
ue7Ih6IR2pas3tlgyAt5Z2zjrBzRKrAN/13dGXPoFH0+/87QxAFQmrdnLteXYx9B
zTxfg/lSCwBZ9p8/Jt/0qzY0eTjl056EEu2eeqUE14JSE+UNoz8ma6af4ZZN6e8d
3g8Hve0qaTdhU/irxAnn8JCqbSa47w4e5vTvj5bCZKOjJPdWzFfcLn70iaH03Oxa
Db1HvgTismpPavV80qgM2RGRC/8s8uTguNfmDchHlgg1A/dWd8LpaRqugde84ZZB
+bx3sJqTJM99WSvqIrzW2xUVwq5A+JyoMz0k5cucFWhDzOvUAXHfzDbmRqexFP2r
+kwVG37sGnj8Pd4gT6m0NojgylLY5OL1h8C2L5RzIvQHfwtYqa+Fe9Aru4lnNOUL
jbRmeXDmjmrFCOyw/6arF7TLiQw9cCkQe3kw76WIh092YkSCJ3HMWTjXl0DGYaFK
mBDx/s9Ej+ZQEKm28uUooijdZseZvN9AzW5MIcvadDd1AMzvm3ESV9CfwHGwOcHd
IemHjfdniS1PaumVuWMEdezwAZ28ElknxHIaYex6w9uw3hPQsbEA5sKMtB9+yiEf
WEIJPc+O481oYfXMW5+g4e0xXHZPPUVbJZTljbi2+8KuUGqBf6eUuCeyI17aKIcQ
MUseXMNoCf9dzur33ELzsAFt1wBpQEkn6iiOl6iVic5vMfjucIYvZ4VS2rI7Ft33
kWFWW2NUmlUQv95NOM3WO+K60pjCkytDloebwHYXs4htY3AOnGAjm0K3z/puXUkm
GFHstdL31ZL84XUpk8EaiWb8YrMbvtBYNg17noVHEpIFlvuf/JbUj4fqDQ30R1/G
0Zfvh+XsJeAjFzg7kGi+/cigIcTttGsNZ29qbIZ2GJBAtCsZf9Oi6N7dV4jRp+d9
97IRUPrBXDdBvDcgZn9FH9SWK0BqMBC25QVPAtvjQSwG0YbYF9D/R/jw2COLyXM9
wqdhloX46iE5mec2gRghonoDyEA4zgulaL5kuFgCJZQ/xVVfK9PrZ/KwbTBwa3HQ
TOJF/pSLOArXc4c1MZIkwIoyB87tgRM6qzM2jsCJIZWPX7/aQWIivwjEKteAnAXR
aDi7SpfSk54G4GLutycPTPd9ni5Qu8446erCP/ABkDkNcoqhvw8YDlKjguW8SIVm
P/rN78dFfOiaqKpOexer8/IFIL5jYukWfXQ9QI/Vl/KX0Qaqjrs5ImzUiW9wxaIp
6UCAGlbC+D74AdYlnSWhQjxcQbZX1uBteOXpbBU5Dskg/0+7u0bX0Lr1+4TxM/xB
xAiWWL7lcY+9LQGdQf+YUMLhuc8HwfcMh6RtXLwv174iqUeSLn9UVz+DsoNohxwB
wT3gi7/ccBwhumt7immhjbJ/oOzxR5JfmOmzJReqOx1mf39DDNYD2JnaznlOPjL7
vSvJAbJ/cCAqhjyUqaRS0uQXn6kHQKXRS7ABcFBF56n/EcGem97hOCjjaGX6hV+T
B/HsffkpAiZ1DEZWCGYmd/Fn1B+/j5jKU5GIV+Vvfo6ih7imQqwLwx8ZVLO6RZ/z
DwFFFSZMpO+hiK+PK41xKm9PCJ4azt1gHDtJ/J11qERktz9ZUNmL7ihEG3fczSNI
Ba9vsYOMgXlcclxgeJXrK/9eITlW14reofPTzKmt8w5rUgKxKsyXWb7+1C7kEY9J
yUHW6c6crIGVxSg3QAE9Qi2eD3j7OuUdFJLnmZ78Xwg0uqYW/yyh7mXlz4OaazOQ
1Vh/Dl9wQfxsynSwuKVxRMcNJnzK9Aj6nftftpoAkK0Ngp5noBIysQYWLPhwAmuP
pdFAva8jVZEjpwDaXevKnd3jsBXxCXPzX44LOdRhkPL5E4k9p9ku1pWyO0JBoaIv
yNBMe/FJJgH3Wqou4K1GI7RH0J0K/WM/MKmlj0B90LnPfJU6EUJTVbfIcaA6ynM0
gspYaljqyxaW4Z5gxLd+2EG+wRIYVGP2hoLMusRbqXjG4lHRxwIO3wyH0TIV+E+O
mjsYWZ5Q5zTlRVHxXTZ715odgZzqHHe9PdPEI8tUi/sGEHJFrC+2yNyj8bOXFjGf
mDnByuda1+LoiUmvRf7yCj8DBbmp8uVqulAAuynSK8eYrH28mSblFbg3y5rA2kri
5/eE8mkDjxAc420bicKvwNxrSw7FQTGDjbXm6PgNeW3T1ZYN7+0ifAGpkrfOTxoQ
+1N4btMKF5DICCXggOAdjyrFOXB76bl451jTuaXkDRd5gam0Pa0rsxqV1SbSl7Fs
DgXRye2PIL//gYqYRn5rHFYRyeXfWvp2BgzMaSeuj0zc6frQsnhImImTdv76wza7
lt3BcRggI62jjFYALNL1mIWf/9iX+Groo1SJVR5XRtOaGSevpSq5ENCyeS0lddAc
Aqcu6UqipPS2imrSe05QZHfwNDRyzpoD/wkpp3q8XJ22X7E6/AP6MEvnIA/4vxjv
qp3pW10ivuRABVRuI1jE3z69zcyDvr46CHL7hz7iXOaWolWq0k2DPAD39Pluh8wO
5uzAjt/L5OTdcHv5lVft9m5Gqc98LTx79GXZ/ENpTsd0SUsK1yCPhLt/5IeyHSeX
EGPYL7z5r/Et/9IX6YaVh2257MV+Qq00xTG76jNwDiKMsprX/0qSwfnWA9gvNT0f
I0+u2HVrqDPfRFW0FgE9QqX6fhFht237WlBgFzw/RGDY+P53ALCUfxhZlRwffTSb
GLMCpPQWyPonf3SkXm6HBgvr4Bga/mjvoVxIzAwoFnpSE6eacQ6D2klz/KC9oRhR
a7QQmZNObJLC264ohMr+1BqARLeofJf7EeWOIr/XHLG47i4qUm2WseEBqvjMYn3H
wlXvy7RZaWCh5ZMxl7DiMChXKm6zSrY4kznepHnKRwEirf6wg5bPYW4bp9LXL1ia
sylvJ2t4F/0g5doKnUNqqxzKJlyC6sHelvIkXK/8QYqi0y6ocAA9wRO9WLdVDEW5
fTD0zX2/dtnGmLGit9istYgEURDnGwZB8Q30cPjWn/SmtgbHUdpPpgqI6iZQvoph
zL2xpqQqrz7FN36e98gQA5DNfFSYSvoqNq6YbJq/8zRSejQQAfUtKSmSWeP3FcKI
2OHZfB4c6YWBQdFeHeeseTkCzTUT8uBsy84cKPLFOf13zUB8cTvlJGi4P24mJULM
UdvWJ7P04uRvF2EIxfze+luiZg7u1vcC1cKLFW2cZXjZ02IsgFByYSisMkjEQ6PC
cnMX0Z0T4R9hat4c46JFciI7/Z0b6f0x/h4dpHeX6s2Lh/ApM2qydshvcUi8Ytrz
0CVXdyNo6al2qEymao6mA+mb8wT/p/HI92WUEI+y3solaKojK6U0HnFfzs4kos7e
oaAzsKAFccOeiGa0LhJWHuqTFqK3Evt6Qxdn5S/CPcqDAJfQTHjRPIzIxCQwMIcu
bE93DDMorW14hqFVb9dSRX+aovhOcnHdG5b0x8MeqaMxBUk6JjEvoVeoe5c9Vr0l
7SEyC+whs4YxF9jvOvDWtHSf1OnRirpNpjmXlAGLdL1gczIrFseNH+cG8aeeSSMi
t6xOZakZbml4lFWMsrHc7BkWlAb4aPQsmgcdywUftP6g0qnlMRrPKV5Z+00q078Y
vMoD70Kb3meMrKduqQyT5fvF5jH0SSn0dyYpLk/EeP/Y+IrOFwFYvI3SDt09jeoi
bzQV6T4shVEP8Et0y7p9PUUvFeH0kA/FZKbYR+MdpkeBxDS1xHSlnJGNqXCXQ+da
3o+Z9umCEaCTXSyQb4gW7ElSeZlxXXLRc/uW9SLmHR3d1Y7NaUhhAXUBSJ8D825u
vUCdnPJiA2xkpr9p/jOXYQgvD1cyFt+mhdPa1y/Fdwcf0Vlx7jq68pSiO0UwjtTA
Di2PIh2EdfXxaed7xDaYYSSCDxkugBiAJGWqg5abjEVp1EO80wxY62mXKcdZYHEe
OgzvxYXMmkpwhMpqQ0p8uOQ2g53ePGuB/kM7ukrvouNJfxdWrtsFmvVSS51/BkA1
fbPF4dYnJ/P/fgiLfXWQCpHsQFRwStx4Irtfx7nL5KE2IcMASeOULnpYlZI6AiYm
Eezr11Kt0jF+YP1MIjKWLTtzvrQwNFvAJJM9t5GlPCSZDd+Xxk/b1sqtcHf8khEA
fcOmyRfG5W4W2HhLpCf8cvPCbtU5vQ+WVDkU7YZOIkq6zmrRFpZ7leG0aEFYYkSp
0GKIrIwReoUi0zpfX6lcqETJ5CEq0qIXIWEmYbUHU7dXVpwiCwMhGI7IrY0hjX5c
47RuToEc4I6hY3KiLancod7TH3YQVDsBsIRtiDtvsMp1oIN++MnIQT36Kh0N5UJB
GW9ytCKJXSkckTgTG9MPaFd53ZRG0OCgKOzR7caFR8Tc+IhDh4IcNQWuNIgowgjq
8Ty996UKnkNipfrsxiOS1rAFc9rgxwO697Y+bkS05L12PnkJwfJjUvBCxE8ov84s
5b0exO4wERfJSQ40YEFl+BNIsOP8xKyjgpjkC1glYl4GTchdACJNvgl4Rxvc8pAq
6pyODkQIc5B3cxPxCbG2mENRQY+3fI6hS11YQRWMzfxZ9TDMPd/rx/cTNZ/fR1qf
vR0zotrTapcWr2zQQY2QzEgx6z3xMbkgSl7CAT+2+TgCsbIoXmvCsqHkAuqMXRer
KSPN2A5WFC432OH5bTwWxhkWWrmXI1PH4UQEvkr7B/gNWu1JL9wJfs8dyNTSptpk
gvXjbvctYqmGUB2tBm+rD05Z6A0Q1BAgE55uXnUX9hzprWLfSMcjXP5kk9k5L3zA
39vF3UUVgea6XKnxUGSJJ7DSckbFqqvTeyHgtEXzSvN8HYwgMfolDCBwZgtUXXAy
GgBVJdbsOU4l0NAKEKtp6qPwJ/2/AEAChpHkOYP64Lss0DKv6im1V+OPG7zjGH2+
EbFjbRJK3TIoOcHLPHzmcd6xKPMz6MNP5G75ISU+AEEs9zk1vCqhpHtxOy1HXDfu
sMA+37c4Q7+RZ2Ldpm/KrZcKCyYJWZ/Ebm3iNDK0wH71SihUo+Fhu6zJXErH4O8L
uoD7/lPzlgaBldHHdK6kR+XowXr/+zdhWeMvXmWsA1+IWKPAyspV0HiTNWhsGWbe
5mFtBd9aTMK5tnsVPuvZqZfFlUYnT4UTTasZlbgK6uNV+kWwHNQzWxapZ6/OxqeF
VBGeE7pYcYHSC4GR+HI3HKxFLdk0kW9gQyLySB5FcXkWjVA9kuIYBW7la2uneta+
qeiRDSPTnFOZgkznBYCHCD7qkiWngANEcZcuPhj8xX59v8FVS5a/DWj8kNtBkZj3
bH4RinDZelvbA1G152kdM6OHWU0i+8o3U+I8Mu/sGjC7dfLmPrferG+bGUnCPQZK
en/EezIXf3FEjZtnuSqBxG3JM76H8ZDLfiFRLiQOJ2hT8gRUxeunM/9zw3E+O0El
G4LWEpWMsamjSC9XrGhPF0tXfj/xYyBR+hjixIORhZcN7qohPwtIhYHkzqsKqVTH
J9KiBCs6gXKvRcIrXviffq9fDBPvd9jJUeExxi3aYriZS92Im9hVw18hLVMKUhQ2
7qbn6wBM20hcFPRKFtY6twBxGU/KDNjFEt3Rn7zZp/N6v4gOy6n5FCmMlrHkwnqV
ufvKOl4G4GwPsGzLzfbcIi0keVJf8yQnj8Moj3nhCQw83YpGdeJujm6eieYg/IQv
wDp8rMfaTpaAXki1oC3vu0d2JCeD32Yqof8cSvKrlNxVgHNQrLunqQUwKoL5SJHm
Yid3/tqoePm7s23CyNPek+Oj27nXZcFuBECnjODNfenglgw2G2sMUUnwtx8cEh4Z
C+H6vZ9/G+rstZuP5TnHndIf4o+YLNYJnn279sy2aqQ58YrIQtrznYCKaywygF/l
h8QKJMvLCvG4ddWhB3qI7PLTyKCgZjixSOAtiCEd1O+rACG5n5YVYwQRHzmhcdQo
9l+GSSc1do3sEvfuaSIYPjf1OuND+K98gO3Y4PxvUzkQmuFF3FEYhhR1ce4YUb+i
apNyrN2+J2FJPeHUrGV+jdHTUAH5lGK2zPBO7MVipJm1Z9BlLZW0w7hIPGy3KpuC
wA7IVNHA5C8ZON0aHPj4en+cpYAhsrL0mqCkX9T9Myhd+oFE+kVSCVDY/sAzqi4S
y2/UQNPW/os43LwvoXfvEZADXc1M8kvIebjiJn/MKxCL4YmTxE+9YndU7ueE18qH
YSgqgh1W8lDU6IFT077uQO19tfBEBoqfwIVD8t2kSysQBiPfjl4kD8FpTtQj+erc
u/yJZj5nPa0QjR/J3cZ5YNy3GYSVyuckvuRxrsqKvJ3bN7+xPbUdXSIfJ4WMSivs
tjYGcSvdXzjK4jFgs5bBAd8VqmDrYkTtIBX0iespqepwPCjH0d0xL5+65FOcZZAa
kKxy8+RO5G8Fs2op0j1ce2mRlmWu0b6VT1374vPBZs2sKpyGcq6W90Q6TQqunSmm
jMRNX96d8HP1sVzjiBybZGxw68yA2I9fDaWhOqkUSsDIHVgflz7V/imwbLd9GyZ3
GSBkbATpki6AVX41fqeOCETGPvN32MmjKWOVcXvPL8p3/+gaRmG2POAXUDnQV6qh
bGOUXdrsSQ6lQdOVflYa5bpPS9cnXI+YhuCEzddL/2IblomTfnOlSWVYzBIq4m+G
66LVgK0hqV+oxSr7BVZJRu5FzzuvzW1ZWuI2hwNTR+uEtijdgEt6+lLVRoogLliq
KiNBu0A864MyTbkVR/7hq0HCXpe5NHmF9yx7ONs2/Huxd9OpM7ieUV6BIgMRJJu4
kCNaOUD5ikSFJU7jRfSfqbwm+ZPJbMDvgHbywWGtwj8FsStXza7VKUtwL5DBXmgP
7MtiztQERLV4t/mmmCmxd1vcy0Wnj1wdoIdwxITt11gQrrUAsrV5KY7LPPH091n2
WluzscH82nXT+E5x+JnRqvRAax7WjQFKLALRtmeDEEdnglSSvIxcA08YsuXIu3k/
ktCO1efIJ5L1kFCipGPIXXel7ZYotyGZjB3piLWfE0hOUQsjZshsmMkN6pVNFfZc
zGgKnPvJSJYSrwZkODqRu7yoKI8bz10VPYqcv1KN+W/gbW18KUCJ0TOGeyarBosc
Rjzaf8RBVZcEeD7O4RgpZsLbdRqY4lvpYmEYT1FIb5+n4PgxJ4FRGR/WB93E9C8k
Twvw+qEeEcwAYDk20KgFdckKaXd10kc5VLSFRoogutQhNwZkLEOwfvw1Cd5MRwHW
3aCNc9L7hBa+6C0NdgMlXLrDUUhbabNP7+U0N6mOHb8VU4i2qfJGlaSMtv20y01X
b/00CrV81ZEmMCSwFk3IY2vv70L2BlXTBLPt9eiz754/h4LnT36a/7TEZs8R3zpE
JR4tatUdODhyg+hB1OBI8WKhnR228Pp4/IX6gxBFGmHfFhK+1z2OPYkC+jYBOgg7
f9prhRaIDQfH5Y19dZm1kelASAScKs3I0Sd2ZAJwTld3/ah+vzQ1XCREloMX2F9p
dKKxnf3frHkAyAVENs6JJMGC9s9x1jY68pwXt5VTBQFJAawwCANjwwqAdkoIWsRK
vn9QYVBFhhBKSO2npvZ3eRFQ5AF7XnisvSHR21NYCOZcmVbhbzlfQcArZkcVM+6V
fwDlKINVxY4bz4SbkNQISI6KqX3p1m1eXo/VwAiZVusHIRM8G8MDDBfk5W2JjVYv
ZY3Z5pBVAYc8hqBGSy11zjnHi7sy5ZGADxngyJo7QYxf9v+YN4Jnz7w5uujRJpmJ
d/qGQBTvPbLsaU7eN0pgD+ac/IeIxnEx7Ahyb1W8/XCR2Az/Nf1kARZ7LD/B0q4t
v0OQVoItDjSIiINeouE7ic6klOenXmMt3AV4o1Xovgsvu3RGKXg8Y+dsSwV8vbik
5Wk14F6JH+LhsoteSoBYcXVM2HDv6ZOzCKDfKTv9ZyVkUVcIXAj1W2NyI1T5oBY4
cwIHzh6aoWreqgGGJ/W+1DuL1bqPr8ZltcB2X/3UpdTlJX+xjSlAC/K/+kx8LHXb
y5PitjxHFBJuoTg5Rn/znyxhqsN+YnqqtscILg3d+Gz63WynjkDJBQUhoZnNXoNr
AE1DygJB3RfYjVuAZ/tJJED1uFBB1/bqVWkd3NxEmsBbVu6gjC8Qn+sWOWaNWuvp
M5+AO5pM4HFWKmxCiLvY8Mg9rs2FWrYp+l5KXPQdm3ZZOdj5IYhxpYR3GmJls7UU
9KlhkBEcJyvfdwJ/s/cYpQ5d8u7ggEFQ8exa4zMpPsoGirLNP0Zus+eCT88PpNDr
8hCc2MvJgy29BOF5wsTUruMLHIi9TN7ccJvrkX8cMv/cg/vi6hPetzRvErOINAZc
JkQ0pIXCzv2S9JkPY9mrW66ZW8kAFnMXPDyJk3DYfL1BuqPdIyFSAGDmdtbDJD5G
UQ5dsu6R2HDkrny5lVXgrLAL0lR0aG5FQfkcLybLWGFucDM5VF6uY2iiJW1sO8nF
c6At3BQKLBVbWGVWOAPGYdcqx0qHXXij/83gDB/oYKhXkasaHc1Lr4qJKtMq7I5j
luvNdjHGDSIPXcXso361XYEK5jVJNLQ4vv82SlIKLY4QTF+dy/fCqxTxKtm6tyMw
Bln/8sg2jn0KndH7RS6dP0SEk26Ac7C/aN/crRhCyUrc2VqPuBu6H6Id7EM/LyE4
l/HGYX+V53Lauq+XsN6SLohuSNy2f8TMJYPWv50UK/Isqpja9bDtCkgwHpDzYOwA
A+Z/qLRKotoufW6wq0jQOTcwbxwQoML3aLQYmpwpaVwaAHYhuDvuuJ5ek7VXlh82
DsEOi3rY+x2OYF8nuYISwttvIbT365vNrX3YHFUXLj90mPSeUlLl/XSBgaCC0RHV
O3KVwmHNlDjeHSDxT8ZN82T6BgEKz9/FMx6GAjowUWE9shoxM2DOUK5VCMpny73s
bz1zYqp8UwJ80ym7vC+u22rD2jZxFge3F6cE7QCoQr7HKHf5Ar95FS/CdgC1Jg6j
OEzNOQ4t4xpc0BvjHU6ZFu0Qkjt1GfrNy5qGFTYgPfXN7d28LH4u4qmfP2sBBGTK
mGKnNVZkvUZfGALZCWHxfHGBBer/91mMeoJxzirub8QYvMQzC/OAEjWn6SAvgjOl
Bf135+uMEc5hG1NYthMUU1B9e6KAHHgwhYvXqofikGnUBI2hj71DfUx4r2ePwg3h
HxxMbpBgvqkd9L6vNHJXYDwnxUfLjzFTWCjqa/uccZXmmnu0okVCKhQB3512JrFZ
K9uqjOluk04TJMQxvhLSi/Ln5+EY19Ke9F8jAA+7iDIT17pWj5IDbs0oY2l4Pa0J
BQLH7UDu9y5S9YHOovHN+KsQOajriDj5uvY2Fa5sDeH+T2BN+ZU14HDJcwxJTmEh
FlVURZ2hHi5PTxGVaU7ETLdYFlWu83wuY5mo1OPkT7RgTI4+XcqHnorDsHJB7SI6
dxx5qG70o7+3pDK7XWARRTkNcsaY83hX11FOwgFtAkTi792xgh3OGPB4lOMS7Rd+
BS65hemJgOJciBV3ZSYEg575E/aLGm9txFa5vCQu2iNkHrEFdyC63DXpbU8JqFWE
OwyDGMLi8By5wP7FhzWiHx3BOHFgLRp+F17/pUaWw+Y7zf1tPrAH3pJDN1zFfiBq
p4EICFJTYA//l3dpiuIgsk0sv56lM2OxbaDZGBGs6DJArkJ6UipomMhI7htanndS
p2e3vtU84isC2+ZdgnZ/Gdk7QfZlbb8J6KLYmRgWtoJVmRxwDTEeKRy7PMLn5COH
grxPpn78fyB1S+6hSIxxeBX4IVH9n8rql/YyejelCZdoyraxYqYdSzUHPDBwP3rs
wrPO1o7+BExn+/inIQuJ1AoKxKQqDMwfyUmwQa1rJZqSrqJgZabx1SKfRjsDjdKQ
vqPr29S2nU7sa6HgiG1Soxuhnx8TZj/AChF62/PYj2/RJFZ3xk7QKNYQldXscFmX
XsSRv4fqx/7+rsh6JVAPO0PGVFo0Ow9rkWG3+nWy/fM46rfCWNqNzNWMSI03+WMk
4qtIA3+a7z8vYMJSU8w0Q6wzQma22C9/JNOHPdQjTWXs69Y4yQQ1V6ooVeTRb/F5
brKaBhmg6J9GuSOPaYFK4zkdp2/T9tEkXhbKXgLxj1ZwQvWc3vIX9ZflKHrfDYZt
fZKAza0XYEiocrZqnkDwGhQE8Lo1P5ijnbWhigL+yQsnOQnLoIrL4SWOfTTcKKry
1UGzj3WUzMvCnYWQ/y5FLiouakogw9oPQNJuyum2MEp07NoK2y2AL5xLqaL24OcT
PUgsf+xeq1zudKDTOP4JA+nOdrVz5L79gYgba22mHsKvMpCW0KcNTIDJbmhLjvmk
vDibQAvaU8+e9JZF6i5VAa+TOtwaj4KKPx0r9B7PzfOKEgbzfphNi93bM/svvdMu
CKd3pUE6ac2VPqPlBX5jalxBamUc+JEMyMjT6oUnevoXr/riN2Q8tJvXykYzp1a5
NrNiDuoQ9EsguXive7DwEw1iog1KqYVJzgfk1BcHezBKRP18QAtPBr4saNKKtq5W
XlZR1WAmePnZvgQW3tDj18eNXzvmxzPzNpUBP7aDxyZvaLA/tS5evN+XLLTXz3JT
IKROr03EzlR2w7hapYttC4gtpawrSphANcNPTjJ4cJSkxc2123Imbv+fqib/Y1n0
eowawq0zPodK/JJLjOVpIAaOEybQWppyDkGtTK83nRkkHR83y+P4Ro29Sxf8kqGC
12wWmrQ+JvtjBsnz7jjWeD7ZBzBgTAYGraAdu4wwmOw+KO5kUo+125GnbY2IY/ZU
L5QaUdW/5dpoUwYlsZmDNUtbbqGQOKAFeho6oH/ZiOU6MkQcKR8sqAxzJMNJCHaQ
khHYbknr1Is37WALUgQ5RgTTCKvfTDKfA3Du45v0Q7JXvERJPI6ov5cdEwYjOd+4
euCX5/F/aA2B/mi8YJnp5ZL259+PdF4QCKiXoqs7pXnKDSJhHh9DnG9WaZrUq6yV
BBjLdL6zhfV0edy+Vy64VZvL/7fiAvfj065Okl3oJlfHuSAzGye5d0NueiTn2Yty
XpQSvCI9R28gjFTCL2+u94oa9M2dn5Ge8eHKG1W4xZJD9tID6YnPdc3buLehEhHJ
csKyk1Q0nyfcir9D77ByJSQQZBamqiG9aIV3rMXZuP2+JrA2sujXFKT/UUUuaOoK
16YzugqgwLbl6Ko5ttoPxo1kyEtW4Me00DXa9/bRbl3L25BCZZk1+Y6pHCVLGxcM
EClJEd2GZ0zDB+WSmQmfaciv3n2ficRtFCLO4buLaYjZi7srEa4ZnWWV4EISE3o3
uke9LIAGWtAunqLUDE+d/C2QWE4oZbXFO+Mtqh5HWBAZXdp1Pp8iqag38i+DaGpu
0JpiwhxG7e84TrfOWiTUU4Sf+7oOCidIV0312ZiJQVaJoF4i1jCkBexqyOcZf+OI
EFXWPjR72SV9KM6F1zqLoVUTWW9auXlQL0kCC0UkP/R/T1Ysra0gRttczTev1ueL
LWQsbjUF5+qAe4ebOX91hRgAiW0lUp06gFjHHuXCaOxXqpw2W5bQR57LRixYasRR
N5wizYbAjvupTVKidalo9z8pa0HBXhuk7c0tWyr8YzjOC9pCTXx+kg+YeadwSNGr
mZts9E2VW4O9c3lVG0xqpMZzGYpPTMYp4K/bsQ0eV4wqtNFEs9wVn373V8ks6/R/
q2gFELB06IkYdAzOeg1UMrFlwbHQXrO0IP25EQi3oIrlmw6MWwwe1/OL5VXXLY8z
axU0lvwNGT7JlmFaR6Pxh8Y+MBH96rhhgPhfLGnIrS2FJDSJ8Q9/5HObpui+sou8
lC0xucU8w8a9GX2zUVKOYH27t4yKt3bWRNZz3JD139JhqtVqjS0j3TKFMjGDK6N+
Lk+pC4KXA4BdKEGl0owlJ8PWL9F25tUphCtK5TyiObbKcwUzchVnfePobxkblsIE
3gc1nNL2OeLc3BxgyJGNj2i0RTbuCVda8OPxSPqgawrhQAYO18nhSmtT/93cXNgA
+UoPtr9EAQn5YMUYPojQVakV6JQ1SXmvkZgshwSqK4wjpwli3FSBo5ZOOxwvOGEv
cIMWw4aS6kdqDdv48aG4H6Yt7lXZMskrcsJhjeFQR4m/lTtnnc9eZR3BJeKO8kw6
ArgeoSSoHsdVEoR5cJ09Vbwj6JdvsXhBE3hdv7z5Q9Y8GCm+5UaqkMQgky5C48ef
xHcOi9UXqayE821E/FzAF+nY4lGnPLlGn3ZOeG46ifDzLo1jGQPaWzG4Jtq6XY6W
IOe5tqJiE0JYm9fJ8ov1g15BQYbrznWTetSkuDs8Wc1FC71+VBxvsKWVEbEBrRLw
w2dJuaKB2s1n0vtFTTqMnhbwKQQaFtzC97zfeh3HGP5nuOoLBwTxRpv5aOHaFJog
rU3Q36MnSxAPxBOVTyDXHg7v64zim6S/+qt1p/aQ/3OhtH2cji/BkGkEFaU1fS19
yxuWd/tP0kEOWO51R2xHn+h7WYTIO6VW3O//LZu6ezL0loGy5z5m/P/W+j26erMN
IGgpgbczxZYO6U64E1fsTwMmubgYjfWOY6rVniud0RyJ9Ax11T0FPulRFFUvZaEk
b1hM3HfPKCAIkxyMjV5BGB19txZ8Ci3ecZJpmB550lF3wji/NO19Smy4fgO/2HNH
CNa/yQuA2RoBKJqCEFwMPd097p5mQ2TfO6lrBJy+2bKEGevWMRVAebb4f1sspTz6
K3bq99GQOADpLe0tO8mdNzJewOIvx1L5r0GaJXPIJne39S1yVCclYFB05Y7K5pxI
V6dJnXmO22htI6/RSLKmryZhVnN4HQL6Ms5EZi9W1+k63C0igpcQyHsPI1ACgvgF
PDMomwrSqHBHEAspu4vJnBGPUJDjIy5P1w7sbS/2krlsavwXLqBalM9VlHHnYGtt
QWVgAwfR9vRb2uVMgG+RTOHD0Fmw/6/4IZapeMxLSkgzsHNZRv2bDML+LcC2LI8a
k2nw3fT9cJqfkOqQdEET+g/M+AIanXi76YEeeFDV2poGkEptSBxRGk4fgGRH9t0d
J780qSYLYoaIC9uuMvgJBQssXH8Q+sB6IIXa8vdUeMhk52RibiPRXv6X1YtrSPv3
dA4BpER48XFQuNZsfFa/OGExl3u8xEME8zz0SfL25cX21e4e6mqv/9sUvwt1i4by
bIqz6GHuH+d3icXpIBEyi2aYknJlU50/N9bQgd5O88UdDLvKdUM3vkSoPa/rlpFV
wus/5gQ4YmDM5OJRG5DIkHJkhASt4pceW+f8jYwpOg2maMVETecBmto3LBbqzCor
fXxegXec/4bJxmiJwwXJqGu8VfCe/mAb6IItbkagz5Yz1PuLezhd9RovIya9J6pu
YKUuZSAJizBsTv0zrUzoHMJAWIJWBUczDmMmwBPxdM9CGBUkCJEZhGaIhsu85ycb
uCTG8xDVW3JWqfan9gP1z4WBX7MV+7U6kKitJ85d+eDmc2v8+QHBsSOO3YycOoVK
tykGwX4ICfLjT/SzH/CRXKGmiGnryCodWldQJGL6Colhn8IaxHdY6wwC/a0HVyJy
585rQLnwt6BOAem3WeuBiRvfeYNNwI+JjM7+NRLBvJTwWZErOck/qEYbYGUQnCg2
zMa++b6zCub72xZHRzzbvUnmKdA8uXroplxT+ILmHbGRYy/ctR0jaUqesaFkrUCG
4VQHT3oudXStehO8JOpbjOe11Z5lMBr2jSO/+gRSS5FXqNSEi8ZpwDuuHCcWoR1s
xMC6VOrr0PFjNGZICz6mIRLVSxi4Le6pYMoPiGIEH2RMtfAlP//d9OrNcqTSBhWP
lROZ+Ae/YFyoary81Lc60dFh/vDKanl7KPULpG55vwCrlpMOaQJfbT3iI5Cb9nDo
OkQXKYhVPigKjoGIfkla9KzP7kLNliul2/o0aHa9b89YdW3opjYUava+XhsfuGjb
ueNe+Yj+nVN8EfJZXPO6yhSWMIbLuLZgIGLArBnnmHNUZQ/mo3Y1SqbOWDfKnLUo
inaByvJ38DURPfNMoOMPVuWOlfB+79/1r5/TeoWI+wVw4fZBXRwHoLO+Zm1m9I1V
XZYsWhKWYbf5JFZ/Pmsnwa89axc9WbQNdUXDNR+QPuYVQgib5euX7X2iYMBMncOP
We8fJYRZrLrqLLpoQZAARdT/PuxxVDv7a6gTBD4xsP3uivB/Sx82qeuBZ/+KswuK
XhDTaBs6MNCjpqZdl3veRruWevDZX0pweNtN7tz4oo2QzLAWd9z6xm9J4Xtke6Qy
Mm0ZRVOiCJfdhDGwdXpf6ol8Kq4BM7AOzWlavp3OUK3dv2FO0jCNi26sFFWUohEB
RMBJ795T9xnG6pXAcfomTsPMXudpZ1fF6rG6dIz/ZEXuyqsDPaC0pPh0Mf6H6WB/
yChLs4zx0pY01kkGyCEEkotdpzXnBAtzhYlNlXlY/0Xo4UT8S/PbWAQx9LMd9DNS
wwddTINGat4Z4vNc23Y0/m1CvoGJcC34I9ebd5SiGLq7WqgCW1PUyVGtIG8m4RFn
8ExPCc09PJTeFxm+lYoVIOfuw70ZPnOyWrV7HJFOwKe6ZsEPL7EQSEtKVQFyVwae
zaxXeakkChYoogr/HDzpcyz5NBSl/xhOTlKEDWoYeTGZYHi43xKgvY88Rje16yjw
+mXmqyv+wM3xYdT8Fnz/DIHoNUr7g3CK0cKLK1KFNA9hGqFkS5r0tkK+fGHrnUeW
YaP/J5QV6/ZDktDzpXd0LRJJDohrA4IcYmE59IMwiBz/rP8mufRzEagbWzR043u1
O54PB5vlpjn60GIGFR0r30YTzxMBJ06KSPcJb9N5OuH+gquHE6udq5cQb1r6P4t8
F+x2VHyXL9p/8xZkOVmrHFRvdEYWkMCQ/NJzAlM804WQ2AHOXzn7fhZTqYo8rIT0
iZ+BI/yahj1Z+GnFL2z2hRbhB5iuciP7ONpy/gmdYsIy6n46aAM4FyWFiGlNrTWN
mtBPlBPylq/xhi57iEmEopkWSbq3pIXUroexymB+zfyHuDriUzL8TWtJW3cqqjst
2VjevT4qtZhq4/VQ74kZYuIa1Wt/JkF1ubCcjMc1cO4bHi68DxJo9ENDedfkjSn9
vQE5tgspkyoKW+SVnFYkuwFlD015TGgme7fF70upNZn6PbQGTmbTMKWn0jekVMGN
TEd1ehre8LJyXUKmelMU39DbjBWfArJtRw6Ns0oP5gwZbyposZdWtG1w2yoswTfh
DPgx+zwq33iQeU4OSFbQPt9dfyT/ZWmktf47dh0dKWaWdl+v8bVMh6y42SYYzMLB
idSZVAeq0plRUEmB5UBHhDKyZ0tUOY4ITMBOqzszTy2LGzCedwwhYnOv/fSAyvvA
/vkjaArEzbvqnOKlftR+gqsz6yqPz68lxrFqI5eMwLc6FOyMiixVWCY/E7C8fku9
a2c6G+brw0G0OfZUc/Uz7CeGgZDQkAiJuKwRy5B+vvs3yzIkRPAsQDTBCX0lALl8
ls+n4pgscendq8LZbLyBI6r7/XlBaOKf6VXHqhF3Llgr4MvxaTlDlMGocKjZQWGP
U7YZM2ARmyJaMyf54GazM9Gj4K2gNzzChlRkgy7oeDc62rs5eVBEKniq+u9v5YDh
Ukt6qdal6sTKxb2G9DhRCpsBFnlpZPmBcuDCaVggLXTeamCM9nbJQFQKzYgVmqgV
ncpS3S1v/x1IkW10nNvj5EGNfNrltnyjpsVPr18rZa35UKAFJ8/OpLqfsy2bn7OP
x/22K+B6sYjZOFbwkHirewMbICPBRp+pFNcM26UPSxtaymn/YE80fT25VuwRobDH
A+4A2YLLKYHTVoABgozCCYrzmUTjkFwdtJuauTUilrVM6kYSoino7SPxvvgvHzha
D98pc3+796YrA/5N0bX1uCnR5GtxBxMrG/4jtV4fspI7S/kA5rmxEFz2lt2AaPm5
rYYFzF0iioeCMT/4+Oz5h9nv+9oODRFjbr19QksaarGZ5GOOogIfDXbHmF0O48/R
asg2VSj49KPbQ5jkvTyq6dVuFyGjqhX7m2/2GVmNKFphK/wfp8xvLz8y5BPHtVXd
DtVTv3pw83cv//mX/kIWiQSrAI9icfhbnSNee7viSBU3ZeTEj1wSzKJQ7DFEwNfo
xoT6eRAU7r1AnBgF1AlcaM6sUTZz5BkB4t09OEEM0to20Llf92XN5gRHFCoasXu6
akzWhXRsyu4gDB44n1MLkDnAv4sJKwnuBKb64Szc3lsGKCvvqztvkZ0uMYfcaWU/
WmBHBSz7BC+A2tAxaJIPJG8svsM9LH8AwWze5bAxbfRqGrtfwOTOdAPhT04Ysg48
YNwUGw5ep89xrHqaUS9I4DGWaixaMU8N6vxya3wfxV2NTwhBMZbqdZihxWkalPfI
iQdfwe8/g3HAjgTBrRmgR+ciXrZDyq+LAeC++BCUAU4IaQxt5QusSa9UKqfH2SMd
AU7LnfLm6okhj+C/4whfd4TvP5PaC5ao+7YxyguYy/8rbyMRDaWhQCA9/ENK5NXU
pQXYRInvo0VcocNR2/vETA82VklHnTHveUEVUGHdyLZ2AC2svZcAt1m5nkkWo2rT
HZ8e3Fjr63yft1Q1TuGVtDMYY+wV4VigSEjvy/4DDgq1mxrnflzSfEatxNj+44Do
2ZPGXZ7+DIywP/pjsM8jBKcnuI8cE+XYs+W7GcJxUIxeOdeCE6JO0fzxpKJtplXF
m1fitmIMYGYMR0moVF0Jj8Oq9sIbXt8mgNeO9/I9apKkomCr66AiyOX6g6/O20IT
BAA63xZ8ye1ztqz4yQgp3ZpJjrXQn0N6K3XSeEGghL2+JwR67T5dgCmRDmylsMiY
kbx85hIBx6j4MxqIsjMyhk6kjlEGw1830jQps7YcI57RLVjbovMtyS/WLmq4FzRN
aGNhcqmV3Jzv+qKUaoMtYjVPhJn2ejsO+PJHzoBs2pL7f3r7saHKX8g57du8PZhu
fyL/BRlifgFTZrIMuaEm1QPwlpyNVH8cI3vBRMVAxiVP/rrMUCDsihWEM6wfwNIy
rUTmM3sm8SKK10oYvensG/IRMwVrGP1GNV7y3Q3I5V0KpVcAP3Dzon1tZQ6T48NY
c/C7sjFscOm+kJq/jpgvxMtU2vtWXl8KBK1lre/26eosMbLDZEbs1aCjRvdoZWcK
3rMk/O+jevsoa6malF1DL+kwRS7KZRsabtcfkfe7co3BPfOpCRkPBiLuINMWAb3t
yiYR1YuJIlauLzisSOrZvZkwmE02u4Flw65Qp3ndx4LkDZvbXbCwJJAEBRNI8S9P
7hvLKEVIa+QdwSZKnY243LcLehX7q9kUtPowzrQnOdXGimnGUnl5c7WsleiIzbWn
bvprEwaYeNPwzPJ8erfl3LND1swEhByFufTygjiLFqUN7xOUEcihGBHwrIGFrnHG
KpR1jH3zzkCeDI5ODxl+8RJSjwF8UpXm1tBvmUibsV06b1G/OPHPUEET6h6ePQca
Dd/imjlaAAZCyeZVbCqAtgO1IWB18/Lzv/QDWKSlnHe/XkUhpn3yMlJSPiXXpbrW
EpLzfzdqoniY+iGbK454XHepQPCu/V9sn2su5/21a9WwkBSCKGEBpCuHqnn0D8tC
1ZA1+qgYWb7WJRI1ks601zElqN1ZrGNtrNjBtZILfhEIBxRGV+MYdy7x0JIOG6td
lA0g+muYd2Sgw4TyWZiiPk6g3Ae0rddLHOWOBngQNlOpdv9AgWGRYcFou+V9wzcZ
FoYT6aXGEYgvMn2MHnNtOeCyZRMUylvHfctEODkLRGSt8saR3iOyP2xw8/MHAkrT
xShZWDmi5Bh7K7Iqf+RWH7mSb8/3S7Xg3hfqa7jm9gm8g45+RWbeQIbFhUB6kE/b
Cm6WjDS8P5nn2oYlBixLg4c1txEiaF//WKrEv/uvSp7Ehv6nSRdmwGAq4xBnjzbP
7sltYsJSZn9w5l6B2JjqXPxdAslcgS9JkToTGG7sDTsIKoOfy8jiRZbS3T3JViOS
wz12m60FPK0FBK3OXP6+xzuG7sXAGBP9lxeMLFFSAc2bxwCtahoW2Gjxyk3yQoay
b/0oO89hTrZWfqT1jzWvJU+rAqJbJzbTCYShvWAlDCrhpBi6gzY/5M12/A/VEDGf
RKlvNrG24bWZrgD8t6sipby4eC0vAEkmnpEpPBfDvItt+NkAtM82Fcy+ojzaHblZ
sbzxiuZmhqi0upWYCo+2GVL7/4kiWKGUm+BK44wmMMuCH5TxIirvVUo9onbB2vBk
QOGEESGzpLJmStEzw52/g2wHUstfSicnboFHyhUNuGf2bbrxfeA9bJPAPAX+nN11
u9HtM6JxXOe5D5CItQl6gUZeGfNfRxMzuOJiGr0SQ5rwZJwojsz+AKtOM5JU+92d
n/bHBq6GLZWcA9Hlm8CUPIUdDKIOOZbpm87VFPxB8LtHzleq3LggYlkzUp3ux2LS
XLvQm95vyyyMXUDu5xhjqPArzk0iuWfk+CiHSfUBfhxcr8lPi6WJIkSiUYLnbqJK
lTGhJlkOgTc6mSWcO6aqW0qMHJjnb1zIokEdz3oCKWg8pmgUVMr9TWU1kO/LEZHJ
yRZtsvKuYUL89udBUGHhDVjWDUCBFKC7KTBPddKBMPwOpZeVwMjqi3U/AcPLWvDG
OQ9ScnCvWDx+GniRCgw5fd4bzHHXnN712nwS5wsFc9DzI2Do50JDWJXXwE40LVDF
SkjthbwfJ4uINfbqZPdy/yJOyq2jXboEZIMJLIS0ncG5crXrm+0nfr9ENCp9FE1s
zOgpPrFESqKwcYmhX/qeDU3X3PeJ1XTT5iij4dhnR/rezEhRBCduf64xni9Xre+F
ksRpz56iawJLHavzKwp9jusZxFgkyEq6sJCHrQdfsHREXMgAawjhYgmTJtsdmDvk
q52MADpqus3U9MFo/x+Ywt0b2NeDQ//ZrrpPao+IG39mIBfCtd8dX0AsfjOK79nu
5f7L/MnnaULoQhQZBAAuPnjY1zfyzhv0lNJvIIMxXCeU7oTUAuMob8PiUl3mBjRN
AddE4l+cRVwcshqOy5qXbnmt0qUIkqaPXLwNsfgNFxtNkYlmCJqq8GlbrICtTSGB
c1fiQt4ymSGX9dibAqUYXpedRL2akPQS1IEMx+Rl1DqZzc6W41eOtbmBxXWU9m/k
4Q3opFhux4MWXlJdXaMCPyWKTjiC3MYP/RmdSOEJMDuct4qdkdHifbKY7NhG7wLb
nrcIfwbXAqgP8ej72VRyib3/5m+wH3Nndfz6Xg89j+uz2F4A+SUy+4cNlrAA/9Qe
C4rJCmmtV42E21ZsoODk0cuOo0tfOCt7rYvPbTp0NzTY5RKAiN1HxnNhZ8Twt/bS
2393VpslndTWE3Y/uDju5vxfzXEvWclbacX3wJV0cDSZkLyQx+xXXTap8kTSZq+P
tfSE4p+hG07i0DuPn7v1CvN3kabWPnGAllwQaAzfNHbVTFxzre6oMComYzmfZp7n
AW89gZsOYikGRLud9LridtwCZGhAJDOHrP37LttWoHEz/YMdQg1JZoFXvk0XQXFB
ExCcjjU0lv3gK5qRf7++TvEcK1LRxiKlMzsS5RcPV25Q27kZ73x2T1+K9L8uEms7
/iwbnHO/uH2FamNp2lthAnpfbZVtpzSFLeg6iRp0HJJUn+yGEQ9G1Di9fDDZIgP+
y2wvB5Xgtrr40K8z7HbpjjMVGV/RMQGJQ2s4j0pbyepVqNNcj8y77iRQ0ieqv3gT
Gk9iDYF5usuNtGJE0FvJFiENRjVvtS+GSfzFjV6U2TxNt9br/lSN/K/lbIbUac77
C2q/SUTg43sWpJy5j3wMFX5rVX9fZwugYJ15/znUnmCa659fhCHrquZnkyBiaHRQ
AjUyRcpT8dog5KMEglNnFK5/zf35GZmFWG45jpkCOTavGP47dVQ76AGJqPl0zTXm
9gbtf9ct8ynaKY0DQbzGzy2g2bNGCzNZvr38V4doEeETiTiLAhL3Ey9XsNR6U4Z8
z7viKwcwf3F4kkZc8aFQtDrzfeIPiAuK9Gg0plecv7D0GcPuqGAs+cp0G8wlWCLi
VfvzLnviTPmcFMD0OucatJw5XwxiQ/M77v4xQe39Iz78Iga7aAogeduN4nj4M19K
/S7ZKr6oBLhP9hJFq9U/V6XCBge+575Uvfs0AKSu7Ye+xfaTMRqa8kfZyV0zrmhA
tk+2kr/mgUh20sosQOKT+X8d39u8k7xEwBfC4cOOiE1ogaDXDFavuusw1UQw9g+V
6UsC0rtzp9Wb64Msh9GsqR4HLzEgYsnaJq74sMr7omiSkZdycaKKLLJFencdOprG
tbQJJpywzW2S1aOkbqKqHCCxH9Px6z0TZdb0GgAWXvxFxoYYAR7AnjvGj3wqB3ZV
1xjgcIwfMy/QsAGzZVwFCgWtOllj2Kg+/GXSIu5Y4Kumn4JlogeIm3NRLgRJwJAE
KK13OO74Ku7vrvvUH4D/zT/QgsnTZyuRdLOsIwjYTjwxD7RlmXnEqCCfIHtOpXZp
VV/w8Ythtbs36sqIxPPnXJPYO0maZe3l0Dxit3l18PL7uHGexcIA4DI6Xno6/3ce
OnG+vNb06q20xScOYWSVdg2tiEhkGSiy9xnsVUHeSd9SdJNuKWXu2FDzD5F/8Zt6
zGeMjuUBi9tGloCIrX1G7gZasFj18Fmou5hbT+/s45ji9mMFhxLugANJpX5Bu1bF
erDYGpUB00aoPlUsBdSgIsi5aKR/KqGGNnrS+xDrXUvJtwCsjKVVWXTFfpOjnIKN
M7JBVd5UMGy7x7MfnbFH1xZmpCO44G+CYMVnJfR/VaF+bdSRhCie7hTbPb2gL3me
Q9C7ZNpqGgwUw83WvoeHGaP6XIlktD/2T4OKwvze7gQKEF6vhZPqjQwDfblyyWGS
Wh2LSccP5NsBfB3CvogIdXFm0t4R/7aI5wzhtb2IbmfVjtP0rSHU/nDJc90kph7Y
bcrANk7tl5tewxwrcTGNqDfA74tmLsNyQTWVh6eIRkqqhmi6uZHYJCemO3VBSAhN
tYbGmIY73RoU+Tr/Cqw6iw5jC+TPEpvtCfgsXZW6NYsRMEyz7M3I5Hld0pXSkwg6
JqWTiYYBb1E6CPXKYVcmcOKqZwJpKacPq8KF9fqXdxuskNipdLfjq+EmqY3/D8B8
ADCBVkCCPPEqCwJbwlklR9z5mp7dGyzfg3CgPZvKEpC1nFxeV5HtHclNWYoKZ3tW
+so4TE6MnYVo0OVkMnu4iC/jbmRWjdngyzPmKt0+sw9lpQM1tmYE9hIXHRQS+FuE
RWPbjZN0xlltcgxHt70AzlSYkR7EtXRLv3cvK7DtkoCovMzQvFh7VIF21LLuSJzS
iPTV32v8kL55fS2YTmaWWdpNGLehWzeAS2S8RUjb+H5VwjdkKPoiXlBNbdWtiDni
c5IdfjWkJ02nuac8Hhmks80uQKg/lM7EJE9h/mIu4wZ4UDXszoDDoHJLSovNIyhd
Wz41dTSvtxEjneVyxa+WlKhNXATldiKhfZrAIFAiAH5BYtRssFUoQ1dCJh1+Ih5G
ROe1AWaaOAqOknBXh9NV8fo0ule4cemmKXU6cgSbCatA83KhOMqYvxti5ShUyF+5
IouAw1rXWBXXBPVHv2HjuoGnombKnSQt7PjynFk2tSd1V0aTS8IbsW9gxsrvesPi
rVSsd2mYkVw6AkuFv3+O0QuNFzjaJqwi1wA6amh7gZOl4Jl7rbnb2BJkT71tbG1u
fG5dXby6fOtfXnyAnrkgt3VqE/CLp9iOhJg3q+zcKxg2gzhb+htjGx8i0rdPmeYd
UGRItk2IGD2MxH7db2vmY5473YMUfhs7T0FEJcvyB3+7PWN4oxfjvK0ysRraOcp0
DrIqECAEZ6JJjm6MNSSTgZwyDMYBnWFAX7ssssC3ZJVlEG4S3uJ1c/oaByl1uatv
WWrXdO2hb9+BpeKbKUSyRmhKxm3PRQZgRna02P2IeYhvyKc8g8/v68Qc2yHXa9XZ
fsDDN05NdJ8/if1y9iHrsAfAeicjrVEJiwFR6oKR0HWy910kmcbmFLWPYOeMUT4v
8UkcOWHzGgCv42NIL6E4u7k+QFmzO9AIRwUNUCeA8zdOAlIokevypGi8VVomkseQ
Gy6jCjCVjG/3Er5EKbIGvZcNSFSCoKgR+flNgdypMDyhnKTzZ/dOaKrm90wy28+n
Mf5mMyhp8RRon+wCBmJcfPz5fPsSGXkv0AJHwubTizTj5cAlA1aGtp0u9RSgGZRK
WmShjX/C9PjOttvHPzf7h/9DyJkRBx9Se08TnLT5an9bWWJV8aidHGOwXM27fLyQ
50opuMUMk/fZKEKMOOkw+YodKx9uA99yju+Li5VCl7IsaI4BtSFD/2NdTfJYSPUG
OwaJ82jUvtNbrSStDnoPxEhY32KqS3GskQ7TkdE0/zSITVSxaxwye742T4d/dIht
COuVGHrkwj+M5Hsuxhydt+0sDklEupC2856nQsp1JfyoONmwYtUFz2Omcihww96b
tnoF7ysWE0nPGISje/QliH8Ujsz41jSVrtrXh8dEx1UWpSU3ZptRJ5HtgSOK/5EE
0om9OFFRqMWbbITi8llm26k6PIlIEuwuBdW9Ro0Mp6yuwEcUcVqD89aVOzkzUyYR
c6mP3U4FfGuHlvMWsGzHZEKlSTW1t+VNs/5iUr++Qu/9ancPCKzmu4ReIOlhWucr
dGZts8cWoxIAS+RbDj9kEnI9mIylQqgoqyc2PpboU10pZe3yGO+rRzdgR6WNDNgW
Jbk6lQU8x9oTk/bVQF8ihAouLkYhhHgF3EAXLQpKYVXD2hpzwTvyigmvUjdbX3aR
uksSBFCQ4cnQ557zh4vhaNuAwGO2VuMhRvqGabzLvWATpn+O6L75mZhv9ZQT8BB0
iN0/IzYlE4FqBQCssMxQy814+wYP883adDIHV0MtasCMTBBMLFSKVAVnGSi1JRS9
GW5tLfSUPA6G+e5nrmj7dNhRXOkcuhd2R2C7U42SYy6eDOfD5+0aUkTVFe5GSEPc
djpvC/cGgjMAP+ZqMaicQfn2/PXv9wwyGw+WH4h4cO8aC6OkIj26iCMk1CangRp2
56/pYq5tFXR6UE3pIhqhnnZIzoFBZtqGM5THSgabiuvVCJf7e4auiHmCK4/TcxxN
7aopOKWQTBD2KES4PtGz96rXb8JalKGmRNx60cWJiDU7kDPos+Xrd3rEhlOIZn+L
zX/CNXQDW13105sceoWw2NGTNgQcOZ9Z5GRtOAnG2DlKap9VJ6RJIyUsbQ2j9KGk
phTojLGqpswIDUlmApqvwxZp7ejQqMaDpNOlceX1EWxhgJ1N5lGcpxr6Qalt8lrA
Lu6ZAJtK87H5PPDiognHume1N6J6PR2ylNi2dfJPm4QtEMV3O0peIYaanOaUXUhZ
eMgSZTRjQrZ8Ilu0w8wsgKrJI9fhH2p2h16lxidVUG+7vtQhx3fnwuO4b1tOiymg
kfFVH+kRv3VddParwCwlYJaLf+jXUyNclJoPPUR0xKYyJRDnzFDIsOfrTbaHpdFs
Z6Erf2VZFObaNkjT3Rh5Tf1H7y7rKG+Dc89Fv7pdYqQ3AdLUkpnOV6bx8fVx3MVR
a6IyVs7aMlnU7Ch61HJU46qWCzfNMN79OwjHaoAV/TkoyAzzfXfQoMGdBfnA6pf4
aDGmiODhJI5mZliDZCQmFFgjrGo1V9n+chvzfO7wuFuRPqBAuklLAdPtV2C1oesL
vtGYlWPZCTuPDeErZ52SHuz5+i8p3j7Lkg6QXXE+N4u3QprISZ5NVsnn03P0A9pc
eUFo35gAim9YbjEsBmyEqA2IZ1yVFqG0u3nbHAPTAcVp+jsV/a9Ntn2WivfdkgQf
RulTskrJuZRcy/yviz1GXHbFBsPUcgUh3C6JPC5QmOIy1fwhjJLJuzco5Yf7HsQV
plDGO4UyxSokX0+f/5GEfj5RBF70ZVn1xkH7aP1rPVPEkiUX+MAFxyMEe2ur3skG
iV6Wh91jeS9ouVcQSq5QINLjXCR9fZPsDR77YiM+0SXuda85JNLs6b2qh307mVR3
lnjX9g84A707wvaEAQX5J13KgbaNMwZWA907DFtMP42a93K3m7PouBrIHFBJP7Ll
WJ/k/zLT+H51s9182U2UiAygTpVlGq+aFU9p8Yq1VO9ofvhsUg/VU9IDcyxVtCgi
tZP7RABdGr5SfZJddvlGfTxHwvwTrgEfy0mR/3eBX8+ADhe8iTC9nws3wxq9S6Ou
j5DeF2yT08+pN494S/F/KQgEk2dDkroKAy6WGQ1Xo3XDPGcJRm2V5BSkJi8hTOMk
1+91QPFnuH0b23jshsyivEsKw5aIWDMHsMDqmT9HxmCQQm3BXlvqYTbXmruDKqG9
TL5QcfwU01SI+Jr/h3CqkbyZb68deaemHtufTwB2cuyAdcGNsn1/slIMLlVDQuhm
MU3pZ3BfhmTusdX5rHeKrnQMI6I1I0batsW5QsexiSvvcc8p5P6ngz4EYWghkUDE
7MGf5D5uiDrPY1pAat0KZyMhbdAA+KUR5MOilhgHa66tFmI36TxNXsXWY6oxQB30
MIE3q/4vukO6NzUY6P/oESG7PDLb771Nm+SqTlkOwWVaXlYB5m3V80fb76O0EyRY
HiW4Dcm9UqEHlBnQBBFuapilaIFs+jbcJ53hxF1oZbWjdYfszMmwp1GFY7tiht6d
95QDNzoFsE9aX1+xj0lzUPrhv9th+ZDTVjuOE7BfQTB2vzTp2V+sGVkkAm3dk6W4
xi/W4RrTmQaPbatJaJ/mZn5NfQLRrq0a4h7L+d2ZreNqTQcPaz48+plxEuQr68A1
35R1ZVqB5yckAhWB68dsrisXMbWkhoIXCA/nDSyVFVkOC2k6oOhQ5nN0DwWGeg2L
ChV59FiEiOg+BQSgJKD+IDWpK9A0YY3Y1F6T778PBDLRNsMHQKSoy76Rq9DjGYUl
L9FaKPbEneTxLlQ3Q8ixZEEqFRavOlgEI8kJUjhx9eIQPAibYyi7kjO3pn/RNbTM
kWcKDiVxqtj3O2LWM5P6DwxORJYZG0acC1RJ5Gu35rsuNvgiMW33xrz511vgpByh
vfPijmUWqZatRskvYjnjfeDCFhgo4uoNMfvnbdA6wcWKLJnuB5GOGKidglLaFMFR
CDknoiQYSQPA5XQKcJ1lpKKbetfLdMdGVEwJ/DcH7hB0skc3RGahYuCKl7tgxyNV
Kwljl9k6OIEVK4UQ3K8wC5t3JO3ZJSya/IrRbPWQSKKt6NtsGcoG97RKZvH8MVeo
X9g+lUDV8vNPE5eqjiebbvLbZ2VyVccjwwZbG5lWt01vNffTjqnkIAEsKDNn0Zaw
nmOuzj2pH1wP43m7dKUCbWhpsat9FcvdXhggQ5BauNYHU/TgnakFNsSoItLQC133
E/S3/Rc5Q6p8R2hedUF/KtR4v9m/+KPO7wbeQoZWdkQ+pOSOK0gTjdj0FlfBpxV/
9RcvfBBJY/w27jJdjK8k9i/Y1j1NeuR5Q633n7SAu/a+KpuzLPLBkUwpiRqEodFm
OOG/UmSoYFhL/X6Jue7H0CLv6cPtkcXQf7egzhUFLWRUsdMZ/FvxWZLxDcHovM5K
SL6/KMGBGfzR6PJkCkPPwn97nqoWdvt5KCeh4lagwkDQu/8Vt4z2znIkoXpy8UIx
ryrghGB9k488bf9oV6GQjrbf1d9xywrEQbR0W3ys4GanhkWGNz2ZVPzrHnbxykXU
XZbiskePy6zQluyl6n+rL/Mf8tvfdgSCWb+4+8TZmTYFsmeNYqyzHe/KVzLceRYF
Va8h/rhEbSPsbODfSO+dVKF5WXre42t7V1VxkXqPTkxSDoHlKb00faBywQKQtQWU
MPbNStCy9ohVHQJn+dy4ldyGNmns4NWECCq3rWvdsiYwlc+403vJdCGebKAEXhp7
tHMIl3JLTCR9itHClmQAPNeMCLsBKD6VgHEeMyUH2ByfzLbKDLyHlgEdcs64/Dfp
xBgKDCN3wJHHi1XXMNtQS7WCJCJsP8Z8d3ebEX5+FcCbyTS445pggW1pV+q5mez3
f7yQFkbPXhuIJN8MvPEHJ8apcDUwx3PA7+8rNH9Ns93Zdt/7YsZWfg27BN2h+Khm
gXsAjAWxlDtcjH8+2LZYJfPocVivry3oHGdW3cOLJA/tspr70p/5M33QCNOk+lre
AV1Gvt9GU744J8b47pQswc9PZX3hjeGMeG2JcraqbwZqElq1V7LebUjaC2yUlAMA
8rqR0c8fY7EUmdz8++QB9bspuNkOcbKQzp6oAekjC8s3Z8U0nBJikFRCOFmF9SdF
lO7WfRoyGNarQjFYr8UoRCtUrfS5bSusBMThtEP3FYtxBzZlWxb9i4GRHuOw8TDV
3gwlm/nqTadxUVgmNDs8nhI9X9nW36glyE0jhTjysmUJmJYX+tOoTThhO5vuw16/
zs28DeK1JxC2Ao9QSzALQ6IQIBVtEsdfWkJG5obXqaM6wdhz5S3O73eF/VbW21Ax
kGes2Zy6oxV+ygDVz6kvQYmCZ7S845bv3Ze1KKRRD8tRW8HOubQdclQ7cTIbzdiR
FNaL0mrGetiSincaAAXsaC0monpb6a/SRBnpws089ZBRIXWzPLUD7524pL/UKUny
qZfkHinysrbom44vL1EBP/pduXjt1bkwCZiHDgsUq3z+28PA9vag0rRrTQc3FZHp
YV1qKNNO5UmUbflYVqA40iqPrOzsJr/u0jyvL8wmGjq6RAbLHH598iq053vXPdg5
14aRmWasq73Zu5fnJNi0Qn3PUbjbN+H0WicdmaDCpdm90RR7RTli2QGRxzW2Re6D
Gj9QLDjanYu6NHzqQmAtL5HCCuGWbFX/Ack6vE97LnuXxSf4Rd1r64gQ3kwd9hUK
L38xOrEo4eg0sWKC+LfTPQUy8tlLRMhaiflchlrSlW3UsSnbRKPE+QEH3UJNrKt1
xQlWpsPKVG2LogYJhw+cUHC2c9Aky2ih4xxlVYU78lX7HF156sLSZ+9IsI3AiHJc
VzgBRyc7vxyqqLEb65NUUG8DPzbij8uZDmJXxTkELZu2cvNJmQPkp80b3K1EoUht
DJaaZR1eQ5D3GrRHbwf1cdh8EfE85oQeqyiAC+2wnlP6wMuEJOVqw+MkWHbCA6fP
NAakQGR1dEAQM+ArpSNseg1tHJIVwmMyZssaYc0fJQuaERPC20CdFCAFbrRAcY89
gy6uLD/psQHZHmeKPg7DYQkcvYpFFQBPZEoi3zJ7lsuFRLs87Rb0yhctY9c8Ap4I
atcveWMTrcwNXsjsyUyMlScSQEPJS8RZ2t7sweyuiSFAIj9K/y9lgDPWhKb6mww3
XBZBZUGqB4yeoH5VHkVq+fykNneLp8UueT+7AUwS4kLuuY3RdKaJjKhVz5MQlbnq
eMV7pakG1Dj5fn6aT2JvDjZZRL9zZDo6AVgiMOIXnsJrK038J9epi7K1KVeHBxzE
AqNsMS7LABZ3GnZctrMTd8CHeOdcxt2L1hiBheA4AiYELsDyx5cnPN2fo9TSVgns
3yFgTS6nBBbwGY1Y6H0+Szbv58HiPClz4YzwsRZe68ofSHgEVmN0deR8BUFPJQp3
Vt1Nr4H0xOdI7tz4iFCyXFrqrTv9eypSzkvTwR8F2bHlmW3T9dn9QiPqN7wL9gm/
Y+ZxjbsiSVGm3VgoZv4oTeAZaia+kIQWIFjpjDtoiAgfDsaBIGjbcZcwszr5XUlD
Psr97Fonem9q/EzBGDD3lm4nz9VcxWFe50nok6tPcCtbY0iL/06rihZrbCN7uM2X
KuqmogoYIixVLZAkwuKc1Vg7Q6/EaptA4mb/aZaKY/hTYh/WwIX11iLWn32INd3g
wGavjolNLOcx5qwquc1dID/NbQ4g6uINwKPbcgV4B5T5kse2NJ6bzb9z9O0/BAOq
PldQdMsAQ1UqxTo5QhP5Dfe3MUCxnEEs+P4P+wOSRQapA7salPe4h6tVi/3bc5jH
Z6Kssx2Gro7yQy9zMh32Qf3dxa4bh7uiRYvWL9JyHNzo42wNxbDAcMgfVk0reoad
UHRslFlQpY2qQYOuM1rVWbs5A7AlTf+VgqsWJwd7iND6CwucNjVD6Xh2gzE9c3nI
pFFWuNF7VQiXYS92bpJKMgya9HiXOrpdgLNv+YoJ45bcd6jNbWyBHBzydWAvNBmv
6gWg1jfFueaZBJyFGwAEAHqf5EDdxiKsAyChRRNL8fgD3Zof8YBxFYN38d+385bw
JaFbef+fh+MGTfw0Ff3yFzVyCHUkwCzv1BAlPJRLimr4ISXtiVsJ7MYD1YTo7Xso
Fy0A1iCU8pcRTFRlcEMC6R1aXK59D/pI1Bja0mnBPZFoVtiISaRwx1LZ/Jp9P3hb
e9hM0+nnl1QPZjJMhmN8TYVClk3wZ/Cdp02DM/Lh1CFieuA/NQQTC4uDap9kMpht
bKYdh2+WqAM1aAGXvjNgnPoXc9lqadOCrgasxAchuI/NWw+sLjMpM1ou7xJ0wFPd
nTKAt35fsxyvBpiDGW7yQAT3g7oD3jX9+CEQui2olCPDqrOK3Exp4wIwS6pQr/8C
78FeVDfd2+6kkJGKNZ9RP4b9TcTmUNzunxHG9yeDH/Zv78FAA5nWazc2o1GAWMrx
bHwSpwS7+IxCKYlXPSMi4/b/94L3pcsbEEYvhapjmOV+vNbeQnnpKInLuHeMh+nA
lkIFMC25407ji0r2gxC2XzM4n6c3xWaoIFWX9oGBo60fZ/0sAz/pylmthkmfD8M+
BJpysR0O0ugRjngQUKCm9UFWztaf7xDHwzNcpndgZapFMA9KrXZqDH0TOJl+4Qyl
tWL0C8LCCZI973b6wGo76961qMLNcESfEXSzgyM/cNPfIGzsKFNKhv5Xqm8z5aAi
CMeLNK4kNDWlAwA66kvAJqDhFu801TBwyOl3eVMQD9YsQEXmmLUJ0//1LQGzMiD+
8G0+pkFCyRCvghYoHp1Kau9z5QS1bGLRAMJTMKfhDqzkRSu27/QkCGNz2uQ6+255
YV31Vn69JzIubmM4DdRa93jD2X9lmwboU8qNiaqRYp1ybKdLxFD7Pz0x2qQ+3coE
s2/wrENm4Eo0mh251Ohluvxh6vtBfFaQXwVJitKArPZXXJsob0MAqNkw3dyJHg/t
7h4L9R7Idj0XQiGQRKJ9v2na5ijP7+rbRIYkWfB5u/ndY8f4DWH0viMwn6oKTWIy
T2fyr11fYojGyDLUsytRqvE/pgVMSdz+w4pDJbfX+Mw9lz/JBNw4/afF3zGk+o7m
dsJPb5DB18DUr7brxpWeZB9YtUBhzQfwjaLT18RFx7KrI3bVAbOtIZn+nlO/lQV/
6An9MVG3ll2234rGO5l1AWtVqS0UeVtuT24Pnuy+dW/PYQCxXnBbZ1Lc6lEEOD8p
4D28RwSkVk+wqH4urPbYd5ZDRhOr8sAYkDRSxQgFrBIOjNSYMYJZSkPt1kaMBRAI
w429LLp8zT0qtdyUjurGR7RHBaAmV5JGdSYj+BYx7vXzFbYdx73/QPYrVV91eor1
s0NhjLDGJywLb1GcMNrYVviARhsDPhPlc+1/u7MXEKLeoG9WBxFrra531A5hv4L8
8MKNrFWs1FDpzmSX4txZgdasAqs4+lYMpyfKSj8sh5viAI4zzGFidvvgshZvekUK
agJEnby1B4CBtsxBt/vHqesIOmpOTfIdGBkKfhKHwhaKOZ3belvhJPRuef+7I/1F
S3YeyfelcI37ujK3wYDwMuvsiepJQCrUpZAyE3ynhK/OeAd9M9pbWOQM6IPzu7j3
VBsNwenZhmqmLSSEBRyYeiWd9Fl1TpAmVpPKrDMhsh5lN1io3WMrdUIVext3rrFv
hN7Bmg0cXFODkclZYBUVB5ZljtYz0JgxMTuTKdJr2ccRGfsc6D1VCub4CYMeCJOb
h08DILYo4mWVLttcOV8IpuEFl/CDGrHBEspMr70TdMj5uABjxm6xnlqOrIgjT12Y
TJbdT3fPnprpNcecuBNfcU375lO/KHFua58xNpcgp7Bd35C+byFSULwcxQXtWdC0
thioJsSSC0GFsVz/uwacftgjAtZVEpFKzMHzUPL3l5pp5oPAphw16xGTVkDJxkUs
0BGHeDJU38b/7i/1pJN63U6iu0YIit6XFyFmzZdDhrgoEkB/5LQ8iRfycci0M7Xq
FBkm+dGpDOwlwQTPokh/qZIEbxxd2PhQ2H13JZhsvHLxuTUZSWAZfnZXCaWq9LSm
uC2JPXz5RuGD8MtVFxJkdy/tspeYpRqx1gAlQzhx0F4gE9FhBY0SLw46mDn0x/Qo
p9quYfJCzKguj2t7dPFw4lN1Vh6BBsed7/6Y9+OIyRGVX4jzSthy/GmMX5rX7wwJ
NVMNdmfxViMGemTzSiR2EnvnfSHOOTlqlykaLB13dLnEdflOZGaeURhP7kInTmwC
Nn2h7B3x00AjijBAYYvt5+QJ4XBAdiuhlhDztb2wa5u8I1ta7SQdc+WcuU2hTtBB
WHhf3rDr63DTKDGT4bG4+46HcdcmVi0kiVvY9yBRexcNIHPKWnvKT0jf95RZi8/H
n92rtZYu8Fi7z0mB2VRsJu9Nj4uojY6zHxE46uxNbxa96FPtL8hZ2V+qaW1neTPz
BdcO77NmcMy6IKC2YVWEiG5EISuy8cLJSyj4SWM52iRzFF90AvP93CZ9kT9i8aqd
wuk5igl77/Na0Dgh6jKmfMwZWCL3ms1eq+hp88VUX9jaSvP93QKFuoCrmqVHjmZG
9p6tk/aX955WA2YczTr6TWUM0aL6GjF1lspRS8FP+2iqH/wWXhfOL2LRBjkm7lzh
/7gceiU2gOHgxitpHVj5oA1KmtCwWB9IFWUXFP3mPHxus0Q2VaBeEHtjtqkLvZRl
arqiur9wNkvWR7KCFdefm012NIP/0HpK/DUJ2CFuY/utRPbF/ImSqnu02nhXQIdF
PRKx7LWyCqdeGz7UO09YNjymxocG9xbc/i95vjH0hXImpg4G8/cJQuP5qRYscuAI
BxCw9/9pzbmsVXYU/oDn4oa9Jb3hMOEs5t+EV26XD4F5nXmx42HN+OaXHAILTO53
oCDMHX6mnMrU+5NYIfLc8MXNlTBqfWIheVwqqIs5EsCQsVw9hK0+xlrPRCCNmfC7
tDLF1Eh5DuzD/iOR3JGSHv9cQ3RP8uJGq3c6DmPFnQxZF3AdYZPFPJEMd0GI91pW
jl8XG+9uKtYPVQ+hkMu4dKSHaxxbNla2SHzwK3YcW1g5wenzXItFuKup/OLNP9j1
7/dE+UNd6vjflaNsuXKHypOaq4YVU+SDN9hS4vP+PIxFBFbX5jd//Wfa7R9DCQlA
zEcU3pf4A3IbP5AcK9lGAXJk49whyNMeRZ5GXDTcZtj2rWUDEuSoGcfdNUlwwDN+
Apxshcb4CvUa+GTO16jD11dBHMy63Vdg69fVJQhvlfZp5x/68HmInfHiSedC4ZmK
LIbK4RGWWHGGBpr8938sNqTG2MwQBDkvfdGjqXic6wXyn0MTm4dz6G+JW+wOEPxx
LjP1qbdyQF37zu+w0SDCxg6DRqieI277zrxyniXcTrMT054wHjR3L21VbvsgCL4R
Of1vh6+VMShkT2wf8gkAkBaBfeIKa2UPoJWMK2bzMpipdLZZQXNlGCvijoYWvIKl
HSw1P/L8YomS6AvMSOMsRbMeylmdbBr0BdNxZkRSDY8gQcU+4rLfWDSIW18AkOjX
F7hyk5drLQGDP6d3T+f9uJQf0q0EgYVt2NfIH4OwkBh4gEcDoe4WUljLYZgBfZ0q
tc3LY+1jOhyAeoDcl8swOJKh/ugaHuJ5GIBx0PhWm2CAS2j03oUxPmDQMiE08anm
yN8oxRpU1yLBGfXHFQOdCrJn3bSphNsSQWiSdls5fsqN9rj+9wYoLQkuUKYtmAvc
iYWzXiEzFW6+j+z42I2JkTfUk+uHi/f75tzS7ssPm4LCIe72mhWYn//5eZSqQWDP
PNus6Upy8r2Fy0FiQ9rAYHz1ILOzm9Qm8ri9ui5fwutBEy4pFJQlSoJaGuzZaXMG
p3DJLRE5i/VMZ7uezhpxt6elFRpVi+A45pLx0tRQAETQJrVZO+ttoulGl7pNu8zV
np9c4XKyzw+nxKFIG2Vwpx3OOneu2Z/6K3u8wweZUuxQQQMQLMsjG+TXyYSLm0up
2UCVbRrOY6DjS5OOzugu5YEaX16P1F9QK31wpDorTDOP/LntdOx0ztlqaISAw4YY
oXECxagF9d7lCVA3D4UAWzKL54fxTN+GVKp6tMBTXu7gSpjipv7V+OLvwHbS6qmR
fjvy8ZxXTPnEEu8VkUXoQKW8yJOToTa5xBMG/RzPOCATZSJDEj0yhLJm9D/Hc6i+
jVxTdSs/2Q4XHbQj5H6ZY3wn8Expuyb6WUy0ERFidLJ6wWM1X5dH1GcNhWv54kA1
T3Rd2obzFnZ1CWUuY7jm7aLbMSBnTuYAa/iU2fz6/vJ/xUWfQTb35LE1yZUJS2Uu
WGRmHK5EhZaT9CNrhYcv0bK2gfaV5KS9qlMJLK+VJ/lCfHdwdtRuEVquibXXI8Kh
vX5t7s4MVs0E4diCiPGp1tqAbvCCD1Xp0ZGb9i7DQmOAdCeP00TbmxDkdoy1hlJV
n/gqn4ByX8rANvhwP8XpnEWmP5IMbRrLwnmq1QGBnDIfrViNrnMQcFhSD6RneDHc
JSFG1nWCLnw5Li3YrYfWK0ukwyGUzdof/vbpGLaUKEqIDmUUy1raZZNkC6uAbH/8
7hpQdzKltYPEg2JzxXALVlvMNdS00IdQoP/O7B5ggb0Rdc9d8jLWMLy5P8uTkb7o
RnUNjm1qNF+r+PPOxmDXou16JOb+/CUfev+b4EZNbf82HnBHdlq80GEnV4TKSSJ2
DLX4Da7a3ayQdMZdm2gu9/6QaFWjEmrWPgZaufy9/x54Z+inPTc9XCPgP8TxWrJd
LhZaX5trQlVNErDmeIsw9/U92gbyQRvDi+D0Qx6Dg2xYjLk83Al0fbpPYYPRjtwE
Ew11EX0xnVypTwZPZjGB0hKN/thVi09IrxQlkY1Qe8zveXQ2N6+ScM9syexnOxn1
O1jZ00LLK+r1fhHwCnE932rPSnZhX6An0XQ9nhGZtrDC3rK9cz32+C4VOUySZYrD
e7Pw7xBnaDqZFHwxaY2pTH/+oY0l0Cvy8SH5zRFpVt0cBGWyIFzgkW6TX6Q0C5uG
fq8ra0qGs9v6hm/+to2kSvL5ltaoL8Zfy4rOC3rXQiibHpFAY+LjvcYomw8hyLmf
Uc43PDjJijEYvw+dn8k/klZHWJSkdRfRzcP5wFXWYlzj1mptF948h7CUfgqQ6gPr
p7zrkRnBgxppQh+h71yf71Fc+QDbJI9P7zTIy15CnJgRRFEqPmJ1ISD1ilyvkNCk
yGyo14VogZqylIrgW9jkVsxIkOcoKsspPskjG/QcpToIW1VYD9qm2HeZwUgjONTz
E+Yjw9UY4tOJ55pLxjqWzZwnyW805FXM2ao+tIjj8o8lg1T35tTJKikX49Kr+HR2
g925FCU29Vy+ji5+jwSX94pSoeUcU6wUyc8Sk8IDvnnPuNLUiYZXfCTvuGswtE1B
ZF3edgFHLZ532rYcQ8RzVze+9rlrrTxRtvdEeGG6bADWQ2CvYlMxRePbmRxvT5aM
AOX+8vYtPJBoYSRJH2PcKVpEBz9LWIiPFMOA0rgRFZCqW3Mw3cg0hqk6Gskk66hq
rQBbLkVITqWy41m0BtVZh8DDxD33ihLLKWuubSqru9itN2h2I6M3PBRxSqsmxrf8
vF6kkkjEoAS0RhQqxDqDkBJz5kDWSb5iRthipW19a8ErtMjnhXbtIhyaAM34n+g/
6mO8xLXNOiOHD3BFD1mTgBvSMBr4NBcFZm9cWW2eScWlGXXYGwmNpkUa6bW8eA0p
9rqwNjjb8Pv21BXZ0NbdxAwhroSU8SZGEyuV12UtiIOa1+MwZjBHQBRlwT/+Lv2B
t93QnrvbtmGxmiSIRaWJi01Pm90IxNEgC35DZ8vUpFa+aGrxBOhiLElakt8mpqRZ
X6MtXD6uwgqbtRGknjseyyUy4x9Tiqw9tupKw127EheBj6+y3RIzpHJtDk5AAbqM
xs0e+6F9qTV9knBBOGXBGvgccrR2pjlCiARml5c7NAEebcwtTrNe1izNsfA3bAvg
c9VXOcMof+tIrB6o2yKO8jZI9UMJpfe7FT5Z6FjvKoUW/asIMczK+v18HUaME1Vi
SkpSlIizyxNr4sfWpDVgvNistiU5bI2vTaU+aBUmqx3uTnVl+OE7G2NZUjg+sIK3
v5TzMiCWq3VjHVOQS4SDYT8PpiJ4bDu2MMRwB7+vzZapJTFhATomjZx9S2wnLIfg
Q8HE+xppMaaRdDipslEoQ7xaIJMlw0zM64cGrE/gbqou1b9FdCAvZmjjBrcyniFk
2UPmdpCZAQlVA15zfCjC37Ay4NMuRBhriYV0cdP8Uk2xddUofE9s1NE1La0Ya4Nd
+9rJxaQD2uts71W+pbHCNrP3ENu+jCdOIk4FWgYOtyrTmKZk1Bg4U78snHKOBb5J
I3TlWE0FGdIbvr7W0f/jrPlmA6/puxpF3b/5oWlrpLaYVGe58dNMXJB9ElgOkp64
PVZjTXFYqC7boaBwIwSWsT/GGdOCEy5yTrj81bd4xei1st11D0Pu1dBIX9CfC1JP
/KnuOlqC/avtcjEqKGW87XGY5pMOjFljH9m5ILmSy8j8eQ4aaEdAj3X2Pe44VgAi
BSFiFaPijNQsOutlaH4sAhst6HhJSH6on9m/gkqwhcyIwMwF42ppwAvfaETeIgpW
0BJFpsmwNI4yMMPcTLykleAQlcfoIZ2vt15mkaYb+8RT0WH4VQcm2iNX3ZUwXBOm
z0vvPSycaU3/GkjG9ZxvoY2pU35zOncnic4s/094YZ/CzR8W1tb69HxVVlk/QPOo
hsj96p7q6hVmJfHAZQ1xmxPZOm1cl1ySdruYq0JUhYqvVXur/5UwgFxTDk2YKlo4
+snzWRRSqyuWr+B1DYsyg1tfG0fA4bBY0nLTGd39hTKwMsEalJ1JLjN9XplmG9k+
MRvM1rpeltAqk1pXvlpeDYGXvFhx5lJybUdUeV82JBYYoMttoEtquw3kUnVCfRoM
Y4T/o8ViJ0gauM2RO7cQdw8n6wK2SbHKHt3f2+sv15OX1CPeEO/jTyhz+ddke/J2
J4wideAhs0T7+nyqRpJD2rbzIA9WF/jlRId9oZXePYTUXPQNwtsH5V8IbDaIakUs
2ZEb+L7Rrc1Ri9t7g3JGKYKyq5Zu1z7LBdZ2Jj5jCciW2O8qMSORKMJX9eW33882
w5TMyLuAD2NMPyfG7EuLxx3mV17yHoLKy/zu1ApRAPxL9vTL2ZFjT5LM9SnR90L5
z68RcNA/Sa2Z6OL1htTAtla0evjheLfbtTgmgiCtox4GqaCJ/FLZnZn9AowLZXIA
WaohF0Kokf64yUGOJ5/RnjHz9DLyh1C+PLAAAajyadj+qRJnU5COaCXXhDoqPZDO
FiyhuBVWoPxn5nKUR19JDTpb2TcFKqU5zK9kEjyQzl/S/5k7NKwCWqwYZFev11w+
RWgytj1Uzayj0/vm8aXgt4s9C6oS4kSZVCwkiqCemG+vKxtzspfO7JVInOm+9+v1
F/EBgsHMy2Ap9XKVxyXcbLkJSruG4E6QgosUhzAKKUD9HPIXbtJFLzdGiP/a35IH
KC59F15VIbGBwMDwGHVk6tLPM6N4f2a0YNtBN6YHnQP/zKWzd5wQUkA9z1eIifma
RYNjZ7TM1aAjTJ2O51alhzjzo8cjjjvHyRj9Bt6jUFh7w8HOmTzvbvChemFl8QwF
ubSOvxaueT3Y805YSh3R7H5z2imiGJxBmsURTrbtl3RG4ageycr/b8RLhWoYxQSb
G0Zu0s8LUWTL1UCAuBeVeQ5IC+Ehfpsf7dELelJuqmKFnMrygeLAW1MeXn5mCq1s
tj3uhDlrpp4NJBNH1a6eljRYNOUwwYsVhmgZCHznYjsVjpSRCRNLrIATxlMxbp6A
nENmRRkviQfeRIZuamj1CxOzwps5r8hdCxsIcxm4IOwW4ud7Ehadnsvj/tqh9XV7
Y/uPjFkmwhYDT9LMOTexfyj6xwwt1JMlx9vTrFUFDilZK80ZbfX40gGi1zqXAgd8
jMk95K0cvL/t86mOBO3HWMBIINNV+WixB6Ek63WuF3taZh0VVtROizw9/qXmnlp3
6vmpK+1SwW3X1Zz9hr7m7AYf9QzDvE9p+KCAW7d1wIOxAQFVipluW6CaUZQuYQj+
MYcBaQCMF+ch4AeCKEPLovpzAOp3d8Mu4oaiX5rNKB4y2LQ4EA0d7Hcn0E75vB7c
Bp01ix1cFK4I6/cmtlvBpo0f/mVZjDbhfdg0BjgX962/lYCuOFanma54U0ZTXsNr
LsUVjAc0PulrnG+k04KPycWI0SzBdy+6BN2Vuw5seOYPBrDPghCrlVcFi3AjAzEn
Uoc1UE/5RPJR0jloT0enpQ7dzfcVLaluDhfxGfRyl77WNrin2blggMgOZ7k3T8OG
MvN18iCJSEKapevbC3MSMCMq0teEWBw+2RbrtZ62yLgDOa75RRmnyFlNr/MEqqqs
kLawji5/GNmx37GHNHkqv7X8TXZzbB3V3advAduvsmOgxZ0O5jUjlNsv5W1+ygdb
XIHM72zWCG7YsdiIa67QbNxyHyNCogLQvUF/EtpccxVEhtTZwQHqlF5B0GqAEjq+
W/B7qR+bMp6wSBVal24OZV6Tl92wIVgwf3lSW49jgE+bdNoZCQwPOVT+iyNaiobF
4fi8tHdtouxd35X8S+DIyIFHQNsE6vUo+i7wd6+l+DJdRVE3ECk/fB68o8Cr2+BS
7l/LrsdMryyUZY4VvXDB/AxydVfz+qlKP0gat9Xf4Y997kDhBMqzGokP89vpFsyK
2ta1XlNQcFVeiDzrAHOT9FryzbXyYLscEokN7WJWY+36zIPY6dzlTNPlrAMudWUJ
B1bOpVotmUPSCkLIzM/sWRYEd7sImNbTp9ZYw08VcRPRMqzq4t/tJZ2lABVmY+iP
RHjEW54U8vh6iUteF9avwUWGjxwqIXfSwvybMImUlkFe43I3zrL2yuChfiLona+8
WFQNcwXr4q31Zg+X1kJiwWKAYiRmtbJhl0dG3ZE0V2YL2JJKRpCnm1Ngfm/hvi+3
GLIpWRdnjg/2TOeWU7Or084dTdO9a86XNvQQ3o4pBVJjGUwQy73J5OY8AbLFHZwT
30/EjpX3nDAs7pdigMpkOLcEeWafPUS+kJUVuhfFAOGbqfxg0kvkHnEbDiXPul9S
Prmej43kQ5d0604uxOJjnT/+OTEdEeMeMEOH0RBZRcGQHmf3NDQMI6WmiYr+Uw9a
JcfolI7PmGDxskBX8DE4apUWIJmwnjVRHNQ/nD/BgpWheLYs0/CYz/JK5sKcxlfm
nFn1Ymgf+IMIHtz9AmBywi8VSirWTKpsD+zt2rCHM4/ie0ZQT7W/6hV4L+zS6Sh5
f+7FA2DkNQU5eMml7Wf86nF3IaFnjvn5ZRHrbRiLHyfKc5HMHNaJCvf3o22Leq0M
YGCZqYJH32KkKryIs02/g+4180OtP6G8UW1UoI/ja4P2Gwq0JiZIaDemghjN4XCC
0CC1+bHuirCiqV/wBgV3AWRJFMMb1/FQ5hh+iOPHtbrU69yxJO1x+V5XOoK6ygJo
t8CV3DTfN5HNGFtH0G9iqHQ3vj9+SJOLLfRsIKDj+cguiMFGy8ii1+SNK9bDiOa7
tq2MxzMTNuS2as869T3MQU7TcBBZddiMrRor5bT9tTuWX9gIVQmZ4UPDjvTLVBAc
P9+sfs9hT50v5hzJge7iISgb3rtRF5F5m1T4fLkYud5I1/ArnbIXIHTGqpEYfnSW
PhrIe5J4rw/LoHjZI0KMUTvTxtpdCrmiLsaYu4a6VNntTT2pWZaOT0+Mdmp9QWFR
+r2/pb0hWXSi6uZs1C33gJybReKZ8HUQouo2NnkImRSNpUQkhQfBvqy59fmV2B6k
HaseixCfG60Qopz0B95txHd/UWEQQa+J8EfllKGDg00tskJ1jYvHlZBT2R8NJFha
6DDW3st8juLc7COI8Dbr3az3Bf6wLnVwNRGLh6RWmCMtXdoCTN9Wg+xUqfH/laNO
bX9sRZK3N+zWkBBTlfkwJQgAu0pVh2tnxYt5jMDY+crqrLLjGeHhJY+9t75MsoPm
6lEtMG61qIjhVmjGbrd1tU+Rm4sZ7stmqwj42HX5VG1biUQi8zy7okRdJkza7n4C
YeZzoIplckrv1jOTN/xpUgqUjYUvIdckjV22XLbv6YzxsykBFm03XNsQWzrd5IHA
xrJgHlvPRkZNRCIH2csjE3OCPAJmGx22vPbk1xg6jGEa/3Xmocv7ohdu9twMnYto
0DFO1jG0II0kJGL7x4AksM2jYheZsiyMCfscigszJhUDFHVpaqkPrDqwQaKlix2I
q29N2ING8rbzDZv9wiWZRoNMHyod21L5PwiG4wu7ZpMYLmZvZRLRPDQx98gT8JlZ
XF97sAKIZjhqkQu2fUjKRYJCB9k0pkMEHlU2TnuoHPUt+wldkFpc3oL8lQFHleg9
RgI/0iYJuuZcxGvHdJ1wHThrQnwDMq+4MJeCbDJD6GFAQt3AIBAx9Hunh8utySeR
n8fWP5gxtiiLcfaDlLZNJEbrw29T53MFq4iPf+Jw3J+0iAPEnuWuirSJ1LbaWAf8
f+v3Wp9794ZiMIYDY5QABGXu+bBwXfts2kNgy4S9jRohs+I+sJl8+LUdtLmSFPbU
5aLAnk7HVzxT15yMMH7CIGpbUXaoqe0xdGVTPXjYuUbWLwMOKR214wlsJRt1mik/
PoDLjb8P/9YnIx9NFKM7sCDfE5Z8U52c3N13eljuzucr84E70RNpfTeCn/HC3Wl0
2kQqd3UivHgHYbFnvG00t2cgZqEM8IkZOOUcHMXMaVvoCG/WQ5N7fqt7+D+fW2X6
SKj3Wl9wz+pxB3Jy+DSW9FX3hDyXQpzhCL6Sp/wFCOsHGxoTQXn1WSFpI04X76F1
G0WNXP+yWMii8Ad24H57mcNBAatzUDyywCaBa2HLB+BTEWMMgldPzfy+aprsMbVX
DEpan1MJGtzgpbTfHi96QGDB33P3RVJ19O6NQmat1loFD+nTl7dpVappDAWUDoVZ
6urNjhU1+fDQndL1PPmOtpLlabMKYb7TSuejt17vlxHASj5W26W4C8GJPCssZ5Vc
kQ42TLkhwkSqtFjlPRP9M0UJN9amiGRePN7PigihTKhuNGrefYFlELzutL7cBQ1Z
kw8ca22znCPgeHR37s1KpL0ehIww0Q3od1mYGgvVjyHKj/Vw4ogFnjwwb3IcAlgU
MV2g/LSWN6vFiRVwHllpGrIU/VQu/QdjE7zuYlIK9DHyUme14Y7kU0Tx3ZWMR8/9
xZxTtWESGt886L695JoNIminSvdSmtd34MtbNg/dzH3hih4Vz6wBRT3VmXaznhki
c1ui6J36suJjK2LKWb7A4JfxBfrMgSwGTsmo0E5dLUzjizWJ+piubJypmCbEiLWi
alXxLlFs8LaPTUASqHBYZsS0YixszG8L5H2H2IlA2ZmSUj6QdT+CR1IoJk+VL65H
B0r5BAzgcm0qTNirk549QfN8+3r65LkSyZ4orxEeHf6utmB+EpciRaX3FQtSL8WU
KGxHlsJelP9pPLfUxDHKONxYRip3pbbPytz1PBFb/jQeUnb0xtUuJkAFiFvJ44AF
jvdoukq2rxqx6K4N4t/5xBBGo/9Jg4O2myGPKrYpoBrUc1iqHwqADyugXw/edWd/
IfsJyib9C+GS475pz4wvZyPssB5gfmVqh+1PJPYgCQ9AH69KjUaOyyOqZvAvxNsL
gE0iL4avx+JHukZVBVfvM5oCSih93hVeXibS/Zdwk8ziEiLbRQCKwHsJO77E0dfw
CBbv0UkbQg++qsfDQ71KEg17yeyMc2FxotKggGVg2pNwRcHzl49UEDT42Dt8vkL3
N0693JM+tG/6ZZrUOkq5ELGHL6uSKMW0VbfyeI+bya18FCY4QdkckC+Z5SZix9Dk
+ii95Dp/ysyXTGv1bpnKNdqtUPZOGUAUQprBInxb/MW7luVPKY0b4N92+iqdfFUR
xW1krlHAfoAYIoDFmR60J30n3+P0YdlkqROqUvU66YpSHBUtE+sGjeAIjX/l/ssg
9OFqYsrhq6hIW7lXyz4/sIt+61j3w6zalMIp+tWNw5DxK9Q0ihGBULY/Jrmwjr/Q
d4YfUOwd1HL9Y1BfcqsuEv8VQk5ozaDP4mEKbM89zTarqL1rHcOTcRJyvf7A7VIZ
Hi0PL9k7XbqM5hcPtgvPzfdxPUrmjE8raYpASX/AA7+0RUrEdOtiiiZLHUs98UKH
fPgt5ERm/TngSdtldUIQiAYA53OWuZam82JUhY+fhbAwzrwZkrohU2aa0TrDfOg9
yjE9gBOC8CpFDhIkPuanMJBCZ80R4CJxYpG9okyXZ3CsbAlKZtYbPcdgyaF7Y0iC
JPSG0F8zemgz7bD21yc3fHn6z5okBJd3etccICuR3QGCh5SH5NhPg/A4vnwVKX2o
SW2ZASTZeF+2vePg/LOcvakCuhea+oKBUfD9zkczZ5gtBMAh+s+h+TJRRiSE3CRB
Q/d0okN8wg1nsAQc5o1aT4+ulrJrAfq5aQoco9Rko5fO6FYw/IZOhc4L3tnza3hh
hbS0vUmms7InOpGXJpw7zH425HZWAUxPVYMbpdh/0wcRszVb6I9QA5cyp0eEU+8Q
1GEY1gmBMxtKmoD/4XXoqcHqMub/w1HT/wFpSWoHsEU8COtpMdACUB1OdXo0nCMU
xCkXdD3qH0CGGIqx5Ufoj71ecszlqKy2WA0bWNSHcR9x4Nx5/LjhC9oXfQ4fFKfN
gRloMhIWqTUE+ndDPE6hhqESb1ISoWF7k/x8zCDkomE0jLUAU4F3MMWCN8KyjvV/
EIiCSe8IiVnOnKCzYLCaUoHTOz1k196Dshu5NzlcBR+2O3z/8YTPd55yDvj1ymwC
ZbjwQ7haOhPhIvHso3u2MBb8Oq+74d/wytgZn/fw23J/+Mrw2yVcRWJ6r1W+G4ex
jAKLv1d2cAIegfKeF4lY+N7mUaFQjVBQB3bPcwdL+5XhLpbwX4Ru7hRuknANDjnI
EGJU7PGQLQNvAQLIbhQ6oi4CpxstLK5jy0YQbaZ/g7VmY5FYxbZdpQyOOdux1aiH
qTW2ZKE8sMOjF0YZ3Z43C8/JwAC+CxY79BuexNLwh5kJF3lq8inHDdA666RKH7Ze
s9Bi4iGp497BlJeY7aOBoarWuRyb75mA6ecbpNJhlUvowJ9lvsGy0tM8BhsLKYIn
gNIuEhu9fKiCn8JVq5G3eEUsUlGhPBsVeH8k1C2maTdCYbWaaXIpDbxTvZNkZ1wY
no28IG4f+rF5rCF0xrAUwICjCHscGs0DysVFdfin2/2FojuWN3HlhmZ/OiKjIQb/
snlrSkXZXIISZZiSSpvtDv/o+JokuRHvBue9zAgh98R7juRSO0jqT3QzRMxDiNnC
9HRzkmYvUt0HB54RedtVdCa8cbqSwp53d8+jLGHUNd2TXB3u2GyXrJDwKQ9f8IUB
/HovV0CvKWbo7JosmJTDBUseijcbP/0Xb+kat2JTDOf4UTYuGDAbW9c0i8azG/JN
wU62+HCptQBUNwOjfL/WkV7Kot+UYNYgv7KurmJr6vLw8rMM/8HHBqWfm1jOfQPu
Iv//PtK7vgG4lHC2kQwrgcnP4qrByM32nfZswUzBSH8rfxWTXnAK/cnk9IuUjmeg
AgaNAaBWToI4bAiJi4TEbD2ObqSPOP2H8N6D/DXnhvvgrpqRzbgCKoIaIQR/cviC
3ND8rHA86K67q9m8kq4n232Qf53RlsKXRUlNHIRafEZJzGKlSYQlnAo33qqBh66D
/3Dr0gTj5qXhsgCyOboKzoPinfzJ5uJFnsSfa9ns2WrU6U7R6cdfehgG7D2nFIJX
MokFhzS4Ou6CAMKBoyT339YIqnYTCc9DnQg+0tpFMWe47vJvy+IREWXCc+apBSrN
2u3BsbmcjrD3+EqvFYPCzZsq3ONfBrJbTm8oGvCAMkbfB2MHNbQ/oCSuIcjBHyx0
YxMtZBpZBy1FpjpPZpvwzBpWP31GzZ7aIMYfjPzZCw6yLNJD0kAuv7KJWFujZ3tJ
h+YNtPFcY/ECoU5Rtnm4fFXQEJ3w/mgSao9V2Wy4pyIgoDJ/B10w+wwwKWurrvZw
lYV6Av4KNzsK6xHV/UIAdDn2z0GLoAQLNVgRf2qe1gJrO8gNSbYJhCBvSQHeNGaS
Wof2rbXPa+cvMsUhguefxUqsEm9A26u7hcgu7UNL+vW2vB9ySfodoSZxNY8f/eNs
F5Ucz2eJESnbGxmA7wqWxJ/TEVnWODEULJB3hMks32cF19PLiloVnIpK26l1BL3P
IP6sPzn5QY469SrmicUmqddiY3xWgyZt2cF0UxKDip4nwAF7wKzbZ0IPima5AHty
l77FPsNP89tNafIWdqGX4XDjtAiimsZU5CoZtdZcBlUTxNo7ax+pcWBPuYjGIEJl
wvUC2jugTYMhQ/68vS7k3FNsAtW25WeoOZn+Hr6Xy/mfC9GWarOfMIH94uFW0BSG
GV5Br+jKkPUUmTeYEAQE+0nCHOhbvJS1YshpRprwnqSYLVM9dhLxpiIdIi1gDgPd
sy1Vjt4EWtxePR3iPkC8IVkLGIw1tFZZlKz56J+biC2DOhkKK9/GmGeYeOMUlJdE
N4FJqqSN5f5fjMmFSh6sR4J14a5z0gtk+PE4HuGci28DizuLwzas0vc4jMorDzs2
jAo72vjCnTtZpWFA3s8JEDjwTQq2YkYBxWS2HjXKAKewM6qi1aPOeJiY83CM/7SA
+HJMMS/hgFGXcNRevqVQ+asvkEQzVkttm2VMStifuTu6HhkBcgujFx25XFa+dhxa
VGkBwoIn1Sbd/Y5O7UIcgCPoyxeuw23+7z2L7fEO5Z8/mu0KUlgsaawmNpiSAdy4
cQ33/Q7I6TN5ypVYoe8807QunnuMuEEbWBg0t/1gcI4yRESv3wvbYxjYWXPSeeNf
hZ4NpbsZoajUtJ6pZl/vkddxg7yMdpUTj/ywmCvC81E58VLI113kZvtOZshwEFtV
SQ36O3baakwAMnbPmDhGjzrQWSCSUayIfJaNPH6uRMFEOudZ2naWRk09O72zbzeQ
u2NGZCa53cXChq54pNlK5WOim3fGwoJ+23jiPX64YAxQfaALnLeaOkC0ky7V91za
bTMd+VZir2Y65KiY08CMGXCXfODUN8VflupxntJQ5QnbYliJhu9T1UKNwl+6OajZ
u8Vr4TMS/3XDKZGLbn6y8J17sJtiWM7bzmjJxgwnKCxWVNuoStzxdO0DsE4+sLxZ
xBVt8G8xZZaKqD109RP/EcaIDgYJUYuUkLflEgjfDAtaQ0xoQJRABklAkkkHesmC
Qfi1Zb0mO3HOYY3cZSZbOQqWCwWYlcQoOz6PmSJIHgsIY4sapkthg52eiA34rdGg
ZsiPpb43P3KNijmFpTy204tx7bd92fA8xrd3IivOeV64ZrF6O00EHnTndgOc1mNk
rs4du/F82pbDSym0FQ2riShAM0drMgIv4uHVCfwdmRi/kXTsild6CRzh+dh4tAJm
yvHYIRokGnYurCTXyb8r9fjeU9TsI3d1iza7uT2jOmGbanbiBUKusQJPBAZGaB1q
zEIPfYYtGCOxpmRzNVPoP+f28efz958g08ZB/yeTPQSHxBQl7IuVH6EXG258JELG
ziGkqWwixjFWUj1tJ0YawsDX5vgVnllhwZgUi0nKr5tHwYry8NCsvpzKx3AzAWW0
Euy/J9E5V/oJxB8NGz1eyK1fA1eprYpISi0PzvwrwFMaT8f7e2PaUYSsPe51hUMZ
NQ6OmNGwCPBkseD6taMp+Vhvq73ubnU8xGVZldiFHOag6sFphtn6jcdf//sW4Rln
/LaXrF7oVaRk1dJTCPDaBLmP5D4L2P0aWFkIRg04D0CS6Uunr2T2ufPQLQ0+7LA+
mtare6HZ0Sh+w4D8I157hFTxszFVG7MxL/QnEbnOM+v74Da1r5YHEKFFStTa4UNb
DX+Tl81lmAreeRWeyOsN/o+7Nnv3htaz0ZttVHdtEV/KCP+YhUZx7ZGDhHck4HS2
XIWvs2BZEhmMqSo2/zIEDOG9RhIU3GC1tUODSY13toWb0WQEULMTHlAlr4o+2Zm9
UHWxZgrmOqf0RgQkODQzcjyHnE19XbFh7sHgd4VRHvvi9eE/AO27KWU7Sa82nAEt
fdol3dKGYZop8hAO4tN5h9CayHn1Gf5CUSfg/TUbVni9DkwKLZwzdq4QapKV2IZg
BmYZFxV8qgcFlh8WX76X8DgzZr/8w5yYdqMTwwVLuz1UJki1ASyPuc6AAIRa8hHE
ZnWSOgqJv2BUcmnVWWJvRmAigpHu6FIKLxzP7mfrNFRYsLZNYvxp+vNFG+zA0iBM
kh8yIa9RtLQmVxNNpfQWFQidl/oQtbuoSi9meAD+vm/HuzjkZI+9kcoIjQZm/9Gu
d+ui6EVg3WjaWcNqnSFbMP96wwFm0dVphphEaerTSIVJ4hr30ID6tx6jVazbIrV4
MRR4jJpiEs85Yr4ZbkkzE+0PhkARwG85BH0xhlLd8oiaTRuDbbwQa7+8J/MWGB+p
l0qgmqfzBzlUmR5e6ZcbNQU48yH6o+gpySm6vSMWjbYUrIdi/DMJeGsZiGKJKGqq
OmMTW8yYAYfsZLSXArxODzSiH8oncMnYKjozkDiAzJwfND1ztvv5AKDQdvpHhQrX
FKDom7MLNaA8+C069Mm7xH0Uq79l0J2SBMOqrpkAxER0fL2t/jCfuOBHKPQUbjTc
dIkJoQ71JhAHzq4tmz7UO7L45Yxj7WUAC9IgLwsMv9Eh1C4j4WLd8BgwaidFqAfq
WLMelc380oKvoWQqIFthdsgodptGpwjSgG2f3trthNKvC9C5/x9ONxPEfJiX/Acl
NR3CtnSg6hr6uLjDXiBmVZKeLj/b9DAxarOF/ooGDl//jPGLozGrSo5msj1GvwK3
DBjmUlIATpuNLZYzDiyVHpLXiAfLmNipo8ws3rz3yETs1dSZp1MioRjbal/KI0m/
aJHrV2UfbAXxC6PGRSTJaxy7yXJAZhkswUw36NojrrLEuiuldZy4/lT+SuJtOYm+
l2n0V4I/LH0qJTwZiVxsEPOF6k454d0M8QnPR2Et1l1FY/0GFwoEhqXhdkg9mObM
3dt80MPe7IHdrT8/QpJFXSNYSSTeWJy5430UkJUd+z1wh9TKRndroEaYMZ/InFS4
rRD2kv12j5vVGtXjqKwxD/848s46psj32DOpmnC8Zlhcml5SuuMA/NCbhEqUJMMe
z826f6Oxv7+/DfyuNpQSqT46cTEu4zqZGit2Ve51kS5Dvsw4hO+FcSuuBS4AJ8XE
oaaorNVGg+hd61ZBzGZHEY5adV13CoWdA7EyPmLXurYdLgZV9kjf+BqAzicftSaZ
/dKibDRb/uoBVSqBUgItc88GBh9YaQoAN4RTYmrK8y0VAcKyNaAibgA5keoEXb/L
DWZ7PQ8CHZ27arMhZhWjQ/STjTuZgk3gLgcewCn1PTVfsC8EM8wkX+VAO1VwYqAF
nTYluFMjlxz1FuINEklMPv7SbHrfdNcS8AulRBD5PKb1CZkvSMA+5jqQw4vIa6KS
QtvQ/BtEnS0yZyiIOF+Y79kT+K3S7HAg5cbCrlfE1KH2ovB3eF/0P8zGRu/LCB50
EUCx9Cot9bTBam3QhdsHt9irZ038iNWfRCAQ/iOvxjdEovw4grpcRCqIvxhcqrWr
JLMCG4O+V1JusrDFRCRfepJwLew/YzgKbIPArf/t+lYrbZx3ypR6CnGRGRekL1j6
97PHqdG5xLSk9857LJhKMV5qZXx+e5jKkX40xQmQeSYJj6f2K1tfmtBZOu988s1B
ZfOnOnigHVoI+/ABpthJsxTNgF3h9tUWffw8qPJduwOZzVcKjMLKhZEsguR4BVL0
l/QQTtIxHRsGdcRVuN9m9dEsxKqk5S24d7UakB+1rBjGLPSj5LJtI2SH/n3hiIDQ
W+GWphr3iAIB2hyUCfPe94f8XvKouTerKKrdKLf2UlJIMCH2XUpN9g7YafC8fnD/
Gc+mfdfBQc2+6K8iBtd3CAj6+zKw4o12Ca3z4Cy7ShKxviQBLOdoipDeqXbD5Xs4
dw7Tyeha1HraSXuOPa9iZ4P73YP7UxlhPTgDrP8coOZh71oZ0lKmt4PvV5KS2SYc
RR4iETYDWRh//7TGqkYW8YwkMnbmpS6iMD0l5tuHysc5ZG4BkQv8fqdCVaSWEMan
/lCDe8vyJVMYyY7+O4d+1wuU6McngcL8fWqlKr3rU/5+uYw1YDJ/6XF009aYEBPw
xticmT3H/Z/8RfFodFr8Y89XRkANgJtcTwBrPXs62FIWEYdOuMo+/urF9EjU5Aq8
Uh9VjwpVNf8igzBTbt0JfRtOXwpPdVX2LrJ7G+BcQStqCZumYq6tz6u0UzlqTTQS
4Rjre1OTaFH4fC7I9JAdDw/dXT0TiwbrXk5kmkxpRUdhhGBFN78eEXgAW5b1fSed
kjwAE5vLzR3il8hDiKDKmK5Nd/tBAzfVfGc+k/5bmYRpxddnPwZ5BoMb4iU3VPNj
Q3+5kydWX53A5p98oyB4m+jn2DBymi5E8GKzZymoKvPSfL+IGBc3WBBMlXKo6fls
PFTnh25vdPIb8vUOCahDutWukuYyMkdLHpEkgJ63ke4m9B8kax9o42UxkzNi9WQ/
X057zr2tctmEgWUcmcvpcL/qz/nHZvT04iMge0qjXGJD5h534O6nKboy/0VYPTP0
KuvmcnEie5XXjuHXo/KA/XF+UqBg89/KL+8XU4WJ6DYkIhyIzSyfjhn7wi5DYBlE
2MXcmh+NvQTLBUTsK4gt0RAbzL0/mOm3vTTHQMdBO4DU0ZUhv94GDiKo1dgYBuik
3FQLs7KnOlLGXPNUeapgAAJlYVttbjNMiJQZBGw3kNYM7LYEX12ykFJc32xR6xhm
VA64ujdNAqvtUCQUSGreWtjv0gZ7szroKd8uMJ3O6/eeRvM5GlaAEzngLQy3DLm9
E3IAIc/+8hwNqEzJb7wTByHIU3Q+N3z7VFgrKmMayYJFH4DXWxJEpTW3JBuK5Mds
x2Hio/35eYkD4nNn93cDiJmdCVmhvb4WFs0lqdYbUvNXfJHqdBARXpxWJrltt8ym
8b/mAB2pA62Uq2g+pR0tdhflbE1MKsZg8n4mkoYOE0PB4bz0ph7rjgns+kUqvcaI
/zXqS226PSbiiKbX/tvbAxdf7VhqFIkOrSKC1yJYQFrZn7IXV6v3IKeVL+fH8X1P
s1z4p5Fo9yGIpipoKxPsof1f4EPYurYyu+DCkgUtFVe5aDW02PhOaC5uTjzEqs0W
kvxu86rn+SjqFqDscS8BcmXIuHY7CYDGeoVEufm6nEZ0sRkCbT6TDZok+isCWJAY
vkHOe3FzTju27jivUNNAHjMMcdE6HDDEFo5i9zuevyfcWwShm6y3mX9QZorp90/5
Y+VueVz+m/18KKIF3ghGTF40IJSr6IHiHpvNSXT+hF4tFp9LWPTtDCILdX5ZvoqZ
9X0mZp0TmG6BWH9GAH88jmseuoy1cKv5n8kswFw7Zer2ly2ERBIOjs7zcmc0XNRQ
qv6kuPxmArnar+YiWPVlpq1evwVgj2YaCmoY0lGjCaY72etSEDkGXm+fxZvvapVn
tIFcREdn+C3rh0817Ohp7+Kg64rZVp7Ks1HXXGt1FiSZMSIClbttm+R8loGqrsQt
BiMNxKsIxypD5542Pk9VvjHc7W06vIKszKpu+xn0GZvSMrlJbSVL6+FbxDGrm5Fp
8FftOWqknrgvgo1ReYokVsG1SCUPWcDpvwp+t5YCMzuDp7vTDBkI0t9UbGDHfG5d
I2kHzilCrB8cUqBCcXvnmOsWJ4lrcxgLUwaKyQoGH9vcY7NJwDsP/NZK1nwj4BTj
EZsxIhQfiYeVbq3/xA5Nr1tLRijLgyUTdBU36/oDYeDlfJYD2JOYrYYob8eIb6oD
fsH7lFHN/C52TSmknGNLIHuUZAin+fFW8SHjbtJyk8F+abysUy2Not+Q8ibfyzDR
nsDWGUbUK/ADhPypZbsNCPXajL8e65sWp/G6YcNxy7TGciUYO5WaSYT9crijJtbX
HIccoA475jqAJbFcVg98X1iVJxydMshOPLhyVvVOZO1ybPhZ12tYeoY7f2uXVT4R
AKSpTMdtAvqoO+ZDgNyGqSCLHk+ZMmDrOwM3I9WqOLrBv9TerGBAEBQT3/wx0PWp
zEmXg1poZ9EhbX9AcCnx+wtlE7K9Vl9eTCBkhnlx4G7O34bk00yVH61exhvUq6Nv
iO6RmmTQQYFiMSCSSurOJTAtOotDCyTyyyS7LTMz11T46qI/s2joMitCzkjFYy5o
auXYLL1OBxnoOiDaPzph1FqL3JH6NwF5hoVAD0hnQCJzYeMW9zVJLUP+PmhoGzaz
EvOV31CT9QQlsaHWDlp/tUR2f8DvSSY9HYJGAULOG9TKlv9GL9javV0X8UPpKUwD
Yp5zy37IwyxcRT9vqLqSgkLqVPLRnE6Ot23cBb0Dj6FbzoXU/cnEKLbOe0yP6OoY
jPUq8bmbZ+8s0mnMmtlC8hsQMy9wzOxyrfRuaF+XF4XHUdZvdhuPSVMMJnavMnh/
BQUQqd6uzinEs8ZjxUvo9RYmtYbjlf1xIph+OIGTqMEFUMzLPtl4FDxwapOqXo8n
03cFnBAXQ0Joola0hKQD/6O+wTrUWaXhMY2ye5rnFeCbAai5CLLp2mPbYg6Md8o9
zMUl4uBCxI7YqYo/NLrvrko3PdMux04DgEqafQ6nWzrJCLjWSMahYJFJCnCWWumP
D+6zkJRa0iMLvNP7nkIsScZNHtPcsIZGKlCPq/hKXkVA8U33R6ElC2PDEd4ohOA1
6cvdTpTuwE50G8jIX1q4YCNatbGarnKnV/iZTrZpB8N5M/28m3+RdSEccnHXrOxJ
1XrW3J+DEC4dM5ZjqcdJY0YQ7ZGx5EKmnPA9C0/Cv5+71/3dL+RW0yD2elEqM6oZ
2Z267mtp9gcBz5Wm53X5+8NwFoYHpuHpkSSzScu9y1t85vIqQu7B6OBJwajXqcmB
fKylfXS3wEtMRuowCIZY3YpStEKF+6npV9RbFXc0b2tkSYMElu6z16GMN8R9DGD7
41EOFGTQspPk7e5W4MNHyCynGwMpxrksJckDkUEpNO99CJnoy7qxjdOmey/vk5hV
eavyiwJRq+DDogCqrhBVDYwMYtoKbIbh3kdvQrBvIt7qFnqc32BpuhrHHOkbdmYB
An4gt1QuKTY7fSWGz2ckh1PkeCYKUk5L/b4YhLMQ7ehcvBIJrU0PS1EYvIjXk3BM
R0N1EvznZhUOsZAU4av0t8tF5lBDY0E491k1sT8CuSVXL/ak594aPM9jYWxA8VAT
TlFYuCjRTxVyN5d/JAahm+w/EL85LEsQNpe9i3cIwYsai5pIgMTszDIrjKUZI1y5
ppBe4OIoB4WXtBKMbXr9xPytx4wAGPQJBYrZR9aKPgVKHDaSpNWun9BtCg0Acons
xPVZIzwffZd7N15HdpehmeGSV/l08aj9IVjB/yzfUSC++vkXRJeUkwUwGvxWMrGd
QJQqKKnuQMmJzyE8xihg/nDLx4X7+nUIv7BKOzxooCJfNCLyVfT8jHd3rTfHSWTp
bQWfVXYZA8UTjuC8O5B+EiQTtRVswOdlqHIf5gFqQK2PfJ7omNckFCS7vDTLSgh6
Qdk7xEpAGQSlmuDSWFeNkNQTb9C1119ffypg21D9WlKz5U/kitdHpKvBSu9j6+gj
xT76lfyyNabfGbLjqDWWPt00EqUsYSd9q4EXjWqJ8G9UbISUKEAjCLBJd8AmB+e7
X8/Cmz8gNfGUaUk7I7rv1aq5E8r/jSD7StO8SoxejsN2bD5djKyISuxzNW5usqin
XpY+UB8esEZwgSpdzeXuFX5TCLmp8tv22FpII41AQ8bYUKRtzJcOQCWsjYeUWuZs
66isvswj98dfW8KFrRhwo2Uuz9kgKkise8RCCdCbcfRG7fV7pX1LhHxnNo9m/V37
fT3KDfzIr1Bnn52D8a+rn/v2hdwvlavCVbu1DZAU1zb8zzYXrloQairrjgOwCcqv
Hz4ufr10Iij//1HR5x4Ka2uJxynHSKpgGwT8PDmGlAVTYxlBrxHaMxcBiQB+L0pa
v01Y4Mj3Es3xY0Lwgub2FFDyH+Hjm6q9QiLEgm54UBqFtdJl3vf1H1GaHy/eCOpj
FxBFqP9BwH/3+6XbHvn9eLHC13gFAmN1b2t3dwSz0rAmS6hbES7f48Jxj043kjUf
q4Vqh7f1HHV8ERHXVwKBnwebH8gpbc2BPfg4ViqiAXf70YLRGy/cYy+E+c7VwKOP
zRFsTd20qHE+it3mbs028ymAbzZfqCQV+NH5H3jClVU3inzbiuXZ25BUxZv+PT9D
7I5s+CT0V9H8av/WdrSTpU0R2sX7V/qTunk+0mx5LyhBpZsecmf56X4jIEaLvu49
pDJEHsCtZnLH+8yQwP4gkx7Du4d4HPoCkJw0YAnrD8KWK46V+m8FjlehKAmKOaQj
XX8dTBVEYKYw7cgM2K8Y2cIHO3B5WrjsBgkls48McH9m7r6Ts+wJThDhL0phL91/
gftkVJG2SEFrpF6ME3mShiC/rzzsj4mjgz3RRzosD60mbi5BGBwLec6Ucl8vjQ6j
s6vMUWJ5IX+xNlTW+mQct4eikEfR3epxZLEqevDEXMJ1DASm30X5v3l6iMwnl6ER
/BhnFbEf+LAkm8ZGccXGJ2l9tiycAhgcnFs0MO1sR0ndtZ7vwfl9tJnT2+JsUe+h
0EoECZdkOoUtkGW2zAUSpvNIdeyM4uK06h/KEF5+SN2tq+mvN7k4PDYUuny/kCIL
lV7uhI4m79EaMPEgV/o5ZRVqfsi1zTzfoCVDOyoztQCXe2GrUQCLAueSC6J2VoeY
4FHKJrH4h2Irshua5+jb9wHblrS94WXyjoaanH+eQaLuNWJJ4KTVHb7uXazUOz8u
VoECYNEBVi11RWHENr82Mg6VNSZFcx0DpwD8+6V0hmGUa+CtGRp/Opol26LJ0chL
ka1OEU3+DcoSOdMBWG1f951MDx3wX5M6A3iOpsLpxm5XY5g+M6qiBYNtcteBEY5A
vdQ52r3ogwPkro51++bCntR5tosFtLH5AynzKijcFw/xlZ6NuIfFGi/DWz2X5zPd
dTeVADKcyu09KLAX/MCPXyAWsabsqH+ptlcSmMwKY2kzalYzmd/NM0NfGsuD63vU
2kGQbMhlBFzEin/TQPwOWF2YmDb7M+PEEQXpY152nTxPQPfCnzFQxAEAKYZ/QWIM
GTHVAw7J93zsAEh/svTWYssWemayDEOIAqwhfI68cjydF1qEfnK9hBHRpKVfAXBb
O/EWhRvOvv/GpDlG5zp5mPO3BH9o7zNhkoaQHeUOJmZXcGGSyCB3EfNiRqp6V/SR
1rfZTO2Jfd23BKsO83FXxIN7+JE09NJC5VdU562O54wZA4ROmsG8fCAth151AUYl
wMKnaPEZdKNPPy9Q1jLpxTllqKkZ52pkvS55AQoR5Sqjj18e2DatLcKMI2VBDV4b
+kRefLfsvggPCO9ONz28jEC4tVDx1UproltBr51pG/wV1CQy6zRBSSJtv+BuIFJ7
MCpNYIAy+Eb2t65Eccj4TeSLINCVBPhPng5CkwYgzKImOGUXoSq9EdbR//6WSBJ/
zVL8quHINI729mRC27a4MoWxTIEnAPCv3n2E8vn/q+Gs0Tw8qZOP8hZAhkkb8X8J
bRusngp699pkE7rrIETsxw3EXp4YrPewohH22SJQGiUxxktODlVJ2h4ugUoR6wfy
6XYr0fgVCNkMX7KGAH2+876nzlI3CbJTkF0p/kKqwyS3lMH89sLUqIzH/qsyIT5J
+gRL0EnioXe9Y9aeHwS9n7M02pYBP4K/Kzq9MPqX+MavP8SlOk3z5MgZ6AT46+yi
MZTFRBf6AmBLPbR1a45SqiIf66OvDArqpjVBlIW8qX2+OfiBwIOXif/aRmY3fL4t
jHvlqoYISRefql8qc2Oi5RmResP7bqEgexLqP7sYIQ7ycBSVRD/6F+Iw+NVGDXDv
N4F+ujEStYPeXgGJKYoRDdRFNXWL2iGFpYpGAl9eTinCr05EfymxW3Sdqp2269Mg
vN6nfFPefl5y+yBUxtV04TS+BrSfv+8wTfvZXBVnwnTq4C61myWJd32Ss+6/4wA3
OGLLGjmGq7c53LtxAOcDEePMTI1VqqRrxvslKGYCgJfQmBHW1XmKtp9JS0hxgNrw
WTsCLrQAImjq7keDU98JgjhtrF+sUC0Vzo/YsJUb8hw6w/VemqM8sNHOuebzJmWi
NBR8+R6wD8+34GZSjNMKxYE1225D9Y25nO/03dQ6t7OfmLseaz3gjAHYxyWZ/KOp
qBkbJbm7Mp6VY+JgKrktW72IKKCVim4gBUlL8Tpwx3+Tib1kjQkhtYpA7geLHhCL
ArEC5ngNm5SWXEj6r4cCLMiMXqQiRz8JCcwZ3mxNJ4qUzJhDddbmuTd0iKZP6ZB6
/pnCY9WlN3N6vIKevmfAWw5fzPrsL3NfuAHgSEWN/aHe0p8ZbPYk2oYMtY5QkeAS
ajoMGOgFq3UQ/rodeKdnRmHsdO32cSQ7v5t53Ju7inVlIULeyU/x6xMHeIAFcZM0
3jEEPcaJ20PXudxKB0pJeVeE6JPGl5eKu3AJ8/6FxzisBPIy9ga4KUnwBELGfkf1
D2srlt8UJJF49G15zZ+YuTdOHxOdbOv/i3sk8bp6tliTfpiQ7F7IIJJ3lXD2zNmI
0XrAIcMgnpw6dLKOt5Cl86qwSEXwCQqURtD8yEJe0Fgxq0uVr9Fcskmgdz7uT+1A
dxUSGlu1N2qG4QCh12ASU1T311CrHnxrPQMNRwZBEU8AdHS65u5D4CXvk3aZpJfH
7b/CvSIW2LA7cFNNU5YR5OKacCcy+Njf5YZJLQHwSsI8vgqYqePmIalM9j5T6/Xi
5hd2oEAbRObCAvj/4s2Kxn/z7RlHdlZPSIF+k03P42AD+tMvQBrnV/BSuQfWIdX5
HTn6AQa+5rDNSExEs5GzE/TObGQCJ/gc4jMzjwlysakWJckBnJz+dFKZTGmysLF/
diaArAJ6VDptVz2B/ncWn9kUsvMkFJA1ZBW40RndDacziaoGwugmNQX9VtyHbwqT
3VZEgYpxd/a1avT8RHhjgFblzEAsxEQCJhjFJ3xfKb7AhPuUMTEx4oMy56rBWo93
6Qx9Vx8IIU3Hu1SP8/kzcorK83Sr/2aUnZTTAcFtXJLXJ3QUKG39JyKt1RTllACY
XcdrJiYWCrt+4eAfZ0/W0OGCAUbsBxSQ9cAhULpBK6BtpBhLsgKOyTmr4NiaV4oY
o4AcEBrcvEchYsEahwfV3eyC6pcPIMbjMiUjODTjNwE6YjAXy7MooXeGiYrzeChy
kYU8BvMZ+wN3/OZy6+WJDgLYwpe6aOyBdPOXfXraeq0AEcVL/iwMzOjUr8bLQ6Hk
ahg8Wnop/FsihY1poLkNxivyNY8VeEIfRs+aUIMz/RWBTBHwxD0rp+fi9pjWswEZ
OHFTTycmzenUVdcVVuMeF6oYC5XJjnDZwMSqEDfQsJH0AVii5198Z/KZDL/sQTPe
P8KUlmhXjuOYhdew4O/EnrH6EGVBImtdGYgQ2//DAWeHqNAsMUC5YV/5SC/TMjto
tWkgcfTAmASlo9r5hK4WFR1j0wGnHWSJ0G4rtDckW1HUm8dleY2YSKLjn4pz8dMD
LqXmublmhpAOU3J4c+13NLYOEeQAuP+piD66AXOUYxWY99CPw0IXzJyUioAyKp8n
XJ9LXZCCtFQz9oFmeEcEGX0wGZALNqjgM8jOTT6aPNjdQLYzprzbTkGUpIPYJZrS
W/g/CNCnYRmqUVlDIPcx6umk+l3kzHqJlD3uhyk55Dl6h+1xBn6BtX6O2bhGvjYE
pLdbE8rIX8AXqWsje1Luqdwi9VWuPb4VEicwtMx9OMXePJltA6AmXDT1aO4Dp+qv
CIKXKAQX59t6W24GL1Kfasqc5nJcim7ly2iz8fC/EgbR+OZRgAtpSinjM2QHa+Oj
l9h2Gwqs7DVPnBs5c6gifoeusPHPWMzTD8z86t0Uc8yMuk8loA+QfdFF2pYqGW06
MvMDrzvduc0/UMs+fBfxF3MZ6Nd8LM6I0wTjhpmaZ5W6IQU+axWbc0J0iPvqSMTh
SdOqEw5cLk7pL1m+6X+/64yfn7mhqjRXJ3f7ZkqztFYWNyteMp7GWtmloPlXAb2B
NEu3yufMk+dskYgZ7DtRrA1u20ZEERGtktzYGy3Snu6YPKasbKpW6TMEdgrvsdpv
v1VP/FlhTuZw6yvrybb++n6PngY7hapVJ/HqeX+Bv/Z1kNJZ2eXRs+nMSWgAbBuP
i9KXTvx/5dobjS9nauKCM04JuHRN7PGpggBQLde/mXsokcbqNkaxc8SoURjca0ls
SzrgFVrAMdmhUWbK3FicTzzuNNmg9pWH5lIquDWDgn1KglbPwZAmZmA1ueFW6HE8
46h0kxGTaNNyczbZLHiSI59e71RpSu+6BFt7u8B6auW+dXqWBF9UVUww6kwlOwx0
OgNq2whS50r+FouxJBqu2JMeN1Nck1r3JUxoULhmJ9X8mTjVnCEh3ylq3TPksk9E
LJZpRJ8FKqhCSaSNXRzQwLzFy1YVXdhRcUtquyzWUjDhL0oKxfquYtcr8QEBQGgV
ArPFXYCT8LIh8csFQP6JNpOkXCnsBI6ScM9ZsfyvSShf2FJp1+O3YkS8HgOcJOtQ
6MOhMOjUmiGI3vffDB5bhXp38O7rhOhyV/rosBiPNVF6PmNxjPX97nxXZS3CMGXf
cATEkSXrl6JK5WNHyvEl3nFCsNkPhrtdfF8lKs3n4NxFO7o1+uFo2hrAgvqkMDnE
XjmGq+UjqvpRb88QRkQMe7Yu7Sj5C7SAuXr4Cpge+ZfI9IyxHoNXrI77JerVZOkm
lc25UwgCyIwuxmXmq7wSTjyAbCI9dFIOu0qfGmPbC5rgZEs3c4BKLb3pBYv7C5TB
jDtXG4NpAkQ/FDrQprBfJQrZHNWvjrVyMcSqChTmsVJ3XOmn97CKSLqYG4fc3CTA
g/MvpTF7hGjdy6jeiNflgAUyustldnDkZ6/VL0VfTOwkGkF8gZAkGR95wSE8tdi8
dtrouv4azpWWcpLcVDn9yQ4Vrr/bAVHgs6VKO8FZCPTmemytu/xpSQDhRWM5Yg+P
6Jdr1m9X5dSXxqXT6sq6/08YUmQEKGrWGMC34YooKhP0Rnwpn9S8OlbB59mDdSW9
DqTIPeDN1J9SfsMs9FmbXNvORSF7zLCncR5DfYlsiFFp1WyqkgfpOTi93OomQt8e
mn7ubYC1ryFuVDBzle6poalqHcIKHEXB7zODhuScxO+2w9fuZJV3H+MSXHLx6MGc
OH1hytBqJvXU5R0K3+lFGiB9trd0WWOVGo84oU9OQYD/deAPnXQzq4owVMpT+XGF
8GLNA5Sag2bjw9eZMvneryqrVafQFZr9raRkk3gbBnNUlNWGtFynvNxpFA35UC1N
DAkr1MdyPc9XzSiYvSnbG/vYY0wIOIY2mzYkHLhaV5DjyVlcB91KjnHBe2JJqti/
ros9GaqSjqI9bRtPVT3y6zffSAAoNtj42+lir8S6+WVAhW42OOpgSYTShKVApYg0
Z6/g1ML9WmqgH2rx3HdoodvEGlV57oo0+IbcyUi23Pq3/rYdXTbNwHdkTubSxrno
+TneWP8bElmSiIgTW5Tl1MyJ4TmZz6Bqy1DZBvOMvyVtFhtOVbP5swmnrvGUF+1F
MpoBXq42VTArj2LIUb+3+2kOkxHw1i8GMnsNFAl3vZrDdNAINSV0c7g1y6Xqjyeh
GIBnmJBB5JTJxjW9qY8udtQUSMKOTOVURaNeymgvYcSwQUivxOZEFcNmedPhp71d
d6SC3DZRHsPQdYWBNpz5mgDVeGuRPF0qEtE0jVRxxNzxqTrByr3wLQgQ3r+Eie69
99nqws0aPtU3KFBnuNuEBAZzjZZdA3y86sW6BspMXRkLIW4y2uuNRyTkxyyxe0Te
V1dJRgiEqXdeFwv/Hr+Evy2tfBnLgy9goCYkAKIL8LHPQEhYQr+kUIyaea4MDID8
caBUe+SNmG1AUXzrBMQxZa79GRy5UGg8LgCk+/w5lVjpacP0/EE+CWYAMgVsW3Ig
AHCuo10+YbH6iUKcqubMYvqKIOcIU3W3RpEM3jKDu16lRY8tg0XDlhtsOGpxxivy
EC123wVIcROMVXYfmOun6vC4j5BJ9t6S88NOb+7+BbXC69L8kBbC98m+1UDQHNaY
x7cuCNoBWsJ9fhKSek+/X+fVET02eGaj0LNVw9oftBaPa1LIi6u3Ma0+BoGZEajN
Z9Ripc5TL7LIKUKNI28KxYYSGOJkP/ReUVw0KFhn48yZGsnHINClmzCdPSe/5Ksm
FrPKbVvRJKe7T0IhAqcZQt3hqTcfRtAgcNKXTMKFOxw9dzNZjHD8LvYvSsCRMy4e
6giUvZ0xzMNnaSBwudN6c6gp4RqYFwt9p1Gz399HR9kmeDeX88aENXVa9yQI2nN/
A80XOKpyV6oLq24lEhY0A+6P7r42TSX1UYJ27DRHMc6tx5mhDXDxDv5M1KEcOxL/
hOdmANbElEWfvHxBntC5zZM9EW+vANJip55Wk5dX9+1Knqb02wmShHXfgiMtWgIt
CwsctSLWWBgrBebF7D1QEY0ZEy4WFnJ4n4+sjggx0vJSMBsIXnLi3WKxFvbHOgLS
vtFRHz13Qcgkh3W/wm1TfO76SHV/QE3mUpd+a0/qmm6OpPOOpEKs4K9gtDiZpFLt
W+jL8OcumOMr3M2cL8tWHS47txjTaGf46VbrLnvgD0gSBEnT/IvEu/lnEjzVoQCR
Sapn0+O/9bCrky0JtYq0gv+kW8W3RjP5zZpEtXnSrEw0B8EU0VQ+jAX74CFdIEr3
v6WbVG5MThffv8kqUAXq1JJatKo+7JqbqofgpRD4brWFCtiZlNTIRNNAkWUQjt1E
NHWhNBXi/HhmzeASDWGUdaCbyauCEkMEW+JX28e3ETXf45l7krbuhWxP0iNEbU5i
iYTi9RKnjbgXEHzhXz33kHhxFh9cxEYNr2/mlAituaoMLtzFwGQBQevdx/V4Q0rg
niXtWH6MCpkI6r6n/yNv//AswgsUgZfqNrpra34X77Y8y97lRvUcKfPR97O5VEXC
+9GXA7quv3DOhK0yzAhi2svmJ1u6NxhAeIbneQuJCrAxyHYfTCKTaTjw8owQ5UHt
NSzp37Y5GSYO93liNmnumgkC2zwGVKQcjI6JB7imwmB8GV939x8g8aim/HEosXzt
MefYkHN+HYuMzPiQURu+IQTScsXWCzCJp/ESavRJA9FU07jIofhkGibmL6EiquRS
/HJH/zvfGinflrcTC425/1ltlImWeKST/Z3sztNV/3K+HZVPR3IwF9/zhI+ONg69
IeGjU8vIcT3lRPhWT8cr6Tx8iyhEt+pcYZPT37zffrZoj97bf1SQCf6hcPdruSbe
h5mqs/ci8zt+ZdJEOHKyy0v1TBL4dBJqWBHWN0SvW/ilUu+BeLzXukeLXlNXCN+l
RcY3beKXqyIscF3KgyNbEeln0N/6NYwE91zzM80UCgiWtdIOVIflyxHkhZnhB6Fe
lKCidcVePu084X1S5ZfCjnNpUgNMa94kaxrytQBNeSlq5k2dgJsbww+eDMeiLks/
33S1UT2ryU7yTJd+LdWsnQBAe+SDUYngNwOytpyMuB5UDFl0ZB704v9LrbHeXxXc
90py7kHTXAq6Y70yW0NhO+ev2ztyk8MwsdmFDh13l1uyphRhfdf8hiwAftG253ja
Frl3Peq/xdHVph3f/3fuLaC4d+Oz3D/yIJ9D/hmMIM2WCgW435RXHgz6gRm1FGz0
WcADrLNj3rshGz3CoNzFj9EbolRdZFNJ1gqbB10gbuA0dfMXHBVvLuNP1KgLX87L
a2vcNxxyaWK/SZ0f+gHhtmc4iZaHklmen941T3VIl55GYu2cekU+WV/c7n2g81jb
JvXLpyOLj22oNDPz8eVK+nLc8+H2V/ecXohqbnUGdjumv3EOYJ7pmBQvHNh6pDva
c54KRG5XH4JYX3GLqXf2dMpA0fHOGVf5vYOGnOKbMHrlCqIYTm6VPWUqPBU4/xho
hGWLCJfV0GVXnn3LOMHKKsNwDKtlnKa8in3+snFue5Dz8fXcucNHngxNO/VxsqB2
ezoukDsdAlA8pS99Hsuw4tpjkTSS9XN/9WNPNfKQmnyABa6jI6hgtv0ZjvxQ2BAF
vXYvxwIrO4S478aOVZNtoPGdOj7Rw3Ai/Unn5aFQzEUBth5PIp2h0VH8HrEO3ooM
UANW4TSGArEnqv6DPOi/9dYtqFftS0EjsZA6hdMl0u/psUk0OV0rEorwvA6Hkyu6
PQ7BXQq8fGyqKIob21B7vGZUg2wHO4XhSFGZI4O5U2B9WddAfSAuvG2RvttLj3AQ
t5ea7GCSyWJAUtp9m2Ol4x48P/Mny9PylnWJYdwQVurPEeRmmAqW3VicGMQDYRbX
S314bnB6JSv64LgiNo69HHpl6czxTJwGIFx5ry/cX4ybr4JagX18FnHKEdOrMkl1
wNwKXBrxpzjoEFKmI/SLEV2BQ6NIE3+k6IrjT6sNcqhFWNWNAVEkcIBuDzuVO+mX
/p3HzgKczXlL2frUM/NH9SgaczpKrhr50/RTrmgAspWcJDE0rW3j4bGMbf7jysKp
snhJ654heCMZhC7+3X/6HWq3FImlp1BDu5yaEoICcw2BIz+GtjXz8l9KpsWIwqiR
Kdz+4VfeDOMY7YKUeoWTHocbdNpShjeCYOpoVSnQu8z/2qFPuRLcvAc0tVN4HDb5
Wdm77Aw0TOuagtddayGfD5pOt9Mij42ylVlVl1ILbmOZ+LdrJSh3UxdI17TsKXtm
YPZirEKHxcFLchDwGU7ayenff+YDemtnZGx/ZC5KO0q1rBOGME46l8Ithp3xUz3e
4HubcNbWa/W6dxKc38pAzOMK2LYOEN+5YkqSUrw+tSsAD1mlmhIBDujN3gfmop3a
AreHi8p2qLjI13lFc6dvJpMm5vhGxy/TpoBtRS1oB3NgXwK6gLTZ9IMD3YPd5qvr
E1oxXkDq32067SIb8UmsQGJtWp3V3C1Cn/6+Pair0fCQSZgKHLnXjIJ6+MDeeOMI
kw6mmDyCWOmuwB7nZ3OlsoqhysoBkfXrfnLN8Z4+IO9daG/43lEfPpuRkgyF8LRJ
W4LOecrrk53pXGSjzZVkFAyjoX/1KC94zDmSckgT6D8HQiFzgwJyvzXrMHK0ufXk
QB29qP/2dBSG59bhzFG5lVPbqyi22IXWWh/cFl2LNjjbDYnsOqjOYoC4ATf6C7Md
L6Y1ka+PpIE4zTz4lPEIf+uitWcNjqRp/YqRCoHrlCGo7pzirs5HwFsBibFKo2Zo
dmy/Cf0GMd9oWwlb8Nkyo0BVDzCglbQFI5zpL9eUkbBHXuvhJ59jtLFElntXjlBH
qToogApD65m3+RrtHocaSK1Tdbdqonn/fhjfDGpm3ENo8LgFl3jORhbidj4JptM3
i8NmR9b22gLu6TIE1inQna7JUHdgH6gCBAhqgv4iJ//8tRw9ZN8YIpV7cLRXPNjm
PT35ifV2M7V17fkqmFOdgCZJ0Sxu7AkKETn8dpMHEGJKmjxLK8H1qfVC55YY7fgU
+PQKOS2GXca8KKU/wU7bYywndnC74oVLGqbmkL77DUeA2Bx8bL4c9whhGCFGiVt+
WpoTU8EYVSxWwCggh4Ood8b07fmwOzVC2MP8OG9vVlUFBxF6wPONy2Hdgu/MlvI8
KTV8GGwnyYE1uFRxtBIjYDTGpPHHoYlZm1qASvaPczEc7gAbbdVw9+U3W2cv8LeC
/4gnUWYwYlPiMvIYwyBOQi5Ym3Gjh43Rj0NJZC5B/zw64tTC3XEMLNw5ifRh648k
0BR/FXXfSeg6SYFz6ztyzwsx0nzRL9Mn0MdMSnpLqhH3ONTgdFD0Oem/ktrJDgRH
4Os40xVcuEF4V9ITT93j5YboWJ0OZdKZrjx3RIjmCMzFjw1HecybvTVk1HHDtsgU
4B9fPZdUwFeu37RLR0MkNXOgJgVl/2AetSbpEu2MsyVqyCANXsahs5bNEXOkzJKX
/Zq/7P7hEp+BtEjCd1Nlj/XWAZOvDpVtE8OzegMd0/GVfiUFkcX9d68XqiR61Qnt
lBsAFm5H+/091KzgrzQfPU9jZay8vrT5ANZZKIyhyYacE9waKltIboopqOrEwh1I
wKUiSjoAy8XOOFovxIWBmk5rFpPzIkrEZUkryaTDeSPpUOyHMYaoX9GX9Z2xjUt8
ySEiu3TCa0mYJ6A3dG/Px8tEJ5cQ84EzPjt3jXfFjp8zxX7NT0tgYvS4n/JithVK
bTxjUp0sSu07xBP0QP6xmt+PyD/3yvu424LEhyNWQVaPctXOKR7PljDEb2tuzRqZ
ec3nCHph66aYodDWMPEtT0R+/iifQ6h9YqnMI29LQSgcI5HUURssJmD8jPNiAPpX
2Rr622zVMpiGSkfY5E4hDUzPJVvmcH0pPFAjqeA7xso6UaNz5wJW/TuHpe7THNOw
6ntcFET4Pg7qQ+yWlTvZRyp9ZejNyzAL+MYygX8ouEg5isRHGhkVfQd4lEWqjUJA
wfPZguIs/f2A5O1bG0EwPW+jTfwBh65VzKzv98XGzWAKDK2YcKHKeCbkrqO3C3MY
IDf3uOG8l3/SOe6DxeWmk+S/W95ZDyIw7gKuG7Kr8RT7e59IfNuimR7yyetX8rco
PT2xbD14FqYyaiSo5T4jMafcQga2pNMxAFSHuTka9Dr8fFo8PbCup+hr190MuqH0
viKENt0CuBrq9jNuJF0XycunuFT0LXFQxClXbbIJHCp5wTtIXr99G2xgXDJ4GdUc
Co/rG7wc+Pmb2nfH/IPegxK6fvrRFfAMZa6a9wFQy72RdxTBhKVjxDzG01KncBUw
Fyc1UmRkLuSi3/jwoaLMRbRLodaH0OQAWwXn8feAzZV1RBDYP1tm91B3jyeWsw0p
raIz53rIodQePdFZHzaaAias2wxUXPD7bDBFnYKfEkAl6U5SahTVygXvLn0Ay6UU
06l58qVY67U6rg/UNXJhbCJLMJii3VDFP6ubz5SmQ+7EWOMESUWaQDh6UbW4JMg4
wL1K80oFk3Vf5juLgbM41nc4xSjbGQ+xaHwFewISHD7dOEQxBcVrHsyRYUwMNl0T
t0veTWBwuF5qfgf7+/8auhf7r8jqQDVViWC1Rq98pbJsTgVLbfyk8H1SbHmmYovl
aXLiP13nCgCwDpSTaGMkG+VIIP5/mP2yWuM7x1zQwo88FwuUc5Xc1rg8eqYVIWSn
r2MrEHZ4Rbg+PaRbLx1bA3q47XVu3EDA8VyHmuGDK26SRHLxdormY3IYwMwp41pL
KaMbpJs/J0OdTnnwSGjEhvcekfBQM7I2fbXINqlH5sykexPOeZOc34daxGArMcqB
Rvzb843O4qKcBf/t0exUBNKsZwrfD/gGSX8laMF2bcApm+SY8G52kqAP/GNK+Nfl
aKKGHOvhkmv0Eznix0oWh06xI1m2AI1n0rJdaS0u/jCGRo6QzQLqvo15Tdl1z5km
UsEixxM1nGp04rFY7AdokpgNZR6qhHTwgE8bGY0f2HpeL57Om/NKX7eXr6T5yV7V
uyLD8VxojPYAEsT/z0T2AZkee2ibFlzuugDE4Ge7EY1z+POUM4UOB7DS0cypZWKq
t8QnOr1vsUcNzXGyV+wq4XiLkDSR5x0C02nPYA1lWQc2S+TrAWug2BPvxLRhv1hS
XuN6F2/jDS4RicjxpHKygecbNkIL6aHZ4MpjDmlLcxvjIFD5wYKtDMZ5500hMXTg
75yfn/KmzcpX5vXc/vTVsHD3hWo83doLV9aPXH4XNmBD3AXEEWB0ZEVdtdZuR0Jz
QEyoDxP6kttXsd/50rtybLJpFaNZGRNgwJGEU95lVZnG+TiT1Yy6xQ8kCx+MmlmC
nk3INCstoDEHjqsvOvy2fvOq82E4b8Hwv8M46azUHVN8mRISv5GN6SzgJ95hx2c3
dBlku++owrga7B1LJaf87Klq1nHxkAdKacWy9vgXGOlg0Yj1sethLptInCJZ497u
eKbJaNymkOZGXV1y2madWPrL8Z7R1qxAuSDLuCj4DEaGIqw/GNyqINVvDkKyH46m
7JmbYv0CdPDGtp0R2FCg0X1ktBg8z1chcrWXVZi+Gu2CkWfcVJhGsqkmp2WBx9Cs
RLcfk0wtjRdRWiNnt4GJBSdkwIb1iyHQxb/iLomRzFrrIlzESxiSwLtVwqOF63Hq
RiUSQahtMSYy2khcB00HqFdA6xdw4Dgwl/5+lnUqCgOEJGnDDXnh7fctk6H+5hd9
Eiah8WMYqZC0gxCJWZ9VC0h4nXd6PlHzqGv9wR1KX261QcWHiuM3gORm5oESSZ9O
SljEFPP0h1BzQXBunfVbsXJSDe9UuVemfAmqQjxGujf3yR4au4VRIMZYarPuJKKq
NvtlaT1EkphPhEspUm1UKc6N75++PRzxLTq0T6tHj1qaqKTbpQxIYO0Tv0KawRMo
oTPHhTXSmsIhwi3QsAukCj1I/HEGo31cEl4Upp8XGrGOkpiM1fwsERxuA3slZfQd
S/t9aOYA+vvGSthO1lKxKDZD1tNp4dCE2ey+4rRP2BlhZMUGFTLI6RoDD+xG33Ck
Rj5+gakmjReB/mIT6qdIl1oYkHzQ4iem1+i66FkuJWnHkQ4Z2w3kdiWYwY6LtHpe
EcWgS6YpDs80m9SLOZvl1JwKtc0rgsQ7qP+SECfUaVdJJB5ZCkQVnnEsoLsWN286
I8tm/e9ekcAAOJOxFUCkI+pCNXuRCC3unVI4XfkcZYUcFnNKErc33K6LIEtG/JbK
5aZD+AZSAuh1UHHJum0mZ+VRNnbifxNkKeKWiP0IVRdn0Kw4RS3S+Z1HsPnZ6KRd
De3g7SiDFLih1BJe8Kwg8252sFo3GOHLYHcwZyBTEHRKDJRifSTmn6PHZEPQYx61
FZ4amKpnO2vvWHMUCNor/5mAkt3UmS9zBQph8fp03XenmjcbhiixFR3H/T8DjbHo
+zvjgDwC5213Nql4IxfIRhMnsh9EdZcR8hWK7fTxcteZxMErklGDYhBj/FuBnmT9
i+ygAs1+rm/y0/MtC234W8UrR66OcKr9HSbF/B8U7K88T1tmMzh7WeIZ29js162F
LRVFXtS49DIFXvy+obmAwie1hFdPqYP4iJJ7TG+Mtg+GKkEcCDxDgOw+4L/2Ek8y
PJ2o0sq+iSRRJfQiAHUCJnIyMUxEq22k5qtftnGMXiNifYEQMpAhm3xi2fCQJSJx
SlpqVv0PQfWMfjaHgNzE/G16wISj3y51gKs5HoUj0rhIyBFJajBV/FSU5EYjuJ4O
IrY8QZ0htDWoNW5l/okV5gwOnpdlxK0AEhyasU4Y2iK36M6VCL4TqCwHTn+4LCoH
sqs7vGN+GDEZorWXd6ncNAeYqKveGFsKPpZeI4ETsuBruNB302qX45o1XSJ3T5/a
S8xUUuXGzxhSNQCCd6AL7fNAbHSCYL+oYG7gDwftvLAsZFSua1me3YSlncsQmera
J20vT6bHSkpK1nJZ7zv8pt3Gl4eZTYIkcHdfCHAk1DsDxQI5QxY7gxl4kGj/Ca+q
g0CYkcj0bc0RK2f1+tuA+QABUTswEsxMBIZvubo30Fb0TRPb7R1ASSFEBZKhQRtU
piYGXYI7Urke5+abH69hx+6e3aOhPlAaXG8rVDgzgYLKSVvNl1tgJnq58cfazcnU
IUgSRKhe07xWDf0aG9gXZ/oSr0SLMs4+OpG78YKbz/xzoc0EwlhQZjQssjsI/QJn
e9HVw/Eu/thD2enqoJFqm8qP+VRt6uAkG6vRcme1XweJDYqaq8KtQrprm1kahGD/
vG0J9kawpZB6tHel5nbI5cnyHYaxOv98yFzSN9SzrOLiLmOSYarCwzKdZ/XUF4YI
02HGMfEKk+57o/ilhddBv2MI0OekqZB2a7vF5P/dWikuh7ZUs6pqYnj6JDmXRCx5
19qHGj5BbG4EOy9O6TtECoDQFynAkjLzJobtS1AAp06K0uvgPF62SUkjXgMxsxTe
m+/M+ZDTnQYzc41oDlq9FVTRr1TPQolKTP1TKacFINFEMms+VnF6SZqaPg3p7h7+
itnhyBY7hJikyetoYUqA8Bx0EsT7VnyUZZLWZF0K4qkMq5FSj6t0W+nV0NGjfKgR
Fo9TMudX+qpcPNlPnVfU5WKbLfEUXljF/VXHaE0X9YTpfj5fH5mUr3L7DBhIECDn
e2jCKfgpMObCM6W0yN6gcdIrJEKbUuFsyRtVsegvj4KOQ02XXcWvE27TMSgj7c/0
uLC0aXQ9s58pkyLY3wJ2o/tAxXAxr0QPToLuOaUOwidcsiJiHr3bcOmAeylErW+l
QERNklDFF0bEgNHmDCQOrfvf6384oGhvkymjaUEp/TO/d8SkyJ6A2xWnV3IO8ZWb
wfpixbO8NxEuc5/am4xQ58Ele3JcKwb/V3K+GLg4aEX+IkIWPcjkc1Se0EhU8sdb
RtIgxGHyW6oXV3lBQlmO58ffu+YZUFsN/EYlaiBSNaFLlGlrjFDONpl+Fpo6CjFI
FvI3yU1McvRnUFLC/ZCxGZm9/iOkIlTyZsVL79fiNu6VAtyBHfuqMZ733KqOmic0
zrZzhXmQr6EIxhD4ipySaHOwTlLqPV81lPGn6D6o30Q0EXc4zJTIdqP1xeAx+0/7
McCWY/vadgj5gBd7tSTWTypIY+b75mZ19I38lftG34Qnj6RIiN7YYxAksEO/hRxD
1pSVHjDajpQL/MuSOqcIBOMmd3VyR+vB3vWKfngwPWbNafv8Mx3NBbNoq1LSkn4J
WIeA6DoQ6eV59AAEBBh69/wsRMFqss2gYdjWsegTl/tEDNrXQfgIPvz9Laybzp6m
J4lbBeErTKKND/jP8R3uwAFQBlKusZp9xnOXlSbNlWu6E8vtZpmdVnHFKtvbpDsK
1WAH7ECwgak9Cp9fzvszb9Bw3ryWsD2wuqFiBiGrzmt0NUKRd8/d+VmEK9rTAs4t
6F/ESXHPJI0UqPiEMGOmcabP8m70xKR96Y0o37Wt505l38q0ZdhlzONEjsRLb2CX
wbLF555ukdWLWFPOFzN0hisEA0BAjgDUb2kEug+T13er2h3TgTMHLz0tMH1rMr4K
81lmIkUmush1nVKi+tRAgBhGWBBjFElsgAIXflks4zD6+0nMNSA4IwkExSMtIu6P
YCXcD24vUeGdB/xq2b4DhqsUUrx1Ozvyk1eBBIV2vaqvL9s8MLrCGxP6/IPBBe97
nWPsTqGWGoLfisqIYHsYJMlYS2UihPrnGX0rWGBqudM8sitWf8RvOP9M3eFcVyoO
FmZ2KCKxWkX5PfZKyW8zVKcPzdSgwZtFzJ8kiGNp3SBjAhqxU+U7ThzlR/VA7WdT
WZnftyLDyKTbJ2SsnCOAxkRoJ2IOBgl4rdYxuPRZ88FFaWT78zqji+pdI8IMGt3L
c8n60HQXg+9OVCu1E/BAy7NO0MxlZK1X07UK9lWFGZRQ0LkSnVAgPCS2zRG7ze+e
a07/OCJLGz4rlgD1F7ySJxBQzsopu1TuIHUNIOOuBr0uehQZVrUjOtcvUEl/99ak
cHkX03lJfEgQV/CiDoXClJgBq6QTQLUY39Y+6WHqDDqpuTVFjuEoHL81IvOHsnHK
VtxrBPbDfRWZh89Rx141YFX4c20y3SfaigsAlkJZijc4wmaMrnapm4Gd2zijoaVn
VjcA3h+/I1K0GAOcZzL32c4R0MzxpSvENl/ZLeGHeyCtQTBu769qudnk/ebHGT3x
oy39Z/082QX9vFbUeyrc+UJxAT4SF/LGpffa5ikKr5DqeJpByJuAyOc3MqhCjYNB
WQx7mDNaWWx8DlUueh5TT5LM28V6B+NrY0VB7PcEWXkW98oTkBvEuOuuNGjwBvr4
yvon0xpItcwQHZevkjO3J3L3pVASSo0TY3Er/IXoRs5PsylzBfEOfTOdQlgoPUOc
GXN93dyK8JDvF4yxB6+0geEJqKJNRTO1etuAgSFeGMKSOPJTcIO6SE7uLD7PwwTb
fyUC3xjv0Lq/2odVk2wrBZiyzEGDq1/kGzgd8JXHutr2ceRjWy+S9YZ09DZBhj+Y
v1AySFKhc2+hB9mEiT1GB0lQplYSHF/5kxRrvG3tYV0BjpADAPWRupRNRF/G+05u
58YWjljXT+WKm7+c1DpaVbwj4mvc1V/4NORJBwi5f31m5Db6plIcnsNTSHKFCaS2
kOG1KanitUzLx0a0W6kh00Lw94+aX5fU0qEBR/lIFmaIRPSlMeNUgmDYz+wuqhy2
xv/uSWXZjVLrUbMZbHfTarQ2dmMZDDvz3aUj02UguBXSURGroVMWUrDLBrqiG9eF
fc9JSrLs1I3gkIo2xgIV7AJ2UVHgQn4ZCvM18A4FPHeVvSnkMP4OIFW/MhBH7xsK
KNrDc/uBZ8GErCOOUNKdmgA+ItNKdKghEIeg8r9/D8wsKpidRuAWzkOcVZRHIP40
w0Eti+R/4671yrIUBDyU8KDI+PK/ReAsXu7wB6uLkgEfQ5zZPeZH8mr+Qrvdaqnp
mLMUI7Wi3wkCfcOZ0wKHRXLiVLIwK9ppEgBEQx34IchmeRI2Q7gnQK/ijRiU85iM
0p0B1e9j+kYRYftD4TBNqeQyFGd8XZVkV2wWyvJrJw4GLS5CHLtt7w4fglP778kf
jajPS3GwXvheyJmGWNWN7ELTP4DolkXHUTYmF5WrcLeS9nhmUV5QZOfc2S3JCUdi
BPBeP+vXxIsR0ve7IFTg5lhqOYHDzjAn7IhrCh7JMG0NErkerh2MARJ5LlCjQKRh
+j2hLlLwXOidO6pwqjpPTdce4T8tzkFSmjdvJBfJ+yiynbm0mrrbkArNkJAKeS0C
SW0zyDVQUMSORRG+XrLWBPl5cory9dKNA6tXBuwYODF+oWsRsonI8mKvTgyqpg5j
EcTrvyYufR0o4hwXOwM6TEZP8x48mYqVEnX8bEikOdSZn/3t/jFh0Ir07urxUwXV
10JCJeKW0XvFdJgkQfNDlxVRfNT6z+J/iZjXrzbsSnCe0886MSMyMAWwUTEomnY9
t2fnx+2HVV2vCY1Z8V2XDUxRuFF9X0Y1+E5DuU7sy5x17k2J7ZjY2MqxURA4qlOC
DBj7w48NerpHOQwI0Spc+lQSsE0/pZw+5O5z5m8nvSgH9BOWw73pYpvTsd89V4J1
E3+wnaaxTWbdEscvPGeDGYyciZqwkFvTc9ATAXmHbnazF2tpQ3zFpjHDCLW888hD
S3I5geHR+ZHI5Rbfzdv6s3FQNaV8Z8ZUoL866468e1Y/FiYcHSzJm1/1PcPhPM4A
W7NLUyTSQfqtqWMRUGknrfyHFxT4k/zWxtZiaVKBaEVgsZ87ClqcFSkSoaAQJ/Cl
7zys+iC0WVV/rFo4SErF7mz2+tKyH0dGOsUkWL3PEzZojVZxLYs5LwsOuKvBt1Cs
9nLjac+pUtQlKwEo0JNbGPjOFod4n26R3yvsJ16jY8hvG/QntagXCGsI+66jAt6+
iGW8U9zwnxI+rP4pfpjH+l8rbQh+mC4VubboYZZ4nSETq3P+jJ5b2RJ/ZluuNrnf
X2SSHIZpzOTeUT4Q0Rk/ygTPwSWZUj0TclBZsw9VZqef0hkBkqRVzIsakUO8DQsv
qnx4ekOKi1Ilm2+p2L8HVktZS04TvAhMcSt60e/6WYNRvP7fSeYOJb9f1SDfg3Pb
zErLJUa1AzG/T32TcLnTv4DJHZx1Z338hdVRh8OMDagf0CcjU3wv/yR2cDHhntwg
8A6sprmyeTuj5pi9Z9P2ocULXFfZtE4oCAg/YfHv/D3NnSzqE4nAt93cROJXMmph
lYmf7aQusWO51T+r+ofNLiPFRR4gaOp15t/P9hcVEMKkXl6RuM2Z4Fc8KnkuNMCf
lmLDA8D5ahXnQ40HRMktTs5aB2F4VzBjrDmX8NgmlchnXKbagWWt6vAj2w/GZQzh
TfcOIUVto0wTiIuHEbRD0zfrfqWm6ALxg9KGajjbTs09tWROXLjUGDHwR9Yl9DmO
F5svdvB7Ur+GMKF3bm/5sAXWgfE5f+4VLg2ip5ozdGTtlawYeyOoC6YbGcUdG+ml
oJuhcKfHl8Eq3w4v58PNs92cJRfmoGvpfVIKhpAsmP6uc9Fz0BEPHrsTBXOz2nFP
743mrEanv/lpsNlkTz7QL5OO+rdas/oFR7qSgvfT6R91SztiLyxMytWIvJGiOS7g
Cpj2DicjvM5kwxIpu9qcfA9qRZbq7hpiIgLqceK0d03iajSUYX1unSsg5K9GEjE6
Wi/ywNHCmawQnyTnjZMU9lWVcgbo5kMQrxNR/IBxhJLAhza8qL5CgVTMxIpAXRYq
jWwW/Hzq8QzhtN4mSm/Yz4l90ye5ow9myqB7RIQWzbLliOohd8G6gVi6mZPP4Z5y
RRDoXRlUqfmZdtAf1P9o5co72WiWGkSILJHmAXfl/mJV743e2eMw1xPxlAuJHI8C
zkw2J+uIlOO5MvwfY/mLyWp5BjVvx1RJe6kb9PJSmgarKOXXewjvOvPMz/DttGS+
PNFN+ghzp8nlBZsRbeJyHcxwLJjIe8WnMoylOJCyOiLmiO0/iAIabVe6LFOqZxC8
GTG2ldDiHfC5sMGwMUk+mQVMkYG/dodT0XwQj2ogln9p85Sy1bCXOCDEHRuu5EQq
bmfVy1GhzfbbhGOjlFdhTBCQHzhpBVQx/bG+D8Ob0CUWB/WMtfZMdI14Kwv4+Ch5
//Pxo2vO4ZkM96YdfgbGD20pzIlC91BH23xE+XlJ175xLwlE33noxwlF0E+vS50L
+IKVj0gOj7Q4AwAFhIuRF2WbEQDPhT1lX7v0O13hLmneDHGmxGHBycNROpeNFP+y
KgiY72IN+wISvwzwLCteVPxVoibwJAGulRH/AJYWsTpQr/sMqj9ggkJWtw0I+y0b
phi5+cx441m1boQXaB0vkB5xjI0sdsmzBjZ7jMAdXnJWz/sjlI/8U7Dp8qVYvPH2
hVxjYjrQh0PvU08PCfuSO4IsI6H5rtMYnjyGX5q6EgPVBIx74dDSFPIM5EC6xnuo
ehz6txQCC1Dk/8do4D8NuTXuG/aYar3lCsRID5C9ARrZtFeVH4tH24aAy8YABovh
SlWrL6anX4z3dre3T6Vg4pAul4gQmw1MLT6bfXPxWsRiMPnEU8wWaQHeHnAO+7Lx
eewnEs3GmEhGSn8mnDzn4u4r2QXfWQvdiCcKmIbM0YCWNNv39wY+2+W5BcrmBXvW
xvckeOpMeIOr4Dwp5/9pXy+LGBEZ0Jsqt7O4h5Bpg5zLBalPH+5epHVkbqWTyuqG
Z6aCDkKXOsTsI+VoPC60Bfb3xIvCbWxBAkXFhUqkodsC7IpSI3viy88I9e34OGcb
4GYRTbL+Kk4l3ELSN7L79VMH8mTVSdLr641thV4rx3/pfkU6TOvgMV8Vg6Rg9BV6
GzpcMwPPv7yAWBnEkyxAipcmkvSHbK/UJPhPd6C/w0ZsVu8ZRivqJFtFAPnM244p
xUkdrVAe1G0p03OryYmlNjMp68GSsgO0NnNkBtsVe2SmuT0qsSNYtCGsNscCcRC3
Piq+zASVvrpNgsgUBI99bab7TqF8BpBAnmlJWjMbFOHJr/ohzR4J4+x9zftQ78ZH
oo4D+t57W35Lp0rFt1i+tfvAspwl/KrgKmXn2OFVcFDD6ovFi5O4u3G4goewSF8/
mRVzLqumtW2oVex251CW2n8rPYrW+OAUXln2z9J4hZcuEXoJzxaCknzKBXVgrWxw
2RLyfcsoUqkIA8g1HzlZqnP4VJ4YuEktJOmP51C2WWhxTsSdmxzOWK2HRMMbit5L
JvWfBcn/ruksqbmqJFnLpS5GtEUswUujAET+sdIua/6eaE6FSllwePLhsp7sYwdy
c+yxasdm9QIAxwX7IDa131w3rSrFNxJOaSpKZSMIxYpoGcax7+AVcafOLccUyoAl
lddDnTMf8FjsXkw6zOpfDZ+cL2gizyi1YKEE/fB4+90KqWC2sA3umAPxBwo4ebcj
5e8NER88kAYXS08jTgv8SkiOWarqj/9w4ykRt9kfzYIz4vh9yTtMr/0H8TuMW7UU
4YZuOv04UzcOuJD+Qglg8PjxSkDACghwCRlOdlbrfTcrY3NqaSppkXv1oTBkLqsn
3ECJUWrxjSV8Bksj1mB3Gc2rbda2lqnn2mAMJMYpuqnChj6M8yUFuR/B6ca1bXBw
vKW4P0rNk/5zQuZqWa0+I2aP57tWDKznJWj4IhHoCOE2jn4P2FI/aVxfq5qcuUSM
3n/PJL+Hsv4rlQauEZloH3hZO3p4Q5cvm9dVEEaIf9n40vd/cEl9Ugv56Q49EeZl
mc3MJp4HQQtTWfw6S3HrlCOrb7RSodp8446hu1sPv/GyQvD/8JI22HwELSofeVJP
HS5QvVkInO8p2BmlfmvN3x6iU5jD4LYHOKP0zgPPUpYwCLnVTnMbLQzaqAPDCL+U
+TgSwoFoesmObD81F0A5YZNNWFiDV9FYb768KmzvEln2W6sjIAUu9aeXnO5wejgE
7jek7S4Y/7BeEjq8k75y4IfFyxhM5gDNe8o1NHBeqKS3M8ouyZk7GvfQbJPYR49J
nsDcwJChAGM+A95YxDGrB82xC1ZKPZdRgupw3fIP4vaaaTLAdQHvs/AENTmZ6Jf1
j5YV/RW0erjXC1agouIAGz1G1lomIvJl+s2TJ4CgmViwnepQqqNfXZBVSi9Gm9dM
3J5W32Z5y+dMQ0F+3mlhsoFzcQKChsZXfk9Ak9XGxA3zgaynYoPqI2ZpXqf8NB45
A/Hb178R8BI24yguplKQNa23jbS6nmU9kiz7UYVOii1yX1YOQBnjrT5KrBdkT4UE
P4BpTdLu/0wXXhOecT1kEvhQNICmp7SC82kT6/yvhSv3O2WZZHWhKnU8Cof9VWMw
SsHHNH6XYQBjtpOkg/drOfS8HWkwsAkIb/VrimMMlOsE8G/EZS1kWk6SOIk1YI08
0CdePjSsZ+J6t2nuja4TNXdQrWH96UoOAFwgv8y8x84i1mwJ0JaRlSoHus2g+0KS
XoefdsC6yXYYh7fLVnUglh/bggz2wtIYc1fO5UXS+M+twGDBmSpAcaEGsv5q6ruu
jljD3btFXOupQMaQOscBpWwng7TQoBCBz8UaT6Q1ry72S8Y2J80HmWFcqC5ehhHb
dzT8vpQGqPpvgPuz4UdlV/AmieMMo0wYh/MigZvYMhWWT+3rZSG/iwl0LD8Ohtr1
Rh8OmZxd5aWJ6LrjOfxqpXkynGFFOI3YxHCRWK+QOvN8j/9hahFkXt//+UJ4/+Wn
KH/3FHHcq6XAUmoAB2uzhHmPgSlYBBUkcR29ZV/TINySv+axndTlEHUbtp17IsHl
OXL1plYwxMMMzhnquHj2libxg5Ccmv9g//UYC82KRhrTEwJtRYq3H3Cc9msUOZjM
7mOv/I3TLEYvmmE6VJgZx9ocHstOKCZCrhQG/lLVNFdlDuzvQklyBYw2pGe2BfFr
91UYSjW4KN+N9j0BB0BGtGuqxlYCTHBvF4cxcw1kMpMWkGDjuXQmeKT2SAzN66Iu
TdDm9JK3hFbZGlQJoo8d33nIP2fTuL/c45/vMhyxwredBkjqoN2olmx6nPKTDc9T
XNOM3RfxuzFFt3YQwj8LKy23ZOV8EGgNPBJ5iRprE90hutorig4GXkDZzOj2mVlN
+h0BHllWk1xS8fYg2FCqEuXxhYIS2qhfKDmwlDjTVDp2e/zOCdEI2FTvCit4++qu
Uie3RrzUuI9GNORaksNSOz1/6ml8QrnjwW09ZBhy1mFo4OVarecCDS1L8ZVrpDny
Ql5EDcQeTb9ycj13/psCbABPu05EFAAlPvbM4H9JMl4hlGy7bltrlgn44ION6GTT
ypdxYLaoF0uer1KzQ2yLL0rWsIJ1cXzQKs4a3u3fY2NHc8LEv2CcSt7Vw/9WHYRy
xuuu3kITJjs+3UGehOzmAAjEU7cR/fBJUiV2m+8ENqUFXrz/yC9Y+jXIhwwleENC
/o9z3+eaP6fmwwmB+Rzl9rUK37NmBxFNjsr0Et5N54cBsBTab9mOw0pl2nZlazgy
eMKTDaPKYgLtjK+PBqpIqVqWpNj8S8gBG+BkDRgJr7uKGlkOzEZt1qZ2QTCBPdhl
6aR90ORSrKGjopk+X/pUMQhcwLsPqmW4TLqMg04vPzlSb5/6BN2NKKI8i3OqnXNu
W4GC2wvKke1zubF2mivNyZPRYAcBgV24H0QqojLLFkEoRAvJ75fjRWq5JKL/bQDY
efTRCyDDWsDni2TfRXCuVXTRwIjEpY3Ncr5BLea1qJg2C/Z2Gdp0VvQMDeT1U6Le
AbhgkuyqIWe8ny89TdojTBYSdSHEyQ0A3gxakQo2AhS8zr4Vol+aNzg49XU6FKbA
K5Det3JKd/19zqbXhc27/6WgyUIb8SCN18Ph5uqPkimtQDNTaGHDTs8P8ExQMFhD
g/6qqIzO5iwW9adgE9sEFJhJUm2XDNIFvVT5XX+I69/sn2KIH+UnEyfbqBxvGbRB
RvnyLRvUu+MR82xe2RYQgBYiCr9bsaExo2572ebL3htftHXUlYNAqG2AfP1bBDxN
SxctYoTvaZhl0710xr4fPYC5wY5enhMKhRm2RADrbw2uA3uYRKRXziczKJqEULXJ
o8v16dqmdgSnNaEyqpqRUGiQHzBo6NFPH1DsSAAy+iPyeTwK91RYQ4eqECVF/ikB
fLuHE1uIW3iKSarqfLCHL0LgtRyqkKLQ2pFtPRoCp/ZWVCJ3XUCWs/W+ZlrEWqJM
gQCEGDQCEoVFXqy8uTL7S9l+VWJltb+br8ajWr7sWFiylfzr7sbjT2WBusFxzARV
ZBMpxDrePy84aMhqmDWD+JZ6clXuCRla9qVRvO98mSt3OEfDXmPmTuhxDkecYUpk
Ir35H2hWV1ApmkiboA5RTb3i9gkwVuLrXuDy8zSFQrodiccRDeN/zep2Lz0BRl8I
hUAPT7h9tZchf9phTI45BlkHemHSG0OwOYdYlsV2quHetN75SDHLrkYVW3aG4rE2
H4+uTqDIqqcXIrG9iMdsLrrRfk8pnwTt+tABXB2suneMYijLgtHBpDZpf0D1/J/d
P1gkZR8zM7daqlfBt7ubefPQCWiLh6XPF37ZW8TlzY4GX6iA28mJNIU/7jFh1BiG
nohzB6ROtCE4tFBozLS5uN06GoD5b5EIehr5bd3sddNvq24GEvGyaON/2QPWAIQC
A8w1NLc65m27ZnqVJUAemNbhidIe5DaEzFnViiAqAj0kMvh9Vzwlo6lTqHr0lmpv
PLBpY17dDccBWiXqNDUgs3GkwzNsw8ROFAiQBl476xyv0RU8xbwdjbEDFRFjDvLR
CXYlBUz/CCM4GdLGEkH/jtqJ/p/QnIhJ2IvNEpI1J9A3O2QhGHmmLffOUz6jVxC+
0GTQwIL2JHclN7YRLcYytvVvFOZ8ctLx7UsBqmMZVbKwH47HIKuX9gjjOaXv0XtR
MYuW4mIaLVfoYIDkpobJfZW/UTw/aeH7v/tKEZ4HiuqhhdN1ZAvSmT33H636ha2D
lk3EdyFhqSjmdS/iSdsuiVva91gw+b0JS9Z+BFdVPLmw9JC96T260wVOMlOuuKja
LD9Y6tfwrLquA2hS9P0nzAy64Me1CpmGLx/D3XVwEYEnwN+mb8Y/NLDnx9lg8b/r
X5tPCKZI0u7Vsuutsxa6zXrqJdtxRwA2OYS/FrF+lpObG7Kj31bs4wbfRUuD0f3O
zEpzK1qB4P8y4NhUSaxCiwq82dGwCvYwSysuU/NvTTpFWXA6+Tr0ewiaoRrmoVCH
ZJV8zx9mwa7a71UR/GWIxqblDc0xJ7oF71H8QKRXWgBsntyHulG439mUcKqhXfqE
Xq/8zDPY13Yc7y/Tln0KrUCudGzlE2gVkO1TsSyZMMtIePQwTtRAo6yBLTWDfdPG
SMPnrMF/EJu+aJo6c2/pZ3JT2/GvsWU65LOadwjP0gI3T3BOZDJug1kh8nsi4lZE
asjeZLWHe2KBOOqsBjZ97LONCQ084go8PTBe5QrX8EWVJgFcXBHkGk526MhXsV9e
ma5KGtXg7nhIO3Ksqf7bOvx8+bm5Qu0xmursiqE4azcA8Q8jbMHHv6YJdECJzlCq
eOvTQQXl2/yYbl0uZ1Kzv9YPw69LIqbpt1LxXG97aGNmP39jhXKdha8Rs5nvMalH
zNaTDIy2a+ZkV5cSZt5OlfITx+olndwGzA/B3yUA8FUOB/cLFoEnBA/aWvEGs3Yh
ugDrGqhh/J2DldSHNcE/dX2hKF6nFWBXe3NNdWfwJpOeul+MXSGt02AAUbE8OoWS
CqcDTjXaxeUpFi/n1EB9txtaRsELknEjQPqzOFYPWQAn6IsXTI4n937JvEmfP+as
oxEphU0cQk/1koBSzA+r1mx92ukbCG2y4N9MooNSlwVuGoS/R8lUQlu4MZEOIvJq
KBQdEQol2/+Mdk+6Rot1N8mzNvJ6x6onzVjS1TJgPoWPqp4Ej7vYay3h6JWhV1FN
KdqlqcoGlKRMyOE0OkjBuzcx1K9jGA1c07MjHzTgd8H3YnrPV4ppBbUzYwg9RxYp
wlblsO9TDFwelSe+UXTjJozYdVGL5yXChO8/B5jBHyKA+cQOOnyLQ1fxppLEM5wg
syRC8Cp2pBdStSmLw1MensBiDgBqRCTv8s6Iz9tyQHNJuuLo2eoFpf2S+MFEPl9j
h+Ic3f/Ro3OqrcQMdhH51Yyc2kJeHBj17SfSyME5vymNTQFIEoAKuCdqE+fdkVi7
opA8zuJ49z7jNkg60U3lqysTPtlhed3GdxedzKsIQ8fqs+Z5KWuWwMRlvEA5bEWR
86kvmwp2R6ERjLydl9UiXWapT+OhJ9RDJrovQ1AjQAtPsmFySPO2byNb6vjRM81G
El2++48/xZMDf9TvBK7EcbuFNa2wmXkBRUNqqDooMYzhyw/UoeIjgsN+UJZchnpV
5EuG3D74XTTmL4BCpsPH9rCcCL4EPFlFlGKes/hc4RMMLAAinxHE+uV+X8pYHFu7
DXfYrpTGpqe0GlLr6ZVI8P8+31kpbyerr+JL5jIbKDPOd5IUv5GMHfZOCJFQHhwT
AcAG/bl75Bu1pWGC3EKovx0hv9tX5WDwMdv1NwzkqB4yj06k3W0PVNMEqcoW26XR
OIxUap81eiGOQ2iFFO4H0fe0rMUYWEPDUnRZdhw1LINJheOT7hh0Q1rj8euwtcai
quQPuw+3OXUsOiBpOLsvgmL7NJcEkNsVpRZNgv34wK01Dq+eTicrDRR9ZW1iyqKr
BPQUNWFDHfuURI2L5lWHRvKKRaE72Q2ahjcECSVn0tHoKTCWWp8+kVm5NqNZPQ27
NGZee410LSC0IVyvnQCrLNOBSZq94PMJV4Oj+2AwjWJ5pI06L0BC5OjhDk/aVWzw
L0eHezJwu+cN2tNT3yW7xC3PEOcqzgasJTygSRQMOgd4dUxwuz+ZngKojy5yhQdi
Qyh/y87TfhHJkHpjpela5IwzzBpe8ilj/wtbwWKsvCZjj1H+fWbto9B6SIgZBaqQ
ZzpuVQ3jYO7Hdwvavp2h0FTNdz/tNEIps/kxpfNEAuHYkUqIZzzPfmXdiiyR8mde
DTVea6QBEUI0J0aySAiIFxOLvOQ4AEly4JpkZx33Uv6yfOqjvZJ/iNW8dJYXZ68O
LCfX/hPooGk/uYtX0Il0i5wk05V92NdAyTq7MX3+ojKXd7yXQX4DagVMDQEt6iJM
2SCDSrKRTz8Zl2saC/vLb3y7K5KCVtUGMM9eQZgqKVECw604Fq5EDFJhDpi1tNHH
IkpSILMae4+9Xs4YpWca1nypjt1M7kgfuI7mBaCjvpeTPXr9I8rfSx8xkJvXKhir
AgRxye8RkEHvnJ1bX7reXSzOg/8R39Uq/hVQM/6yCQC6v9XWCcXOQS9PHKdQjJKy
RxAQS85Vh25PwNXIvhqAPgGaoD8fhCSQhXJH15RF7juhrZauYpMkskf5PcSsekmg
fAJCr46tyVueabWFZkNhNU8RjTRIBZoCq3aZP1kND0wPQStuzr/KE9pbv/smYiLw
Gjv07MJUJT9iMoLvtwBZBaTRuS2csoLSDQfiWHYYms0lD7kSExdQbCwQHuDIbX7V
sBAt9c1dfc1p0rGdmjRC+CDMc8CkywQhXBCXMVs9hyCUFwdDiPudKIEVNAENCNxk
rXM1QWR6JecuHoy4y6XyNDAeRTw0hwcXqtKa/o0XKnbryFQYqWOe0zMl84Ztaecz
LMbUg3/dGhdz0mi/az+fLalsYaIEcodRyQ45raXKH9OeKZe7YS72+KmSFGXbJ1aV
OZPA9IwEUmr29t16Yu97gJFTG1QCHJaxKpEgHHUhhHYwhpXUWnoq6tAhsminvQQ0
WB8m5w/fWM/oGfTq3hA1C/49lXdZBU3K2wbTVu5Qigam36Nu1QAURwZEyqoCCoK6
q6bhxLMXLAr1xwSlYSvUGm12KK2cMiunFH7XXW1Oe2BDwsfvRstthKg+Te9L4pXU
6+qZdvJ5Fs+rrh1NE6qPS1qFOUXeHPYDr1biqoM22UXY5FlRICnxAshobJqR+2aZ
Wm4Vrarko+5VlM7tTnoeAofgGKAz9maPQtq3hwupOqaxBDqkkXn/DN7x7+MYKVqb
pKX5eFrCoo0q1xSZYebMYIGQvAFZk8utAoDAXHHcibWKh4SyKWLLiV8FRwfrqmZl
X/PT2qJv7gbtYtH/FFxfQusOto2knZrJRqCUaCFVKres99b1qIGjYGHqmuWdp/ip
ZLK8YXrfPTN+m8kwCbmY9uGLsCP+qMzY5Gf+yp/POD31Zud3A5G+ZxSmJHShCX47
SHnOU7vAHM4rtI2DCnnnabefqcBhngKc1VdYWCJBUfPorF4Da3PzC75BbH8B8/hq
inHGT49J6e0+jIype1L5hBhrEKM5mwH/S8rzoGsQgA9o0ymD0AlRLQG5YYDWWEw7
JGlVBnT9oZ2gT2Nwlssy62GIEnzM1T5yci8aZzcyC2xjD3S6J9QskCxtXH7GxIZj
dAUv6Vf1votWTz/78bt8bmDMSt+Sx5pK+IXlOlFciacUzQHdYP/OhXwFbDueT+w9
Ccm2jDKoJ3ZIcw+rOnA4/aSsWzVoEoF6jxniU2s9zLSwleC4+kT22UNj6RlGRlUK
7t7gpAqCxha5UXv0cfhZex2lhfhOo7mzOEdWkAJsBg9ovsFueHk2jDIynBZC2HVo
FqdNfCs5pNJtew+ofly8xExYOCPla3aleYcA+5m+QWVlGKhOlx/r/9d4+/h28hn3
hXtguYSNyWcl+webxxTaaIE7HzckO+xj6MlJr9FLILAVXCgt+nyM+VC/VvpAaEQ8
+XNmiIA0oZjuTc4WoWyKTLBCKuLVLdmjJxEC7ocWnNXL7TFhfnwn4yYMuersVE3D
ugmuMl+v7M9RLS+Z4wEr27jNT2bSYF8Gs6SrbnbsBGvobki8+h2j5yLou28PbuIe
o1mfTSY3Pw9vjKbBMZ5SPIh6mw2G7G6xR6IqXz4n9q4Psh+bS2jtPV2f5SVWx+Qz
9djkxUL6TjNplRpp+YciNOjNTueh+U0r89mOkayC678TI4OQwyvBvSHLUNghpMKH
9hfeJ7ediONr1yRwemf0b/Oa6FgXECrhpT7WFFW5b2tSVUind/TdLgubTvpVDlmE
aU34mbqlji/7ZDITgA2t37T98slSNH9Kt5/RCAf2tM1gbRQ3OYnlREwMSX13g1yt
m36frJkrkfmA8BxRTJfkA3KngHk7WKf05OrRWd/3DZQdkJp7ACC3/GwVa8lFmo88
C6ZkNCPwvwWuAak1XXzTsJiC+FYA6SqNxfgBvLduh54zPxewYFlyFL17F7vOx/u2
BSmVl5RDXmghuHZr3Qjl+EnH+LzIvHvDOECwkLI2FHFmcCPNNesyLIBW3UuJ6drC
P/zbMFkAtp3ou+IlQw/8GN304rpXfHS5tB6Kr2m4runyirSYaDo2Aha9zRdEVjQx
d9Tvq1VUPP6Vbw+Dv8d9tzexzcqrvSdcVIWaWM/grvPbjPTjJPNDSpL5DRw19QHW
gIRQ8yRF3JSI1Z4RVtmM6NTpPaAt0aj94RpeQ/mEU3hWKNINpAZqcFXz4PJFHOju
eF9ynMfc3gmtLw+vVk+TA37BRNerV7CiNs9ZticGvjYrXqWQq0Wxex8iIdQQTi/g
SnrpYUITB7q6Wxoi14AWEoB1wWkKpxbbuxNQNyo4pB/2sBeRmd5kC95WRh6cRaob
TkoBxW/1np6a2HYM+IEQp8+hjr7zWHtIEE0XwJUhEe0vB+uIgOXeuKltZm3m8Csk
oxOKMWm1fbHjSA0gKctrbM0bDBDaPm8P8N4/Ey8o8wAAg7ILRzA+v+NMCLJSJht/
YjBlFTEqkb/VC4cOBMVVWjUuu6Kf+cXTD7YX40gIkt/K3OYFcuEllhgHPk/v2ZVg
BeKNIyuWyuB9nCwU7w2CcRfvDF8Oc9asxcjkwdEWUCTyFM2ANIlWdX8zPGaP8glH
tkU9CrsP6Q5n49zT64Dg68BTEXaKWIlBxy21WueuaYzpQiOiZQ5e2EqDnQolTW88
D1stxc3hcjAMfBMkZmGF3exqddQnbJqtgp2AtBXCetnStJ+T6G/PxZejXQxXQrte
7bYETALwn2g+TZD7OLNPBJPOwCiFSsYeFyKnWceY4x8yAuxOcaNx4Jb4oVzrbVPl
fbHfQwerv+wC9gSIlyzwGOMbwEsxeepAMnvbwW8v4N+5w3Yc7AYav9RC2xeJmFMd
W+tgI2+apALnsbHvcngUw4Ux+4NUBDoNGaT0g8MWweue0n7sEgvfBIRL4tbpUtjo
UNlkv3m5Lf8XiDJX0VvOmIq86rUvTWiIx/cnzh+WoDSxhg2/Ap/8qIJ3vxiKSFnX
t+o1SnFeGVrSwoiGJw/meyx7jca3o898by4ryfNWg1AoeutJAOFJOiRragNqz52j
WG1LYlYjvUJDTafWfm5YE77Mo7P/7fC1JxEqrd/mwa2KuFMnVcV4wAlDJ+2a15ah
X2XJ6QLqfB9pL/RNbK4MItO1RWBy8rC5qJWbHPBExVjEhGmvzMEU7aonESUwZTFy
/gnsXLyU5FIOsrDWQGMDZ3MSyxO9xjTxgaL27jlEJ9qDZP9XEMfSGgm6PdsHOBbg
NsF3iO1rlX95MsRmL0Q/57wAepCxjRsmg8TqTeYCeufpIwTi/9p6jpZQaeZ/y3As
JpxKDysgcQE1NSf3DSq79p+Iuo8s886A3/ZyxeVH2QzcMeRBL/TjDgXXeyOuoRs4
u7FNZQuzKMllXgyleP7rNsyrSqNCy++kvno3bU97jnCqnO+Uv0lUu4392c87UiO6
tRrwjZFox63ahFTMCldw3LBsNFfCx+ePXalYI51wAr3FzJJfIhzH5doLJimvfMuj
lTG0htddvH5HSQarUscpdufTASdQjF8DhQ4uX+kA7JB2ti48QDUe0vUgXOyjqnLw
QG8Kj6vnaxW1Dls+jGdfXw76TmhmU6XwoY5Tm2PwSsaNQgvKvfRsPl3xN4ifI+fp
HT+dSq5pmqMLfqRnaNrdTcHsKCAZlrnphJm1Ex8Ml0kOIhHO7/NQktme8e19+XOP
A1DhDBijFaE+3tdvVVXcfRZRbKF6cOLmnICI22U445Agk5g4cN/R60XkwacoCwvv
gUnHTYfcwh1CGau5QQxwdKKkJusuwW5DLlHvKMN+l1Ou2IgSTFKvNx25Q1d4CXVy
c1XnZSfzO1UHSKOKk9jggcr80fQDtfz3RqSYzL+Ic0sTUBi5qyO+SkZXhGrk68Cd
t8Or/h8Gz6W8rLaHy/OhpAN1FLOZjurT0psRwcHDyfOREHrxLCQqsXrWK/HDW9bf
0J0QDuPfOScDhJnDVm95sDfCRbfnvQEGDdJS98KAPd+Vd47wN7GNdL8JM5cvf+bZ
yU54qAb9eGHd6k304/b+kCRh4Gwv9DiwwxUCejWfCiRqTaDsaXieXNVrxJbqs5ym
Wq5wC/P43kPHu8yRSNcZ8CWBwAulatS6vtLaoVWUXkAvPwIx5fEa4K5115jcxOQk
RE04VoQsh27XupdEcaWfDKzN0h2QQ5GUq8chkJoMkbqhv3e6wXCgsaQDQ00K9wtM
ViqomVEsmlY/0OX2WCk8PM2Y30rBBzx6lcCBoD7oK1TsmGLtMG1p8aZB4yAjKODJ
0taNhlD2wwea6KtOTqa5tgvwaASlNxVE1BVTUDucN2c5gdvPo9K+thzCmCN1YZOb
6bjb/HxlT7Mpxg60osXhVzOjdhAlaXASSlCGIl/EBB/ReKfqw7e3nFPWu2uED3PC
Lc3Ge/ZEyi9TaQe0+e795TpbTC8SKNR558UdBFIYvR2BSdRLHb/VKw1tv3MY32zg
h2HV8uSDlgfh9pQjGkAsoL0/2M9NwKX9ZJdLLycBoDwibIcmV/fedBG+Y64B5Y91
K7nDppVAaUVMT4bbdP9E7Ku9pwQRvFMzt311UrXt/xP7KNuqHfTBtU7DfEPRmh8r
sdw49gc6SrY8FA1tklZK03859NhaShKr1dua++gEf/pCj3fv7oU8JjiaGm43PreE
G7RlHx2hWEY/Wgh5przGAuinJzjzc/3RbE+m1X9H5i2o73fDB10DuAlLgi+Glmv9
/sWA7fMnJKpQ2DCaw1R2bmFTbplu5iNZVpq+7gxAnT8/Qq2lCZMVojoNOig2MXPo
z5LxTydFzWeKHGBhZ50tkgBfmuOj3vp21oYZr7RtLi6hwHynIQqBsJLc/6XicSc5
E3aqomO3AUvqnNeshOdG7C5hgZYfHpmyRLCP06wF4uzeDR30Azx6PT6WN31aRNPz
HhucqdqZ8l2GfrKe0owWsRkgesBZBakksi00PA6Cp3tpaixcD/d9r8LBjrYZTp2Y
LBQy21VLmPm118vZDwXuOD1i4FUoxS7ZcUs95rhNPa8Y7W4lGwI6RgRcILwJgZMC
qRD0vfaWi0wvL0VFWALdVodFxsmPr66nq+KC3akklRPIuoGdMqp2Tn8Gkh0Lmp1m
g0nrKKyhccMP0SXGefONpf+cBzFKtV/06etOzzf0OEPFTJHlUTz/UBi+hHI9VENM
f21Z8QrVExgPh7kg0VTRqkE1sW+UsSTJaEOMdSJxLq8FHz/tz1xi3XTXFZ/O1B/d
kgnQjcyKouAJMn+DwIzzqDt3X1BoL+e8UmmcAzWbbwWMQbtou99ccx2SUg6hGHBf
XWHznafhdKR1k+2aBJ1i5WfFr7j9tCKUaSGxt551AByd3Y7P+zDPYpVCvr5xm6r8
Bg/TqvTao3EDHKrQ68CslZ+hXHMhPzzuLundGzohothFXfRm2Z/6TazL7N83Shlx
TExSIoCfcrPXs51649Mei2JDOCg0vRCCRVrqy5vMqTX/AiXxAqCd81prnOa9YyvZ
E2bU02YGRdsf72j6BOF5gAZvNtSDqtDNM2KpYd5hwmHLoZ/VyGLpfkWeVlLJhXgk
LxfjAvFy6mstuxWFQEeN3cyhpc3m0Nsq7rU8BWG0mSarpfcudEt3l/CUgZy1vg+i
YSUfp7ndT3oqXSmCNadAVwPVTnzhpqt3e8gXhXQnSx5R5pmCsf1Autp1mBS7Cwxm
GODwkO4vFrQ0rJw32V2562f8OGjRMRrCfXoKy6lSXQA67K00rIsku5tHETO+/uxv
7fgkvi4eF73tmLn12fFz7MfiuCfJGW8CGxz/v/5d+FApXb+Wz+JtgwmrSUNQGKsQ
Adz7xBw8WZnn2oq/5y3BC+688S1pBBRQoTIpx+8cUJ4zarXe2E3Ju3InsJr2yyAV
txgPS/gNfmLpeIXgtSOPaBFC823NxaDASgQeYCx8OPgOIwyD/sPbMIxqafGMqtug
2VnFdNF9Ui+qztoC2h2vC+97AcXJlg5PfEB3zBYVuab+/Jw9fZlkK4wh95OODkl+
+gAGOFnqu7kGNXZaSnjY5p6vEEqX5q2NqhrZwzSIdOQwH63AYI6OiqEcQxKiimIh
/hoewApUbH1lS0jpxpxAduJ2g0Dyepah0lGYe7ysz28STUwWP91RfjrcIsFKf4DK
W3mC4f0/AFNGZed0pzzCbgOQ922DDJZyBpEz9V8b5cXMIh87Qv78bmYSlTRghR/G
ypsK0i9B6z5f5WvjDLo3h2YXVaMF08DKu54Z2tJnXZwwbxy8OyjfDF6O1RK7jFJ7
XGAcaB39hmzwYBUCBtNDdgiEO8Bf/auAcknIaPkIM40JYqXaxujNsmM2buFhR3Dq
58ZMdfS4+d0k+yFPnhLD4zDDsqxE8AENVwCNOdsC+tlilL1b4vTFCgFNNc6tfpEk
iypCml0sh2dtaFWQ1SLpkpXhGQ544qknTZbPO6vFI2uZCSqPW8HNdm8C6t5asUtN
oDFRncun8KpC0drhDeMzRn2HmEOv1VmTBzuJQjaLRwsrRNQCoGkxEprjP/vU0126
ZgCMXC9Q9El4DpAYx2UxzYckr7XtwZaTF+RYt0Ki2kOys03YVJHfpAlhqfNBSP6P
pHclSlJ2NjYEQ+YAmv8mPKEy4e/lKZmiAe5oCuBSHKugWPyi8Cx2AOkej1ozJMU2
gm3dun7NP/5smbNUdIty0JyxMDw21JBbF0fcyDRdsl1U3qaI/MlP5WTwp4LqpP/K
3f6hvgYZd1IOPVkN8ys8L/BbaPAAgEFA5k+c5L0x55HDIjJkgVa/5+UPqzNhCGcP
R3vBquMCllVJgzjux6DyOJLdlIxxY8sgAxaQMewTl073z7DpwpJgdhNKv7qvWBOn
BR4LsoQFRsyGRrid4WE2n9BRqI2PSMkYUECqm4qNTYvQpS8nBPE7bWpZLB1zKT7N
ir7K6loam3iw6Kpo8RCSypCDgJI8kUAdwmVRvP8kC6LvQOx0aQhyzv5fAYX6oESh
7fLQPXs14VB61KC4ZSMaOjFIOBGl6288EZaWCOcDFAelKAOKt9uIPDuwjnhXL7uN
ql6L3QGYGKLKbM9h9ea3hFc5Jg+oD7p7EjSDs23s5v9+CdVFi6Paw5zNah90jNsP
bJxlIZkF0V+b51/B22reoYOwLBMAz5CVLVgp3xbwOmCC/8RStH31wjpBZMzZlZxd
H4mgBMnnlJjFrIlE5zyGgLLWNiH8l4TcOCC0+kut3247Zo6WofNgUdGXas0PuS97
rMe9uR5BxEJYl/WSd2Db5e/CbAn09IQtivMJaFxVXXcpktFNTN2AaZ7opcXBU1FG
ToCm07LFhHBJf0ddAxBbN7ShdnGuQYaQ9Xgh0HSIfOT5lT5W9fh6+y7EXf+wI3MM
QizXwZPGiIxppmfx+gwe8KlrGdaDIZiHmBCjeNbiBxiBPe14mq+aI5iHXwYSFBE/
8n7XUaC6jkvN36q8MdhqrvvMAlWn1OkSEiS21egbFMtDIBDNk1PJGZt0A9xOlX4A
NcdILTWXaxmANSaWe8brg/rh9GkwemOUGHHoLqs7c2oa0cxfMD2eLJ4Po4TbBRZW
6dyoqo5uPMe5bT2NAKzDIsKSmqx/Hq1SpZ1UFr5h6eZFNC/XDT6Evr65QWT85ysm
fAATgRh2UY6W77DR4PWtX1FQc+uRkL8WmPb1nJoW6pvOrkPrNO1Srz1Xr8jkCrqr
LUcHWOO+zFkCyF0Ao/3PgGMdGU0SEI6CL/t5KUvmxmCenSRBNV4ssgBtEi9qqCfQ
1HK9lF4uJ6MvG6b0Slo7/UWmXMP3IkUCFcYQoVkPtyIMz6AsI4Yu7Ql1ZP+jqsvV
2TNFp1Xqf5mOZZp48nwLKFMuMGfLWY29wa5GxlrbMKTVhnl1w5JQFtxixkElPIAx
4x2Jkq9G/v8p3UZYooBmJ2FaQUnCyCueYMGjJyJi4OdkUuz/tEf65yiHTM0wS5Wc
lfnTMAY9lfP5es05PGnEnV2bE4NLZZXS0sXvFJqdOLIBDgCb9QTvRvLzKe1/puDd
Fn6Y09dhkry7SPpi8AFUdGPeCix6ge86rlUeIDU0B2K0yvaC6IxpSvqvuXpAyLw5
GQ5093+jwVMWEgjATXCsAi5jgG7AjsjROI9C2irxohoBxFCRIN/vsU9Roteqv2OG
jXn0JoD1519KU55pXkCODuOdmE+uDmFKujRjVpHq1I2WY8GaPwpJB7YfnC1NrviC
TJjUZy2WUXjG3eBdBOxv8CMzPoPFHWFAzseG7tonLiK8OdXZN6p5oIWQXfPHU0mH
fdocw5T2OK16ZssIFaI5B111yECF/P6PsVsxYil0aG/upuxFRPJ7zbtESjljU0RZ
sbnpuheiSsWyTUXCYmk0LBXgXFsmGO+5Lm/JP/sjxp8xLH5D7KSyrlfKxVifU9Jj
GhNGQhTXxxLlLWcZyITJuBoFvJdQWrS8X/dft+8+7vNutkUyaRmAOgLOeKp+gRPd
byIBrjgUvKxb9p8ue3GVog/q/ke0Wseb+rN+kBrQ9h7ROboNimEk71xy0ki80MMY
WgLJYEE1Paf/4VQvBsQM+LfNL+fS3ZthizEaorukw30qxzTLMHOA6Da+EhOWWAgv
FxLMFckuKGidAEfYhiseFMkJKHjwPSgtIQxI82fEPdtLpq4bAT7K7idvZSbe7PnD
YKfe5xoO0HHSaw4wv5jdZXqcCRAqOJ8GZe9Js5peGLRDdefgghzxsB54MCwXbVc1
MfpeoNzgQQ5BFB9TNW8PVrIpk6tMm6/7ucRqWONmF4328EMQru6btlTIWYkppYgz
vFG4gM23nySAR8uL+2dODtMO7CuOyaMyFa8Eicc4gcndWZfswEMzG1H+ubOkMYHj
7Hj4g83fcN7rliOZwUNAL1fGRAM9QZQyJSg8wZd4avyVzT5it0jYE1xb2Owt8alE
Stn1UuWb29Dhi5AMSWW7eWKyYjX1DHkOhymQ3LsGyKMUcyOonsp5wKv+6jRVL6d5
Oj7+MVB9OAAoN2sr/amd+iDCsF3MZJgsCn9gYNGAVSZ4051RzbfEw4UUcKkaJ13m
JeLr0YK/xgjVYMU/nM16P+L5QnFXXmEM8RXW4ybdt77Z2vEuY4T5LDd8T9TGG8TI
l0JeTkxd2XTR9ftLR3qbfX4VDnY+kZSfKoMDN59i3LbVAZqmCQpgTB6ywiN9ePmg
rJ7f43BvReFlbblRpR+P7Jc0SxQrGPvAs5Z71/xi+553IjGB3ONo3SmG+TylSHTP
AZHXpve1khh7/qbhgYfom5csKxy4ob0GkrGKn0OlXr+xRL9D7OAfjBB13FsErtkQ
YEh1vVRD4SrbO8Ycs+R9mtOwr/VHnvxDhHCRVtf2yf18EQir5boE+AL12n8NcyLS
CzL/0+D5rKNR7ktNSXQHOHSblDG2W7mCR+kzADdEYWuj7ajI6jQ2kRNwnmVD7kW2
+L8pf26YHnVPLGQBCinpr2HNK9fWhTBeJMeRTfkc+wQ5ZA0+Tb+yld7JYpYm/ebM
pftMMyDSEDVx5gckK1lxbLVnLbnZpgwb31MJKB+qzVWU1Grza+XVtGZ4fzqGGhN1
f3499p3cvjN4b7sU0HGvLV9DZZVdJ62/Ouaa2pS7OwLn+0QC2hbYKngbNR71zcqN
v65JUACEsB83EbVo7n0H1YrOJkTtzF3aicPHc+2odb+wp9VYTOr4H4f/EqsoqEO2
h6l0w7pLepp3TWxwMQUKWJWJmYscZAAa+CRfLDXuiCBAzY7qEwZlflMXu5X15YaR
OplXjybKhRYibpH+9xdoqKEfeHU+1bB2q7dz0BhscgXFXnYyMyse6KPYD5jOXUqx
jXvFOmc572JpUPBpLOiZpM9hkXTjgnHDvCTY6L5mNraKwo/HW7alufECAO6nCIwK
jx4rYKc6PG4zMlFJUakAnkKB5d86WOKP4oIQyLKMmh2VP5eoWhNdIgWJj+eCRoO8
nZ81NQUhZEJGktKCdgiopDGk3XUb5UOpfQf4uEkW1a9SG7zViyAYHA7dqNVui5sg
+YBHGv6Lph6fvTpr3OXXE20z5KynRbB0SZzInFsRmCMeqfCHDS1khwX1antdmSza
4dih7fuHr1C8UahL2PL1HwkXbTwpTndwsSsxJqFACNtKI0rwp6FSTYWKSflxdEy7
LQmGQ0NHdTvgNx3hwa/4kqKk89CGMZc+Y40kfOGqxLwFdLA9LNRPdmBJsEjpl9T+
N2CTPpR+qv2VSQUb3LSmDKFWONVulwNCMmbxsEf5CrpQhD1bQkg87qZptcbnqlR0
QkgM6SubzUAxAu+k+V+Fk4BijTZJCgMDq+2k+ffWy38uvZckMMcGoX1rr+xqiZR4
xbY6NRsvwuCYJCsn6JAn/KA5FPCDAX1d0cQ23PIRmu0R62jXlwO75j7kerek7J8I
yr8X2FPkk4zOkSGlpU0JmevcgwTdVP3yXwGyn7xC64g8Z8/8P4v5r+yeI3AstuHU
B/AMoi+AFLKNXFIjUhIfoEZIgKee3ojecJwAeTp7QKz6qHpu4DgAZWrE4iYnhXD4
5ywwNkq0m3b1xZBfXkkZzao66z1PT9GJ7S5xiYZfBA0JCumWo/dn6Uf3YMiXhj8N
8vs1qjlgpAxYVFXhwzXGeWI9HGCi7m4G2L91dUoiQgQbavWSl9ynYQ6Jaf6oxj2y
56D6hm2lRxbc5qj2XDBYZA4k89kW3sjV559ozzM6SLv/Jm/TkjCQrcuLG7rPP0vH
Ax7m0icte817qim8hDhaho6ThfNJ5Y9g0JXiY1xoudBppbDVGN181/WTxAFA9TYR
Datrw9aSamWlzh/uuV7WTw1gzE1L5xTn/5ZdbRV5/XpoOeGIKur4ReL3jm0DKyXO
Is2hH1ndY4EXf6xNUwlnJgjbNW3Fy0ky7joO2Zdo/NRGijvNgErVRLaq2XezIxEf
QasNazn9NTpY39+o8iMRLZIttziRtolakICAz+/wU3pvPoWFzE90SuhKKrO1LDB3
5oqSXBnTwfks9qiLtM+WhTXw9etCieM7b90lzebeON7BIrH+z3DcEt/Vs/wJE4Qa
fzFw0wdswyhKjByaFwRqek60syZ1yFL0TxVqoGthA23Cd0xgudoHMYy8VL+LTRKW
2enJLXPkWudUTvU5KiiOcafoEsCX+Jcs0n5Bmdfc+8hum8rU+6n7+mv0B5/zeAYF
59hwHCBBo2WZN1Y72ti6Zvd2osOq71SgrDmB8z/KhAzcC0990wEr5QfQ6pf8v40y
AzQrSoXYRT+S4cKz1c+o3sSxLeVTGOVEwrSsST8OADnoIwHBydWHmUQrYT8xEIZx
zGGG8OISU0lFGkaOzsnlTEUET2bNzWDbTxK2+o2pnmsUe5/BNhYQl4Q9y5Uhxi+y
3DjZ5UVQk4r7iMn+4SAbi2iQ1MOmtWOYn1la+xZzdL5iWI1oW1M/8wwMU7naAAQg
bnq1TAcIrSodzz1zakzT140jBShwEoa1h2wjUPvu2OgIToqXVTZJ63eWygfWPtYn
0bpKWvLv6+noFmrM6L1jMhioMaAwgQ2UO5AXVOLlNUA5DL6FBZ0MKWoFuEiBJ5zO
f2I2IhyhosHLl044KVVc/Zdp5InhVW2jd7up5EkaBvTii8OVGfu/A3ljmi+qXqFr
pFvurUfuOLWIy1a2YiZaUVm8jf0szwXeNZvPhhITu/oESYvrvfN/7oSSqHrnngok
TuU/fF04x+jwKSRY6oVuxzdZtQCx3Ec5d4XI7C7mppXsTKrHzxJjDPbvBsrkhIGt
+Q8YKvog2iFjda1xsCciSttrhWKU1xezfhvzlF7D1Y8k+biDB6/LGqZ+EIMxXzFr
skKrlaEFpyrzV9BhldtfJxFkCrKpVH1E6z7y4ZEr0TNgnb0XP+XHzlW7chIUzciv
L0LQ0MfuzNmrktaOGXeBr+pb6u4830nKosltex4wDMHe+3VAmsYcnq+bsXErfjAM
WtWELtvkbjnQPOyATJeCssI+FJaSV0fphz4eo6OCwvM3CbK//TOSKd5wS7KOHqWH
WJcILakMPQiy01nBnvzKsaf1s3fJN8xlmTUjVx7Jeq9kB1AtFh6ASOKXkw4SvDml
r2UhJoINdnf4sobMMRqWTGxlnbu1/koZ7KoHyRNTSNjIcO+71iMDm0x3sd9uP73X
uel0kWFE/GqFHrd7qsvoONHPX8mVEL1AiqIxqXBOzMZaI4hNtIeHHwEEXid6mv34
pCptgWJ6tVbB8Fi5fQqrg0U/+jUUDq/rykBFC0H6JFnZ0OyMDLLAnyjaszksjJw5
y27R2qai+e451/nXSQ3aDEScF0jswG0uebyX08AyHqoVPFfTcBeg6gBd70j7k/Ob
hwlo0EBn0stUEKHFnZpa9+PAh9JDfX1I2YrIJK0AnhKv4fZVSGNUZLczyDHktolN
7UbJ9rtuRR8La3mgMBUYBcr5jdTPho/AMxLp6tDfzIVrFba3MGBpjTjLZXtpqjRF
bvH2WpoxGVcba6bSziGz/2Z3oJXT6uYD8It4HtfDYuzSJh5ntmjsYhGvKn3xIcWc
TU6HQKdPc2PFVU9vszfI4HXvKEerucpPpKAaJ8BtvUPebpSx2TmUgxmi9XQsMLK6
ETysoJHWU5by/3v47KLyQmwjqsRRjGJEevtFf/DRhIeCwe6ahSxp3VWrPSSbmATP
yhO5/eyNv3NyhpG3LU2IUq8CtAf0XZ0zDt/ZGaFazSI6l036DDsd39RzAI1UnxSW
EofGC0w88QCx71u3YEd/NHYc3E/TL8/KbaWeSx8IaUfKj5rXjBcPuvXxzHrX6KV6
P+e7yj/yYc8nD8E/PT6MYf0dbd4P16nzBHRKGnrxKuNrx/raQYUw6TrIjs54CAbN
J4JA9WVjELhb/TeFBADpmO/vPcbFpvtWP3uP9L4UTFycHpBlpUB7qJvh67n6Yvnx
h5dghrZbxh2Noh9t2MLrxYShTdswZvJypfoSdye1RLCWgm88YUKyNXbfd9DaApZl
8lWFPyM7/3Rvc5hUxOrFoxeAyzBD6mmNKUtCs5PWm6DHXl1tfqlbFVzyMeVelyPe
GEaUL/0RQAI+bpCqcAvOfXap4Z9p9w3Mg82riPHrMotXxZjDjuM02dfooUw0ORYk
dEhpwoF2XO5Xtxagx2abFnPqG34s5MZJ6LCAE3/3uiKvbbm1hcBBtCOU2H21LSCw
ulRcf5PHZGicINfxSUYo5RDWEui5dHBbfxY0jQ2l1Rx8y2Uuoc1NFP3YK9dEcsXn
yq1YBeCYVDLtI6G2d7NbqtnvDPjugIwFV524upssfWwQjRPj2tuaSj8spRoSvJyB
d+VBmppL8m06bxlXDJgEnVD3CetQ95a5P0uj4cfDQoDufjsa1u6cUSELT9m7sywV
Zy21MfC0I8fUdBa3vxX4Zh+GFxjCK8Gz19hsI9JexdLRDJ+9wEdutwfy7Sxohh/t
pKUnL0HdB5Om4B+GyLNfngbNLpcCaBWUqIi/Ve5pN4UbKa20N8A7GbCYMz80oKXY
rC3cSb7luMXILEWGoNJBCKx7SKUp4rQdAwcYh7pxWnWMN6p33Z+3Xdb1NTq+VhlU
TcnceKXABRMizOYVg4gWTp4COrnNvYbJUMn2g7NSiwrC6OqkSlWMgWyf6+pWkrqv
zTJjSNvdQ2LeR0NlmVYnBHm3P93GAIIKlcubk8FqUOGtne0YbGKSFUqlz2QlWKty
lQBe+Apem15zhMMgJwc/d8pCHZR2UauOc7ntyLcNAMbpFxpPGJTZyUBwFzIptAHX
eNvH7bcZXpI8pTU32Iae7HZhG1/XCv7/tA+NjYUeoMcvga/QsNwnxo/75DyaL92S
Zut+pVFY7wPQrNC+XTJvgfiYQr8UzYRVYcVnIs6pibVStVnTIspAWke3ePE5s40Q
6LCuGxqsK7uno+cdm8bWLx4/qOuGGe4DYJ1Rc1YE0wynPOrJXmQOC92c2wak4YM8
L/sx0BgJYmafy7GkiuDkIJOBm7GnYmbWkL4lbDJL+Fhtine5VWtYzyMHTGeZVdsJ
89K0G6AYCrY47pgyvsBhscDEAAdUHhVv7xwBT4z+oo5/nRCAhgNUVqxhD98usNGK
ckAn7QlEA6l7/nnxpXfJW/1QlZOyW2NBoEjdmOg0sQrW0HAXBtAgX/KJeEADMBW5
e4pVU24PRgq4tqrVmkRqAPRgkHblH02DYtR4YVzSzVtKKKbWTm9lmk7MGnADh1t2
fldHAtq8vsCRDT94ZreS+ZV1e63vhBL72mr71auOkC5Dq4riRdWxexoU+IlrATZS
NAuImC4JmO9HDsZdgK+ucX8cTVOdN50mXibNjaRpo1uTmVvuDqR4hg4y2ezDdTyx
1oKEz7pRXPyfTsjMjTkeBKeiTg81kC4cpOPEp9w8MENVsynKDRHOrWFWL1IYS2id
j3e9295i2KWFnrJA5w9MKxupysowyiEw3F2LL53Ohy6JpvGqMrUfBsctKrnnBnJN
e7TX4YM4zX8ei2s4ZGXfjNqGeT6j/BcpHl82OOt5t/6adPAFJ+URnfXhom753BdG
zi/jcQaQXC6DM5/lz3J1m8xxj+8Rn7Lf0jpIMaLom4VPFWg5tMJG2gQ7OnkRHMKY
8Y+3fVJp81RSI9lthzB1FPHxepmdqaCLv5NVW+RLu47GXjk6J4K6YV5Wqe0IeyNw
iDn7QPZeATGhfMTMChrZ8n4tF4eyF2eaD8aLmUoP2wtdT4ZvB9Ar6d7Qsj8v6DDO
gBhlcps+Q7qsJFqexDu5UQBEMAPftbjt03fIWlQoiRKs9X/xg+UpRqypGx13Zj/S
8OyhLfSog9fqhmmbc/Q48J8BB8LAgVpAUFR3mnk3rKPkRtw/gxgyWcKZlxCG454z
AGxJekIIyqmO2+u1WLPqWELHyYGQuBJjKW0I1uKieWLo6v9M4XF46IiVI82wKrsb
hHIEeNtJ2rjUX+vrUg+2qXAErfqY5PZnivqfZ5UUgZn3Y1Xn2AgYpk2cHXEcHyGV
sRVcf/bXwv32CeVenjGPcRi9lEgcEK1I11vtmlNPEpYa7RI3XaLxOmOxI0Aj/MyU
fo3sCTIDRSRSjS2lOZ27Xyh5lpMKCnhnzzUOIdSC3XcRCGxZRyVBbIMUi4tB+WiN
BtGPw3+JcQ1LClvs51ho7XTi/wD+6bU4a/f/ayfA7ghpjr8T6yeUnjpaoDr52tFr
SrPh2yrjjZQS7CViX1yzaMEksUuR+XgEnqj/AgymtAadRVLqrlm0O+fYN6nL43XH
9C524qW6e8L9m/pXfBe1P1mduGzXO/v+5E5za01EbawEQsx7et4jYbbTXgEXiR4x
OG4mME4FXh2ZzoY/KEkDY64XcZ7v9lmKfqTlVrLOOpqEXd5MkYbzq2O+O0fTgqeT
cBCUB2KeSvPXTIf4q1qcE6p+nHCzoLg4Onx2fqht7xIB/G0tJViGMiDeUJ9Kp19f
BXhO8sM6Mhj6CyB90bqCgBfOXXBjAz2hxdV50XVuhA0wxA+b/1JG7JAEflr5PSjp
ZsA5hJsikNKEE6d+eZuYP1uDLc7Rzk3MPvtsv5LzAXdRWY3O+uvTvtQ0ay2pAjuG
GvBSyt5d2Loq6vpiS8rfsiLeT7xG5gLtLrM1Cd516zkP4qOJ6WUjeo6hF4jjpPLT
1JnP3ablGK2c9jSgQWIQ9de6ZNV9ICFo8XubZIJn/ucBsYofaJkOk3KGCt/Y91l7
61BPPGxq0cpnPt10KcDU0bwqb2rYYgIYElA8TDyLQkhCAM16UpA/ee/x4cZkZBAo
xY8JbLwtSlQKVw9YCAnsx2aoUDrqqv/H1Nz0uv5Ky7OYh2W1UU49edKgomX0YLuS
Y5z8v9BFbBtxta+A1HQhG0fJg+WyUizZKCgTTXrrzqWaYvS1U/nSwWXPp1B0H164
cvQpcOcI0vkjXpMxdhT38BSaVgHV2F3cAUqT7AxEpnOuXNgsh/43bC17fx9+BI4E
ZjS01nbXUEz+78TcR+aataWLL1vdTbppZ1yxMjJAEsEv3zJER9yqwDLYfNOpWBwP
9s6b5U2SSN6LerMUOrL6qU601LIopnr6dmIfNbxg8VM9rdKJ6LX1T+4DIsTmKj1n
HXG06pIq0YpXs7a7Ok/ejLimuIRAP55Q/179XHd1a+0/XEfs3uG3T1S+AnSkhaOM
1Tq2u48XqTY9Td6YraC2v9xM9uxu26c5C7oO6SZ2RNOOR20e7feWzdECjju/av5l
y9v+PFTx2bS9X4RDEZVncKnWhtTlpE18l9AKUNw1LVn6t9QK0fOw6oqLn0dxs6Nm
NBkbUPed7KLxgNRTKL567Em6eCzrjOWad80VdPT28CiZ7AZn62JyCXVDvMmHO+D/
Imo5PTU8h5g/ySWoOzSOq5iYVQck53g0EBmf/SOnyBBnRMalQRBU5/sYWkt82L3n
JaOriBgSeG65KYPVESfdeQQWTFydG2HIBBG1kPyNGqBN90Xg/nLVqBX8Vy9UjK06
/mkKgtdRFn+AhPfo7ow6xLTLhYUv4lfmiEqjyp8hedpdCa5xIOVf+iUPVMQ76SZO
iDKa4JoXLzSJorpLmrWxuKqfJEtqyrNLm58HG2qH6MAMilHe4TJ+l3Ao0W9JK3rs
/jk5izyvwQDC0zWa8M3AiibsIGjKDR6PTZhm8ODBGmk9k8HAZsEtV6ih8sIGineG
189lsb0gFUZT/NZGDGwyhgol0se2LKhNK27+iHInkHTGMWAlL3W/k6EFQ/MbeCPa
BOuuLfcqibDTutyZZpRioGun9Tf1VObXK4+kHy9cfdTONAOVTMVx+pf3WgCKgSUl
ZDQRNIx7S+73epPtcJJCBVjj7T3t8vMcY7bUj9MJ8vtE3aubI6TwmULusnzBFHbT
vxd5hvHQWIfQm0PYPESIH8h5UH+9Msw3pZirGuPaheRPlOnLjt7p7pEKN+/xUYXP
hK/Zx3lNW33qO4OLix4Y4mlXcTcxoq4xf4sOp9oBw3/zc5DMcvDEkVXKS2E00jnz
l8UJ2GY4jW4HsTCTcyog7Sc5EhPzUxFc/TSIW4ZmuCdgK8+rlFmxCPulwGzied+3
Me5zaXqQyJ9aK5R8bXiNbi4lECk8G1hlGfPep1+XSSFm0T5APgzeVApWjh3ktJlI
XLI4pdM354OchtDlcEJ8jsmo8MVmnD6VSxRCM5KiqT2YVVaouqLuFdHwxsxqwqzL
oAquVSNBmdviwcAytzzyUJLKHCb+9kET6X8sWluYquMnJ8z6SkS29HYLijI4at9K
E8YpxAmzH8M1o12LSCqOiSUIctR5a05RGoBvks7sJ+zCHqWI3Ece4kT0aJTuFzYu
ulsjX3V9TWW3LULvAHqyEDHj6IPdahVpMIdIUNPmnYO+IwWNHxjAk8ccMWqroPb/
n0ucaC7Q+fa99TxNNz6Ikteqj8DiNTruRzCjNW13yWNYBlQCNBp5e60JcdbqvYHl
r0pHj1vLE+orvsfjiI/fvgfZwn9f6FgXr/7kAxYopxYMBS2RgT7h66wvn7gLU5PC
wBW9WIMSQ2WssPFf8Niaf1aRKMXK1P/IXc8WO616l9vQBQMyg5S+iiZ05rOuTKWs
LXt3wSWPSKVm09lWnM3EQ/59ha/DBAY2pMkBNIllu0+56UcPd6NR1c7ZxxsPuxi0
srIJUc2kmYzI1Zx8G+E9Ro9DocqO5DGcS6NtYOa5R+NXuFw4Ry5B/3R7D1vn2bLZ
kxjuPzgFWfdj99bofupWOgjkE0hg4V5YrU2aEABD0EvWsiePiNudXYmOTeQc7CXL
ZEAISzDVPJVQHz87ceRNJh6lZf5ut7zx0OpXG8nBcZlYnwOOgHIdxXTAn66ugMwH
8IzjNFQ13JMBq93SWPk4LmKRRlHyYiaKiognlE1XjuEFqhF4dAanQucU4gbPrSZN
ABoMPbEBa+59qPXEKB0kmhM6cI1DBFPYRjyOC1MhSmLCr9pXf2qaCp/ySZTm0Fh1
PXJ7QeVSzy+2FkHavvm2Q01cTbJJxpTbdkErvjTVseL9nRrZVJBrlMmVp6xqkIGv
nhL7yYi76IvLf+r3v51MZdAeE7n1zL1xQp57rAGSWUmYF0acCVEcoJjXMnUmWnhg
xDis09QmCdA5d+Qab40Sm3S8TIkQ8314f3xNucElbMs/qf5goYm5i+UlYWeeejPa
sDChz2+CCCMDgZ1v9zkmz3pfgQ6O38ccF0OX5anfGPF23pnA0bdYLK71/QCsKAhn
sF83ZqzxtEgY4GaoSs6Y6uG//fouQUMXsW/Y9dr23u+k595XSWJq6SQXkD3wBfEh
eR2BRimAdaGc8UNxXCbSbrVf3qPDHZxWp3OOgt1IGlWhTbMDMp+4oEbodQjHkz54
RzaT6sZcvAep1E20EbHdPtLobfXzJ1ROWZ5ZI51zUNnJ03CHLCkJFZpga/GP8iVX
speBlqvlNRUkr7P1U77sA5Y7XNKnawvFTgoyyMPelZ75IioRLsbLsWnHoU8RBjKn
ZZcNUeRCwsgdgZ11rMsnYQdk4Uo2FiccOHgo7oEsx0MFUzJtKKOEyGfXodCSr9n8
Os2N5whnOiMuTPgV2xG6ZUCyjR8QFTUjhERXwJpronM4cAICiP22lmH7INf44z4I
v1UADuJVDaAAct1K5U17/fyDhHPUI4TMSJwpY/CWPxbT2SAw64tOEQxd/jl4SxKx
ESwJzaZrdIaNX6d2m3wsRLPaHGMtJoX8CQwjwi7LCXjSbkf8mMPXr3OxpR8jaHz3
IH546I7nEo/+exqNF7TITqUJgsHm2kX7I7N2bHnmbmeVck7sr1cGXWO1THJpKWzI
3/Y9Yum74NVgVEhPAIKWT5Ug1zUIv1mKeTyczaf+/+ry90+UdXk5q29cg19CCBl2
5L1J0Av6r92Lm87zRqgNERfe7mrDPqQGsLxuhPLKfifQSZsgYecYA5gp0Bg3wweC
P8oXOV4jXFEgW7Er4nHLHV3O3tnuhqEI14VCwQP+glDd4TrUDATeeP4v+iKZLhVR
vYn+vUxNZriJ1/keiSC/iIx40o48wZ56xz1FJdLXfQe5mf2y4sqlVqrU718kV04R
2+4biN0M4d7enPFOdf+VGMuxZqiaXGC4VVGyYtTfw7ZDQUZdzl0YtZOAE8y/lPHU
H67Jo3Hq787UNR+AR3mbiGHK3eZlxjNhhx3vRfma0SsVEAE0YDpPM86I27LzhPCV
TVDhVU30CzDlhsPIz4PDY9BPSJhGi3/NqaH7iweJ85BiRwAMeGMu50tmxp3Q/Rk2
k/EeGB/tnJRKxeZwY8u7gbiqZZPfLVqOGev4dlWsd6RjypEji08NY45IzWA0XbEj
y9eRhBvIlIy47QUe6PmKzWjhE5A8/qehYKa2Cpu8smbS51+U3W9RYOLtNd25w8wM
9+s3MSp6VOCg9F9mDUJ5RnTZ686eyTSu5ivLuCCu6tW6FHME3dSeI0ea2d8wwmpB
dcAZ43l3pS9Y/IZa1z618Qf+hiMPGs7yT83lgMFUwvBaWQSNoU8ffz8hHDAvh5WJ
QQy9kNrsvmlTNM0jqaSfC+RNTDpp3I1BuBYzrhRvQTYYVPW5aCjLck3jbmw84HbJ
TUh86VYBbm0MGMoifABjn8vD8uQo9Y2VEoAYy82CmhJLGfdy3xRiPBB+eOUaa30l
2DqFxCaZ9kucfmAqlx/ZvtWnkpqGI/iHaijx0+DVIMYN7OjgCGpquzItAgDDotIn
rHMkI2+51KTOW24hqOPdscxUnTZRoYmayQVQcZWqvnROidZYQFhYmvhyY8YYOdji
KAELAiOnpXA/vgI45WEI+47po8uLQWs3JncYHT5BKXr/lkNzsBSntoEJ6lnLmQML
RIGjTAZiXL4HExw7N5TaKvTNC5kPDl8CaRZy/CGUeipvFjVe6llobQsBO404G+Zj
tQAhoagQZuBkSOdCU6hycNOP87AYs1HaYAx0d7TJLbfMx2OCCtZpXpU9eDnye1na
SeUmlTs0MlBEV47TiJ2xz64C/nflsFjzykj6Ww38cyV4uyfCtvBwQEAwq9nB7HNV
t36S1qJFDPGhS6vMSQ/Z/TaIAAnSZygx72WVXgE76VY4aiKxaoe4zrWBw2JM72fD
mG2KYuQRfhE+U+GMvhPkKmCbggDGtqmC7g0RxB1SPH6aV3g/zZwTLh+SoXDtOJH6
1u/Aq3GGiNkjxKQqyXa1Zrm8p5tneznKROd9lz3Scz7Y8cqdvAQyxQ7OtkKh/km0
t48MsMmpjaStYY8LNnrUAAi64dLN/lphu4c73QkRbBwus/pdaqWPE0daReZV1ug1
ZX1eZZjssTyDzyUY/eOj3x7oXJclO+6HgZ6DLQqkY+7ZuHyVzX8FgYxlOz33xwV3
Bs2tWeIBE+8ccaMQK3ok4QrblYh2sNRZOHeW9l985KBHLsJf48tNIPag5B5kqnba
ixwJbGy/+i9mlOVwjjv3aUYzVUeN7tNKZqcQEY3FJnpdokrlTIuWg1KsAT4vv1GV
t906chYHb/Uh0+aq/DW4lpV98SAdJ7Ldb5NVKnRDvhPEXqtXBxzzu5PrS8s8+WpR
S4YGG2Q7vXC7emjNo6af4rys799wH6Vz5iah8xeAQpvaoufjk8+bqkmQUyyKqWBt
VHt7RFM/2pUmD2qWKXj7xBE4VO1SIUj/Ah1KMdHDgrWEElGZvs2W5s4ifNBfRwPN
9x/isn7tW3RFL9csShAKFw2RvWjameCed0zt8Vh0Vy1fE4M63pxa78p70QAUDr6o
eLUMz8Q0nJCvgphyThdRA5ohzjijXjI88gDzss3VUcIhuLipXYld9/ZgMMAEFMY3
WCCvTmVKr8UHctQYvgWAFbHQ/dXN71oIEno9i9I2ZxuKOjM84t2pzrO3NBjDF1Sh
t6lzO7VEz+FuJQB/3T5/MMCM5tFOXYPqdhxx6xOoMR3bneT89g/GjhscMSaKFC5u
ynAhdmLh6X6JLGBHiIf3QVqwguvDn/hZQpKdy5gc/RkxnaJzVZZ3KpXQb9KJbCMo
it2wRt1bxd5tmUw7cE2s7RMD3i0iXZl1Iw/Wp4BIs1ELYVaNgkdhGkQG7z+7VuC2
35Jan/rUF3eScvIFc9eFWJEDNQub2GnyZSRcL63xyJa/l+wGYAODHhhGywxVRNoB
quYsdU8tcQ/z/NmaHywnTRA0XjLpdfgROVub8gdEt3SIXCHgDDzWt9oNQ3yn/sE/
GpR83hxMEuMi9TcCibeuySxy2oc9dcQFR7OXJc6083qbi1A7/LSKB/VhxG8A1W8s
9GNDwXi+y/tZwFdOivSJ/JyOD7mE2ZgntpXjj75Z+WZaoI1mjLrSF2eAfchN9mtU
4vHVJuMfxKzyw/USutJ+oLZQfN9MgSI/R4U8pM/3DXsNAjK6rITwXgFlBgSnveFb
nS8rICsMwu0lcDWeq0J3TYmx70GCZQia0xrE+ElK/eFAgnBn6oLGB2bUSVe4+hIv
qE787Kr3C8X4jhF+6L4aNv6SPqWoG56UPX6wyoBst5l+wsY7246YhNB7xoa86zui
BfBWWwNHnCORfZ5GsCayp9YaI5UnKIQFKZ2DH30L/EdFeusq2QBR11XjAA8Bp45x
75hss9h32/uWUfM7HxBdTDexMTW6JgQi4Cn3zEQrd9/Bi2z84TFpbWCT6gxhXb53
8L6aAq9r9ABlcvnMU8t2orXMSeVIznLCKdWgFEo8Z+vgiSkI4xORIgBUxE0e/Aez
iFkm9RS9pm/G6fsugxt/MQ5bmBQO8PtES9npeE2r7CU2F3iq9RCfJpUPrC1xnhYj
Vm4brZkoeq56tJNjIO9qpiTVRvYL13ehiQy+0QNk66jN8Ck5BRGFUTdnnBjq8KHu
AKM3pWEJorYjs/NY/5qX3BRKL5oSr4qj40QJUVN9A/SfnlH8/quvU1sJe/hEtySr
9uxjwbqURaL6wma6Gq5lsxuJYwAvxDg8N+qcvFNUonLqdUEoHNYccrwRuq/BYZ2+
cD4h6N1iAgnPbQcL9hAJaBYj90KZobOOkFBhmWIv8k7Lp+UzWA5yVk6dlooMBOKY
w9XQ50Ltzfah5YRJfK5LH1nBHzfZaTnc8/ayHYlDnqu2lNpKirRDrw70B3VELoN/
cJdTtPV6qdVbyjrEzEwRTtkz8hGep/pXtQiQcDeQhb2E8dF6e/MtmgI9uzOYy5kl
7oncEA/9GoIodXiXymYBNUWAwuhCPLWBPVUJnRVxXyuJUEYULcT+5BgD6orplYhK
UzCHXko7bL76k0bap5H3f9WKfSD/Jdf/0ERHMgsfwEzbhrX0sKLdAlv2ESMjbpdS
QazaDdy4Fc4cH4zMDLYoBv6ymaR+VU6SNWeqzCxI9uCRfZti9ABst+lUt9C6fU6K
CEahSP2GA46JibPz3qHgdrxNTeY9B5mi1cC1yiDr167d7erVtp4r7OtwsS6eqjrw
TOEhJnFtVGqUIb4tPFY/HLWK9wZ1WkhxW7Mr8RcEvQ220pjqvHOdVuxmALPlZMxL
mhXR63UJp3JIrw+DtHN8YqE0yvWCOOB7kUh/p3pCXeLLVEDruAGo3+yxqNNWoKQc
9sPxS0qmaRDxfzS6GJLQm6va9clgOCU16McVTB3wh0nq4L/hHq+u9pEC96v5fHYV
eREKYaeHZNvo496yglWLbqvq2AB29r8xSfuzIqptO8zOlOtIQetC4Jd7ZFuil4pc
wVVTtrkPqpPwplQwb49pkHqE2XPQUG8L0pKaNECcLbc48TQuN590zO6J5aZcRRFf
rQoaIv5Bx89/g2yOO06PZUQ/dtx+d720nocxU7MRfayQl+A3/ztvBpdcS8ZJd8R4
nA+VWhwof61jkU/pB0ZB4H8+LLOCbSV3PtOEnOZNfMTvS+7YI0iZNRaWEV/V2mpm
atBP0ujRnpsmfZe2io3qH0mX1T3O42ies+hcf6TPeNXJ8xu/iS4bTixqrJxafaCc
CjoVxtIfI2K5NYbKM3YblIdpdqyZKMKFI4BURWnfukvTrzdAjwpUUSnm02UfaQX/
JFrJ200yJ01EGUqiuUTGfURDs9SkfRFb0u3c5SfRLc+4vf5FZWoKimXHJ5I/acwB
NRoMgRngy9/LZ1YyBA0xXjJQnSNQdaQs3Oer1xnAmerCxP0qFrB4cwHR4w/W8Tif
UBdCND1kkWYSFjA421o6xRPOiVTqmVp8ZVFCOQx1wTsm6vu0HYwlXA9z5a8Tg+Ch
c+JPUSpMwup7OsmH1j7+1DEQq+sreyMb9djve8MI909Efw2nPTeAZMHweByINvSL
Xb7g6ixb2Q0cG7ZnYhnouvLaulALNTCNlr6uQ4TjuNEjl9hKMj2LpJNhusg8Dztz
69Y+PvdTEe+SLgmiaewWQPX/UV8GKPxvD7fSrf05tbF+BoSWEjlHiFX+ube2f5fy
uecwu04/5vcQIiZT6tCFXhj8Fn7n/78al6TzyR79p7jSCzzRSYgY8hjbo8SItgO6
3FKnTEw6Rcl7cqh6ye8qEaUnCoNEo7kb9piW9gr4A4jXAFCffhb9MbKKT83O5HN3
SNemMSkwGCZaFA+v5c2DS7B6SxAue96VzP42whDSKKQMLyvRKo2Nvcyd5U4PwuN3
eDMBlrPclxcWBcGT0tRG/VzzaxdGgUADoB7h1lULVStunNekEmQXgkPRUlAkqzCH
WZO1oqZbow6AEJWTTfyVs1tvLuIHgcQH44n9aZwLpF9buQqxYvqn7hJauamlY9CE
GK+YvsKZqC4gv21Hi+Kjt4j1llXRvYXrRv1BFk330cTRQ3lfZuIeO6HC2WADpAeJ
VU2Pf8pUO11zcGE0dzMK2TFged5rTOI6d2xhYsm7nX6m/MjdJV6tWBmrLNoKjf9u
2B7kMYN1bwaqqCfGuxoKTNypxpOJptC3L4/PIUp4rB/FpU7Olwqw4BZUzT4vpHie
GSQTqU/HloqX9bXwG0M4DK6ye+2RgIw829M4K+caGFdTlidPtCMwIOiyzRcTmX0F
ygCXBpTswtuHgoU2RuZZVv15TvkJsVzn1lRfAU0044rvbI8DYC6RoTlA+ZrSZ0Es
Qv9iR6furZvAolnx4oh0nC8X+zrb/kWp8CGqqHZnUUEtnKoZ1eApAXSxZv5vkC5B
cXNqxQyZeQWNVE4Hn71G6pWI3zgb46y0xCbknBB4ko4o9YF1k3Kq2GvAiD+Y4ZNg
boh92TzsDy9fmtVk+WwibHr12KOJNk77VeMMyPIYLYt0FRb/aVcRsdhXtWTtNuxz
iX+pkcwk5d1mMa43ck9QNfeKNB8/5DsUbXqsOgaSS3IlXbEEJJDQtG9P3Jv2S21i
+v/ES3chcIJKAvwAzukEjSnsEeZDVYVz6bNpH8cASoySTU28R7/Jxm9Jf5G382Tx
ZxjVL7lfOsopAAE+7siLoGiSV1PSsBA2EsSWVIxYMVedenQOPSqQqBGUtx7b+EU4
qTuRSY/ey2F+vibUYL0IerhS5d7RbADpP/LBJx/VvrSglMZyNNV9jG2kpnju0YCu
3PAjuufe/dDXWMWgTAMaImqM/oy9mwNIzfb4K3sw2AHzIx01xpmBh5KEHmsYBpXb
Z5lWudVM/OSqO+vLOAZtduxiqMdJ41kgwfuB6yWiazsbFrf52vQJiK0psUZms4zb
a+AzAp9Yzkhw6lxvxQr3n1tj6+LQMIqaQJVPH+Pf65RSdHmB8j49mA3DJNlwv/hD
tL/U/qdSTVkCI3iSBnt2MpDMb+c08f+K1/hxJ+9C2MkANRfJQTyZ+7/rb6+J+qGS
ud5YjW0/X1asvznZWC/vDZN6XkixgJLbGboKBj3JHTsmWWlZHNZo9NGLAzECZXwO
PkSaUqSeDbA8vC3ZDq2eagtpyWz9Yw8bQVZsYnLV6rmEVWqnqpIMtKqaiG5pHIQ/
SFNUKgUDturpkIoFwu/XCxgZeLAAhLVx2pV8dpQxA8JdEdDkUGT+9V9qHXy9JPii
yLOqxF+K8WW2ZjKtRG0qhxiz8JFmCAPXLjv7FPmPpDZlJynRNPE+0N1Tx1Ac5ApW
rEktLhWRJoggUf29OfsuQVIrWhhDojCv9EI26WoL1diIWdJeir6qQS1uLUiSYgtY
RTtU0O5v+NsD5sZe0VxJzYkUeyO+KEgjZK/AE0NKx3N8c7PBHsdbKLR0qb3LYsIa
srl+vLMIDKNY6Q0GGJ2L7jMECFJQm/vyueFwToJtYrwch0UaO2ZGRDBdh9Ay7u5v
uCQwy3FuJeijIG7P1y7wFfDzzuJml1DGqRnUPG5V/pzrCaIfySFHa+SRrAnA9XGt
4KHbIY127zS46JtToSfsfqbG6uuM4L+oUsUBcAgDz4dcUY0wNpudoQZcWjAeBhkB
jasm9tuccxLbe+PKCXO5HWey1J9Lv37kNX1yw5TVu11OkpVvcORJAZSdqiD7F0q6
vVsnI4PA+pbR6rA+mXmksZRTUlDWufyGRNin2+Ld3Pavq79YdzbmGKaoxnWUKxSQ
UIi+AYxndShFPVD0bee8VcvumkWOetWJdk323qdICcJ2e/eUniuSMYtbuwfmZxaQ
RFqAOKuLnxVUp3KEySE2niv31lxKanwRx6WUR7/JzViw0pqDXfBUyz2mruPPT4dG
+Tgo6XTUaYQlT57Bs9zfW0BVRVBauhTpBiar0RIYzBHyqW+O3FCaJZ7o3+YV32MN
9dZ/Ztm3P9PRNSQQYHtmbCo9eTHFlTPUUdXUBB6cDbA0OCkPx7O7wj/qFJRGhGBC
amimzpVlgWOQRyZoK1Q6U4wnbguiZ9o+1FP8TjHv/iOfBy3yxGlh9JFJ9wtGAC/N
1YSJ6q6c5YZR9FT+c1zbqtloZye4cSSac4VpuUgeqet9N9svob5sfim0mDdnXjLB
AL5amqYnlHPtWb2E6NtaM/S/DIpOLtJTJEQuFoY04VRlhM3EaPk59xayLf17v4Id
36NTtdqSyL5q2mETH1mI1eiw1+3WQZZm9Y9cQIpV2mtdXvWWQSIiQ/kTrR053gXR
7VG9k6LK2a7FXlpGEnEo0f57ty8Qt55qICKQ7LwZdwO//FNERYH6uSwDF6G+PwNO
uGJWySPvmmboeEYqC4Wala0M+GbcafwlhxUNB1stNUsHyz7EnZqWoNKiBCLZkp5B
Vtd3SEyIPyrm+n8Hjk8uJEp8WcSD3eXezo9BRiUXNnhdz31v9YCxS0u1BHlLnCzz
1I6DkCOWO4WTpL196r4tKPWDb7WF91XhlCP02IT50xglGPeoU3i/uFayaKGwXt6S
JJiejDzwiTQMEILFyJFJt+jY8mTuj3ue4Ed3hekGUUVXxYhiB0ev6jch2TWaoKu8
Ue3wTX/DABh9pb6JDFnij2wLPXYfkWc89tWL59IP92bvheDDUaxbyaZEedmZP0Sa
UFpgZPp75+vn3US0l1nQvvlcZNQP4Jnoxd/SVfS9cZ7rLNz+n8SaPRuOlCsRBeqR
PsxgOtL61hUS78lCNGEceyI6ia9N1CLua9DCcu0Ml9fMMvYIATHouHGiF7TF5pyx
qKnbzO1GaFoalKtTCj5nv16ZHZ4hL+DQa2HDfCv8tjFe4BYrQkaAGEFxbfQUZ1Un
QrZYkBIEvyHb3U+CEK9iFhzQ12VcVKLP3224lLP31HPU0Z5cf6RSa9sL3c5uxDRY
B4p7m50uEn9NC6Knd4ejUWrurRTq/iSrr0Y7Abdz5gwZSD0qHkBelgklPe6ufny1
eOs5inE6KUTORYGr7LyT4WJhwKXw3dAig7pAxzQBLrF8tlGI60dkW1QkfT9va4nN
vJ3Lnd3KTPV8se4OxfRUe0EjMWRdOMmy1tQRg2rYnEnIfYvrja77ji+A3NfkazV4
8AHY6/w1YjhREc3PLYwXygJVHdCRmcCHUnRklKMZeuxLOqnvTUQx80i8vh1mTDVN
hTAZjo5uichNqVhdDpT6t7/mvr55FMJTXTBXC9espBhbqrPbAju2w25n6mfoISdj
fZFgclOkYinesMR+vhPYh7gDCxjRZR+AGLJTzKQ5uXcryYRIwz5Kc7Wnv/IVX7gW
RRP+My5D4KZ32rYvjAMzHpewiIDtJFuVnlUR/L4NgRC43Pmwzvi6y3g0j+DJt88x
eIBRh0v6/BZRqvQTVnlvKWG79BVWN+bTw7z8NMpv+6np8Qahln2h0zWkyfQVHaow
A/RYpyvVEAvtD9dCd76NQZRNWGFNPZ5OFJfi0Kg/XID41ISt7Nt8rMmjPeh1Pw5t
+MAoRrU4TysXM/0CA8c2MhZSLBNyNdOZwo0cjV9olgR/OgeYtpI1XOshpz5/t73z
JbMb9ccqeEa5hOxJo4gDq88+uum55krmhuZ5Guqpjv/+IEbAU4wa6pi9eenv/bHy
K8WojWQ4azS/DRaLOKwQxKF8r3DyKzgZcr61PiEw6YLfS1tir921H1YfK++lj3u6
xvTkSNOqpN88pcMSYcPqluCLRedtVkY5E+LxfP8vROV5011BrE4B8t8X7rGahA4D
HH+swYj8njrUEZn8qt2AzfAhYGjeR0fw2jRVD4NX9TAw9ItAtFKFMhZtR0K4/Vjm
fcMLx8XrcG6mGxKemMWIKKrhhfpz1W589GonYh31wFiqWedszGvhkXP22awpmQl+
kH/tltmeGRsvhLykJlcx94VebOU3j75aBHhmBuZlLNSM/sgBKUM5pN5S/4NNc0gm
gYt3fCjdQfVZxT7rK1OTm4VXhUCM3I1DtMsq1OnvRcUWhqxFrUMq8P0NVtwx7a6y
WAS4IA5cQ70tne+/fX7O9KnncLJnzlBcqyGpmRXZKq9fCfbFaYx2Rqqu9GnhkOEI
Hk6BzG8RYbiJ5c6TYOVJIb5vDWPG6yJdiCd+JLNq0IBrMzEEGhmTInTK2kufPtlm
BMKNukMdLJPgOsSxtknChNr0xPHDj04291M6JdRci9ETVPkfAJgK79ptES2cAR47
iE0OQ+FLO/VpjfByEwKKC8bF5viyRNECCmwHpaFLyHG7Uhly7stGPDzudpjxDb+x
bmt2UOD1/GTnDsowp2gX8DoY5MJQJceKYDkd5EJJdSky2DqwUNnjaSrZflikoZ51
hsaF3bDvSisb2SJ0A+SG1pqRbFsinxI/I8g1ANaqjQBc3YZUub3ZzrJnrlLqQ86d
k+D5reF3sri4YwhZ1yc4LHuhtGV5uqyUz9biqmLf6oFJ+Lc64zeWKQxKB6xWdThZ
jIuFumhvO6q6qacQWMCoLywCn+Ygb6LwBhkQsP0afSa5Wj/T15pe2WXOZdsFCb97
zQ6dOmBe6+XFnU/ZKSbaEMvXLiMjGfcwFCOeHRRVwSl3XIQ15wzQ+Y3CXwUZal1p
3BBPVxeaviXL2tesoIVzlA9auyFAxfiPHuKTDdJ8LmElWt0b7ErrKSP4rWP61KX8
/iu2qh8FsCDkmIy4MazYPsUwhK3ZzSbQ9YOjkSjF5w0UdDHXL1KjnjKHL9zF5wew
9ose5hXiUVeWF1gI0xrxjVprwgQ+PmuDS30cETlo496wf29/lOAwiR3sAbJhKpyg
EO2/phUgIpZC0/WwwQqVvBwQKfi+VS74HlrRPtVuB+bEbD048gU+wVJg4N0zEjYL
SxJWvjj7diWuTe90RQQrqX3IJTQweNNf/JVxBZIywvoqyzKDbWyKgunAV5sN3LXG
Y8VQCckNDCPOT2YYy2FQL/QyNpOtQmbSjWrLQ/VEaHjBB//mgi+Knz7b3kzcupY4
VwUj32lhA3gXgj9GxXOghQ8P6YZvuIQVVnrSWsQ9cvpFpHH8ybFfy6ecn4xS3ZKj
E6xXqJC04OeayJ0sumjfvS2XfnO+dV694OaZ/SWEsLweSWOf+1ykdlGbMBHLl/F5
pGahf7Er0/N2YKjiThIlgfu5akl5n+Q/qtLcp839eKodO6ghpsQVEd18JnjCSP0M
OHQvTGayQ1O0oalmCGnhJK+b9yYtexHdrIl/IbQetW8v00xgjmV0jqiq8Jg07qZ1
UFol1N+BPe6MX6UeqIGJeECY5xtgFzAA1/OcqUBKUDnHVLLPyKtdqHFq8OrF3Hvh
2ghNaN/dFk5spH0wcHsJfjrCcFQVL4sJ6MW5em7RVwdY07JiVc76svU36ieQhNCw
i04T9tZerimCv7ZhgH+WUZa0Vwfs6fm86lgkITyUT4xd/8WucF4/7yofYaNVpZOG
NR1UAyKdK4ZsYmv6UiGbxYu7N96/V4+pteecGbdM62qM8CkVD1ysxscYfsMFxV4c
rhtIhs10TgrM8TGpgy36q8IZFvK5R6yFnpQ++yJbkZQviKKOas3HKkqq2+HBuR13
P0jVLv4eOPRWzZn3aA+OSgMO9nBP4O8ePDYwnrJEFFSA2kzLe3YuI1zyOBS7KPvM
0062c+auNqLrbUqRrJH++uM46iUTitmExSMZcKiikOHtELO7Bta/4kV2UFB1IfnG
F+wdJgvBQkkHK0B9twnTzoeUJgkipVNlNe33zMwVJcGai4hntRT4VDE1L9iQigcP
vIixS2s0WtcvGv4zX2sotqe3ag0dTN6WZ4d94GyaRaQgMSZsB5vBLXqWShJ54p6h
Kdu4Rqtbpc7OX6YrNVpwuPM9gUtjDO5gBtB2VtJ3nWDSMw+LBeWXjdBlYVmczkVj
yXENOlXTncfpaC3lqSnGIGLxA7t5O2U7kBrSJ35VpUAzvehXoeGkkp2EjZgaUUAW
93TvpyG0wPBPxkh2NLm9DPzcMUgfnpOTKAgCmTcsYEa3fOc4pYx4tMrpzef1kBWR
JiTbw/Cu5RVVfqq18tLO4DFDVYxipQEemIBTlOAtx/Gfw3CkPhN2U03lGJiqdrTp
62GGrRss3zXPV4PPqTW1ZcY0hj/0Mr4DeXZ/OU6HQtXciOyGqOndvHTHi5a0OdbJ
OqdoOmcRlCG9KdRn8fM79vMid02EjgGyoyKP4tmVbLYnvPN1ntRiT/+Ok21lYQkF
Tkr6ST7nsdx917ulLxgnmwla+lR+VinGDZJHv4vf7AQi2eGB2wURm50WdiWkD+J9
ZUWGHuDvv8K99JB1A7Oo1xggR15lRgc/t23feqYy2aY+kfXlLXe7UJKUaRczHiYR
uUDJ8IhPJTdV7zUZjXAeXgjsCOF88mJ937Q902rc1A2fthYguDJJnxjKVYzcGe3j
xDkkTwhTW2LBok8PPRlxqoZkKxCd14PeBuOoPglk8FpPQRUBHoGhUwm8LibwN5TP
/XwxrhkwbB27wq+bQQ9cXMwh2E+sQ5uWZuNh85LebgVFWNs4EmmYjN7vCKURvsfu
5fwRXhY6pkwkt5cqMfjL0nDuZf8kcj6dMxKR5HmtEt5wJPuYth2SBwXU9mWgx+Xr
BOdEHnoTrLkdLQpCMer4Snq7u7ZxMAwdZERXtARqH9Au+4gWNjip8gbK+iPJMQPJ
3QC5Lrk0k/D8ONjQfBRwrX/37MbCVJVlq9MXyq2/8EjqLg8Wqh17WTg5oMgxO6O/
avMD0KCF0PfFtG81WeVWmI+S1UPrQEV9Ce1aRBE0am1qR1Xv/2SRnB+flBr1iSa8
0XTTs6UYM/qEf+LLTxSttqCUASbcbJjUSDq3G8P5IA3KCicFtcr34KLTxsnA7P1W
AiKMmgCoGX3/XIhdphEljvGng5Zre4Kt6NkRwsStWBKyDeLBLQVZZ3m9H+RPUWj0
Aswj19DFi8D5lGOQUnNiby57ooeXpj2qWkX0k9tYlrzhVKQvp6APPAG3EwLrWE2m
iShd6CyyRXrinZrtCebxnc58dkFTTANTAlH2zD9PJaxiKqyNMrpP2nP9JtGKunuC
TJOIlDCDwB7qg/zeOWVoDnqZw0qvsWLMfoRNnZYg0yQyi50brhE+6UXqDwOc7drT
+EQF2Un7IrWVysji8BkbeXbYb/kqpCAUXJbDwxgjSZ+amMku53oLxVTaqc1rAAbp
+KYm8SYvphNBktrzPGNQ24uQ50du3d3B4xDjjqsJ9/CeLLznMjTYmZvdZBEdZMEi
26n+d3lvYeh0sWPWRyh6RzTyi1GfRk+/tXMM0KZu9J1Yn1OCUn5wLWUA+5WJGHZN
p40X6yNnkPoLFerEkSBl8zR2EwTt2qi+2dyLT+AIdYRc78sTrGHec392XVldrrzK
Nidq3NdxmtVmZBnmPwuOAW45CYPRFBSQUd/X34M2DrVIVOrLUgFj0Qb+SWYtiyf3
C2zhlk2T4ddSpVPvpphWax/YZKUCjrc3ficYpPNn++xyFbQJlUbyCIFGGBZHdJkg
z1JFkOxYGSXCdcLg+J0Lq98UWpu4VBX+smZaJoNKLDFbYfp4m516+OtBvEXzl+Cs
9SOpfYTmfecF/qWCx3rqxi240XNdxlneWF25RmJ8DXQZphb3aI2VemEqOdGPfIm3
8NCG/kY1xaqEYp6pXxfrfcoyJrR2xuu337PWq1zumZpKxxdwuZMjpwQWNQmFcJqu
bDL+pD9qFk7ZkPhTC4LoAoOapIoLhe8P0YT9ES6xMKJ8qu5lC3dxEk3FcuY+ga7p
Xp1lPbqRMfwh9Yyu4xruNjx4uRkuekfFWPRo2/z0N2FYnpUysgR2WfCWEvj3riD2
lxru4ZriDuWbwFcdghE7VoqWltovxbUp7/O5iD1aKBLUy1o4Iwiefins3QZ7ETIU
l7kberPBBOoaQc83mIBhJFSuQEh4oqXX1+/nHQzledi5kGTT655ZawKKZvaGEYYq
rXkip3vBYVh8HynWCvkCHoJzA7ztTI34P9SlRhOs9TxLR8ke67vyHO59rk34WrSH
UidvfHrQL7R58J3REoAztZKw6kVDIMb4uph7hAjBM17VzCla3YyfxpoGLLZzU1zY
7VsW8Y5PWhen/Nm+m9aNWsLLSmZknijYIUsSdHOmCH0S+ZQbRcuhDGJQRaIlJkn5
Yez2vK3VkfkP71BdLnAtAKeBS2W97dggfEpLGBgzqkIA5K/p1u0BDQ//0Jvho2Wu
YiXqz3xN67zVa1K2+KX8J6jfNtrsaDThMYzULnNJgQxTgtZ7zY3u+ToL/VlReiF+
jHcobRyLKG5od85uFyXIvBa6S7/Pu01vHaEMSMddLoUBteJb48pUJHmd/WwHigZs
W65pvD70s45DFcuEIYSZ5rsH0mUhvSxpKSWgRQIgxFuRIOWEnquCnEJ08hfldEQf
pKSIeRg5eEd5YB7H8o3ZWakZE91eu2P6T+4FXlQcnvs+mg38VOroS876F9zDj3Aw
N5rgdPQ8KK5anhFy5tZ1YbaxO+cUxfHNlwil2JWKx/+jZxz1oyKR5M1gPi3sdjJ3
8zlt1F5Os6GiSHC8Siea1yt2feKqhVlGCBANwcZ+sU33C1D8mDZX7wqroJL0TDO+
xHiIBtfR/NtVo5mMFKroVELFcinWBt+w2oks4Fn1rWsDRpkTwEL1nF8BPWsglybp
M6wEG4aoREQ3ku7Uzaxn0l8SenW1YrXSX6kk0sQ4QpVXTDEhtWIBjfvgPvLkd8v5
2GvFLwOXukGTjZ3HgDO5MSxJsGRDwFXz5jdb6LYtvfjBsA+fH9uaPZRBFbij6p3v
kWyYQsqDxLj40hVD0VGM5BBGCq2VhoMaPfmUjbKEIg/eK2YKUZw4BBbYCPx0AFJu
M+MUZOeONYAbOlQxD+85hR637Rb7vDTV5zJr52yhcAkzLIHC3AvJ3OV89+q9MOoB
H2g84Tmi173RYH3NCskMhs+no3CL4AdAUGNKGvcHxPid7E0HS05AiSAFuM/eb1g8
ORFEDsKIJL22+BU/ysQGmAzJZ2PWOcuurLejjveNx7DsoqPI5zkbS8ucPf3pl4fe
hVI3dMQxJyyMd3DM046G6kL5nPyTyYhqLe8ZsRO3MGN30BygEoESZc+qq85U9hIJ
J716xZ49Xwdjr7Hig8pBkEsDvg6pwHTZi6r7mskjM86BcOvuF95J4OM0XyncNxA4
BprhcAeOYH6kyPhf8q26c0tl08wQuT6P6bZ9saXTfltKBpFCfm409viHTNJr0gyr
HcPDnE3XWiSHuAOBgfgE1hPdRQE+9buU4tb4W1S98/EiblgedabTtrecBnTGNwSd
EUdGNfRG8NGMRilDv2SAreb8ehVzUgQa2VP0wTQB8GIUrpoXnLRXJoaHN7nhSQqu
3THURf1KLnRkHkRPlnHPap8O8mJt0ixAlqGeBxQa4O6sWwJs954pU8/bC0Sl+Sxb
C8v2H5sOLenxcGsN0JpEm7NDqLIALz5TVAlxe27mT0SZmKGJ8O7/UKLd2+S48CL5
CuR3bFqd7dWIuFG7C2nVG2YoD8qCpdEGqF5G+Djfqs+incmbG06C8iOLIZpuIMLD
oMoFBl44Lc/RCmX6VxrSCRBNLZrkWjiXZV4wqujbie2fGAcJO6J7JsGAgWaZqv+5
sm6EE9C6CynNJv8lN8vZaxLYvWJkjNHjuhzF/ATgknn9l+m+t0gY/SgnQKbNann6
v2GROAEi3Wtm0qoAyBTnqFdWTPuNgAHtQm1NY4nQlh6sCVf57826ElDR656pJJta
bAJuNdhtfm+pxuwHDPIJsOYR60zcgMXMY+0tL2qCpitWoLOswll25/UpYUpiMrql
TlsmBRSQwrWYcLY950FlEJeKyRQMC0elGHfpzeqydl9XqkYbYI1qYOkAvQupROl+
jN/FAfhsjAA0+9pBXdSPJKUa/Th7tqQvwq6b08vL1nZtn/PPBDWQc0H47LiqA/7h
psknqMp+Odw55axSDX/idH/bIkj70hpLeGEZJTAgp5Z9Yl5f37u7zNuizfVHP7Gt
0gBW4SGOM9Hb9TDUgYyqJtwUL9uWRsz40lmhMBKxQavQach8boms/u72jFWn8UNL
iQWljS/kE3p8cyo5RpF/9c+1AjQFt5yIebXmxTyZXL7tk+/GuPK6VmKmdEZbxLeV
u7QuM/iWjZDE+r1hdBJM1QIFiOnaJo92E/DjQrt/UcGrbB5TvVViRSYC0IgRSp/x
0iKtMPVE5Rpwzy//hneoMJxvInKjNiJAybzP8ILedqFZIen4PRLH4kujR+1eWcKh
yN3RtMTHHmecaKfzBHnKydLh7LMd3LupkTpkMxlcb0HkS448ks0Yvn+3T13w1T8a
hR0hGLKnD+a0UBr+3664pfWsCGhm0cD54OKQxjojv1Oggu/X6N/NINSWwYZpO8TJ
ZEBnssUa9VbKSn2WtiUWCt9KUD/PhTadCNG1QK06gGPzjewG41TxyCQ1koTdVwMD
XJwmyhKfyL+w8nDr00G7Jk2mazqmDjSkG/NIMxJohdtTfGYL+bZIj92ZrZ8fsrPy
Zr3D3swRyboaoA8MTnYoAJu8SHvrYHRHOQFX95jV+8WN8eZAeUvSmRdSiadvY3wU
/6q+sgmNprNgJFWC0E7V1TAamSVWL6Yw+H8rROwdnr5BoNMpwTWilUJRmpjRHNsg
QpOJBZjhg9TU/p00sviI3sTS/BE2T5NAVfA+IcYJ3aVUr5YcjnCRb5C2qnLoiDzi
/UVE+T1OVpOUYvth/QH3VcSU2IYMgYEj/BRujrnabOz9Wx6aFJ6KSuormOCQ/at0
oXDMuh2exoiTEXOeDeFOp/8EZf4HNmi6ibefN3mRZQm3DUo2qhvxOlG8WoYJmJCb
jRO2EBAHCbpSVszYIj0GXBiloCsrtljHjrgrcCOJad9nP2ZjTVKLIKR/JsKS1NF+
kHMGUS+ky2wv/Vi1Q8WiOGsnpM7EeBS3mIUduAUW6UBHaXyZbvnE/OcwZ77qeZ8t
YWrG/K7CTnaBxEGGrzdQYptshQXHlSSFhpMPHORZ7Zchscp8Lb5XqjKNwaGxO07R
ZMljkAcletGeQtK2fojt8X8lnt7PsY6NNVE3ET2v5md8xmaswXa1LaxZdncnjSnz
eaUEtAMhtJmdcCxrXwmKzKWkLcWwy2OAdQ4G+Y2Zjqx7CZRAYYapatJba9ZsYg3l
klRqwWXv+JiiEpPBXZFr0SfWOtIkojmtLTaFnf8Y7eiWCsif3jJdTHh+UOX3FXFR
/gpKOWXUGnPA4uHdk8ouBEu2X/fv2IB7Qb9CBkTfAbzJOdrXkuhfVDkdLepn/03/
y58sybAE54OBmfszacZ/9oKD7ItioGg5jOQVR2kalj3MwgMHJGn3thm7Gb2Q210m
cW98JBGFKs3s4KEM9VeTlicShHRqV0kIqovtdIssPbouD+6kSx+tMfonnUb9FM6C
mVDH64sXoDTy2qcGcV0J32VUYlWByaIpfuwbaEpr0jP7m+ak2ugR/qTqX0+aTtfI
MVZ/Io8c654wLfbKhOJ28t7Yh7unwuUK9E3TKrxF4PWI3v9L2NPcvfqWknkiZkfX
tHIgULWZircIScglioSWpaObgr9lqO25MD6Bw9WgdV5EpKWHhEqyALJK1+uldajw
f+5U1kHZ0qvo4Pcpcd6QJ3dvMNrIQTbbT+ANqkY2CwbXqxQNX2L1dmuMSXjPUSAZ
h1oMgiqzjWMTCxYfzUZooWtFqJB3K+yKuO73VC6dtdIxtVg5P6lxuaY59maVicYN
UqljNTG9uziSptBFW4DdMqfB8yAOo7+XN9VNaFniPr9Ko4jsCTN6VG8RtjI0pC3s
x5nS0+yZ2GxolhG8pF7ZxqAcYvXlfuIDiA1Z1CoKolgRxM+gwsZs9DtVUMq8vZye
1BjThz3MNg2BNsp35ZYk87kGXpyiQxOW7rKK5jwSjaLUPaOoHt5qWc3o43HUFawZ
w6vOOwQXNuwdb/2KODhr1hCyg1byAQnhM1juc3ClTa30VOVSE1JDQ0OfhkMfkR5I
p2dtMJwSTtE42nQkoR6tqkFPYn3M2PJe/8GoweEhWhZT0sY1j9vOfawKO0JaC1GV
jtpBCDDz9E1dtehKcNzKzcGh3Jzbj1UHZziyMV7em9abXV3sJ5NxYFXbmQSvw0LP
1G0r3etyEErpAxYsz3/7QK2NJ8I8fmBlvydHhnqmOnYYd08BN6qSJNKUF7cO+tqb
ZgI4mv1KvjE4AfFLCh5C7Hz9G2b3AxVllhNYbaBHbGDYN0QDGKmkiOXvugHbA2ef
O1J7E1c+P6mkGzanRTAHA9Gkw9f7TALK4WA3n6V8oa5zRt54tzZy12Tk6fxSmeLY
VXlyKP/5mw301YyBZiFjq5F0sijRtDEeN24FFHFiQlKxbLceiTnoqfJTw+1UKahg
XDr2/0N6iP4GssG3LKkVDBbaPv3hZ9D0UEMFANp4hZ8NahcEumr+Gr5JQWYMUy1V
ci2idRXlBuSUPXicTU6WisyLjwgoSrTbroQXVVbJbGiACLpxg+ym0704oJXlgPLW
FTORuuQfBPdsZRj9Q/ELYtxCywHZm1tVGDxd1ibKJPZM5j3gAtL8w7TPlTvy4rRU
VpEXFGzhCN8GqjviZXdStlFq3p0td0Uoa5PDMTU3s2dLW4gZuAMiEofcp+2vtMJO
gPkpljrydAYkNFtSYGZV44LZQOsa8Sp53CLQ2tp2MjCNTv9KoEjMa1o36jxvUINt
R8d7WAYwRrfdMPFZUupixQsIEBb3ulqAYKZoEGra4kxBlKXVjlFibumOKDX3XmJ8
fwdlZY5qd/SRO1Pa7btPsaTeEkBy4cqw9iqQaydu4vid5I7VjtXoz5IervN+PLLP
dtOAAjKxVNZBY4aALj2D4Mx8uHwxW3BfJOBqzvUBWiwpgdLsA7Gqc+PQIi1vd0ew
OKVqWeqGmHMzBJFNFR6gA+uSgm/viaPhViqxg+ldkIbChSjJkxxx/LaQRoj4a6C4
QXS6aX6M7QCYKyuHoUYHImivybjUiVVkMx32FmBlfzkHe6RI+if7jdjda+LPWchy
nncGhIkkA97jwYcFNoKRfMiHWEqeIlUNMQMIum517yAcrWbQ8O0FPN9plbqHLuw+
pm1VEAtjeb9/UL+4yqVk9dVXPLbdrp7axozOhV54ZNRIRhVYvsfyB44b3Rcl37tr
pcUeI9enEnzvxkAbEhSOMhqDEkb/aqyy+48QcyTnL6C5XaPcA2Qf+DWiBtEkFSX3
9h/URZneVrmxxSiuswsO/BsxOlJZBnuheeWWkd3jC2ZmgackVfnX6dx/8GoJVbg8
j/kSL/LHw85M0mDoX36UW4vas5Tdvq8aS+4PdXU74x++IiESaUP1FwnnAyWb8ElM
Q+i4TnKqo4iNKtxustpu6+fpntrot86p3p64jysgpmw3ydrV8pXXR7UQnQL9TDiD
uIT5SVlXhBso073WN4pO2DFBOCLePUp+sMiBv0LcNCLsfw6G0GGMwwTtBPHGB/Rv
aA71VnUs2bamUZ/VJv6i2pu9of+WugRz8Mf7aFOtSynLn6obLWQc5H6NWw2is7hs
ylyj1e4F0PjLGLQGHeUFIVrKBTg47nSK7o5zgpOXResbUMGBoA85bTZie91Cy1Pf
Lf/BQ7O1fhQucnpAVQY4DOKi/X58CFnAPxN2KTG0gzW6rWtwoJAJ61kBFLIWsA1z
gWYqO560jJXOfi0gyzwkLNkIAaodF8VR5DntjR4C+X31I6mBqBCe+kPHyh1DkCmW
i8Or32NehNJhxmFyieJp8hEYzBaLyFAC3Y3vrfAdwGQvCGPBGlzLEUB+E8pyb9/P
d6AXnuEYt+g5CaS4T3JNa2iJD64caF3/qAmqL4H+hLaE+jWN5HWNRi1FjMoSLk/T
2feVAIgQmMwc2+LUhBSHO6SoAiWC8+Gggk79Uiuyl+NO4FDoOkeGujSSuwFHy9HK
/xfZgfu+c7ZjHa/MBVU0t7+CBVFjWnHhD4stYpRb92nrhKXNfh2/3BnfhjCjmjgC
TibGv9LMqm/i8UhhnLibSMYSHx0wR4J37nRuAJtuEdfXpgWwkBuUU222Vkw6aMcn
8/Dw+v+HGUtGBuV/XpF0TQlqjs6C6j66MX7KEBQ0raR4v7YB/ag038XeS9n935RC
nF8nAxOrKfDSKHmJq59IbPGkPWWRAu7HaEpowgJtsBHiwXdVhPIggM1i5076H+JG
ccACaDtbGssmVEj+GqaTD/4DALkRLCBGWazLpfr1ts0ldwp+boYhzJjg3xzG0fsP
51619ue+eYsfBhvlryP5cMpdS/AelYmmKq+RMMrpsEJuK+vpXcH/z41SNseTh3j/
WYJ6xXkiGLeI3lhSHNnfFdML0bczLHqmeu1LPFcRFSElTfrvKlXxNvBvPmYdfGcQ
UvsciUnyJN+uTIY0tEweQ0TN7yVug2FloURKT1EyE5DI9VQucvjbALiqrtkQtGVk
WO+ZpEl0rF50lUAqFuaZnfCqIEoyDy5lcn1HlpH/xP28iMxuitmXbjmpX3CIgXR/
VxuVS/easUxOC/Q5hZMQbyvxQost+mCgff/TirYYWgKDkuFtQFqJZsWEHp6bOaio
4jJqOVepi3CWvFwuC+Ghg36NWLs8wzURM1IeERzq7MeH5BW0quZx3DLG8N0AqXMY
2eN3/8gwex7facJU72XriX5D+mIxR71jWsEuvwu8wMQA5QcRETSPJVe42EkDeCEl
cQPku/Cw4002/rrwn6kOIkbZpq9pQGe1vKAWtKwSwCh2LtD4MDz8ocAv8zyQjuI+
zCuS6Tg6p3ji3EBYtExK6uB0vlq2rIY2hJG7kT6zwAwrwSBCax8I/fCQCk4tgIO1
WsFnk6Rr2U8e9SXFkPUIbjTdUUfhjwoc3YvkmlteVnEe7yxRZEjPgYh0ujlhJzhr
Wjr0JfYrXd0PEsMVN0LwZpqKDd/b88ACjlOCVMD4xeMxAw+mxQTpZbBc568i/HiV
cFdOa6cTcwK3nKnbdF4jPtviMlOg4EOkJykl4wCm2jwMYiirlZx5PtstYDS/VM+r
iuMLthiR5Jbbez8Ir8tAFfsBxDKOHWjeBMKCcbJUKkrbTfu2uZXMyDVwe2jT0sgv
uOS5kXUeJd5CvcvL5GPcRQfL4RKtgAE+NXSEI15wu4AP5l1Wo2Ckm2Faw4Jh+MVB
LB94RaS83onRoVzvXRhub7aiDK71FztZe/C70uDtaw0d3bEStLILgEtogUaQUVz4
qyJagxZBLq90N+LvpzWNNvVGHMKJCihvs2dVGrkR5X5PP1apedeQCTwrukEeq9y3
tAyV9+WHch+63vsa2V2h3a6j4bLu7TktiXMoJTdSnIDBHnaWRFr5SUUiPa0lYySD
BowzVpKx24pcKMXpRw7nAO3oBHNi8UD/hzxgAitklPZULdrZd7SKcZmwNfxm6HO4
CZMGN14WMmxvrg94CkJycgL19K+01Rh12SwPN9J4IUn7HAjTr+r6EeR0l830lp6g
ah/uR3oxL3+ZRes5Q2dY3Krq/yqjYAo6xNOl2v4hdHd5KU2orIAxt8TYYpB7t81/
oByLzEsNQ90XlrEfut9xHeLYKj35XtFcqaeV3N28q0DXpTOVaHUZizrUuajCSOUO
nlYenQvcWANQQzC4MQEVQTumofYB9xqspxghLxQEHmdRDWBolOI2nslcV00Y3/5C
7d2tBNsoGjxnuX393GV2iltIA8gZu/owSNgJr/PxrGsBQt4PTrSVNUauOVjAh83B
oYiHxTmsbbuA6mCyv3nMZ7mNW71aVF6E68gdZTLz01nGPfHU56rWwHhr+jSsQ+RW
nNd727TSX03ZwlPBbk8jdLSkgvDAz1FkBDKsm0nBwkuZIhYY19tzw/6lEHmUpFiE
7D7RoJbca1Fg6DQxw9q7QaJhS9jxK5jdYdFZrBSDz86TVGR0OHS9uQqvWsAyq+jU
QXiyAbHAeobnUBlQ7A+qenBq7QwdFe7M6b9l19oMPSJArrXIeOkt3O+TQFJARlUb
MJLGTKFkyMLPGCV72qD6/rCKNsUbLTjr1wXSoFWcjzscJxdU2yuLLj6vbtQuMJPD
n/1MFOAeLJmFX1SMm/ejQoFq6pmztdVO4iSyYzlDCDSbxCkvdEzams+bDf9hY/qo
7sKH0CokKaIb34Gk/+m4sd1tYVIGaOYNJ9TocZyMzyGypI7M0ohhnckNpGcUfT6p
yiN5WjFlNO0HZoKZhrWcVmuwV435g+gCKer2xNjO8VqbLZhjhWYjVrhdNRImxdPL
7YmM9w/dijN5ZkhtzNweVdvqnXmFoPhpk8Sp9W+Nao9oFII/4/VoDdof8PUDFzoX
o6iJ1fxhKzVwiMDU0UhWaqG1pACL/tKujyczEg5/GDQavnXNGzMDLIICHslO8QzS
PlqFoUPO6SYvUMt8zkNojCI6GFtuh1kK9oIz/amiJZhLl5zlOjFzH94BIwEZ/WO6
r/mjiqPCRE6ecuMJMh2l0jTnV/pJXgXOrVnkFpy4s628Ml/aopns3xGMf0D6POU6
DiLLhUsgsH088Q5WBAJmO0OSmMlL+qr4WIp1BgAwCtrHbk9u7KV4BBjk95B7thcF
L3K5gnfSX2Cwkuh8aLGe/GXcE6AMBfOSSumBLXmzvZVo/pOXWO+mI+93s35YXq2T
FF77zfJkAaAKz+5Hwh+1Mp/u+T/8r4pJsG5wb1gnVLxypNIsdroPI2rKGwTI/J2d
bTpyDXLy8X36ipVMQFEkQ6FU7rzFgrei147GU75o6jnfKe85WAHwrjqh4qvHoG2M
gyJmRgKwJlRuSVaS76pMGl/OXu4c8QaQufDcGR47TmWBAdXTUbbXbxa7CgOoOdfD
eNZ8aXeeQPsN56yAP+y3VmHfen7bifRKBg4xb9GBAWVLLNwJf40rhwisO3kLrHAs
LgmH8jB+CbEY8qFQKdU3tNCt7PeOzteL0KIVzehzs3ymOtv6UPlx8WVgUswFLPES
mlYg4ESdZ8g0l3GRxQhE+iv9KeXXazZB7fjIzUNV+fPRtkf4cSMNhArMo4jby1hS
84PE0pxXLSFHEYFcpUdlVUvNDLxsAgJ3SOLprl3WkHAWgporESoimzSuLACakOqq
teBzqW+bvh/dMm91RueNvYA7417+VUkNbI761O32TvdcvkoUKgVN+urKaSm7xG/1
+GG4GMLMNaOYgFfm1N/hcZLPjBAMuHmy3xtGrDnwQGTU1jStWixoPn+tgQL8uP/Q
Ru+YTbQc6hb+M45/F1uqaSZYoQHY2bLJcuug0nQ/t6fPXg56LzPakK9nE7YFNF38
mNei+l24cSHnA4vzb91mN3UbpvfS1KihOcg+ByRnA7PZAVQFqWriMRN5c+APXB7K
pflRZqEdFQAf9XxAjfRTQqDiCgKFej/EIo9P///v7AOyjQUkBhEMFogZJspF8FPY
0zhtANAH008kAnvI02Lc2cJo5TDbV6PT+8BsZ9CR6rHKH6B41E5UJqE40iEMPeFh
5DPSvJKk0/ssT3EQgC32wmo/nXGRSqdOPkNBz1uwTDjtYDn+BPCMppUSZ4btTO+r
SejWrB+hEWl8nnavfx/n6y3bAA1hx1wEnivF428K/Gel9+dKbqnQC7Rlxa37yEpv
NQrtaei6PaBnXUmjy+WUCC1//VdAkjtL+t+Ojtp7V9ug62dZyn5j9doWMOTxUx3u
LFV13sPvkrxVmeNb0q7UhUbP9M+3leb2A1yXMaQcs7cjqqmsm7xoNSAbhzxvTGaj
1MflPCFJ4zGOBbQYk8F+g6xjE3oGvqGCz3S6CaZvM9igc/vhLPokap5ukdGnHoTB
tuaDTJqT2BJbQOLAIxDOMo7txAk+DgF1DgSeSh9rXW4OjxFMMY7JMO8Km+VJZ/RN
SeDYeTHBMBV+KvbCo6RKDbbvAHT5PIgJxdN1Gleyy6wrR4BQft9EjZ7GIWz1rk5U
gk10IIEYaE/Od3dwyzG/Wgki4hUVxo+IZJbrWo1f2Rf1YBSTTFK27+yfhErSioNM
EQWlnPQzSrKKKmAgyZvz+wJMCgqO1Iwq0pY5q6yttabQ17Z+QzmdX+SLYIeB9Ck/
BunqJy1U82abZIGL1aXhSzr50FnUihPkQJVchy+ZjLhPRgcOUteS/yNDjaJfqwQU
gNHP+UvblOaG3XwRzTGpdwPoSTNUHS3WhPNPVCzKl5YLwOkUgFkOwbhM+1Ki9QnJ
eNCpJco3sMDm/GSnL3M8gkKte1Z3GmEGigh/EXih6EwB+SIxHKEWnbUh9bOOKEvn
mcStapYyeJeSzEkCqb5c3P3PJnzJJ4HRcj0L2HXeL9pm0eeLrcCCHq0xlFrSPTIf
i/R1IEyCFboMWeqqwpzxsoDM4sv9D7syc3i9fYBTm34Y6WaRSmNeVIdaHz8mWydv
p7oL9Lufkv+vEIVzfSFn3DJ2YeyTQ+k3VfIQcWN70u8tzal/ps2FRkFbtddviI2f
p9HRNclVn/SE9mSwUe7vkybN2n86RXo6eShDnqGvOs8q/tnRcCSprx6WqTKv2Gyi
nPfuP161tRX9fSXvy8kf3VkKKQZhO2YTv4jQa2kJenSiNAaxqfTsjcplatiBFvHR
ItWEa6RXkqIy1aTiyKnAohnVMZ/U8D53R++rEjV08CcZP1cVUvp30E0jb2WqgC6C
A8qXsGCyyxvtNyAenNhBaP+gw4eiQdoOuhXrr25EGRJvlD6WnP+OSUOM4j5ZCbXu
S9GtxEIEPabQmuIyhqCYYeJ37+NZHB3Yq5TISLSUwNGNFqvCj2sGy58Xjvx/mAo5
Oo7jyHGtSxybOfaLVtJgZvTygtkMgWN7y5Sse09q2PWGEuJagrIVlT38lCxMLoAY
B8bv3WcFlD3RBxXKVo3XkLyhvE9Lb3+wS+qXkBtGC20FtEJJ49tmFHotqBtAbeg0
g0dxpzTYcMrL90E8MEgQegqJpb6ug7cfh+UZu5lrUeNu8r39GMiU5GLcIRvt8zCf
4zA5ccCc/4sIsSf8H3zGEQqOxpPyhXDY8BY06sbVG5O37CNkRNZQ5gUMVup4M7J/
PClQ44jb0wYqrK7Mbb7hIDhp1JsXgZKkyS+MCRK6kr2mqnUhIwPYr4nlLzBNb/sH
LBnixt8fK9eRcnNngQy2nJM+Reh7MFu6P+WzkcmbvZtTxGNlAdcA2LQwYYImYu/s
Td00qf418G/G7RigIkcGx1Ms2lHeGwynzZzbZ4/1UgP5trgA/EnlyCM/TY7wFozQ
FKYhEFwavqGP3x7BMKK+wtHM20iGGHwF8QbSdvDFxy3lepbB581VH7RZiCrLvBV+
cZjyT5f/PtbOq2+voNTtJ56gSE2earVXx3f3XrXWBFnXi6920GjvTR1o5YcbSKlt
hAAKj0drN4dnTugenh2RLkmEM56SJmhnfvqbiAFKvnP6Wxo4rTjhThm3CM2L4FGe
fPEiO27TGUDYO98s6L8P117Uhs1H1hfDBSJFdWFpMOy/tC6FRt3XbWWqbtBS7ogR
4nb8fjL1IrCLXaGw2FYVB1Wm14Mbe4mElchHV7hI93CTU2s6Mp15nZPO/38UeEae
ddiJD5uZ5SHtbP0EZMg8CgK64W7o15Fcti0rZ4OpItIRBKiI6jWeoOiPzCpLy1r3
+Vvto/8hlYjuHkAy7Z9dPRXD08V5GLljbNXfvDPC/yZtyOpK7VsWY3Trewi5LGlz
TtnHytundTH11oWx7Gdlqn1HI0kiL9wswjrIOK70GBAe2aiv7IXXSQpZ1nfm+5XV
5+e/CwoUEkFSi8CHXcT3nX+Y2uE3DbxsQeNbbwEsYMqF2dCThkolRiX2baFxfzki
dx607jWceMIwSrQaddSNdW44e/pgxxHn9akUiOEv+KfOfqglQJ++5IBybJbUulfy
m2MlgNBZvmf1Bf+lADLDfnyU3V1/T5yEMZGRzFfuaMOd3LrGzxKzkn0jgZKbhGVM
2RHQ1qLavUXsvQJ6fe2TwQ+Xlel5yvraCLyxQ0DBD2G/p9vIOKi1dOz/PEpTn7t/
1TlosBNSmSb2QOw9keej9a0ECfVtpjAK3YbFG6elUcZo6oalZPnigHJ5OxD9ZEdC
zGhXV0dLHhslwxrPII2ec2vtwOrCyx3LEyh75WZcP/7fcALI2Z8xXCRV6RjJ1bhl
NTTKZ5IFP8YxAlFXUyXfQSTimhKOmplXgai43Ix9s5oxf5EUhjYwzqqimzVMqEYY
2QEO5ZBNM4e0TtkXVrHYZ/LbyvDfR6efiPaGyoJM6FHmapArqirrsDAyOqqqN3pA
Z4cKNp38Ca7E8ilPzAZp/sb15ElPIlvBbjnpwPxOxi0Zeio5su9LiRGe/iDWvbLB
Ouwnu5L9+xGRrfEy2W4vP2ovYqOIGw3kUts0qP/DepaBsA9t7cHWXXPmqE8CA8Sf
LvsnrIGP++hKi2yOcgsldHTglY/2ETTVvDdDcl+DHJf3e5WJCR1Z9F/FHgfhAd2J
eeI3bRiQYdyIo5KjqGdKmY4MNBbo1nldOXpQeZu9PaQ0DFbEbChLWfByRLRaIQNk
R7o3UMSr923sNlWI9QV7bwcxRBrbEOCtoRJa1s4pwdmZj5ZaVqIW1BLcGpk3N6zY
iS/D4TOHBQ7gsoWtyjUoC1d0mcxPOmmht3sjr2wahpXDbMtkm+b7PtA+zuXc13rQ
o1sKUhl7rq34LSofU/ahF8xwaqDbaPPL4RKCxSxPhiHNKdZ6TWSDUOyYf2GqlM22
rg5kyBDJNqZwpGYUgrpgoJrK4Nte+YORcqlVIupFv1MSafiJXKdQuemN/pWkLduT
7uXgkFOBPT/cDlhbjvQuQnUqP5moqm9kliwY0v4STEgQVPlWovklwhMa8v1iH6ZG
l4djxzgwptcXq6tIo5NpPQVLm9dmsf9UeH+QvxHtvVJ5dosShKpQ3utdeT+1d1qJ
9P8vcfYl+nRNmQvvKzv/QwxGH7XpYDsZ0G38NZ5cZDyJEDtjNs8MF5cUaiqhF/Ak
/kJgONCj951IjmXw5PKmLUhHqCIdvfX6Sso42ZOzX0eyHAs+B2IYa3Gl5gsy4WAD
gsY9aCGo8k7Hf7uiaiuCbjD12n9a1WHNX5/uuo7IVzmDAhWu1lzz5+v/pAV2tPCG
j+tO7L+a4SzQF7s1MFRrBRqQfpfTpvHQogD48Ju6+Eb56l2WflHpRaQHpC6MhHRE
zOuE0/rjk9zglPO9CtozaETFAgmVvAWTDLZ5LX24eFPaSJup1HLHJsRXgAtLbDJC
DXPcwgD6b25Fk17TkHO5YURYar4wRmlkXcbukL9ijYrRhHWm1ZqpKN/nsLRCTK3k
RqG68mQzJJZuUYT2MArU7auQR9iJ18Cv/3hABFuJ2WoVl3MrV6BMt3YLCZ4XfUtP
kCnd/nAXn/crWBWawv4B5ZBIP56PZE0gZvK4ARIHlLLdA7yzxKPwVJ0gpXBmZ960
1WaIHmRQguRLddweLbaSrc1mcyvA0d1Ia7x2zfHwdJsn7RJOIVywHGw0xSkOfKx7
6bFD1sFAhSaTk3HFLS3L8RRf45t89q7Ot7KkmZveUnmaiLmtKKNI34/NBx3YqEKC
zuA/1CQhgvuq/30h/VISzDdmBLQv8lnZzH64CthJlo9ipRQVTg1PBVieQqfMy5+B
gf2tkb6YXXTJ9f/LIh0f8VF8st3JwVtX46j+qZ2ouIDbXG/kplAOah6gSnsrY/8l
K6EfZT4Fc3MmJ58/ehPZ9e7yKzO/Gpccsn9oYtPkyA5o717b94G677h2e4sPsfM7
KYR1uYWBa0+lvOWTfIeZjHqAKiEZ3NIqBy6SJ40i4+NYcOZqqvS/fsGNKD0PCST2
s2KdXb6zGccRQgA0bGWJ5pETrH3xIEf8xUPZXvyhZ5nIB/AV4VPr5EcCDCsrTJ5o
StbbmIIDsWxawoNhAY5jbcGbLkOZYQGHPSVlUzWYz1sjYIxCcWyUTSbriYxlAu9F
6aa8gqrwT+x/oqrncW6eC6EQRcXPWWflxNF9b8o82oOAmbfCYwZq2MRTJ8NlE/2C
CKhmzNnD+4+2wcXgyymL4yS+y51yM7zaaD5m4N1d1HZVdZ5mMy52MMYi1Ddrh8PI
G7JVV7tKc0p7If8NP97c9jiXdald2NltmdexrGGrtomeN+46OMYaOymGMGcctwVQ
24fI6DewDxxLv9JyHPt3PEKySU/2c+fUi7tOsnT2eOH4+XYsTes8CkVG0IQ4dJ2m
8csnEIypd3GR4DUJWgYSJqXNP3Ou7T76qs2dbxFQmzMSoeabHsHfx7nblwoqWhcQ
ZcWRY8pobiDky6opbm3FRZoLY6EAvlO6WQzgWA3XehdZlNcjFTPOvU730qFKpDuj
kazJPj+mODJO3InYzduCch/hmU8tv/qMa5i2g1uTTsa/oU4ieMo63LZSv0a7WmSu
Bn1i3RdoI2GrzfxBVj5u/xIO+sdZqWJjnD9BAqbIImaNs+5Uw7+KgSZsoK90UrO9
G03j3AwDqiD+VIfVthOkAVoG6N6ltZcnZ9AxTb9fUVCCVuqNfBiA4d79FfHPov+Z
d2AQqymujiEr+8kFi9pvFXzgjgKxafEELqUJ9wYlYIQlLwIZOQIB/FBfdDY/fYr7
VVXVe/zWWzw2gbfEqeJFV16jfWFXkEqbrnIwaMxHeS2sumD7m/w/eIsyVssTQ55h
1rrLos1J/gALBz/dn+9twK9+WQomBG34VaPtKopV01qOaYk8TVHvb06nriNwCRFC
IS/eG8zt9ZO3D3vM79XlvREPMHm/BoBfX939FiOKcyZKXKXvqhQ4yn3YVXz9YDDR
O/xSF8yqMi6DoyBZEuCXbbb73mYeQUZK1T+2FRuKbQH71PkAoq/Mx6IULxjjJN8M
+Og+dsMkvpyUoHA7N5fUtM++1kqIwm6ib8WNAMoonlldpP/meE3wgu56xD438cyI
8QD0g/ypiBS39Vf4el5EaYIuYIP5MSaPdLy6DNsSzr2OLaLRn+04qynaKLvwfn9+
l3G3PgG56HDbMCNtMVS9YfzyVE4BwyhFeBxtwDRTm8BUOfDWIeIVphASBZF67oAe
ICojVBmWizdG/EwuuxRSwkRq8nzHVhloE6Ipftr9/nDstO4p60mEj5HUKVvs9DVv
GFeo6Elk2Nr1dwDPACWgIpH/jUeQjgfqo9uOuw3qgcch4BEcw3YKtTJoOW8C/Ksk
EsxT4s9rg/BPa0B2LMtepKcb9tiuXNM0mVSRHqoUvTd6BT3mmwSGdClcusLPYmXJ
3BokTQGNqaSv1WDQR0kyCXC5tQu7La6V6NgsfJb+G38KnK0QmWui7T+AHsYilFGX
dZSRYhnBbtvOCNMK3/gKcaugI5puZjWvCyZXvRaVP2dlss3TJnfCELUjZIOpeklP
86nIMC/48cL85M/HvhbrUUpyA0WRn1l/OqXrBiJLNfefKtEpRYugbqJlT6Yr8p6S
YZ8/HlxOCd4EyEJxMeAr+nYkAkfPnuKIwssKXI+gwIf0D4exijs4Hrr78pmzWXUx
c/AoDW7iq8L5ojRItuxuO6Icg+1tj9uUHzZaxumkw1lDQ8NlkEPQYpvTfSzAFziS
xNoKBhG87fhQQShF5/Z2usfOFyKPtYhQ6UlKRdYOJLDJ98Sr8QPvtgx2LgsyNNLT
svt4kshjoNSuOOWWAV7pCNk6XJOf3tWV5jVPV+KEH0yDWn2nFzbxi/V5kYLdQDeC
J0QpVcg6sbARQ1gCaI6+NQsaJI27s2oqSsicVTBSXbmBv6D+9dtDHS22MqX3fR0g
FB2+kW7EN7/HeXuX7du0u8CMr/rA2cdQSK9DQ14XUkR27BFk3WGYJslRoEmrT1aQ
KS6km3N+DsOWFxmpvgPIlp422F5iP4cqdWu2ZpeOrFIX5XcXJowXq8WfWy0EpQkT
cIQkT26ljrhRyTaIO5JK/0v0Yj7AoHSYStxtLnBVurSkH/yp8rIUi8EEtueJr8X2
KSmGfKoDU44LgjLjZELGsj/lWhYjpNEFHUjYJuvj2ttWMl5AG8vQknMVbAZknU/m
VBFCiT8YyWElJ/P+N2gmC9ycv4NpOZW6WqdUkuvQansocVodb1Nw+slMXQ6FUXfu
alNr2IgN7jdvFnCpCLPKtsDqAvSmJBKhOqBZJ94L0QQPxcMVisp7tvzUM4zm8Gxj
zE1yvHSvgd0pZ8PXyJpqDVvBU7PtqYLrLe5veUgvImuc8PNFiAA+SWEmzc/feVlr
RWn4vipZ3KdaXPoE718of6sXcdOKeCYRdDVn7aocIG5wudyXQ1ypyG2qqWezA3UW
43Yhwn7VJh0I9rqrVcjumjqKa8pYSr5ZvKUUIZem3hVRsAxYj1oxSK2jApRjNAlR
9eKHFiUQMcF9/hzVik7WPNTRJglyWAi9VodIig0l6AYRlIORPXNXcxHoGrIj280O
NiOmUAydTgtucDlfrKGpBXHkeK38BEv14N7yYAaTCSo02HCiDc0+krmvPuiiuINJ
QBcdlg+MuArUlYsxw5V+cx1KpDIV8uid45rDn8wL3yDFviwhZtzftj8nTDESuTOI
i69E6CI97d749l79x6lnvJGtiZvi7bbGi+OY7EOnQPzWN/heZy8HBsbdyRn3VHQY
N3o9obRF/hNmXERYBg/myuySJDM+oK3gDNQvvY1cE9PYKORRtABD/uARgBedL9wu
mKsuhndWQ/2OiKkUybXkBOGlxVEwZWfala5DCl/WQhazRqju1Z5T1f0BCKQt524S
ONeUBI3tleV63IQvVP7vCG9qbpBiGiDzhyKqugaMpxT5W6kFcyXJ4Twbi/95IvpK
ofEwq0XFNSz3FflTwKyJF6BWzHgMsSC+d0PNJ6pclv1hzvWvaLVX2uFoWIBswNH3
B86R1caVZfPY4hob6TD+0lToLZu033ejduBJ+4sh8NeLDKTV2M0ZPegYHdAO5oa7
rIAO5IifWHIeajPBpKLtWgZrKlkgHUeUZlJg9xz2ixU30DwbHSaK5h+tFrmZ1GpO
cxezIbEzoK3HMxTp+z8FSXYGI7jnZhZUcNhreBaSsILw1I+OinZV9XcccSOIwMDW
fdCbH9nF5jg1WWi0WSbiFe7hyWdUyM7Y7Ecs+/3QALd5NYaRuAX9fsvM2+bpk7mF
+4rr80bL5h9jPuMZRBrO31V9garvnKJaJWTcA0i/Ov3skW+ZsUcIUjjQy4pMSLVO
mr/qgdHWtzD2kY8WtFconbJ2gNFVagH/qsN7inHy12Yl1kFBj0pJzWWf0vpkJjRN
pQrG454jeeear9KCvNWGkBwDq49BmozIJ5Aex9YNQmc+1+6/fhCZIeZ7oNsTI8aP
gsJJDs2w79RNVC7IJl3zIiTvcGIzmSSCuCyyjiY8kij0+UVh3RLzEk+tvVmGElfM
tKkLrjTHc2ayQzlshF+u3Ay7EyptJR4ihXiRNZm0/9VBQOuMR/E5+Xxu0XGrMB+E
pG8VtikaCX7OQEcVlDx1cUrNj4P2Nm/RXxVmrMZC/ASVAdUxslpMQY7hfQwNDCkI
/Kf/O4yBu3sZoIgJcRHJC6nFfy7c81+9K/IPCwLD7PMpRemed2K9jbeJNnwE1Ywa
F1nGhlVmT9m0SgIuOXYGNe8SSDo6ZbDbETI6AT1GuN3NeAqp2P5pr5QUi+IrbtU1
fToMw7EPYFXWEcV/O2YtSsXS179TV7+4Yp0TqogUKckuQSHqMun9Hq5q95rxhivl
iBZe+e+sckrZxI5mOT1eaLTHU59dEgkO+R/OPw5qTMNOWqOfzqMxZTX7ulSu3Wm7
39KhkQPOQ26DIaHOM6fiZXlAPfvXkORXOQ1NsB83F7v+B1LaAt311K//ai5GKw5d
HOv0d0QdiAD2GERfg5Pw4uAWKtXE9IpDEbdwnKHiQO6z48FP2j3nxnJw+S+HtmVq
Yd+/xuAJ2gwGzP+D18/8l3o+s5lf228J/VIkH8cXdWniItWO2ZpuFT1IOL7+9ML0
A+xzUhLPmlduSEjhyidsAWI8vAO0ZstxA/C3d35S1nZmpiTf4GYiABmgUpvaRaRV
jRGpZB7yilsjjpFOUaQLk+LYpXqe3xyZEI1n45nI4s1+kY19EWh7pflu9mzCs3+i
cEh6uchN4PRqAAaezi6ja5OOMqnkYpz/UkxVJ6XdIXupJfVj8X/8z5G83yByBxui
GaXf4zRoJ96FM6PlJjIpyqzPSRD/tVbzU31osqIOHV6MmgUpjHreVRutBpOpTM/m
82AhCc430VbGLDGAA8AGLq8vS4ZROciBzst2NT8SMFh9qSjdXMNROU/vmdquA/zw
zhybfsNZERSqhRHgBuldV4C5YKieTsptVWEv97/YQqD0Lg6ISFLfl1Zg+e9BD/I2
ofXM1+tt+L6rhF/B6O0WOlDDEdRQVPH6mgzpPc1YPt7TX2pVdWhLvUoeygcBYkUA
qgM+4br8GCBGVP9oTg6sr56iMh4X9USROCVc23Ejzs1jlhGjbcU4wYZ1C5OBH+2E
OLE0ZlXTqSzIZFEZlZqD850shml3fiMJVRGkF/8ZpT4Vbr6PEHErrZAS1cHDUV0U
4FA1fy45BX9b1M6ib34vD3WX+2KfTuYJ5Vd3X8EuR4+RVQBmpMw10yWJHiLhTCZx
VO/20CGkhEZHgkNUk1MXq7JowjFXZmL8Qx2JuO4ECkedLDLkoKv+3jdLbqQUO5+u
dY1i8zJDQdHg4HejJ46O/wWDz+GC87Gxy8MfQpoEwKpoBJnO7J/e9hLn6xMTjAFb
YN4c2K4bEPf9VYMoW7Gxf6PPLs+uro01JltwdSR9R/opAIi1+z3+CkpnlHmW0ZHh
lDigACFyIU7G5iGM0unJXRRFJH0mmaohQ6BRLUz5r6R5vZpVZOIwHEJGYiXFiM5k
EKUoXQQAPdl9uV3e6r9D1w97uFfMfXPEDLBxXmOM1qgAFTqPzsh1a0z7g5FefyGo
iYmNnEM2P3aLUlZHvVYSQKapMQwCFo8uICAftTAevXpc/159uVd9T40CCXndIdh7
mou/QxepNPH8rRILIKB2nefzc2gr2IdBUYBI2R+CONqxIALwtakGBeup7OTDHe+P
vGWXYm6W61ts/vDM3NDTeiHhP40xiaqErWptyEqSxH0xbow97IuxwcRnvb2FfyfX
VWFasjLHY0/F+k/eHvbJyzmGYpYloREMShIKJ0ET6mWdqb3jxZdgLu4DFLXjaAqw
Y/EXY4aGjbAte0hkV/NXsuEb5baXMMHGOM+1I6/0PJcHVdHn5ci3x2HvJBPMGp+P
OAwy7hsyCMciGLHeDFRMm1HDHBZI9aVn932OFprSs85eLCq3lcHJu5GbXf4O9Ua7
kelyL3spc+FyHjYVrUO6okp25Qkqp0EUZJjSO4YEaLB0jxre8eEZF0KqNkZzubiH
3W1BJHVvsZ/FtUq8dmJQDeVgQ6f3sSUQKD0nkewl1OmRsrAZBwRfZL4lJqHLmgBD
mvsnK+ulTnhiLrmTkohZCe6TYWIUE0730g2uJtFjjXcrMhdwqNe/axU5R1ZWbkoS
qYM/4qOslpB6Gm0Z0Mcz53T3p91nzDU5NdlxbJpH0GK6YdhJclDI/X/jTUGGInzO
drygFHGA3iRWeA3L1slAunm/QIxkUNMi9U0VAdoRuJjcfFL9zitwZaed5y9i+RbG
skP+DQemk37AzGmFbAc9fqCLTsm3Ccux254/1BM6Wnm1qVKFJsHuR5uYByjswWE7
Xrz5gq2gwsYk4g0gWr6Iq3sHjKDxpryhwT98kcSeCJVznYCBgPSvfK0iFoctw75q
n3ha/IY5D5TtcrWrxCeUUIqDKFRGPlcRyX84iWZDnPWK+mKvvYRaLgsZGzi2wPy8
iwadvgiGbO19GkDtNp1mu09i2xZQqYHM3IjnEBgfnniUyVeR7BbUcRIFA+nJUz/L
upI9e/BgVvKxwtNNLEwsPJzbhM/Lva/QCszDSQLBqPEikc2H6yyg7kazJl81xm+y
+OhqcMGo+3asaRuRjP/35+O4rek6Q84O7ICgcKV2wFvyvyD0yNBTZbVQ8V85QklZ
p6oV1nu865sbrhAW9177tJdas00gc7TChfJmyYljo6mAcT+XYFg4o2cocuFXdPzj
3nhPonO8DvePJh+HPuS1Omwn1qU0v9fMHLxPbyMfUbFilzLUBeYE5z47ve5nTCRK
w6m8JvsIZfzIaDIdBUcVknDqFPMTbEo1Ov8AmHE3lIvxAEj485rOZBlvDuWvOLq2
BvukJjfEQ/Ayl1Xx+ndeUzw3wZrSTXv8+A8t5xtzbmR8MoxYnjsFyxk9ikHXHG/w
x9Ixnp1jNMUBZkLNtgXEb30purAU7vDVqoJtYNPhyUn1VIyvRxefAuZ0Pk1Aw3Ph
zy4yLgFW7nGycIB07jgbv0Tf3BcSOBCF+vsyNMxN5uTfNrEs7S2uuOQT6yV3C66A
8V3FmSqggswH6aJPTzpbvcKjNjhUyzHYLZInhJbn6fCd5BnR3gfEk4A5OrbOgz38
3hz88/iTmqQHn16tJaxwLVnO2veTJeE+WYnuQbn9fTbx8HXCq6itJ49M3QPClbeA
MdKlXf0jYaAdcegit1Rk1Zo9rH/BoZEnTSo70mZMQY6CHs36fnlMlD1QDLShit7f
ytCpg+me/3bBNfJ+bZaU4A1U+0DTw8+3dAgSszhF3mmI3QSp5GGbrzSKZXXDI3eQ
LCemDw70kdCwDMEG7fQsSXQlDV7lhfot5jzYk5IT2+y/kzy2/BZNL2O1kSpSPjce
vRvRDMCFwaYGu+aelkkEsazeYxx73OpS/nMTilLpS0ZJ8kGhhvlfh0nqMsP52WfQ
NLhofmuzePHYw8SP65GGt/bM14COMVP4HaNQuJUTvHvOj+QiWsu1kTOONd0FnVav
vJ/QFrFTQLTdvbekbG7p1T4TKkPNiuAXXIhyljXknZxce1HSTWaUSG8+FyTMt3wm
97fc0zqIUeu2drDDI3jrebolDa3+Ao3AZntj4V7wjESpUgui4F7nmG8eqeu241BC
AZ7faOBkz4bOMwuUWhQK2qbUEgnYyAPFkP6qLCtq2fWOEYqqbY7GfpAVuoDAuPk7
Xiv3wSRIE5dKffCft7byuW/DrvErZlrfE6OZeuNIGk9sYwVajl9Jfjf9OdI40B8V
YLz1B+TMZO2chWa5Nc+s9l200ZZc5AKmNBuFDquP0NC1gBT++kE+S6lFNMZtkfZA
hRr+cFHk+0YMU2QPHSW6csspSQLABEHF5dYM6g1XPj2BahuLXpJA8+qKY5jmpq7G
8wGBPLMrPWtkoyucLCd/z12MYTi9jV0avjzKPImWdsgNHmP9KxJlpcrQv+hTWyvV
ePr9CWwkT9ptk4TUyHHYJZ881qSV56fCzePPX7Kay8+sTNjhpQka7hfILpsSI1Z8
Jd8+NIBOt8UriBgj8q35QenVtaK+EVuycZapUr/mQCpTbAz+Dboami4bClMdAwWL
np+2uOdPtM8U7IbPRQXHNXmFnQpJ3uih2lvlyuztshmcMXnGRw53Wpo/Eglg3g3Y
WspL4GSViAPZ+eNzXKbzZ0MpYrtI4/1FH8gQaiIQPMN80kkA0I1Rd4jTI3+QoQAO
DewOIEEGarU/OO4jKW4iBKphogFTRX9fBZ3EFofk779iGlFH3rp+1nbTT83TxGa8
BwfUltIGxMbICN28LDcBGpThtJ5uU+ZpPpUePzywCmr1/j6oqB9E6+7RQ+/t4ueH
pNTH5doMff2cCr3u8c4RLNBZTEhGhLMedkUp3sNJ5VEYapFc6MyWGzUHQnhVFVMQ
LDWNxOsnH4H8Ls73TAk6RDU9tRpBlUfjXy77q1JUuuQzZewrXijsfrvV54m+JFxN
6hCR1ZuIcjmkMZZpLFNF1zbdRcJ2RR0pU86oCwJO6JZQVfOIYsYHscN08YUlc4bb
pERyafP24pYd4B/OaflRjyGDvs2hMA4c/TlXZ08NGEQORxMbuwvFzsa0ZrxqeX9N
gpxzsrNbPhpVW/RnVWjOf3afkF2har+tyKMy+62mwNR9ad+J2nztrioZlujZtNrC
PWSGX+sJSvH5mxUhIXfXJZnbUrZMLOEyhmS0r0TIe3DEQjIxTtzILDwGRKM06tc5
zNBpU+fIgJlayUDiqJ/kJdmRWwLaucRgb0EhrfPAVLovSKlnxw74nebxBo0W8g+8
UJ8AngrHPtZEtJPc+Ex0nsT9iuamtDJBcmuHOwZmpbsT5VZNuvmV49ihYO7IdGyP
x4v2JzdjdbwijOo03zABkJcCM2SCmonDCs/GpHHuI3DVT6yvCAD+pHfFB2dw36X6
jDyfJ4xfMDipmKe9jAC/t+hQvTG6dXtw0dGsWzDSLjlaiyPWT/vbZSQpmoYTXNip
ZJ3/ZNXCdMUD8kuuHxAwbAuxUsJXSu9qHaip6muMKGf8SCvVDLNpXZ5W0VRiua1i
xW3XYbxjlZL1a8CHpBcLhVprpHpcmFCWM71zSTz43VBi/TIuJtZlb5pMNtTGTJkJ
qOBLyp6BmjDUNMgXhGQaCXvey88hMQZlBPEMIuXTfPXBZ5wtJTQwoBJ67TsYGCuY
LXHny/qVlMU+o+8/EVPY3DLzSbZUxIdyexPtuBN71Jvh3P2sm4u1nGJGSfYEWNsM
XhvefWWfdcjdEtDeDLfpqqqZJPDV30iN6j7LCB8tNCDmVO3jVyHm5X4PFQo/IUdW
Nvxoi3Tr0t57CMpYoe2TKX1ra9jjm1O5LjarBx1YAQo0AE27Fnk2ASuNyQaQ6f0q
VOuOJv+kdBdokM2qLOolPNF4sboUcz11afojKMwyMVApWzISOt5NrW2vTiZHXhzB
BQRcMXEe73XVtqjzklk1mX+YlGKx80n+ccgN+wcSjwMEvi7mnjjiYPYxaP4VPZpZ
lk4Y0mX88SQhfRIQjWZX8T24Q3LtL7WVFm9UegNh+vuA8WgNXcyqiYgErwdgu0Z5
/mMf3GbphQDYEUcObiaZV60mqxyxx3U7CNX/zwWemxmAOwrlmJNLcVzg20mMhFSk
qj7X6StFhtCGnU5NX9vX9ftn2ofWCrP30VF8coJSfI3UsJeRNEdV83vwtSUO8rAr
A23DeXkp3jSDn5M72W2KnE0QJFS31vIvjkGz8vhQed7YU/0K79QXyhu94ANK9ryM
5B9smvrHfgLfSCfGiIZOmVnHuDueBfpMAjMMOuQ0mBu0TL6yGcJdSTtyiY9UaTPF
OUv2BSJNqjC8laXvjzZAZXEQqQ13V4NYnJsCNNBjLhDpVgMXJY+k/68yTL653S6l
PfSpFpuwJp6PgnXrhjlFxPDA4OMMI1laq21NT96437qmy8isluO1WbGxxFGfcDx7
GYDEQEudEX15d8B5EVWnW6DfUr3XmMpkrBqmAOcgUrU25oG3JlPrHBx3BEh1rfGQ
laF2sGijl+/D2tqcz6dxGTJwQQ4MtyedTnBNUPRrIy/e1h0BBL7XkepgZRxwKOkk
6RfG8JD4IWpu8QvvfP2LZDtEUzz4+3fvNdzWkGuiemyPM8iCsFEqQsFVmeK/Gqop
6pX5znth8aDHJ+eRUrAqynrXtf9s1vVKDHXFJSEDaR7fpVZ1VhqIs71lJI9H8gbH
wfWEciLegSkfODggtJwj7P4LWqY1etJsHPCcEKuv5a0Uec63iuxnYWnBXdETsMjD
mK7QwN5QbKQclhbzvqfbhpszLHUxiEK2tABauD0s7UkhRkN4L1KN4x7KMBa3qJoq
mCkKlk5apC57hQ88acp/MKKskfdMgZvkgmmLeE9VLzHtiCEYnm08sqxq62LnYdGR
9D84lJiH537Mqv3hOnXjqtTbQ3DyyismG+kVeStKCWcNpzICZmkrVLn8iOxFo3XL
0AdNXacROtUCPJAdQhZ98UARJFvMUHQX4M93W8iK7OwC8SCurtBMVEFDUBcCRtYv
nPcUbx6sgVf++U0wGQgMzQ+x6xIXIbAm+IHISi5k33XRz62nU3iEve58+LwOwAsL
oEnmBX/R/3OmeUuuYmOVCos40RqubmHx2YG3sOvNxBNWlMWGON8eJT/7I+yo0oFb
Miu3JqfGlUe6Yn0/Pvlwxt/hE0t6FezbmsM/uWKQlY+KA57ngIb0eExdHjH3e1tE
a/p6elhKDYyaWwjmaVbFSNEEBYde3gQzBCjcdsp4YEzbxc/3HXEYDHp6rCYPtcaO
mnsAUAOTKCbaZvkrAwPTFaoFBZc6pXmVPbS2ALsQNCTuy1FPVz5wMZdyrMTULkKy
YZNvI2FrbDYqMWx+WAatuOiQcrxb2lwH7IW05vuHxv767RcAERGcfKt15ijfoJUB
wgdGtDQhyNUVcyjgVKE8nXlytHswlm1MmUK5QJ79kD4oaPDYmS8/UuIUwgeQtGZ5
GvmYP31KdOi/fgfBNmY/xTV13fUDcMRXFFKZ7hlowKr5hsk/I7ObEQ//TpVSSiNk
DU7PPYfkgj1yyx3aD6gkHku/2vEPRvW0imqZwmOiA63C+D6iZldhiQQlF8ZqZx27
kXhq6279UcTU5FQWCh3V6njOs3Objv088Xrj5wMbnkb0D0099YXPE4sx4YBhUgK7
fEO6JBN525tbrxMGf/vkp4pA8EIqBCJG1l0ZyxgQw4YSoSsYTBzzaBEjAt2VUxO0
61NzBbGTkyl+ANqThpZpF8hwtMV2xiOTbJkzRUYoI2Vi01QalwUXtA3QdltLlfsW
ZxC8m3C/bOjgM12dk0TsVrMGZKfL/VwAZ8Vw7ujc5yxemOLzF02pgj2dqM/NhNtv
p57wtybOkQ9e/AqZQ4G2P8CNtVsGIzPrRhP0Ff0SLS4aokL/Ke+CeCBO9VAPCqNb
tOkHuTbhhqkT6mEp1z2TCqSLyawnbb/N1k9WJxx4BmUWg2UbonfPmQM7HhUdnjgs
q/tfDlhg9PrVfqfBKcnd3Hg0EDMAYL/b40OiFw2UcpLk9B4lq4TedBFIF7ns3uzN
NQ70jbTZ7moiSKZd8klaIcacgflLiExtaabdglLCsuLfEyvYBm6MmzJsCO/0WCsv
lQEhqQp0slFHswIS4wvfAE7h5cJEJf8KvKnF042V8fBoy0xiBpPYQXyac6JlDcW7
U2dDA8oh3pXqWYAkmG1uxQUyvy4qC6+hOEHjP5KirwPqaCc12ZI3fsQcCpBtxqeM
VOR3W9NIsDRjV5d2HMLP8fDipjNFyBmOUTEuQ0dbjbIU+hYtjtHShyjeHtzLVuE0
vN8ik6nigXAn1WOxICSyXYc2uXhj24TluQR1Md7AXUX/JyYLmXS1Iwsw2nfKiCtc
3wmRls+ExlJ2Z9gU2ASPuDNm03unS/4qw1AwaWXUJoRFrfV0CzbeU+TQPD5NDNjT
EcueL9jVfpC8GcHhWnoe6dGDAXWUbn3opCzBfKHSprBuv6e7yWvkeVhbHGZtxipE
vmspgRxhe/BwCxGtIhDsj2GvCz8hCnEm4BHos1rDwxYYypZ7etBaZZ5P3bj8Jiyt
iK0jO51KKejOiJ1fSL2CQPnd1uOXAaawc5cWh4jdX2lfXIR7bu691kHvk8bmDMot
ayLXL1OFbg1fOu9k6u+6cZh9aiw2s48vrs4SDBgzPjKD4odyslzaT9bf3ELqwReX
e3YBvHKtGPsdl06R1NRYiqeqw7GaRYIQ4+QNCGd7E19vXOGS0DFpQU5cl4CV0Fgk
36a1lNH68JJSkE/rVnCujjA56BDZvemrEa8hj6Iygt/XY4E+cMcSbmBf1tisbGRt
RJbFxDmRaBpJ3ALT70YG+vwOlVJ888tekljKIqg84FGZVOVTEF2yvF6fZps5HnQh
ItCk2lnxX1qu30BnY+0qqu2tBqPo3TCGbn5TwcOktvqBJ8/JfwIDBYu44eGKYvqR
dyQZBUejkhRsNQQdQTWFkknhAbAqRhbljZLoQHzvg9/OeWjoeLW2QlAMbDUciU0y
fpJTk2u2R/EGQet/4xbmWViuKsePmUmLL3ORNvLZRFN8fS60eB6vt1HzlqwBbE36
1/nCG5s7lJQvqmD/dWjPhjaZCRX0ceFcsbtoYnWGTkIrWLFdCLrlAPs/oSpiD9yj
MHPv2JxMEKudlNyHZTO0o/mH1Y4OW6U/gAw1rd5SMgcDLojopgUP7T7NcWm2rMHM
z1fSbwXrcAbiYQQf8YEpIyEzzJogYZ3oDdgNJPFvUAdTXDo/S5gxhZCMDGTR0z3I
g1rSKhURT6gAmBgNpfcCgcuogWJzBZ7AReQKePxjAAkGtYAB2vS5e/Jsp9luh6zt
0auHnaAOiHzwABbJBnb31L4fw//GceDvsGpmCPpuyN7yulFBWBzMNm/vxHTPFgkc
b0HjRrzJTStP7IFmiZBjOcTgjXycl5HzPF5V8rhxf5+eR2KlAtT4WA+N6zVI1tIj
ogNc4LnRDrSQm6w7zQRjMjmYP97ui9EKcnI86WHIglbwUOBjRuvxpDSPbywIkEHM
xo9vvNGNKXHvbOiiXADTNsMH09w0lp+L9O00/kzPJo8qWXIXRwts04zQ1noEJTaF
kCRn1eWgXCgR2pFRyOmTIGcaJ9dCBGNC/DfHerZKIivZbDoP08SgQoYlPjxmFbGD
jiiTNXWR2TQruHZ/lSbf0agmG4rk3fJxmDeO/WOOMsPxjBoU676QblMOmXGHbwhX
9DNNGiuhFFeyl/mga/xkrINbqTAXBWKMKM2RRjbBElTdenVfPWCK0lyFNSOkAvXh
6BljLfnwa2ahdXXMmakQjkzX8UkwsrQhvs7yiLAPdXLaord7bVJ8FB6pzNRe01Mg
Y18bGOYwxnMGcHOGerWzlyNfAGoO+o+THP7VTgox9AfIaemQuP+xBgx6/L0ugtqn
YuBXTHvifI41GjpGzHMqjirvItaQJzS2BN28m039H847S9crwETvaTqOr8G9goU3
aWgNrqJjPqWgzopNPO9H80509QcprzTEmZj4qIUqflE1vGCcwWYhMWaZfS9OX18X
BOFaSpZPyZ4pU3CVR8JK0y+dTX1EVV6qjhpnMdIYwza+cjwo5qvcVOgZo8hkZV6A
ChRlz/YjWyYdkQVumdUQ1tw0v9MY/63LzYrIVLw/nhv0CXGX8PuTGvsuhB8D2f1Q
/ZnwnK4Ny3KDngvFuLspt2+HV75J0qdi/j6/QqULnT4c0F9kf0EhoHVoeaYCKpeo
Ia1xgCLTQCTn0wKc10OSXRLTpeeFJtg1TZa9ngitqWZQonrW0OADrj2M0G3kU5hj
HDjLEdfJAAmPAwTIQhs4b2yTB2TzUCOKcHkfVHJcxId9maQeGQUdz7PG1UZNlyPv
oRZzwtCqsjRNNagjejTOdP2hTfHz8u+jLUQx4+/7ShSj2eE7OTVj2qDssuME4p0X
skmvr4SYmYIaxEnfoX0A4/MIijjhwKEEkK0CqQFHiEW/i0wVhTPfhC77NhYVoLJu
xOJ3bvpDL/2i3X8bZwgShmtfBdDpq8+/kLAFNAmiQ8e96aQRHEr0hLubYKln9nFI
ZTuw0yaPzr2xdvATY17jKCA/XUKe79NYZMxPuS/i23PqqsCs7rjnXXjZ1E2aWgcP
Y3cqbuBgVKCqDoOa8D1KgBqncBILjwdsQvypbIaBoLGL7xHjI/xwjVLEjtcdOa5N
J5dvi6282osBKNrk9MJNnUaKzxHWNpkhjeDSY2xIxo7yzX8AbyQ32+fs6URU1+l9
Z1k7L+rrDxxO2rFydFpnyM8Xi3XDpyPApPke+0pb3O9f5udxp38sM30AqJs98mjR
qTxLqeSyY+1nXXjRLjnvrpXU8lZyjklNjPciPM3ZV0EXQWDPaCeuubn30K2Hm0fq
kQTOe1VbApG6FojsBtm6URdw6ROxbagiotsjGDF9agxlZDztg+2tKODoI3wlBkzL
Bz3b6/R2Y34y5BygOrEO3Lt0btMazTVdFh5zDxmD9BFyCOiHZG7b9Fd5GykSBcoS
obpa+4BSvH2AWQG5TxnvWTpWDQEo44YClog5exqXq48WzT7Xnd54I4Obtad/8FZo
RNB0RDid8/ZDdMoxCdq6z1iXTS6YZ0pP5ugBsiYfnCjhVF6vvvr1JlutdKkxKeag
YIU5auIUGTU3I8Lgzux4BccCom1ofYOooV02m58Af8GqKQ6vTySe0k8okoJrs/O0
CZ+RKGoOT7g7chgvmn9ogpmd1+mZdQXOi9TtonuWT9oLsV42cn1fuxd4cUGKD04s
VBbkeTMUgAd5neftHV86mGJaau6gVeM47Q8WbpBblGuidacRYLkNv+lx/amZlbA0
OGo1L0O9uFBq3y/6Bsv4AA6Ra8xaLxVnVZ4p3dL0xh8wMmBunjsSmIOeo2gy8IBn
UNWo93wD/qnDrQJL2DAEZgtCTQ59uYmzpzquQ4IOfHZ4/jt6dDsmhb765zYcdDOR
Fal7MD/wZ9dS8tgH1WS4yV1cUP0hugx1oUFAXLfRqjjXWw2cMb9abwerMRhid+ZV
Rbfilh0M8Yy0eQdNc17TtFIJuigoHiwiuRV0/rhg4OBV75FvZ39iRZtsKcc0dZi8
uuoDtoimMZVNiET8n2dk1dXdB2QL6/4RoB1ycxAWWdCa80ABy3Pd20Af2OCIm+y+
TCwxCdBNZWcl7+L/48jwo+MrAcN59YfrUf+FaLO6+why2tQPEHVu53P0e8YxZjD7
KA2dZnk6ectNwGRCNeRmsva4mtaQopCbrWJ6hqvn7dWM3Et7tiRlqGYkpS1uwXst
b0jKHZB/0PFFq9VC/tz4CNjWj3wlzjBx5XVuHm3KMhY1+qlNuimWkjfN31lAQ8uf
tIWH0cJH/OtIrDT6XgWVTNs3QYz+j143hIUoFAx9WroH43IkBXs2YiDRed/9gFV0
R0sBeJHQKDhGnRtKw11le9wmgKNlB39i+0lxsqUm5KTlszOVyYm7r/mC7YBcrwQZ
MEGfhHeHJudJgExz69Nni02rBu6iXYRy+kyfQlnMUKAy1Y1X2ML1xJaNFtCgA3hK
Ajf7B0OPVNUlBFScknMotIvXQvqQULihomyzPojiDe2YGrlbq6LfJuz326pLE2Gm
GfmAFjvur1pKYwRS9niElkeASwpoOBzjv1tCxHthcSZ8sDDnQPrDgLucwerNAoZC
4UtxBVO0ZX4c7jDCPwLODuMppm3vRDFQMHhj5CjqiCgwLTZG8zCaaxZpVet24tvf
naJMrJfAI3UqGJJThIRkhfFao1lk8iQH22E7WDo+aTf7RgyVPdgnkAO2CDcRTtYb
238Qp/7Uehk9pXpjWWf9/W7RV5nUA2W5qDOk6EdvqlRTpjk7Dmq/w/GZlVCifkNr
VTbZsoQrrKHqxnZyHQMLPQiGbCD0KDb7+Miu3Jn7ME51L2/kcIR9wL/+FR3klP2z
drDYt1RmfQyjN8knhMwknUiCgX+RR+7djgxmYICMW85ukHGtX9eTgTVDc5mlHDaO
0mG3HAvyiNkjuhWzTbmKwV7q0g9KG0yzu7DMoIFIAmfdyPU/TOQeUFu4h2mAjjrD
yW6b82kY/e61Yn0eL8SYw0Tf1VfR93fJrWlGqpw3W2SWRUbfEbvaVdFJ2jG9Y+00
1hKL74q3aN1R30fJstDDggrKHeolUMHeL+/Nh7XXNh2dvWCTYFDtV/S1KfrBNm/b
+MTrHFMo+0pT4jt83cU6zI8+ypwj04s8ype+SRdDgeubVSg9fUANrYwpNM02mLcw
VPIcbZxjp+bb7A6V4ZpdgumL9/hv3WKtPG5Bcko41yuWHWY5+s4xrpLnCXPG1bnW
TFyFnWZnYprrJMqhPlqQDACC/i54z4ey1HYlBouECqR2jDdDLUjsamNGpgpnI99B
O8QhxdmXpl48QniRBDYHAKURlIVtuJT2u7pn0L4ccgd9jFgoIM/0o6GlrJJMxV7N
KUts1fz64HdiOxpXpaSjNGKf9MWlyrbrdfhqzPaXg0Kb2QBxwSffkeEg3UwrB9or
BAsTJfwRZGMJfQoLozp3Y7oc9P5HkWG5nQBW//3E9gOtQChthYsUFdrxYtt/c65A
rNv7el3dgKmaqw06KquQraW7P4lrCq3zVFhp1y6UpNWW+0qbR4YbL1vMLAJIfYKA
drk323oszuX0ukCRB6w7VFEiSwBp/wul18Ym59EiScZrz2Nvd8fbZ1k0gDDaFb1U
V4cyNelhWyh4jWa0aosdvhIfb2iuPcIvKswFZDOZIM6UGaKh9xymNEVauZFfXEVk
b0V0eCF8sfZh3D2PLzFsnSF1FptuAfi54Rq3g9JDiHItnk5llAbS/ltCHBASQtqW
Nnt7clVgheJX+KsaVagmT8gDkqvmiMUu4cGW3Kf/fdyCMdbdBIyppL21JjQD83n4
SOMwg72n61rCird9IkNApm+/LHK5jEX/IPZ4Ib5cWiPvCsCw8fYWc7X8zoYj+AXU
UoqELLGx//7fD1LPe1NvDSUo15wjFg5gc0zfzu8e7138ZnrAWs3RBTPdE3Ptx60W
hJMrUI1gZFPSaMhbTuPydHpzy/I1w14Ow2eyj5Vmh4xCNQSf+vGfRJ82k6o2jwXt
N6DmE1llIckheuKjQdiwE+rhReecVRdjFjvuwuibiapLMX19kpTMyTKa3WUKqPHt
/7ykpkieUpO5kdq9mMzWTLYxhcUlYWyyrYj8ha/NNWavmtgvwAKfvic0DQ8sCdtW
O3iv//Xq/qv3cLH4qo7RvPn0wv2wEoQmrAuzwyE6rM+lgdBAr67qdsI9DjXePPrn
txS6cgbW4UJNiB0JATu+AScDj/KA4IViqPAAcWpyFJYIIPO5MbXUVMbsOrrgQm3l
aP+yZCIkA4MWJ6vHCRtiXXBcaTuib/YUdSdsZ3UqtE1lLbEcwylu18GHFTgp4wZ4
OAv86iADF+XxHD0HlCml2AUx6DHbtv1/xbNGbtileqOx/SSKcPO2oUWH/p2jxCYH
bfWiKqYlyOESVvQXm/sx+WFwalxR1qssX7snq3O3zUjSL5Va4Os0JLQB1SR/o5Lo
dZsUJwLPJO8KWbNQX8VM33LUnwBu7n8K9qoT/JoHxsH9MVGeUyck/2zWKgR+XMHt
oZRC/7RNmFWx0fNDaTSqKd6b90t/HR4MFPQGMLO0pfLO8BrHdbK9mQLVtFhL/tYU
6vbOaODMJ+nNBqcYpMkDnuSOFQsuPituzkQqxotXOBTbpXvXgzK6G99envsh/ZQ7
Vs05DAdxfC6z6nwxiWuAagvJnAfA4Qv445uoakZyFjgL4dt7VoSmYgwx0TFTmDsR
MNOxweSXjaBfBb2IShWtsrIbPAnXk4fRSTHX5901rEInoS4yjg2DS/w7BEaBPNm2
8Gk15lMZVzcp1FjykcBTa253fdXLaUYF89pMgm8SDCqcxFE244VTIqsfOASDbmFa
TFFrX7kJTmTJTrVBmcw1QcxFy1q/WDKzF0FNrkcFcgGVl4Kk5XdrpibtM2X/PAe8
BCZyCIiPdUVyVFXr9w0IIRTJbuU8Vy2e7mBv7YQIe1I2v6v6MYOPcQv4xXCFRt9s
f6dMxEzyf74gOX8RdDhhhPgy4mPiRwPfPktrpWkAwF4ibyRbmLsKN8tTLGJvuoPK
JYG5+wVWXxFz8tDzAMSwro0SufE0Y2fgMBQzNdZ4J+I4az65wZTpnLAA4EBPUrcP
oEuJRrcZBA0W5Vhu4VqNY7XRzO2XlLaz7Zqc99w1gn26H6lH6N+4+4Sk+/WsUzbZ
SXq+BvHmzFrRHe9Z16LkYiHU+2gqlRAObBxEHYoYCHQGGZ4rCUOOBwYfxK0ATKWf
9/6dztqO5tjRBNAIfekA581Zk2xPcBTvmJg3v5VBebFLOzsFf5DTHjofU6AMjdDu
iwTHJx1AoMy9J6inUAQK1VwnR9GXtCIzyoevD2yMTxApWdN7ydhyATQlLoTg8CIb
hw+jzogSNDEeqlNW/7s36P2ix+xZ+uR6iilII4LAuFYJ6TNl/P/5ciqkTZlfDic8
NAqrvQm53u3S8BQh1TctayAnrxDe7Lrn5h1MSqyjHabJZbTpkAZFuIHRYEnUoKTT
oaLNOGN12FkVvsa84aa79mrbmIYmONihEhYcV8gc53CJtWvZpOboCG/tgQnEUpdw
FreNIKwGIvDb8ohChd97/I+M+35gk/us8VylxFjYS1yw08gzWis1CZZeL0upkdMF
R0QjewS+Oss1A4lmHwY3IKMNCK+3ZyolubBDm2gy6VF1JudHeBP4/OhOKZ7CFN8X
3ZsmcDvKsFX8y+JS2Ak2+SLbpKkNod2et7D8aUmmn+n3RXfGSdcTCOmU+VACDopk
l5BAfzMdFcfxNmB1uAEl4Em311YRwo29UuckIYjMNK0dPw0K9g2xgEsizo74Dqkc
CVo1r3IS9Z90aJ0/4xgzCOFdPU8gbtUGjPOCq1vCVcfsIT8r0gzGgQKjT6pGNJQq
FrYiREOu2w3XqVNAFqS1JyGg1mW3cTlHbBX4Icm7VkBL7xgsT7V0LH5wJaWO933f
WiC9i/hOxAf6uldsrMlmgrhGBljFGadAchkmEz5J5TScbwcLisov+YNc4HOOtVXW
AA8/KH5SuQNcNx6Yw7JhIBR1ekPat+YzV0oJJ5ckO0QwdyONuNrC3MB9WYaWXi+e
DujG7U091DU3qwfA7Yepm8rqxnk7mcrHuxE5UHQD4wI+ski8qAdRtuqpavAOb4/u
huWsJ17DkhqVU39m8S/DYzGTnIrHb/oNu+qEwwiD+3AU1PYRg7P1U5VCxIwRvp3n
jGk2P0yshUgjZ5rPSTSM0l76M4Nv+3fX/DlAFHba559hcJZhF0X4b3cFF2i26P8Q
/ZeloEpLkrwu/mTo5WiM/KMK/fyVKMrprXwPoXBYYPmsqsnfkxWMo+/i72G1FJYp
q8uWsi8WryroRNY084otaz2v/V0sWLl412tnq8FTVbRuN1/Rmf5pyLZTL+jAIm5W
TNznvarLgzgMhkA2GN7AuKevmoD1yXTc7k8pwR+SzqPtSZKUATJ+1YbXIRF6TuaK
N76163fYUXNx0mf9EcLR1UctT3wm5ayaFp9oKmN1z8X/g6PPVqw99XAlYjgTb2Ax
B+hr7TZI7osRoiI1VPTPxgBj222MYJXR7c2iMzAbJAYjrLkObsFTqltogYx97fXI
jtGlcma7GP9V46aRpBnlzPaGk8vssAskSCV066+S3lLLj/+NMY6k6swxu4O14OU8
eyUYVgtvXq7eNxsdhWbzhhjgQSXEVaAJlY2BXUC4g+MqXgMm5LOWX73r9TJ7vPs7
rYG4oqCxeNSm1gl1kQR/XJmU5BqRWVP96YaK1Qy/Oa6WBV5CZPRxekL57+GkpltR
TV5s040ujN8s1c4b7H99JHjpdfo7iXr+U/3reFRD43DFTxYO7M2XH+Y82vrQ/3dQ
LBC7xqvs5VvYKd79UL1szMpqc3/5AISrNuRFOFImw9pZe1s2eWEXrg/mn8dnSKNt
5rtZH+D8wPQ0AC/0H4q2FvvfVmnY9aHK5vrTpv+LG5o92FPpHyVMCrD+14tSQIM2
evkvmGOFGKMeFvIiGt8aC2sIXARW4IT3ct+T3BXXGldd/3Rh1XXav64mieJD8vNX
t/UqXK3TrmAlMZt3q8gJx5MVzmAqdgPWlCo6+3QunRnSCvaDkbnVhI8fv3CUi2Sx
6miFKAltG4f/GY3W4N6GLKceZJTiOshrbLBM2bFPu6El8ih1whfq2u5EqSC3Kk2s
j3iaDt0LOY9WLNTIqWxFjNhjqU4oEAQdKmp2OR4CVVDB5ixcYg3oDR+wl5EDN12S
7MGqJy9gUl9H93JKyjt/95Tz9kySdRdOsUu0xXiNLtS9TNzhkjFlMXgV9WXvDlDo
RSYr5ycO6nykPjua/mySIksg7B/D6BtUfBgAd5EELep7aufWi2x99KC145HCwlTE
9S+joIvHO6qeHdUyEH8RIbVqknNUx4ckZkSihcf0JMXkR7QLlOJa0WSyGCI0OmgR
xvDkwgGDNEJKLI49H8R6Z0oNYmC2+p69H9uuQ3tHldcn4BPFiqyy+ID5MLnGjgv0
kNE78VCI6cVXWth7yD18P+OKRFR+tbI+iBoAa2Pt6AQvYtvRYoL2PoHV09Cx1Ufw
ozH8+44SVPLv+Y1dFDBb21zvtFPeA0cQs1nrwKRcbLminStq8R8NKilW0FKWg3ll
TkvSrVEgy6k3qgovmd6C4qYgrCvmAP9QJGtGBSvt/sDSJElJXNuq2Hjzdr+3cYql
CPzU0LnBpYhZEhSXOYd5qQF+DMR/VN7DG11XtKr3q2LLIKksLjHaGoKKBvNCry9J
uAkwb6xNl+q093n8VSZa/MWdZFAiv1/4Y8TKcaHLuBiYBmAK3jTgDPnBX+va10rD
XIAKYCw95Iq38e6xIXhBpJgeKsIdO7m4GQzV5qYE4OlS8Yypp+CbDFnBl+KXOmaN
i9B0zRljOBuD3iV/RxN5US9vZe4SVLyCCMS2LLrCCzzrOsI/Loz3Dsnlguq1IAGs
FYXAX5xqVoxCHJ42vlvF2DO/x+eqRPa0/n/YQd3o8CRiUflbky0I0B+G1U1UzksF
dbKQHWDd19JegeyS3PTZkkRg6oytWQClDRjxqZJCIC6+QvJxmZjCk/xY4ewlob0+
AAJcfS2GAcoNfSuxR5wqkC43Re4dF04fiJ/y7OB+WRy8Vc2J/NRF/CsoPWGA/4oQ
/GoAF8HiG52t5TWv7tVnYCUcMYjVDLWhGICOppcnVuV2KJxtD7BFGzLyuQIeKmYY
2bKXLrmh/ezRgSNlX3hXbC2J4erLGaYFA75OilUFeKF1wvVLztUrL6YxlPqdf5+h
85zSvZobSaORSJIKU/LAUM2wlTZG3RAl4YHx9MinZ7ghMhiUWuUo1qGNO6sRFgGV
e6E7Qj94kl/4AzfmDh7JDOsH7FefSXhUSahg3O9Rztx7JkXxgqrXeRVjmYcUrECd
WMaKhMHDeWcj4C1uwTBIGhVsyTfdHG9LmF0HQNQaf2iIvj+TWukFyEEISGOs+/LZ
SKcbIUI69MJceNJeBLJtc0LGuaKWOgFwHEX1l3ZBYyW33AUcz1A28sHZ+dBTZWoc
wp7PRC2KcbgRPlbiS1xnu9/tunxJDJXxv05gH6iWozY+A6gVE4z7LBe4jDpPnkIH
PYUzgrHViDgO/xT30IDy8E+ndGOa4UYzGoYR5MeJENHA+4POJOkBM5owkoRGzAaS
DGW0Fk5mn46PCYsjfE+AZL2pnsI63ATTxbSx01xbxLgEzgz9zcvaCC7gw6ldV8kH
KwBCu/4zrNgmFUcxq4NdJuPlTRZn6uXMbqe2IHGeIprZoMXP6HWTCBYyWksEMuzT
rWp9Xg2mkExiT6jLPQZv/GrKsgIDgtvO/yrS0CGutO7fGJYcXO1bUCltJvqiRdkj
SWYPtCIK8/Ncr4/NPnSMyynnDSShRHX+9LW+q4NyLq0pXSEr96w1LaIuOu38UZXX
u5ArMPfaaT94M/WqsSw2eeI9BVbTnqm+FaznQ7+N7pGUKz7WyC+R7BkV2gMKPYg7
sV9dXuZmPHgbuSRzCl8hNWtGqGCgH2+MdEn2xFrmti1un6qYOZCzN1pSK9aJEixm
Pc5kwkbhA5Wi88jfEgm4tU95dfumfcd2BU/HoorcXG7CuLLDkKlE1oQWOI6oSjT+
ZoSjit16JWLJ1+hSPliOthL0Ih4AcvidlXZO7Vb0UBMJaYhB78oqm6UTkDmXCJJv
/5hVXVdS4uLPvoHBCdbgwPZOUIPF5o74N4/2rPQY6UrihRWiLAuCfjPy4SIe0a2M
mU9cm5arQWWN40C3pHL+sv4Qb1tWWE2ELv4D/FFCQ5x2sZmga7CgXuC2czbohN9D
hA0WX+p1rXO9AGCMixoSnZ53D+eHjvwHnVnfy+zx/F6VbGgYkuFB6Z274Wk+Xenq
199t4fpjhmlJ6+GWzQBOUY+P29J/Fmr82gwBGZ0h4YoqbexkwndBuRxq++UV8JDb
NOC2M83zNcTF+vb1Qr7VAPhEMCxwFp6pV0piPeafioGsCDWPpTetmFCliim1Kmsj
03dxVJgt/uCYtj94rY1Qf7Kki06h0tTh4SDUp6wOMoJjuC0M+9QY2dxLxO8eUo5a
+Lh6qJB2NLCr5Cn+jYBmoFlkBWVmemPD0cTLfTb0RyhNnIfYb+rsyNri8oDcKNEh
01/Vr4DKCU4rU/7tK5lb4mTpYm6Xr35q+i6JTh5kFVSyqA3oQcDLE+MjNPji9lP0
3D2gQxWYOGh9CJG1JA4pJycXiD8u7P6+5qJCx7KZsEruiCj4vaR62+r8EejmtpgC
qxV+6jAAcGBAXNnOl0gHIe91FpzClahAiIWRU8vvc6NjhcXIgU+XMx1LwKkrW9uV
j9FAAtppAgUqkVm4XFP4LMAiRZ5MrS018uGUppA4FjFmLjIwDiA/krQ9Ae8E9nGv
R9wn5CQa2Z0AFiJE3KuzeCl48smee6alw3qxOMfiKo3snE75yg8N2wucuRPofgLu
/dJmJwxi5JA/PVPFpSBOp2Zp0uB8jl6MzFj8PxRFWU0AyoaT6bB3xlJbZ3N5VZUa
FkdH3X5DIomjm8EhZsSl2IKNfOAdRtiwAS0Evatx84YxrydBx1KX2/QTcWzcJAB6
Z7DYfSGhfB7Zcua9pd4+MNsciJ9ta9U7qxxSXXKADhzQt1Np9rZu/QhKiZTq9zq3
gCbXC6sp3JHOjqmj5gdJbLvJAdJwO37iSdxy0LTrcWwkHCUA+xW2hxDbfUb39gGE
qbFClrvQYW7Df/QHEMrSpshyaEirjfi8mRFJYdLElZg1F2guRtSpiMbE6DYQNv2R
DMOlpekfLIapxst3Fb46tMQGXZxjqEcM3ltZULNhdIEVSGkcT6tNeeddUVM1k46w
RFAqGcY3UXlqPKZf/LUjGUUxsnVvi7ke9STI5oRntSOmu11RZYM3lY2wWF/Fl0xc
VDNt3xM5eN0EKDrRQBaeEDg54E6+Dc+6aRM/h6IGlMSQDrRRhybql8XsOXEC95ID
fAXgQbVKS7NOht+TqLFRDTf8aZacwPnl1bikszlwI2NZeUk/pnXQdOzrLzVvxCSw
SK/tSla60qTsFAjP2JemwqxG57rq/7a+sxN8s08COcr2amny+umIq32/LnVN+RLK
SawgMFyqO8LRsnJp727M3kdTRq0hS7g1pcVWJHgzGm3FmcjvsKv12tzXGylGoCXG
tuFqK5OdfX5jHfVjg6c3tnI31nx+/6HQshVDGZ3pKDv2sKc4IiIFWZycaOL04qAT
l6A3Czlddt9uc601UBBHqTmcNIYPacINOUuqEpop/rEqYFrHg+gzBvbUQqYloP/3
y1HjSdpELbzdXL4iCa0KHCQNamYij36c/LD1AxJ4VFsFNdd4ytpySvJgCeSpVr/N
2pyfIbcPOE7F0KEfJB34sG1oQKLHywqAzKFUyE9rD57cr3aKQk57wplLIZLZZbaG
W1KToQd5SEzBhW9D16yr2nPhxRtC0i2An4iPuzL4ETXBfaQjr4IqRkNE0rxC+MUs
ffHwbf5HlcuU3H9Pe5FSkK6fNgWUTo3Ht0X1td6IRn8PNQfD8wodUELoyMScNo3R
+5AFotlbFBB7vLh3p+XnVpIkWYRn35JC7YS79kjp1XOEDegevZrCr8L4CAxqTZFt
Avp4Gg/yqXHHEUBYoc18YNqT8ozWJ7LK4wZI7Ytl4XuEoqUzQoYEQo695Of8LDf3
RlbnIui/rFPfTKuID0/DglzlZfdhxihf7yfZU8+FXUE0/pPUZFl/i8vHCSDEEB/T
W+5l2VAqpdqgp1aJNLIc4tgNyN2AcTyN/aVEDymRTY1FJoYmCFxvTY35IJM3gJFz
Grpowue2PmRxI4WWz+f2KITGUOX6Obm832fV+uUBtTIGGmzoozQMJp6Z0pJwNR39
ptkDDlzKWqGZcwWq2vg+Vt4GV2EbZsp3jG+x38QEJhhdyZp/wj/LVVYnYo43gu+e
EgxoJLfqkQOYxGDyHTE+9M5FexlN5X0ld2bZXEd4duX3FVo98l+dEGIxfuMhlLM3
cZX39Y4TrI2Ka5OBBi0KK/Kd2AVy7c9EciLYa6aFW9OS1jXVPGa/2Sn7lh/DxGgb
wh/rEjMORaEnE/FOJ6sCSrvw2NF59aq9+phpkzUhTTFkWOi+R6klzxSwDQ2Yw3dP
LRhp0RK3/WzT3I9mjgm3lxNvXGy3KD9Mu+i4XkcxPe29ZwZomYxveB/u9sPpYcFA
wnWuthjhSDqqE6I+6q/IBKribpga/UIQUz1fOyINQCrWV8w9DZSsHcLInQp/Ul/Y
VScPlQ2AIu5uhTwCaxTw10v4ilF3PU3cdk/d7cWzhve/WAlTeMmHhBckOJWWIi9s
ClU35OovUGK9k4N/eQT07fFJrd6KvFqBenCDKVqBEj4Wq/cumEmb+fw4fIpYRbcd
aasAY/7jcbJv1L3D7UJ5RU+AEILb1GXxXO2uEBZY4Ksqd6ty+lpGIThzMuPiAroQ
NwRm0GZ7tCFEZU0ul6I7rc8R/LBPNqVn6uPU78fhBOsuAPmxPaIVbJTHpZhMPoUK
p2gfHaA/I6Z+TI3ZJzhW2imRbfvjdUAxDdOIRXGmJC2709BuR7evdbLQO8l5q6+d
oFhdVxQ69NlK20ABgfmv2M5PD/x9+OrEWd08fcFV/FG/YkBYoKZ/nz1VghBsJXnd
zC74QmFN47RmuLWL7jgalY31UxaOUCjpCOHOFIz6+cny4a5LBvOolDVafQeWJCho
+1BEnY0vzdbNNWesEgKNP4ReeFU6rRvhheNneSQ/cvkuaBYzeNJQS0epx6JwDRSY
0e3ObMXDjhbnSTik0COX/4M7ko878Fk7yVn8qMdWZ9MbeqDXdKVzQT36PzE0FXL0
HRmkogBZRzJPO0O9rbDgGCDhe4i5fxkUPwbp7IAuuzH0o5rYHrUnAn+Gt9ZMiUDs
tQSne8AO9pjykYc0XBMrW3pcYmWEIs8Z4zdCVsA7/gxPY/s+Sk17nk7pCVxSCMHw
9wDJkv+vysHJkybTyzSBOgi2/Ml5+N8Qe6/XOByrfyhPMkhNkDbjFophcQY2q6TV
/KxmU+5y+8+CI9DTEqcSxLvuf4YxlJRKGNDwYQ8BiN+lPS/dJsLn5AsuMjEis/Bs
ZUsRLIb2eCeBWiuhvffcUj0UnXeUqWguZ0iW33HanxttiBIpX+/JuL493jcSEON8
ZOVbG5hw/skezvDyRLZsIjKRxUeopEsZhrbHJgDb4yCumWqwDFNfxwR/85yJNHIA
rQ8HNlXVV7LopgNdSvI9Wag3EX5HD0MB+ZxCoWMvl/ftKiWxuuf9DTVr9jVtpS0m
S5B5gEnqdDhXyskb9+7zUvqOFtWrrFzoUxMIEenMPRFWb9l8vakjxSdpTUN6OfTb
/yMs+HyqQY9VhlcW5zQZZJVe8nFwnKDQLMKaHVzSwm6qoguaiCQKBjLnJ0smN/Kt
7dHxrgfAtKBKLfDdOYjKe5ZMAa28dy22OE9HcixhuznyZlngQ40QF2hsgEzoOWwN
Bg5NXTth+BqkhCPYEjDEIDqQhDI4Zr3hPEQFsoKpSx0Uq5dbp3eNJeXZOWVjhxWQ
kcJj0PfqHiv2V190rWPteDiWVg+LDJdLpKa3SWI11GFRwV4baPvXlvEfWAiRB17f
rp7Wfb4GDRqa+pLDM+lanfVyd5f5Iiduo5Vb01yzFeAMBa0dg0c9cVT8cTpX/Idf
so+DD0Ey3PIClhbWnEmrw8d1UGLerSr99E2bWPswEI9VlmK41jMnsZYHd5cJe/Cf
ossHe7xNznkV3VyxTy08ZgM3pX15xYDPmSX8mR+FSteo4FTeJc8R3UDHohP54jpq
6UMxPKNHWFhrbDECtP0QjbLd5QU667vl8CnJh2okOP9kyynYLDYfj1X5LSgKyJED
eGTz8ADrw8ADQn7fzqoB6S6WFgJaQSssqPEyobbnf76rIbFJw/APLts9/2gd2yIn
AJtxdifaV6f4+dG0S+PO4qixnOBtbDse4PmiChQMGDh2o+9BKxhguAsP+ak1U8cd
lrL8RcjFTMPyth6m9dEufCDVEOYUtcHjc8d4TTXoburUOYcT9myplHWpBe3CKlzC
SgH6f7KuLw3OSxFkrxn9bhEPwH+1IU7cALIPqLMMPrC3ZwXJ7jIkS/R5f6k7hfYn
TRDFZtxgNeJAjUwQgdqGuera0Qs6F3P0HT4OlzcWInQlcRR/ln5YfSI7t84S9AOQ
/P1rcxZZox9GvkZf41ow4jp8Q/9hVfX+PyIQHb2+k6IGphgqkbfnpl4WimiC2gAB
Pozel6xglVoBES6DnY9h59k1Wp3RjdXgI0/pAxdQNB0tMPdnRUAl2OfN8gWIeQX8
I4sjikvGj7g4VHTS5sHnRGgx6psOYSIN6Y1EJK29vpephvtyh7sQXvKT9VW9GNRd
+NLVULoDC1wM3pgQ6U8Y6TawRZVK6vrf0fHd4ngdlJeMv1Ou5r2UFGIIzKIOeqXN
pq+gK5rfuk+EYTnj1UH3LpConr3czzy3XnU+NR6hpvLbTXAISxfp9NMlcus6gToq
Szryvu7YODa4EB+HaZnI5BNps7AgQjmVcY/of7KYFiar4Z5rID7fv/lUFFY4MMXt
qsugQdQU62e472O9RN43ORwa+fWpOVFMmvUiC/PS+R1rrDNHc8SeabLRHmm0BXBF
CW5cXI6PAW0HtPIryVoeHxBEhHJ56rrPO80TW59Roiss0qMb7+ZV591DVo8eTEAS
Rolv6K9+S6xXPeOmu8y296X5n+PhCdu4oXNBeC8WYknn6c41mZYz2SCnePpwnl2u
4PtfkkWg0RrHk4GZONw0CG2C6UAfrd8BFbSH4Lk0v3yIR140rDjvvEhxCPhclHts
O6rvxrKORGgxbFfT26uHsJg4ONRN2QH9evYC4TndDJ5wBAJIEQsFsIusoJtXw0UJ
Iu2ZT4zgs0vR7fwTdT+GYlOBKL8/xTfu6wBO+Y/a6aFGGdS/Cwd4zqhOkorwjUXf
4AhRsVWXi/XZI5nPGd7XdMxjDimbWWVw02R1A4DIkqyGs1Rx07fOLaEwjPnDEPn5
zC19cBtc4YfTvgP49yX00fXxIi1eWJbEMpqXoME3Dv6dFbmEwYFXSg4O56syqan3
KLDUE2MQKqrkyi2yA4iANiJ58hb7MD4Jf5gez3cVX4/aaF2oTKSVCxg9Vxg5/m+T
vMwOBeEON2Igm3G0t1nPUzxZamAHrT71CPnjYflshKvwWpVaQbfeUwhooSVc3hPu
yIk4SrWn33YfmeBhknIG2PXS4NN6P0FQ9klp57oX90UCtJUXYzctwalWAyjHegnY
cD/fzlEP6mX3GOqc+6fEEKi6Se3ftejItg8PKBm6vl0AFgTZG6ysidyF3aZWc5/a
+sn0SieNkwXxGTL1W3JajBzSl9ZEBawuV1UjXMe461+ldZMjk+tCcB3PxtaB04Tb
9lBToFj2CltVBa2lBids955sQCwpbSdcMagQUcHimQF+EIJnvCkFrWWTzTaUp2lA
oeqajGTpu+Vh13qF9OYNizcilINp6prS9MRj0OliYuRHx0f4lfjHdVmeh5jVRM8s
lvFZj5nAvpQUu+7OoHpNjUDEngooL2Cigv3cgr1js982jrdVHgdAMFedIm2bH0EN
fK35CuxNot4lYPDwLopDxUWU9naC7BCI8Smgp4s7P6XKZrUg1K6Yid0G9p5ICuhg
cJwl+xev6oLivq5DZ9VdLJcnsV2PWYzswktlox8YB65/F+WCyHL2nQRjfMNUqhNB
kQf+cQksdBzwJrIUPcd+spt4/59v0lNHC8bJQvTVbGeijkNWv7YjwjSb6uo+RndU
iPIeUFM/4ISdKlDTvuYHOgqczsF78HURvJ2aqx+h1shwrJ2/W7qqiPBCyoUTPfSt
Z0cxS+gbH7NNeUe4r7AQl/bBT/xlxvLZblVIsbBLlolthNOX+qWU31uzxpHDAVfo
RVvsJNnwsi35n6hvfYRnu9dP6rKhJwRdAK3iuox+ACySBW3xBn3Wk2yys07wK2WB
JEwzPO9ZF0H6aEkT9PzhO+Ih7dQJyM+nB/e0LglkQJ2GJfo+wbON9hzEkJY457s6
9FvJee556V0Rh1Mqh27i1JxsZ8pE9FbbFRwgsOKGvvA98hoVg4ukByta8Ua7TKTf
T2HPBDBmMDXe8YqVZAYu8Jyqw3yWQ2gH/UGfPqMO49Gee8WC8+g589s4hETLAfBL
4yzZdXPdkySpCDGhPYnSilaDKyQFhpiM2o0Vvu4pcMbJeHGkoxEj16kltuRva0bY
SFXLB/C0vBssaSsGoPpBBA7vW4GoA7+pKB0G0R8j2Rs1tbVjLnTz7uTRog0c/ZcO
e9e04Bomcv9U9MdcEMMKLXrGwvYAtBEwQaipFh52cmaLu+nvLNogACrThmR3wp45
I4C8sKSkhZSkzDlFJxhMQsJ0uwPqpjBN3whaGsXX8AFAYjBVveFBzNvI7g4xJFra
Dqxw67SurSffh1XZVwYsZXb7BT/OK1eplFDYNcJqgO4/B3F+DrFvFHCmOHrZU6rq
YbcJNM/crPm279LfMu5UNcDZPY+y1G+fKr3ddogExIOc5Svq7PTdWV6pKlRBKCTy
7VHdpOr6oOZMSUpI2fW0+xPR5pN31c0vK+ZA99DPjP5W2r4E5dmiTV1jyw3Ia42u
Cue8jLujQSlVB5jyfdQNLNI+bndAk3IFW63fEUQOYBdeAKIp6bCEpQ520aE2uFVm
MhgOY4pBE43UJJApmGjphKndhCHR1F2eicagO3h/0X+67zqxEkX7PIAspotF9uYI
gHERITVWYVYTQNiC0BE4DFvvb/3MBYeM7nItvVNQ9gKDwndwE6a/Oz44mVF1Nbof
9Nn5Ztqtl2Y9cJ38QwvGi9oPEGOZYyJedKv4e0qyI8//D1QsdyD1osqkGWshMofY
8f6XGKNtbOGWzZ1S3Ig+6ETMUBxs1ERPXcalzMMt/3ohHnYwu97rqErsFnYLgYzL
Qhhp/UWycDP4WYUfNuDvgCSyETbRVv0JXzO1AT8aMj28oXfcpqHvZxTt8nlwV0se
n3TTzjXidPjUVoBO2qu2TUrUYVcqVZpssfowdPle1QeRcjVLeE2N2DMsP76iYNxt
iOemYGShgOErWU247P7R5Y6J6/xehQsV6uA0+fGmOEiFuznMeAeSDSbolE/TenkQ
EK/UD5ehoxo2DmKn3gZikzMnYzBN1Ka1dh+dlLnKLG8XWTL4CHzYeU9dvyqpZbLF
F7WtH2H2SVXwUI3CS3cF2WyqhLGGFq/1fdNHbffdUp2Nwmsc2i06W5zqLrQiM4Vx
9M3YzQgAlF6H7mkghszWvU5XyJQfDIag4tZlpoIyQb8NbxjnNXeurWWsDJ9xGwoW
L9azXUy4dKx5e7UnSSk5MIhLKVqArMOTxzHxM88RTCCqQd0d+rxlntSC6Hv7t67F
o91VovdV5UNOCXrIQFavS5pRDfmDxyG4bi3V1/GhmVdZg/MBu+bYjpylg/3e+ZI1
ia9U27/+IIK3SvZvGdTrhMgkrq9FFKabYszb/AdUxBsbOftqB/kxe+kslfwEJjpT
RVIaBGeNh9W6voB09VOhHfMAYTGzIcYJZxXWc+u4FeyoBRlAWg1djoEifdNXnR75
IYuzr4UpDfv24zmZ5LKCrx600Cd7K8A1+BoMuKCutrBnTChjIZZ2f9wSIpNPBPzx
lm3x1ct4DgMBbmoG0ht2wdaS160UKOVIyZqSlbFzU5YFbU6Rm35IiVL44isG4DSr
EeJHKZwb7a6U0ak+NlTRYr59pFY7RkagBIIDcxlSPIpu1rv9y3R6aidGBgUadQlm
lELw611hEdhfzoe7dm0oeMFWvEGUT+KIMgtA5SMAmVPshv2DUFVHhsU/7iivHPLE
pUIhyVwsKxREfet12TVzswHAsgvvqEoLOHreSWaPQgaUiI+MraVz3x50aA8p31Os
GKoM10qfhTHz8kXn3p/6pCbxFBiSVbVtwEXetQtHCL1vQVX9shxgPUIPvtfRFuMG
jnxiLX7t9ISmdQfdKdYUYAT+XNDZo0Ms8lNBSthI0f7In7WGDaPDhGnCca/kafPr
8J0ZSBxpTwT4DeiRNMK7vO8RWSBXLLWSMkJuQAtSMLxInVbB99Vn7cTkTCkIjU0H
YitVXp+QmDXGefQXbCYnDtEJMAVGUkrUmwIW9RVu0rNaWTOD1JAjnmDIiUS3OM9d
O4MTxofNScaZTgkw9Dm/VlOmtAqeIeuM8BasLpXPuznEKTe7Mm1R05C+ws5ZqUs9
zgYjQKPsRjrzFVrhlSy0js6JwMvmXXUg6Dq5+gGlKvzlPtoY7p7AOhXCPVa9Yrnc
EiGBAHVkCg/GDbeECRtV0P8wl9cjovPDXQ3JSaRW5QXGCTp9yoGb2e+3eyboH0sl
HdyE8uiNH4VbxbulLzVRP+BbG2qlydUivp7Um7G1LkrEdT/cPcK4KMPlsxiBogr/
fxgASl7gMXmmZUSfea9H97Rme1TVc1/sE32ADXTRxfm2wIk8zEc23ji9nWLmvoO+
CSuadq9rC0m+44cJC6FJBsyZpAEQIYI2eKuqdS9Od20Ym1PotW56Wi2/768UDfYu
U3DpUv/PcoHSEKFawAD2v0yyNoSPINOFPwJt9p4tDYpN0uvae21L1zDZSlJznZjd
seoBcS37xLqIDiID5kifCATLr2khjtCrY3e0NFCt9Z1FnuNezgh9ih7LzbN2eO7U
EnufYFLknOIyBsAklKcghzX28rD8VHi7KxDGuzb/WJlOh+oAlTZXhIuXAmnbJhcc
oP2ZVvnu5N8eMY/fyX5DHLWS2T++ucCIgwKAAFpiAMx9Rtb0jtamDq/GpA0ESSyX
SZJK8PkhbT7RWp8iC+kISqlvxPegYPmRiHDIEgN4AD+F+FJ9qPnY54Rm3yQ0w64/
6dywiywKNu4yTjCGhcR8oNypqoGvjxknyl4QhoxbRVsMIAnNKla3lPhsNxhpVjoB
TPEDg1Vjrndnn8/PJszGIow1INu9mwHtz+GqSQyarYHTFnagMVO7JdJjP1Caww0F
OmcqNC03Vy1+B0vXFtetGQxkjZC7JEAbqMKtSFeW3PcnSV2ZSgAZIrKkuh1QYPuY
x64zIeKX7scmQpWna2E8dPT6c/SkqsNc3CNgvbbgYDbX+lcmQJCRHII/UrLLWw4/
VmH90VXC5Bx+h335a4WvIgLVybP0yy4P21b/lCi//aHgsrl+MAPDZUYiwMQi5t42
R9RxS/TIeCWcoLizyx2mTZZQ1ge/Fc2nFjB0qa6F8ZIBQRL4xXzJwffiqnfKcsB/
BILr+0AaLf8um6zeK49rMID2ecMTHRXlXN+cDf9t18H2rBoqnDxVtBNYNNONXoPK
G2NFi+sdtKyQLhXosy1jaMsGFZtA7/AKDJdkj+l5R4Umj8lt/R9lx7HsJQl+VMV5
zVjI/XSnakk16mVbyejveEZKGYA+c7m1ks3nCfTQF0lrA0uRN7IuJ1dFDed4lTVC
mCVuvAXmAlLCcb109Xl7Q4aB/3o9LaTL9zjpImGCDEPz4AgEw/mbyaL/MivjoTyH
UqqBSPZmAgYhrmgbh8E24JGPhVwE+s85MXh4S0+a2/dPbmpNbZ9DP5+QYu8RKUtO
6a33gdlFW/q0URTi2qzEP1PAvdUl5SWLLmZ+bS7lkIclzcCCIKRBy0YLVJDe2uNu
7LJbN7lAJ7ySkhmQI30NbxlIthRNqWQv8nCmbL6eGSiR2Pamto5Q4/lXtY21rWwP
ycaH5M0kE+dh1Mlf8f7CbYoS3WVl+Ci0ey5CaA12N2nKckjumqTsb9WHL+v3K9YQ
AMU9bZI7oYrDHZPIkpV0YuL47o0ntq42D3scHysU0UKgnSHgtpu+SzAdLBzMvCL5
Zkxp6LRKRuuChfbUQun/qzMisYDH7M+EPjgliGMvDGs7N06thPfPZ6/Vm8uD3l+H
o1QIjCuqudMU3Db+bczF0EU7dfN1k2xEKJp/Ts58dYEAOLCa4lf4xyb2LlGc+7zq
X63/Ht6fhNSGIaIkBJ4Ic5FOr9pEWz8LcZzVRbx9NQ9ExbK55j4rMpAPtNzRkZi1
Vvs+A0QW+rbKIvBObdFVTxOYPr7AkAYZKpp50eWe/hNMHE3BijuTxdWTQk1/36P4
kU1e4ofV79M/ucXvRC0SQG2+UgrDm/IkivTLT9rlFixrv+KDrx+3D1NI9K4yEHRa
gb0HGVGb0ZHV6ow5xI+ER1ZlJ5CffLPpSzuWNV4MX1We6Flzh6GapKB3xHViYHoq
Fh+TZ0QubsWzlW+gHv8MRwMJlW2ikUSfckVNleLBeFPXJ3zHraXBJK/y54O46sN6
VYNM44m3e+9TLS5pgBi0QyMnjLF8ziRSsGsmCIXQ3tox1OhqPcpyBxneE2LhXpLd
ZcwlihKA2WdkVBYkbHx8tKZKc4/rYnV9BtlMN1soiFQTnnYZoumhxHOdzOOtoZG6
9dFzi3mHeDhOynz2vEEp3EVDxOUZdLoGeAymC/Z7ViFFOVf7svszBpG39qkInetD
tFOQJrVp2II49C64T7dcxaFHMi2L6/Bl1kgaeqOL7AyZuDoIZwQH1jXjES0YJ7of
4agyK01+cvI/N2cIv6LUC80szNvJBeBe49Cx+DHTCPpvV6EHPpKC6v8tLhDrhCXI
4ISvIegK+GxEp8arY36iZVJyeNvweOS6UjqHI3bm0tqNcbhAk2qg8IkV++ovi9+6
0oOubCOhfG7zjPQk1Zl+PIepWlQl5DL+krJyd6vdwgy++oPkRDSwyWyT3f67h8FR
AtWYH/VcfvIlFsZVtINxfcytW8UQGFPmicWvBc+q0z/fJZi14sAGLGDREz5A/nkQ
uyYSYJzplhcdbgYd4OxYcuysRJ/Yx7eeTPTO7wKYJ89ciS14d+tYtNT4bnYEXD9S
QCqhCmb6IQr3qEaLfWz3gA3/5ymq2JRj4/tCKDiJ8nvy+rWfviWIwocf6jQCoPSb
O1poSBVP/n3MsG1U/Y8UjHKee37aVWr2nYKOj/pj3sTDgCizsuEOOi/U0cdZP+hz
sSDw0d8luqzToxVdjuDLpDvLQUP6hm6deIKQZt70tv9Sb52w4CvmSVmrCByq2BeD
GfvhhxmHt8bShyXzneI6RLVKpXjIwvpfls+u62Y9rrvFZm8CED8KBOEdLt/RA9pw
tT3AG/qk6qxMx+YMxTVvousdchMFKleVeRCU9ViquoT9+7/g4gP6IqH4fdZpryry
CJqNX4eJnqNeKySGSzyukd4RlE4gnlb71Litm7JSIlHXG5eiaacVH3gvBUWFR6pY
9box14D4yhFc6R9ar7gA1FoQ3uM8HNEjJUNyd2GdebblpG2K3wLnkGVvt6JY32xt
+c6bc1gOj5Yxew0GGqeqSVhzGkOU3R0k0VGuyzd6puhpXVm8u8Qu7wf7os2tClA2
Bcwj+Ov4VWxL7n3UcDwi0dHkFqT+GIQ6bPOkzHm+IX4N8XggYpFko8UgDJ8rFuBX
JYFYuJQSDZ7JrwI+UsjMOSGN64ihLISqnbTTPsE1Cz/ZYLUiS17RQ5AcKwTVnei4
2ZAr3EktSZAQK6tquvDfIiySDFaGkMAuo0ePrh3X4wbFupFMaMryYru5q1UtHJUW
sLTTY15W8KxUxNUINWZmZtqsxxzLuOG9CHvJr55L1dRTG9tlK3FP06NeNFc+rt2C
dz1uqOe1URwXIACSFdowOgUSjV5CkQYDkZ3e1J/FYIU7yoghS9W4rwzcoDEz/Vmo
AY9+Kv+Jnv3JON1KXtBy5cF5a8RxSCrWHnptMSGDN6TeqP2MwSB07ljCGjnHWoVQ
uFuXM8wJooO//wS74AjcwQYDuiYkPHpmcb1SDN06/1ruGeA4YwwAA/xUvjboV21w
L62PPL4PNPVezN9IbO8ml4zm1n1V4RLrZLf6/XblM8BHTftp3WHx76j2aotkicON
UWsJDK45pL4teAzTM+cvgNb0XnLjq+6njMuFOj6wGVAv8cGmVJnS57jjxxYYHHFx
zV9uk0tao6u6S3xNu+SGmpXEbOReYPJ6e+2Y0raz+ss6bqKvCK481wJNhGXfZkzr
L6yJLGmmbnICLeoNXg0kpeJbawEA9DJeE6zuzquzk8feRoGYcFFGuwpw+S99QoCE
pMFlom11jGERNKF/+HzdvS7bZ2KgrQoFEbRik1hRpwywwiv5/CD57Rh9Hm4SH4iv
fQ5dHfiU1cFz/dbxaicRJwErmsguNAiF2misFBV5y5TWrFkO9dwSlxLo5DINBqJE
OENpuOsrh6Yi1dZeSCVzhpHX9get8Kesr1gqDuEWlZq5lNV8QQobpHk27CBMmRB8
609gHelM2ie6kquTZHzzN3fuAk0UzqamwNen2uX69BslbOdD0kAf9S/+hLQC/dRk
itBHrMjv2QSijnpboYxcvXTWSL1/N539zR/uuYT7Mw09+yjHzx+piTGC1NiyBCRS
4eLGUgxUVtL+QmvhTKFwf1GCKirfr39qA/6WIBjTq05w8347GuESqqj2fwDMSBMz
Ejkw7dU4ExQJEKmbz3lpc0cR4b+uamUmFbZjlZnrlzAecGS21neK9AAjTg+A6CVf
89Fqmt52W/rIdOkZBUOSSbTz3uBP79eksYjU7qmi04Q6gnZxAf8oxnbMdHIaMtI4
NL1UidZmDxqpQhzDVRTQDi6PcsjzEBkbvVTURmEwleWgOwtG/ZqOQyN7DWtzK8E5
O3h4TUpKyIw66Q/sbvEmXBKt0cARdud4K3PQWCzqjy7liuSyWaP9uHJ8JuaGyt9y
jhN31uT5iRZjGKrPpT1ZlVBfDdO4pVQhtFu13nqwZ1yBnqPyjwCmQFXscyYJYD52
RatOh9XAFGG1ZDIEpNCUfdkD5KXOUmlxooZOos28xFg1NM7+GzIvGkEku5XGbM/V
YSAVNgbynNZLHS04Hl0WWMt4fPaIMN4bHqMAZai3czgn3UzGeM4I+yC0kilSrFEn
6bLvhROU7OfLPovS+j7kOfr+djHmd/c9XmWVScimXaTrGQdPp1qBSd2JOKaehG4v
aG4iHNbMJGlRwsus0MK12YqQKgbBUiOtZuqhSn+MUlnZd881yzgNIx77OiL6hCB2
C4gBosJT0Wxk7YLHmlzQ+Ar1U59Krlt4s879wAKd5txIZ0O1ThoxJPaJwOm59b0Z
7yzDPwIPW0vXwDqpgRVcLWKm1U7V8X2hORW+c8KnyUWGu8oJ9qagCuP/LxdibFKE
evGwU9xGsVeae8gfUMdJ2Wf1j6pvF/QLQxqSEgl2Ge6Vau4GmXrZKkbkMl+Ny1Ls
D/vZPN+i3GxMXDKJ4KzSWM/8AXfUORmHG/qZQLGxYIY+rWhlkixqDwP68b2saZV9
AfxHRl2om6KED7aabSQ8rtQJqwHs0qPHOwDFFDpUVSx3zhI2MnNzsQqAAXT0fGJJ
NaIMMo2r1c4eFPg1RI67MpiB3DH6XIWBmkrAwEHzr5BnlrHLOiYGw/fVm8DfDI0N
lE/SC8mDeFoRFV75YYk0HwnSpU1AHwqKhpp8JaatMDcu1qXL4Eh1f5E15ZtuaLsW
rC402SWUNrq+5HswtM31JEqBp+EyGhXCFknn3XfgJpH4nMTLG7Vy5TWgZA25KHM5
ibs9kkQT0wQ9jQjqOIBxQtrjcCig6UzS/1A8NyPSSUS02N2JLKLFISa6Y0s5UPqe
UjRDFHcIXyzarigL2XLqaWlw8+cV1MNwtU8ju2X6zjM4dp6AZ6pbREnMSi/VkfZo
r4MtE1DNg0EnK/RpqIxc4UTDmYQeSjJO7A+HYenii7OrU/bb8D4/bgWuRw+hWbRa
rxCvcCGVnVvWHKM5wpmzsV+eWkomxS3j6G2Q46xaonL/SxFiS1IWg+AO+dB4jZrD
FhWim7RA/FtJMwjheoKzVAw2Abfha4BlN2V2I1zM+/em3aej0kxoqyh9ub1dnOhX
Qgg1Y9zDqQpI6GplnCEzoLIY+ltDECN0F4NLm1ifOON7YU15O90jN2VVjEPjWwG8
Hbt20eeDmPM/6Wk+pZ4Uf3acrLlTQnBvtIdAhc48Uo4dCc6vSUZedBbJ6/mSYWkN
R00g11lHN5LYL2EsBzhM6Y9QgtFp0YE5Q162TWJuKhUsbGhda+BNlCrITExc/BO8
RmUKxFgks2iOkSno9gjMJr2+j0T4+JuwDQkkMKq1fw8iBwy6ALnB2lbRZWY33hBQ
F7q6CfzpIZ2qCZtYz1vNGCC8ffAI1wU61yr/7auTV6fb4jCF887TE6ig6s+JWkXt
+zHA+vq1wbHMwgMQvGeb9TWPHdiX+d/VfVu+8SE2hDuODE0rcEUYoLyccg+9+XP9
hB9GE/gdS+H30Bdaz60Wy3BwuDIv5PQGYAThYhjM+iSNB/EqG05qOQFUUx302G5F
xq8GbXYTInauHt/jq4WGaclxvCjJPVt6al/gniI8rQuR1Ggav46EMofjrlZ7A/zM
4WpMRXo511fBGntXT2ZxMrw9jLYGnCiizOpO1sB1LhMWg38qgXILOLREiM6KWjwJ
4n1S8P0S+BLGAmPUhIYM+5CmmHPreosFLvWO07cptkwpfXa58CM2pYD5/QyBTKX4
G5OIhOrsHDsZD478vF8Ylo4xBcsFhyayuTeqmid3OYPfjOjdURVb9W72SmPYtOCI
rMweUCE2o6CJMNqm/Fo84sjjqreFHFYS2d3MsRM4+veX0i7r9DatwvUEoXc9gXjt
qumGLDZ/0I4PBVnsTVTyaD55JCSTHUaP2cLZloRmIHdmN5DEQrUjVpII5OEQWUde
Ri8AJZ1ZogLj4LoDh+yCo2A1EGpEmxHqamD5BP8Bg3wn/4Eq9OYCU8qx4yf/Fv63
23JL5c0Im/QQhGY87QYgwX+Dp6RuAGajbQyr4mgbHSgBw/DZHwEKmOqbdBM3xsg8
oGaW4BEVB4CL0TRIqTwe3Ne8rePmQHoDPka7/15DwxNbqH3EO//m1Ab2X+r1Aiku
HTlVnQjXL3Tn1ykJDjaFHtvoTpqjr7nRkr2j7ynskQ2OxXdTRfpCV1r5X49h9dZW
/+7yMvOYrcEmI4n5Fd4kAYC1G6JhU0NqM2+XlsrQE6h04kVwVjMCVEpwslqQ7GXB
uBW8vMO9fUEOuq/Ej25fvlhS37uEF+53iYm1Hr6F0FqBEEPSOZQ7uPXYcxnSiO1+
00aEs81ArfkzXlUU4dt7CPLLLVW7eyVxOWJDUujSrOidJzbTQLNJswH2BKiDY8aK
XUfEqK+gW65gUm+kW0e/yuzQBGDzluqGLi9CdFVEA0HSRjAB7d+ldFigE8JmDzdc
LI6eSWIttP/87F3tZvSS9oOmW9A6r5SlZDR4UgkKc1hmBdX4fNNsXnbf1M1ofTrh
yf0QAQkgg60piVS0fYLsWSNLaaR4ylQ1DRfBXKKPIe5DTtjc0PhsfDZupfWqagyl
tiO6r7o5eGEA5O+N8AShWhGjifv+Swfio5QVp6qRtE+/RIrFm+JaP1Jvr7zVGwbs
AkMLf78W+4uIiTBlTUpzWY3SrRXBpiuqEiWhpyj5nu1f9Px20hAp1kLloRc+hvIR
nZtVOCTLrmbf6TP0NsBQoelLNDUiJUB9AfkT8b2BldCjmq22PrCZCS09da49K9Nd
G29LMUgS2DUh2XlncDV6/35ro9MEi9qNINC0zLk5RqjN/txNFG2g9PD8gRQfGbFM
zgDaiyp9SrSlo1FscYGiCWts+1TEk/K+AgN4KTaXXahe9gHn1VKkbymg7DGMWk+a
pmBkQLMnhNVfkK9NaIlwp1LQ7BTI7S2Z9YKSeCA9kNHo5+GxglXPH5CLw+UYFS3c
9chP1YJiAy8VlhU1vqtVnDbxURv5crwZDNyCXjVCx6U3gdlIUmXk2s/dKZk63h1J
zCElFnhqPBDShtysigz3hAi/REaWpBypJFD7eDt0Yqalt0rdA4MRKqbfP3DumjAX
JBSmG3L1TkTcWYC3D2R9NiM2Juzi0QgvCRiriRgfAcrLbRBuSo8sAX435WFaopUJ
dgiSrrIBupSAzDUyT4J+W3znHV6hEt1hxIob7Qr0OKRHKB4SCCYISjOs+24JTcNm
NPRhYqZ+16ldhl+gVKm4fdZ1b6utFtlG9ZghWgRX8q3GiwiGXe9ptcebgxX11dw3
kS6n8NQFJWrnws/nbN8IiEbE6gpAy8KLDasU83+AaQhnY5lmpJj3U4ll9lcLnGCM
tsvEIeEeSa+8oJwmTYK9YDn85CDMIrs8UP5P4uFBFYCnLbb8mjXdOBf/3H0CFGeu
yiVL5X+StefwIpiCjF+lIiChFs+VYfqCmXi1taSAO8Pr66fDCNj47EPRabTKc3jl
0+rU4RpdZKdlZcD7tCNbA8xC9euXPbOArI2pFPN3iyTzdXIB/7HmrYR6YfwwrNRA
R1pNfcrLzO/dGBcDjLNMzMgQoGbXfXIPp05N/ySb0c4GN4gEihHEsUbK3oF4i9gN
JqyvlVLE9DHGi5QERZ1FTVvXTMrmOGgwp6Ji0dj17D2h2xLfoNvgLS3Uq6YmJP22
D6Ed3gjsSYOvVPGG5chO2ht6ZJgBZckFK6y79+6piRslSYMmFUCDZsG26kF8Cqe8
YgMFGHVrEL5aksPIEH3i/csXwZpt3JDvy2f2/aoJQ50o5kcuTvr5EhZ9UGI4D/RZ
rbnEacKBYCkAU4JMml022yRrJrCSQDzN2AY89RzWG2MknycTXqCvvOsa1pWzYZl8
o2597CMMakhrISGDIn8xyx/6ltIzrzk5si5nd53U45k0Yr1N3E+wSIpsRrFBjl2m
CiRV8rfbpo3EczZ4oLhqLAZahAPgAyEdnAuHnmzMD/cDMzpdY1II9kh3sGCPQh35
c3P4MTU6ADte86v1CoYB0JiSySmzEXhDsu+nnOK5iUuMST3pFrsAFpIzeyl7ioWQ
iEdNdckGDmm75ai5NFAjVNl6K+uxW7kIMwZxKMNdhYjZaVPfijLV3x3VCtIyxv9h
wIwxNTSIuEk9deh1uk92hanb1ZvHbdbA/0e/yAHfIG5HgEvSTX+DZqBA53KnawmH
/KM+qx71Nwwz3pgE/duwhnkIBl9zrVK0uzGPu3Lzc1w6TIlRwZC6+gbNQKidHpeN
dT86dSyQHdApEEDS1i6Syb8fxRWKoVZELESjrmbWoRpHYh4suvacoaJuoVR6QEls
Zey9RY5Wp01Lg4iXUMwa3hZd6zPhjvwOZWDqbINd9DcNIabTjxW+BA+cqoUxRtA8
GMAZ6giu9R8QCeYEUgV9Bhe+Mr7V6XqTgDWQNtZcxewlgsA8vqiKEBVfc3gj/1R/
e38czmx/+9kLiRuvwfjrliiBAXQRZMCfuWfdyWXj1OwyJEAHnp3qGHpwni34ugIl
hbI6x/VHgldFhJ0fIGkVIkhngFk2Do7Yftc5ukDxhVgrnFN+FbnnAbHksUU4/AFx
4358+TN9euw+9QG8fW9ue4C15rg2FB74OVS4vZgp4hKHZUbO8dvv/GFu4QZIKYEw
RNnbMRVbHsvPUUD8h6KIR7TPQDsdk5xyM6cwQT89XXH/OaFU45091MiEPSovWEnq
31LigHRlP/lGU+J6rhWHmv8k4Y9LJ32B6yP7EQljQYt9Hb1lRA7Y6nKUUxqrjRnz
kdZ5MboNQ4MfaROEeP6Q/K67/4BvvceLZ9YtbI72v4YR9UwZKsCNntvOHxJ3V/ZU
ygdKJRyesUbKy994LZp5uJUZUXiezsupd0wPIt9ULQ539aRte1Ifyfa4Y4Ko9Iu6
yrI6w45RqytOqsk+fj/3Viis5CsvUBN8qGgktV/9If7FvrOw43ELH/DO8C3MDhGR
LAI/5y31BmsbQdr9rOYSX+5mb87A4yluVgfP/MNicSPBR6KoXIfwthmLl4TF/jCk
om8ngzsAYbMpdHFkJDnz0rZd0Uc98THZSrYvg+R925/WgIOrteZ+3fpU0PPoG8HV
oY8+yqnAaPlzKKZQue1s1gd3hhCp2I3yGDRDlTzVNmxYrsFXAdlz8iadMMWPaWBZ
p6OcoDiRpwWGd+6CnZM8VAmSSBOxXgCCL8OaeukfgNGKhsgdgHW/NtkmRl4gUteT
1THThYD+fROX/iogNRxA8X+NPC0j8/Ey7/LCDpi21plGXE/c77SGDE4StIbTu/xW
szvO4P4oeMBV/YJNiNJOubVnnxYGBHC0NhX+7I6pvxEYw+JYRUbzitEagkn4lJ+R
BdxSsMI7Vo1lper+WHd5mYqm6GLs7NDmKsnvdxuZHDs56dH2GsPLeH168fZCh9G8
X+yKasCrUQK2w5RmzJHAuBMgd7b0av1KcOoPpDRXlNQrjc7/eAQ/xPNJ+C5wRgfW
xjPM6Eb1zQVKtJe0MvSFdnyMawRoCZ1/9KTnNTI3i2yDLrgpZPjxt49Hy+C/xe1l
rdK1/tefhialuLdui3SYtieZYwThE2vPSBztV4Y6kkrjpb1nPrHg/ndl+rGBAR/r
ZMNQX+Psmegm7mZUq17U4oMTu4lHjgaeFEhC+Ai52OVMGHn9bBW+GHRm6Umq1eAy
ZGMwQZq3mEUQQhG8bs0r8Cwic6VtKd/YEpyao6EpM25dZqhpYUV86OTpfwKgAOU2
5TfzJLd6GSOU+EFMghKxjH0iFoZQj0eVrBcLJusRfZEYRZG7f31My6rxGPpSb5gn
KYRoJaki4XmeuJjkqDwIXAEzu2R/MMhFCbVTGZQRiPJRbFwc7lYmtnsAs+5WQAVf
3Q3xTFUIJgg2Ejx286DDvk3nxW7BnJkxlVv7/QslljkLRKTOd/SGKDqlRDkuRn5s
kAXo42MxI//NZvxaGuXomMNn+iOtFEp7p3n7zIQu83ErIFth8FrR3x5T3v2aZ70E
pJTFGjF+Nx6dnDxpxHrpte/SgljgmbjQfg20Okt/GaAqsj++CYTtYqm5lo/wiCYU
+1iD+OrvwRRIetzVfUad7Vf2Kbm6HRN+rIXJaTlcNZFVacP/ybuD/VLV/fNoxVR6
EHTNHGhvhPe/ryFETstrXzZl7P7UtLD9TfE+XPHCN3KTkFGTVGX2W7nwIaCU1ZLu
wOl6lX4mq8EJPhkf0RrBSk1P1PmPwITCCBXVLMImz6iRuu8xsPQSVby92egGE83s
VL1r3Y13KfllFWqz42NZNPY89kBhFah0zhhWcOfvB+Yxbqke1inPGbXOprqpvCi5
zR+w+0TJAP6OOWBxu/gwmf/71MH86MAlJJD+r9oWVJ+4Gwn2abC6YSQD/rAKZEtH
FnRv3aZvd1By1IbSW8/2CORPAxJgVOTfrd9KXC/WKuiocsG22/XlgIbtWaI+l+LC
2OorzgF3Lap9QMlwb0Y1SQdxRkOciY063n2H2XLs1Ef2JNlIH3lPwMJvpZuJUlTs
XQkrSGo5ooO9vQaRWzW5ghI4GornuTEWKE4VPd+6MPbkurMzlP4u2tjk2YZHAXq6
4/pggqjK0+3UJd6VtXsKXoswF0G004aYnmni8a9FLnhNMrLC4Ge43+UiO7UEOHwI
c093jdIk4L0yiL+L8WDy7EbdGv/ebsfHsU/kElLvEzctLHDBcN4XpFkhxf8GJhKA
LEy7tKLQKAAPLMtjYEXsNkK31wNew2uOQsR/OirzqAIEio8kpV/Ieev6Clgp4YdF
qQjgX1Gaq7Al0+YLIPqmdZ1Bka2kN6ioCutotNotYbclTgO7S+pUBx+gb7AO/8Yv
Usc6SiGKgGAOSCYvk9LH+2nEoqdIZJXqjk/88UtiQKZ16qRp6cSft/wEinajJ8Xx
mxrEwTeHVkeONWOm7vap2MzgrdrwkGDQhlU5Xk1WtxQMDEEIFqhTxKdG3cM7/aEz
lnSpLoexQ2vX0sOclRDWNmJDjNQaw1UIWKGdePKzS4bl72bF5Qp2pye/wEZxHglq
wDMjkBpdkQCKaxU8IWBMO5ZwZzrcmyTwMiw3GoM7wt016RU+XnVqfeA80tv9Xnj2
LzQeCvudJRLfnh47awQVcJwblqB5c4qxBBFLAbmxcHe0DOV4ZAixsBovq9zBEe86
UMKrhyAlox3oWq5zjMrQn1xmnOt2c5HdbZlwvvhI86S+l1FRl+5gXnrtD5BGGa1u
+bE/GHAcYl/KvvFeQ5plA2lu56tZw/da6NyEkg9QOttaPAy3z5j5CBEj6FRwND0B
ARtWieAoxCioVOcE+ffBYesGRxdQ1kmleo+9/TOOtBrHHmB+U4bvx9HJ/YKEqJws
gFz9k/TFgjsR03+WEYvySslPbTlvW7dS5dZ8DMYNAj4AwprsCklI+dricL3mC7go
ov1GRcwnauiqC5nGQmoCJ5w1bg8eTESaHSe2rEkOTEMkgiYOrbH+wtBxP7I132hQ
ZZ/mdYVkhfb1OYoKVKPRn8/RsuWjwiEtAgh2zPPxTyH6FmR5kENzJkZgXIiOK4sg
PiL9vMRxbbiX5Vn8XDa6V6d8sxaiVKwdIrcgzcneT97mUAiIVO8rjAortvQIDRd5
K3BpG2TUWiAEiCPRt7GW/5ZTtwILUXKRmfIzLCgwy8zvNsW2m0+cBUBnPMv7o13N
Q84c/bqOOLd7iCIENVfTJW2xX3HM2nopqeFBzUH/jScsgMVvkdBp0p8FSsr5/UgK
CKlwv4gl8B24B/HoBXgEXuXX3qhSsCVjREtWX3sDHQHOzbs5LJCue6BKEq2dykXk
Mt/S3dMgF+BaJq9l6xVi27tCMovnGeDPwiyHtuGJRRUAtGIbDibxRxn4aJRnpQ+0
VpG85V9Bfj5/1gXG3NMVCSxbbdipdyTp2ze5QTpmycP0wmnYGSqjvybMzmUp+kn4
SJUbtBXhlt0XThDvnAaDhkDI5BNrNk26CSR5bw0N1U5gLiE2wyjtsCZszuk6s4uZ
z6W0ci8iHhCHRHCj58aWxLoeZHUirxv1B1TSocM1QBw0ccYqa9YhyPiK86MACbdT
6hhCvVn86ft8QBzBvRC+nR4sb4hyhp6xLG6nZ2tVLRx4uomlxGhrAXYISG7bsDRa
9I6YyiJEeSIaFbV10cC7RdcQFgt1+l8jX6+zC/WDiwg7BieSGe5JGkrk6Cdk7WOS
xWEfIPF2umBfzI1AAac+UgYsG1EpT4WSLpVyM/VvaoDoepjovfYwV17/tqkx6QBZ
gz7LPXqbO4LuGP0PrUCwhIzFdQZOWdJ2PTyeSgCAZDlkhJm6k35rCgBxzQ3OmYpb
cTJfmXf6EYzpyH8blWFcd10JCMlVxxxG82jxKDAtvJCJQj2Tk8+RSDQ2F4Saz31E
qLRkKaFsaurmiPH4J+Izw4+kw5ty9UU+41YqUrd2vE8f1Gvk+HyPAwsHLDqUhAw6
vrw7VkvnbspeLLfPS0LGc4AnVml06cmrhz4nExtQDrJFtmWK+igTazptlSH1gEzO
M3Q3o/XE9JK2ZYjAFG0gZW0JxE2V2g2tY8xiRAAqoyxmwaD1Rd1c93m5hb59MapZ
C4WckTtJmQS23PRNHh1n/6sLrZgi0R3bk7ee9Dac5eAuQmvaFcW04sK8EzC1ofL1
d6xKKGHbS+PGcj2DpPm0A7NgdTDBUceNCj5GmLotSnofJTy3My9g9X4CTBL7jHRv
1qMr5VRPjgjR7Qov9sfRyJv7pp1DJ20SI9O8SIHZWxoN/ygV1v50ePLfhw7spgxA
Oht4BhXbJkreJ3t9SwV5z09Wz/mlTI/HKgPLVnTwNtyNQrtwKoPTZ4U++75Jc8fB
8NJVEdvPpLQtkcr1C8C//klYUD0rm+bQ/xPz2wxkpq2ugTuVZ1pFv+n7cSeo0YNs
JIpnbgZ9cipaXalyxMSIdnILlDYGgC0ZDmSpe0pwL6H1wWJdYwYlZixyz+6HQoaI
EilePQFAirywA9erhUMEezEebXOW0v7GrLXrOQPCdGNK0Z2ut45Re1ddQU6XMj7P
UDYIQLaKSIPCZNyG4BFrqKa95/RS0pMFfFzXepwojcncchLjufrzPwuLNNHbqU6x
e74MhqeTWHDYBxFlCeigCLAUx0dmHPF+XoM2WS7pXZhU8tb2EzgphN8InbGmgTgm
Qvcrw5jQ09ZUDZB10LIIxDMThBenjy1InKDk6TeICvxxw36SL127flFadX4q9TEL
1U5bOmU4NOhmls4htHf5shPnSfbo1vT3tx9yiviMqV5n55ZBuLg00hgKhZ+2vuRw
Sz3TdoEGsRHI8+7A12KFy2qCYhCr/EwJhn3OoGoKoN/hnt3+iuioEvH0rqsGLNk5
NANu4mgmd3hihxfzavPAvE1fdUhei5yTXARFXF+tGAp8HRfgDDsmRHVVYas2n93q
VIZ+IFq0YmH1uth0wOCc6YBA/jpFoatztURkqTMFNhbB3NthQQN6mgAgwVqb4NQx
RtFY07OSZQooAdw7WquyX0w0rssVuVestahaTX0RCzwuzRZiaBqy6ppgwTOtNIzF
mEu23ScPe9PTUIwZ2EAF36NVIBjYP41QNhBgmF41RkSmLOAzXUhNxhfjeBIQFrTT
s6L9eUaIg+QtxA5fjc87XYgIwslOSY9AtfWq31ZJ/vBt3k46w8U4kCh3R6xhofID
EgHXQCaH/m93HtHx/TrXekuhCAZ55z2npD4FwbnckOqQX8lCPIyzwXjQ6DW+6Ech
hk5AFL8fv4SigIl8LuEnrv2s/kk95P+zP5DnAbrbWXpxTkS4T31fDBglnKR6pAgg
SYQLplIXaxZ+LJiF9W1PDE+NsVqjuh6sSEwOfU5BcMUJOEW51YHfBgo2lBBwgAwq
qbtT2jC1i66RbgyMzwD06pMRBhcETiUj1FaIWePzvj43Ma7G3EfgwIrr2yVZ9pG9
vZ3TIRYYrAIxjsdv7bLXyVIdj0dCi8/WXROmqaZOYUGTx72Px3SzjTsD0XIqIeLT
q7StMAApaUKNWYX3iI0vdwDVYdX3YLKC2NwnJnBrY4T+WA8OCAFQj0CuS30YTaKz
qhoFkxZ74uCvEFaFu8ezdExuHweYjPcprPRcxOW83MlD04x6mwAGhJvUKkcKiYwo
X7uT+/gEoqiEg8lQRDhd+JWLeE2i466mTQUCWgIy+1M0aMlTlkmU/6pLVWkpHMv0
SF4avyTyuLEs83KG8s3PNNF5dr3s0EerlzH1s29zKqj43QtVp7bEOUYAHhpMIwi2
G4oVVlSIDm4pDGoPGK3tIBKVaA0g7MU37T3MSpNJJUFueh5odWBaHgdESKS8T7Mg
n8YdVctza5Zxy1i1M+uGqqKGA67Pcjk75vyhlsmdaxCzIULgpqbhl5T0IpMcl33q
IYM3C+mGa83NZ6Rb3s6x/HvQ42LnnLJ+GUqDHS/BN669MDQ/AkC4UY+reWZtjs60
stdlDDizMjH91UEpMsZ3jlWqYP9dzhaiKngQtmmyYBdyHGQqsByyDTbuCUdop5Ao
PcmMQOylNsq1U8NHqSGk6WtbCYr9bTXp4akg171t/5wwb/uBWOvm/kXunHfTZ3kg
VPdZvjP696pIuDmisWXFzFBc8+qjq1x4JLxJ9DfMgKIjIiGeZQmKbrHElNlOi59Q
+q6yr0wtQCniyEdf26TfFZw6QTgkFamkkQgi3WrdKr+NcRVPBjY2BgNEc8+8h6Yx
ifumzhjHWt/XNtye3P13dm3xtZ47jzLZ2B9hFrIlfFzpBY00N5Rx8IoA0FNsaPVJ
kx7DB7LKiCG/daOS84NfGcY6IdnClFKW304LgLeSfSW4jCH/Pcf6V4TNR3vPDaV6
CGFQUfCCTw5vGGq0dqkTVMWpV7TtKFlDX/bJwnOthUzxUH8+9SEG75tNRaMpYk5F
gLpWV5mxSCopiMGuUk+O+0pOQ2xfvcR58fMNN4t2+j4Fc/TiqflX3ZRYGya9rP6x
pMhbIMZaQr0jRrp2zk8U3zFvAsBankYA45ZAPGMiHbubqQ6U/PbW2eEzNx/sNFVm
yyB7s2LrbuUguK0jb/hfvlb0vHDWuFCkbPjLIQPqW3RvMiKK9KxY7ssuAmwxJCZI
/NRrz3CH1TEjgPpHmkVIWPJL1icKJMesFdUEVX3ITyeVZ7JX1YHcI32wQRfHW4dm
pgVkwMq5sdokpqMO1LYc8PGnvBhRFkwXNsO0cwylDYVvhz+HJ88aLKTt+p3vljRJ
aPm5QHVezbLGmhiU437j138s6hIzb/s1N2ixvDMd29F0OZk7keRUK+InYRpkcYV4
OhMgZD7Jb+sT1d0hHDnPEiGJl46vc/dPSq64hsDwfDZ0VBjDdZAVkmB6iadosfjQ
WzZ07rRwGE8SgSr/eTNqUZ/XovucfyuJcAkhaFLuCgwQjqGoQ4wTRypc+lIyM7Ws
hJ7DECH81ZCe6KSB+Se5AZd2KwKJyk3LQL5i5/VJs58dDH8LByFqWniMgMgNratg
578VicSyMdA1TTmVUzyn8HrO9YsRCH6/Ceemb556Tg3h/DK0wDG+NXdD4KSHVtE5
ZHZEg9xxaTnfpArWvUp5sbcUrqQk6OFq2JR4KyqFSlsmMuZrTNeWrubxSQmq/7Wq
Y2vupbUwGlmMopW96TFsuiPsgAWVp7LbnuqYtjLJ6EhkigGYPUNxnj7Q7KAFL3gu
Tq3Q0IEql95IyuSIYaiAFoGPqdodgFv1IfanZspGoHoUGMDuT37O2GnrrlcCeMCG
azRUkhjCEQt1NiE70wo0dXmm2PyuKmqCdvnpKtws2U5y/X5amVW5mc1UtaH5jxRK
ifHSJcuI82NLZJxOz1PnyVsjuBDezIy+MKgDGvJ8JSbB+lW9Udnd+siDuE9OuqkU
KA48hQrwkjlo3AwPC27Uj/+1GvMibzAQ8/p1MRN8QARDOh1Mfu22BxlkGi9tb2zu
XPUkFGcnJYBDFGd1AmEZJ2WijJM0BlrM5Q6q/rzYeM2a0PCJcwuhPH4YyMRs0d66
AOTyE1xdNxmmtSe6XVU+CqXbx5CCgagOoObklOExW2J69w0m0Ozk6lpyN8X7hVKS
ZxGa+NBgJPrAj17j/I4lfGpDwEY58cu4GeBcAnNG2ilWtKSL++cIZdva/1z7v0km
O5aH3AXNkVddwghRwt8CLznEgeI47bc/np7/TYiS2whmhY77WFHwhl+Xl1B5KDhI
mGSCha78SuX25+pWOFq+JpNqcRgKgjtry5SGvwB5Iol2SfEiRSfnIeNrYU9rCUaA
9tTLCmdvQYPhUhrRUxzAOPvZ6Uir1ASE2TRyMOlJbr08948EoGMx12vE///6x5VH
uToRHRO7W2SP8OMC2vYnFP0kPrqcg3fcahlVABYLZ0m1pc51Adargjva8vSlNM37
4c5vapBnehOVwP4jfyUc168ZlZz8ExqWBG2/JzCthalI0v9e8C/IoNcHEYlQuVM9
8zSxlL51/GClGWG24zQxIyhJTwNJwYmSigIfKL3zuWeGPN3EbObU8ci7qWzV7rTL
ZY2KHulsDxiJJSpdgeYJgCWOgcTx3COEPVKxWf9ZLsxsTxfWBFpI4Yu/Fc9EQ4gC
7S2KltGb1+tdgp0WWPfKzcXXSQdw6PVvsQ9pai+DeTF3z2sksSOmYWJv29ysQtZU
LHEIuTSI4AdZHCouHSa0UU5UXpH+yBxtgnbaf+LpV2WmcvhpqBBp2JKEAHa2NcXa
AP6ysLQ/E/KxHqJOeUX2Zn3XW5Keql+xmb9WghpxHft7zsDYOo0LdfW0+AF+H88f
gxe1cf9vmTBo6J0g9+djZw0GYEbEahfJsFi28z5c4UG4YAwE1N29eWtMVg1NzMBy
fzQ6gSOeSFiZMnJOIPmqCLTpnaLy7RByfzRzjYVJHd+70JWKwkfo6oJbG63UGICr
zxgXrA+vzbwfPnpt4QsaYQFcPa8NjzvQ0/hkOxnbLhwMXnKAbR7x1QzAN3VZFH+5
K+Rag9zj9kXApGnh+0n+Xy/nGMuuaqgh/Eaxg/48n2zm77a08O3vQ6wfiPTLXptL
jOYcbXaUItM1MfhUAtWFXqTi1X+R69VP8YwJJuDMO59p4bqBwKhoQts6IFZ4caEZ
j7zwbNni7JFwtRFLJxxB0Gbn2zb4z4cBH5uw4P4/IJJYSP9Q0AXQ9t5scmuqKfKp
LbfbI1owhms4enT2GDF+UrWz+oeliOqO4UfDb/QafwlNE/cj7kLagMWuitNypvzl
PW7R+SywcDfyC7tJ72yNVgJHYeJVwodOJvFGDikPC1ucTvaKBep2rtNmL8/dpgJC
HWsEGRa9jcWN9EenTBjN1S9wlWeYTjE0IqMML+xXQQh6wxGJjOjUjEQnNzadCAZg
puxLC6j6kK15lHn2DMXUnShmCbEvyWNq1MDnAh3R5UWG70I8OonCFs3+ugMu9IZz
3fJRQ0osybmh0HICBDBbPGIHOqIJa4ghzS1m2U7n/w/UO6TDNkhtg2nW835SStWp
zELTh1XwVf9sXgU1B2qUTfM272R22zDCyNhq/k2ky0B9/wDNSl2Hfc1Vxn+dsx2T
QO/v/Xx1mEf2JfvOCx5f4NDThOmF9ZfrHt8TYFxhvE/KuArfzPdmSZhH79YMW/Gr
NyBcAeM/OaR3ihZJ7ixIXujRqEDptEAWeaBGYg2H+NUOdp41EFb0mHLMyr+gs7cx
hjC3Rpk2mLZ4yOoj7HIIeogjnQ95HtiAj0GaoBwGxxTbr44dEGU0pQKbkaOjYl3K
vY9B55MAPwfz8jyKBcPosGFF1OKz7GQiD7LSm1UbPZT57aQqwqX4rYBZ+S1HUpEz
R8vXIRu/RM2bPfCMXaVpe3Kcd5IqEEM9WggqQmgr5q0FJ8KXHnTkLzn+RmRhNOC4
5bDalGZwEgMRvjeYN44SKm+ff84qqKNvylzWk6wmlRPjb/2PEaIboXy+KJQIU0X0
4eDDuJPMH9QPHUalvfijGIxt/VIdRYp+6BCe5xFsFPrzv++/uHECOAp/EXH5lmwf
hhVrqzLc8Tx/JaSuGifrEeN0Bn3AxBaJovu//9pOaPxG8N0C2xEFY8q9KUWMz4On
kXpGItv4E5J1xt1a4J6p2Hfl5d0aPQwcoSGsi8lu5vn5uHzvj+Z642c5QZg20/So
+z4n/uua8sWHTKxGk1KRJdT8/htMraE9KUojQD96tskcxUxXOirnnnmra2pcZ5se
tKfFsBMaxtX0MMpF2+VnRz4gmxfiiBQxZDuiKpRsvCsJTKa35GK19PirxsUuz+lp
PtLCabJXKOwFI1gEfJVFR7xO+D7+xGSldL73sC5vRjTuyxPR/DGe0I5M1uZq7Zgb
Jud5ERmk35pcePxmknGTD0rQ2uWADHZgPHyor84GvYlKbzxaCTYzvyZ4IulLQLI2
xoZP5FGI/JqJUNDzrods5qWQFTJiQkVzwSxjukFqTFIxR7zo9yCFK53oe31ydogY
TvUUBJFf1wRE93JkkGqoBpvUU5PS2/kDR6WIHeXqTxwKqtZSD+vPjksgsFUSLSyU
bmDxWErv4RVF2a4Ar/bdABSMDpa8WOx2+SoZaOLT7pZWIvPGGrOeKLEMIvkr2PyQ
X1p12dEIKSgSWm5dfFWgTzxRsACa6PR1rpmpkbze0WeIPTrorVIgTNm6TlT+muAN
yU2z19RALdtItZ9fwH5QCbzPj0VaOQvWtOMbNJzgy2EqP2C0ip5mMV03ZQtYP4Wf
v+kVj+kB1IWbuMUg1NIbKUCE2ua5Uv9HnbP3Tk0SrNeuuWULWc+nwL0jvB4JTni4
06KI8ngXKsxAFDJ1trNUt34Fq3PmXOTKYMmKwSAcOKkSV0yQRGVTdqhAaRnsfzee
uzVGuQzdwpQjf4eM2dYRow6vtXpMmUAkLCdW5eobXwn0Qbz/WF3N3uVhnf0QPDjl
hCUz0Ou11fhq2eEj9nNxGenMN3aeXGXDBwGBRkT0HUYg7xP+pkVDUPVsm+PWTgin
X6xVl0Yc2mM8LGTl8koI5tRzqDFOnXo8s/afHs3rUAeDHa4sNyyGxYWUW5pq9tDA
G0IFfXttq7aECuJxfvXyaPfaOJYFFkbHFlLTW00hGUo0w9jX3Lko5tGCmHcY/FHk
2Vs4bxXZsXyhzqPGU8KAFHgCXmJc6JH1n/q7xitNdlV6cBQVUpm+rl8xi/h6y5pq
JhofLGIG+bwT5GbPLlXro98d2I2w7W9XSG/Wd76FqMkK+62Ft9WYPDnsk8AhNIKT
j6xP5cQugRPMUj7hv+Yo501fO1oZcBpIj1r+8hnZki8EVIAGmwQtYoahT9spiPT3
2eETwe4eoUmtPKa8lmXM/uRow95VGX5cyi/hu9sjZGqyAfqjJVAAT9vIBfPUsl9B
MzFFeLy15QcbIES87HDMiQLlF7jr3tFRwaH9YR5cshUpGVBog2CSkQU+oULSHMJg
UY41RckVvpghA7yFpKSDCRW/qkgUqeSoiVD1mjNo0VBJ2YSnkKjeAECmPghby30a
tlp94PWGkvgU8RjbCYfs/PxtdJewp8ZfKPNwjjk1St7Fy7lyYAl+G2CvwJbZ2Pdr
70YBUorxv3kWrup5UVkp73ETp8UJ8QGjZoFN3I+GAV2ow9jUourE6CrbQ2V/vj8F
F/9ff2jW4cH3SFzTnOOGIecIcfIiPybNxbKTGdj031aUYwsY2qFUqsC+jxDWRz82
4ooPulSQUUA1vp4NaMUUsG6Hj069lsxEvZGY8xMKRHpcKrYNb4BOuel4BwA3YlX1
wC+jsC6d/XEDjubz/8tzhCMfPloqrppLJn9kSyhL5iy5K1Fbp0N3e9JvBdaytqEV
BWdAzhYGsGS/v5YthKV2y2nfur6YaA3mNIaXF0Cjo6mcCWMHemPbOyK4UvTe6pal
VCTvA3F0Bbc2CRp/O89aqW/df4uQhFNHCTCExfStYrmIfOLzdZfU7DwTDKv/T5jE
CBDlkXFR0BZSUukVnWEbNVtGrMr6yI0idIOECWSk+8wwQsJzE8AFjdSJpGhe1GE1
vMIJN9XauXXpmLIkJX0OPbRN6VKCIPPRkhp9J3xfrmLSa3yCIB0eq9paE0uQLM8j
p0bhwcC/fumz1GiUOe0erwK8aONc7elRC1dF4tm/yKPW8Ac9453OvLMGoHeCPdET
euSA8RozFesw3lyS6bcZIwLha3syTC64aprVcV81Q02MdLAWawF/OIlAyfzxKhRR
dl09Qk4s26uiMD6wANooB9ibQU5I9qurRBukHhvNcMEtB0/gz7J/3nJOm2lRpQyr
+DvvafB4O1bvE8U2P3rlh4iZ7xmTWKiihkOHSTXyhVkVqmMcI/H4ZpAcFxIFBdPU
B6tv9LUYlIq3t3En7VMyymQ44x5s13Qyo4PDdKkQHveMsm8fdFYy3Hr4W/kVk7Q1
M0pvBZo76ewgumBf6f+gE5QvBnCxLSjS9hwxborIGCJmuw6oAY8AeuJwYkGLakR9
O0whRQ4hU3A/XUK/hGmpI2KWLTGggeqn8nlz/a2nmKOMMsCasDmkAIbuQhPDz6/x
bUTvSWRVM2QZMY17sE0nADshqlvsPwf9W1T+Nw2ErSLW37r/frE1swfOornsQQKz
jTUeHv5vlKYk6Gu0RrqwXPN8NmXQWyia7FWKdiviKX5ycb8l3dFFPMPoS+RY59pX
hLjdyXMMDytE+W1WAlq+5JzzvDpxY4HvfrSGcctpSaIi60S6Ba7TeWRBIWzAyBql
ujaMhtdhxAVx/2KY0sN5mTos/QKNSNzNZe6hv2wMhlELzl1X4mCZiy2/rssANPD9
Oyp8xTnyyfkl6qWYJQ7bmDBsJT97TUap0nBB2+Uqfy7doTVR+Pd00lfaMfThTTq6
TvKQHWeU/fogjfYIrnQCMEM70v/pZrWrW5X1w3mE6bk1i/bsKMINZBSXq0chP3WT
/2XAb1we0y5dun5E/CJ9p8YRC3VrD7MshRYGET3uV65kNkrzBX/VKLaA7j+j21Fm
b1KfM5jxnaLJAmwp0/DOxhMlvFxrioeWAutLZ2ZEyS6kNIDP3LdMIoQTkD2+dbmt
DDrAVlx6q8krSi6J0aUPCpXbqrBOO9l6vmHbpVEdYvk4oR21LgdWrTWDggqdjOck
nCpLnueSHljFtDQKgsdoFZfneFLXwXfOlfzMLovxpVg7XURuppwsuoypzRGkY9DL
AfqFUQlH3AX6XyCnwtXkOgSBYUqIuVA66Er/KL+bSA0MnTsGPVqAGUal/D3+9wlG
nQbzM9kZ3odoPmoNxfq8iDUZ7NekDDyMIIPkpsnOc9BZJ1HCdPJRULBcF/b6VTOH
U7J8HLiNSHpOAy7Ua8sNzcY35Z8vb0h0y+EGxS4+G2rTVQOAJZyZ9tgwjisV0GIC
zfWuahKD11C2tCDCajMUnkficT1aQaZlyL5G+7Ue+V1N5Vw6S88sCrhILvDzewGi
TDij3X0NPmw+vih7PxjhhAIAeoYjCUY5+INmeYG9a2hNxSJl/mx1XhVrotePTulV
McN0I2fI54CDc5USk7cpUTG64CiaiK2mVw4BPSL5TXaTD/m9SRrzpRceK7JvFxC7
ox4Fr8cE6vFN/KdGypp39Ai8RrX1o1fUqRnCqIiS0ShbwvixBjgVt1pVMWFNbCf1
eP3/XNzLB40aEfWVyuxBmgez9AXa0JW92OlMC7v1wyAWhMhulkTHh5Fh3870Qlrv
gFFTpDz86CVP/rmRpizYHBUohtxrW+27POvi551K4NjHabJmFinbs5oOKYa/P6bM
i+4y4ZUvFvBqj/A43kVEGrOXooRxqlpD2Rcpnq02DHS5LtU7J/ln0wPlRCKmY/h4
uREkW2z/8p0omdOow4+yJ5tt47Yx465DEZiuGedjiAyG/L6cP+0WDckxLpNgZFMb
glqsdKc8ouustEIDBBKq22ZmJlanlpR6g6PcJocYY+szREbF5SpaUCCwoxRPJpnm
24f8WKQOoDkTTZPV+5/bEDqTZVJaWFQUNEQ1fayB6cNVWYY4sKExix7qH7C9sk4n
1KMRI3e8k5NI2zeOZnNqUTUwrW6GpQ2EoIq3RGaHhfiQMQI1pZPSpLsFFCbN+Zpp
WKilSom6PSd6S1KJSzOkpxlDXhZF6Hh34AH9MlOWFHsscO7ibMWtEkHw6eCpuwBC
KVrV2jwn3tM35N/5SUDisQ0r9qFKUqJ2tMVd0d4BHpTcgX247Kn8FVBiPG6SEFXX
scgv1iGZEg6zeQAPNU3bgUMw0Zn0JohrhoTbilAKgztDDWz/6fcqeA2MrZch5lsb
K8cOVTKpu1Vr4ChBCCLd9j0hYLqpaBue1Dj+0kGOH22U4K8NOn7RAINplPI5O68z
LkWgcdxyDVCOFitjEVvraAsLHGvH+gLqgPfMoShcehCB9fwNe+mn4sELeAzOXJLi
B4srhTVCR/90Qfe6telNPhbJDxVpAIB8YgQwVhDYZKD7moI6HRu1bOQvvJ4dKeH1
O3HWqpNuWvwTsNZsWs8VTWVz/kryBOb1kqXgDCSoAAkLkC+MHTYVKkNNBLUCujxp
sY3ayw4YmMvXlpzjLt5wUPIk5GYpf29gHvmzxKYfOFrawVvUtFT1pbUHW4VMnbOf
0dthzbO+WJfGgiYX+dT1yJRePlVnlytitQA61CUZ9iy6vTzQwgOF1QH250gOyQ7c
Y5J8/tSWiJITEhzZnq0Pd8MctXcMZf85fz742MbYZX+HzxdvsauYvCC+u1wTOJ6r
7hjLbRn79STkTdGwQiP0PJ3lgJm8TONGqgLh0BuxUrTFci+mHfu1uJQF09FV00qM
WiM+ICI95zjLUw6rDQvZWRRKYuIxhYWpu2aO4kz88ny2612eXcSix0fxTAf1Ropa
yUa3SglShJ4z8ShKQ5gX7lROx/kzhUqOQOEbmcTaVKwI4pKMipzoKXP48asoNXCw
qSKNgpTlU2u8dYMee2P9pCXxJ+pzE8kqAcRX/KddOql4sUxpdIMlICchscwnORUy
AIIgPFtVZjWCstcX+cuVQIS7UGuD7pPVtpMexAabSpk/YSxlkEIyjHkN5LD1LOgx
ZBZSWmNLQdByMNBfQxRWHJtQ/glV8htYwhN5huG5O3EJK831UAm/Wbv7YYJQ1aIW
q6RsXLyySNbyTrbzNiN05rHdQcKNjxN8GUU+oL/l7vu+oc6UxPGhlEarRPItNW0q
b20pHu2n1LnEqy6+1tIYsPhCKvjH67B3r+zGJCloO/TGye8h1Cnis9pX/Gw1hLT/
WHgMtn744GI/+HVwKFGFe6MnS0rwJG89nN2rHy2JATsskMgwUVANUP2D1Dd5W6h4
A2Ax6PRJcR3Ao/XZDxcquakYy5jSgw3i84oRz8jit0utz9wuLhmMWEeyiOxYrwoK
rWnjNhx3ALPJI+a9dRIZMnvzysgHOIMktOQ12PPNNx6K9PICBPifzv3Bh3hfFaV5
V3q18dwtdhEP4kU1crvps13P7yo7FE+EZpLgsve5Ez6KyvpWTZMEmg2s/ENh+Cep
D1K3cbt6xMX/BnOgjUn2/zIBhQ4VHhaOxIZOrpQNAoZOBQyy9AVj4yAZoLVWpoAV
x8X2znou8GnFANTijTKmUM1DODuxnwZzF+vLb9zSXBS5mEAIiXREEz3vZQH2nx7p
6nfUE3MjkK0Lnkii1qN/4dBOC7mBQcPAnDCFbMn6kuSjQzPzGmLn2mZjORPSxdmg
i0DBXxpMKYnThrkZpJiOXDEaJJ+nxJC3ieDFT1/SlXzjRuPkXFN+7mRiADhnFN8U
W9RJKq6PjnZIPUJkIP2Loq3HLVi2voZgZ4mXbkDTlpwaQ+SlxHAEvTB8YkliPyTs
xoGVBw9mJY8Lhzlx32wt0KoYTu/76QdV5x+ofhYKaMhNf7rWe3NfcBSTOil82Su7
EkGhaajnIySh6wENAzTmxv7Q/ujn0PIcpHWWVuSGwehhvUM/ClLevP20WdDHL5MK
KlPaUtv6Yiwe8bdaNjVXGsSoiOFNzurtx8GyVOjL718YxM4x0Xr64MRrhdzmkkg5
BjpuewJLWt60lK7GQJKpsTEppRnyIPjCo9ugkveyVdaghpafpIO/ZmJUY2llxk34
qdnTXHxfIqXYK9inFmyK9J4IQ9EYGig+V+XvnDx8fwxYxoVtYo63oxsWmi6SFgti
4tXZF+WR0ZDhepHaOg17+euRHKsPxQiqg8GfjDGcMhGIDXnM6BMoKlrVEZpbM7Yw
W4J+toiTPnqG8JV5+5pOjWLnfiULgwwrdzTckzkdr6+MCHszMEn24H5qVhPSgpLF
1cx8DRGEp7PeIbCMFioF1NfwXup0DZnHd6Iyu6EKdgreo+NGE9aPOZlngE4lp8Q1
x2foZZ5npkSN2fsO5eX/1Ddk2NCY0D0ZeaG7cfGoJBn6yVI5bcr7BYqmEhDwDGdp
bi2apVitwTMOJ7lQ1a5M8AcBy45tX4zrDfu8HbI4JCgmxaV1baz4Y3O2dDAe89TF
4/x7pOCVSZbZkafjLECEEoRabxHupo6VY4P9wkr20NL6KRXKE4KgH9S9f4QdWTF2
l6vPbmh7eFzMjFEz9OSz1FBzWmz1ScJfLcv5DgIkWvCYeUncNGJx70nMar3CYneZ
chqRNgMfS0ajOpIjrd6dKP43e7tKgmo8IpUUBEpYjzOIqidPiur1ytJBBt4gHjTX
gEeaximrFkIEhJharXVOt7vtsa7VU0XQDlkbYZPI0lAadN16SZ4fbsswXEbIc8b8
jQ/iTmeEGcPBJiHKkCYaEkStFM0Y7vNrjmdPI7V8Sn+5eQG8gZS4tUJrIM19xxjz
j+VJvx5uq7CbcGisVR/xM8lzK++b/to/2r7e6in6ZybrvZrxOj03RISQnyDYj24X
Mf2kSPhoN7iNdLprmQEa1nZj1WBxD73RymuxRPEmLWm6m7Tl0RtLaJG5EhWM3lMd
C2sQxM9wd/z2KuFjjQeEnu/R2qPLtN50Mw+QazdB8lJhxFinQcY2ZZ4XDAXfiD1/
jJlN/MBXB6ZvLrvsPN4PlGhO8RgliVXAyicDOVuDlhEPFPty9IqPZdOIFIvHpnGn
fo7XTitfLIlP5wPcXWbQkAv3A/yiwgY37Hy8oUvQ3kzBv9xRR+9ryuMRtdgPn+hn
WffN1MFVo41V0NFzbUKrmYxOJehLfd12vLvM74e5Vya+RbXuBoT4n7Fq3pzpAP/n
xFMdcbDYl3/W1w+Y/+jIsHDOC0ranCx+dO1B9ljTXMKkh+2WH+aK/ZH7iab1JEKL
m55Jo3/YkC6yOMvoHWOkkcWC7hsuTdQYd4mZKwrCopvJQq4GBacAu560AruX5Nx9
Y6LlKGbRNEJuOOLYNL7irTgDwu8t457pKLM6EEibhvJzzkzjUAZM2OVyVaLVlKwn
1UwxgzR8i7AYrOJo9YO+xFsS8PMHBTmaHZXjoY97UFRJ9yHdrrNiwPG/BvFUyocB
l8JPz0U2lh91HF/q1g3VqfbUzF7kW8nlNtH29yo3ntsQSYc3pr0o925NqDxfG4bk
dNpfqG68vBdxg/TKAtz8xfbEATNE77GMro0E5yC2nGZPGXzbEYs7Mv4713zxLco/
00cA5oml+jVQ4f2Ek3wQLqKrdmj6Wy2LGeWAxIyPnykPWQ1xOAd2SIhP2NIKRlci
XBgOL7zl5WufhQUeMUf85VzaKvWRrVi9Drgx2qZgdS3nkhfplZRYf6l/y+D5eUIs
50760ahujSdW1Xarwh82B6VnRx1LTd8HZbvnsmGbWxaMezgcRCkXvzeKpTFd0R4/
Olc6ncle3U2TwXjLTGp99Kt196lOsNiv2d5qZuoFR+GaCNOtI0c4l89lR+etWhDG
uHN3dcc8YRbEvVYmnEg5PI+1AYQouCCayQWh5cWks+IfpKD/6aQvApRs6xPFS2ws
hqXeahKs2amW8IqjT5CX18nTEJ+7SqGbkIrQeS9V0XfAFRBjdxXi8yY4nlwKnKXD
ILFgTrzs8BR+9TyNo0P8YdI4VpLHQd6dq1xophZYMHrIORrOV+1I3Gqdrn40I5FA
bvQRwZf2u51rvgN1qUk54dcwo/mCAlxYLNCO/QkqZ2gTzRVIXTf3wbV4+ozwE94J
K/cxBc+BKrvjqDxUkWaEjhjNd73nANNhXeY3APZTLlQecDHLT4i/I8w9NtsCGMZs
l7zEG459yVaisPts04iYCKzWqCZdld/FRcAhy+kMjsPZuBj61LZJfHfy6KZaUkUh
wgqB+Zu90EaCqWu2dNUVadRjEWthrlx8TewxWRPRypWf/KFL2Lu26xTWMMI3zLGd
Ur6sn7Ua5VjdKNH2AgeoRkeClfRvDJbVS4ALhr5z0iJQU0HYNhbqa67QWT7vwaXL
Yy5GJjIs2ee43s0sSeM24Lczy1WzBmwulTsmFk5eq4U4pZKW6c9kkHEaLirvstky
3dqsx+aco7lVjmY7PuquGt+zr5TvmS3OuCo4zABVM5VGSnehvAY/pgpI2QDCG+lz
gYWks63b7TZAS3e1f5QBwSl0JXiX+mNyppOiB6y5pw/0HHjVJlSAZvAfiszR3svG
QWBYjICwlbUJKRJYDjr4Zh/KzOYMupi8YyGcO05BbQL8xmwW3RbeKFbLZsYqtKgS
S5zjzCJDV+pdcR0jEkA0FTSDJ1ckZTEJ5fPp0zUZOArahM7tN+gsQD47AfUzCcmt
cJpSIPA/0T+jIWPl+RQPiddKaBAA3fNjw+asGKreRK/svbfyZJqE/lPlbPWA2Ton
2gtj3gUcs4hgiW3nor9o2pjMBBRlLbT7sxXSqJq174AU9ISyZ3QQiGoImSFySrQ4
/C4nPCp79KYyth4G6MjsVovM+hge6rW3HuWKZstz9dVa9S+J+aqGI0Fojoc3cdvE
fujvnHRznrF8ZNxNGFuPW4s1R2vXp6AxVughm7qeEI58eLVvPcSwRYnUnVmPtGXc
2yiZAW9mUjtmQ0rnp1OwMf9/tMxlaMxcNMJoUNalCaZFDTmglitc3cnMc/Zq8Neb
MsXAa/TJSSLdiQ64O9qIILD5MyIxhj3Wz2VUHkkJAInhe0N96DNy7pdKR5GIg/wh
IUQTPbg8CPnAnSUwGHPV+DcfgXAfslxMlEz0vskkA+zKk0cghboUs6YuxSuzgcXS
6zr/aTJIhgoLOqX2OyAsmE9r5bow7j+eysO9y2H0AqH18M7EuY2KmJgGQrAyLMCp
QBNTXjJEwQmnP59CDG2v5G830xeZxdEEChKX72noy3XcowSUN64kOpOb1YaTzGEs
ZXlwOQ8LcsoydlNsCmj3JIZFtRIHhuwt73taC/SfjuvJDFSyl5Jc7OODBRNTf5RA
h2pLBrecVM8OZIF6Ed2U2MNrZdWingMVOiyJ73lMhxopYc38bodDx4uzfrH8yFnL
xSdL0M2r4FqmzpbnsgjMj2pRdymW9JyWxcGhdq9620+mYKo+hsJbk/V8QnOJUYTq
Z7pwSF4v6mw9iivZQDQB9nPQne1sh9embL++XjOHhII7W7Gu6oysf5vAj6M6KePV
76r4IW7/pROgyMZqRNYfAW/Rcd0utgF3/VqyNAhq/5L/hpbpiAjkBowNAGY7ROh0
qXIgZ8zpD02fDntAx6LWtwnthB38Ap/rOE405BJi7wWHxxBSH3cL7pnIBSPWBjXS
zAD6Hq+F2yLVnzeq/ybtRkIlIkDkHCCqGWzMn8vv1aMcZrjTCk14mXfZoZiq3azp
oBO/14W1vLmsEuer5H+axxuSaR0L+FUP7oTkDviu8tWAlp0uJgTlIYq6IsO6at5H
jkl7o/5rzuKJl/K7I5HGH8ck2DqxlmIvX3iKVDYJovKjLNK9zEnNdKT9irwEFcML
KS1d0+lg5S7dNc7DZmLnfLEWU8mNmMDz2bOjvHlx9hxBsBCJa+k9JTbKb0ng6pbe
XVB4gHTuavCVOJul7sYwfC8bcFEPo8aVwOKSMTBK5L2ilDnAMFkS76O1bH9QzuPE
KWxFXr4EwBQPJBZfIBLH/p6DwSFAQUxf5/4r2BFZeU0TnFq52QJovTy47+F2irII
l0vcyCBt8RmUcBqXblupHnJO0Y4Ej61rLz9DkCctOa0R+D1FPTGYpY6e8IY/uML2
0ovLS9HcRzmbYwxovEUg8KA+VZFFzaU5HNcRjSUeHslOdYd4V2QE20ppWTIv3up7
wnLv3d5Z5MGWVkeg/su5YtQQOFBIudTuyBrYZ4XsJCmnhAVaUseHtiAvbHauY9P5
3bVCSG6G3l5Gf4MVHOubTQpFuRLaPUfw5LEAR+mDw/UjjFR0ZfrOMCglmMWuqj0k
sY6T69u/V24oUb529UVzkCvvF84u6U8Fn0VxdoNiwQqMi94ZzmaNvg2Hy/wa4mfN
/yHgV3IkVB7ZtjDYfnTAG1JPY8QKTIRJPDrp7gv5yr5v7zo3GF8sSLXbccvkpJij
B1kUqgu3+/IPws8haeLQufEITwpzgK9AFuBIoELgNXy3W6DTO2sM9R23LwjahI5e
V1U8rsSg8gVAhOQw0uVdCuDNt66sI7LFQ1pZ04wywUUjyUKs7XBoc0QAkQIkuTh2
WTGHdcn62FLkQfC2wRd7UNlP09Xkr3QTji23PJGJLBrToEdn7uD9ThdyT26PvYHr
uV8lxGzVF1YDMnE4e7LJ65jUMbIY7uMzSY+0V0BGUOFc9ehT2qLsgE2NoyyyxOJI
vOvWpT5x4XiBsAxeFVAxynEaBWI+rnq5x6as7N/FuvyjuwwE22ftZJBzIlyOPrxe
TLlPFXOk7SZbqhpWeqD5ffCgU99/SPq2tFxwN7H0SFBATFvcP5e79buYWkqdB/wZ
jA+czwog5JGbPF7XijSsmkvioIw84xB4Q3MxkfN845rTSuYt49LIZPcNZS+/r5Cm
Z3xxIGdZjIcXRQUhqy9HbYyUoGAePp8fTTBe0SlYyPUXnnCnI9ks7/d2f/YEiBCd
TlbYodqNIG0NYRibToh3hKIJk8kL/WVlktEQF4gzEedLO0Ofg39HNw4iRWKFChlr
21HjVE1GaG8kVbK8RR1V405KiBQDMFgVW9PUVbmDEnJUl0W2DAJOssXYaD27GBcH
Y+fnpVXCPx0pgwjs7f+kBCSjVaGN+YdOy+3urBTsnp9ufJMcLgdv9e2gPZFnqTYb
orDxpEin9aXqs8CujxK9qsizUJ67kPLcgNYNuw+2oR1pQcV+4as7eHegtLDg26Ds
qa+WCjKXPmaHZ0W+i0dEDtlI51fbMeeiMYJEDQDLhlPAjrC2Rhfu13fFkiU8+dSA
G86r0pyA1WCmVg3Bkw6M7+8ttykHMkFvf0rI3Cx+Xhp3AhrrVZUSxYYdPc/u0iFH
0UJy//x3voWytNej/PTrMdJmj4sugXed6g6njYdFgn8mu+ARoqwjYIitFxtTOzxE
SAWBl/FZWkZJVA6CnZGXva7Pfj4ZR2NuYKzIqE/6SUcSZHIyhfOuD09auXYSJL2R
oLPBYua2jf4ePvMzKKsv9g8VVb81xaRe/QmgnvmBFAh2xwg05pgwSe5N60JHteSP
4P2vYtRGcA8usgo4H4VazyyIsamawpEdsaLG4qIBugP/IDXGacYW6TnUu4K5t6qy
C61V3CWJTufbX6eD6nEawTDQlqJNPGRnUoPcZaOFUTVYBgQ7prViv6pti9jqk0Ia
m+0TaZd5iSvRvezJk+d8QKlC18NDzAjGs/WdQtItGeu++ZPrXA2Icyl8k9lYjdpF
wvF+Eld16yi2waaHO0zeUKBUwpIC8G8PgYtyGaoX9zF51KvmwbVDwm2crE3NvgmY
k0QDIj7v8TtqH4MnL74kXeW3QKjHs4mcEeL2/25fC/9niRoODdwC6EJaq9hIhcRc
MQadAoVgQLM2G+ACM1r9xxsDPu7ovTLBnCZOxJV2+Bn95fla5wOJ1cUpobE8ljDK
VhfjDTRyiRZoZ8eQzHvZYnN9sB+7tffvG3yZ+IAdyTYCHvV3NfbwWZF7kosj5uxm
Ytx+gzngfNS0+dv318HyVdemyCv17uceCVxG7y63v7uW4sIvHXm6mXH8zal3REmI
az5rtyHNJrlidqwwygbaPk26wYswm+uXH9Ifw0g59TONH/nQe//61wooJhKrY9r1
F6I9Ta4TMlFL7KUYhSaq2+D2euaISDIFNDzND0kxTpZNpnd6/+W9oOI6UgKqRaq/
F4fviO+aqiLmRzwIvmgLM+0Pg9bsK3CF46fuC3/rk1LcVAwMTX2gu+8BJWyo5YqP
JQ8HxbBUaKbahtAuGltcxN44AWMd8dHhxK0+HH36/o6EdTMAnODty4tEH+Kbckof
i2yVRhyVPuLINjMYuHWyIOj0vAfEPXBqW8zMQndjIGpq9f3lMD2Lz5yd6wJ0Hyv3
H1/IgBzAUm9algkyOoN6MR2ABZbuCDq97u+dQ73NnYTXR65cJZE9K9CcPQ8E5DGF
aK5gfqUYHMe+jnhOup+1FUZx5VjwrCjyv619mEa3kEUPId3zWRPMH3Y4wZkAUY7f
u3bHFO+NxxVPLGDdavw0rq51sVAOJcmhCm5IkMQyt6J6J7Vc+2srrfz/mYD+foNu
9wjJTnvbwv9qKlyivhdAWODs1TJvXlEfDErKWdLrhzXf9q/V8nkRgcxVt4bU5Vue
BJsSJmycXL6dc+ZsMMBWe2z8RqotTW6zrs7a5be49nBtKeWJo0IdXAXsCvWQGqJl
IvLcGF6c8NDo8l/z8OUnsYmx5IZMHIoXMvllm4mPIR6wA1X4So7JoYoTnRNpp8vp
s5oy56utKjTe824vMT7NeKeWtDs85DdMf/X6zMH1FOFCo58p4N2HBqWiBc5YNxtV
SeyNDhWF/uLnej+Hf60cPGoVi/O1nTJczZQwIkEFo1+Y9txW5+SNWGD6gvaUBgde
6HxJlOejSs2KeQrHxhdR28MigLB8ua5+ejyF5QN3DkGiAPBPu+UUI7Q63bOMCZoC
+w3cKm16rLcbBBKflpyHNXmOhuk+2P2Eq+CjMLh7wlTBSJW3qyOrNAPLnq39x4I1
vD0CSUARl/vKAdzbfPkN+dO8ejFUOwwa4tvGR55vtoe0nwI34IXpeupf/g954e6O
mk3ex90MpaQaDuy5bvyRsaY52YksF8BkzYI5xOvCIdk0zJtoT6EWkSfvQWzTEk18
iICxhXdFbyKlNTjtA/snMMg6iN5eLWqs8NUSMDrBqaM17ep+FX4lpjSoWt80G+A+
xnsWczfC9l1UQhsVJbBNyTC8XCSfgJMQin4trJy/+ZpsUWISb+OskLLJruIJ/S5Y
1XMy7j66idJbe2CTljjt/xKrTXk0LbJVuvzs/2yqHmGZcM56jZtTCrjA+YE6Y3/o
3AgWyMx2v5R4KthvjbYxWt66uEsCBsf5za6WXqDnIt5uZhx0rqC4YTQ4tiTVurgt
0+Ip9muIS/DQ9XMf7Fe6vd/nAcE5pd4EONSQtlyEVTcDHgzrIdFme6/bQfcMNCEX
EO4jLpvMDXQcxMtPMyXOfHBncgPBfNOgEJEDh88ol/XU59F+MLxhmz3vg0GIuuds
m7tFSb3TZHLxreZdYmHC4i61VUkrcMugQ24upD8Gs1dvWkp40kOTL8tKVKGqM/db
7p6XJie7k/OFR9I+JLQD0qqI2iU0yXbttGUVV6LtWudiprzWxkmi1l8wVE7y263X
UJHI6xXmzD4Sqf4/BE3+JDMCM4ZHoi/NsUTC+DHxZm2mvQDOnaWUT5pglzUcYxxK
Yf8C4hmJXt2vpOlbOKQnFCkHO6n87I9LhhDSS4G6Y8bnEZ+lRSHgGWtDHvjNr9Bm
FVATa1rkIvWG7qh++BtL40dvB2UW21T4JfnZlVCMBxrIL7Doxt0XXFHYHRkadU/Y
dsTNwp5hQ1f7rn4s7NsIIznjaafN67/IMZJJX7WJRNowOe6h5HrU11KA2/uW2Pby
ojwpU7hSKqrpq8YYUF4vobnE4DqRmgJNlkmk1q58ZUY5ejH7lzNX1hyhLguvxo/0
teQla+uaWkORnfH76IBCj4QDDT/rWpFy1DQLHqM94pLhqvQEE+7iZ5ha+DJ0adHZ
09zBG3XkPp2+FG1+rgWnBr9FQ3wWYb+TY6u6rDKunxruR7k7khwNGN/+oH+TxAS2
Wo71SOpG0WfAZqB1Jeet+cIqga/G/eu0r8v5exqjtJhSmsXXKFJqNg5uoU5nzQXT
hhzmbgnKg1bAlCy1VBKOu105hRw1ZjcgcGdHk/jDVhOK/LV/LrWUYV9ME8ESelaE
ZUieX1mDCoJ/gzYCSIeHM4oNmDmd4n1ocELC5pgUF9I+dj8AUqNDJvlDH4NQWRYt
bEXbUqw2m8PrSqvSDIIr79AEBVipCuyXaaHMGD0LJZU9YTk3LwTFomwnI9cw+XmB
nFf7CBL3jIhq2tHaGaEltBwLg859mdT2/IUrUqVnTyR/vdEmriFtbtCUHDLHWCNP
QBYbAyMOCGZVEC1/6XuNI9xN2MfXfykBFNAmgvoY+0Fh83OBfYL3xA4vEOHl6A1I
ip42eMCm2HU9QJKCrnRAwEggJP6/ScwTwXGWlkQII3iTaRs4qEuVj9Hxbiw95TGO
E/W3Wockkv76O4YRo8uZOQmNGaLDQF54HCnTjKy7C+zsRwype5c1Yd+gZa1CEALi
qPHJDfPYTOAfrpYe8tN/eUJCSU+ChciTMDvyDl/S7Hsjgxlr9bETEWRR7G43+1vH
C4G6Zuk/rYMK1km8LsetPV9jJd4Q306DBNTNaNoTbI8042wcBQS07+/fJuVMlpzM
AZINFyFnFtWmIhapOK/H8XJ0Oi0opBv23OsZMm1lU5ioQweWvIUjXDh65+kre9bC
debPPcvvkI78XAsjyct44u20VhAzTvmuMCYqJDHCKrBqYOlACJP6qSqv6ngr9C3N
G6R/hfWNO2XCoLqplNiD9oVfAUObF59JbqAP7kJzf9se7WfBxe7RCMxYhhfLuL0a
OXRWZTvpiC8X4q7Ev2ghZ1UNphYZUFF7aUcuNoBMPOTs+/mh9z0mj2IGR1tK3I8M
BCgUB0B7KMiouj19N2OkLdot77vzxtt6+ni33iZ46oRx45z3HvD90ILRicv2/b4d
iuzrYGbh2bBWR3we2SysiL+OeurWfpnMtLSF71K7uM52rcIoYo2qNaRhUX/XF5en
tTeb7SbwF5cUBQTMufDlorHEHk583VyHky/gkVV9H8KRPZbDAiY21lZmKNYAzFbw
p5c/m24lQ8IgPvlyWwBEEVp+B6WmBVbDfURu3AhZrwrBayrkb6EGAGDNIuariGle
KHnkpohGBwxzTfRbTlAK+vBbnQ7uL5heRq6So6A6bV9Y1LTgQaC4G2WK5Am2a9uc
8GvP03bsV7IajPyDC2ZSAOi1+lsa2S5XhrlZ8A92z1OgzWFkyMzUGzRc4L96b/mC
o++Eq+xe/LTLXnk4+9KGVs5VHLBROJJa5vz+rlquTo+UKVG9HWv5s9PBZQQGFB2V
OFDP+hEwBea3SKOC7tCEZwunpdN7D9fndvI/LV7cNqZbrwoJXCMCIj0+J/9LdyI/
bvCyieJVYwjOtY2DBw+6F//hbTdTLwtMcs/vWMWtnkJzTZNEVenMqFyY+q+FNhEm
BppnEOt7ZIjtsZRuHQCbsWoaZwa4iS3ztjGBT6lMQa3gklZLdScLQ2OkKtA7b2CO
lhnYQNzybhspFQXv9+fOQBMvRI5UNu/n6RcjKWFirS+dzmwJHFHb6PuHdpvD21yY
bi1jdQ7e2UwNWXQPUTxflXzMzMKlJwGgqMrBmq9/H12fVZkiI8HJRUzK7/DAePLc
r1GjCEDus0Q7j96siWobwvJancbF62jiIqjlQxnzfI32XaUpqb3itZ3XIkFwoJ2z
HB53q14ZAzl7/s06STYMZW2bFXdH1hOjsyJ1hfxnKavIhX5IudepXBI5DQtii/w3
zTfR5U+8ivPW9xTlLPrUFE8hPonVU/IOmMPCSshLEKAN6VFlrA/s8+0vlEr/TmOQ
6XQm0qdkTBmNJk9F8erng5JIN3JTIBCNNNB6K8w87t1U2qt8K5Dxz76NwKPBNqRq
9cj7yK1N9iHw6xt7//GANnpViiYOj2BCNLjG0nLCHM295WKwXZjFYi66OWYORvrM
mjziYTEVz4F90NSiZdb2pZY0bTSDuO34WuKubkVi8mVnBjBmUyBn32PqfM9+vdK8
LDITq6JW2xrb0L6z0jYyo27TL1wJjtLQ93KhrC5LCipI/e3P25Qg75E2w2jgJvhe
euOtNimKMenspPc1Tga2Rbr63QSuRB4hjgucdVZu5107BsHw8+Nj2pypQNd7K1wQ
hvG/ZQLLB7eD07UZbIxro196Rv7iWvsjXjYdF7rfd0x2VBFL9qIi+rU+CDZuEGOY
GvvqIsx9ASb6d5+7Sm+pnJFHDeThJv/B7vDb1aJW0WZCD88Ly5rnfHpoVNmL1VcV
13H/jf5MrL+Cl9URvTEAHXDM3lz6R6ATy7hsvalGKgDaQFehsYhZKLmMB5KW9RWm
HjpcCcNUvS+MIN/KhPb72AqT/be8eL45PWSeEnV14/CeNp9g8J/iP3uHMwVshhOp
HNclaXkRwBo7Oka70Eehokg9aAv1BTMetP9gMdzUd/qU4axW8cxQhWpMzbB6q617
5skxYP4btYiyhZHbUVzpWUlPXWyWrKfIdYb/dFni+osqjceYk2Unp428UhMX/wAq
AS3SHMXYeFm/EGAQi3kmBH2VS652JgshY3iMguy1bvmWRFWVlwhQntfSSCyUgnHY
3XL7ihdXczdN5SWzOGJZOru967S+S33W4TbTq3riwDVcBjouRf9hzpm2lB0Y6zSV
0e4gvWXOUSqnrSmtUccj2vWfYQSUBWYgeLRRJNcwT49f1mDCYJo4CT3XknvgD7UW
afqX83jRTxMk7ZYncCBErNVj7LDO5NKJKPqtIxXPFf+ZrcIkpb7SrQJ/ekpaxsQ8
9JlPmxyHmmaaPqcaOaTpbv2Cf3dvr2phiDF4uGC7CegIuxC7lHf/as0UIvYKyG0J
8HZnqX1sYxhlDQxdlBlPfUQWdtgrqEGkGo2Y64/vvmgO1HfHa/Se3TvJaoB+HvQf
P0HLZnK4nyQNhcPhs6I+8KmkBLQ1EKZAOJNQ9nIOmp9Tot1Eg3nB1fQhPEL+YX5X
vf2Gu+6YCnAh1tnnVcWfCr6LHobjp6LnVREDvbq89XDB7JVW+J+5TibiZw2fMGbQ
KiQOijEKy4Ky3Y5g7diRwZuzR5tzB+BgMJiJmh72T1Ept8FXyBWlMc3gFW8QhDj+
uSqY/Kz37oXpWAYENFLrh/MNS8l3BelqSt95Y0drE7MOYy2fVBTXwWY7gqLOE9Ez
MTQae2Y/3oRQoNjdsoBMlcrraROmJsjKqZRP8DDw6azSET9eZjoWy9EXsrUY78d5
kEn0R6WsQw5PQInjasaBxRalbTQigrRVI10Qz+wUOTP16ACPjuKfqtfPrCL/YVOr
PLD6QScW1TVf5OdQ+qlwHBr/oo4N4wy42Ulubxf0eXvl/CFV/TJnoht4AK8aDOyy
+wnjZwGu+xAc+55xNIs14OjkFPEBHGm+DsPOjwfEvkHC8p5AKcnml9JPnkjPPHnz
4I2kSFFhqG42hjyE9VCqb+meO2GDOf6lHTrP/vsT/VerZjjYTm0VUecSAK+vKW5Q
40QRuFsO20WvruHuL9+YkQ3GV9vC7UJgS9PZjlT+8j6wYJmv0bUI3zyiDd/2lTJX
ZhanB/HN8pBCDOrb71HDOR3IEWgr3NANiilk8mAaCDBlPS+9EFaAy6AxWaOAA99f
QBwj7DTFY20/oTM7saT9UfNAgzaZOAHVo/T5YEhisJ4tubQwelpBCvwemxS3EuQ9
zY6Gy9WG9Q4XVeMdFzZYtPwawUXbseN/QqJWtnG4Sf+LpB5At8Qx4yFMpm3ovSlk
MTNL5pQ9GRfoUvg1ixz0dGKkNxiAZ6Vbp/9equUBehpc2iZ81fZ+vK14ix7sii0W
3R3oFYZdwI9LziuHiuBX1AAkvB2kazIpBONByYkGzROwHigHnkLVJck2Jck6brqg
AXSsVmymRKEcvkpKISEiDyQJ16k905q6q5090LfMrRZgq3nHO9TcKmoWT+QgAvGd
u+e1v0QkoHjYpvazuBCMFfhoW9YPEN89OeixKw4EjethOZuG0vHFW5ozRKY1lxaP
OQFQyRtSSJFyZ8VpgMDuW2sUMAS2/7rBabrGHN8b+iQ6gCobm6MFrcn+gFcNEbca
hbRXlzkJmrVNwPkwvJMWfyLECD4gOVYXxCIRJog6qbI2+3+T09P/Vuy9wInSHfoC
G7FPxsAEodXkV8+v9i/kyhgnjxhV6bX+X/iaDbx5FiV2YAhydTs4bxJQX9o5+m+Y
hR6ARuUFCfwnVKi385xWuhki0+HNI6h3UP5BRKB5p71cRWUMmJvIMiRgBv2Tnmq6
RcXWXnDaFFl2fxc38YtenX15wQ+uIvX73SH4rERc1nfvltMWCefnyoCHAKnbFDMj
3DoieyupX6xjn8lPL13Uo3TWaWi73veiRHlW2MXNnJPlhOZ39BxtKqQdpHyzgu6H
7Gik4b1I9fpaaXx8prssYi5G2NhcRl2cnIPcnXLO0ZEHwX/f7/JGd/iUvx12VoD8
qSe2Sj/FtV4evjLmO4yGhVsSLiV6Lj47cTtfd8e5jPaDSNLksiy0vAtPTR90K4J0
XTjNZruR2I3qyETHxxTlHvbQikkaLmvFZPF4Pr3WhyOjQFEsp6TX+OOp96cqUF8Z
WfW4bb83kJ8PN+RR580ZIxURNMuaDdptdkMvM07jGY6fgq8Tvz+JWXO4OYQXQ8py
b2xZ6oJ8y8xFa3DG7t3+bFpfM+NqUgLlblZ9gz3tZufmSfslGMbbHOgarNiX0UCu
/9dGgVfl+7JK8WPyqs9KNZVVQXR9q1qQ9llDZ/4E8FCH2ITv3rUTKEMzGaXat3uV
z07Bl0/as2uF5iP1/BHYcsaG/YxrQ0hNsxGpPpDJonFBq7cN4od3yvGLsFIGAt2I
O6xKoAvEcp1s0e+H6PEgYKx0duxhpRpYap+bBdJVHVZzXFXZgcOF0OcT3ckkfVcU
Vo6evU8yKwJ9pWXlqos6hHWZpjlwAtIRpBFeLSBOjv0YwVI8BEcDrnrG1Dg9xRu8
1bBHlAylALvBfOAN3ciglyjzQWFBu7lPccsEc6iWqePr8lA56+UhpUpOal8V+eF1
Y2/YmxHJbuJRkw7X1xhqzHEVXZ/W2Q1rQyy2fUesVRfxLrJ/Uc32we76CYYYo90h
dQ0bxZetKXFfoVX7Un1EwChhfavwY+7VqgPU7Z7Zil0Iu18Qng9klxggsPxuYu7F
HNeWokiOfhvllezDNvPVZNjNQDal+q/DRZ5sYPEJPDeluFAKAnJ/BXF0KJ411mHh
ukMA9riIORuJix5A8x86RlNTpyZf5L0VjUe5AWymZQ7uYQmr/BDXeLmS+JpwtTca
rX15K1pYi7gj8dFeX6eOvyrqy+P/z1740urRBIhhAZa7XUYJB2gTGOQcSOdrN5tQ
VZhjVxjKM8vKfBxYqm6ZCfVBhnuZaiDJwiZUPUPMl1OG1Q+qbCLBGrttw2iWJccd
sB1m+E9JGTCrF/nFMXyi7BVwaF+3Tf/OGSe0O08RYeZOdjyNJfKyLnQBpyoxPoA9
Me3ovWSF6Ol/At20VOqqlo34Fer2zZhse6MxsJK2wo798hOmd/uzE9PJ4WexdmAA
3biJKXCXabTzpo5k2bhXN79iZKWLDUTnVAbjQft+R0zpR3HaCgqHuaOuNnjn0g+b
NS2AyeK9epnMFj45u8OKdn4P8mykXL3mnF1YIg3zySGxf4pruR4s9+6yLFljBGoS
TjthYDeoEtXchzqw+tIRLcNhjjoQ2Un8G1ryUO6+rOIqxRmT/K5Od5YhuIiKYfP0
KvnjLZ7GIrYIT0xuu7k+BiBGnzWxOIG9xu69fj5BYPQ7zvNRrzjw4AILzfKMDBMc
HQPl3+hvKHc1sGYFflPxqbEDxcJZSUtlGn7WQm6hRNWEtNNWeg9qv961EkjTRgfv
wA7UxW3WwB/LKHZhwJ25PTPTFD3wmU+FkB7M1co5zSO0w1sBUu2++wU2tFPI6kOp
7LaIvX/oLJthjVWv3pmndawNtaqq6Po+rhAk5q9I0Ju9wsMEOYXT8JiSp55kG/hg
mL7/ydIe4IKcExKt9ssmPqwD4yFrtxwqcF+yjiY5w3fn/i3o2bDohdmZ8t8Ssudt
TsAivbhbWd62iWUWjIUXJmLSbOqjMey5JMckaeRzEhCixB55a+m7GU436TB/6JH4
Bd66klq4DNmPTKRk8vs69fo4Qn/Qu+9fDwVMsvXYB2Q1fPcsslIfRDWaCxWreSxe
2YrPXtrt0YdYXKYKFciH5/CYqOOfcfibo4S2786QqniOqFPNo9G11OWr7Y2tZ/W8
mBo7RN5+KQMTM0TVEDpxCuZGUKJsbaXpD8aw02pS2cqYsUa8RJpFUtMASYhreMur
sy9FXPxapz+ezl0dUYLBabE/eFLHGKJuFH65LwxnM+kOI1oeJ8emeJgne9m/vKge
1qXTXZFmq5JKLoSM2iXn4ZVp+LUfV5rc9tprPoxH85Ch8OF+nc6ODgc4Qk/b+wbV
pqWgMO3pu/REgSO1ajVu2ewzi5wNN+YH9TMnnOhDVds0msaxZB/lDuuDGVvtHfYJ
nKPeDteWo7vYZI6M//rI0FWwKBJzUuVrxs/khI+1JGgHnCStnuQMAr6jIPOyxeG6
R367OnFnwR1ZQrH7o/Tx/7fLfB3JPg2za0fcwRlB0XhUEdsidU3fTLNjyJxS9IsX
fv8/phBW377yOl2fA2Hql1UTqEvoVTjCbSPf47XcRUMfFItVFo+DvC4pbg66IK+a
cWv3nPlXtMD/qjiTLfFap34wlM3sXNGZeuWK+DneRAhiUVhhU6kl5xhveUI7Rj/Q
HCQru2hkISSFNs9d7h599+cFovcWRGhRFhCFM2cyJHd/mXEiQrixTshUbY0/nvI+
LdyyfWC+MoxJX5C/FxC7hAMOCNISw8i1pkxlBQdhcUqGhNdEQkhNEWi7ee7bE7ga
nvHqpnWJksljC5DLYhmOW8ZNJfDMB/ZwVse3C67eX1NdN7QQOTXIwLXs1trFXc5d
MlHeVBON2Tz7ykm7tULTpuJgQshZtawmaXiYoOsWty3TP7Xjf+9X1kSQryPTh7as
V1n8hWF4gPtwxbEf4SnhNiujdFI8293LDvGO2mlW2zM3j/ym8VDiQ9dLqOj2A26w
Q4nkeUQFHkorVoVB48PFFnFRnDD97h2DAoa6RJlnzvrKqVsiS23Xe8qFCC49g0S2
nh8Lu00BorbqG5sh150YAWEb2C/ShiM9kRlJAVhcKPGmeUPDPa/YNzYpxGzm8+7Z
IOR6vf0XrT5XPLzJA+dlLB3WEyFAza+8/QmS3kDDuUlf6ZEQYDdJC3pWfMicSwPs
hkV6bGe+Dd5EfLP2GlGBh2CdmZluum7tnin+8PXO7q64hMPcgCuxlX6BGeQFmn8i
ZFohdG5qZ8KAREczKIQoKI3M9JrNN8tKlNhmNfNsJSpr1SmXEG/5FAAEli1ado63
7cc8TvkPLgQU8xGsQ2hUUc51StHX1XXMiF9rZElB2USLyFcp9CMRGSd0vTgZsKmq
AU1ekclgI8xcoiVhQmBEry9ytwbWS1lAoXikZTw3ihDAUwbTdBN0TGVIaQct0WKR
osvkGehi50xrpdcnLFrIxKtUovZfwR/cuaWMXWmET4xGaI2r06UbSj2RmEClyO9B
EvZS83cR2mlweVIny2hOB4NAmw3zvST7t/oCqOuqEetHd2sHQRcJzvoivLKqAF2C
s8hRlJjH5VZIzi9v4k5eF3bfCkDiaCaE2uA3rv2xHRVjaIRXjhIo0MSaf41hPDSJ
qm4p/c8UC0+SP5P7wwGq44Kj/5qGonvHLWxeOxpcFnTrZE1k+QboLF4f2ThpArcX
4ak39a1BNiw0lI+Rehs3INZ9wdRgmwKTna4ICW7KAnTc9ABasvzIP98TNFzD8ZEW
QnNENCdiOVxVRftSwfOZA63eZX+hHgI1Ehe5/7gLmWZQmbFFmXLfLYm3rXt0yzFp
En3J9Z+wf1QKrMIu2ylMBJfmpEY5rcEH1yA9PN5W9Yt4ovd4H6AMziOkdVQrN3r9
xdidpedyCCSuTJwi9hSb1VDNfZgFG8K5jMzSVu1upNu+s2qROMx97ZORXhW2BWIz
zNnqbmXNjDGcae+a1teY3nKBDQ/mOJIBgT3W6TQwUf4qfEFtOAcAr0iSJb5jXgst
ObhKlJfqu8HMAs3/hzBcydVYweiBUfM2+hqJz16wA8VkSBcCePVsrgR021/OrxZt
1QDTKHcy+33NgyZMde6PuWZ8lcXfi5/1DBLBoKn/Se8rUlb0Cm0413gQSOIwoAfB
p+rkp9pSiNk4LaB6XsYlNn36PnrQcW8DPTP9mlEIxct0Qvp9uEdfpH7Pwhojb4eR
oW7VM/FOUFVs1deJowoD2E5jy68A+3qoRX5URuXCjU3x/d0yLKmsFSyW/WxQbjxJ
/xl2lM/JQBpl6rz+Tm6Pp4pjvjpo1YvVwHckJXRnjfEvEV9Mq7LkL5A+ndf2vvxl
/7sISieTPPPL6oZYv5xh9h+f/uj8UHKGNsXEntmKYgDlOc/nLITPLDYSk1wx/FX2
33keDMhw5zTsjhTdTzr8lAE1L8UJm4jSJC5KSz56NPqGDzaRbV1h48K0xlolX02U
ZZNG5SJjHXwwim7ifnHcUhH78fIMoPvuTfQ4v4Rsc3zOiGWGDa4p00e7pDT+PKFc
nxxdzgBje879njOlOdW+YCcYisQuJRzbEACUX6lodGLu3+8xfCLZA8TkHMNvAqRz
jkhHSbU18eGl2MJ46eLzEe/zTvvYlanlERFzVhAysLchI/O+aZEFzjpZzh6641xO
VP7S0aNwh6ThmXpuz075qF45caDReczWGxdYegioB7xQX5W7dk/6mTOFPGoqHknt
Uc5870kG11ueNRgz1bOt9PMuWv6DsAjsEx/Rk6r62AIfEOGLvJIJwguJfDUcYVv9
5OsYaTb2dX7Zl9GAl2PyysJtmOiPBeYYy4nZVfcSUSokIQkAlHFQmlaDqW+joEUJ
FgUzHw+Jqn/KzQ96TAZTByMxxs15k//zQRCe7ka+LPM/FYWm5r3fdDIJFbsqioYl
AAmyhJiXcqkTuCiupYmr3ZcWaGT1pXRLjNUXiHNS2qKG7roNW2TgOd4RAa1iCagZ
zcdFScLFFKgcCzGrsCLCN4YVP30tlzS5WAP7CFB32MW3wyNj2M0vYba0kuWsKEpp
nDgLWVLTHgOHraUNpo3N1QY6cbSWRW+kyqtOwJZFJaixk7atJP0zJIyi3yNEOWfJ
x0iOUR+r5uk5KyqIte6BZeXz8JTnYoxeHgWiAt0S7Ti+4CD3AnvRbEpLdTTqDeWb
GWUhXUpDAsQpdwBwmrWCN2VydJk6NvZsc9wqfUQDqGRnAH30Na3JYY13T6WxOu38
hrXwVLrzOfPdfHbLAoMTiN2YUSi9u4NvT2ejPmZBosmjWMVujLkBFD9/C9Iu6uTY
0R2di6hF59BKb03NnDSGjXI38zv2j3LQaVjxkx5SjiBF5kwqvSJ6EXx2zyNGewRU
gki5tQPUGMUBiFRqYloH5S/3O4NMUk97fRMzXC4aMT/+XzFOPY1/rNbvrUltFx+d
vdu8feeO+gZbYK+ylaObc/YAZOMmTLIlM56rOBgiPvacAidIlkgeEUuTtFPCQaxn
elNUjkuvi3iBaJ0SEVb5EGdFraX14BBvWwjZUFH2bnTXs9kw/lfwPihqv6b+VPo6
cBc5o8g6BfDdVTsnr3QekxivIM13q3kClhtPcYvJHVeGHkmGslNGQ16FckuGJn+d
IPj6o5Za7VunD3EzoUc7yOSpoKJcweaKGT3iYRXEjLHIaBzqgR9bspdlNp3jGoEb
BUdR4II12x0+e9P/VE+oNYt6PZKPyObuTD+rlBG3etYd1L4cMmTIKXDplg+7ZqYu
a7Hh/lLVegOjbQmS8EIbLWMoYKkiYrn65aPvuo2BrpJZTYLfbEwp9dbnXISlrQ+z
CdRn7CyTRVq5e7slcPJJ5b3vs9klCJ4et8RnHh1ZFmybf23nWmFQZtJVtDaPUWMe
b3mnio6+oUTVDIHrJQjJ798sByFT1uj+PAayQzoOoOp2jwaZBtUiSoZSp1lWEhdT
WAZfpC+IswS6rLxfr1ebCKFKUlEvCfSEUXnQiHGiGwBh0RnpS6XpCmhkj0NFB/6n
H16OU2d+Ra+TxTF9uEzlgRmlAvMYgsh/qi7ibtg+fewWXxwZGYZztIpZF66XVlAS
W7khcltHHDye4EQp9etq9KPg2w4cgFsVdoYyJH24Cl3upVdL/JPHT+RdlKaHxE1w
zlhD87kYS/s5o2Dn0qMd5pa3kelCR/KoFP+AZew7ao07qCCEHudlGyCEjILylOO6
hmOxW5TRBSxdOi7IgJqLS1+vgBuyT6SPX0pRrHvS3IHlpRBDXr25+y2SmM1+/Eax
AAmHeVfZRqOV20hZf8qFK8dTuVtMR31hw8H9GxN9MPjupzn6TM9u/6z7sAAppf46
pmUd+3Za3ZxuNKpT9laEYE558KbsAKVTodxGwJZR2jw78Qklh+wgt6L9mbraa/xv
ok5UbNsUGGl4rzrb5Da05ltZJS+2I64wUwmGi7tVpnzgoZOrBiaALnXGKakTK790
7Ke85Zkev1E4C4WHYRipuhiq4OKK4iy1YhF4jsdk3l3i9nh5u8ZBqumm6JVtczer
ZP8ejBeTi/jnp4ntx+AhQ+H43xKxso3j1DrP2uQPAvCEEfyEuXva7IoWvP2TLhcb
eSLrCvUCdJa41L0RveVZMqhwqsPafDHqyKXIF8xAgSwTE0jpKEPEjkBH51+y3UVg
IMFy9PM52pQZsKHoJWWCl5CY+Seib/QAyoRG1jUTRlxVsWYC15J9QvvSkEjlFb9A
pVdSQEdyGIjhIqsT4HF216S5Y0fu229j/WcSUAE7d7PkcfSDLXpUdT1gWr9xUD2D
uogF2PXdb0jKo5SevEaCpQTJyPXDolgQ73mijy0k+fmrC9CgIo8DL/gfTbecJu27
TX1GUJHDPfS0rawzWxxU5WJIJeXRg1I4KFpN7Y6qgQu5Hh8VgIK7z+UG496pqv/q
Hy+EEd+4MXh3MovzoGtJjTfYlIWXBWItpLvbJO0SthAIO+hYtJWVsSAeW5yHpeV7
19vrfjCXdGie3iUajWj27AKkqsb65freHEirSwhMK27MQrI/+KjrZD4tsPdWIFKU
JWUcf6DR9FrzpddLNH9z9DJXlRwrL+4hKkuggXQwu5kaH/xjOTrhmEm0LfpZ4L0Y
QfISjG+B5zT34AUkbKpG070DnusH6SDMQPRsZSC6aaQSFPyLv2JYualw2ezDfDvx
IlR5mLrC+44NliOGghZRS3fyd1994Suc7oK7fuYrUbHbEI1n/s9oJfQaHHpuBm2R
iRVBoxbUQJQwKvTSI8AJcstf/Tm7GhqE7q5Ps9E4AmbwjoU52ZVuoZsJmXSrYwR2
HtiUkvATaBHtXYv+v5g2Evqut5RYIIXajjWzUlL6j9PvQ7UNsu/+1sxBOGgNWBGF
AHlB2D8kKtafz4ZQYdAC4crvBlabldqB4ZzCZB5Qhl7IMNxr9wPoWfoEf8jWphOq
mOvowl08D7325dOIosUxIn9NpPxK8CYq0ZNmqxjblcSjmBeLSXh3g4ehmzOyU23k
IUhgNxXGOXYN+rHzzUwStO68Q2INCCZOYOY3K9TBdcJ6kS3ihdNXhsDFVeUbwlkb
vzRRO1NLkxprmxmW/E7mJ+5HjQnZ2qeWLCLDhtqXknYMXPHv97TDZnEbGgjUH/kZ
nrJ8dEgZBOfyLoswhIqBRl26ee84Z1PnBVXn+tWhaEGhmCvt2gAYDi38t7tO9c6g
1rxV1ITHvee0CccHqLJ1ptoZ8kQQ9is9X+LKHx2tRlhTfSyVKh56fiWNfdXLL3v0
Tp3DYQKXNU5qvgDAmvTpDoP4OCSAga5QRW7yf4s/WPYyw4UJ4w1qGej4HeRQx7G8
CW0tas4jBFnnmvuzC6OLWvaZZM4Df5QONYD3KlNiMayahs2elC0Dzt8VqN5KP5IL
ZF7tct8A0bnzlZuUL06i82giPGHw6QL59D3W8aTCy2OIOqwJNojhfiTJSmYHETZL
ugQaN7uzdmGQkhhSmLNFS9YUgd1zh03NJMxVmzGuqzuiWKqj4YbtKnM4MUc2Avl2
KOFNf2ECwHgrB5SCdbIh90+YnZxnfFgdRxZAenodtOeDkSU52Hr6rtmLjHxqc+1x
TLWxdz8iV6n6nASHBs2TICnugy0bI+X5AL/kIprQvB5TaAYq4IN3vuQ4ypS+U0xL
KGj9/+IHeB6lxCVQriD5B7bmKi9oC20zd+hv7RBMeHIFqbdHVjeXtuT66R2qHaXu
RKpid4MbBirUcA+Ika3uQN07usGjm2gf91fu2FEmaOyUcG5ZNoSOasXyjFFR29zV
xcNFUPzDCVMYeEAmPADtzMJp05PBJCfTySWV1ldLvOO7peg0jLA9NJJ9e5kT1SYk
Nhzl8hdWcYMHRJfxRsD4YvCGOEor8Hk90OjJiYzHpjZzE3Q4+gvYNEKBNEIHOwOp
oDuj2IdZnanthUjz3DFMu2yC07PBfLiWOU7iHC5LukS3zqk/K5PzCCoNjKPgQ5Mh
NM0VJO6tW9xKjd4WHs1v/QqHMZEn1QT4J3zoXGh+PDZjLQIReqG+sNu+sWXyL/6f
X/5mIY2PX3kcSwKZ9M2Tj27KxpWGJmAG6Vp7qBRNKxI56HmC5XCTEjNJ3oEF8TmL
Rw1dj8PxtfhI4DHIK1pe/AYtsGcihgtSAjNJCq+VrJB32Y7tUCDHH+dVCBB9Fim0
pLqpO8zDwp3YgpI5CQ0Vq34giVytXRNjXCMs5HWO5qow3s4rwAYVhPHAgOxy9myT
PoK9lAU9Rxnx94XMuEcrPgDUMk5Les2Mo+mPbhKZOHt6NfJ9gFe2isRLh4bIS7Rj
EBUvBSi5ryXFS2hdK97itO+pfdvJ5pG2QF06buSaGGop6FZW51RddmzhbyGTS6ms
KjOdCdXwmkaS28vRLkB6Ni7ZDnzNrzQhOe1cCfr6M/BZTcacNc3kHQCPOXSPA9MU
085J9v6G8tYXMmbRI6vSZzId8ofv1tDvsRRRGjmmW7gZ+T8TVOfwUxt423zejXOf
0Fp7YzK0OCVtiK8tB44/qzggOUryllo7iWqN8MfYsxqDpVuVyu3o/zP9cSz7XmXZ
+dNTLYiRw0hvuf/PQMmL5ZjgAIwKsM8r7HvuYr7ztmTWbxKNul4IwDI7MwGRrq1T
fgUHlw5696PZLYdFQ9qfXNE3l3w50IclGem5vGZt2p64HTeE10nzUJUY65708FAD
UssL4VUZVlECkDaiy7fv9OnGs1koFk5jxtzA2RflvAjZTUmKHBbu9ctDGA2MOTml
2Dmau4HGQGvL9bFEmI8nqCe/ihO7OEbM4T09cqAGd2iO1dwXchzMO9Dh8PTAQ5MX
JYOmz9SbRdDI6HkiAAzlxqyfy90iNa6nY6Hj9NZL5orxeaO04x4Ag+VCBk7XFWcZ
9uH2jQ1o0Jhvt53H95qY5HfnbPc45Ie7NDeMF+JDRoixZVa/BPXp2QXFIlmDluQz
QTxsegryjoSJyIpEmgPQNyvof817Nep5QHBCU4gpxEL8RHime/J8Vk+4UhUAzyvt
IzNoJtaeOGYYB+It/eIP0nAxP0hTrnWJ7k/NpdBPRziw6vyTE6Sdl/1rdY5J8puv
ztL6l8jsn/k35xt09IzKN5fN08eha1jEwfn7T0q+EF7QgjuSYTKBDUQtMKjkyho0
9hjcL4kCcYtZHF2Dpi/XPyky1pPRdWhl5do6MQQYys+qghyjUUB64UDDROBfgnSq
pL172cN9SqL+8aY3UkyNkzuSCZtJcREjzj792tMkyrpFnQ58ORRwWRqkbWMF2W9w
9PawTG4LWUqgo0B7gzjOUmGeYOQJVMB5XGG2NWUlp0S3zcyVMTRQ0PnVqbHB60zM
kY+bUvEHLAXqk3szDNOLq8Dl1GQQcr3xHO801CVuoPk7NimfRTxZ2lwOP4B8v428
bMOeBZC8nHeCyw6eEQ3TqhpS7qSMZmqYXKQiiPF9Jlqg4Z9WjMyEOqXvA/S26/1p
rlBs+ItXXnoK9uH6CwOe2VX/3GGsTGouVcvv/KY26URdp0OlQhFQ3Kh8yQUxkgY5
eYgoy0PO+RAdUKbmPnkbFi675/HM35bnVq/gsBInpNznAoMpF9j7Ew2+lXbRJ5fD
pHiRcHXSVvnJmsr9y944siHmrMFVb5Dr6Ply5nkXPyZ2YoTP33t5kf/selcahErJ
nxy+egrfbwPiejMC8Ms1kgCQS1HaqE20ed3CMcfcvsom9xVd03LoAhEIpS1bqwu/
wQ/PMceM/pOw/2rVxdBk8n0rTCq8iS82uWQle4x02fPjqwk5s5zSCGRlswh6NZk8
+npBFvNbaUfUxiScRc4qXJy8yP6CN0lpvFHKP2WU/9z7sgonj1EQIWkoYf6vK1bJ
JcDnUURiFkwF30SAB2arw7IdCVHYQOfwyk0xwHREVHfkVm1YWsdeN3cQAq376MQ5
Y4GzNiwCRMVMbx82wY347HapweeGi9gpsmlbhKgYsdzAKc8q2MMqZm8QaD4phCze
krzcOtxzZ1pvrF1ZQSjkZuQtGWqvLuCz9XuKcmEpc7mg26l0UqoPfj+BBOxUQjhA
8xePotoeqoZC+JDZsC2y9LJJe8Osz95cFnKP4ZP2hTagTrDJKaiaxqL+4ibu0EnW
Qr3o+Bq0dJHTou7TOblZ36fILYM2BK6PiVsWCsXRcP/FmuoNoteNYLQcGfMVHQ/9
C/A+YsmsbkGdjhNjCcY+jCD0ipHsYCSgSRwIg7+3n1gXD1n8/P2Xl/Mo2OQ5WS58
aVDokekOiH6wKZFrePXUMRxaFlEytp+xdk0gXqGQqeIGyo4ywKxZNca07uCHLK+b
c/YerHWLXQN0tc3ilz7bYFPckoEiUINhr0eUBffHS9Gn0wZsaVVIcRhwuCC2pA+9
ZIUCoooDt2Yq+Ht0OP0GIkW6ju1Xg6c2F9SBfISpWqIsHpOQHESVkwGTlCbW/GIv
fNDPBhLfBPwkZHo/YX1q/T++E9lsOAE/JjdZOTFlmq4cFr0m9p/2cmKTPiOmJfBB
sMSKc5rSbTyULXKHU8zxV31Bv5IoI1J4lsbXf2dNH/YI5ow3aRbu+dBHjFV/e7Cf
gMhDbGJCtgrkE1+fZW+rIZs/Ft5j4h3Cdho9Mg35qr1pA1ADgYDX6ONHoMZsxMcF
l6yQXSXHoVY8uO5aMEtq/mBE3unDalv6SfQft1H1ppd7moXrVxHe5bPSXt+2tQZ1
afXEHsWHnUa7T48unHd7LWZhI01AHap2nfWXtYbjpDWMAHekZyhH6bJqe0U1Eq8F
fZ0juTTV0wsWrkcrARyy6b4hf6wVPOnXldcD37muPVHsHdfh2QltGr/k5L9txbZZ
1IemHtnhcNzsvcQrfq3oirnWchPAqe0j5M04V8XapZuq1FxMAQE5gp7RzoUEx4XM
XrzxQ6joyXTlTYrcpTe7UQSXWqDhPAbwcAq4bHjCqxoQ0fNwMmLKOvhcledGZqvx
9ZSTOg3Nq1G5KqeTt7dpevEtGYEt++WXLjvgfLMGzvL9PHds9Y/gecO7D4nyEyFX
vgqhriQcQg3yP62cX83o6VxQOsCcb1HnS0R1CHgnoNc95Z1GMo6D4w/EODwssrHH
ItU2wV2nz3vAom9itZprChOkWZ/4agJ+1I6eKY6yTSK8SVemlfvS/4eNjYbUcbkm
z+Ipw32/WqsNbS1kWlE2j64hlFrFrohJtl5AFQSo+sfLBjcmgsDFp+gq3lNaqznI
uVhL6sY2P5DM6/w8ggQXMO8fO0uk9UvEKeC8eQM54CiLI8LbLJZ7ZwqKbE+9krW8
R4EzEG/VNRXtJ66hrDye1ASooiJEazKVDCcmXymzZcrGtJ9jyY1y0LgiNAN80hXQ
qMHbCBgq+yfZFymGBQk45+S5VbtnI7yh0TOvdkMZDwNt4dW4tTfhGu59+M9vHO2i
moTN+Xyt9gX00gLlzrQlKtW0nlX1gS0WZZbhdJeeyVKWFvX14ClSt3n6da3K0QkO
DWeHxd2KI5gFEEPNhWWl9VgwfkVlGN7CMdlLow4xQLK5S7BEqREJwgyFQfg1bIIW
CuDW4g7tB2Sdq4x7q+W9YHOmwuXANCc1xqiG+7X7HS/ea7nzS1TTMMfdggBB/xhh
VrIGAPvCz4Fz51Bm8MhbPDVcIXB1VwsXLv+apXkfehN4v5jSKivG/m9026suyGqu
TIyknkCuaDt4qduPJuLHd9HJ81jZqWKZdHMqFTiahKLHAV4XkTUAoLfHw1EP85fo
Fnmv+H2f0v12MxhOeAG93nGN0PF+lm4+wwCVhlZIZu5ZJtwTaEuQv7VHoMVRVHHi
WZBX1s9IcyUEa5fjn5m/oOsvRZIh2CZ+lEvaI7DfjPsRzCzmClvfb0ebxFrCiGX0
4yyWydnfRwBPZYXgWwAehrbFqmY5dRU6Tnz46hpxKzNKZ4H+YSjOjkM5BRNci8l4
C1ZkmwUyDRoRcdU6X7Aji7YwIIx9+furFDfakINW8S5wsv30ObKSsRh5NDeDenWq
5Lj1Wm9VYbMDRfyjCkDxpQtCVelaEgF2XU6zBbW69dd1SGe85/AA9bh14n6YIm+C
YInWPFGnAISLSsm72/63OI8Zt94GL7SR353wOK1tetWH2ZrLo8/3TQzMnpl6V/7j
vHMXKVcCNtp96/VAFmOhxl4wJ0KuPwDlg8+d3hTNSw4x2pkJePMn6A3RbMM7aHf2
0ji/Oqzkx48EyRHdiRKSP735ejUarDznsgYIZiYkyRNayW+P8mZntALXzeP32cGk
WNyLr/wQOTbf1BQzr/BCBUsRoxA4G1CN7Ed1kVt9hiVBIl88flkThMq4L2bU1wZi
dajQx4VAHKeYY+dqWe3PZLbnHBDvlw93HZJj7ye6kQUxJekcDRDzdph8Gtdjk5EH
lFeaohqSD7ZhIsWDq+F1s8LQeB8pB6BRlYa/MkgqOJavNvU/Da4UkhE2K+bCYw93
ilHrfMTQokdQySuL0swvM+wcZfF0bQkTeuM9DAr1871gNAvzASh8+1ej4YuxXgfJ
ptih34rfXzTrL1PXWbsRR3nlYrmLrFlKqNGjHFqu0ppVmSfutNGNWKk0PqWBMGPv
RR9CNs8J3DVHECKe4I8YlIml4lZgnfW3HpD08+IdNsrE4Zs6MeSrGctM0PsDt4/e
qxH5ysbEvlBO5QDrohFTyKNnoiu0YVo5h9jLLteXL7tavst4/alU88nwQ2kTC7ER
9Gq24Elvnjzhp0a9xdr4c7pJYV2Io3G8t4HjFUpmPUBFDsjggaOsKD5Hb9Vy/ZnF
S2xxBUbwx+/r2xinCLT12Tx0flcCTMX1pdnYQ9aQloIS0sFDJsLrT+dBlnHTOh/I
tNpVzXulsW21SBR3qUdhwIGytbTx1N9WFTRdUlI/SwrP1SSaZxg+0hh5oFG3VXmo
ut/5ocGz5cHXkqW4e2u3SLzYerzJTvDJPZ8WsEtfnWvERIWbPsgDeZefo8wSWsCN
wiwjxueMso2Ovhwu7D9aTblz/v9ahzJ6Hsx4SX8tGELaK21zKeKTm7vZd5penGwd
s0o1uFPAxo1CmvIk6rGNHiE9DWiC24UewXPl3/61HokDd1daO6r0C89r/PJJ9PE1
8AMLqUK6lJpVgVAas5SQvumERV9hYc/RjuVcGrCPkUx7uVZVOiKd+WsMlSym0yZo
tEiwzGW7IBSRtqy/9WQaqa0cOvOROhaKejjsHNwDIAiIRr/mXRiLwDml1lslVRY1
yvMLgxG2sJUwixHx0JYXFkZ0P56dtR2uA5uwp75e2OPnsKo00T3OOQaxqD51z0MQ
EDGBX6Vl3ocWj8ichiEamnePa00840EwKrs5/1O39+RiIAJR8/4K5gdP1vU6pDaA
zllQhQ/NlICSSy/qyjEhUkJX62eekeYc/FGToSssTiBFTewsXlPDWdQ9issOrUl6
KBGO+/Oibt8yHKdYBv7CmphNYqfT2OY29MrW5l9bXjnWrRGYeMOmZra5YhJOTGii
9PT7C7TY5MsaJQiDrmooAHDZnSWL25w2l0cA6arRYk0AXoDKgU9GgfAnyOocYGNI
uF+2rPcOfaLC0zV9kC/ZT+Td2sZvGdx/PqPFn/+YEvmCKK0rXX6hNhAUImi/sypM
gLcmHTpDrtrB+gtZUD2Vlr+4sVPBkm28l5CjJe9KDaKBh0+kGJs086ITgrUC5Edn
VKFC9opESRsmHq+5jNcmJz8NxtolLInmNLFI044CgmAao+TC8BfE2zvEpCCMRoQL
KnFbKZaB+HsanCFIBgL6SV+oQAKoW0zadIeD2BNvmlfbNi+D+WIQGt1VKjMtpBqA
ngkJUfMsWA423isfB1zZZW4Ck9DOySd8zmMXgBGbDbD8bfCrd0JkcBQ1SsrlHQLy
+D6QtDU4N7gBkNebzbkheyoS2iUk304clw+CiRZvjURaW6PDdK+fDMoPbaJ8oFja
sh4tLmTWVUi7PtjrIqBkVnQHdooKQnDgVtoAjEyhpU5KJ+m3mPQxIzVOcVw0JaE+
VnNzTEXSfWFP52JvjvIipW5xFX146k5oaWKnTDbP7ErF5mKaGxMGB48AthJ7Si0r
uqhgZ4/uzfVTA2yyVbzAHII/Ilq4ncznD2ATIWjBFXd5UTXgCBG156F9OLu6SEKs
STPYd44kq4yhxIxNUQUe0iwXrJO99ZgVBqeDGqL9GXtzjmEngbKNz+CLyy46rN2C
HED08I3DuXcAZHPQaDHWqsRe/+4i1GIxFfzBfN8dwVA2de7kmxAxtAg7i3yKpa2O
Tz0ac5QCGYISGw+TXSTHNQGJrCR2F0U7i5R5DDK1STZwDNYfR6T7TSBkZfvnyytP
d5R2F3M2VnRFWVBEnwDmCVNoI8UNwpASXDErvlDHiaxfoRAL+UrC7mtDtU2LoUQf
H3W3eSxXrV7qf38l4WJKcU+C/l79DLE/oTv0ChPtft/G+TTIBxVsWQ/0zDhpnjgE
iZK93214u+R5yQ+KHZASxi6msamSBhSYImZKBeYWwS1jaBT4ZtinI4N0SFeu4wHt
f1P/YyXPDo/nAcAG/rUGlsXgXYQrUWghecOO1c1rXlBGmmysVUx8S5Tb0lLxg+BW
xugOR/QKXSIFww7mgT6Y+ny8aS5w157uVzncuEGCdlH8FOmxTEAYt8R2HhVT29FK
sFx6bHCGUbHu3IEJPOjgRQhK0Gx20F6GWEfNlSYvlf5nvzZ0H4lKyW/QWG8TyMxR
5AJIPtFxkYG4l0aPu1su1FN1Kynbq6mi1sOcywtrXN6JpjbJQvuW+hVjSFRs7nYg
+yLjcyyu11I5n0rrZp0xLetPy3EyoxbXwCnUzDhduHs/2euFPrvNjsa6TxNA5q/V
twQZMOwJXM9n1A8H3IApLpZaRyG0R7qVH0tV4BJp8/CGfqLg4/OOpsmmmOjpseE+
eZojvQMysq9p/axj+G/iQOSFaaFumOy1hV+SYp+68mxIyGL3sbgHE9TsvMVd0xeu
o/DypF/Q0OVJHT1CduQR7VLJOQaM2t0yPPW64fVbVg80CCJfYV3XRYBX5Xa0xM43
HeoenDX+Opg/ZunFttIT/aDMbHxmeqdasrHp17Rfk6K4OU7tIk7w8OevLarUEyaZ
nqHNgTLP8x6ck82cZnijlr7kt4zphxJPZY77Qgd2dlTWQftVj58GTPV3gxBxR2xa
q97qZsa1dWvn9F1oEoKgw3oEtpYlr/TfCbLfDHlPZ0VPlhLoVorxJonjvunOpRaW
DgZelzRCt1P8sZCN4lW/4+7hA6LWaDh3LcnlzAj4KikbkitIgE+Qyy0T88lzqD36
ruh9fui0IhyojUagmWAILjxu8a0gHYqtRMzZi3h32zo46hBE6vqVv/alOLAyrUoA
hpN8w7KJIU84Ue+Y4sU3om3ZJIqCx1xbAdrklR992LxQ7Z+8Lr1+bXdNbUtk8/pf
6PUO6+raZptVeASa/BOWtGiLALljSWi/iWzvdT2VL52ISRNdRt22E/9BAr6N34l+
RKjegpbdHLehe7++M+nN5rv5rTdZk0Kl+3UXJ702zJWzJ8Nw4i32m/X7OC1eMYcu
4uuwr8kd8qb3lMS0JvlFfJ6MU8UzNJvr+bg6uPAMX2aYkVf3ZYFL2y0abZjQANps
bp/+Udj/k2SGxwTOJX+wzKUqD7Q9kbJkZeysUzMPXAtzU0vZFhYLGuZyoKgJTKSv
zwtGC90RLZkwb+HfOUZbaWe82wRR9whhsYf+AyzHiTR7GP1fs3YF3c9YPRPYylSJ
r1AmHrdPgavjkuOu8wPxqCLPAtyp4xLMxfNRVYEK44glHLOtEGdmCKzQV8FWg1uI
FmriALa4BsvDXVV3REZjY+SNDq0+AWJA3rJxly7B+Y/tlBcdToBzoQ9IRcxDp5NH
24WYhHOPpa7kyiE88luqgRLAuNBa/vfevN+EBsgpMdrPqDFzbzkbjyHF8b+ovAET
epu86UmQvs8+ng91RCEvKIqYNNJfuc9IS06m4V4lLudckQTTESxuHhLD13wWlV5y
71TwtfhWCI9yAHyQiZVu+ET04f2YAJK5vEUgbJvHQuJV36oEHMCJWXPKhmlVi+HD
KEs5kLzwO2Xj7QMUomLQgZnyyz+nZndBQ2fOr62FeUTtjCPko4xlWZHF3EyYL6Th
Slavya5GqYPgfGzel5xrEdsUw603hSLpklnJPGv/CnT/eMsAYBPiovc9QbBoKCaM
V0Q7ylPx72mtWe83h+5HwU2jz6qy2rcC686ky8yL+fLp9x4c3JsVgnRNpJmLrLs6
u2ID3Bphn+2OhJvXIoBlUqphRIvsJK9Hh8WIPwOkhtoQDyJiq2biy7KU3rS0Wrdh
iHfvadNDQ52UGmfcvtk1/07Rq26WoOzfGmyNaZjVjD57p+VHO1hv8sGZd3mykwy9
JajVaUhd3RiHCJyUPz6Csk6N7BYplBjElzwwWB2HaR6NLFNoWTG7ToK9eub2Uvdq
FhSCzCpslu2VNidmb4+86yUd0VDZDXTX1ff4LRVavIFaO974VL1k6iN26JSJFCb3
F2iZGwfaBKUI3L1CFRyeu9S4YlxLnWbv7oxZBE3LjhbMP99YG37v1BL/6Maic8zy
wRjYCLLsFJPwIgyAUdWHDkf/2icV0gZU/96MXPQN1sSnZVuWBUb3hkhl1m4qDu3G
fB5g/cVnCwzWkUaGyxvWmd+7Pce3dMRq2m1Cnuvswet7/e04FHgnxJk4260soCBG
R/DsuGr5rcvyQaiEVPmb7fyD2+E4Hs9w8PjYdfzcoJ13AVZswtgiYjREORBYtoyo
r/GmzGtVU7zQe6wkH4484N25bbUQiqr4JkFxNWcssfbztDX6j/NV3EJdaLYj9Hss
tBptQI43uH8H8e6F1IsGecy+MDw50iV8j8fd8UZvHxhja2VC+sG1shuHsFOxasv0
F4gXcPgc9sc4WdZBkYSIUaI7PQs4dNJMvryPT5attGQ5T/R8DvZV2/c+8uvA5lkx
N0EAqhhF1csBlYI49HVT3QyF8qz4sJKrjOMN0mG7TO7RnYn1q2XPTs99AU38mcxo
Egtid5zCdXTw+Oz5MT4JVn9Z+ABoAGR7LRLiSyLr2lQpbi53tUAjiwnTx1NK4DRZ
RCexCxp5IqVpNN16dpmnosLLRwzorurY56GS96wDwtdd9usLFgUCBSvhe22htw9D
5LK0BkBcs2fliRAUOIlv+DGwjZPRJ0X5HZ4aYloRDp/O4ZZvVKbsO9cVUbo3XIRC
v/4PC+cpTaG/KwtpDI0B1NQeFvi8cfzWHlTytNNp6LDczQdxxiPLeKE8kLlHjvq5
/JKrtxCHDhDL+cLSGo9JBQMMww+5H7QNq9+q2p0Q36w3ppP9NHsNUN3LwGhXak9F
0pElu7p52dJkEqsr4vEw+pB0Zxq9hN4rejEnG2IBkDXcYOfyZVcCfQlEj8YC/9hg
NuaxFTARQv1lm62TwmI8k2oCHhsy1RVEbFRACidMgyml/jBaFUGGGcFnD5+7BPmi
y/GnbBnnFRsCm4N4HghE3hoLRD6CDCXS8jwZcfCou58SJQozxDjJDDV/o7txcSzb
ukGjPxn5dUHUzgcHHHMIdGSleZZLXvaWtVgKEYmP79BCTZG6zW6GjkM26mX8bFC9
2ioelMgcCG53qp9QECPeRp9WtabbXHeHrsiflP723vSNbFviqA1sB5Z3ow9K8y/z
+4sZ+LjzJtF46epxJIgpUwVjrSUwm+5PeGBfy8NJ8gAWVfcj5BwdU4UncSgW2eY5
r0b53m5PathXzaBR2Vklmxs0KyUygeLuAt6ZGBwqINUuuBCXSin4WGkDwFzWGbko
DInfXfXLmYl4WmU90I234RbE+ZTks0fYLpUCB1kNEpmDuANltKVRZb5DIRWqdQhu
1Yj2gKE9GN2lCaoAwBemCSed45GG5ZPJkbtvEeaAdbXWySSZ7OQs4rRa5hAhxWkl
utJ3MVoww9lHgE/LlmYZc/csJ7Z9ma5mLr9MaJZyhwiYjBG1xpow/CpOahBGvI25
dnDTRc9y1Im3J95YVNJPFjxQV3AqOxELFAgNZPMdnK11YJnErcCedACbD7HeR9Z8
xpAYFWSJA5FjlKb1Nu96RpwXgEPCA1N/u7R3fOc9SazZyzksWCJFbUfgBP8XYDFf
NHhN/slCOyiSyFlMYCDbDPHI1+FWncl/s4wxGIVb6ksLdUS5rSGmWT9O6ZXxCIRG
y2nbv6ZK30t4k21Wwd66ajJ/BehL94Lgsy8oADL2yDnqkm6DnjNoX4xzLEyb++Pb
vpOTFEd/9ppRUp4rmRz6RlBQs/stnYzdWknRM3TICNvPHs73a1NRcue5AM1cxNCL
mpd8J+fxcfeEhAW6X1Ey91IPRmihHZHYQ0ozQq/HD6q6oAE3mcgfx1m1BEpqFCJ5
ZWw77/dR484pxiCvEtj+OU3nnEk5e1RhQuE/E230Q87Nk6a1mIzlacwpDKeGuTd7
bXcRlvx3LBogk+AEB0nzxtBrKAGwUK3e9sV6sFfNA2LFFEWaOSHAB3L16CMfdYEI
DL2nKwtRStYGBWXxkWX53yOk5fCbAUs0YR3U1NpZdobH2rWqPMtHTxngQ7CCfKrZ
zmN0ox5wp71tzlrKzkC0BlYeIqBRCICLDvkQTJjrQHe0sfudelOS39z6JIrcRGHw
HXQJaHvj62Lllyh1WbX6iTISGZ6TqpUbvTI8DOWa+3a5yAO7TEys+1yofu3ku1+d
u009cez6/JGPWQVFQAjrEw5H6qiK8zc25fkY8mIZQUHTqYVGcZxV/lMnLMqZwcQs
xmPgWALs7Gz2cXzY+OfTqWVSijWtsagnV03bSM8DbvU2vnyGvOWJavZ5989A7Zj1
fI/+4pf2PAlP1a4+4QLYfL9+ne47aGoQe+FptrepXHkuJEeTdnz+SHpKLuLPXCJC
Ai84g1jqshEaxnXHFcTJDlxXeDxkiLk9tKsB/78yGUplw5dVhoBhtjNUf9YWvoHN
UhVqp+8VJJ3o2OGzcAeswprD1hby886egABZNF5qqd/lDpRqLc+p4LcihvLseY3n
o0k5L+X/Mc4OnueSdKuvIPrYwLTHFwl5fmPLzr4JXn58gjhT5MHXgt4/NBKh/NuA
j0qw53T0VYKibidLXh/lVECI7HkDyeeOlgExeT68Vll9YzkWYQfw3jocagoWMv/Z
HbvXC8gouFEfqMs+Oe8d1NfL5bvUD67vxx6EoTEOKe/4CgKEZJ/+PEVcCgOi3EM8
cJyJLXb2v/9Fk2ee5zGE150ma2RO5LS4H2rCZd1bgcXGMo8XPNFdHDg287kK5wYC
783VbmnFQueIlaANoxaaLlhThhGufws3nnQ1bV96W9pygsLAv8qFBjZJQwSqGXbe
j7d1p3qlUdcVche5ZNySXotKkuN6b/SQYizZpivhkl3iYhV4W9A+lT3jwyG8n5cg
DG9OiQotK+Xs1kg8NtvN59xNz3P47EygvZpfThVGoAFPo3obU5kDfTXTZeTcJjVq
vNIn/DHqnZ7pPOF4NXnOgLg4uO1XsFpx5L3gSZ+AiOJa7cvDHQQrcQxcnBm+rA+g
MHlYfRDfX4OR4u5apbUSVs4GJrpMLUcSntSHXfJwjTJB0DmgM8mbIWTmiYCf6XGe
5F8pVKjrU2spXM42ffkWfti3CfSUZW0RVTgLagbiwu0gV1vyK336/nfDu8GSgbto
dRIdYtCGH1ms7V8iiuQcTEo/3QkvWFQBdQOdi2jjmTAfnOdwtgXNgs/WzBQ6AkH+
tDPkNHR2LnZMQRrzns3cu8vbM0y3VLGtX67tRNcloBFm6hmeOvYwPrh7dMz5LrtJ
1neg0+jUVTyu+B3k4S563JWKPkVUPMXiQIGN2NQ8xBcqcGAuw4jrfj+bB4f/eU6S
0r7PEIUzAMpP8AmNA2uIHwVRpPLgBpyHMwZFnqEwgvH4xOLDpqNEl65iiaihzm9+
wx458fSb4Rudxmm/nijJ254zMH2C1j8e9o1oF1bJV1Cd8hXLsjcjdbP5kfoqekWb
5GuxNSfUX/4C/jLihrkpBpxSKt3EWk3zFK1eBZLnmk3h/DQjcyzctGC20XXQ+d8j
W+xl3LklSvX6ovlMlQANJq6Bqs+Rbz4r2fMbXS3pq5tEqSKQPuV9yx81J1fUeeyJ
S1UdUoScr8eSTcFMGoP1w6SusbpGb3B62X6NRAvbG9QxcnYW5j+f0Kg29gN7P7pE
68CmfOWCLsJjI8kBDaVSHJ+McnJDCqI4X/+LffmumkN0AJj2At7q37gJadqhiOb0
tcH+k0EXdOhEnc6H9XhUh6oAlt8XZ7vmV43SHWpUjAkORckYJtIe7u+FzUCbA7Y3
z0u2iwEw9jpEGvfPHt+5vDs7V4pBrCKVQ9Kzsjzw6ccl4LjLM1CalsUQVY6Q7MZS
2BZrhlmxPJMTzYYgVMREmBXI7x7ajC1SaDJjvYwPIAxAefufTb3feYdjAPhIyDdh
VQ/3N90h+PiRSHHVpzMWsuNinEWsWrzfDn5TxflJVMleDvkmRBdKTuWpw3NhTyD2
276+31cmkZB68UvMQJGbncA0Ve0OMR8ue4pd7v5oGsFArXRjWzVKS3g5v2HODRrT
PbU7i4CWuoNyiGom3ffH2d0UBBGSBOzn3UMv7GIviAS7QMl0WU+RsQGw+jzmzre/
euTk4AnlJsvfukkhhBRR+IcAEFl6RtoA9MhF8Tjj5T+QtTwSCSNq2iTjfCl6ln8n
fMzU+OhcFu2w6Q2V7jFFU+MZzCfK7YjGeptIuuMUs0knV4fpCenv2hcSr/oh9lRR
EwTRhDIZpgciQMpUI+pJcqf4FRLclAheEEngWmcBc+Q6nmN6QfaR0mkjGUtvoIly
W23GWsYzLEOhXPEguMPL3rXhHSg59QOfWYmthk58IWN/w0qKWIgQYPdrUisMvpCo
JZ6ES0t0tRYv4xYaVFGRznI8WKUOhb1CptpCPVw/6PLKbpMZ4VgpJDWzuK8Z9CEw
wDvmjJ2S12Lgf/8JyAwIVbfH+iaTtfnoUYoxJz6kBi/6TJ0oA51IlvFzlwdT5yd2
mKjlMRr/Xy9n0f6gMMSuJ3+hXKhUaTATV3cjlk4ibIEI6a/M4qdUcYiveCdn99/j
+iTTyoFhuVcG894N16huv7cf4zminXWCWgsLrR7gFpb3O/Z9GGA4HIDL6yf8HLZX
3//DyJN2VbCEpnbT3naS2jY5HDmJKNBV+LBFgSppS5p8xgbG7qGHALPxyQ/0ssNt
+lyMa8eSlIzrcJdUURaKoXt/Di8n0VtCOQi8k67XOrTeQb9R6v6tIOiUgaFM03TK
ShVJz5VaUhVn+AOzJdNh+vU6blsi+NpzF1oFITgsD8mSbJi+bUTIlt1ObjEKAmVy
Gsoc9zacNVi2i+KUj1EC2nC1CH6n4ho4X744ReVWpU8ND/BuDje+rFjf2kN8YYqO
c2lEyA9rwULWu5/TM4vIKOhlxG0xBLe+WtUpnFpmOTrH9VrX4+vUA0cqC0deQbdw
qYWXAHDIA+6AEIooQ9x0OOG8By/bhJyf7tjPcUyT/Gxt5jIFigM+9/+VSnNTDI6b
WpoxoSh+rJKDphH8vG5jxB/EChtKFR8E1+i9ocL3TIJs+BYBtkzoLsz/AYVtrCSL
pYPmKdy3MMGX3kM0s1XWSbHqIBy6W2sbb0kQPg+oFnra6CUr5pYyMdGqjmmWDtcp
me4dpybX9gJfcCGD/BlVUNHrWnBZ8REuoIjmkb6wJx9KpCGKm4TPp/LEt2cvZRmc
tyN9BzxWbFb/uWxkJJCwuMBCnEFGrsVzCwsTauJvazOwbZQnTVpKKr5mKTOtM8GO
OPhyREKQC1RQvcPhNOtceDbR0wlLufDVUV/dysiI36z6pdOBAtgxpQKM1wn5tfF2
s4ITgFNiFilypwYdWY0MNbvECC/Ik0tuc30alLWZzyZaacSMuK/gbMQ1I9n2V1/2
0hY1A51aHLlBwo1LwQduSsNm+gT6kjrZr/GNiJjMrhaPBPYXeBdJeZnoZ7fpWHQT
b8wunGiRY8tD+Y7P0eZRUXWw4LMJFR9sfpdfRQT/pm0alkZ3DVqP5DG+soBRdDYO
RL5sXdCf807HQXhgh6y7zMgjJT5yy3MbHXUKmSuMy97e7AFFNAhE+JsAqShjm6Ih
KFJup6UTnWw8RmznWhV0gtqG8V1nXtcSdomjwUnVwcK4ngzHDDtIdNRy3abkcJmb
Bo5sF5cBghBefq3SL4q7kdaTkw2MK2wDzNYGq2fmz6f/Dz/KzWSSzdeH+DGAlaVg
dGWnj5PMSIG7inpP6/DtirODlVn5LzL+m8F//3BLhVJsUfgWcIj6qclmM4cwkNTT
IQEN0KMJKcJ5dzm1Ds48yUphe6ApJ4b2kfHEsd20BICoKcK87lNI5FQ0zO0ylloV
h04MqH86LuHs6nTwtCAddZQlvcUL0fslauPfPbquYu7qtXOjMomoy1czsQgFRe/M
/oPrWT5RdShzaJOplxIW1OJsl6YS9IldRBNFIJaogscyZvx6bjMccC20jrlTG4ab
LVGEIMGnR0hbR2G+4WgWtcbMjT62PifnWi3oSmW5I4ldyl9ioA0JJ2OiKmH1NTFb
gVU6ZHxI0I3pXvW0PaUGBUyc29Job/P54wvZ3Jnbbqd2JlapkNimxl9xb+MjxTYy
rcMOCutJa3ZXk+2Q/tcEIs5uE0JYelIIqX09R1NyM4Q0Ze0a+dHTnVbVBTTGOV0N
fb6Clfa897xQ0TlVley2yUuBQXvoAL3cLgcetNIS+9KvRvWAIXHOy1OicY1dPVq7
1d04RBSZqRYdoonnuFqVdXzq8lkTeW8X0/56W6mZsRrdE9O5yAnhf9SDVxa/EjXk
choqNz63cGYhocG13UzUuPFZ1fAjE5mWf+FL0xkrY4+rmfcCFORQLzzKibqJNXet
Ns6gft7bBr8B8hfWewHyBP17Er+kLy8pZf74+CayJU95dOkiEiY6fcYyem70ii2+
nanOvRz7zEvOFgWh5xf57c891DYbzJGiouWLpEwW4hnNZuSVZRw1Tx+NK0OgHVSv
jyed3c+QSSkFYTfaIEpO5BcPe98bFat/EWzPjff6aLIIk/p84vx2yTy13PSRvFXP
nRS6VruDswwbDRso5wGY5rqwo2HHHDs9+ziGQfQNcZud2s6pn9zePvOH0nsUGPvv
se9+lz2i0npD3WrwRqBgfGbjJdbW6O1kUBpb8fS1GntpVjgwBSm0awDp+nztRWGi
1msdMnh4I3pYHrzjN8gh+eutk0liKeS4J9iadJHDbZmmc1anVOG1Dmht4LJEm9aV
b/ABNlcr91S+GfBCrI/qG0ziILtujclwY7SftvkzQrEOJCN5dYBiuZHichAjz8bh
yfo4HDisesJ3iV2iI3ks6RlGEhUKHEvoLUWJhFzKXPQrRV/iLtOP5W+cihPgLTeg
VG45Pg3/WYDMqPo3WHWFuMmAdVvVbWYamtbSAYFLHegoyZyvBLWc527Tm7oiNgQa
UxqKyBRWAKvuWIvM6fzv2KfSzMoTsNyz0NbkukuM0EqEOzNUEbo/7JVDDNksIEh6
F0K9yrFJYR2engKSYX3g5a3DJwnymMX8/7hhAXis/J+X2MSP28pfmVj+Ff77+k3C
zv91pm9LXRp0g1vImBwLSJIZYFitSIvIjJxIODk0DlX4jFKJgn/OZuVAwfGbi0Nm
kOvwega7vq1rnGuGEa52IVIjE0ELmy9miO1JsLCfFPOwRUVKS6JzFdwcrcNqmIXH
LTqxFtEB0YwR4E9rnpUp1LO2Vwl67hMtgaLIoRRATwZEaAH+qgM6OMgWrfvAJTbt
lASWt+HNR6h43xn4i9Pjf+a+4+eWSS65qgPv65qY+CC2jMZ+OnEtCKAOsZzBnxQV
V0UFXMPCuL/l2KUu4EOSJN6L0rNwViEZ8l3um5WUOQ9QwaVCQvmkVR1gRg8tbrGC
d/eIi/qL8iQibrlWNF3MVaqTIbj8KJBZLioZDfGZVtZq4yJQ+evj2n4Jok3INnpt
F+142LZ16Thurgw2n3ZiIrKbqsL8NwQIeRxx8cRAd8j6Fn+utzBOzHMJJXszylJu
/Zmysdqqgp1ek6X/LNBQaM7Q+Q5/ff0sEURd5LmmoAe2BNvLlsYz69t1yO8/Yreq
VWx/XWHKt5SXN1jomq6TGgGwOR1duIB5w7I1Lsuo6Yhg1BQ2FBMlFVRczUiqLNVk
fLjI+7TyF6bLu9677ksZX5pB4c42T9TZiVjKxxHll+rV2hS3QJCUkZYpAdjsAnVm
/NrtJhPpYFMpPUb4TWmhgM+XXNrz06S16EPbzJe17hxXmyzMzNWqL9tibOnHLLDN
pDRCVdzakMer8YV5RCsv3KvwEyzRCm9CyGF75sNZLTqT0lF5gQqirR3A08TOwdHq
8/I1h8sOns3h08kN0vTHz4LSlM9FaULM7qWpC1K5j0VjqyeHu7JvIs72Hu/5igdM
2muVHOzHKaiGsTqUHpO526y6raCt5T28C7oJFUiCb9HMytDErXXtG6e98uomwh6Q
dHS7tvKY6sZdPASLNSpm1tM5vKoTUgPiBlFQRSBTyK0i5RyuTQCsdoTvqU7lKis7
jgksflx33vw1VeuBBI490rreD9kHMs4ErhdxZ1RFAZM9LqC4w/DOAEcgxIyp/ZfW
AGEoScfW5OjRm5Av4yCBH6+Mm2zyIr2kUBxS/+CbEcyCUF6T844JOiRk+DANlxYO
7dhIRzRBQni08RThUaHe/2rWrAVTSZEaRoR00Tz/Ynp8ve6UObhKDX1UGyka3nqW
cPJqRTKJ38lS4puC+2Xhw7k9Apz1rfvX+xQSNxZ4lRtpJ3KRHQz4Br7o7A7miAIZ
vwwlj9VileEe5bb6hAtmc3SJl478pqapNcz2Ew1ITmdsQBy8AYLE5n2HA2gHHVp/
YtwYAWydTTj0jQL/iVZD20ca7qz4Eb6jC5MVsGb+9q9IAmQR8qYzy6WY/T+iuVPq
Ri8WVQOzEnWXAHRCPQicT1q2Us5PAbBBgR8MAerpinkEY4GtJy+wWpswEcbvzRUZ
KmP2898LCT87cnYrKFuA5xQGAecmQO6OnrVP2n1bdYN1A+7aoJrgi3c9rf6mRGBD
OvW64FCjdI+AAbqUwMxmMX9jXK9P5T+UVhOxlHeBjA1/oaUAWEFtcnR/tbXcZN1Q
+VRZnTM58lLUIV2rlLIZUQ2icFbGEPnmJE21Pn9MmuUvze331q8STRRkNCRC1s7O
0ofPU3uZzDPOCr2WmZxbgl7exto/fVqLRKZlB3qx0VzT/TbTO5shP5+YwLU6DlRH
6WUrOjDYewjiaMfY/Bd+WCGiMfbMT5uwjojDLJdanIJf2vsXOrC80JTxD1BOQdFV
7ndgIvksdmunCnTie/b+z7lZTC5JqjNAGdKRU5taYpq4qnKqYtDk52Usuecc/M9Z
xAibZvd2U7YGI6Iw6HjquQdzuMHrI3b3D4ctOsQClNpjvtruAbtkuhPZrehmuqgL
E3cwiNpUCuyrV7CwzO1md4lWVygJJc3b+DIcw2ZquhszgQG7J1TPRqVxn6MyrgRc
t10Dk4MjuvzWMNq+RCfl5cSumgc2WEFItv4xSwnz/sPiCvMXd+ScIVDjJy++4o3c
InP14GGqQhnL8ZTc54AUzLDLQAmK/LfCV4inZmYbNbN2btyEVDU6AmmUch3umbb1
4MJrH3McbHrQR4p2Nyw+2IxNrylTLxFV+UCpyKvYnObuz+v2rir78X7NvJ8aQ81j
n+rZSFv+6Et+pOfwCofXD0r7pjuGXnFkaD+5thYOlFmj48UpygJHchYZVgUBBleK
EaNT3X1tiPerCWBpEF+mZcRaOM/HrvXFUbZGfCREJUEzHB5f2UF80McgYh/djrBH
+dfv3GCbtraKZWhp7kdYF882mkI1jul8c6i9zme7oiGT3uQOxDnRGzVZYJ0lmvdV
8SLUdEz63Q5SOsrk9rJXnKzpUsF9v9LfaJwr6bOmMrKZP++08CyCFxajSUydzP9+
7VSZR1Z4sc+q1Cg96+4jrOG8QsnX/iwkijVQpP0oaA9JsfrsFD74dWhcgprhG4Pq
eLulMBcGCAbUxKCacV8syOYbDUc15YM3cjv9UNTLrO6FNsojSDBS6IDcdgkiuTJT
rd1XTb8bn7+K6AOmKJl5sfLXrIjmFsAhaoTBlXiYvpDGpI88oaV1kSX91M7DA56S
FIemm+cQvBYxNfVecB7d3oJMDvqoRsVEdyXQN5SPOQGA52nF+8iA3jMayL0sSXjB
ncD5MMXqgcJXeFleOIO6pK3m8bGZQqnPT0qJo75+JoUrzIUSpGaa1PB95Qd0cZnH
R1EuULSYfrmtB/VmZOEh2rQTKwMXtJOqtCs4JO2bNWOKtbDjR/JgXzdkCO79CRBN
5joD/xCGL0KJnTkmHzl3bNnK+iHKbvYOJdBkbzYTI9llCsj5utzVhhbXzglMQkCU
LvGYgjbQtTLoZTfw4hL4w8B0RO9F/Vdpl2eQ/xp6xXexZblbIYkouCogu7C8CE2w
TyA+UVHiqDX3Ro1ubWSRHJ4dUGYa5KgkNycRbF0vRq2CpbyiYPJIgPaWJuyKiKRd
hhbgKRqVl14TItellp1aY/cTKywE5J0NQxLf6BqqaBjHF5CS8zR0nBbVfUb6XXkF
1fPkOOl/03b9CTmsVXFCbrHCzm/OwvaEZCRtG8E6uQpgLGJPJQrSObeB4E3RyXly
HTR/8WamC57B10tir/LTuBQzRnuYB39AguhPZiB8X7RAkyrkWTdwZynajz6+w/Gj
kdN76wyzxAPwY/0riDbgKf+n6CGIiAsyqBB2CJhQnvVBvjdh9x7X4WmxEA0ny3AE
gut7D6MClx9eIvxrGymJDT+N1Su71JPHcF4uRU4bZF/s0CXmkZwKRvWTedU5htjb
ScOQRNjbd8lilEea15BjsjB6pBlHNPph6lQRpZKv8a4lcGxo5aJ6i1sGkl6OTxU2
m/3VSK33dM/ooDLx0SF3hYZYYp2896iCo4+h7mywDDQYbp/aH352CwYlhEFMliO0
IZ1XJInwbGTNAI4gQ0UCAoEkwUfmQgyeqayCqtUmn8f3kGhoCe3BaDnbuFJCF94o
HIK5wEe1WMXL49ndl8cATN46KdSw+9BDaHdzBATRaF2pWmzO3FDzotGTc1Xr0be/
RXnT75q5d2d5jkU8+D/6EMeblFRipHGySDv1FpcDo22l3hQFaoS5B2wkOoJFl1CD
uMEvvbm7XUYTv1COh5vqKx+rnWJJjJwmj3LMj+k6qMUW025LmBRdyzEJzHEyhkH3
IEII/9Ak+pPd+yDT7aEOTq4E7+uncDDxVNfp8Z+KGS9ht0VjEd4o/AtBFtuYpL/1
f/54i5ENS61GsFLTRF9Zl3SGONA6M4Ka0EsPbEsEGHkUO/ZrG8h7znkcX2Eoig/Y
0dbbolgkY2PEJR01sYj4Q6iDnRdAU+/mH+pGz/xJTDOPv1sHzrFYRwLw9NLTgZFt
IAtoOpTpMw0IM7OwSQxkkLsRorO80GGI19/L5m3BSLa7WD2Le5eiGQ9RoDsCC7h3
0DZtu4gCsRE+GVjDUYvSNCM1SaaNYYO3UehOxCX8w4jlcLmD/pJiU/4ZHsF7SRvo
BpnokgU3mrT7rkgErUH7RI0h4o0AiIDaEkaVSxGUmk8AGJe5Dt6wi0fIikHQTJWE
nG4cyg43LuDtV7XYF+jFPvaB1y+kc8ifJNdbB/+O7EIR8p9BrYEPoY7zAIlY2wKJ
BWNjO3OA+IfegYK26I+Y4KjvESqMrtz9yVq2qeVTDHpHr625fN6sgnuyNiH1md86
393Zpzs8Y8B3x6s87+8zxVWQnUK5sL8lK2VhRO+39swq+4Dy0gRArCc99MaTdKNf
nxI9pAIMiU3OE8zyn0K1y2T0GmPhePI/wSC1i+7UNyEMNyQmWD76l7bu9f7wkHuk
cX4NdkHU6WZrGlY+NsxrGkgBR1SXD6u+5N6Wz+YBbZdo0+viYjbm0LgOb8ZpKVSQ
pTlQrag/eqXbEKM/AXT1BrhBcTdcq3IdxrILpJqYjm0+jCdOUGanC60my7NaBOOO
txjSzv9rd3c6Zd0gT4FnYlPnqStJSlw/SQJA9l20Qx5eF+7s1OqHhpQJFzme9Bto
PNCnePVb7QGU5dFAXhaldKPziEPfCoPYFOV8kuUPt0poQei22rvWIYqMcOzIXpCx
kbyOXtNTVWIlR/fXQj+Um1nn97cFMtDbftgRVmu/FugZjPdwRRWRht9ms6z3xBSG
WrZKlVt9FXUElgpo3MzQV4yvdbiDDFVwwb5dAmG/TS3lr/NNkiC+qtBM9yO5DHfO
cRvfk3mYXDdlQFkXPMyR3Pk+AuaRZKjtXai5QiDSMlcxP6TtFx4Lc3T/oX3czd8G
6P9ABKlv15UxjajBibvPGSmkG6yg8ApjCWABfeD0TwY+Sp917FEGwR0c63YPLENo
xiFJ4cVxEvfcy55qpBJEDuQcvR56zY+97VgXxlzv1xstNdd7rZr+w4qie68uV0nv
e41kxANror5FsEu5NWit6bUj0SImAFg5vDN3OfvbHb+WSwLBqTCrYIywzcnZtK7g
8Lbppit8aJAc8XQSa0ShBh6lpnZZypakHzS/9XmpF+o3Gdpdj+Epb1RL3vY2GIK0
R1WqywTFaqPobREfzTRyr8yTlpy8IauBQ+GvLT6BaZYX4kf4At45BpX9SLYL5+Za
L97dUK/90VSKQWg/lAmWV5hScFi+cI0WI4BxFwg5tj397nCJDLFj0HUOIc8uAVuR
1d4Y8UD47ZN4NqfKxNeWdT7b1wGXOEupFbSRkCjwSoWBvaiqYHnuNqsHGJboh9oH
FO09b1IKkRWJ7bcEMqU/zEB3c5r4XWyIIDbq7+ZVJln7AAcdnkHvW2IV5WJ9STEy
9dA+bvAcEm2zw5SjY9qX9ESlzBth/6tciPvMtB5kMBzuyUmuXqcnM8dXqWDXWowL
vYq1m2q0nsfvJcTP4hmy5w6L7vQBY65rfBP65lCbu1YKPqOMQ5YJhyFyu4zrEXiv
/z048LLqEsbNIp9SuRe+w6bcXs3JP5jrUF/6cwG0QcFZNpKDpkEdn96lj6lQw4vO
czujBH85kYY5/An/7oIYsHm3STrfIJsE88hEGtwFMxWT3zh25izxQB9n1bbmqUBy
pNtGIHQ/9HqCT7KiltC9+LLpuhtL/Yw+gnKN+1KQmEMUeDNWmo6wISUrrPAVPH2M
DvaS7m3+S4hSM2Lm2r4+9GYg/vZGVjdUEtenPAdAM/+ewjecLanKX55LdulaFPPq
rGA4Xe5gGeZbVFb+2x7DXUXNLK0WlIRQlNY3+HmtdQu1SMWDwzRSU8Q7BbnriFAt
ll8KVYSWOKqh6xy/j3LwsOlH6uOPFrnipCEbGzanvC4LVR+xroSW5jKEsIRp/kvz
SuVtZepiRUM44c0Xbeg0XB62QYHYbtmNUWvpjaiIc+WksGKuC+FASh/Zo09AdJPS
OxZwGqfneHPAicqSuyEbjbCU/r1ElfMwOsv+2iXJRygvvQs1yPYK4CuGoRoCRyFD
YpW40nmKI+i9ONUyKy9VNvJshTVPcs/ULgLFZs3f+eSU5uG63cEcoZe//es9SRS+
XkIJeGGTlTL7uXrJ4U4fIYD5nwcrOA6KK31wdjo4USmsArvSLI5Srmsa3n4Y2Q0h
//ChvBPy7320CPzDMTqz7sUNOmy5F+j16Uj4ukGO6w3UMW+o4I283hk96Tr3usxS
JlbaJOTuMpYXquedAo5n8J9Ff5LAMIKoKED4w+k710kUsRt/E1kl7ZGb8kMiJ2jh
19Zivzh6NHfjKl8iF61KE5SkfD3qlHdmQ5rgn71GF8FLk7iLPp1sxI5FiJSQdcux
xXb8/tX8wbXziZtE3CE3ZwOFoIEHiGHWmhszKrSWh75Swljy8LrOxKJtv5hqNLMs
N9sGHyExi1KtqoQfRox+7MUXg1AvJP1gJHpfU55XBwxXMddcQ1eG9mYvx6GgfhPl
Be3ATNUXK6LF9D9KecNLgmGnyXQ7Rx5n6D0yfiFqT4aIj99Wl3ddv/VJVGASKf8g
hiX2zaRlSdkkZPGoBr+F/zGGy8M1fLuqYZtfX/cnwA9kIUCFgOgFSG+pkKPs3naP
qCLQ2XUdNSkinF7ii8iRpTRXNEDhbQbvkpin4nUbXqdaYc58diSO6sfrmBxNJaVY
TamS2Cvum4kR611CMTcHDq6bH+0UDZyoGSnmOfvE1Ezv8A1lYAScM1yN3f0ksW/O
kssyMdZOt2ZdavR3Ey7ASFpKUkFoIR6VQsapskJzuXYl2dmFlJ3j8DfXzR+NJ6w0
9varZVAOtId/HvO7O8uI6lt/rnD8LI+dxlL5XFn/MjNF2mLuz3l+jvfq4f86VpnU
rPDE0heRwT6qiVWBQ90bf2ELi3shYnO4tDKcCzZqq1qCExKV8+0jyTko0cIsbniN
DOUnXu/QEqs5bCX2yAJVQDTdISHA4UPso+0DtVySCawAqVGVMx8xuLpcsNWoUunL
xN5P+QQvGSpwbBdzo4ZOZknmFotiE6uyL8l+7veEpYrJDbGOueckV9Etie82NUMa
ceJRlgSNJd7+R5w17EeSDp48kxsiDr4bnVqx8nUiZaPjZ2PoZ0lr3SFBJd3ubSfm
L4cOgAvhVg7JDTxR/C5lnHpVhvp07gwX/PBUYgRXivkZQgP+GIUQXEM0aE566SSO
G7/L8gRVKhgN0A1HUqh/LoNkJRCDWW/LFoWNEgw1AEwieU7q+oC51b7MKS0AqryM
g4SNGJftB4h+WPEq+nrlH7rjz80/WQG/kUwMspw4KAJPNI/51KV1XksW6U/I1c6U
UukmbcqOnRu6uHGW2/eTk7fZrRqvW2hPhu2/4UZDIx4t1gwhS701pHgbAUfQ4KnK
aHLqLv2z2mWs3P3DHM0L/RRlPIgdsLpIiaJW8ZvxM80TrgNFFRSRGkFtojw9NVqM
jZcPFMz5u7RDf+9wMS55UVXsYUQCJu+rspbtKDI/YaOgIzIug1yN4Q0CNQOrfJPR
j+TSvGzy3LpZr4r4FlygVo8YNE39azEqRm2wKjPSC2b4LmceFCUdLX4fCwKPCcgq
T6i3bmiI6+lx4TpgEEp+QjOlRv2lQaS7K/qCnhYS21BspkEHdnOBJIvSNoFyzI/K
8wGIj956tAmoyyiM7JOct6mMY78Ru1/VZgHF6gZj7T+Dsps6egbb6eu3qw+14m3g
MozrN/6ml7KREWUUygllFVCK6ZNtJaGFOz97O+LrHh5S0GBgbEEo1N6Ss6V3gMrX
Psu3KKwQmX+LzNyCHrj94ueuabfFC+3ZH52C00JQSMgliE8/Iw78AW8nFE9Mqb/e
zATbZe1E/fBFs+PtPuvGm7CPW8MXEldgTXes9xdYx6TDQ4WHXhcKOrIhwm3HQ5Sd
AvtBqfeWW+DBlTjix9nCIsW+755xRpRyIKq5sVPo20pD+cTeox2Nv5a12qinpnEX
kGfbI4WZO30rb4IWjUlkjF7Quu1hOi6TQsgF7NUO+h/ludjb2JYgWFjkEggbZTHv
HoMpFh1tsutw2tXiZ+r/L/s4BXX7rBhOerKYmxdpHvn/mIhREGREoDgM9gEdYTcD
kCJhSvfmAEpz5xV/8InwWgfVZ2dVq2Eh+Gwc1HBR85VbhVcR46jJtZV81jJtuen7
qFc5bDq/WYlFdqen289j5GPU+vwe3qkOtOudGBUO45HSX63tbur1bgvxBMBcKMNu
a+3elO7/KdG+zXZ+sybeAm8kIlMkxXebSsxgLpZWTSv0xANJQ2DhIPmrw0DgFMuV
2WaXtqY5MAU3haPwuE841Mmab3FIVjTJ+eIYJPescjlLJBs5CJukY8cr5qfFFjOL
Ca5bsviNIS49wa9MM/KVW8O22IbbywI0IYSEL7LWfDAhXERzXtBRTxqpC0w4Fp7a
d2BLyA7OIEejE4KjYb7rU4qA8neEhXLGS7x9fBANTSTyhhC7/oYGDUlv764qkRCV
ZbXtmly3BjHF2tProGOfqLyBOI20r3T35Jc8Le0xeoFico64MNDdB6BHEz7kSOXY
Ot/HYuksziddW4zUI95EeOFU0xewjqwvSdrKUd/mR18YRuv7QY0DXKRaLBlDwLXf
ph4gi5eYLivyjJxpIWo49mIWRqxFPKImkCQo6POmlIdnrMT0cynVbFK1AY/eNZ6Z
ud/0Ml/vgV6cn+8liIsmJ+NfL1sLwhIVbtz0h5aQ9sER81OcJaMliq4gkcJnyw1m
WCIl//xBoXqIX3yzC10seOr9KyGUHiOgMRHqLEzxdHhN51L9V5wYpsz1xmD8OJwr
wmaj0BZxnb1gatHxGUPhBzngX0Hb/8rtFPajWYheP2ivy+e/tmk2fFg6AVFie6kA
dr8rpL7kUrDWdb+3vW+F1seOag0m1kVpVrZ9Vz59NOpCOn5d75MRBCOV1+2FCjsQ
1HrnLO/eA8k7E+HbHaYUNFaKXz6XN2B7SLZM6iXAI21LN/79pAnIivICcRegxrEI
kwFFNMrVgvGaBZfJBfC+Zo0wtkfg/I+DKUlnw0izKdEFX8bQ43sde/U57SoLiJAN
FnZYL/e9cFSA+fUvUSMP0BM8uxcqXGS23pzO0Oq7fX/7f4X/MQY1L4xiTQ1rXHe+
mYdPTTcw6FdNbxgatB9rTlPXkqbpWjUqZvX89QQ8AVKV6uQtvZ6EQ5UTEYmnwKhe
GSRid0VQQdIp/wVZVkkh+yShiK5MTD+9BD3+DPU41Lnn1ndK4lac5Wg711u9DWM5
fxbbZP5a5JVUD1Oe8uY1G5z24XB+Ic/iPsJ72mQDDJNV0F0x7ztTpnNfwuHVsbGP
lDWa2eXSMzOjJzPFwVhLlS1iz+/OATWCtjx2PJvcPHf8eUwhvISp+IeHo2QFDU80
sIHywd+G3T0InFOfbw/xXJ5G7SRru1+yLF0ut5AwILS1/0NDIlVRbAnAGbdKxkNn
6neBzxM2TDBBjt3PibvWQiyc9ruyFpHKo6udwvyitdp2ZhMRqxqQ4yWoj6lEMXf8
QedRduEjpY0xas13eB+7PcuN3GvNKLhbnJODMX7J5d1j76imqqNEA/L43mKAB56Z
EafoIL1mqDeefS4xt5o8da30MdgUbaKYMRmrVzKxEHu10fRXqY+DfQPy8lfHC66z
XZg72ZUrzk6hwGE3lkFm4sGOiEtCVQhcz3TQUb4SFfgytkbNVmERpZFON6zJRlZZ
mi6wtu+c3wRFHQ18D0T8bky+TjdwgSxxPO84YaUXYHaFJUY5vrCXSAWHQjDxjD9Q
0+Yx/J5dPc1sSVKQUKb21PEjhpJkZWmL/KwS8RAjv7pgNzwa8k8o2zuZghJtmX1Z
ZmF4sE57e+mQI4QNi8S8gQ7XN4gATsS/1wdWbJODOAIlgAsp8VIkgPAuJqKbEI+2
gqQSwCPSjiqZcLwmk0JBXNB90fNotNzk6fiRqjeZ9IQ29AogB4N6gWig1UyIgX6Y
PiL9T4J7G4JJnNzuTgLNHJegETdUUmW/FMo+MUUY3DpPSl0VLH7XSx6zKO/sdtvJ
sq9YSZtNlplM4k0vCw57YBwwTSJT1Cb6AIZHCbEQOVFMF0JcrNGx9DhIgwz2sb2e
/k9YO8hoiSZ4iLwneoom5asBYRXRvJ2l1ZoNhNndhPuJkQlOKcI5JoVesJ/Kf5Xj
qL86rrzDtnMBuy46gm5RDubcir3Bit8hE2lXAztWSz4d1UYk8h1RgOYRC62++F3u
gietNwuEner4YS4cZxSw6oa5A7G7KKeYTsBxwQHGRAYM0cCqhzSbpFkxb/xbkafh
pJDIFtRZkLmQCpBQZenNEVW/Ib4tF6CDOdu7/346PGgpvc/ijInQuY1/LROE0htz
WHllI9gfpHS8Lcba2RizKUfVXdHwNsyAnBLiIYYp34NZqbZFOkptcSHDBNZR+UfN
ewdvgp1Lcin5fVAP6g8ppaqP6lRdVP8XEFYGxn4lUnHwBrNjZt3P5qNyODl4tno5
sGROOufOiCRR3AZ1sqWZ7WzStEX/y5cPz1uoVcZUN8ze4CjP5zJttx2nNtjidxBf
Cr+xY4ktNMB4CwsJ55+gJltT6BZ+eoJtoaQkBaXEHby+30/U53fdeUCs8aOrGowG
lNYVb9mzvYDncIJHrSWaaHLf27yc1erbYvDiZtotnoRWe4kY21cBLuhsXWljvm0n
RlKX9hImxoNR6NlAfe1HeOTynnZTbU/Tdye8dve3MHgB4NGzva1B8vyU7O5+x9Lb
RRV0RboGwJrgITtVyCBvBdzhgeuE5iwNfIT4xJVOUDq8bb+CG3yQ1lOBFieoTvf9
J3nLGOCD3s9fWpvTc7FAVotHrTEWWEkfTL7a+CqvPkLbjrHgrIyOrJ0cXjNhUAbn
fqxG3ZvSIN7QXl+EMQO3RReHwICFiAARZ97hy9QFAP9KiMHhS9uIXAzH8VpyX1nz
EJInzgrD25vTGgrw1kcUOCK3e0SbDRiGcoDJSC2A4exWlPN02pOsHFCEdF04lGgh
CSLSLGalR9cWGc1Jb5fvFaBw7MZNXSDPAJB4FgwoGj6uqYCjyIwkZKWUPcjfmRWt
WnPAbqJQ8uIMl0o16OyTLtDr5w263VtNrn62ymGIVWpTnk0xxos0Vk4ShWhINZaT
Du/+cEbFyvNDPtWnc1bozfPfSeCEXMD3zBjU60b7zju1CParzLoHJa/kkq/0B2Pb
N5Xa5fxK4exbkBmOqEVKl1hCOWxSijKeW5Sqn8nx5a2KLXPr8+79AEO2Y9wCujyJ
46C5V7BhWQQFpcOSoPegS/xFCvX13CGuTmYl0qNdDfSLjEeUTnD3/lmkYsCiS1kn
Qt9N0LLHGULD/CGWYMw3wNum2W2JJsqK/5BFoLOu8noRWCUevM5aTAFzV7g1gaL3
pULIGOJzorF8N5ZBbxBKtish55bJGDp5shI2uLALWDlBmLSu4NvdiDPFnZlnFP1t
LRnBn0flrFmWxKV4DO8N29B9utylmaRmoGwvgPDxK6tDPGx6WNGJeNulTQnM1MUD
8lkI5cexh66AVT0aGkCz8jwTtuc3bGLEB8mRhzLjnzQftA9pEO6b0pGXEJTCEipT
Oy0N4fkXFA6rqU6QeVUX25AUt36QbRJ+Bvzic0FT7PM3xgb9Isz86/g/v8w/w6U7
wv4veT+j2T1vc04lMiqAeVF9MjiF5w5TLfk2oFx8vW8q52fVxVudRILBN1++rKCz
I/QlxrXDmyEy7hOHFoAbwg+Kb/Zd2pDT3QPwbPVc0uORcfghfiSZJa4EbXxH3MQs
12xEDZZp5XyXVQLy/jSPELUW6MNSt0chO3jaPp6urF44GOnoWPGLstRuuEjna5+7
IYTN8fWw/Bxt+m1ZlYhjp9QYmco6ie0M5Pc7gEkq3H5CuB/zbpq6c78AQir4HGgH
NyRxlwGMddxoKpjiOQ+JbbtFd0Rm3jFLqkF0g7xF9AQE8Vgk1kAbbMl9i0eIMyej
gSafmTqSNcP+z6xfXVycEsVLF0y2aqvevuh44D5Q2Qd3vdm5w79qmnxk1nbntIT5
ml69QKqYjdpL/3y77otok5lPzqCNF34br5ODvgljFfHu+PYkaVsJaofpcVJ4NDEV
qi8jWX721bR9+vGYKXwZ4BOA4v0d6U1bfrttYbLtWlFu5Q7+C4hOXYK4XVsr7qDK
A3rnCMfPzqIwhtjPSxX/WsqqtVAiQL6/ydcghTZ0dIfWRkkMusX2ZG3qhSMHH4Jj
hQm4MzhQi9XyZLyvcOVeK0riXlxfTEffYBA+uYmePf+BJRv+dVb/ssSxyBw7X8Rm
mc0HEoovz/kghPH9hhSbb365ngkoGDTuKSyYmGe/s9k+LBWSEZZcVxvqRRLHXyvg
sAMLZ67i9aMSYhXcXiY8fdi+CKY5G/UcuEL1uNDsl7KR48zrpNnoaw+TgNr8h+w/
y663Sb4KR6Q7CRilC4a9zlhknQf+P1XRPnGB9SErYyoXsCtLTZ8WFf9U8MUYHiHi
19JPub1o9UfIh+CDhDJnUE5c3b2LAmkq7A1cwN98QzS4bVR+RfDj23SofsCME109
fkODgAvszfP1pXrMVjJfczM7GXWwnAQQQ2Ea+d/we9LbjEKWlJTEzRq5YlnIJIIp
YQISxCYCdoGf9hHaNT+2FJTcYjXLnNu8k0LlMStD4MImGwaCO2Uxexb+mbDDvojF
OLjqU7hbqV7sGY1vq/E33gnp7G/yFKCjb5VGjERxpv6Ei7lo/LMI7mDqCa0TlQhX
vz/u+0fr8qRG022Q75Z63gpl8Wnc2en3nJe/VjvBMkzfZxv+KaAyY/IulF2jPtZo
hTGjrpP9gqTksyXsjbgGrsPk+SBLt9uBNdtm6Xb7Z01uB0d6v2WONqWk+67PNk3S
j3Kd/e7pKDTzqX3fVGCUOxTCQWnwdWe6ZjYDsfIkBGB7b4qLrEk7PiL/ddBOOU5k
jzTT7ZVqxuN/GxVsj0ZJU7kFx7dE05yYOqHL2z68LIZbnOo4bUaLVoMgFWTZ/jDX
RgFIM2HidqyYz/jY8mW6kYFobRuN4i/+OZ6UKEbKWYjabyqKPYnjiArRzqebi68O
RxYjtUHTuUrBhYFUNuDJMY2nwMe7962nQUSe+s2FBXR3KiEwgg05MDsvGfD4IYdD
p2i0+gdPB/TLCyrAP+0k3z38rb/MhK8YeN8nOKF8pqcGureKkWdQsC63sn4ixfJi
w9tD6DbkcZH8U20YYkidIKfQEhLmeG+/99NvWYqJ88ldcT8H85VyfiaktHGqywUM
1xnyGQbxrgbLjd2u03bVrNYCaGHitM9EjXeK0nSokyR5hv4GWl6IHBPONcEiNU4p
8htQDGE9w1pJaI6lk1AwdwssMT/jS+99d3D7cmdcf++X1r4RqRITfOOvF3JDg4PD
S+6qb//No3RAF2CFmmq4c8DOaRD1toRBjdrDqw/BarY7mGDSHtKc5mm2knBuDAVN
sLCVFTGuPRotsohmvyOkX7/o5sAFBvg1bUvmhkxbwVtxZhL1T/MGIlPUKcq6kwVQ
ToWk2mtrWSdw0Ep3cYmPZ+sx4AgXHfYtM0uZHf6xMBfKlO95jXZpVm/M+GfwMH0L
K4VI0fXIXJG3iusHFW9RdcRUUSmFqVwfigMS1Dj0MeWqwZHQCRYbeIGnJIM5JcBi
4GT1OcFrJXIFUsitMcVytGK2HKkMm43mAKJYzmzeMaDB6mtZqqtaKNx4sE7sdWyu
vQNB/oMIvtvjLZ5W/QtCUl6AHUiCXEvysKuZCOYkuTi56MEQQ3A3gY9Ptc50jfLf
E9gqMACuZnBaSmr7Zzrk7I1MntuyM3tPgVE9wWs3i/oV3K3oUmrN3uVeUVsxE/NR
PHr8/GoE00crXQKP6vTlS0bboj8sTQS8jtt2YpnrRXigNMrhEqLyDNXwGrDYDWWY
W96Si7Fu7nrsYIZxFacxfGXGlIAUkcjSm0RVUyRwg9XUcXT7e6DxCfQIcAptpicQ
FGvCCO3ym3Q8gTH7nniKb0v6Luwx1YmzPTltikC3jylKl8IgE7bU0OZWdcWFz68k
nZxrlUJjWB7Tv3GBbc3hgT9FQGwtI1bBxdS77fu6bjsmrCkBI/AkNcNCEwMIYlOa
Vxe3pJmC6vnJ4ajk+rqeKVnPB98k914LFaSdlEobzCmKWKVCyNOsPdPidx+Fvb36
XqveJJ15cxscYnTZLG1EavLHlahevcn8jKws1FWYXUByNHOBH3/VbxBzHWtKFbCr
7O5PM5PvF7M6dho28A2rkvgj3O2J+WBu3vYrj6MmCpHKrV+QKisqx8sbUebIvlV0
KDuiVuyBUDxAhDqKWESXJKq7qwGjlVAKerFYy6vXx/6GW5MEsUJhtCPDftdNDyHH
DkjhMG3WMiLImwDnhJqs5NuxISGX+kjqbvtTTI3KEEn7JsipFS2T1DLd/C+l6QBL
Kg4yknY+NZA6qYQaLixg+2ggxHWuiMmE6yDFIxu8LwOa+gxSGm2Lo5+Y5aiSx7R4
KayicGTv4wdRrIpezRPQ52IVORVHTgpzFiUt2Q8DFZ6eyCrZSVOBqoEh0zhXAHGc
hBXEQGHjnf0Y6q1MvpaNGR+WfIEbWtY7L3WfKsClvHnP8nIs2fbBBJ54bz4sSLs/
dTzw6UvFg4uOEjb8/YJ+iqH19+37ImEaAbkd6cARk5Lee8U2olPZKhGz0KJ6eUgo
UBV5XcFKLefpoKHh+vwkPZzCgcBGEh0aunk1Cgc8xkpf3UmAMNLNSoEke3T5JHJm
epTGVvg20fDRjuJd2VQ9DS9p7hIqncFm3YprAQCLlCdBwKeyOfG45wfRBHe0/Tle
dUkxXHwc4r6xwMocTwQem8MEaf+mYAer0BUSjUUp4XVjK+TZyslULwXNLFkBF8vT
IiAzocvwPoLRU6az4SShtrg7oYviac0xqLebvUyMOj5xbrann7giTTE7QcyxkF6l
SLYlGfI2KDp/fJD9J7akUbeds8NPl+w3RrUKOz7j9mBx4IlbzUT7DY9vMfqwBhAf
YKPqCpomVg7Y2oOaEk70+y+Zt86uXkKI+keYG+MZGP8IpzctqHAxoqP92l/lSl2i
7fjE/VCvfHAcrg004yCxMqB7rozMr0GhlE1bjBeah3HRwlxo5Lxa7csqlAEesdqq
92tnDoGPdSvJX8vTysCJqKWw3ec6lB0QrOQ/YnwvZCSAqDoilETAgVuKRe4mf4kD
dYOuViDkg66iMUsr8olT76DhYhXVnl6YFhpPbGJpPM/+9fM53RiEdvu7gwWsJcSX
bbTIruMrFNJsYyp5rPqOzYRKu2o39SbRR7OPyNLidvxS+CjiGjBLETg7LN5KQpXW
o5ewyQh9klRfh4jriWftZmerq/72fwK7HBbm37baN/ND5lUKPd8t2e1zxNKR2Byf
LYGtpzXwwEGR2GATR+x2Z3XMKYPYzQ79sVIxEykUqiH0r7qACKRGTeCC4BvSJNBw
LnummD0izxO2ArAjb/MQYP7N9FW19+QSm4remZS9wIytXBzxsdNtb9+/2u+sXiKc
Kj7UOflu1O8OsKwRcMpsrtS/0lTHL7h5K0a/eGYYyIWqHpDXnAXd4AkOhZJyvjOe
N/qCdcna4LpW3fa5p5HsVBTRd3CpeljrSFo5dCB9AVUImHxK/FbWK3jV2RJ3gj7p
qHpI+NDSbMJnf7KnH4Fx22A0yTOaXtbTw/YLJrn73Ml2PriO8GIQswWDINbP0cmD
05DCf+2QpwwFhXe6Su/82TN3fLUuT8T0okmRU79efhwiYh/xA0gT9UU0JWiyAMis
OvfsrdULJJg1o4yOvRvQJaAs5lMsHjUTwETEzmYh99kCeaItI2QoTI4sIc9mehyx
Dd2D4JcfGjkiviMrNLXszCv+/f1TgNulKD+eHZtao30aNsUfekyiwksx3nSJOgqO
wD0aLWEM+cT9cIcECbBfWeCoEwjh0ZoIukY6qG82iRjxLH7BaU/71aNEAYSVB9LE
Rib/xOOSkV+vKADT4joICRaeBj+jOhjdUa/VePdPME3CqSr+DT8acGTWsAcExuQQ
awVdDmic63U4DvITe7hfEr2bE3PL8/Xumc03aoFrjomrXcxiEIGPyfp4BfRiBwe4
Twl6yTONezQ+qDwYMCRHe/8IlQYxzB96YCiM8BFVfTjQTA/bip92XPzwYMR9KUFj
X+ve0gI2ptDcNolvt/mc3hhLqbzPUNZpqA+UX0AvlHfuEcHGrU0CzHgr8rtCC3MJ
UjRF5liGawqBh8+bvOmrVvftOmShbWkiFxrBJ1lKsjf8aRSKrO+PYFwEJplu38j5
jERwLNlpp3bVD5pHGOL7d0RTOQUz59gL3gp2oTLsiglVIr8DLJPKyOc+37UAxkOT
iAn4TKvIimajjcKDA1dFxsnq30TH/chyTHJZIeCWUYnTUmSpyhIjah3ovpSQWBP8
XKgLENkvqObzsICBJOCPJN7YbC3xt4FKW+KM1xjBuwRmpWQHBMZKQ0D8cDz6UCFp
sQaRjVExHRXQjb599Eo3vPlSlQGwx4gJ8HtEZzjcVWGSKeTR4wYK5T+xMMTsOPEb
QUpfNgbtSMr7FTbqKa6TSvUyxoPvzBU4PeVu7eq38b36XneOF+qihim8yW1Irz0a
IofGJ05hOSXf/qRvbJzXsWlkWbuM9EpGnuJTBQeJEs1OAmNv9lX0QccOIIbnCKi7
ojRnqP9evWH1vF9rpdTN4oI+A7vd/IC1QGgGxdN8+/Gq0LhuUqFQQC2bTc2aC3FB
+fFLD8lY8ihlL1xHjbBgBFH+VPIkUOPUrlZLHm8eoTUAbNg7Fqko6fL0kn9JTioC
cmcA1vIJHPTBhlEi2s/mBlJWOHqisP94E/e4tGPwZ2l0BudHj+bSXxc1wLjXUohS
L6ywVZ22T0rrlfMIEj2zk+lTOBs/1UNX7yq8X3/pbs9oY351wNasCsclbNQINUSQ
H0ro0pCihPDkHDgNOrrnoC6sWxQ+KuFJrrNxG7QvF9vwC39OfxsZjdNklizXddie
qaig6U8oFQOC4ztHSC14qAevcsDhbKEkifCKVklIYNcopkbNvIjmIn/pC+0Ecocx
HaJLGEMO6oh0InYUfQozRWYTqXZfNqs8MobDv2gDywr6iCt+W8zD2xX+cyDl2aDW
yZI+OHclZ8lenmO+ORvTVfww+Fgn//OUyIGdF4GFKeIZPgvHm9YWnSBqnflvMiZR
aTQl7Wp7kXb4XWjEiLuPlXOGnHq8g23fOOCc8gzdtg4RRLRYPe7cQFwXaWFY41KH
w52yAkbRc1aqWk3mmULg/VJ+56HiNzOUEXfxdvba0g9fxbwnn0ufaBWbly10A5VG
5g3NtqkVOBXIVEWRyWiMlp5aAGzE451uiZB6TGfAQjbKVBFz5wpZ1ImPrKdz5LmE
zQOQpypVRdSjMUHVMLcreZncxrnK41jSKWo93caWZyIMDjoe1absNjBDSrln1ata
MDnf9whlWaj+e01AYIqTgHgyhIXIl+dfvUZUlkW0dgk1fgTJDcKFKkkRMIUMy6Py
kcJ//J+Kwh4BrBAs0mb0x+EIpLnu0u4KQLKk7xZXDhSxSZK1jbfDU+RlQf6UCEuw
YkhmhWD9u5R7mIRJhYyCL9eA92LLcRdMA57Gkjt4c1f83LsuL/itosW1OyEi1hmR
SuhwQtiVUuiZ3Kys92BfK76ywIsCVgPr2HHq7QfBQNV6LbXLJja0XB77xUftdmI0
Wsir9tY8I1A9pteVf2ukZveEJl9EUEU4cuMB4AtkLJ5W8IgxPs33qa4scZ80Qczi
wKJJrJw3EvXGYdvVECFw0ZnZAWhkan/2AIUUBoj/G4tTy1DDCsXBPh/XBso87rDy
AyPmivhfRb6cXK0e4M6hWskGf5+a3nUmYncKNEOsQoWBgjR2wuFd6juODgX5tepO
/VYrTvC2C/IrWHDAifHax8lvYT+O+GBp6yawJZQcCsqTnqfBbEV6KvEr7kmtzOQH
SxvZNJ7M1M/Gx2jocVI2mwdFm3RmLKR+T1tLVa8ixTtVXW2j5d8YT6b4HGcQgACL
gIrBB1OPXnLiJWtlV92Sx0wezq6i8hH4UKrDKPdd6Ea0ofJz9trwExA6Vzb1GXui
JjrjMZ6pINjfkXBTxXGYn39KVBljTuzRbOUuqy3OI5lBHO2y/b1ZZhYyKSN4ZOwd
ShQYOI4T2kDG6L1KPqYo5qOwyCVc96QwE125zpA/zt5O/vjBBqbCCM1rskeuJYkA
ndrZlfDUU8gvKJ74v1MBLnhpH2xUXhJDfroav7c93QhilXJLZtHynhUSXBcjJIPu
Z0oa1MdJ2sHzslM9udc0O6sBWWVM/BB4tqE6CS7okgpvo3zXandY/NJE/sKWpD4R
tQjogUI1eE1y9OeXKd8afKCjkYFhObbpmIq2EIAufCWgvhCph94v+CCn/NTGnk1o
L0N2BpL2j9VqisHuVk8UlC9FOAUP/D3SwZWqmJE1VklXRrT8bYnPEiP/a5q33k/e
4RYkLh5MIGka2zgb5iFT2EuN1TOXjA6QX11Udw0EbfLe1VTuGltw1t6Z73y/FEFf
RzsP/qG8nksKaiwP1pv6GFLtA3vagazehHaFErFzx26JVvmjvksXUxE7taWQJsXm
T9ZT8S24tLbjFSX+F13pN7ifYHUtPB86+RK5bnuCt6Xv/is2JR8UUYIRT+Gf6gl+
OH27nJzz3UzjoRa0CLhPxLGJ4rrZQx4S3tjHtneavfWQh3xb/zLBw3hkQZWa89mJ
MkkbgEyWsZpTyj/cDDan3dTyuTOdzL0qxkGFCvysdZZjqZKHeHfMVsZFHB9dhzPy
/thxmwVg9f8XFDzBXPXTkDcM93MfsA6Xec4E7pxBbQTP0+o2lhk3Q5pZKplmON9a
1fq+/IYvI3ycep3I4fx8413LTDM4srhrUNWIBuwITO5vO8lfmqXnvsM2tI+2aq33
t8cfpt9NWKns/TAYqbSTJoIDqbka60pmrUKb8uIjpRakcmN4cfskkGJRiZZ/H2mN
zZrSSe8GFYkI3Ft2y5KJWdJHlO95OJmCixqbDsqnNpKOHbV/0Pp2Sl+IkT+v69m8
wLN1/hpUI86qQUTWVsNK8Ar1Mddani+dfZlxc93aRWG5VVbF8pYzFzQOCpG6JgId
+diFvIXqjiL1FSfwLZRPH65Gn0Fe94aohXaP+g9ikntppY3sQZcNBREkR62RCTuA
5e9MNJ5HtlcPvJtf+fvIJFI6aXxuPKR9z7r10y+BHkoBPV4y2lZlE2O3vAu0ByU7
ELmgje3FB2zgcqT9K9f8FW72PlwyF6XPgJWj27Ew7djB0gsAnCpw9ND01uU9GT1V
d0DppoooWJ2Jn9A8Vhw4OKGUkWeeBkWdFV3qBffw0EjSpYz6YZTgWG/XgtbFHlmV
IRCS+NGNHLiq/yn9rZdfFvwAylWtiTYjVvnpZNG/oAkpPMO4biVdDOY0Zh6ahvdk
dH4wNuTz6VYfWOID3P/DYvIEXnaYps8Ktn3fOhFgrvNtOFiRbXADyhb299naOuxH
VEcYb7b9NjXveHBtf9HS8e3QIQ17fYVY1JQaw4/FP2qujj9D9K4/0taebjRTdPzp
oua2IOdfkGbiW/CcDjEL6jpteFWRku3hgEATwXIFMg+NHXJ88v6AM5cGIPopwuxq
Px/Rbs+NIaH1h5KbJx0t4VbZ/3dF89Uw+D1a/KUUQviIVDhwCnCxEG5S5GQohH7/
LCtm1Uv4b+crResMVmDQHAdQj/SBKpfPnI14CsCB76pFhLNWMWz7767iFB99j/hd
y8F7t26Nze56qou+37mT3KCP3rXj9ejmpOw1iCeoxQGH5LLHvAss+XM/QmUOWZHI
wWhOY46nEJqNkwIqN0U3cNyI4pERODnd10JKhEocWKcRl3vB4N1WS1W93VyMOkaV
xnIqMMEe6BfxzjwpbPT5sLjkf36xTZnHqdOe+R0OKfp5g1Hz+8NWfi4amTKiKQ1N
wkNpznrc5DGGb3cCCQMRx83V2M33OZqpKboLmLIql5yNjadKJH3tvoAJYHS28vrG
Dl0l9X6WYDyXvYJ5J2nHU6LmzM87igpMMP/cRw4RporbkEHU9sL2PCTPvzQh4S85
LGyohoe0RsL1wsGtUlVNHJg6rWLD7dYkOQI0Ouoszt06tzOHIyhebiBxWPjxo/9I
N0PMMALIh4NTPNA0U6S1XW6xBWORQYFMXsN4a5jF0Pu2zqwRk1fDGq/tEma+U+ze
NtvqY9kz05Mu8DVdvRSck7zE2W42VYsSrDsgcZN7vtxKSYf0bMpOSMW0J03d9rnB
56tdzH7QGim9r3NHl7O9gMjOBZldLL+reavUzF6Cmrf92pvTSil7hx/0Cf/m3VLT
eulmtP99m23Pesq7T/PJHq4KCwCKr3UXrieh0HlVOjRyI97UHMoq5xZJ4O+6IUyc
JGdmTrjvjchgroVNISpFb0t+RaSEr7AgHkC44eW3nypcKFzlT2kgecfKq7rWJsRs
eF0QDg+O39auiOKSx/RwnEu2SUo11ObK8DUrzNRFRpTymSsQEEqbIDrQBplD46RV
RdnsSzubeT8WCeDrcPDll9MXfMJnIjy4kpUoxkbpKqqZukE98O/hhJmt4+De2btO
cBdWxHOmDeP3C5y9FKoEy6a4yfKk9KP+KYiXQMjdGphvFVq5GbQMOlKyvOlc5LMU
sM2//kNgXi7cPhjWzfo5CJdnvCFwnbmAqiHAUUSgZTEvkoE6sS/U3xxEiN633pBX
h3/GEq/BvQDZDulIwsG7uQiKfnO2Oc+mim1fNr/zpFVj+TZ6Au0tuxh3A+A7j8c3
87apAtYIAHho0wXe0IwBLg3DCaDrYDkuLNDMvNEv20C00nhLtHT2byCiv0zs3/pH
zp5Ivxg6/A93IoK/KFbbZJsAgRrmgtG/60T4aohDM3IW3zZIY8jQJ8UW9Fn9x2/4
XGnqhdVlKoizXIeZxiGdOl2tvTcJxHmeZQvOZRS0jmUR3i6p1ZIHvolPnAzk3yVC
RZAaIOsL10kUTy5crWagpeQink751glVjSIeHuFI9aBur3h3dqXlFNnIiaToSz+z
1mSJK/AKxXiK5RediIUS7sgff+GRip4uKFHHwmVS7MRyRnOYnsGtzNsz3IB2xOjw
K8kc9FjzbFhqM+ayw8McobtAo5/MFEd9RSoxGEhW343JvaG3xyJtXRlTcVlJRs6k
PLqEmzTTxY6BaPyttKzH1MpKx8/Oj2stgtp/Z4/JezEE9ijREUa6y2BReBHhO7Vp
FFNQoKSHCH2SQ3b4AM/2s5l+hzEmr+jH3nXGZVSJYB150vEd2uByrgDzMm5PjkRd
FVsql1e9D3fdQf/pOyJpPKoxrTlt7A2CLFdUmco1DzNToV+cPGnNGfml4Kz3Y+Tl
ASCWpA2AC1iHiCYcbZzOkFmgCny0mD9qrekeySBT6QRX3aEBtrcRKGifpwQn1zle
zfL2xgJ9xTJmUrdNDfIYUYn4wsI245IE+JnzSQC1H0wMn/zbe/5XlqLpnm5BDes5
DJFX++Paj6bQm4OWjJMdjhPgK9dePcWRjv1xNLsZWiP5TwZG+G1yGHg0I1KdlvTe
F8sQt6SByA0L7wlQxxxH6CYTsSCrBqnAI6DkOtOcUrM0D37i/X6+9ngQh2E1EqYv
u7qxgHoRAskHGNWJ2uL71KT8M7HWHTXDxROz7soKkw9gKNmp2w340zRoEFHdvClO
P8LuUDlOZJzQvJgbtNFTd1BoZa1mW9+2NcEjA45Lfu+NSTkQ69pCtxBYWwcwwn+p
XXmaEZv1fCtQxigitCMZqPhCHY2yzvugtX4yU+ItbF7M6ly1kF5PJnlcjmD3Ld35
86MAxyCHRt+LhfBqpIhqdktxaKeQMuwCh3C12tdBhOx0vCeMojrsOJQt4Eb6xCFZ
V/2jSWw7hXNbP0Ov4jLZuTRDbRFGxbi6Tm4kHSIK+MTGMNCmnDac182E8IiMNm1H
6UxwheCP3gX5w32NxDXJH+IDPUnagPKsViwwtbcG4slR058DhQ8Tq7dCDMHdGI9A
sV/NQ8BsKheebBfyqF9/dsvpjlRE29PPOLTCjkXa0CJNda5psb43ZALVmbURFqf4
Ca+xO1LKPV1UblicgC1s6Wb7WhvehnmN9FwpLrqup+NrS/dWOPGXdzK2iTJJ1/nL
nVhO/pEJwr07KuVQf0lVm38qkM56LchxQpSq1P40OG1vF913tuU5BpzHn+0PSgz7
rtnmS9fgPztnLTARr/Sarj0HJctD9GVfmeGZBV57PoWeFf0vbwzSAmy1znZcMjSd
FljK6FSZNVsvOQPjQQXFKZWqv5zVb3j43NicbX0ofyflBhDTj4YDukseosJaKLt4
xbYdGk9h2ui2OrGLQ6tboNUAghfKDzUBDpFr/Dy7vyZn8rhEqCtL/iSoHPitQu9I
83m8b9MPaka8lSR+51JABYYSK0QH5CgnE9i0CbSshonnabCCc6YMvwsyJA+um7e4
oR7fk/KoQ4KHUEr59MZsGBcO8rFmRY4Q2685GUJf/Nzb4URRa/W/JfLVKohX+IZW
RWLxBj7FaPsT8zeJKhuWrACM2mzegFD785i55uT4mODmprKzdRRWdPEoidSOTCAT
nqIy1NVx585dhn+sodeYF/l5gQtx7MavCvHa/I8s2QuRiVec+akIeIsMJhjdoaB+
mcsigskR5uCIFlbrEVv886+wWmvf/DjAAHcB9ICZSidyB5CfcWoampWGEuuXIYJz
GAgAzYjFOb6e8V9kkNp0X44ynooBu94rIsotG/QnZAqLgzfUiFhHCuP0Ok80tBVw
H0vJmvmgxPsYPFs05gc/WFid1ztzgh4kcIMGBYO8jlNkGzAQ7ShH1u1fVF8wpnj5
ZurbkxyZ0nx3xm6kNOOSyrEmDtTwcyCf/p2dyyCXMzcWJZ2gtZ0WK9nE920J15s3
QtX+e6B/YYL6i51LAUDs0hP3UmtMl+YEaZY8EmnTre1HFSwGcGofy8kekt4FDw0V
EAHOnUhQjNTERVfAGuilLAZNfDOK0qGl+YLZdw0utBcJtQZLO6A2owor39creV0Q
D2ENhZBD0IPPbv6KUm0Itpsn0RkcC9AelV07YtGe+EzT9kykeNU+Gd49/qutTlyV
w09GpCCb7eZqe4VydMb4Yu2ZR+30sX2eZUF0npGYKS5XcVi9piRVXTWRNiKvc7Z4
cDxeREiAIcyA8+/Q+G9DVIrUk5ZfuUHdUvg3Bz9SLSslUVwlVi3s8eu8eU6Z3Gg0
Pf2kzb2br5zTAUY1VBMgO46GaPj4sEsNHdgLhpWmQo9eqUIHweOwqi2Lpi7mmgF7
0sdA2O/syvNHkP8jj5EAvOs/G7ueC0aC8600gazy1zyqK/DweMPyRMHYCaUWZY0C
hyXaorz/znDHUIhL6pQGDktiTh4uVukcNLmXsaLhrqkZKVdnLMCrHoD0GlQkKLA8
4qt245jYPYBBhjxBu5443A+4ybhzFB4jJ2ioYNabJzRDdqwa5zYpLfSrKBiWaSyo
78srYXGJKwCSAgoSgfoZ6vsvIg8k6V9JZp7AHFu7fK9WDEpUwS2y9ojPz4uNH6VF
gKRecFN9jHuERQcQk0xJleoaewcUKJ5aN+XyoJf+P43tlGBQNiN/+fZ3BoqX1rYI
VgjvVnuisPcwPyHy99JmXLboTWH4eUXOzy9LVCu+d53fLlsIFsPXSfU1mEuZ+BCV
cVMi1RT8X1+7+5s1uFlpPfTinuMEx0Lz2j+ZHTNyl5UaCUvr02FCjMK7sv/ydMlf
8FHkUFDPV6vgl01aCa1L2slBG1oRs7GiuW+VCtoRvguJ/v9gv26Z3xX4BuD0NDhv
FzXf6YuY7iunIYkNxJVrPPX4KN0PzfynjP6M6uMJwshylase+UKeavCx1pjwXvCS
UsBNkYvGBUqWXpopAymZnY8DkHxCbn8RgIxcP2Sa3rsCCG2TlPLXtnAC7cho08V6
7Hn1bvRM9wWdx5BmvQql91kKxUs/FZwqW5CnkbRAj4HyzgAD1Ry6Bf0PkqEf/eui
q6p7sQmCZdNzPECLrjUd1cfUnpRbQi+UdvgVAcSBVuh0ioxhHw23YOxC/HXqYInQ
z3KnDS8kPONoeDicquJIdzSzbvKcIj5eyE77hr/39IiHphOIIYchvLQdz6fdOBqy
6MVJQOUpJdtca6FPlqR6QBAoDrvd4lEIjwKyIFPqJHx6XQOL+Y8aa7ai636EG2u0
WgnbWxzpDPYrJ9pRyNuol8B0YSvUgDxNEIzHzjh9A1LAdvJxkHm++0qXa7fnPuok
gd0g+3W6A4fAKKQLn+GP6Z21x4t2bhNheG/RJ4jxT3BKgyzVvvKRsM8zB0nuaDXZ
42WTc4ubiQ70ughuZRxZs0Cm3kP+wEEChpK4PaeDkCUqKzqfOPRZ9raz8w+8AcrC
rjAWRkvk+Fn6NeQpGTjg0nLYGpHmimuGgzj/cego+zZhHZ5uSite91bXrnjxgqbN
/EtDy1Pd1RtOOHG/dK9ZwGtbr8apgHVrl/MkTUlrjj70hYeZZ/b8sfL+IsUHMrIs
Kq3uYRKdR7evf3kxwGeqh8ysie9NpRk2f0cmltN6gU8ZW4hMtETXpGlS37y2gX4X
ScJHAq6svfImc0kEBGQI0CvTnImnpXsNd44xzZeqmIyhb6cenG5yJ66uB9Wm97CW
C9PeQE+QmTMkKvSmNIwVf7SILcL8GYbAhCluKvd1DTyWdIa3F0yB4whn1G0gz/QN
m4Szl5kyd9kP8gK3j2Owk1gY4M1LKdD3vDtQ4wkZQPX4W25ElRK5Nc0J40jwxwfM
yr/KOYYGtZhzhYoCcAsyyQLQdP998M5C6Ws56hiKFqKb8lF4slJAQr2DaUn2qFRK
oH/OM9R3V9zKIeKajuSEj/GH4PO3EyfBlX8RKkegbPchqxoieV8E3ioPf2bAHKlM
l3mgU0kKx/J4PE58NHsCEL+X/ml3tcGEURe4KDPBSrKF6UdeKR55FBxtG2uYCWZo
LFY4/1HW/lBMwYZlv96R4Gom2uEgebg2KOoqeviEafbXRyHTLM22QL7oK5AbiYib
lTzBubDes7JfRuEG4jefXGrXmEZ6ZSJzj8dNk1Vl1TsLfzpuHA3znGKs9Wgwf5HY
VyEUk1YgPZlIDmi/+WbXH7zD5R46MqqzxyyJwqlXSxbYk/o7107u6Mfnp1+WtgOK
szo3KJE6q6Aj89OLupwy9PH5j5DgC5Phrd+urPbXBqydTlY4cL4ZvLzOBg15/3Mi
t25uar+zGQDKUd2I5q0gJT4VAEjxR9ClzvKkvAf2gpWgLBnthaX+eM6vBkR7nwxg
9jPhQoSYE5M/6Cs7m063LE4WVhO7Ph7utv6kT94v5euzzyvBJA+OjmbXtAGXwcIF
lXsH8o3GZ6r/oYeSXbid0oVmZvv5BwVdIfNNRkGfDwXlj441Q3zONp2mhoJ0Vh/U
V3uBBNeZqr5wFtCnN/7wA99jtd48cFGc9h5/ypMWT07m2lmV4v83ZzJBObdIdbgJ
HGqC+yT0UG76tD0xOpHAy5LBCWUZdi5KAwwC6M3VijsR4bik0iAPQdfpRz/ZLPQI
4AFLNrsCV5JGzNfQM9y9dpj5LaVS72vua/hq1z/ipd8NmDrRNMs3vAOVq3zJVNvp
0cV9T2htBTdt5ZLqocoSVAFZ4FA/iGn6SE4DANBBxEK4f2vrtYq1xENCxqIQoQwr
LfPMx7WgHeuVArIfRE2ArXFQrpXN19/Ue7IzHT1faqcNaKKfn+iu+dou58kecYER
s0IovXMCKoAkYDEpjkiXR+hgsi9cj1UTyhacGI39fhelibYoFLEAbpT7QZsZDjJz
m+pK9NILjWt5Uxow7vYpcI1az1fJsYfEABlVFOp7e05UrbN1vB6SiFsBdl/RFgai
XVaz1M33UJQHyMy2UvRihkE0w+wNsSgv8/p6LO/XX6piReMr8CS/c9fo2LSf6g11
2IjENS+EqXIWjQTcWt9ivQBMf+2qcQtBmYld/q3ICsctcfr2nf9w15GXtApqA0WH
8T3gpQ1bNUHUiSORYKnF4f0T2V5/CbwHNQyzDh9ccjPActDaLbtnWQ0olYGWy4tK
bLiGKl7lECpHJf91V7OpZcwRwxUeYWculGX50P8J2DkvL5QKxlESe/EKpC/8T4IE
Eef8d0MkxRYi8z83VkZ3qmCjOb5Ug2Ox/yt2INUTWKBMMJeW1Bzcll55zjzlD4eh
8XMajfkS6DLYzHoPQNSWyHnJIhIQxv6m8CilbFE3LpH4FPoTBIHbT/6Gu67amAaZ
sRaH/CEZi53oTzF74OM9u2OUlCtMBsklOwlk3L/pIM964x9giR0uCXzug/85KjzO
c2jg2QHFqnf0ZsFpsw9XTPoYqvFq4JE2+KNbcn3GoxhZFCT3qhef+LrbF7yYC9Hz
JK1zYgOP23yJ7EfqmIVHlkkSHn6d2W6nwClrm2VpC9LbZevqY7bO77OTqj8nl2nf
lIax146y2ukz/1cyh2WXOo6kb05utY6j548TBUEexBcoS7JlVcLZ+SVDFgAmbOGF
C4mPiclmm45EwjI6VSP/eAH3mIgivQR2azF1t4J23emScE84cS2IfFFjlGsp92Cz
EzZa41015fURhC5uNr2qhZKXRnrqdKH5dRTVeYn+AMjJ/LrCu96B1HWWMiOJf+5p
qmOxKhdCG9axm0s7urAlU5xluDF4Zp3LgGuo1oUg7QDJOYYE45I6rq/NAGE8eFtL
FtisGDSNbQRDNJ97x9NZ5etNcb9nBVEiKQhAPm6SubhJnhk3jNvPd6rNt9OVHv6s
UKG4yiAC3LNlalNGdcInZ1RPNBuzdelpWHNk6g2HpaB7OIdr0VNF5LRiMEAN0br8
+elUp8daqsNvbQxCNXEO2n23fBSgRJi+GOliP4+AUk/zJL/aZWfFJSaXNXup4zed
uuCnq2VPnCoeslyGfGTwcGZSCevTC5fvG8E2SF+bEKK0t+zU5NGolma8bSPsiSqg
Mp4TYf25Bi9oXsD7absmExOsSg88ZofHMsojCMLDXCICnipvz4ViO8GQSPVAz0go
fV2MtxzWStQ3gMSRRO5VDUB/qX28v7LekbfQXaDa100G1okjBMgtR1+QOgnIoBPv
0u7DKfDVmY2+/Hu836MAnt2ip3y9GT9o7kVX2qkTd5S0Yu3laJ1Kz6kZ45HuLzjz
kDlJlqvk35ytFwG9VdEH/SaTNYhyKP/M2DK4rQHkHCFBAn/uicCVsv3ubNT2oAPc
PNig5wqf8IsXn8XYBBWeCQhJZ0CWaEu2bv33qk3y56W+OJiJb4VZfOwRwLlmC0je
j9JWR0BDsVG+sOOGJTNp91j/vFr0CQfXHf1KlnzLb7J41AT3NekquOEeVHKxdjBK
2hV1WUKkhzY01boVebb8ouKt0CSOHc2W0V/PEeuwAmFlqBNmU2Cw27NCuONaZb13
9TAObmKY+sDnCkdjsfGvDzADxxEfMu3Q/xFUyXOxNGhA2iAV+zDHc1EB1TfQVXSx
8VUrDrN9Jo/IUKE+JI9aCAWRZcctF2kpU74oHDKM5eP9342Ow7171mgCoOoJD6GI
eDNwespz4MlU07C9h5kW1bU17WFKADT1m/61IJtx0BRxJcACM1MRw4oklgaPQalL
X1UwipSQEFtJiKPZpuNUGGE60G0cn0fiOTLvGygINI3w/fGdOtPk/8f+7Pj+6+JB
IIsEUHh+6dAgAZTvpi5F0N5DEX2679hi2JuG7sr9c2w5bjgMDEF9eRPZ6M8L7Erh
jAYAaRHp3m5Gj6nYLHjBB4EkbxtMEaboTRHFwrJsyYh9kF/Epztl76EmHbuR1up7
6gQr2piL/jucTXodmgyAqvyZ8xbGF0s0S7JcjWOoedfU8YJ4D38A89ucAhx4Rfhn
Oxz72c4x9dFMykeuvOzP7CNRNsM7MFWik3i6sAmEPR9U5BKvh/rcW+ej5Md7vdBW
BhkuKO3aAn8tLFfm2Tn6gGTiP4RZnmwlka/lOrJiO5g0Q2rncwRw1rXaQct7GRMC
7Wl3YgIZr3cLTZDnRbVC1JmcJ47E6ckg4dYPkUllEwD4FqiG5lk/MRB1vxP3Jnwk
5Y8bf20HQyT8SFZSgFUCC1usuR/uH3iFiZ1Gcwe3iYNkmGUq9bRWYP+1ngnb3mUP
xXM47vbIMEgg0LJ2kE2g5kfsiej/n8U9Yjo8qBLLexY7UN39SqHJvT1o+8PD+zSC
RvnDpHmnceFi8+GYfe1Q+oxnKJQLGsZB6tuHQUaGVm+rrBHBvFFWv/5Msy7FgFbf
4HjkxGo5VL3VudXw8XGBbc1uYYbUCirSHI7HVKtXwsC8FL74QmgjF9dTglLi5sdQ
gcFh0O/Vpp30MUXRigGWBottq05VU1HcvnALlvlUY4Y0Txnb586bpP/lJS2X4E25
r3o0vKIMrLl6Ru077FVdOKFEumCqqF+vft8rHvPywNQHUKr35cCVDpihMwtJKknZ
4VkrCgk+V/gsFq8BwvTCcvK2EwEnrW9Pxj9viijyzH/83HatEHVYUUZIGTtDpPRI
sUnijx4pN54e0PlGsjgpeMUmyjsHZ7zPfUvTX4efzGr90wTtcIBXmGcy1k2CKYM0
28qBs3ucJOfZ7lGjF3qXiY/qrEWgTQETB+QjKLM/lnHVF3ko1DAFvZV+aA05qfc8
j7cwqbrNAFNNwwZuxMWMs6n7l6of6Jd+67v7Pl6naJP8kS+HcwBzT9Z+bIpCaGWg
Zo54+LyQl/C3c5/AoJt3RAH1Zl01cMLneBO8KHBMUFPlbEhsXiT1QG5gUAoT6KzY
SSWbL+T0kujc1ogZ1nHWzaQupPRwQFSSq86VEXFHFdqenF6W7VEIqJ/RMjQrLDeU
bv6UTGGqdHjZuV+itHPW973NlqY1vCMyc8Me6XCDt5fCwWZl2CTCzX5ZpLUD0jub
GAezQ+CbWmrm9TBtwZyGQNGN7gO0XH2eO0HpJFlb9d3O5ccadLE9lvWQw3vowgpK
6FhZflbE3YfNwQWL1LCKGhGRzWTZZ2EVDv8ayT8T9tW7BLbXJHohSf2Q2UQy4nwb
DDLkx3KlzaciRoFzClGlGw3iJNnnHz9N0boNJUfPD+prtitmmPWqhXtUn9Y3TTe4
zVcmgGBl1Kx/qyO24IX26VItAbrRdu43NB6rsoqRdFFBioxapvbC7nRog7uPbvcJ
RpsoSYbVFqpcWIIwMyjv/iwUtClhXMdU/iUdP983fOij9KG0dcilyYD/Ivc+Ut0N
2XZwFj8Pjjxz8yiAtp1AUogHXzs8fz4Z3qVbzm6PvqeLP3lz3QTY7cHN8+cg6mvP
V/9LeBTdZf9iN/Th45i450adKaBqmfWkYFFIU1DZZuAgS76aAbGaNS7ulGLqEKZu
dp7+5uXhYMuzasyHLmqrY9jluaz3K9KkPtQT+LBFZgMt6RdEtMJRo+JHqnUBsH+3
TQvswDjqQP2n4c9lo8SXKQdHvCcYTA0GRNjf0gPPPNBi4Ra2P6QLF4OFiylS3asW
gZCNAncP3xcKVgtylqU4OmYpn/W3uEEq1QoZEEkbxNwSAVYHtWrykd0fcacXZjVX
o4IAWj+M/AZHy5Ivc8YqYvpm2nLnRi6s/4TDdEXc2/fFP07kbhdEC4mC9G9sgZwn
NTaJ4x2Q6nIjbKMiA2Gr3NcpRGBOFbUaC462/TZ/ZjW880USRH0CfyHcTwenGtgZ
iOEkIXlrU7o0O+aOZjZAeyc1iGise49bh2FA/IuDSBJ+mR+t3yfaiC+d+3bV4oCT
yoh/Jnr7/AjGe1gGwUnDvmD5VgXKGZWTLqzWxfaQT7JY1AwwScDOB6976PhmCGH8
+d7qRI7vOGCZ79H5/B+QEqKJN5T0p6y+XAWFNudP/zukUK3XoOkUfvQeWW3uHjfI
6bDRdifMQEde6yHX7cqX0Ek20GcvaMcPG3KAKT6L2puKouo9cjlv7IOrdGkX/8Nc
DhYOWbpJ94gFhHH+3zNFXXvz9AcBZgVVlUYtliszYr29FdsHM8hLotiCa/E70Yp4
gi6nd0ztLjJURCLva9d5YQ0DvYO73AGx1o81/wPsTHmOTO0df88eV1z2itfjMil/
IAEGb24NG+bL6fQkvlZH5LgObCxDj+8szGLq/ZbgUi5JyfZt0VkJs9mmG+Q5ttHq
fGEFkqUwI9108ih79IATkeq9A9iJBTvQf4Uy2xO4jgnqORYBW0O9DQveZa05c5dt
FlDG2+ftKZm57oBXNocTaAEEv8EXuDY9gIK/qmnN0W+AHG7JjxUYVPFV5a9xW/Z4
nB9uTQc15XbOlsdrjhIj3wL+HZfmxgI56Qm4SeXSNxARIU5sCV2MYl6MithwzEMj
lLFaVWvNASSRJtfzW3yLrrExOsEB5sfovNqVwgCkbXVohDHaq9wJd0v+Cyf0QERk
ffrN+jxbAF7VtrgGkQtIpCNln03P2TIuxl91ouJayVz15UgWdGvvbYlPhlaSf1qy
qzD1vlsExl9T8DkRIzR6adLNANMc7ceXNmXLkuR8W8mksiPsZWkHOjwVHrzgI64Y
lYtag+jpJergSZ35WR4tiZodZrsT8BYraY8wXFqZjTW7hWdPl1Hp1fPv73ZwiFFK
BQqiigRj4NwrcBZ+dUStH/0cgTMtwT9lRy7Bi4zQqcEVX0fyfEq6IffEFjntojl2
9L3Do3wnCKVC2Ir5mIr5H2GD6flurjzIdm4aPInxeFOJUum9EE6HlcaKVx+eIJ4a
yPS9XuSN2AVRZ+kEDQSQnI7fw64bcJw8LTyD3mOMDXBovEm3womixor7nB7lj+Kn
tHPNRc/qzkinL2KS4WX1W8Fkci/GCo66TaaHGOzf79Dv1RONEOjb42wSVihL2Yeg
4FhWgvBOCxRMpAtCx3GdCH09vWqAOQ4JwHkbx1BCYPYMp04v/AQGvUDqccrd/u/h
kP7OdUtbhdIUv5MG4Mrb52lgpVeQCKf4ackeKeEbmCmqpKqWzaXCXld7sUkoKwvD
mPtLntly35sM1GLugcmlKunNAhDdsLrtK5hkumb1Yg3LL+/3Apl2DMlaJFXSVlBF
B3uFFdemNKlwKJj54Y1ftuSt52QaWUwk2CS1r+xe6DYm9uVQZWSZphVCSDIWEuxQ
tMOah2QFLekdTqO0liFUvWiNV5mm8siwV+VsA+d/RypEO3pxpGkqmU077WJ9MkZn
JPvRDDYIW8jTAlAjhHaP7LL4q3TQrjI0rWCXvzdgqt6RkTpmZjypZ+3GercuKPzR
Rj4IEpqoeBDqwzpmoTncP8+EmU2zRRc6dU5Iwr1yO/3c+qKYLYsPGgJXzER8ORBG
3e9B1siZ9qCzcSJiuw/iDMgrmPqibFnvxT7htATZfB3lQJ4dJHScW7aa5XGrrMoG
CmvnnCGIECKng1TJDsrxkV91si4bgZ4qZeze4oZq1W1A1wL215rxbAU5bQwbI4+M
8VXjLDtMzCyZzGKNU4NzCApfTkA/0wpC/LKEpbTVyNLvXV9rEzcrf6qHw2X0lQzJ
+xeJQnJrHKS252sX6RcZOc1FF2mxhnJtVbXBrhYXtEwvZV4f1uLsks/sZzkLaErk
fnpdbGugoZ8s+w1KHqWaEnQEKu8dQcdlfN/5csgkwdhFDAFDkiiyOf2zYPD/WQl0
iUE075wJU+JMa5uUsvaZBn9WVKcTojhTHHra4Sb8udv2YcgrXyJGLle8/vNDPwJ7
3oEZgtxWyKnvPJEQdGQSuPFlWMS4OurOorOCit0OzvySw44m14pYfelAifu7PSjc
PKcn0Gd0MndfZpfnFBil6fjhCs5uyg7vIdZvkPrTyU91BcjHuYnHaXgu7KeXqFFF
SW85HN4TLVcALaMgw7mw3W4C0C2ZGRaO+FGMFlKy4qrtBsS07AH1iHwdp9y3blDJ
/VDrgMyxPviCzG70CzDZCDkc6uhCHH9kbNOvRrL02UQt3RAxQOSF8+3MV79ft7ZY
nfoLxLQdwYmUKEtCiEXHkN3cjTxRYgSMq4NRJyrxJW9PRbDU1kkpn26qPYADtTxA
qDhZgn5yLyY0MRsdRCrUCzYLr3Q69FXpEk2zmb5HGTp7/5idViFp4/CoqNiniLLH
G+xVz0sIICiec/sxZnir2wTgUGieptBzThyr1L9/WuZx+99wmeXviyh1o4eveX2S
A3glksG9+hJPBHjm+qSmUzq+3cNjT+VF7ZuYdVg8yOCjB/rbeGcRtZQP5YdcUCur
gkOIb/dMIVFZELyn3giV3aMOlts0rrq+TaL/H4DRnf0dhXxAU9h4RMALuzJ5kAkR
EVe7gvL35NCxufVCB9799nRfG/xMCdWcIZ3ZImZ1+VDPu7kiq014xd/cY8krRiL2
SxJqz4A+U/9s4j3gcZTEWSNI4TRUfMcVPF1rQ+N+X0Ed+nHe5MuwF9BUpJpRBC9U
r+1DL3X7OO3miQcPCZ0RzStP3cG2KDHYrLmkVpBu2KJth7eMhk5Gyj0ytT9JPVS5
2DDvpob/RdlIqmqFhpxkC8064OiW20CswUOY/JP/n91lZVWr0Tyaz75eM/9F525w
7OrI7kME+DzvrBJjsgti63ks7zJixxJTL6cS79MRABxbvibOHyaHIg4GHF9hCUro
adsiENDMSHUFyGLGtNfFzcgkuZuA6Pbz8UIFN1OiSbvPD0NeO2u3MOcEkjAeQ4og
5hBfW4KoXnjvnTkBDz6IbxRW/ATSYiwC/jTl3F58DEMOLhioep89gLB8hdYWGXtg
1lcwvF/sPUsyDNhAHzpMkPsWhXpGbZ3mhDMmTJVpd9wXaw7iaSllj63Xb7qGmg1j
CEZS5uxzfOpqQc725pBNwsIhNgXUy9Lts5B7nI0B7iiPrkyALZC96AewpeKjOzTL
IYNlUzP/3q2LhW7RtRhWEW3g0Pn34a0SfRMB7puysHF4ME+6WzHTJf/VbG5qTl/y
9NsvFRFCOJ+i6v3qYZTCJZNmgYAs4ADkWmmplWBlP34DrGJgc7JbH9h5vN2dDP9m
uRrM7CLH8FND5BxKXj5/gkdk3o9DJqB8RDy5oCxrHWHlyCc2W6Q4sAvxDuXEHyqd
EOQ1mqsqpJTkfjNmCrNDA+wuEseE9Chd8vLEr5lpjfasOHrDeBd3rx4KHjghiYyb
kyEwVK9Sd29tyEp37PpEtmflZ+KWyTL14AZPNyUW/+t9toOxQAtw6AcjQL2AvyEV
qI/uNMHje7ukgKmAmZ86ZfEwsuTZdhhVZqE/6ywq/bp4R5bFs7SsrHWxED61kcCJ
iYn7X1fCVhWBB8z2NxBBfBcq9UPIxRzgo3wh2nOxoj0d3y+HuaacaeF83FEG797z
1uTD/pA1ztvjXiufHz/OSKhqDkSYJURlxUpXN72K9lzK7AB1RodjxfXysIx5dmxc
hM+ER1iOnHJRzrn9EnuWQjXdF9INSlaJDx69OQLBYJJ1NluF71+cknYYUpw/uxEC
LvqzdjvOK8+LIu7gK85oJ7T4wE/Mz95hayxS4a2Ws6GrTjVeSV46gDwukL0K+d0B
J21h/szxpPYmHFImuUy1Y0G6Br48f4CqO+NhIbsLmN0LBj5upRrIwre0WCZKbl8U
D1t+KDpRsmKoAHohxHIAkWXjJvQwCu51T7drfXpOx13d6Z15ZkqvXiAf9ZLrOw6p
7QD6f5gcTI6xgf0EdBT2fENP7gcXaET29WmghtVF8HP1VvcxsGxTp6ABS2GpVy5q
LJM8vgU6r8Ehp+94cRF5cMnSizCbVC/oXQw5jn/OZHscQZL81AIT2taXtj6blp4c
iY+o6vFQPSutnD+eaFaNWIH0xfB287oqBDisle7kd4Tz+GmU+8oDBZKl8+F+XB6u
u0QaNKkfG0w39sM//pu54D7GOwFzAo1G0GFiSqmf6Z0pWVgxL1F/zJ3SQvZvmY2m
Czp/dRUns5vzaJy01fUKO3hAQZBJS/JHFdEk4CDkEZm8ps8q7F/uD0p8FOl5lDih
tVE0tq8H998/0HhP0PqEnVkRLzC3ZTYZVC/IClxDSOlHZGnwsYd6C/SBhZqwL82O
DuTFB8g2wbcNTquZBe6xpktN8ynG1OgDOw+MoCS0eoG+ok3KZS35DqkabBKtlQc4
W3L+2Fs5zdrI2DV3vuba7dUV+mkMf88zm9LkZEDRfjeHWLOqQX/lxtz3xJMQgWaa
nLWlxFeLRZQXex0+2UNwdFzf4R8lhKKQMcoh5PHTdNX/GhnmFyL1p9GPGeVQ05JN
7lJbu3CZfoBXTqQInC+aDpdLiO6CSTpy1YSIRl2E058JS1RzA3aGqmmmKte+CpCA
kg39tJv99I09aH+h2EDQNoXu3oq1Ay4uT0/nb93DJirQH3xPSBxDYteWR9EIBkAb
T1qWrZAZCbZvzzb+RHRQ0i5K5cDeUZIeoX5sN5ubwi/RLVFqHQXpTSSdgUCAMq+s
O3UiV8r+j22YV4H6r/4f7rhwqLvY9QmPntLr6Zgxfl/g2/FGYMwK8V1gAc5yf/pv
PsGgNgXRQIlHKEkbpn37wijAjNNL6koyxUZcyYeZ4qLwUuNe245ZYi3p6NAg0Xo6
FKQYLKlehYJ5oLIbPnak84SPiHXKbLWnHCUP4JGfkLEsoLOPpzsCScQWSwz9fyQg
lvFFpWjkl1Rc49Wb3kdDLgECrDNKPKzlaGoyfD3GvwLNehrmVZD77rP/r85ysgyf
C4LhM2a5MMhwgz6mj8Qw8QLqTeO7vBrEPhxC3cZ6cJAi3GZbQz8s5rb3SaRj+7eW
QjvXlX9JB3hjdjFeUTL/N4Jzv5TWCFAsx8lqtydj5Flibmj/Dn2l7K9xAx+ldR2W
1EhZDB6MHzoBuafR15MIIFhXVHvBlS4Ms0XV122WWf+5SMPneC+2q9IKnrIKZ1Cr
0PqZZfOlZAfqWncPK9lefFLA50XnkiflEaQPIM/efLYCt5zksdKP5EES51F4nXTg
wgSEHKuyZKF7nduZ8Gm+R2YMA+oc6mlRMZ6R7vwvtQsLH+gXTHQGsDbtbUZnE5G5
ZZeSSDRhCwG1UipYc986uB+MCTGKMExShfYj9TJjTNi9waoK002x79Ng8S/JY+9m
1/NlUXsxH0ry55NtdcU7C0sCKecPQujdS3uEheSnEyxm3H2GJP83zdNgHi8aktA9
gx2/luf8S/+ITRYbmcFNIRN2DXOfi94uRLuHMiRMlP36YBd1ULxYLuRtBko8nD6+
ynZ7pjsyEAUziRhzAWiTCJQ/Z4ARYsSBYmaSseCozk4j4AGw5L2zAqS7QDYdhjlp
ql8G7jXDE0K6OyTU1kxoqNTEQwweNIPiLYEsegRYdQmCvDgaE6hRDSFX61RqeH/t
UT0xmBeyo9O7iWi0bJqTWAAZ+D/s/9bpOtKnTpC1txzdEHLtgnJdbiFrGAkhZutO
5he2W+C1ehgh22C5B4VpsvFG5aiOL05X7iXlLVli9vvPM9eOGiwvfXi30ZV9sK5o
iDD55MdAV8XDcZYS3IM5ah6vG2mJE5hy2zBGHVJ6dLvd56r4aRiiIA9ZG5TskZ9G
PRW1Z52zbSyN6JZtALACW/OfVPvAt4EBPAelB7+gm6MfmC3roTl9SvincPgJdwaq
cvC9uDIyHjxbJxw6u1yho5ayd3Bft/0sGMh6yUwqNYxh8B+q53f2SAJcW2ugIrwQ
9CJHofv/OJyYnZ8mtWm0GCqXm/wZ/VBmk2RqgakpJiSt2s5XWmpRTm1sRzmYVUoC
W17prMRT9Hc5tFoC5L6atovu/J4FqOFkJCouRli/nz9p0ib4X6FHqakD2crfGeGE
abpBrdCL6BA2Qmr5swkhhv8EKqUPSEW8QNlDrj9njwDm/aU+qjPclOPcsey+afLh
1WfHYAAyIBpcbbwgq+ODVfE/NkYCkDYKhWUJ67omiXXaNq0GJVBFoxbBZqTsfkk2
nlB2hKCq5wEV2lmLQbSLESbtfxUJuT8p7I1NFS8cRnIiJh+Eiil9r3oy5tfEwGEi
hJlf25jD2e5nqmviWJIi0kcdZ5Id1FoSRTZev7GzmLuank4tdV1SZa6BJQo7T+Ku
pD8yfHnP/vlZVKBasMYOb7gJsJ3vVgY0tnaHn3hbKM5k6n7n0VmZvo3Nr1xL1Rey
+zOVnpd+BLhF9Va0tvK0+/sg24l0J2/3hJymAi/Ou3TqfNd2gl8jBg9XHrE1VgC7
+PbZduVZsAix36fGqMcSOgSV5J/N//WsQPuvNcGpst4SUVnTKh/nDNoZEtUNPkAa
BNMij93fJi51pkgwVL0RSKfuQHlWmn1akpEgL6jro5G0Mm7wwxdktY83gt5JUyJD
cJ+haFONaYNh7JhZVIWMuXpSMUY3sQDBXFvOHx2+RaTjqtMmwyxQYDSly3G0/WHM
5jFZY6NOh1dafNTAc5NShANAwQGHV2bYKGBo1jfZEZj2XX6Kd/iu/SpFBk/HV4+S
A/lTOrHbh5lN48tjAff12v2Tys4rrtI7F0605PRYTdCT/thsizKQ5d1wXCASi9I2
WSUGLnoCtOuZiM6c3rwUAN2Vbjkf6o7flj1CTkyarlb7fGP7ZmAtzDfiOtWX4kQb
hEzSCXrwMZUn0PUhNnhrL/1o6Dc+ZHpLCMmGNLaL7gQAAv5grMTx8mlPTx2dRXML
5tEdNULo6f6MwI43mplWLJROs3GtAp6Uu+LkWnqx94tYhS+DJACRsAjdYezI/iYG
lqqaTlm6DA9MPUtBmGGGq17raF8SO7NHxk0+2/+SHVYeERNTr17gF2Y5iqKv/N9x
iY7Yi88+hBVJX59LavP/AY+i5upsbmm+D1MkSVT0te8vFT+VUnHfWSfapTYLOlVr
5Djk4q87/Oq3Apcy1myd4Pgyfjtc1DCQRyo/1DmvAm6d8VUzT+umLSlQ5MYXeN8h
vVP1eMVGL5rCtWeF9vwkw9DZ3jcne+DszegosjgN4RyDYWoe6UuUnUuZHFH7bGL6
2PGB7WDOEzdJQM/mlE00RNVgpmnB72dm4QGGdW/+/op1MaIuxTKdTh+AoPYBM04N
VVRFtdhrXXoiJxwE1D2/MHXN9oJjBy5YK82vYRTEVSWGf0ohgnVHN1T9oKLNXqcu
JUjetCUkh81yuhuX0wRKyJL0gM/EqojrBYsICpMgA/p/S5GMJ4BoEYjnqTdKlSyx
ELx59QHXnYhz2pFlYY6ZT7XI2zqspECEkwCNz7B3EhzRoXnEAHp+oEFMAOWXeyBj
DLZexq5zIza6Vo5feVbDaFQ03+ZFX/hLNsc+t5CsmW1Tqm8jmGnsblreKt6qrYNM
ZoOIJp8klrh7QLw14KWaXlMppfIhDlf88dF7VoZlYihnnXFXBP0KyOuwLK2zCKAw
AON1+YYw79LYdnGrJaKhkTgN2ngvErenAnNTCXax6gOdiIL4p2GyA0iT9SWO0fey
CqFMDBvtmL8DnPEHOSpYzEhQQtrFibIcSBGBVlTeLC6hcvZwixUC78kXCopp3+WX
0qGxq9/S6zvKw/Q+rduU73lu/HOgB0n6cky7CZGUuRSXQvCSd/4cGUpGVp9dPRzz
WAysjYJTEyaO37TWvf/5tKEaBZLpvralZPsZzxkLzRU8F9fHmxUFl4IdIpvR7StD
mSanL1VpgK7tTwmzNuNHD1KoMZLBCLTaeHV6/MsbeWDLTZru1loMggtn4zQe+qif
DGzJtjXyq8Hb9L2tKGVXNFzYdeD/2roFwNwKhFl9+2iU0/S0WcPF9VBbkK04VqE3
Y0BUCV45j7blreSn659YNSPzfa5/2pX5xm+2sxD84qp7SsxJXoJx+f1RAT+Px/Bo
SaTCukejQ5UxGVbgaKv0uGfWd+8GPn3wdY+OlY0zYU/ityStdfEVyW97mf2PvisF
s7xZtcMx04APx4wIj8TsJBl2jyWmHKdh76sFKz8bd33qCFrPjWN8GD7WQR40P9Ep
wuDghwyXuss/GyAruNFdB8MKSfpEPfsJfsAQdhspWhwKloZ4ey1F8CqahjK/iyL3
5HbjY2j7EijG/mgKkALzrpuQzvLhWiEcvG1rvLnKrQBunmq4CHdY5bW3cUJpLVCG
rzpiORbuKqv9Ndgc8nb45p6XEnljYia0hVf3l56UA6WhxZ/72xzUXU3WMZ8CMlUs
mHbri774FYo21NR8RRiDKqkYLuvsCDzxyexSLewsWP5S0dnmGDvzEV/fRPrxv6Ed
LKvI10JqQ/zVo1ft9+i8umYIcF9aVzTO6cQXjEjlBwB4S1YNjF6rptKXL/413Z3s
2GKD+gWWN1787rG9b8MV3glI4NA9qbdMNxqMT5ejh4wzHxwnG7QoLOnDdzGxwRlt
QwYqT2sMS321Hz2c4smMzG+zvvWtopbId8DByS+O8kJJKd/yyjVk8AEb//4uKo1O
zbU7EQtPsK3C7jHzxPyKu1TnPZvgxvHxMyXDVOSh6evj+k3cP/linHy9vFhCCzSY
pfoTquz5QxwBcDUBu254Qb55cQguXdjj+FeBFvmyt1aAn39mAN+sPqg3MDipcLIE
ZCEe4NwBsq1ggDTWISdCbMbmsmqeJwqaiBRcUW+reLTVvn0Aqv+eaXPj1cmnYqlf
Jc4d+SUC1iMHCaErR69fc2UIeOO47rnKLbSUYLzbWuZUz54kYKWa89LBwdbMXOM1
54NMGGxyjsHE6yPs6AGiFP9ophrrNBO5tRfE5Vcb+mvc8V9+BSTE8HRG+KBffKxV
2zibvZjCUHTAgMt2OVvwZAHmUX+Ef1xaxEmyvPNv3uevF2nSe9epTudAVwW/Os17
n7ne/OX5l0YhadVDOARg8/1jcE8ueDNOqNfV4Wz83H9l6HMo7FADb+W4KZBmUxQb
rUZHR7ShK6lY9CdzwQYzYke3Yxks7P3dwDpFQJ3UXOoAXSYxDOtlm+LBgQYDavvn
uVbjddCDBUhDmWt35Pf143CqG4WliZ401oRxYsIqeVqcbknb6oTCPIzxHyRrmCla
ir5fQruABBxsRBJisI7O8NkUXhWl0EwmtxsAlUHJCySkDpk9rDnpFGaVHr4/KEVh
GEM4CCCIuWT2yv1do39YcDe9QlCzz7HNiOyRgjvEHmloC0012ThU4KVw6K4OWgMX
2dOQIRxVocaJU0XBxiI+tc+kbYBqKKGngzYIpcY4hNKb7IpLu7k879s/aFlX/Qac
H1KtD38zI3VJFxPEzyX0TEvQK9ZbhkRjlumDiloCqIqH0gIwqi85Dv4QP+NULuqj
t8ou0bu1qyq16KPJpUavodZunN8yAOIRPTgW5KIHrhH/vc2wKbz5smYUWZZ7xKFs
oF/osiU8ZE+UTkWYe7093YoP/A2EaU8O5fYi33p4Yt5Xh/grUf26RGzEGvd/DBCk
wW+tNb5m94Ld/Dt9xddsbM+aH0U+z/PVvrZVPuqckhSZidaI6El2IYjsJvrZ031k
jGskVho1TvPDwasd4+W41dE9bmFrz2qro3/XVDu5ETOttM2PI3JjA4+IpJtYNzHF
/r0NoHz8n4uF8xUB+1qBRBISaPfgg+tEmPIPPb7S27ZotyNgRCTosZBxonabBno7
RUUgB32ea67MTop2uKN8bVUVunH078SaJ+/smjIYhy6IxikVT4ng8drqRPRCg8K6
6ag8mML1M4PZDDCUnZNwGdm4IIDQs7mvH1uy4M78r3PFuc+TGNz7KgxMgG6zM/uR
l+V5FcPzUorxU6f4wizkw8oYWESLhvE+5C2JHmpiKwxZ8KqCoqDMoN/b9V1HCxVp
r8Oy72hrqBSvrSMJrnSB3Mwl/3l+1k4w7X9U53C66ZTSIQ7F+yeRbbHjEvL7Sg3+
lcX5VOMdZoBohcPFrldFUy0AEc3G980ZyfePJbLZ5v3xAKsdIuf5nI/gdixJdY4r
YRuL2IFfz84ERdwZ5g77mSUYDjB3km2/gBaoVc+NLMj735K3rhPCTAAJdAht6cMW
3qX0gDF5E4ohFTfEsatjho1HHPfp5jaSqj7X6Ox5kbWvF04OLE12A//BRU3cNH3Q
jbkqHdi1deiCM/J7FJeMPnjLSR/Eqr/0acspf+fGMzjsXxmFg0+WqOmCDTNXjSXn
VkZWtJ5dn0TB/QVrpbT8IrDd9xPaukShhw0LyladAWMCgHMSWTvqfk1DCUN70ND4
duV88l5ASn8elyXYmDnhuaQQLA14ACG5MMT7kqkOX5/eQVQ6UdL9BxNAARx5kJY8
dg+CKkAbeZlJC8OKEeFGGFSooo7+wXozVhhg32lUrNXs90DMBuBsDBPnmSkOxyBg
/zLpq77GuXyeMOtHRukQjwOwtzNcTke0KmetIk5gXAstWeiAGr0HDb1xMOIHIFSK
Vbn11dnmkpSk2W8xb3T+KIdfIa8M/RqS4Hk+vwbWJxT9bqsvD0gUDh8LSEA4LwoD
p8W4koPwbBEz76pbncHeguk9f9TfpbOMLzbgRG2IIA/wGygrD3rMAmVZSQNTDQnt
oSn8XMAZdr1uljR3sCuR7+WBcnUD/NqbHHE+Qjgx5CD5DjFIs1Sd6Y9m4qlCcAD6
qGOVHqpisCKAtIzRQvHYCZIJuuLSZvbMf65oD/sOY1kUf7y4LSxhczVS7dPjhUR6
NWsoA3l3wInBVS+pOsLKB/1BdJbcc5thdFER4gaH+da6x95yvp+i10zCUPs8hnZM
4eRbMIOLT321OUYnTi7pI8dyX7FjbuLk8LShu1xOKI8wqIqZNXt9nuJ27YOAOqlY
zFdiqx1BsnjVTMr3//COdlN5Lzn3ntFt2CfxfEGIzrPsNjXIGn3WKlmvJVMMOxaQ
DlyxGPeDW7WUqFRblHB8ZGdFHcPaoqzbZwPhs6tLg+kF8qXwv5Xv/jC2V4ucclvs
s5lnxHyxJwcy3zH3UA6r+mK3tFus1bcGWbbbT+AuLG7d82YCtbNhNr+lPX+EA6Na
vQpL63lq0/28R508qUl3pTd/GsPYAmisdKAvMSJPYJk6syE2lzyc8X7WjMB+YsI+
5b46yjVuYK09mgS7Ap63atSkwRaua+dOVnD2xmiKSjZEq+w71lewORzNmIF7ow2R
Y1b8fjJXYvxEm9WI5FCf20HlxS2FE5ZajCIb7d3c8UQBcHJJFu0d5WxpJNGiS/Ev
Gb0f9naejaj2BjYkOV+WOItcUaAl1GE7cEREWPBF5grn4TakLVRnMHHk6g5BFY7d
YRHELng0KbTNmI+4iKLcrPBYbWOpvgPHXhFzUdKEkQHdG5r/H0PrWc2/W637+GiP
eufTlyHMk8tput22xSUIEx0N5VRvtEUVGz6yPhhYJ3jGTnpznYh5je7EfqGZrd+Z
gUuVpLh7e2I27zv0RVmarzqV5P8I8OxmSQRox/hghhL6dc248MoTqcP9yYIKFPsP
1Z8pdmaWuOBfeSZRnfsAaPUgyve28X+ojCZo5D324o93zZvpEBnbLyP5EJZIqrn4
30nUGHmYlnUYy+ymE7fuYiZbEdNXfIfkKpQJwcz3xG1h6QhXxxXR3jd8z9An5djb
PX0A8l06U+9Fwe+LhGNHZQM7laQnLqipiuUFonS/eWyZfkLq1D7kyhrOor2rv9jv
JiGWFfJ3eyH2qxAlhjX58WOUhCG7pUpjWvOHawl6ixvEUH+gXg9ue5TjwJNzuutS
FFWsr9vb9IQRnS/8dIzuwc5QWCiWVP2O/rZigbbZaxkU920qmS/fsSU5gIUXoY6y
4+SgpBGFwGfSpi0R/q5cf5j6o7ZqQuxEOfWOdXcxxGEFEO5X9euujLPRUZohCjAf
PXegpmfmOKgUr/2ZzVaftEwAYWiNRxvrxW/HpFSiTlJyDSsLGXZCK8CoHqY7wX/A
Sr955wfoVD20swO3XRPBo+WF6hogQqjsV91A0VS4Giv1HWyv9VQ6loUIOyrwhJ72
5rLZZmkR+VoVD3LN7JE/4oTgOoRBs3y43g2OEJRdPIAsTlc7jDXLAUaRnPkNraw7
nLzbbbA6oudkw28kCYqgcGYmV0IV3wL4i9XMQ3Mbqq0oIsIEZ1y5Odt6aRN84lzv
1c4kyWc/8W7jQiTbj+q8VX7hbZgswXoBvaFiaSj9a8LQuBZNsJxXif0G/QOQG7W1
++snwVVgdBf0Y91oOuEa66OswKEDZCyAVHL+cWIg7V1/zQsSA2YZItkmcmsAfDh6
wIbVEgcIYOyxUclEux3XeAdlAtuFulN3+sqvrUYnLplrE9ePU+gOSS9gaZV1qSPd
mgoZBt/7KbL1/IjSRmzjLJcVTKSYxx9h4veH1Gey5s2HjqJcdkMlAqeKhnR0z1Ia
uhKcjVI23dGj1ApEO/SRwHADiM6qbU6+5tHegYFAvDVvhel5TG6KXtURI1c7tj5O
Y/5TF0QuHya4BzJS/gvwphZyKpmoScv8ZlO8gIgcZLpw4knNFcEyGvAAuj2RWTk5
SkTVBpL7uMe+nSZw9BbVH/wews7lKekO8Jncr/934St4OMKlQim3Bk52XjAhJZOl
Ec0e/Kyeg0/XiiOiHEWCXyofkBSgW0asKYwhzQH88LvFSegyKJLZO2EUITnCjb/2
4jVJVyPKTI25KDgMSXCZgapCFoF0qJJUhILe53QUw0bOdhOozVVvhvDfa9mAHkLe
oOeqRf6HgEP8K3NJeEha+V1r0xyY+AVRqP/fp/AlUoX2XiJ1xiP+MoZACts2fpTT
Dy3nTBNT9wHxvSTUufJEYsl523P6v9zaz/jYoOATOo6xgQ5ZD9AyGAM13jbTZbf6
k5o0EusHml6kXp/f4IBM1QGvu/cUCpFvGNdEWxP+UB/vCL1mcs1KtudQGf3BzSwL
eK/tUYz7ZD0Ss+oNMEtJ00VMZaAA42E5eCFewe0AmRABOrg9RYyH59DtMF+PWN+c
yZoD2NCTellf6vFWt7qtp3F5YrC+pTMW1vGgBvVhsUAIrqhm/rjRyiDgJFzOPJfR
sU/0O9z71arRV9R7Sii+cboTliPv5uMyfwvQWASXxrdJEU+6btNsPnmZv4obSrwx
X/QYIv0a1UxOyE855k87B7J50xWDB1CGWaDuoZWieZh7u+8xdFt96+qhuKoTXiow
37nAIK4HnJFSX7MirNbsa5LyMLDVxbhiXDR1orPzWU6PU7jon43UK7/IR0L6m0Vu
xMULWHgf8gQXzjygM6F7DWdY2/q83D/38CpnW3OjePqad6Ef+CxqnE+4FAovhTGg
Hwx/VEcvIhJ9NDOKlpVtL7ZbeAS/oPHmAD2e4xcOcKHjKWvTom7ubEpSrdGouAii
D9oDxVWW8+FsIY0NuSBbPdD7dpxTs9qf9XRabFMjD1JGcXelRTul9xbi9rEMIQp+
RnfOZ4oeMHJmhpokHx50ihUfm+pc/HsKiazQa7jr694+kZ7XfJDjEyCGCSR01/ri
xrnNsCNi74vYb4DVB+ojejCGnhOz/ZA3cchIiPxoCPtu/bubLwb66dpqp2Kj0gPS
FhFoRX3Hy4Va2kJB/jJaMQ273u0BcTtTlxThp0TuGe3n4wTqPz4GVTRmtNau06GP
r3AnkrfCVRVfDWpKVnP2RJGnvjyRZ/0wHUwkFxkAw1a6uTXb/flauyyDaaSzuLWg
pMaVken4tImTwiG1T7r6orEvdGwCXsSE45SOPuF0nWoH91atBkTSyhiz5l82plN/
3CIsV2Wh96p61HnXzs0STsl4Zso0q+qwx/MH5xWHyxAMjADbgrp0vOkkWlSOtO27
w8RMgBSFHvxem4fW0poaChEUDIcrFiqiY8JgA7dTP3p6grZgTFcEhjFtc5NGIXhs
/5CtDkIfKNvUdqUvXQNte7Texrm9tpM0pJ5Af/vK/i54T7tRr0Vyex5X/9iF/Jv3
1vzkK6mnTOj0tPMsa6ICsFIxdE+ltgjs1wMdKQVunyv0oyq7sCjDS02mkD7rTYVT
k4xdVSBPIDl2Hk4zq5aDVfFgxPrxDVxnHrUyLpijgZ34JT96XHvrJa9pzIqxXn5J
TeSo0VsPJaDXgAblg1n7f0ic7OfShh5jEVv4x0j1IfDrt0X0j/4YAtXh/XUEQtXF
2zKi245w0Ql2l7cRj/+t3c6SehlHX3rmpyrUYCQWNxFAn1JmQPBMdIIesFc+qsCb
ugXQnTTI107a+r0LpoQ+c4cwUxvIlj/Gv/gUKCXj7Jg9iC0sh5IyHqnA0LJSNEyb
2l2G/6jRlPvJwK8ANXgLFcn/n0gTYB/v5khaTkc97FTUhMd2pc4tplDXcT0sA4RY
mYnlLilRJnswv2Mi45qTT2kfKiIriXmEllG19Tr+h/SDTnOqgfge4oLpiOPQwmVw
eSAZ94jWLSYTV3i6LGduQPIcW9LCSg9Qzs7P4TjXv5IhGQhwOkSBp4hEMikMItn0
Ozv7HkaM9dqsHacW9+6SLYLc0PCv/IgUSSWqTPMuijDIkzweedIOHVTBGYEPoVrY
/xKc5SHNHGSYXql1euyvz11uhApAU2fGnEsayumB0F8CpR7dOWNd9ynxfh9ur461
bXmNdKTLWEKOUNpS6OsvlDHBj/qN7VS2tL+pLzA+KCBM6Bm/we772hy0bMsnEADN
jKz3TH9aqeIMF9TZSfgS097cZagPWVXbtvJ1xJCyR3X3wuRWAwV7/prMMLUZNnuC
sNzXKkitvF0UQ4iWXwWpm7UG/LZ6TZ7nzEyiI1jH44FH2vaucUkuEFcxlGp0gS4k
NYTRo9ZNTPH66MbZPg+vT3acJVcG2qLDVdYBBQOThVLTIaZmZJZ1d9smcS+QrmZB
BuEf5DPLx7HcymUuj0d9RRX7BoxkrjYdyta19519ya3AlbtnUwVdbjUhD0D70/m0
zf3wrZNN9dKRqKcTl8MpWvSqfR3hGPYJj5mafRssZ9iNvJvRLZVToyUVNXnsLJwn
dcfkhM2DXiVEz8XWqZCWLcU3C/facJYv5Hp1AqssJqrSNHkW3Je2eEfysLbsG3R4
r3wT1pW25GNRWFcn5c9AzDHxsCI276e7xInUW3sKVW3TPYHtRAgGaCLr1N4qmS6H
Yb4TfkNUkJ3cToaDchA69w9LOGimadQEYOLj41JZ1FDXSp9KVR53rx/qQbcKAH/T
vo+X/NOrfBs4rWLiqBlGre+s/5myWsVdURL0ch4uC6ye9vFaPSCRhG3sKixTRPMb
vUtWk+GeVDdqoZ4zawulIkxbmTk8BdZio3rJtry96Fs3l0TNESiXLz9uaeCxAw72
ejJuAl5cxtlmQI4K+ShqcS5mJp3bCLTF/YCP9QByXPwtfQN9Wu2n3TgaxKcvQmNo
slATOd1TutXNkE7HKFbBq4HzVvFs1y3jTcjeDnOr/F7CG+0x2P+oSk6cqZ9obbcD
9IA6JRF+tiUhwyzG9rM5VfZNhRfb07XVgPHD0iCGUPNhO7D4R8c04+Urm+/dd/f+
VGl7ssNssyB5Jt0ZnJc5KpQS/MqchsU1NKDOuo/t5Q0c2ID0MlxqzBENGNadk81z
aWM6oiiYmPbgN0vc3d6ZsbY3/k9Hf+pfbHvN4lTDyDJANNlLdG62/8LvwwDw8cOa
FQ0dZ/TnASNb3V1UF0OEKoi3igdcz9S7r6WidZnrKxz7R0qptKUON/uPiblYzqxk
HdzHwzNOZFI731UoRly4NCnsllmaKYNDXlusWF4se3ecT5rTW+vD6jDxQ+U9FmAI
uzI/DKgb4DdjxhQJ6U65++pVq0EhsB0j1wq0yJ9K0Kpvrr0Aic2+YLl/8ILg9oDF
2OJ+p0/Go1w1tM1yk81I9xbHconYbOErV4n7zGtoQ4hQk5t50UB9lHIgDeJrcCRY
B6qSgSZDcGHL9Fdeg6WY/GtamQEnVmAhZ9zw9WZeR7IsP53OkduDJpIB5oWG4zzL
ytZi2mfy1Asc0tXE/ugMvx5hBvTpVxUVh9o2o07kJZjeCjwEGQIlSoFSEcugmaut
vmvodKmeVAEl2C1gSz0/bMNRN4j1x5sZUCRgrDNLa/HHdcr3jUWM+qfUCm6D4nJw
mNvB+Fq6U2azYR1AxMM4GCP8Y2jC7mCalcdBm+Bss6y8kVVGIf2vge/xHj/mxnaf
fzGi2wsdnjMIlWZaMoagUmcBtBbQ8Tei6ktDMLK0s97NcOgOb3drhziBqlzFtaIT
MkHOErBCJ+yrieIIf9/HNPgCUuw93Sg/S1nT9HvYjidBKp8C01cI2RsOWMvDXRui
JNzSmIgpivJJY/DmsBPngdoiLK0oW9IafAy9IvYhdCe4na1AG8EZfW/5aiUYahuh
mo2GeYnvg1u5YRg2M24BOHGpslU11ztvCzVaMcSrIf2LkiSHmK+zvqJBDlEesvrn
EaT1XgCLqJW2aCt3VIhHetmDAvyd+eYeMF8IeNuH2Iy2bzciis2GKfaVHpIVuQWu
wL4Q2SRkIDDopKyWJGxW6fdCVZyLKKgzImjY8djpElx/LmYFIlSBpGYuPfh5HdwM
fbXsKa4lSkG6XRj8wpWCsrx2t+86CV0cb0iwKqz3D5diC6aqFr2An8DxXbQd3asQ
ctpzKSzBv9Nosh9Zq1EcmrpZ48fMLEAFDDaZTkbhTxJcsA3WQ/cSAgu2D4+4MbJF
Ff9tUSH9ABzzeKhdN/wDjssYxL8XyxXLSSkpD1fjlZrMP1igA2rPhzO8uZCTd2Pv
W0nc1Zv8bulsJYziMHf7DCvBxMmHdlT22/SZz6xh46NnL7Fm4LrpCLk5LkKaNUSl
zhEgQJnmkR5xIWgGzQR1lgbD3cpl7FfWyKTVnU4tfol3Vj95ayYgcE0suDD65xpu
IXcCIpPzmI8dlMi4KpKsM4tQR+NS7wc1C9mXRESTbYuNzlpfDldty5+vBi0pk+/e
Nv1fJ5CBXu22x/PLnbf6X0cCmkGS3H6ldC1Ne8DcYNF3a9Rz+T9hikg1t/OyO9o8
UY6eignulDmA8OcxSkfJDwkqxOf8XXzTwihO+7kht9ByLbfGRPwgY9H8IcOdUU1G
4PS9VlRmpRe9Lvj7Imhaud2aCqoyTSJ/q+wXfXerdudo+VdGJC3Ac6UX3fQw5EZ6
Fr4GrW0ZaL/BD1iF9Lgh9p2YOBEz6kyQxh8dZP/z/jqdS01pr4IZQrSSnQded92S
16xeKX9EdLeuwapfrQVu8I6hHhEyUNYr9+/mzdRyTyK92KmTVVGi73eoX7eSt3RP
GiRyweTCM41WaOr1op+Ad8H7lAQ3rMbD/VjvdfRamVLmVOAZBXKkrTBgRmB0VA4S
YNM5Bq6D+GyWzZSOQ4E8Mr2H4R3oxuXfPnMybxDmdHGwx39ZgJ0ED/p9soZ4CQ0a
Iwe5qYWYlVlYewjubSqrQnd3DHSmA4yNpm6M7GgVap0JdKNGHgwd52cw2UgetLFc
8iHaDhV8gjje0FEb/+ZKurJpxr0NBkRqKKY1lquz2ssvyzuhpd4PmbtrnAH5E/ge
8z/+yr9fetGOXbgK8ZBMpRpPHDdMcKFB9WmxUdH5a/nLUuaK6yNso1T0l4GdSFMW
3C1OL2lUJMyv9E+1rmM6O1UlwjxynddDEJec7/jEmPO7WP6PYyXTRITWdaJkLYtW
jS1Wnc/jRW4cM5LEalVnNltHL4kHE7Fx4wHA9SX3jSNyB/zVU/KpNDvUaxuJp932
dAJnGAvRbodbveBEE/44YeytZeHgUr3l7pBSK2F6dNDexmprfaPiVcePkdHYry/4
r2+qifrpmvXPZM5TZd+O86tiH7Itcsg+uJ07ZbHLykERdIvEDRwPloj0ZFxe3NzD
mfF0CrhnTLVJR6Ha78XKNTAVHbgZyiAFjjORF3dK4iuy9KUC6O6Q8x5lS/36C4ax
helgJIFdOAt7rmU+ywyv1xK6Nclr71hDmZ+gvu4LoDVQQjQqjGH2EL99wXD0/Cmr
1KKLC5mtOZetD4RRMuZZ8lECFmEWceyILAzIsV1tb7j9sQI0NAV0bFSBmUVhTfgc
qACY5C1zb1mR1GdgD7UvkYBqu3pcNRge9MiX3d4EF/uPYK2s76fJk8t63kmADy4J
OiWeLQgVsdEGUoPfyGH6B7rxgUGDysgnuVy/sLn71yvsMMzbzWBEbndaGZIZiDXd
xZ46AbIq0QngKOh+nzidtpbTaiEda9yfsy2EmDNGdeRnCkYheepRLTLvVYW2O1M6
AvfvxyR3GLncfxVpiL0TDyRzg8/K9rFWusO/AlE53yFp2IUrfXqCORxKx/oBPKlT
TdaPbedOXDeMKZztPMTEsurFXj3kv3ZLt0pJ/uEZExzHV5oKSJHKJZ3YyQMlXyWr
he/mEO/2opELHQ4nuv6pF4FfIBfFl3TxOoirVCWaQlF9iL2Gei+MmzD3Jxt8znVd
XAuppQTirTMaUVgYTb8UPbOpv24ygfLFluETw8lAHTG5jfU+1pwCh3GenpeLKxJk
fipSpD8OJR0hCaxzuKZoHWWmiH1jpzJNtmSlmQhxePB3TcUJn0VguXirYlhu8jMS
3mnqqN1tRQ5puUN4d7Ia/CyIimNTD0ZcM38OzQSBz0FbQtyjdwoJ4aYnMy8e3NHX
/S/lywedburZdEautnqCP6DVSxREQuEy0A3P4a7NSWxzMDRB11kVdH1PsBlvRYk4
n2Y+X8TT+NOu6YcsVFzvvIR2Z1d2xZgv6lREd6UbKQg2QVXqDkT7pFyhTL+f9usP
WKs1Tp1YL0G0MCg8PGDOK7T55OK3RoNaxzq6vfhV36LP+GwnC204kttglEMuh8Co
s7gQnI0Zj4bkoUR410z/gPQngc6TcoquxRDc6sUuES1uBigNoQH1B9AP/K3R7hk4
HnDzxxjx2VKIVC3NiVWR/cof9ka9a1nJt9svtXQCl35IvqCLCSkvIv0UhLjDDvMR
KbjKPaz6pHj782i0V7Kt6gsBMdoOUnzsSe1K2pmEsf/EdskliZ5tqvZa+EPZ7VhD
v8rtj6Er7DPpmgoJD8dxVV9GZD/dj+pFLxVKbL6cH4YKPpJOFmpUfLMbn3R/UqnE
7Vy+ZMgSj5ea7VAQo9LEQoloIJ0HTV5ETXFELYItW3+hmYpwnhqPX0s9O+tRgU/5
An/pg0zkZflLJ+MI6NBRqXaEZfttErifN6Hvmpiz3xmfWScLcz0v99bKw+M3YEAf
ZgtnGKGQ2EfHbyX6UtpF71ho9b1AEvTdbl8FJkIbt+Z6s6oOxtxodLkZUm+rNmyp
A58j1DPgematyuUjVOE56rEu3zvRfOVB3kJYpB76Zx5OV/hIHL7+jiTQNqlYwZMd
4oaJtHnrYlBHjlMbELwbYlKCIviOOw2o8YR4dcf9bmRhYAJNg9ONoy4Kgwsvzrs1
+5jxPJK2lnhnHqBB1OdyunFqTD3U0pYwoGN1qdM60cyYPA+V84cKmVtEk7Bl1RQ8
bhaq9LSS9ENTabWC1ABhSWFIhbgflzxEtWhYsnDUUgKB/mlTFmSbxMMWjTnIaGQG
SD7CMNONDDU716bUk5JdF/a1ppe7b4UrgfaZvmKa+CleMZoqrpz+vkxPfbWYPiMm
sKaM0I0AFE9OmXJLrr4KCRA4FJSxqQsw1wayPdDouCLKv3iMhW8HL5FuUlv8ditn
eiy62CJfwgHL82pnEMCP11abjUxmmQHfk5Wt+liS17QJHrLKiIQVUF0wU4z8XfxN
nTmb0Gb2FOLed4exqdkjvBPc3WGaC3W57z6JwjGTpnXbbCfNHCxwuXalkcGM3qc6
/pEeydZ7fh62OBF74TN1TNCQvGkzsCZw3ZmozxHhHukGUQxV7i7rC5VOxAC/V6Ki
IjAKIERwJNiJk6ZjngOcVeWTO08ps6NUfnSg4SPpUSw12M/RjgCpuPHlzZlgquHc
r6S6h0XxmQ7q6kj17MnAMFgC+a9+Y8DRUUTop/ofk3OpFJORpJotDV2FfkLYs8Lr
EyA1OebUOUa0cYlTeLUfzGMutQ/ENXeXvunjuHTDLQWYDK6blRDIr8KsAB1bCXKF
1K/+JvNJNPXKcP+mXTWaioOvcXTpFrthZxbJCaJwEW8MtkzOQxLqBRDI6DUSmCuZ
mqwD8av4fTJ8GIVKnZOxgVQKo2FtgLNRGTADUy8as05s4sjkDSsk2YFxcRJ2TAn4
wcESnZtrZ/O7rfYKCLe/sC7W/rEu7JFeAKoODTmlzOBrYrwMrYoj6nLprJE58+vk
Py5vJBY4aKm/oz6vngy+ZTU9BIj/ewMcPuUG5fzpchQrzPf/VqlIRY8eA4pshVew
hQJt/IfQUSqawMvZJvL7H2SGBm/OfEK1TCLtnUEe6bqzhZpVrjB2mgXOXylJ/C81
tdruZEKiXlEH0Qgh4/xh5BWzntrchR89t1kwXYHITcXyxRDWx60HwclDBCTZ3v1A
LEInow+tJ/XkIldOjkByvlXMd8M7zlqsB+Jf6+bxzwC0JCSAC+A2bRTX961v9or6
QGZz+4+kp/bk0JonMCgk+vZ1J0hSqnAJmx4OfkwCixvzl9vodW1LzcHJGufV850h
XENFmhRNU3h+bSANb1nTOMKBJ5XZl2fsrgLEN4jdSW25DVWBuUfsUPKfBrS0uJuk
fC4mQdKfkG1IiIf4LO2Uo95/wuh7w38sKqqT1bJ/QGIqm46c/ixbOgxpNhnPuxO1
7q4iPbLVEJdaLfGVozC5WVlJ9gS77zrP4ag32g/x24eZ/uVSMD6xhkyuy5pr30PE
viWGXTqe73/xIOXMcvs9G1jvEomjca5KM83Tg1DBerY2Qde7TT/M0F+widfdZVZT
3dgU7f5wi4fZyW7Rn+q0ub8j5FcgtXbiQ8HcQBauj3xY748NRqfTQadRfcNKZJki
CjCg5noYlZq4aIZ17HX2i5q0Hx0IBIUXMsI8oJLgazu/ABjExs3yVmKHOrqhEvWN
5bFWELKZKXDVnNTy3gURRPNN8NxKmmkyimfK1b5ZR9j6bSu6mHnRXXqhlLQ7duXp
CIE8HWRXgT3O4ABQVlips52bpe58oFoSoWEbluT8WcXEt0gcKMAGqDQpfSnZYueQ
uEWslNjBJYBOxOAshIom++aDWxOZOXulLWMQhCMVvc6LReCnf8OAYf8coyv3rdue
IGWs1PIehIK0iUFEAkglx9pqiOb1vvUGDkzVc6MHwOaZ65s14nXP6q9PSRgLTuo2
8wFrTMrTdZ3kykPDaQkO2aiII7YHKRWJCbUoS9J6nJJ0esRBE6Jv8dAzUFds1kMY
apAEIbggTLOc+8w01vwk7C79jFdz+7LUQkCXOBKNeqcgwUpXOIh89759iLAyLb0L
vKsU1DC0SpQL+gdi7dmY79SkOEptijZa2ZfztVGgg1utiMIRC/rY/uqEs3v0MDMY
KMqzk5n19FjYss2EkjaX8zhn8qgpSNtZZDnPSbaZmougV66kS4OZgqIqn44fCgAE
cdsU8RdUSXJmgFD0EHO2uo7SaHzIyI2hEifx1r9PugGqlJwCgEl7HkaPf4dGFgKn
sv+NA4y45ztiK4irXNnPais4okrl6UshgWUb318yfh2HNolWoJ8xF7OZb3xQzrIO
/B+jmfTn80S50GwzJM+N5mr9tKKo3z78DY67dYQt0+bBPgcreT34m2ABm9vlAt5Q
srSUf0GgxaiZEITB/lyVI2kaWVkwB6zxWKWn0riSWRkBKh6NJHARLicVcJKbJMmB
KtZh7xVZkHhF3Fq704IKIKMYKBVdFM0vR8J4hgmROzuHYRuxVUNnFTCVNADOF1tx
PhSUduWqNkSW7KoED5BcpDL0O+WZjjO4Mnu6oH29Hx6WczUAMrHV747xVi+nRSEY
2xcC4bQkiaMioRNtQXHOulv2SHkpvQqJXME/2YEM+vfwP1CRojcSbs4iYshQ214a
J1E6pCBlDSIwjQdVoUxN7DDkGyWPeSvsXTtEhXr/TZbVU5bjhH6pzg7YAdlUG7Rl
fnhNRPL2h86qfacno0WiJleOYbUjZ7W7FdySUjBMHSa/zHQCqd0VK3b8Jc1+r0eu
zfGINYIy15qQHgxRXNbL69fl3zCCkRUb1NsMUy4ilCDH01p8cxBbVaJiADgQV4ex
A2jlB69eP5MI3pJmWi1AthssRJ6Qw9hc5kwBblrNFhgqKEIn+DLa+FksITeIv5FS
2iNgCXdrmGm9tKgwL/zFuUt8XJzr1gimL6XxaxOkkrB2Ok/fp1D6j2ot25rMLni3
b3xL9lRNwPws7D99e8vNXj16b17HHqi9YBldhi74mxTebNMBL7WfaeGTtxRJzUlT
qKv/+VVzIpRS9aXjst5novOmCn9jqS82GRIGUo5pfSgXLo7eOo57jp1dozjfi3nV
DvUM3J7mjrsYbYqrw/izi81Edka/zWym8OjbxdYBNMLc3BvH9XqmQLGQGDrOTMQa
gxQKtdJD4aycZTtMbMqLUKJj20FSpujjeg0/zArOWqryHFfIVueEJngO8xam7DDN
WpgiP1l9s+KkkGp5JY1RKh84buImLFOYOgcIW+ImleTJZH5Vjda8UG30XZPcYikw
mumP74SNjVI0K479lIghRcyxIzN/fAkU3tjguEQ5Ml9LsmxlmIUbpmaGZ/C16Bq9
YK+WRpnuVlp401nlcfbzbuP7cFjMmTsN+YPmfXdEY4XvpPEGHHFthPnbAhEEZLtP
hbsjxAb0QjcD72NMemV6soNn/xsniwWTvnXblG2vF033AGXGhb9gVIfd0eu56KdI
jv2Uhgi5aEzpOI62VZo3DXbqImiHAnfRO76vXAaGR7VY8T8fGkHTIrMirqtxDCMg
+h893d6MzXphWEJ900LlIos0odnu7EqQTztODX0ZYrC5aLADYUPB8fPpQsUScnHD
vxxqmQod5rAT/fwWGKdlQyXtcCsgL1rt2I4VWsMDSS71cXRIRJRqd/ezyejwbMLs
j+isqSsH3jZS8o7L/CP1rN/gJ1awKCLAgbYd9RVDuEsS0KAzPgKm3zeE1dNTPZz/
2YYzZ4rDwxk6LXfCwL8VSvwaSOx7lwdlcciOhOHMuKjfp2X7wA9Oqa5GaSQsYdbS
K5jC5JUMqMMu+9nnlLJJAXvgZrZ8FcbzoFj5GlhJ32KG5lklEwKw1UwnGWxKA5sz
MwaCAnz56DblpUNimKndUTsPN3EyojIFzYs9WXn7CrkorNRvCCW42YhWkiPfAYHD
MXFUi91iquRdsP1fGFISMjjprT5TUIuQA5gzoQEIy0LyU8YmJR6QM9S3cmeSEIWD
rXn/mlYyzRznoqnvgr1nIwb+pj4c1agmos2AKE+JeL+zOFgtohcUdvUtVxlPam91
p5OfH9ymCWFtafMMbcSO7p0/SUA0LDCq7L+Ej+SqLEdxXQs4GJJLnErlJGiE3Mcg
TCsyyBVLiq4rFUK/teRLxp4shVmowBQOoP8KpAC77BFVMX/wzFE7hMLAIB035mc+
++RhPkD52UePzauMAzxCDINOdyFcAQkFRLQjIIMO9NPJ6JYFWxbLFYI5jVASn+Ba
/dwSEEt4GE7OEVtHnV4z1v9jNV9wtmcpCsgKDSbiPh4ChdNOiXpEZYeOvAJKr/7u
d2UNZ4UsqhX5Nk8vkYT+FWPg9+/eqLLQslmPfTuhkBolb5YIGZ0jjpWD2NhBOx7N
BjmU+TxsqQpc8yJN/PiO+lYrI3g5AaxpFS7ybm7HaisA+mjx5X83TkT0jnmU5nTa
uOABTKjlbhXSOtEH3Qpy/T2UZp+3Jr73ZcVtF8692NBjvo1SZN5uJ8NAJOXov71A
YTQmoV8x9zoOo56UUZN1jINRKxZd6+PcWt19ISzTNvgRUyNPakGRU2A4Kpd1vm5f
WQS1712XWlbTqaD3P3c4lvnXz4IfgeS/Kcuh/BkyrG5wKSlZkwLcp026woN7V6HA
bSpldtiMi0J5s/CJVbjJ6lspmT84/o5pEDDZpcFkyVhWxoj21TUgfn3dfk83kytI
s7EpvuW4EDJskrAVE+FPP6T12YW19ISkEZo69nyqo1EKrXepbQLRhEIbYw+F5Z2d
KwEpxI/twjbxSOb4uc8G204OhRF5/xxX3GlGzcfgLqnCTzD1rvEgovaX691buMuK
pKfCIKkuURT68BXW/tq0l9Bd/yGG4Hks2uY0cN3lqaJFNn7KE7jZcRwzfaJKVExN
iunn2xLHp3QX5u4m7bU5pLbKs1cO94arzYVhMoN+G4Qef/N6wH/0iPflSYcumv2e
hxfwglHb3foT7VZVLsYtVetnVAHixP3b4Xkf6G9mT3cbPd4fDQbL5N+nrJj7c9qJ
TLX+u64TIXh9eeCaxDTKAPbGzUV82PbUyyFSNIWBfA/KbuC8hLaCg6tBauJH5LSI
A0o1AbeOjXLIemV3v31P7UBfKdEeb2O09BqWM5zzJf/BDErvjW0vBLzs7UzbcbxD
pC/PfvQt6Q5Y5/TWFqScwELNzHEwriCwQ4eLjosG0ggBqIoCi8bf0K+nYyGLymgk
q1qB3ydBL/Sv/xtTV1eCXEyeDlu/2UJuT8C47hrYM6/ycGXjld13YYqSBJBzKs6O
rGoWhtzIkdCUXsl0uvS5dTpzeDKT0ED66ViutNdapfrQXJwBZQNC5BjsGE50mdqq
uFcPsBCgTrsmaPj/OikjEB9NKmjHf8QorusfUVoFGogb1LWW9B2uOK+ZNpTS8oeL
nUmZxykvjAyBd1nje1DycefHTKIYLoHV4jcwyxS6yBBmbbbQT3f+312fppsf8WzN
wWqAjiCpboYdwREsq7YPJ0ISJms4lRVED6r9SmzumROJs5k7VgPErmuRz4A5vHUX
B5vClvZ7T1hEvYHEB4L/CRJxuvzHYAk8dbR7N5jbeZPY8kJQtFaEEfhawjs6jE+r
AeaNotFLYyUJJX7Qpy3IzqOhs7tQZHXWHvslHHJmTB8lAq01tzuZ83v3vaTbC7Y1
bGQfq2YGeke+y7du96l4fuZ/n9LZw+1WIx9c4jHWYU3Cbfk4DHmfwOl3/DYIU9cz
vrGTU4Xzs8ZUaWCBg+Ot2szXm1e0tjYCCkI226icIK2vAZywDCi3BN1hWscdsXyF
6xMexSnWG5u+ozucF+74+RIE3XrpTpDhEKxmXoI+qHp13hhuDsn7eMgW5DwLqFxW
LMFCutPAkmcc6Ku7zGN3jPAF48vJujRWe57I9GOZO76jxqF+4A9PljmNZkdb6dzk
duk3oHqep8MbknkeBFCqoP9diA9//qKDuvHC0vivn2aK5dHD4xNEbaOwYkdf/wp5
EJ33Iq1TCnFsj+Yt3yElQ3Fjb3CoLsI1HDSQI1Snp9nC1I/Nz90IDelGFB5vwzsS
ePh6Epv2I5As8wM3pc9FM5z7D0E8NUTnIBi7SBKtHzzTvsQCpQfklCKQHWJshtGp
lSrL6nnh9Cd1sWypiAO1cvm77bgdkRXnC6GmF4PyrHRRzbmT/wYolAdhPDsMnxwR
7EiM4UAwtTMYWSCsg7x1OeWOGpcRbTqUznAK8eut6lSIR+rRYSsTtO4JKljCHpxs
Wv+F7ywRsctPF83qICM8IsDbn1meB/nGCaknYs1CH8aH1aAd1uRkZH8fT2zTLjph
fd8Lqhby9x4y3x1iyWPmOVVwZnNRTX8NUd5nKqtrN5Vb9Ep0FUeeKJF+ydTHNj8p
SkSOPvD6LVKw9wanP6sC2xHT80DpNP4OWSNCB08xKBEoCL7S5Oa2yttkDgbekr30
e27/P5iwZH2Kb5TJNGE1iqU4d9v3jMnDEpcFwSVDf2lqTc92c47NiewaMemSLNyJ
sijoaJnCxNkL8vKtD0CLKx7CEwgjB5c/qm0nIeomJgTpeWohdlUhIqy5Sk8o0lmH
3I9We9v9Lol581qz0KRsqfUgFjcK/7K6QtM0dw0JL6dMZbsRnemPtCexNNTeSkHM
K4Z5WzfGAgMzrgMRoaHcem+jNmNTT+pRMCQ4azwurmR1eXuDE+b5prTvyRLgtuxd
ehMDRHZbKWoTPQBFFzd3Gzhr34HKVZE4K2yvmRjtp44gRz7VFbiRB4l0RbNPNVFo
mYbGagyX5rK3zyXXv5KpSsUrYagPIDsA2z9/EAYq+dwEdEfdOk8FB1JbanZQ/uit
8ci1wDU84gyO2FaYPjSgE59NHPZVI96Q5FUv5AZfSz8l/+iR6zLaxbSWPcStUPNg
nfF2SplGEvDi6FBk8fAyI74J7HlIQ1lTpLRRL+w8MWDJx/voxY5O8zA46TlxS+9U
EGtD+JUAmfRTjEP6wlA2UeY6lw/ZYVmGaO3m/e7+z33fWvtG6lzYjRoS0ZtBNkiY
X7cBuoQ7QKAc2ukVQD/j1MS4KctaUaOowGh9qxtqsFMJ45tS9YCxj3mHhXqJnZCe
IUs2Zg1NxeGZs62lUORFbuIOmaOYtve+X8Gt5XPoInp0kBAeys44TOLnbS4toi6r
fZZRwPn+aPsAr2Q5cSxARb5w6LiHw39QDul2Y0fgtebHY1hjrQhfhm6xFHdBo0NY
IEdN7POa681zAq3ibXCuUITgEoS331xTnNFP8GZj5YWaPiCQrcwuX2Dwe317jxJl
O/nssSM5Q93+wi0GyjNt6SF8mXdb1KEiLb7B7m1AOJEq4IoeO0/e/LQlWt+N9bvn
96ZOQ1Jj46K+r5zgya62rdETzjpD0pFS5Wj3pt/JxS3YhC0bNseV6YBW1Ajb/lBe
t/m+7FvxZJggFVw4YYG0pJiTQec1+gEchZitPJ9/JuAJ5r7OeSzhlpzhv73Kem3S
xBKcDZHplauok/o3iCxJ5whEtOFyXl+Z80tlCL8hYvKYqfcnALPZQCCCRT+JluoC
hWE64w5HrcCnj3YucaH84GtVqcmKrPfEI0xClbPzevE9aZmU9FLJrWsp0nyJsq3V
OqqiYY14O3qaYAsDpRin31CY21SzjqpR2LEr5dRx2aBqYQadG8XrV4Mv74FxHBiB
xSYcvvlEStwiu9MV0IrqIPhu8PdK8f3APPDZtFzQNUgFctie9L2q99SPMOpV1CUn
vRNf/hz+mRDWEL+6mqphOySUXPRskNIS+Npqj6h+bnPiqgCNAp9lEN2jc3ezyr6m
d7eQAiTPEtZzteT+s6BLK8u7saaJ8S1qNKSIRvUbjBDSuho9o+y7um94xNFLdiqZ
1/F+sRVTf/zffW5qwIn+qKdswoz/BvJNVMPpEqJl2WFMePS9Lo8nR8vwASt9NKxf
QqGWaQdebVy1awq0+r/7Y8MlSOfTyq8W2LHhsq54XbyxxT5FNrrmXfkjaE/7PfgF
lb3+3acnwdZxez1IlOkkP19NK3zT0tH+3MPFDSBsIjkiq+VfscuA2xgGtC3mK/no
w0f4xr9EhztIG4/gH//sNDzvLm+Sz8uQd9RnTY9b7hSG+745myIa3NO99bJKHVFg
7opsfI0a+L7Dg2QOnJInNEjgcjqtYxrju91fvPanw/IoqIuRbghB+g4sMZd6fXDA
8y02QKLseS7Ev/OagpRRxBu+BodxFz9svvqmHTwXiIO2sysld6k2/xOHx3EyDnUe
U8KHqsLZ9XXoTbIk0s/iGYtUmZnvfY8hmxflt4mdYOWgm5lWgH9N6Xn8SGCXPef9
ZKPO8hdict40K4uYWYIKnoDHIrrLkX8hOBIxyqpozEGuMyKjzlyOMBqqNlzjW1MS
Zb7/amje9pBqvdFxNdJ1+wUigUOyfqd57qj4JkEZARjvPFCptLNa4lfTSscv9cCj
9g/u55Eg8/J0Y78nK6s3cDd4iNpehLYfEgbuySA7OHJZW1/TKp+GuJxWOEyBqUBA
CLfkwRxR2RjLxDwTV2Geli0QU5jnUf3vN++doj6jRbcZgkaH+Tv1HJxr45dpM6Hw
A2VW+bvuJNHbePY+m3yvOQlJVFIV1E0tpA1XZXT/TYtUVncp3IQuSC0T3i8fr0tF
abUkaFhNLhfQa4TJKCVxmNSgmcelqpz/RBAVteNEpalJFu04t78AIqmiLmW8kiLm
97Wqx9/Cl0zO2gECEkm71K/zYnLq92VU20WDvvA+yACYaNLlaX0wGCmBlbTMHR52
e4eQ95lPpDnqUM3g53QszCT16Z0sKT+PMlwG+b2wPdAHdvlMB11kpBsMTmi1ErKd
XoyvQveugCLQQz9NgqqQGS9N+/2YdF3S7R4Nx+c14v+M0IaKLz+e1i6vcYEy1Pgk
t+xuMGfB86M54DAppptfcMjZhFBimUkfcMNx3o01T5Rfb60Sa40nDXb6cKOVNhVC
R/ycqqcD3ch+ojqMlY7SyoSvZ3boviZaFVgWFw4OMLphgufwedkZrGf9tqLP+gQa
Rip5abJxa8/mFJp1L3gL9zckMeLNgSTupIWtGWyPFRzr95/OpOQbj19Zt2UhV5VH
+kcC3spPYhPGSqJHgokX31pdxqMrUoH3xfAoxCxKLgdj3VEAjGteaHMGXIaHP9+P
K/OTAPVNREfdn0LOyKr3H52PEoAjxBUeyaQ+4UCo9bYDst/nvwEMYo71dzB1xsGJ
V132l/4fwkmndb7pL7BvLPG3E40LRX6mvad9Nb/iVUZ9Yns3Z8LgrK7Nspbc8lNr
cH0S4UZgso8E6vy6cmi/u+lrVTHZZ4kvsjX6snyhP4CbqS0rC9cnZvTdGeA+6R1R
Pg2TPw8pDZMY78NgsXI3TZ9ApC23l73s8G+Mz+XaLoj9CWOlJ93vRXSCF4Tc+SCQ
HrkUJzKoCOTgfjVKMTny0W3dOg2TB51uCFF5hlo4yn85buaiVDy6HEo0K47TUfgq
kyxBoJcBKif12ZqTIsBC73pxEfzMYeFplcAfEMTAyi/SfBq7VtbkreM5dXk2VFCe
qzxs+AgB7W/WLIx0tQXNacJVNAO4siI+GNEh8qDO5JkuEwgt+U6Yxqr+PqmC9DwD
ySFdadwABSUkYzjryKQw35BqAoWF0nHE/4lf4ekFW8V7vDttGd+IC898tiYWIF8g
3bMnado2Djt7lMPOOIPa7wDD+a/Jqdi5fQtZuk4e0wxG9mHEtyNWi8oCRvSBeXaz
Jqc7Q2omgl36/HJm4B7Y13g5sd/zL+JYr+3z8Iekd5bI7ztlAZqJTU8AXStzvdi1
9yre5UckFnGUR9HO4uKVCNmth+Xe6OuabP7q4Sx5BAaaPv+2uNIlNHwDAD89sisZ
2Unrr033gKi2Safc262IffRXhJO01bHYdWxRTxwm+DiYj64qV+upaQSFLmhb8vE8
jVBlm+s348Klr1aYRW89Pe10c8zwvEgwLAc6r9JWEvL+2irjTX7WLS0ftUNxmvwb
1lU7rC99MuLfGFCILsqJcS9ibdhNmwOXRmS8C6NsiQ7cR+19ldQfBxyLRVYmT/eD
MBEVPvNZp3848ckWM3pySZfTDwmw38aQ6sqnnbvnwsBrreoS6haJMAQXcq+W0YKZ
ly0ii1aPBcoLKBh0arPj0WuSGD21CpgO3bwQVCCHYCdsMRdTkfvfwxIg4zSP3mcI
bBtcRzOmEl7ubwsJaK2CtfF4H9fyWGkfxwVMiWPPDCon994JE4XHG56tziQOFoBJ
ar8uwdG6Bw4tyTikrqna+nPlW5QVEhyPWQGeAgfVIRSOFaBkbPVJNW4Onk+bN7nS
YqQ9kEaq973CApWVxDrfa7Be/W4o1u29nTMbmlTcg0wvN7CDPYeQ3BdGWeFF2U62
Ba6hZT5G1nuN9kfLi09A4JOKzU3dGcHM8Ef1fRBU9XH4OSU45EizrF2OkgoG6o4y
fL2kBrSdmBOTYv9+sMjIvwYV6mFh9B4XKDR12IaXDfJy7r1e23hHY+5nA2aRwsAQ
JpZBoR2TuBX7+WybeU6eBF2tJ+6r2uEDefuDWpYeyMT501kbV/twBRblGnDUaAlr
RmutWPRDpqIFFr18UaLRmxpPJpDMVzWWZt1JwvS0XG6nd9cZv5ro2G8uCytvXxAA
1tc7eqOfmvhxMSY64JV8jZ5WE+rPjkRl6BlW7nM1zDPcu4qNAkjWN5XXhaSsRWHt
J9Up9Neuh7mweBR8pLqK2QW7dv/sgKV5VkDZq3kvfoJbpwaVOK8n5a2FegGe9IvV
n78e++eSNGlPxaRsL5+51N23NqgzE5IzizipCCfHVvG849oEZA0+0ZnLRIwDG+xH
rr9Ul16ARJAoU2r2K3+bCbuAzfXFQ/drMc3HxA0q5LyAhavQGnPwwEWBMtw9b2Zc
3AWMtqO70G2To51FJzx8y6TdrQYMVWPAggazbEvNO1ohs0t+Zf3ZiJzeBo30ta7S
cfzhUKsjh8ymKRmT4obQyI1wY3fEpWAW9QLJqASyH6XD8CvxGfgszfngKHqj1TAB
wrZbBArqK6zTDpGHmD9Py8y7PtWl1/TopZJxNl0u/0cOm2jf5JS3azRQi5qy4eOi
frOmZeKHvb8/DEG5jP9ChrtbqS1dOtQT3F2OcXd0WY7eufj+P0kro+3OEcyfrk/U
yADSAckzpmWMQyMJ6bxR3CiBSsJodqB4M+vzOwP/ONiT4u7r357F9lg0Zv9t3BIa
QFvZKp8Yw9sNI6TuuqiYYMYVAq/6FTL23+YxPGyXI/yyGWUaWPvnBotu+0R78RI2
hHt+izxC2MJwe47dJ5BR8eEKea9kPhQPmgZ9lJG8S+oC9T6lIF6ISoEmm4XfMeQg
N+uv88ZHQGweqtcflwuxZaLfHp/u5oxtP+W0dwfs9kozQUYZ/R728Iya8Hy140dp
pxmvdgfm+arAndYBjaywepLDlS/1SjKZOns3NhNc4LTTbZyKmReoNjT1wlcCYR5a
5Dwe0RBOrzq6m21lqSoFHYl4UHn6b+ZrNbElW6YGxHeXJvrOA8JaixMkmh+v/ZQn
pg0oQdkhnLDhMDFURU4tCX97EEQLB70TxcvaUH6ricsdbbDSbtUL13NtFI7VQ+2y
aM5+mGAXppR+p3asPToigRDJwa7nnFJvADlffxq8Qz5JhL74oVxT78AkB5t8+Pdb
AHz2avby7uACcDLGZ0r/JNZR0xbVclm0Ay9JWrBuZEdNvw2/hK+Su8aM5toQrfZq
BOy3SvffMPcdEPF6d3faZ/llJzV/rSI3J6u+0oSXM/cqn/z29JftpP6KrrrZ+a2Q
Kl5SK7PWykZHUufyE/ByXDVo/u3Zh1uzq2Ui5tmyXckTABr/Ai0ZsgU9Uedh0Cbr
6KuDbmhOWJh/R7LPDr34zaex9ACWsL/zpCE+a8SzQrJg79QHpID3DCux2HAyrVUz
fl/VQVkqOq5/bc5uksaSMTN6W0vhPTuZf6L5uJ3vBGQQw60PkpIT6Eh74IfgU6HQ
JcTsMINUwyVYPxTE/ezq6yCqOH7xuSu2ywTmpW2Hx0zvWUebe3yjV9OcFA09/pmw
/Pc+Aonlliy3j4asOSCZ1mpiOV21jEvh9z/FwJP4vDxBEwVsQdCzbuN/090kRMch
z8MSE9OoGvLvE6hLeJOXbnRenzKVfMjM/LbFtMBIiy6cbBQda86aFZtX607+ukl4
JXMKZBV0l17sAFCgH1jmdEt4u37zp2DR06A9MFI71NnprvwHV0Nve03WAijFyIOZ
rlP0WAGftUjQJb6BcP7Rj+ZNT90/EpPo1rx0epB1sgu2NUkcvg2IkHdarMHcE+0C
ziCBtvXjdIMD4I1ZXqTOVTrSaResIlmJG9KLGSt5TdJNXae6in0C+5dCFWXU3omW
gmhf/KfbEsvIsQIDesfMbl25OEFqS99aZLdiO4HzwLTi5zOEtsY+8qKp7FOEKonG
1gOFBl0WH48cXjQIaAeoCea9S3gTdmEyDdmcVcSwcS21qIeijIqyyxxVovcdbJw8
RffF7rNODLc2fNQl5KTh7M6vPdTBoqj6+wUIVCN4UB3DrW56h4lpdlEawrK/Uzdg
yRDa/EnwTE//XPuPDx2b7Rfn/7z6aJFeuqCWueNI/NimgCf/rTBG6zRgkDYMAC3q
PTJU6gukFjlWiVLEMmCZbfq0FF9rQHROkS8eirv1TSLp8sP9N+XiUQb9L6Ye1DE7
5BduwPhbKMs29E73/KeaY36XmVYv0aviB2RywAdzqB4JvMC43q5cgx4Gjp3Fwebz
YQ9aa1ns9MYrYbCCuzdNduIqPaHHi1V9pFLzriAGdQV/7KEmhKQDOhdeACLggUhV
v0WeQUqq/U2ee5ujgk1diuKkpXrrp+uAyswllFX6CQuqyG9kKVc30VYkSZaDHYAa
PR0EqmdM3IIwspb219Y7gBPx1Bqv7fHS8UpXR3DL6Mc0XLFrWsvlJrPLJpS9bSH6
QhI/uN/kOLN9OyLMg7hlaOAMRSoqgx1QXwAWcbQMYuwEGtDZ734aNmPdlIhjORSB
TfHWdohXICexVvUN698yrmk626m5ZAcVlqwr+MyaFv8lGW6PzCs/kJicENEHGAJY
4a0jRwW6OvBRwofR4huuDQFcvqbzFCj7mPMo4DRP2mEASPD7KiHghr6Ae/KhnH2o
3+dZmLHBmZF0QQS7yK6nCmzwyTOPNUmzGawG2KEgWy7Ydake5BMQLA37owFypDO/
F74h2hMc6kZHuSmUrBZp4ak4zZVhtlWIXOLq2xykcNmKWfetecBuaT7jT1KlKDAp
2P5d+Jnt22urRsiIN25oUnrKak5UNCmQZXmvWS+zKNlT/qTwMLWo4OyOZMyaxNwa
g9TqS9OGmiOgAWkOF6LXXW3WMRJG19Y3Q/irtffCMutsGOF86peEKSUZ0L/455dA
1oZrUkqtEQjXP1if5WA+Qo4XD7lCyYM5gk8gSzha57/FjAsNKpuAzRg4aJ9Xk/5/
hPEdl7YbkfjpWcB/U0qkLUx1F6SiIUK69F5SzouaXQWjIvUXIq63Tk3KSIj1/Wrd
IC0IQNn2fT8AhwoZ6Y8gO6grSxMvk0dO82eht3BwRG7TLR/zon2juHq1x3a0vqNH
EIGUTGovFxWf9scvAd1vRQ04CXDVCl9KTzgsuX3YPwLdAP8CSFEKy/1AxY5ananB
iZtxqpmpGzRIDLHIaNr0d9wBZC89CmkJoUFxiefY1NoIOaQlIw37VJIxeijMbZdg
qMu1umFOEdR2oUBJN06xzH8CdhW4kh91vdy0NLlpcpllF7joZdqbKmZCTJXqwvoP
+eMKxyrvCD4UExLEdzFV+m159OQnqksdJHze6RIMNCjpBGpG1DAEMSDrS7et+PnB
Rs7UcMnxzsG95RPDOavZgkSP0+GBy+J31E1rnkB3Ium8aCyTQLHKCYbsQCj9XJLU
VnY8V6NF1Vhy72CXub/8OA40YatoxhEQBBVekv3J8/HBCmpSNeZeyJFSna7G7SA5
3SLjq8FORZiA5JaqVSD0I6cNUVZFQY51B5Opeh8cmG6w7teo2+R++E5VQUEDIdTU
7v9mUspiVPWcR47uL7XthO6FSingJQkns913O7HV81NSRiWcUFWwW/uizCKwOxeF
iKTmQL0LcYY7VeXiuWazlHjNt/YvQBQygiZ/WMa7HfkuOecEp4DXdRXQlCrQuLRh
ETZOaomlekNIcyNkezlKusdoVI1pC6cnLkvr7wipMQW8sUUijIM1HfcMxyq8xxk4
s3EWYnq/1ZWwHJn8JMlDfulfOJA38YxiQGM0KalCprW86dIzXuBqXoBBu7rOBGkW
hp5XUyAVDBoHqqunRu4DeQfcLZnzmEJp/+dij/q0UKa7/sEVNLOklHHh7/JrR1P2
KHl49wekMXVLrmkdb2WFesKRpyyzIEgxzaZ80/OTwKXr+ArYhPzb/uP4aN69knje
SUmhqeT7wbgEbB8ICPjdkDmLheY7d7kDj4opsr2khM52rECXxFEN2VETJUJkH+L1
YRi1OAXWd+d4ZG04+q1FQt0GNZlr05mIYPV0fNFwWREHz3ilS2BPCxkppgle56To
3pZZu2IUc+7Y2gtCoK3GIb01cMqA5emv73mnc5azehczRNuT10OXBH+GOUTUoGq8
tedVj4jt/XChbailFnnXpXuIALuMFVEu4mXIzp77uSN6gR2bYlFT+0YmhbuEvb0o
sGogumk8kFiA7zhHPYNq/3TZ4PAkbc8UYNrNkVVRuuedACV0UbTjLeiJxxP8mdOO
im7HpV0eraOzhq9L26aA9kbxQwS/TNY8HuudCCbtMZ/T+bd5loV2g+2vjD9vklrg
vIyTxSLEMf9IpxNroW2/NKdvNNV/ORFtjr1VFL0JSiurYDnbTzx/8C5k5k5xZtF/
OEjUOzXdY8cbfTALBEoHXTIM9UZ4B2f82pNqZmLrNIw9MP4EYCL+nSIa3ICvvqaK
iwHgPbX/rhhacj8TnSx/d9e/cFYll3PAM8WaFN1m3mlbO3Ktj0hAvuqv2+vZ1L9e
xBGM2fdK2P+N4eiz0LtCUijRYnnncKKmWzOCAXqCAvbMEZcirNf75J13JvKO57FF
X2vYAjkKdkkUlQ3pTbPebgPoDk6dEH7MVMzpZ8CvMLfd8lsYACxGJTlygci8cZSr
guDFniNpoBsByWz4vS6kJTWK0ZJiQHx1p0fNzOUUL0hcpdB0qxuNAye0eSun7wC3
Z84hDf0+JqaNXF5pC+PbdXa2cgfn3mRp+70tq6DBP46vHfDBgxoB4zI/8gy2oD6d
NJl0kO7LdZk4ewJ4i82WjsSEmE6LCcYfplrxh3sIOYTGaaXGG+yYWwiIngRN8QXh
abckRxjKt+EH9dAcoNsVikG8g71j1iqTKfzdrcsWooEWGzV8VGHPPmtfVUKV/lQ6
95wCn8BBBT7wsEqcyYtDAtKUa8CiLMM+FcOtTroPMixNo0NpbjyqyhIKP+qqzbDm
0kpoFO2lxeBq8OCJR8R+DujjUC7LpFmw8/ujqmhKzQPPPdiq3oOMdfqVSUMOufcz
Up06xprjb+JTHJf+1ih1a9HXHYPSy/MRaBVStTiS5MXoXljRfbNOXjQUWt2+tLH6
OV8Z7cp9jTJ0L2zQHKd5qySLtaajW6VLwKMO1cpC28Xgz/jjMWvgO+P9wwD+zhN8
v6Eg0u/aB7nPkEtGXWCLToV3Cdlaiva+9w0aWH5zi2PdYxKqdsNWjky/elvSetq2
2ex5vaDxZsYEqd8dUfsaw74RVgjnXLOXt5gd7w9LbxmwazRngw7DAwr21fVO8RIe
7nMmxn9LALvFtRI5oroIWyU3Fvg7qea1YEAaMQsNYd0lx+zRzoblvkAHyGiQIIM5
2jv7imuhPCBqKIZMAmhyAKQ4wQZcxqt+QkFmXAcX8gVI6nSL7X+MmF1K5gWSU39K
yj3JXuditFOQxElozN9XvS0n7RcKimX6uEc0T5v8kVQUhuabBTiXacUCosXXDWg6
26HY7hakjsmFuz9lrDHSjcfSlgb8K3Yd6ngIFD7ALeIM0GROZjOyKGO962zk8Y6B
NNSdthgy70cdmNBGze/uq4PRHMJdwfqbPpEP1FDkszLNSZ4iZhzlhATj9p+AYjPh
X/TFHfzzLawwYToTQibVkbuRUtJZb1hxk76if0NLK03ppTrL3bhZrN6A6PRXkmkB
9JKMd95XSv5FAZev0I4OTIiIZKo+kvIG9mCsZ0/n42AbkJiFwPWxvWC+BPRugA0w
uqTKdLi0P1hfBoa1lLPtYH89Zv1Dl/p2blIvr5I5erK2tk96ZqVRKZuIrzAa5XcQ
mwgj+8fMr9Y9NmUioe4IDUK3sHrkLlaUyuczgpt+GYdi2vIbPdbgobe0NljiqAWZ
Rrj73Rzej1PlNfd3CA3f0qxNrKlCuJUkvP9OWe6jOR0qb8sojXjYsGX2aLRgcn17
utjYd0lCm990s6KUZ0IstSwMwldaVRBlSMv2UcWspnnI4fV9PDFvpI/M7Hi3SJ5j
ZJS1iil7hK3v01FnJHFPXtFoNR9VtiFptvRUtZs9HB/Tj+7o6X0HqXpCooYL0QBD
mEq8KDDlmhF5OfvXfBYTr2SrIXLcptVbv5hYR7gu2paFiDivxnrpSAj0zc0WruGB
e3hrn/xTDArG3A6cs9RVdG77iBfcQJbLVBi20lMGIyy1o6zFGp9htZGkvUVmkNxY
vcp0M9SRTRWUS7cBqBBOcmVNb2Dh4UCREYcXv7I7aVJVxuRIe+470hh+DIeaqCxw
/tfeoplwNSUYMk1aKOEFgfbFfX04tmN0B5qpbtdTn6esVwmv80N8ADD9cfm43bVi
lK0XK+mKoOyku76HlzTttM3zx02hxp7SOgzgShWoN6ESjgk+aIiuiw7fWNjnAEAq
32qL9uatIQr4He9xzYbo4MaZGj/CP/PprvqoO35v4+kFFf3WKkOm4GQoRZg8wNo6
G8XtbFhVX/fQsDJBjoL/Orhfyn6H182welnCsNHPSDz5sDMgnCZF5NylNgLCoKGa
sFbefMIC7a9BVhGspMg4RQZ0ZaSAzxGo91xJqCRdlbhfVCTH8i00O4oHUyRw9O1a
a6dFqubG4xL/v1Jp7Qh3ee8GT3n18TOWA7oODlFWagcC2Cm1ERBz838/4zciQBxO
DTC38zaPN7uY8E4vTa2Rx5wNHhrYA+BDg9nUhNyKZ73HIU0VkCI74r+Y4wsfCi0G
u0L1QkVFq8aZVP7Av7gt8n8H7oM+QgutRq/nS1SZTMTnvJ5NsnHMRdeLMeT9Cp1R
pF6Dysgjt7KQjXsqVBN4o4dPPrKt1+wQNwkJVyAZTukeXfdMTcpH3tIqMLVF/kq/
oiccqpkgX3Ebbd+FoFgbrURL1BbWZ+LL8kk6iODdLcBhVrQFtiDfnk/0KI7PT2Df
ZjQW5LXotgRVe6VvJTUDAoxyvj07EhZyqkkiIwfqJqTWjQ6mep8JI7RTbcWXt/DY
kjFrf73Fzdk/Bt1xB+FUB8S4/j6KQg/2KcmsEZv1NP97g4h4vLFsKUw5fR2Pz5U/
bo2WvAmXCRBcmAR5CxD+mLsGdCiLth5JH97aqbqXYBZTtCkcVNnEOBbteYdeQ+sf
/TDuxrmIn10gCjkt6dWFINSPZpDIvqRgJY9Eqy30njuBBynrzfnccaiNl+calmDu
at7DJrGbvsT/TnwwEEgygHimbz0N1DMqC7p/97EnpmgxV/apNFCgk/pU8se/681E
6fVD7w2/HVPBnt4ahEQbxXERAVzwpJgB1syJPSADmXV7ewYZuSwy1sUX/WKBitY0
wwkQcuGEBfiKdU9QSNgbPc+fkVZEKG4E3bl2Z1aFdQsXYfdXDO3ndCo6edmo3E1z
yVJasm98DxuxOzMOW4vQD/NiK31NKiSCa2hh2aEuXpH4TuNbe+TNO6xQfgJngSEk
gKb3qOX0+ZsbrxPUw3F/x3rWP+M4FtmIRyv9iv3kOHXkJce/jYP1Tj7CgbvNxwMc
e+O3lfeQxwgbZkvlHR3Q552luP8YaaDu4LGK9s+GXzwNkfJ83J1zQvBeNmWNx2aO
YBKcm1fu8RgZ/zf3dduhpHi7U4G/MtbmyK0eqyJ6cp3t72gqx2ckzA1cQ7HF7Mot
1Ztqim9QmGAg3dx3tnusFCPXmZj/Qz+8p09MJS3V1wjlCg3wPLW6LWlWscaqh2tX
ePqBIdbdVMHYJBgTdOUJSqm3AwC75pWVVn+hgfnMHFI27GQcqaau7fowrGpxhVWg
5VOyXSBT6odFQTUIzj+d8WYKgawb+PwxpuidMCeijFVhM7zqAiG5HzWSj0VsY0FX
lyS6XsvCiNxrMeM2dnd4qlmu/2IWpCHauML54YVoDQT79AU9tMJBEDCoaJSVV+rl
d51gY8GrsBGJC4t2sxYBr1f8OqFTcj5UYxl8RGPAjGbsSF1UuPf6YvrcMdSSF1bc
+x+cQ6kO5T2JIwUMDyG9fxAfkfXRnhnLKTI17Hhx1m4bMHf9AoxFdIrQSEyoulFb
/j8alEp6o/8MjhFdbEY1NPI/pvh+Iy1b/+hpnz3vmAAgJQbliOE2tcgKgPQ+Lh0S
4nd/GLwkUB8pCJgRKEofDp2yzf56W7Px753Bjsur2p4JVOGnainwEX4OPday3NZi
p8g9GkGya9VP76EftRHRAj+0jjIXiea5qKoyV8wJBwrMIaa3p8y2ZtfCqnL2STg5
CWMeQlFcEa331rygZ9p/9hgQuVoFZ+R4PUfCHGnwll0vOrCRc8ISgGahimqZJqh2
Eq54qfhtk0zP39oMZIgiiufmcmI92CWXdxORX6OoPKi3MrbQnKmsRHL+V7DFxJqH
JiNw6cmxxOm2otQc6jXsKLOl1h6t2STXsvsSsq/s9D/p7aiH9hxVdyTwfpy4jqAa
YiVK24c2vUpgFhNGXjut85bJvObwWrbJMAl7CARhGJTw4fH85neTaTxnauA4PhGt
DR8cTgH2JAITUWllNNhwyAQr57ISZLlMrbjuTZhcgyAUj9MPs3JB7GSEtyFQv2sZ
AHW34yQpIvTh1rX3LMZTjdpToR3LCGRVGHyG6NnPcWkZAoApaJOwplQZNWd83qfK
veI2k0STXc5jOlhnq0rUkLtmdtHB3TXGKIib69Ugr0APEVpCbY5KH4fVNBUgfGQK
8ES4HMNH2xHPcSdaXK7CvaxIamVGgB/xkQqbsF9708qIR+jz+eQWLuHfV6gXR/O7
qKgBOkFOLP9+Lk+Uhqq4TwIATVX75M9B7gvhHSou8nyH1PlU6WhtCk3qQ9F2PVK4
PbmjM3axZ1nkRlaqgfXNqG1YvstwrWfIcmmIEE3CpaJkDb3AqOlpa9Bd3a84lwf4
J5MmuUKGeLOyDhSsxLZx6E/2TBe9fAn17fsXW7fstRvIa2wsRxYKqisxwmcurGfx
NqkaoowRXF7A8GJOVSEmTcsqKAQjUCe1ciD7SoQi4JDvAOF/QWo4HWuuj21Sy7In
gpRZyoQiU+n/V/rnHT7NEptfKJ9RlcmJamGkIWfIBQfvnJrbhXdENx8QGXVbtFpc
BfEFBgjtCZVOG6hZLHuBu5HZjY5W0xQ/ory/Oiqmy9V/8AtOc4PfuxPC69DS4eU5
egOdgS/7SZvbCecCtkbe/hlWy5e5NXuzZFDmxOSxQZMc+8v1sUNuqiSZNhlmiFRq
BiRBGNVg3XDfszB2ysKFRzD0KN8feOsU+LSPEUW6e+iIEluRrCkP4+vXIr/rv7V8
WM3c7VwlPWWgRrdeyhtTO3bDhqw/DSR5PLWB+FQsgefz/hOO3fFrW+Ic2cDMe+DS
XTy39WlbZC67/DqX5s3pBRGOxApW+VlHcLmkfJUftKdmbgJm7bx5aG6K5wkDva+I
SbtUz+umJAuUz1v7Op30zV3O2hUyYGvVGOwNQ5dfcuPLQCr+iDxqxlmwunRjpA6q
6QPpidsL2Klbqs/2LJA1n/xBQ/ow3doVnwfejy4OlI112GkzFdLczfCJxqQ1+x8o
mtf8Utsj1+JEbOMppkNhXkTQaAVUWap+vDdCyPX7XwHi3Axn1LH6LmCe6K/+w/G7
OCR5EAqYS4U3JXdiPKTDK/02/NhisCcwC72HY6+5vxXfYni7/RUWNoH0LCp08jvl
IaQjmIKVTIhsQeFuA/AGbIPKq4WM4QbGyHRf6daEAgxkVzvMU2qlo5pWOyHjRSqo
6nPHBuUE/2MO2Z8wD9gDwO9xGgt35JXkzh8sU+id3VJEHLfzCluYbnTGKILjE0OR
nXz2sXRdBksYM5LOghwe7CK2AVbE6dd6x/fGnMebIiIa66y4mQAgCESwOyoEZlAb
OKJECrgeFMMTbPKQf517dmo6RKIrP+FhK//+Iva2O9FVIRFPBjt5aUAnZlTNgLlI
17PZRhMwGxdXFkO2zedJR0w/zqaUsKqRca+yO0JHFxcaCCVIVXPUwYsLi5X4xoX0
Gc6C9X5dnshUPdf9RaeiRHW4o0Xn+IBe4gITRpu3YroFk2gR7fiDoMu92altfF+3
/NolgoDUbCrS8X4szteUrl+qrUVG4B/SeQVbk0vgYwniRstItTzTF1m0m7mYDEEl
wFi9SPe61tE4dzLIWPoPAoRWOSSOmwF8IfemOrwJEH1tnmyzPjfubdO/KJIO340C
D64rl0luPnJvSAJvo7y3xdjRHRfuFETJMcamPB9oYYoFQJ7Tydzzn69ByABQ8Gy2
IEWI/EBqsVfgxaRjwYnGab0s2xTQ54FwnsmuIN2n9HHUVCjNaIk3/9yCkogRRIHZ
HNRdzcEmeMg55OSIgeni1Msybl+QC/WrBcfdX0G6tVF7TaOTgPeMr7OtOlLW+30i
PGSjEUhAl8n6dhIwZ1Fh3AGyZzFgExOJDDdOtwJGXHWrW5HcRaBVGL79JA8JSDn/
CzfHvGlpKrzT2y/mEGeFKRhEVA+1Fcpk+0Vc6qzTkz2yUuZITA2Ln5FWrCPgn9Zd
hIs406YcaTL0upl3R8T3VAJKRNHKamZRpxaIckJiAO8qG5JFzvOGjJAGLtsayjGB
QolSlTc3LWlGx58luKASDh9zf5MF0st+Wnt2pgW1lMeAXCX0bM8vJqCQgpD6pvi/
VQq7raOJYOSgWMVLsImmDgEMTQoJ5jXvykGK/DtiLVSVvZsvbz7SjBHXaoakO6AR
6Uzmg2wjW5XVDVvlV5s2xo1U8XTVSPTP6kLpvh+yIIOmPb+CuMNRmS7fN+hKH9rb
rIjkVGB2Y7LYg+u38Lyj+uc8YGK5TO0m7n370aD8BHda3EFIiERxInquMKKDzV0y
5BkjfWP3jaDJiHnG0Ka65f6yPlmf8PvnVUeBZxrI3/APNbdXFIUm5hnC4QyGY5ev
AewsrJpJKl8NJvH43iJXh8wXOtPWvMPTJkTNwJaMD0uEtU492iQW2nq+k+BNHH7/
3lmWmmTtjsr20qKiI/FZ+d6BekwOSmzUfHWfFKCAz9eqbijUfc+b2vEDEcKyWVSg
7J3PBT893ykDDwskQ0yTnp1mQ1lUJLZ30nfiPzu57TjJ7Glg3/sOC7O9d8edkc7c
6BIA/nDKZU0uGlgocXpN9YQgFHEhn7cBekUOEBugOIm5utXCvoQIulE4CAqjSnP0
UvSGaCmflYLujfh2xgyWwx3K/N8iJhgYhrC3l9TOPPqtcjft+FRY4EPec68W81Bk
NzYUqLFsBY5JzX5An23Pd+stPrxuteIfHLSYF5nqX8sP53PTAfTY0NINVqID19CS
G00DUGijxc4X5+8Le0vgaggL0C8rsz9+T/6ZpPa2SYj3wNFOx3nskB0TdZPRqRyo
LtEWZEIJeI0zxmVTfKTwYpOLdvOw5fjy5SjDUTyTaFV9lMp8miF5+MkTg0HlrIIz
REvdfWu4vHppOlCef6gMaFcTuCzaKPBmPsOICPTztY3ES9zcjeO9QT71eXcSauq5
xDiKbgU6kLG1FEBBpm106fAUQKk6P3Meh3293tzExhW2se29kpooN5LWwCu3fblb
a2OnGrtBPW3L4jdHEJuSDfBgejoCG7Hj8wCJAHHd4Hc3/seTTAvfDAarUPWhmo+H
sNucZ4tVglaMYDUxTSEOy3w/ogLeQySlGzGs3I5F7qTxZwhTJ3LQ38uBRt6rRig6
I2b9vzk418QY88WslhE0dfzbihGBx7qG1M5UJjw84UYD+nAsBG6009VMKns0BCgL
ZnXbOsvWFVQMvUeCCZPku0oxQfpKUMSE69cGKQG07jfJQuAYaTyKNNwFlwCWjY9t
AKQGx8WIHB9YlMjifrAY+9FaqGthKpZZOsKJeUvBTMwTGKuBZevkzo3UOdx23tav
MsZy/Jok5AyaQoReGET5izmX8cqutz8Y5oJrOW7Q0S0Pj2Vagr3i1BvIH63+yvOq
bh++Q2hCQYfnTqfV80GaJN8xIbCYrbs/kWwXJfYpFsCUyvAvdsheoQnZtVTSghO2
TVCpXf3ouZtlETWUXcP0ZVJLVWDGgSR/tvbwEEuU1mJ7eXlBvYQZgqvDQyhPFDyz
217sOSdCNAu1hLcotSCQvIb6+WS6C+OTiZngeg4rsqLHvw/cvzmQ13Py+8VviRZS
1MXpb6/zSTMj8IMDHdOV9soWb//Ddsjb7Wk61LMtsNlLkHT42IDJ/ex610EBpteH
IOkMeBSiiJtG0v5UTvim47SPiuStm+pziaJQ2PH03+AtE1FYm/a3OAga1CS9bRPv
DZ71hhbourfJuRKSSLqc5vPAXobm+WCPAVwGdwRx4nAIQ0It/JjGiAQKoNiBkPjo
5BsrYntENqWQZ0nwGFNEh/s8Y6jLjagIu/5xprRWBAvczFdaoY23vjJu9JWCt+iL
cROT87jHO/tcLjDsMqjKk/nZJxf3GJgbtfWmnzMF0o1/haUpUeiJBV3NZMD+ateq
ZIBCsur5YQzxEYF8XWwFQ0k8H6HradefH27sRZ5qJXHeusCvIRkCuA84X0fBHWxY
GJ4NIsg/d8XBWiq19ZB+3Am7nMlYSCfzRZoT8oMOo22aRuKyYrPpKIWOp7dl/T0j
yddLMvm32t7J60AV5ilfgs/ZiLbgwquG6G2Lwtshj8xhEM9P36bQ5HjbOb9vlYnD
6wXS8Ay28KcIN6Qz0jp+6noHvduGHwujHvUj2itcHPKnjj5zAecyjWP1Z5aBi+DL
OSLZRlJ15E/dBNxUd4c+HLGUXL4A6g4l3GNRQ67SDr4yppLpGD4h4kt3fLyHoLXn
wiEas8KnTkbV/5XsnHFrHGz8IpJ07qtAc4pPy9HY1e2MEuGXFe9euRxpLmG01pxe
Kap0rzXBXrFJKxIdUp+bY2U4Y+K54EisHNLiRqZHIahT9AZlNEVZtZnOraTF7HAf
kPFSYgmdeg4YnORyBCeFmo2Hzud4UMyYdNZmv4Yg1WmG0gA3nLP63Z62++jhebrv
ojscZHOseGFqdjivwbt3s8h3z7xnTe+ZRpFX/MDs5zOtRAkfcAyCOWQ9LVufQzNs
I04mZ2J1ev0i9RFeJcOMDPkftrLGtVtY8HCB6fpelL7jeNBaVLNK7Lf81Nq3QQ1u
kjPb52nBKdIDSCYLDNmfqrUKOc5onPZIgnoeQdZKqx7DK4BqZ43gZHLax9M/UgT8
QeEESCNsMcScOzyO5iMhJaR4Vw0IQFaoX6c61MU8CZaGMI464UUBqzPhPIFXYQ2N
mB93gqXh+9q7E3+ESKx8H/7eqr5+N9616GEb1MxtmOqR49bDeYzE19uWWs9Nar7v
6NmVbc7vFSSdOvQqCfCMS5FTPANIbUYz0YTxZP5d6nnPl38v/21rRRqkPPzNtlb1
KFit6cL6hbs7jLG1euX6yfVAYDE7qHPNEXNpWvg62fUHvQ180hXT+hukUX8PxY1S
46hMCoh29Sc/opmDCDMTVmCtr/GXk8fdWf2F/HuXLns0S77GsfXVmuiTnByxRzHN
Jjfc/XPLOeZubbdGtnYz9brJimNq+3wPSt0FvSEnqQMuJVxY6cjUzZ2GxgjLQsjT
+OVLYWZ1XrSb1bXzpk4bP/zbopTn/Nxg6iDrowZKoUtKRyv8fJNLkjOnkUf1I46d
VCToqAJqwv0VJGLvzrXRGPrbBIMjIFyeSwUK92Cznum7yzsLJl8UbKFrfPh1zS65
ggEHXoNF8gIOYWwxt6a5soqngxZG07LlNIO87IZDAkBC4z+MNGjsKMAtCu5J8/Ew
CWxZi2lI5Z+Qryh/zAa3iSE6eVkLUtC4E5/73AkILgBncMqphaNzSf0TM3DVqXto
/kR+2ThoWhCCP4QrfQ6V9C1ZqC82xZ7eYziKBQxZCYvEBHHM9iQ3bJanCU9UYEY6
42zVnEeKdaRAqK6JFLcVJRS9lvaYuRbdO4Myoj65/yzLQdQY5imJfdT9LDUb6G6d
AeWnfWZLX0UYpCT5/7iiDXB1+Q/S9KB9CfM9QhF2FwBa0wNT33hrik/md/YFUtQA
uwoJnCaVXnEQR79sMkCp3neG/Q2TilFywj7WYF95aZ4eu2mtVLjAU+0XRq7KayK6
7/21rbGa9JbI4zWBTV2ZHc7+LPZVLI+Zy216TrrAhtxaJvR3bm2G5GTlulgkjAsq
NrEUSMjmQw2Q90OY7tGlsGNkYUICEzgCWjGGp5YAY9gm+klH33KGzWuVSEjHufzs
KTbyfcHv6kuYCM1CqgnfGmMvNeom6CEiM7eYIcNXAJESSgkNI7FJ75pRvlc45JmE
zP+fsiKEkfaFayz9GWzVfrvD2E9KeFkPdSv+G7MpDbr4Qk8Yp9p0PMIo8/UMw0Kh
8tPBDiuyMoDY40jen3dRUBqAsI+NIa6g5iZtmUgN6NGlF5PPIEJEfZL+cz1nzGRV
Jy8IzjIvGrMs3joY8E69I3nEjMgsFj2Ly3+4yRIni5RUX+NKfYgQjriNf+jxealO
9XDXxs0+WDvPl/8J/VLcKpRf6Gz9rnjipKHl0tU7g1UMNuDa1oP9gcylgRii63df
8GHVwdkhE7h/XhTul9YtNVPfzgVCwoDSJGu7UWZjrBPJOy4nwOYX7x1veAdVORTi
HLTU+eNVYMqRx5CZZPYpU2O2d43w/Gq+VZdtv3ehwRHO+d9lfQFahx1fpIuiY4XH
nRyqa93Mj4lYJFyLYKIWxwLI+35dfoi4BTGFJQyFAQDHamMGddUSuf3DpC6SSb00
rF31grk++bq7kAieaC+WnGvLpijKeWvFIZS9kg7jdhuiBRh7RS7VLTxnvJkx+T7V
T8HEwatuwE6oo6wl6PkdQzPcVZvw5044pGz/+hx2pndQ9J3t2VxaMCJ/V50SVaHi
q9QqHDsXEfIDiss8Zp9+gr4v5KsdlxgPrs2sZ/x0hnpcTxQqFzwoJhCBoAP6UZtO
S7VrtNdBRSW9hEomF7nx9brostqh9QUkWaRGCeBCwuCbKv2XFIDyIHznh33/f8qR
1wXwWUPGdWzUv6PUKuA5/99iQAfUsV2W5QG/WdjllODS6U/JpVwZY90MQbfpmPIe
eiPLQO5C0jugg5X9JLd3ZzgXd8DCZZi4Kevdl26Xhhq9ndKHPo2nop6NkIkF5unK
3KhCWfJ1zQD3pGcWyzPEp5Earo068bluh3qkmsrq12/SqfA6G+mHwvDgEJj99SzA
8IGzP1drH1qI4pFi2IX7jC5w7zrM+9O0J1qNe0uNI12TctiTEZKV0T+egaUPErto
HTVjbUC20xiT+elMjvbQ+oJrRfu/TjZtu1HnFzrHt1OOdJiMRODMJMQCs3dxXpLd
QYd+kP07BiF0IlUfzafRw2j5deBXH34a2uxOeqiTi2Kz/M2u2wTxZsq+V6hljP6U
2Zc0F88wJzZk1o43/v1Fqp2Hk18k/h2vglJmufwOcxFfYXMWvDloUo0AaQdXC4cZ
4td8E0uej9vCvdCXews6/LxU0BhKXuRirv2T00Lwv813K9G4nu5Pg2v7JOyfgmve
1H46I34EqjCbC+rEGUYpWC810y4F+NClEB7mGYMO027E0YzUoCDIEqhN1vbfPZe9
tLpZzn5+2kpPEv9HE21mc0a7aQcH9TisjNqx31aBlcZFFfz3SBUdCkqgkRlky5yj
b2wKhuznS74tNxZnWlaqlNvPeoM0LHAb5IR4ScarkOUtzWdBm08aLUrPrr7+C07F
fiEk6SvLJqF+f/vTLKqBm5Xl3h3E8AUiTAWD4y59Mq+4+3ko32+7S3w9cWWL2/so
ryKtPj6ToUje8F3EsFPYeh+NjpJLulHt+uIN1vup3tG/EBD27OhbB7LhLcna9j2b
tNszOgBpLSksV9U8hxG2W5xStVbwBOX8b5+S8vxxXcQtez2TS1Yx2mc2NcaUnkuv
5A5ln9Su8vPFLVLu66KM6Dq0DNdil4dT2zGnqYOfKH3Q8HQLaaM8RCSMm4ODOwYp
vVvmoxas97eqNreJkH74jCNVblvYwzsa5iySwLmRrLvlhhqkgQm13k4M7wgqCxgo
f/XdBk7ou82Hs/5agYl3tzzkN9B4zhkZe4uoeUUQVl5Wm3iAZcTzpqnQYYuVTT5s
PqN85MeFoHeq+4C0gGi06WkUhx04G4UVgcCJDDMD+n25pwPPyf+K1ibkobqbhMph
zsOyNi2FBhSFjKT7BCB28RI2LtacBm1LAWIt8u6agS9UFewx6X2iCTAz9wYSU+Nx
H6p0VGKWsmc6PfJKjIgHakNSd3vPToEr7Nzzu8o7/1KcXjImnaCtsuxe5TPysp+Y
3t+hUSeGO8s0M1/QosWw5TVNENK3wGzpgF8Yv1JmpIi4xZMuNTKu/pCYuinzsFk3
djW+Ef7+Ngyb+zCaMzmLip7EONN9KxwaHGAPyKM4g9Ri+WvgyEbkIQ17KIll3i0Z
lKrbhqGmG3R7tvfkH2NgftNb0tSgSJD7Jlvf17DJAPTn3vmeCMBDVjwhqX+jPr4S
1NM+I6WTHzgYFAwQNYp9cu/WoDu7gJru4HrpVrraC3b9YZSNQVfa9g4CKpzwcJiR
jy8Tfsg4SdL7pLti8dgLTEawkfDy1S5JrjjCJH6buMyrRLA9wbKzueecc4e973iw
kxzCjwn+OfZ95UJVd+ODJ0E17DDPyqQS0vsyiRiyjjdO7g1P58yLsW903li5qpL5
k8XSCDmVi2FGP4D3GYxk3O9SkPg+bN8jeQzqV90cOcbVKSmtn0PF5y0fsc0Ag3jj
35MBnwP8PWk9tJVDZZY94sV4bIL6BhSjt5n0O70f4pC70rNia/J3XVl+ZwzILFx4
kKhMiNHgXVihYFGe/2TAMshaw7L+nnwq/v3yHkZDrzGxmvoliiM6m83eeab2IxCi
7Ai+YWke7is8gVK9wmkqZU8PNVsq8Z96HUxVWqTDT8YdFh6RveTyfKJwFiNFJBt6
OdErkeSvm3wjMQLZVLeP76gfat8DJjXJkgvjGTXukhpC4fhWD7F2DPRjXeIf9J4x
3tkaelb9EpX2QRtxc2D5eQYGjBLo4Jrxj1mCiTEW3hjgPNPYPHSoIq8NBemoqR1L
ZxxPK+z78T2ttbH2deuBNIo1w/3G2AWdgxDfkBvqHjLTKqhvtzdj3Ktv2RzHbqpE
68me2bMy6XZCDz6VVHO64LLSDCu2LlBLsboXA+DnqRiMO3o4WnZzy+ItDFJk6hNZ
MhXXU1yaDwsj7Az3IFiy1UNQOWMDKVlXCDkCZatEevQTqg5syJykLUrMQ7qHiLBE
JAqqQaXM1LGeHpsLvgpZA8fyVFU3QMaEk5SNhvq2MaSLhqEGz/X2FosbEJsLyVbL
Mxp+640VVvda4xud7hKchuRm+5x819yMFFZbvfkvhL/vHHmsYbf4Gta35qwxz5Qd
ExgZ6UKDc4TG9wObQDT87i+qLvgPVw7yNWCSHFrlTrO+sYBwU2v7vBDMop/jRVOR
ISRKGRbYjQxa6r4j0o5jPC/YXuQyKGl6AIQ+JOi7ZgG1yK0tarUbGwCY7ScchFgz
dzusZmhGW4Jc5sKUO8X8xK0LyqcbHmgPVHL1myRHvm1gI/z/L3CaqfrxevtpuYxY
hMaRHFaymAg5M7Ks4/yJTig0guabzJTxIwjqg1XcY6fd6uzW0L+ySTnsziAODSv6
5KSKE7r3hktx3xG2sFm//Zlwh5+VbTAgCTXv0pzjIpgojaWz13HoUK2/K/mVq3H/
ZLDs3D/lvsDodEbMmqTrvocgF0qkexTVUbp8KLNRJcT/fJaUDF7wk9RkCmpOyHey
x+DDwadL/53byK33fs0+zkRwLMUwInYGv0s3AmxEk+e7MDG7yuJnlkRfIQl23NFQ
iaIr5OJCXCOdX8PoHudgfzJU75iaX4QqPTUMz4uYAzsM3xuUJQfDhvTNegjfj+Mf
bZ3cJZRy2c0gnA/Iv3NwIBQlj0mz+Q2J+IqI69t65yTjcUAalKYNSYsG9kj6AKmv
z/SKGCYK7oJGGGnJGx9t1YAUAYK9xiO9+Ph6aUf715Cl360Axn9M485ytyg9s4FE
P6UXucrgbPkUZc9gkylC2ZxMjDAUWsIKhInrXPzRcfQLlcMU9/lx+U/Kb1jzmqgY
gPapYq2xGu2omkWDvtH8Bmlwqt2JCAXrQ2iSNE9WflFB3nXoF+BYO/95veS3kgUr
Ji4J9pZdM8ct2w22UB9093mCoHOgSj/BxCConZmqC3B85g2s/RRUPiqg/g5X5vCh
nXDBaoLtsi3/1Tyc/FwNmjcJDJ/5Cp8e2dDV37XBSPtci7xgvH8rrAqo8XEE9kcx
dDeWsHiizOOTzUCv6VhYJO3ZpPCUCabMDQRFnZPXzc5dohhhPevBcTVNL1FpwjCu
ZqMljl2kgZEJMOYnO+9xpJDrMI4/IlDKjfO7Ku44TfTuLK5uEj7dBnDMYEr7P7H7
DZrv3ZtsDZyTmplQsg85CrU2KFyMJpPbPlck5o1C/kn1WNhTxCHr3Jn/coxOBEkE
0rLaNoaaZ7diT51inxq/UfrQQ2codFPVcywev6If8yF7PjorqlKKYF7lp8FXVJ5N
IOMK28lP20va0AR+lrfzi3+9944mczkYIaroIxr4fgHITHdbS82gGoN1lPh53dW4
txrvUjDtLWvXbWAeURFXammoGXz0z/LQkfgVjwwjUeo71ErW4yIAzwD+hs5aRB67
3RXAhcEv0oOjsUSdvKcO0Y2GJZNQb3n4b+vMDwfXLdXS1zTB2NaYNCJVRStO+0y9
zIQxu4v3rXdMCSfOF6BZKEoSZA+h9aIuRv7r1q39Y4r249gDQyzXcb1qoGXXhcGx
GsuzhDps9cFmzCE7YVuEGLaywaoW/J/62lEeWec/2CyH4pTyg3eBcIaqmxHKOqp2
a1rzZ4OxWEADnPgN3mrfnWZQLK8ewbrK0fx1YKM5QrWRNw3fB4uWtyqyHkQN5Vrz
bokOtIYQFerPGrfp2Zimq1JT1d4JVEr5iwTPkHp0Xpe5yLqBVOcfwureqhxFZgrz
kKdW3HqWbQFy29JfDgFPZYzjzxxjl/00GrfpiRR9vRtJmU1Y/uG93CiJ1zKYnhnc
cXZbkeK7IDqNfrSRcCxMeKd4ckjwtv6BoEl4RIPVDfhj0Nm03vN4wHlZH2XFmHGa
6JvQT+AOlcfoqlKgGNdKHK51IlDaFPrJHCJ/p7DM8fR7Nw6T6VMKZBe78ha24D2j
7a9XgUK5B7jt3+ENDiwYJImuUfsdfJLxiEtuNNFVqstnu8OHQ6PSRoaSpgd6R0dF
kR6S49PVF3tECFKVwWqXArBzNt3ZqFl4mOwkgq0dC76bpdqhUKwcOnkbJwAnbSzn
VbdOWHjUVmw5XAs4Q8UHS2uwHxoYAY/WVaM/Kqj8q+wHgEAe0VhGJGcjFNsMT4D5
Hj2aoeVirU6MBFh89FWVA+3jh6ctAZSNP1XoIXVkDfFL7SASZo1hX88DVpl1cuyt
pXmuI84wCzUJ/tlrFdSb348C1GlZPBOEQo6CigmWPM5PCzHPZbetq2uAzfUAgYIh
nfT3LaBro6vDmHaRtwFDek0Wp4ls5F/QPKgckbizcPXZP4dXA1PFKHyihNmaB2PP
4CmSilJ9iYoFN0+RKmz1POqtLyb1itjNebb1Qpp8LZNMCprfJ40B5Tzge0UGftE9
mY6K7HQ7XPE3gNu9ZwKNeX4N+L6gX7aOkzs7fVPpuKvX5JmE7dQGruvXRQ9sgpEO
wSuKpstYMgqrl/96uxqV+5Wd/O9eDdnTBNcny6O4vL428UfgEjx9TY+90PooE4zf
I3grkziohwRA0et3K17CEPbhGm4skEuuvuCfLaNBifB8PLQLrbCx4C/krf0tHMGu
cCKNn8WMwqT7sAfOGbMal21FdAgIOpVCXJecTuunjpnC57Stis6DTijwjuE9nZOd
oC0OVcF03hHfiAk43w0zg2ovpRMH6KxsSYM/J2sNxL3XtJKLlkrnBZElOdns/ryP
jgVHZQeSoFoCz8//Fl/Bu5T9XxDnveJAtM+3jucxgWy/c1l1ungmLcj1LvlSpZVs
BULw8K5GipHD3PFaxXtp3gJIw0tR2oQ9NaGxzVlGX/Pge7B7jzYhlCG0Bjti7kX1
xqoZudCuOGDN7VYCkE/ktngqZPr8DPQ/V1/a/koWMFYpT51eTb31XwLvQZGGCxRQ
/AFU8vdfNc4Yddf9fBrstruo1h2W3+c7BSjAqqdQe5kdHO7QLBlELOPQmnag7IMr
ddlnhz8ZYiKxcs/n40bQCs0BUIhfvvZPs6OdPA1jXeZg4o3d+ds7X7SKqtQziO8w
Co4RKkdcc+SbxbyemRNORaua7uHv6hLNXBLbzCma7xoUE6OnS0zrfKF02lk8/TOC
jZlnL4sYivDxARqrgPx1q0WpfO3wYJlims7m5EtO9/Vy2h1C+/ZrJNp3FfbQGgiH
zbyb2Y4KpyZXOH9Jb1kLw0iA997OnyY/Z7wmkadjt5WMOq0kAPKVC6FmpsGv8OpB
dK5cLYZhyLsL/0L88nWkboG4NTP094EY78NZYgfeZUWPV748eFRVvbM1ZUJTjOmO
zo4+XAXa6kRuUPoSt4zCAEi1aHw3iqG8n0EVPRUKOIErVZDPqKwhKNfmAAx/h2b+
fHfAEdzr0nXiPCADXDZbyFw9k/AoSY1TMgl4ku9rDdCYkKeci7Aoe1zomDR/qD91
YGH9usz86c99zlpwsX97o49dOHGg/95Nuc8lC5BDK5bGHuX5ms194lZr25s7vyDb
jCAxjoZI2B347oZOLiS6hfccVSXklKCLcfoOuXcoXh/LDV8ijoHrNh95Z4bE8IFw
CxfQgPksNH4NRwkn+zwwfa82zVbghE/XvY7q/SNMcXO87AYpmc03y9T7J5KR62si
/EnstE1c/MRFKoOOSX52ujYvK7VulsQ5tfryowJ92Mdm0M0g3gpg2XcPeZC3CA3a
5Ro6y2awfQ7FJrbSYxHpLf2Fpp/w8A9/oxEMsiIBear/0JK5CMeiqEyZrevjbLb+
I27/Xx7WDFL1OXPNW1TzmvS1G36L/UVr7XQcwfMLx+6WJ2avVb14e+6ZoAwvBd7p
9GB2KlKZxTAD/QZEB1AsbuVqxnT9UGZK5E1wMfQXqIQFMged/FqKr9tQyA4rzkKy
cYbwpFTogL3SouA3kkDBPdWeguGgLuuQySc/w3YZrdrFlGZWxzlYz9VPO43D8i1U
7qGLQCxE/FGrOBKtXdamP6f/07xlRM+/7qXqXGUk1D5ijAKDzVwYD/gEF35YXq3H
Q6WiXu6ZCA5gBFXDRhd0RTAO++zoJY1mYbZ/d4OU6wZMA3/YLmjqUT9C/rCJnKKB
Ds5zuQVvqixBHHBBa7j3XA5WikdHxu4KNqOBA6YbahgHDDOtvRlTmcv7gBsKNR5y
ae7N5qIQHl0Ds7Ze3lWKP4/aSInrHPrYDrcDecd48rplgk0epnDlR53FLIu0+GYY
x0P2N21GHaD5bZu3yi677HL7H4ex4QTU2NO5dVZeTb/X8kJVT1CODQk3CA62+EqS
1dw8Piuwots4VRmLvZq7Ln20fEEWymTs+Ba1aphzHG9+LRRpcE3zWSJl6FSi8Xmh
A02WI3iWfFggaQWdGnzqDBTemUFFI2A8q26WGqslxRhGsQg63XJS/5++82wUolfm
yOCJeu9w0VWkMy9vNtRwdpQqzQWTErdzt/Ly7AqeHzyZPCVa1r1kDsE/qbDdszCw
3I2RS88Zr7Rws0clB6vaGtyqPv8cZMDXpy2kfblFVrZEOYNel5K/606REPwWcN4U
VL9MjlTqeMk9FVg9flc86WbsAugtsZFlbbVS6Rue/wkPH04LDVByqhQe4CQVf0+D
2WWIr8WXk7LKvYNXRAPPsSuwU32Q8mR4titdBB4LFUNy/B751QOOdC57UG79zHHb
tZPgOWAkWUanVtO0FyVxIJXZUp1MsNqVFUbHLGWnrTLOxYipDKt5RKUe0Es25Gkr
4ozA/Ci/9S1aHqo8cRV7zHeIDl47bTzGsOuhmFZMBDlpTRIfC6h1HU4JMvtIGOWr
gDGUdaG0IPnoYQcQP5xSiFfZSvDYNIMJmXi+rmdD9vnSzgMqATr6FO4v2VN5QdHh
hi8+ohTTcQavdtaX4xvCQWQMgEBv4bMzMAJgbdUlkrPh5bmKDgUfsjPgYRomWhYr
W+VOjogqqrRSnhxsdk9gtAXf+jtNPH5VpNoRcFnYjhZIhKFv6qYb9kF3lYzRbopg
RI3GHhiycTVsCRjeQk8zB8eue0YBpYcpKHia+I1GgPH1PnErO60p3g1Wfu9PfCxb
c3+eyA+OaVAIf91xZ4WSrkh9fVn8fT7+h1KB01FZwYuSLjhjz/F6vBSMU9GNc74L
2Xug/ahEahISCZVoayu92a9M7HQ+PKVq1yCFRYFpGwrsWs+Q4rZVGwpEL84fbTXY
/XV1VQq7pEcpbANq2/PlpDxcquWJGev0d1rpqS/CYBSl+fQJWl1lHQfaOYn+CU/U
LcPUgf43hhnjwzHLNiMDW0VfnoEj4Gmf2ss8xA81yG9g5JmHuVk8fC07g/qYLH2R
nrVcuW1gnsKCIHJr/+hl+xwfaNe3W07FPs2VKjk0YAt46dIlTgsZRhlcqIWkGOi1
Rw0P9NNmUCmr4K7XhP8qif2ipDfVxW2kBn4D7dLf8Y+QYmUTNCfWefJ7jMuAYc4P
vmpMCj/kAjE7QxWJ6/GKuqqtBUaTH61dosZSCyGyTSgCUi41OWi+eReXuBhSHr9W
v2Sl3HgULIvz+GDqcyRoLbAtubMK/rrV9X9uy2qOPnYl6blxWNoAavouyRUCMJm7
pNKqc4IXUpY7/zLODdpbsm8PdLSG8maNuRa93N+NscWCbTO+Ty+fanSzFVMpzRBP
Nx6Y4SAAKl0DvunCmJvrK3CrsI+91k7FQdoGarwqU6Mo1CPJfzYmzlqiYysJkEzF
0sHTCB6mmcs+7OD4x4gh0o9ViObW0s5JzCEPPOwYq0/eQYywyJRf99Dqk/WyZlDw
9wQ+R/wvW/jhkwWuXgXJXXSBrG01M1m7MkJ1rzy2T7bjx4ujFKGT+oqduiJH1wxP
Ru2PlPDAcgfXA+rfWetqpfQDE9YwCnOvLLiEtfbTweazDLiey2oHTU1lKNpWjbX1
eva9lPk2JmCX+31DM2Br2/pu63+aC60lvl5tuHBXG4XAHujyizWjOuKRSPReaG6t
UE69q6gvGC9RwGfq6wI47nYC0h1zpk2yvORubdS9ahPUY4rKNPWCQYKuIE492jhK
Ew6MXm5qkrwfGo063Dp214UH+r898HhCPLGWBgZSNLyKKJoaFVmxMTN60i4m95BH
pqx8pl2d8bWseDZU3mwTy8V1oqFt7zV+z9CCbBiuhPQnxo1MJN5BF8HeFZ2/ir3V
1fdhufpM0ImjySwziAjfcupzHZgTnevxrivFRRoLdBtApQHZ9Ry6LBn705lM11Ow
xTkXM0YvIQCKQMQ75OKPv9rYjtaEXrW65H0VrujYVYwwaA8lQm4iwapxeJ4PfQOH
bJIl9UwygqBCbKmdA2AlOtvMnQnOpj+/TIQ28Svz7eCZtuglO6ZPxhc7pZvuWt+4
+4FT5iSLX29BEtuKQjBkhMMwnW9QsKuMXw2CbM2LPprFpYeHTnvCr63fr5BhnGvz
p5homdONLu59DpjEb7DJNFHTRcYwTPDi8tLZ1up0dh+Cooe0lrZ8U9AQ+xVifady
L7wbYlzTSkcuWu7N9gHtcVPf3Cv5sej/GDIymBfRydhAEmGeA7dQKNf4HDtBM1c7
9sKoLmz7B48p/9+fX+JrIt8Cmt+JgAV0FpicBqOLWqZ+tnkF/WP5UD/Raq5KVIVM
oxNLaHmWmDNRtBbVdBVZuH46EfSJAFvsFyA8DZy9+TqCrOi89USp8ILnWoOf7+1a
BKG3SBqqewMwwF7QPLlRECyKhFpQfSKpvJ2lmM/TLXgjzIkAZRIbvLvTdFykcis5
iemAkll9ILqmc4hhwe7hyZV1GswCkGYO43nHtrXchgzNthez0eRn8JalKCi81U6a
CszdtLlEA9NyOgI3uR/sh/qDONM/C8KSdcsU//QwUDc4LLsCzjGKXjnrrqRU+y3q
nuWEatvaY6mYU3FVNBUHZweepJHqVFhukHd5k16ZUaDQJv0Eo7iqLuahbfxD8Keq
vB1WJouwaKZYfplsWxKi4CScX3Vt+NkeY4axElS5+uq8kXVUDF31lELqNZxygntO
GoGVk/ZkVpeQuRjev1UBIIgQ2ionwNCHg9b1CZ8UWytSvyTjHVkiXTCi/aWdavkG
fmLw8gmOkZNy3y/yGelC42Ej4wQpa8qTol2poB014Ic87VWpvUz8AdwEvhzeFmvU
mSb8J9MpfkRuNhTwD6DSbfhGo3sXG9gfBW+5BRpzmQAb2Q1Xx1EZoCpb1JjW/Wg6
p/By4kR44uWS5DOaE8cecWshXjwL1AAaGGlRNZ31r29gKw7h1oyFF6B8wVmrOTs3
6VROne1pcLIsjD7vBi7UpVFX3X8BISNv4P9yb/3kDqtFDUvoTfA+lCgXIQ2Pmq2g
2ogeDbtJ8gf1mkNIcusPPAVMsWYg6soA8UNNmELiftXXlpXW4bGZ2iJ+wPagd9yu
ljyPpvJS2VTKilOeS+dSkLsXCabmIBhBV7jvFeFKGvSrZRLbg6bzzSeoBnA8k3bs
vWMA46G76ObAA0RK/XtvNMrt+MIWYXJKlp1LJifpid0U5NRAy5xm3EVvVg5VkTLg
iLpBDm3wm6j49hPJuu6NhjtjM4JgKJkZ8pixgQGUaQMELA8WnfjYINT39miA9iiN
j6s8SWAdRSzYNL2vG447hSpwWBHPsdY6uAztt1SSpsjiQ5kX5mZ3bo7odSOPjnvJ
CkSKwY7ta+iREcJmU95RoleU7gXuBvrbpgJLiwyJEaDMO5J/GT1lIr3dv3QA/MBa
pfoblrHm7wP+by8UMhQQtl8HpqgzZx3DbI03uP+VfZKbqipu5s4qbnYfNOj027Ja
1qvn+tkUgEZ+qptChkcEfAFqc1jtnJ1aX8hlh0YeqUTpZXgR38hk8gkhqzCUCqOC
wVehdpt1VtHDjNXk4K8EsqmxoeqpZrqEw0z38WgDpRs6mRuDcluCXFs0GTuLC9oC
GZ7GFetHe18YNivP3vu7tYRsIenZHVfEt0UkiBZ+nnYGEDtk4e2j5m7x7/PB675u
gFjS1ALfMcpgIiVnKPEmlLuiOUps2xWV1IkvjNE+Kn2WD5MwRG8z2JUrtKCQQWIA
i40rb8vMygdGGWXDSiT0BXZUP5Cp4S5kmo82zJFrhilcaztYrxDiY6YJkf+e78xB
HddYnHOPg2FoQ8lG/mIzqxib0K8TUWgXiG2r87DVSuPZsaoLS7FjK7ZzbU+AvpEh
4ysu5sKTpDfe9Df7FiVY+yD4ZydKqOuxvb/De6k49ovF6QisFy2iVUJytzdKN5oi
YwiSG85PKmleWm/29rYylQ9ICSUX4W4UL3aJ6wQTShmjQynHMmbeFjisC1drahK+
jObnU6eISedPmyitm9W3/yQ208OLmxObNRJJyu2L3BSVuaTLPAV40tkLQOuqjqTx
Lj4L6kHKGnI0zJ2ZIMdVpR372H6s7HvfeBQfin9l3Yf83mwxvM8C//6Tn+6TQ7UE
pUoHpQJEkkSPm4CtAciHZiJOTZS+Aqok5MXF1o93784DpatoPqpmPAQS0GaZBw6e
etvKOmMi+g+Fs80ZqXV0ULvyhmAuTSLc4+rCQRYglU0ZTljhJtHs+57Dtu+POx1u
CTOjiDV0JvC5K0zZrflms6mSvfKk992IFKYhcFlauv93AkLfXB8ZGB66PuozFwOq
1zemrHPsWzupPeDVnuHpoAhPc5DukeY8xYWQt00ObH+IH4WvJG3PjLFRt5eHYiHf
IR6ekQYtu1WJWI1Ii1JOOr1BS+0lw3lelXwQ02EZoOVfo5+Ot9OJWZHg50uutdq/
k+nC9NM/kPcxBBU/Ka70SarUDMrml2dzorIX0bQuUjuLU9fgcnDFkFuT/QVXYkBW
xaXvFNiK3aCpBYZSBBNfCtO3EkDK0hAWBiu6YlXdl4dpTJZKvZecOH/Ylh+Lxq+s
Hocc7On4ASgk34pj4IC+Y1PVHhbmzR78ykSAUjCOBx2SLIlx4/KTvqBz6HJWQShh
/bJIicj5o25OySizaPKajhSd8t1U0SkZill2iWaRsezjgpF41fkhB5IXyEukoT2p
dyoap5R1TuNrYNUu6pN6NnRcWpGz99BCU3bOFX3o+IfSkIC7GR7RX3edLdi6Gh6E
yiQQ/2PR6bVR3ovF0rKbTkETcE9Yn/XYl5sXkdrn9lH7DboJ/nb/8mM9VAaNBvM/
GKP+PTIf5CqvVK60BF7CQSeSvFPzyuqIbzLvnbW0M5BxnCRwkBufQpD6AAEQeP3F
9zhWXvqIIDsggJIUrb7smAdvJ7DvaZS3JMEko81XVmtSqanjUuNPmHxkUZUastqK
l0Y56ch1f0io/rPZiu0658Y95yzTSB7ixpYsSdE+AmJ7ut+b2iqalX2Vu3U5urn2
/ouD3WX7C+2BXZqaNIPvGoG63Yl/+7DMp4bKcewwBk70U85ZWKCAn/2cLlQWU6b6
jb6A6fffWHHhHUutH0Z1wVofpcNGXG0TNAw49rHjZeU3Fro6fzPDW5u6yKGlm/hz
DDUChr6u7JtH3BxZFNRkBpq7yMYx/INboIXWwTOYb2tA6XAVYR1kaiMF5gOOmD5l
R71J2wCfaGilaHey8k8ku5do38Ku3E5EApAJ8XIfF+EhIzEB3xBMSXMjJd6J8WVD
tmgk4GY7xS9two/cILBBYrvDOYdCTtnWfXmxAWmF9Ga5QeXsXP8iYBbvuogQnMqw
lS0UOcj+jZhNDjRFjk0MzGkngb081AArvZ9vciji23H15J/3YAeTA3I7l13cnvMy
LUQHaPQgzLan5B6ylrXhNcsBAwlXAMq7WUogaHyuULFlRqUyEspYzDBurq2ZQerR
Wpa0Q5AXBVEH1A2jUWc0am7ebZoO0KjIlaoQtK/PJKGgakOxsVrq7IgtfT4Vtu9s
nTQbHOUoIiAovfigJGS3sx4HoDueSdykYtt2cv27utX9Y4N3KEdNnm7LMR/wpZjj
fSODLPzabfVHS6a2YN6Yb8R07s5Qhox3iflDOVvUgQY6ft0efYbyxCIvjqKVKf7q
UrhxZhlZf9aGyVn9/5ufvSTt3aX52+nVEZhbw3flw73pQJ02iWNC85TFi3XV2UUD
eKkEgZxKnFdbydxDcHBRrdKHS2iYaRWAI1qRmmGhQopugoVY8foZard5/A7Opx8d
v9eQ3392TW/b2LvzxdSu4XliBjFOVTDbVV4cqNdAUFCQV4ekoQl9tBnk65vGZi0c
aaiAuo75j6BwHhV70siWNZeMZKW8OlUszhFUoibdXM8bQDJN6jCT6Mzm3eFcGWLV
FmmQkJj2GOwomsfE1nzATKZ4uasqmZQnoxHxpp7jnHHoVzUnKwO2Qyz+38aPsYNY
Lb3tVErcH+PPQqcK/ZFq9CQA74GmE4Z6P5AgJ6sOpGfUintczy2F7lSmtG8evQUe
hx31/Ms5XDoRIFK7YkSjv50FVTx9Qvp/jnLxu6Ol6zfEdfH97aMwxFGei/MfstUL
/HrNzpWDtNuiKmrhU4CzIGzpkZ4XLKjBjPTBeWfc2wQnh7gAFIDiXuOeCe6gT9ZL
f4GkNTOHEz2869V4RZVBHTR0ayM/6bmSLZ1k31Jo9T0cjxEI+RRb9PyI6PYuEFhL
9iKF3KLYQyqijN0nsZwwekp+M1Kq12onxLXKLBZ/7rEP6Q6Fx4Qdn3yax0RouWNA
4QHatl9c01Mptyhihfor4Yzxqj/EORoNoDMT1XcZztigQLNL6FWLGQTg6guJ5pbK
GR2g9EkF7KGjJkOZ494UJX7fwDb7rB2bFtuVFBUFuSXqh2Lz1Ve74FVJ22WE9GvA
B2fBIqi80a//61fRNlnSu2D/mrp3YAZmEQv6xMKy/yK2hpaJMdGG+gNv4md8aVUX
ESBDQgvzRQwoLh6C5sriN5TfR34bXsC+JgM0PQPOylX2MqNiuZIQ7lmV3zOt2qYV
clzyF4cqpBAfdwcKVfymK/RbHIstX+q800g6tu9t4+n/00TFN+gVyMcsLYC+3tTy
4HzueK0Ua2MkrjT8mq6VhecOeaJFB1RxMnRWerm/dp/i4tv+Lj5+iQNsiIVYC/is
/9zg4auyO1PGELFDhsWZFFtcvi6GV6EAZQp6ccYqFVRbtUHq2vuuyCo07RotQXmH
Q3C9BVNkR5FYmyV6sRYRKrTSuA9f5PhDq2u20fMGXaaVVNPmFUsI1oQJWDrDh+cL
nAYs/471p5NsOeYzptbhshaGwtWLPdEyR3791DvmEyH+BjyyBQlaP1Krh55nAgw1
YQywKZ3+Rnsy9oxpW9X7HeEBp4rH02FI8O93kDKraO5NcDwwGVGpb7sI7hHrXiUH
ECym6W7SC1t2yVSONB7dvLa+vz7ZksQYPzZE7rGCeteGkEh3MOcL3BCMHs2cNzDT
v7bIDgSMNJfrh3ij2P/+TWKz22NNHh1p+K7XBB3CyMlJSJnSCGHmFwhwMthdZr+a
Dsu5RPB271mloaRWrNNFE+uPCpnMwC0NTkK1q6Oeai0oD7qAGgeQV8alO1tfRtYJ
WULt/9Stt7z/6xvCE3TJZmXqsIjqSmgcuFkeGL7pc4dOewioy5Jl7zMeHevmdqgE
HCopE5w2noiMCYq8YljFKYy7VnoubATD/k5lvK0mg/MMKfb9tp3G69M1i3whpZrO
/hVBe/dZ8diWsa46n0wF4Acvq/iqq+OQfWBS4p8WYzVss5d3QMnb5hLY9tg940Ok
HUZoCoS1JEP1lJjwjdsoEnzYdOkqZYG+cAYnJVJlpt+vGTUu/YxX7mYgUcqpEfh9
36FQd+7fpKUsupfdJONzjd7TrxEwVaV2rBFItrDzINKEXDURT/rtnB1JBdDV2hPK
m6Qs4l3Z2ljiNM3u21C+4R54XKFlCoNkqc5tbTXC33rDScc9eVKdiBWpxzmsbSIE
ROkVu6VraqL6VvUhpdvtPOipumBjFWdOptMb4wWjhhVpKGPJWL6W8a7rgfbwkBGd
/BnCHVpf3E2B2257OoCo86CWwUwHMrZxKlLo8XEder6L5bRD3qBWPAVylfKZ7IWp
ksx83KLwg4wApFGsE+AnmNd/9VO+Qei5q4Ervz/IrJbi9wv8LWZ2IZ72nbihpkEi
O2G7hrS9GXy9n/r0Q6RKT0VHeJJiNFK6Kc5VDMtItM1O7j4/FsuAKTTkPUiJu4yR
5kAT7IUrJFyoXas5OZzB4/w/KDR8qY1ZPqjuNmcHfQWk6MTgXFyaJajYY2cyPatI
mPbJgc4Mu6cGdIRuYYF5CHhGrnustKoA/bihp+JQE9k2bgfG43RKcW6cGsIDQrp2
nckeFIR3GnCqJmwng3fCEs4Zrl8OQTCgGigZI0Ctss6pYi2ctfDlTgTSxQ3/wkBa
FQFDdg00Pe/DpN8l48vuQxP9H5obrunC01axDD7cQ1UOKF4Z4qw0Lly4bbdgqldk
VZA7mLT5E0pNvnjEERtBNM/1vi2mu5yS1ab198tMX5wiv4ZAYNk1HVKX7698HSnL
R8fAZgqQcT8bwHM7tHCBPkegVwfszJWgfgFk2+BKupmOVTGx0E0Yg+hAfM1dz1ja
wS13FajA/ARpwVbpZSA3H6geVSweP9+MmwcOmbjaEtZy5CrD8FFfNvHeTBbkCJjG
iIa3/mNNHp4KvKH5iuuv2AqXcGiKIMfW3ZWrawmvADALNLxv36dnLgN4mX0/f1sq
ZFwK78q8WT3M4avvzo68hmSQmBgWoxpAL7woTJUj1Fjtr7eB2m31vojIfLBKwnUk
Q8NEkysG65EHdQ3/+nc0hEzUulkbtVa47wDTR5xbYT8QwzzeQ4F60VOY2LMubPWG
Rg/ragL9GYAFXEJRQdcPj0ZBx7s74FopJwm6EJrRkEGFm00eTJJ7nknE5gIQoa97
ftcd2g5/99+hN/RH7gUO7yHXOU1hZbGUCLcTXrY8V6av98fkBDiR/zQWxw+rKPb6
geHxRbtoNgmkzJgmJR9vGJdaaFwPeOgSUOWN01rSIc3UW0znt1xJUdLP85v7FnV2
nubloL+m1sbygMbzTWggEnohatUFDuXh0sAZ3O5vnUmYoATC2kb0I63NfguZLtAF
DTkWmaZCu6kPIUjsIwlPzV7ZYU0HiThsGhX+o4rCRQ3A4DIFsVifJtVKl4BGAHMb
pFEdbJUpBp93JKD0GyVm09WOoIR6ig9kpVUq+lqyj3uxNPKry2FROLIPAGh/j1p3
RB+q6cGg6LYoUd2d3Xy1Hs5qYLd1MAJWRG8HvzyJjImczkMNIcE6eV0lRgfm2d4k
sPOx+RB63jWcE+kfrKB7m20m9DgjibztH7rt25EVDNicLm/oDG52tvG+2GY5dW9f
jG3Bv1Eph/YCIjKYwIWUfgVLca0WltLrM7EC/TmjJGsVbepZHZyXYOMumuf/B5na
WQ2+/NffYieWkSejB2reqVi9R4naf/c8S4OTuFnHKNOx3FNCBxpX82OFyakHc9n0
ckzw28LYvpFRtkS5+vw0cI4pFkuwnMn1/J6ZIjctnWU4FjWpEwQsWkz6ZgowJear
GnQZf7j6CozVHq+xsJqgmGv5zYvA3zzXhVCzLI1+x4Axdur0ePMrUWUted+vmTPx
bW+N7KneO6z+mFnhWg871jve19r/u/DQ0Mn1DntLsbsW0HhFinL7kQ4x9p+xgjEy
+hTWehA9CHr/Fm5tGlANqPZafnPX02xtnJxI6/9LGZsm4mHx7NZCY9I/86xXj7i9
eZ9Jun2Gii3aOujWway7R7rb41ypri5qPdOksMsuiHo0Z0VGDgJRqEFqRGVp1JxH
VRXzKsFdVuPjjzHSzSCe2AtDMz1x1Hza7S5tsbNsLjsByvPVo20CvlB/Pda+V0Oe
9KpZEu7mgWm8WL/gNd9MLV7BF1U+C5kiezWOzeMh8abTLnKGFHYriCm1IUGP8GlQ
tWRcbmPCaYxEwOLv8ZTYglkG3WEvIPyRaTCoDmoJdomxDysK1bmB7UlPXFFVOqCQ
fxwPMfxSfv9BQGgfnX7CBrzVHfgq7RvkqBVg7EIEH36iBIf50QpzZHV19WyhcwIQ
K9KiJZMfi/OnmsMDZYtHrh+pWIAecg72cnsmyFFDyO33bK3rJOa5n5Nf7seMgqrg
2S+PLNCDt6kt0qD+uVsuyIXTaAFpKc2eE1mKutqD8cvSUZ+Ry2gFvTg0VjueiRsh
GdmSMlZvikZ/xZWVqI6d8UGXfc8JkM9GrN5+T9XE3B0VztECeQ52dysbrnAiSWzJ
/YU4S2Qs0kPYHW323rFb+0ukFdWrxhfAIyOy/5RivYDLkpkDvpAZ2u72KPC+nNDh
OAvyGRePNRzU0h3wivTQZsHXKWxOCisFt3CLAzli3+ZUElrLthrMrTDUW1goF/YU
/XuarElCrwA0hSvfnEAeoyRPm6dqLy5V7Zw6aOQxK50uiX6KE5GjGgYUNRpMvfdW
9R15e2qKYuOhf9hxqClsHdz0lw78vH5jtn+oM+7PPU+07KQrb10GLVmRTE9Io1BY
m5909ZfJW5JPDF2p7slVX7tWJLehJRVk5zh9Q5y1VppSR4pzkYosKzZh6nflXsiQ
dY89E9kgzec3y8KUGt489wToKpuNpUO8Xcyml6cE2iDqwtaFaj5gyslc3qjb9z31
Nr04vpd0z5K2m3DreXNQ3zJJP4W4JIjCn41e3S/JNhHmwBO2H0/JfmKsCvClqtb0
8YVYFz+YKVdcM2RSwr3LgPiKKDNyqVUUzx7QJKXnfQZ7Cff9UvVU204cvYTitrMh
peXVs0difCmFE5Gijv30wdQ3fwS4m7ajQo0feIkLJV6FZuXHNZ2Yoq+KgeYupgT9
3NZmWy5rzBBlNbxMHC0nghsW3YQ30WY9+S5+xjUrLL5pLeECTFkGOxjZAj8L+QUU
8T4R/Yc9sxX7edLZ47caf/yUSfaVCo//FjIaZlm659golh0a7hmdI1cfI5YC8BGy
XcbqCSgVw86wrupD74kzXusa+fYUkaWYNf1j+y1dO+Ix/ub7aIsxYTcrO3oVpBhs
9poPxj9xLlhWs0z7YnfpsnQ+hSRx3v1B/xbS2FTnMFzrPjeHFU0AxufJytI5Sx67
2dtjQGmbsJQ4WYrDx7Dd14wqMQ/flsjsqPWCJFoIBygVnDXLP33FUW+cshLFj2MI
nCWkn2nuaGSZv93uxS1Juo16KQcWWCOJOB6hniarA9rfAA8FqxxHNKOkZ5LND/XD
idkgWpy3t277WFpKNteDTgrOqqKFUi89cfM+fV2gdNSvfR45WZo228AfNFq+aKeY
scp2l0dhj8Moo6DYaOOH1DnhRAHda1m8OoOqZNd1ublf0xMgfgolvhDbpZ83bJJF
y5K1e7FQgcJEqfvT0MlPR/IeEGzWflnoLMD93kjZg+nV1esK48IYt0EeG7AnZ1DD
fNCMvGGx9xtcbcYp1+skMC7bY4bboc5SkivH7ykI2PAcZqa2uvNN9iGxjUp/vVus
hJV/RQ7UDk0GHgERCPOXqK8wnEQqWiBwDt/JXskMPQHboBoiYoF3hTG40c1LPmHr
xvZn3b5pQkN3cCL9Wk3MLIG3/NH+vr1pLq2PcSb6yI9in1PEduWhnXbQ4LmwBIlN
xTNYm8UT0f6+yWhEl/DhJNg/0UuhpMQQFMVic3nnOaPOaiOWA7ILaJHvGSmEhxJ3
Kku91FKI3JW2V6msCWt3Nk809tbkG3z7bPT0Cq361nXKKNpNX8xBEZKdYHjVP6M0
Yu9prvV1YGWNoLhx5CINOP8vjSzSanAiSZLvSGUNbP5dxVVomtcjns3VokPMw2XB
gUv1lBDJF2YUanEoEoYw7klP/4EYcmZG1dIXC0why7IhgCpeEsgbDm1pZcyIOHar
wsCQKtz8Ggdk/S+vkinBVwaq5kXAxWM9GwEIK8YWQCy0TnHEmDMNhtfPDS25jyai
NhOJ+uUrhzjMCipe5qS5Xw0SqZ1v01uawCogA7yFuQc697isT5VegHd8Ta54oi1P
SJHMn1p34rIWZEeW49UJTWLxgf9BIq0nYYJGIUkZm9Mb2kAqxTR6cLmumY+dKYw7
Ru7OHoUutCnmCoUZM3VcbsJLPrdMdUlScfKFEcKFzBbmjAvNkfXjKM+daFXgE7Gi
E5kZP2M9QcAELyh6cqwZGv2tvHsxyao+zIh4hSFrg5mpN/oQPEnuQqGF0W0CPo+p
HVTcTluLMoSsydvxK/QuxxMtbeATjHTKj86AKBdFJcrMcBlsUBW4NNJujbDmWQfW
+8/ptt20AMmRjZDSjzmSp5d34ZFIqhdrDp2BwxIVep3lHu09e9ol7/pzWkL5CKEI
IRP4NQ4yTmGzX/zPfs4BXB2igte6KclAhdx4uAOmSoO65PP4TgixJXnLUgmuuGlY
ssqGt15C5iGVVaAv2+Y2cFAZmBNB8+gcnEXfZv/9VuUa1llq4S8tKZFD2A4MTeeH
5rwyy8EM6Ht7DKK+cP+j7yW/9aJszY51yac8/30c6EZFEZHRpVeVRhbjsODmVawb
IfAC7Fyjwclk8+G6RV2TNQu5WaWTOzx4YOpH1WaON1Q+xfUfYjBxllXMaKDIOPwC
jLIWkEP2TV2dbPp9BoW3hvSg5owGMAHVqo0DEflhxERMTM/yzCRsP3HJtco9tioo
+kV4jpEARhG7afYtaPVvHv4zJX8SCyG0thopXrIOUwhWz5b5D7VopkaqKtl017ui
EdvBiTwsm3MIKqYKmWsRst4TJBQRIFH9TTcy6UIIEVmmwGVJLRXWBevdOutU9q2J
UDl28/Z/SzQg9WIrrzP1qa+5qrhff/mLi7E8KZK+ttuwV0lMkIkPUzjyK8TTj3ic
7oIf7XpAryKky+MicRs0JC1I31X/giXgyipFRcZ/Dn/uY3e+sExb17rnpMdA/WPW
kVBzCUqQTzHmr+NggLGm3riXOEifsacapy1HV5TU5hu5iuTKqOcQ5p08+ZmUKOP5
c+7vLFxDnH+dPUR8rw3ZYsqtk1wp1i7P//24F9+p7buldXx1RuEx1Pgls941FwHO
G8xT1fDpcyZM6YhxFhOo1eBzIsy45aNGZ7E3U8M8T8CpAoQLbs+p76Q1xzLjl4TI
PoyjXDvOHBUhehYyJws0FcLY9cIIBsbvh2beN4aMhwG5Pgm2DpP3QBdJ/yGGXPN/
WCLgb6+rFzYdOtE5brOJHgKkKWuBCe5t/EbO33laB9lMqxTFh8RBV9aJWdoJqY1y
1lX3RN8s3OdZx7gLRQkfmDgXKa++55J9zMJaoVEuNoRT/InC0pFCITy3F6wOewmE
I099i++qTt40jJqafpIEKrlcR4h+hS8LekumFwg6t2Cx9QvUglWLTEv/Tddvf05X
WJW0k2TLfpiy5a3ITMx56hjqLShNJzuV/+sVEmZ1H9o49be3wVtP7UTQ1nnJ4wa5
m4hExxBz8bD1Nky+vxJtqyxcAYMiSZd1TxT46OJ6Bv6TdNUSZElU18KmdpghxaKH
GNgppGkjag50wKmvmIhTP3Hv6xadcdReGDu5Imr9bU4/8tU5DtVRDs0CSuVHBZOa
fFXbBpzm9k4YSM335MU9zT/IkQALb7gXqB3ysnicLNxrZ36rInd6HAwRIJuvSOw6
aAVFSDGuel9M4Ten4GqkuSCDEFCiOrKdjCDlxebIpKI2S5QpFWBrKz7D61XreQo+
O6qKjPA4vagUfrqJ07EPM9hFJLGD8y3tak6YV7rFQQwnTmnwuL2yAVI8dcsAt2nz
gc4BVx/pjls4fnfXGBFuAbL389OcOj5eaPdIrMvdtqZw/oh+FO6gahxsh7wXqadh
IgBrLHGW54rI/SZaxRq/z/LKxWDUfP2ryHbMKUvthYS4yTPAvzm2IzIh+2pV89w0
p4LBhUeZGk3cvvEYUfiLuyexubOxpkG1BgNbP1EFqLwRiP2PTbiApoIAd7zsLkls
D39HoK3nMxUL5grc+FXqczhBRvRMOVc5/oM9Olvn7NzdeDlFOyDDlBMHmLnySdtn
LkXj+J3ZIl7lDra5C23GGM/np8bakvkr+wvrFkFeh64lzYR2z5VR7ESOnZhE18CN
qoC8wtMeCPN5CfmN6PMDJ2Pw0UgK807NJIKSOH6qBQpiBMKYeYAyd3jm2rBZoNrh
YqhSLtqCxZ4PdGGXBJ2u+knyr7WGDDJ3aWzL1hZC6f6GjYNuHQvmFgcMhUbSlJai
a0dOJprShaBFWRaHaGXJBf+ycxnRsVDfsiFHVWmB1Np9/1rCHihNvHUMcbFqVGq7
klIxV3bO0NQaFJgGkIphIzikyGj99U8C+rkRyMtnhUKm4ShgnpFGRPKs0IwKrX/J
NqvHMO1ngABr6+CYnJkoTpht/kYE0iah7Mhcrit1U2l9WvJ7XX/JVdH5cS2+G51W
/+c0yV1xZiDSNMvdy6dsdcUWEAk/uf8fpCLowE+OaLPyO9wNV+EGTpyOQebLBUWH
mRmJzBOxPOsUi2nQYQ4kHiPkViGM8JscPHhp21RdiyztwSM2My+XfKgm9+Jc6n5t
vl+K2zBi3Ql2DT9Zy2/o3ScPcush6crsyVgq5QRWDCTHg4MLMWD+dbUV2zhwlPNh
iwEijaaSN3rXBqNblkaEzCcaQqf8Iqbf6kI5/9rq7IlsdIb7O5pLKY04gCOydiBN
Q6KDNFxHY4Tdi0lZJUrEefGytATVRmwi2UmZgJHM+VwwCygxsKaBiZ4U9YIEWlGR
wX4jxnZPnQBUjUSdGCwSVnfGtn3mDdMPxA6BzeEmfm1NTYlbH8NETVE954P8X6pq
hZ7qI+wa5XwSIcoIDEP7GKIVLnHLV0hZft80Lx+RhONqOHHKJzV+tPXekD5Is6Pm
SzRCMNw+CMoyH1K+ItoRSV+80bKD43ED92JHE2KDPUSOmNVyMnZYvGYyQeEfI+/L
vSyaPpmChows5gUMev5Rr1I3j3D+9wpJ8elslgqFz2K3w/78HbSg1vnWU0Ny8qpN
YlBM5z6qTtnwq/V2KIDEEdx/YU62vB8Ob7SRs14at5y+WY0EHZLW260ECmL6pCwB
izvOHf8UDAXSNlrVSO+0hGW9Raoz298gwT9Kf8ikc93fuErGZDwgVS7g1IXWXDEb
E1k7qJ6bHMJcOKBAM0UAWU/a3Hqz8ITbGDrl6C8Q6/vSzH4hIIQ4rSBqHWKtwzkZ
LreNdvb9uzTZBDt+Co1SxyQdbkk8fNXBxay7uSFtOIa2WeJt7PyWeC4I47DjVVK6
+uEi2EI9JNvz9snC6WiUl4X6sVcYJ2rzdhe5vnbhY9WR0KUMQ9SoMYVS3Ps5Zxgd
L4pYsp7GB4uy4htoxxjLTTqKcXSOAkyr/G42FDC6wYS0e1pVL7lvjbMyb0STZPJR
AWwgYVNaorixueV5uJHdSW1Cuvbwgo6yNuyn0xNXLaK8D0dxEyGzjINIszgWx/dM
NJolwdrYgkfczJrAjeYsmhD+gbxTT1SLN/KobgIe7LNvohyaDqe/P2kWTAWXcXUO
pyheopZa/kB+iN9cEM1+5bqIx6D07wXjZLq1qqCb8vLEdVQnKn8EQ406fKe0LjbN
slXiVzKUYcMDRKtoIEZVVnm1YeVOR0b2Wpetj2A0Ar/y+FIH1+PYqrooFC4FLH/B
ir5qcyIP2AlQYp8oZrX/sVAtIYDGYi3H6sjwgfZRK5OBUKQQrjmgfR9mBSy/YoY6
QlgX/sUdzRKiSOUoU3VqSRpI7MDA+SgaIvKogsGVxAd9BwraJqNSMO0dtHnPQA96
T+InWawsZQHI3OiLf5aDp+XvqoBQVifOIR09Rx8efgFN5rHQhrdYF3aOyHhb9F27
wvEfVtAzg4aKoXs3DXdgEUn50fkEmwhPMuWMfK2fq2Zpec86ufsydxOt2AbdXJQ4
+rTm3+jVVeoxiLjazws0tiko1MDM3BRrbH5dVZtuTIhEW8vTtHIIOLV5O4jhunXR
2iVil/q5pwMma9Vqo+C+5xzpJtNg7L7WxNmoeA0+Izs0s8XYaP1FNCXyypJRAjdQ
IRiajYsUW+7+ygMj11Hhm6EOnnh3lcf9l1qKL2KnvB31QpYhyMr5zcpOh6NfTG3a
TpKoC5zZpfcixEvvT8I6WuTssMa9GTPbFMv3E+x+tT7f++5H3hrST7ZoEeunf7uO
pu68g8vzQixN04OsuFWzJtgUjSb9vnj++GOweaksvHVqIetXNFalimNeRZ0ClTY0
eBcCCkpQ0HK8c27zcVF36WVTSh+Gcb28SA6OZe2KsGIpDLkmG2ba87Dlh8e5KYmo
LPH2HqUcgARJVnNX5l+lxuqHAkibvORBmZ0W9i8rHsEOtHF7jx97lWPgL/C+S1IF
w10v4GW1xmcEPJg86fnljDaodKnfKGYvse6Tum1F5p0SXUnVQ9lwFpGs/QcMROTx
KEhelt1bmG96b3pwIZrYTTcqchrdySBuvypqHZbXagrUTsEbafY29ZhWdYlFrEu4
nxFcVzrHc74XdPxWu1sXhgoXlzbuHkxwSjrkn8JYOwBGNuZFWbRvkMrdsGGVEduM
uS3xFTTIAmMMtS23usuAgaOBO6EuzueEfedN6aPbAyJAtkajwgdMs4CH14Eqn/jc
vhQq5/gxdRbZZ3NAe7zTo2HDVVNjPDvPQpl2JaOmLy3PCSN+pG84TSzGP0V68jS3
KPcK9hkHfMuoKcTj9jeyZnhR92cagBmXUjmosrK2QHbtvOcsiJd3bFi43wXvwlqy
qYhEvWariHkWgPVspRL31qbroL6ymxVdwyjuqje+T8Lc+7BkVmTCpfUzqDBuo0qo
omTDBuvkPBStCOpf3QizkEdV6o4gdjA65nOh5hoQ7CHYjOVuZaWyTeRJdSzzPcBB
pYHaDExpqnZUeinbILtRF4IRlcJold0FfxOpMYEuH380vxrWgP6We1q4fHEqrAeh
ADE1cVvK2Dua9bmpl6530354Ywi97NBIbWnzdLsC253lyVpU1IlIoUgyQGcSyfsS
OvsNaaNBK3HKchAEpWXun2GpKsGso6OmoyjOh+4aCQEXbHy/AhtcAzstNMzFPAAT
eV+n6TIqfYFMGBBnHRKwXwVpHfSXlNErSVj8S7eWP+ZfwXlD8M+McQl56RCEOz5Z
NES67Cq8hYZ131NvOQwQqFMSXDSaceYnJUm0xGIW1PgtNyEggTw8J9H26G4R9ffx
LjGhViSAUJIFEUwWvY7Wkm1l4msBFMI0jvFXYpMjNLFJXMsbCea9elTRHoWDquxf
OEsTCyWp9qEUMM7GU6ODkG8UP1Sk2e9dugvx/QIeoesw26L4ZgRWXC++fU0k/KP/
f46ipfLIK6USsLnipvUFKP9bb39LsjFJHqy/dQFNZ4GiIw9Y+Xdvs4IKPERfMl4P
8vUmWAyt+jBdskeA3KG2qa3iXtef7FUmoOa1+U5NIEJV+RBcBxUbqaQMx8myMgKG
JOxnyYkjdk0gTL1yNxVevTsCnBfJcZ5Rdq8W6xFslSOWr44f2cL+tfPDgR0seP4M
/VstjonjGZTB5p5Z73W0aD+JBR99hrapihVYlWawJ50Y+3YXVPkEKNgj2rDMASc0
qiiv2qzJvxgqf6xGfnoBDjRk6oNEdvqSLjczEoCc1xX2HJgovaM1s/fLG8aDzEh9
HXDwrsNC2j7WkdbbG23h1ZJqndBCZwJEjZQ5+aU/kS2y6hZ8T6ec9OgmEAuONYgn
47Ys8i4X9OgE0SL0VwJsBzBNhfmPbE90iZ0FtggNRw/rXTuL933g5z0YJFLpyN8k
/yLSnWcbfkPL2KfdSW8KeCxcIcBpxm342Jm3UAwZH8+hgVcVbxNHHa0j6WJWOHg2
xzJJ8oPP5siMO8EkJHsiiK7gUaw+5FVCveJETUD0TYUq0stYl8Ir3v1ZUoGvchPE
H2ECLbLfZz7KkwWw+gNpKcA1cfkgPT5iXVlXCaPpmkskEt/qM7WME2R15M6vwwbw
yX7lNiQbQAiqLW2PxhsedxJGnNtatO0XcKwZ3YHWfAP8qIB/6iG7p8zUQGo6kDDE
5pPgS4FM+0m6ZcwGPFl9Ugy/pyhQKxpiFneSUc0LdOtZ9NtNjFRLNnxJBc+AkxbD
i7Q4mv+sA70+fvsv/DxUNS92d0Bv8ZlPLdN22+HZGe3rf9LEdexmijwo15YO5C0x
7tUP3+gyB88ES/TlWen/3hrqyRkqo+BKJrcaG27kN11B9hPgTjvJ7chkh+qSOpN/
b2fCf8GMQvZCFxn4Duo3yly5GyKWuqtFuvlwIjUUOEgZJpiBQgqzx8plNe33aSA3
KNQc3EzjbOrPF1NYCVdPH/6nSBFP+dhrKhZhiDIHDnGOjre5jHw5BjsLnbP/O8bn
N4jPlWU/GcFUjOnWrsdj7inHUqtzk+oZb9jAkbPxhSB6wiSkaSwinSfrSXpQlLnt
BFf9hZhBxs7Jk/LJPQFBLOx/xcNfLCS0zsr5o9TkzyY9AkUoyb/v8KcX/80pQtpU
0HBXnJobiX+OwtLZjQvTj36L04ERV+W75sETh2DrWdnPOv2ASeElb56Vi3wCHI7O
QlfD464zlVSg9Cx1gFeAUdf1mdU8477rAs2dz5c0+VuV+I7Ia/FbND7qTOAsU3BP
qYHPWCGvFY+uHkIZzYnw4Mxkx/h1MNMx1JBRpAn24braFbF94lxdWntmsNC8h1OI
s+N3iBmWPQXewFzdbLw+5KuKzd6PTGqHfhie2MP2STPZ5CjJ2D9+ZgKR0ik9zfVk
v7xtisudPCaXKpLDkA8LSIT6kJyIyupYLm2jJd0xlV5hRSV0QBPyRoxo01u6lz9u
fEPoPjTC29Bb7zz90IZ/MEubZfOwThSFttj3JWkQX/tv7sMrALN/pLHTbfiWwX2r
ZOYk1iDnTU3Baji+CXtS0v4Nda5QHsHLaMNa3ZZfl45qUP/5uV758Ly23ZWciVPP
7b8dSjnYL82fvSwdwGmCtbCTQYAurPKRXyMinjzuY+fanSnhpfr+UM5xpQ8PKcRO
44fSKNyKTguZyb0tVj6fy+DozIggZU9mx/VU8I3XsBYcYEzbRjk85yQbBfPA3uAP
EiQWLmN1/bh4KbKcA9bc9ur1ZjwUpSi7DY8yh4fpXf7Hg8GFQ9Ji3XvpXlENuaFW
2ApymTXD75DH8we3nGZ7LGJHzlj7+uCpgf0HJRbsivcIK3u9Veu/77PDSaajy9/f
ZXt4HwWW18fXpLfoWaHfFKaa4k56lyfRN61nJwcTWqlF+MxxQDGmlVagXX1Hl0UR
RbtlrCGLGR7RP7DLENfVkR2uO8/MNoXAJEMKY3vyRoCag54/9GVwoDuQ9aHVkKgD
UD2iuCG9d6TQtx6XL8g8ONP92qn/Ek6iL6td1q0IVzDB7NfQDV9+rDqVihvA/YMR
pRjOdQRD9E0lwudHMREoxHqtGKW8l5Yx2B1IGjODgrIY3Q6LQ/gK/lemwieWDLHW
Dkm5J3e3TB6n6KjjcSukVoJmfWy5p/a9TwF5RBRgkcH0R9uk9XCJMxh238Uu25sI
MPJPUuI9FZv5ZfRWR3zbO+QDRQNPcnmBUAjaatyhL82gVVJa2YbqNzG2vmptPHHH
RJJ4SQOi1lrwl37dN9C7XUgpYX3JWCV5ErBBt13WjcdF53kfDDplrASJ7OWRcOTk
R9qeECntaIAAhUT4X0cHLMJ4oPzRwsU/g2KKop/N6ajVkFw4ZKXD/2MpEe8q7zO5
KcU+7y1y6UB2IdgxnfYE3poGrl+xNME/TyEWUiB/2GUNtW6gpzbtxZh87RwLVagS
b5JWQ3iB1EZUpmV29+1WKHm1W9b6ztW1RPlECTE9jPd60ML1FpOFCc10SL5mTFZw
jGrTo9btLhJ/mNCnXfgdJUt0PsxlLUBI2/S8D44l8Ut7EcR5ERJCr7de+nVepTrg
1f6b23+3XU0K2FFfBWZli8tlLwS5/iH7K1B656IFhggu48sXrO62ai0xV/QyReBS
pN1FeAn2d1MhRZy7I69UBdE4WsUdtXbhVXIx4bDRxuaL+oF7TpyVBRrhjBU7BY9a
8oMO0BEw9dcbkw2fJIg7x4Ipy0qvJBlh0TCTE0ezgFJU552sId1yXhN69kKxoau1
0+Fk/sjVM9HwUZ5DfYkv6Lebz/ScwhxcPzHO5VzKUEMLq2CYvmhFkqH8UTzuKAvo
eefgqoDysjFIIau88cAGA6onorcd/WxlnaQBVyZVI2xrlnWvUseBmK31pAwvh9J8
WDwV7lM19fb6WnpnbVepKQVOPE8qGeZR3uSkQK5CAdhxYlcHWAcB5LwKLAxS0PKN
h4dX9kDXghsvYQe6i6+nTqABQfc6SxWs1NBWL4y6+t+blC+XbFbb6OaMu8WPeHtU
TwJ3YToShUPFcR5WHt9cGb2TgLJm/iMX4X+Y/ZpP2m2PVSv9YN0ioG2UBlXtuTkp
Jjna6goi4CqajXsmsZiaCcKvC/WEYYJE2NGbi8W+myWVTg3twUnwss9EH1wdV0Da
zpOJJgxJgKgYMMP2Zpqa5WaGwvgmnjeYHjuK0JwG2HTvKPLRiOTz6uedg+p/aigK
ZOeGIya3nDp1MMV9y7WDqkcWfa3q2RbR2jxSmEnn26t2zQlZ1U1wveRvSLrhTzrS
GTIuQGsf1NiobskOk0dBm5FivUm15VyWveLJAE2BIsTBG16bXhGN5K5MeK7oKRRA
FJr2RHDIzoLV9EsUR6OdLPazaWhJy3m2kWXOypzg59LhIqNVSIc6YzNBIvACJn3b
vwwuJsCqj4GEqnuEgZSg3ePVDpfC9ka8Rk6QcTvVjIj0cKzb6Oh35dVMpo9/yHH3
sgMuETet0+Bz8+uKRdS9xNISugsjn09uLncUlD3g0zuwdp+IE4nBYDhnQjNZ0oVY
4fz69cNeZDRmH+zX5UPG0vajB8i7dsm6aBqeVUKrwqMCvWbqRlKuNy/SErVl3acK
r30pt7zhTDkboMG+Jz/Pg7eGvQmGGk7MDxvX9Fk/LLpE/ZF5/ICE9i01nCn0JH1C
lZ2dQo9W6CjJPdDSpVa9VQ8FLqRlNXZyXAThK6LsBQrYV2eCPOVPjR/uQTKVTaQZ
ZX4zjHjh7xrkZpwxwSTF8PXjPI2YtJHz17xVoXUj/Tfpp7+iELTDundAsYvth9Xu
9cxuuRscTrL8M6Hz0GwHrXgtwDkYrFGDut/Xun8kSY6t5SdKCOeEqgA99OkEDSgP
k6epTTN6tRQpg8e6iChd4TVps/okCBmw6/LZTWHHX3gOEygH+wFsbesmWwSzBEYb
mGcHb8ca55ToaChKDdBUgx46ElQjvtCtK3IMVHfNmhR+35aBag/9J+7Xl09AWUdK
o8zMZ3r96XZoxthw//f3mxbwTs3lNAE2F6k7LzD4wl77tI9PCAgMB3v0jqJp/jVj
DPM1VE/IE0xALEQwzyF8u77PQK+vmFj0zghkMwoLALxDlkVIGL4bJTYz5WU1NwZf
dnkt/fUU0mzv8lRNXhZzF4d9lWHPRXPVobVhioJh3eFYniw1VMd2EQBTWMuIYsVU
z4LUaKW+R42wMQ/hACIQjD/iR73vswvv0F1hHhzkJEs3ZaqF2gtseZpdS5rvB7sJ
dfospcmsp6LQPpeh6EMXNzK0AR1/u6Kfob04fVLtHwmZP0/1bbFLWPfAXJbjNUDd
8ZM4/mibUoO3YJFmaGHTaXipScD2kE83MWvpHAlTzEA9XiY4WBh345gOofoY0Gjl
sl5bvp9xi+7Du1nSu+7mYJILaJuoj1whUUpGkxbGV2zxqWDmZrzFdHQ1PUlvW+mN
+cRSoLjOwJ04Ueo+JczLHpTnSxttWXK2o4ntlmDIwsSWdkcw7Y5Tn5iUNzEc21rR
ymeSlXbp81a2AEydVv1qys4d7RxFRNsCHxmFi8fT23SzXUIgy3n9k0eKvIoobXlb
mIfNsKaM4Vure/F0FTrYChVUfEAz8XnLGp17V6AbL23F/PEshnxwEWg29n8tVcnE
llsA3fkoZ0eGkdW1OzKtaRtdgvKwvICK/xuezuXI4udxEVRRhLKnALMD+yQP0YFj
d5r3gqLS7BsDKw71FUVoDlMfalOZ9PAOKgJzjwJFG1qRYnGdC7cmawVayBTvUDZF
kYo1nbWQQ++ZAH/XiyaEDl6EHxVCqA8evYDHXoUOpjS84tW8/NZ4F4lE0J3kNRzj
ulqYtOcNcKc56cLjndCOsZHxOzEOylEB/oHHt23LpGT+0oiNL7g43uwdW6MgpxWI
IRbvfONnvZ1Hi10ETD4EArOoGvGjpFibZ7V2oWilycfd1pALI2F+IlYZxIC/lKMt
VZstFwoFw8pUvlc0pIewqhAmrxGUWI5KKeVDKAFb/xX49cy5LBP9OrxpGblv1Alt
iLTHpp0Y/JEdRGz2ml6Yny2xvSFbjrsiQveaygPe8IX66JtuVshGIDUZ7qb02tEU
Jc4FlA/c9qAiygy5/jxLp3g3XMFHze6Py146ybxIcXH/L2N98/oLDW8JnldnTlgJ
bLkb027iGFEKcB0TFAhGWjMy7j+Dgq5zgxOu/mCOnAKSQ5cLL9qjDuy62gygU2LT
mM2gB8LhVf6eZrL3YdPOup5hUBhs3KtazyjFf/GAuhpD5YEdC6LCH5qXpAa8JA5H
6XHQlhxTgyHrQdk3AYoCXcgDpkKLVozvzYWAQCVyb5UAyOLQeist34EPyxJXK6+v
UZfljmSDy3lvg+AbQVjN2kYZ2+vvwGQAfSPI8zL1EyYdTtKjf0HLlX1A6lKQDyza
K+s34pGQm4i5qGlnIGFadh30Kop2OfjnEoxDhBvqDZIDG3Z9J857icBWYRT9t7aM
nRY2HE+1d02c7BcZ/t/XPTGDdDiXzDhUJu3YAm6UUaU32GkwVBAUtwLWI0iv2oEN
RmRmnOmRP6HtpncXGQK56KX3TSRDPJu3GoFIFqPByrcH+/L7/fQy8Al1rAm8aH2/
bPYXaD9KdLzOUe4U9pDYfPkMSucn3Tx0y8hx5JtIDxgVpEGHzXvNmpYSNTxfwYyd
6y4vkaRdEHJ35gJHwPIX7rZ454InXx+yaVyi3jWB0loBBmZu+EpKgzv2Q3CTmGJa
t3BZQAspOZ9WBJa1xeYSoOxVB37CypbWYE2f03ruqPZIReyQhDiDk3jld9QSUx3l
BTVCXHghZmxVvBGkEHC20zkSQTteKqr0uAmqsWMGr3bmcsqkfwYVA8Exs9QaBwIH
CGg979MoNlyCv31mI+0BJtPz/G14gT1b3oy1a6tA9GqQ9w8E4c2/NT/hMANvyAgt
BAdILdvFJp6EqpY1kooouOOXBToNv4uFrS53r49j4HbM/rk7YLr16X2MQdKCkZfa
ZaTblWpmOfHgCWltWi9RyjgTIRITn0lTk8uEcdR9lvVVh9kiDcvd7Sb0qtD6SdQx
Xq2sOhH0VyRmHwOf4rGLAYkqpOLfZE9Vki9pnTEBt0frhDyKwVBrsui8INIW5X0q
3tQPfjdUH+5FrLiJIBC2rni2kUOz0mjWILMLaCqW8cWLenncaVHeLiSDh5ntffcv
i1LnhYvO94+t47hOun/S/Pt3CCpr1kElIg4gUPnbV5Mp4RZ0Q1HntZ2q5XJ9vstN
SOi3zjxoyu4QJJpl+WEklzwRCE2zOfkOMHPBFOh28E2BxKqVOiBT9YH141yHXxgZ
M5bY49j5/b75CXVGICSaU7yhnea9T/lM4/kXIcQrobsizVRvJLPEnnuyYNLxpmyh
r0YsdNjS90rlHvCl+G1S9gQSXbz027P4/t+Hcsb7KyY4xxpK6RiZY9dAxR/M5S0S
9O3hTl9DBO6UvgXdfvweYAty0LCDqVXVunYQNqduE7LV7Xu/HXJ4kUysMfF3dpet
C1YfYZ3NjCOtDKBhqHBpY0D98qc382Y1y5kIECGKQogH4I0tPetmdz3MHfld/MbO
38y3uZ0UBMCc3fRdqG0LPkUgoqgFQMZwNR5PPmDCh+oxiJQYTokqlF+dyA94psqb
wntpi44AJhs9syQWBnK+KZ66SES98J1qdTCt4aMGM8olBtg2AEIpk0Z9a4LWQoER
gT1iin73v4shVr4gVBuLBPkcvBFjAT8degcWw/qw65xfF/ZDxvn2raoT/iAB/hec
lvrHqqZaETIQky+eRIcV4SdGaNXOB+Rz3mstDokTrBYRMt64gGV3TksDC6Ww5RuM
oJxsVxUbh7/VTz8l9T0hk/B9K834MfJun505hPmmh29lCyDjHdys0/3pfxHsOq/F
1LJrMclBq+zi1pj1CqymN79kdxgy4bo/thNvvowqi3PJQ6wW79S0sb8EW5k9poh4
w+M4tSgT+JNmeCqCus07ZPzCLU9YVAAv7Fw6omEeL9WzfHJVzpErI1i+Kzp+6iYV
+d4FxogJkExlNlceAI1Edc7Q6Fwu7Sh8QA1n3CQlYhPbKhU8/GFnwJJwit70wbBm
JN5xIdve8fYr1luXsvp3CF6RhZDZMdJLoPuQ8QByKVfldtc/zHJJl8HIYMOog2BO
uKftAfpwREeToTPenO3vw8fCc3yDdXn+OY9OgbAvac+lS+8vVKlFdHKTb/S45zBG
IW7lX0W4UFq7YbZNQTNl0cH6owECDXfAbRkgliAcXwCLMGrUQmX3Y2FkD2b70ua1
UQDDKZq6pw5MAxeERCfNg6vP/01wTv0IhoxEvTqEel2GRANLu5WFur/E70EhIVIn
QpA9+EcUn6I0juXGkKj89hrcY0xL1yuui8XMSL48ZJY8LqYfB2i7+FBxvFKW8CTf
DY7gGleDSPh0M2ii0vYVUN4hFcpo3jMGTi9BOFzNSj1pQLUNkCkSwKwdMTF4ycVz
6NqePjJkTazwSrUWdOSk9Ir4wOP7q62iUjzxG5Uv3k+qOEI4y8Z+T2oM2Msq++9P
O49gZGxba21ivwd9tPP1UxmxOTHt0qsrxtjqAWkT3UUPH0YrCPLYKcuJcXnmgV0J
ltXpzLaN0bpOyRZtyhQZwbr0geiJQYokA26aMJhHVmkNjPF2hvavyUwqO8mnRySY
/7ExrBNc1CHy8X7i4hFenBPRR8vhvc/236VYfT9tAInOkXQON+bOq24qW0cgooow
SxYiSpSYmJqWfMaVOOqfRiTR/gtqtFqrLXTWZQRyiQnbtK2iiAbhtzh4So8abzLO
tc0KyEyATgS7GaEHxUL7iELGoyUWajjjiwHhNK5lK0n571/3eiXhccqLPYVzaRz3
l9RjDzE4K200J/2tHn+9TAHRXYrt4ywcqUP8/T4HIyBns44C3Trpg3gOcdxrK2dA
ecLDSRJkd75oFC/QS51kbAntzk6lYErYu0Pq/GBZKuZEJ0Le9kPPxYhqvQMaAbbj
iDVS8aMZH2hZmlYsE+iWCq708N/QccUv15tkrNZo73GPyqSIgJOvRrvHF5Mtb4G+
Wn3DiyxWejdWSiOshI3GNjtiI3UrKenrxn1jnCDpAY9PdZJKT2fHUJ11B1EWffTA
Ya1cj52g8Vyc8lRqTw2oxBMteEVWtcFA6ZT4naKa0m4bJXfOL3EAWnrPybtyx1Im
jNOltT2yrSxay4mqLULS8JntVBefQExXEYfE1mupC6UNk8msPfXUo3Y5xFcf1cHT
G7SA7As/UykDqt5A5YRXNX3GTcCyuDfQsf+X/4Yr0z6uPIVh8hTk2OOa02CpRVQ7
UgrTR8z9GDGzOv9GoLtTmS7xNk0dmCYpaBiAyCH5z7JLrsSW+2Tuh/9zhyFeNbH5
dMikEJbKFYWmVn2fyLw+J+MaXC8G1frDH8v4L4gdQPLxwqDqnR3gHypOtXOYSJR+
xuY6J8zdVk9Luvi8Jc98ZDumW4O7/XiG/iCqgDw08cEPCqMuLp0FRYPNg/rfMO2E
rIog+oApJCdzWCOc05ogkuUSYe1cur4VxadXTkIrNNXQQGUwsbauix7kXp8PMOgz
8OMMYejlAlXmNXGgKhIMHc9izDkqbo869AMssroegCGCIhXYZAgqebq2IqaWBgVl
Cqcd1UlWYQnSe8xABj12GnR7c9v+RIzlPsV7FnWPWzb0riSfD2Nq4piCciAoWY50
WKSN3UTVJGwi69NCgQLcFmHIUQqVXeF21NdTC+r3h8qvEzyXp6lVT0yAqjLzYMbw
tNRwywdyM/zgpHiuiGWYXhIHdTPIYwOtZ9y8uNdJTJpmJqHBrx/u2UgCx0ckR/ys
Jrq+IdUJbBUQMR+UHNsAiB8x/zYrSPxCnEuVY4INNIdD4SfF7ZnHtrjsXBsXQhTp
m895HoD0/43TNT12I50eg5oOIKKzYVrod9FaIK21zMvFeDhBSf1thdZQTxdQeNJI
GNzFI0ci4wANsUcqOnp/csZnKoemxzMPCcieNUmB6EgG9BsbEfNkLACN3ysZcQp6
VgKVL18RO+6WMBIE5b6G0AIoL/qDq3QxL104DAAYFr5DMoiV/oA/wgkL7XDX05AQ
UIDQ0QVxG2StM4Eg9UKz+oV3dnQ6q0LEqf8MaV1LmyjJH9o9ObJaDFv39473XLj9
XTCa9t3KuVLIZETq+E9Jh9dZDGcGfXBq6z2UtKmyNV0jgpmzciV5hjRe4mNSAJ/M
AzhUKey1HBp5xUMK/sNcuacir+Sw6PicVcHw61Mux5xgiMjuYmytxn3LHJ2Dq9oV
fxo7jzBX+Bo6p1Kqkz9awxjt7/cOcNfKdR5HdeX4eLCFk8RjnGHaQpD963G9l4R+
Id6rxKk3f6+ohgAho4Mb6W4zSRP8iPmIJ1w2SmdnIOrmJaJF7P89lI8fubC87Fri
Y275PvHOVtCBqzjLnbP6RHbmetoa+999dHRMjCNFO5O+Z5CyBSvphajvqdaQuHc6
7mzbDMQZoSwzDWcPeXzY0N10Gp513M/20JHkvc4FEWgBY5jlPTbGb5lObr3rxAuP
g5Uukl9ep+LhQ7hlGG6GybFpYbDEft3kbpFHppZmpJ21JTGws1UE/nClcC47EjtG
ybtZNmobHTct3wGnfl5W4a8f0pam+090o/3bbLyjZgd7FpmjYMB2hNOGJ+RzhBaz
S1WlTnv/e0htlXXnCErS67PzyaPfGXJN8vLDvGikfVDB1BoyBapqGLiyBT3bMoMN
ARYQ3gu22X1dnCEU4jC8JDwP9iqoUO3JgA1KSuIs74N8xKxnSMnvezBJ6BmV9Ikg
PfLOu9Bhrhv04q403hpqARujL+d2lPIVGeCuYOdIT0DTtpgPAZ902CM49MGBdklZ
FL50kV7qkb1prAL/lbEpf9h3EuzouET4GU6wvCtyFoHrlYBwoZgDjN61WiNpZs+J
3RVTn4jUybRWJBe02GMTkm7iyDABhiHEvLQBpMHiuJpaaAeSrvPhoGrtZrsfFXjs
C32LePj8cO4BygnQWzgVbCFLldBGUdFuVWGKfWCRx8o9fx73Aa91fRu4HrhYdESk
BhlAz8/nZfm1wXsL4wS9jy6N+ASIkSUBpyvWuBfgMydCDOihrpCh2M57n3NUutm9
/fEFwX1z7NsBc8GYq/xMaQZpdvnIur4SpiAm8pHupuomD4o+N+TFcWVbu+1yvNtX
uZ6wYKSHpcXbXWXYNxl3pj3LnMHy7HO1m/fTsD6DujMT0Onvw5v46sxcGzP1K5pd
+gkemdt7FNTlx/niJKLtSTVI5DpLXjAQESQCo1+xKWwWPFQzmjqFCYhY994H9zI2
Y8u5wTsVKMP7DDKmKe2DNy9bcuv7fV4NqJ+q2t/4dp+FYdgeLYuR8XxhCPxtdS5y
DfOMYE0AQnGt4E4uQKgtsYqw7wtnIBYoZ7BLWL0/x1SDEGoKZNrOLmwtMYaHuIdE
cjToG0IBB7ZJFM8EOlO9dpjOioMXlNKeb8Qkorer5bk81vYR0guekt/DMtUZlpqE
nRuXfp+UQygzewsRTJ112d5JJCizNCzhS+DxCk2lgBaIsqywXapXEsxOBNOETvt1
4FKbiv/z6Jx3ZHtCoGiDPYaqHOF46+JXMTzbLkcaU+0BIBkGAGB7sLUkxbVT9FS9
6Tfp0dZ3pEYewbCBm7A7dxh/5U+Ik11n0HpMHoFbwBbm3HQr09ZGqKsM8xh591a2
oZuzGGixcue5wTcjG8iC0HscK/yC6PWn5H6A2pHUYGKyo7wkum2tEaYNUm/GVeCk
LrFESOzExISR8A4OslhO4/2LPpLYktNgaF2j30hPx4oYLn+p7pzXcxkL2jERDyRo
1y3G19XP9g5HFs8gpwSxenhIIPFwufwidQJAn2BETS/XH0+W+nOGTk1SPWPFXwfg
IWezJiYUmUKwXoqS/sPtnhsgZZpo9DDx8lXGDc0DsyCRGzm8x5snfp11QAKq1cM7
Ze57OlMNgEJQct1Ybu1yuwcOIOG+DPInePcmkg/LUuPdY/HMYPOjMxnKzgudmW1L
sM0Rvsrk1/Ja4LDqvXegflul0cVvXLmi4ktxrBo7VcYt4MbbbvwECqhelGmcY+6c
BzhqorNrwuwqmgD9qnEJTearWJtl/4y3pHGqxk/VxoxlZELs8Sx1yQxVjThXDxgw
JF/LoYwCXcGf0yusjMZIOyvZQyOFnfjvEYytBo5hugXNu0ITkLTWw54kUtYPt4cS
VPCEXRIm7QUW/quWa2HHLWeFMDY4vBrh9SEYwnKV4uT4DCxSCh3j/hCGRBpC60JT
s9z8rDxzBwkkLIcdCOUSH5rRmRZxx/2s5v4m8IyohNVMysFVPS+U3dJQzALRFLgf
xnzG2Bn3qQV3/6kcwDGcj2Mr1ZmtAVRtjfl2acQJ80GzWc9LchTmkO+lCr9M0nPG
rz8rnzCg3EkxX1+2mHSLvwEtnpgxt6VfPWrZt/gl+Nk5nGKCEadn6zcuQHGP2Vsk
INrruEFraQh3dQ6lcmF7x1B97/DNjQ8WzMvo32940qknGgTD9jCWdxCj7gbg35r8
afoPXcQJKsry6xfsZFw0lQhzWhNJx/jJ0JqJiSLOUlV5dBcgxVagLxqv9ZA4i4ZP
EYEi9W9ahZPfrPonAbAo565lVMu52sx2IUPagzPJNLwZV5zSRk2ioE5VK+pAqu57
sdu5cLqCWhdr0qdyWuB9vTznvz+gm4wFd6XQWpPCB2y21I3Z3yPiaIRkOw4rTSca
axiccJQUnsZIycA0v567n0RunO+L5EBL4KYjYXuRq4/bAX7YifKP9qiYe+NPQ7Sl
+Dk19JJbx1evqo9JKpjXrhgoEEFRNR4m4uxFUSHKWp9iFc8zxyNa/e/GmUNMp9cI
oDJ9HaBqZG2mRAhOf+30rrAHqHBE8XIELfxaoQmxliRLv3opxsFDVdeP4t4QDxGu
JjZpwE/KhIn2f58LLQIrbVDqPi+II12mjeXYveTBcuG9pDnhx0VtK1VW4PmZWXhc
GE9HdVg99u9If5HUFJQXma/ph39aAbV2C3A6v2nMUzQe8rTZC+cSzfyi4uxxpWSW
6cL0iFoVOxp4xC7QzpXEZp+VcBpdPDgM08rfoCXsznYVYKneHzYlt03CBH8gX9Sx
AsjEVs/3wUwzupcPUNhzs1jJ+tiqNcys+xsxonnkNpw0uH28y6pSiM38vQfcydTo
z9a+RrgtVhUo9Zw/PuU3hfQuir4TYvtv/OIxU/VFp0ue1H75jpmfvZSbDV9KuOeZ
woV9aM383SzQc/hKkLePLFTjTRxtWvpmUeV3wjQR4CDzbDkS/IP9gsa1OKlutbXP
GfrZrWCgoE+YMnpZI4cLybnZ24TUOKnQAU09SXqOEiz4ewia2JNTNhbxd7i+GBAV
/tmxkkKbMjw8nwaDQHoM0ykZdcZ/gWWFnSl43hYSGSqkU1FlVoUKZf05TEsapQ3T
Y8OcnBmKXSKp8NxY9J+7scN76GBoteeMnQe/+6Uk/Raq1hu0908DMMZ2vZVWrBrB
HdwDrGf82mHc6lJVH9MyILGS1ZjFevH+XPNjZelcTJMOaWXJNwQbh1GtiZGUmnQd
Yodq5ZqJkYsRZhT4exW/snkDB2EKmJMskWVbCSe4Ywz9IfnjSzuqCpl8VI1aMOkt
0fQxy0EsnzVqNQcezBtqJVx/m95lW+RViXL8AYXqiqslxVwQR5u/81RXOJ1plem9
H85YRl2UI57SO5dkV46PlBTiJp3Ax/f1Ilx2+ENieaRApsuRBn6TyC+msBI9zQt1
Ns5F/sGyC/OZY4hZkWYH0HWnNCDqMX4OuWb0bT+o/rITxIfS+b7sOcgcAOXMGsMH
fbMxnZ9aqHXJMMHxRxKOXmkrj/RnmO1pfftmWBFgUToClbpw30e3A8MbGmbUnni/
zfVvNjinjVspUc3YF+DLSIfEvLqOIvn9V6wYmtSMlMDXJW80s8GtNjGezGr6xY7v
ME26yJ1DOzXPd0Osj7lUK+BvQmxscTNsOKGuUDsP8USxn7CLWI7/MyVlaofVfBeZ
+x2txYTtsTwQPEfXeTyZzuRKeDjTiDflT9V43qWP1337vsSDSQqoxna909Ndaxy0
PhB//Mz+MQRFxgyvjFGvQ8vA4Rlg8ej34lgx95eamboMVFjEnEpHuol4ExxDjTmV
l7+tYXpnWHaR7TC3UBwVoOZMYoqVaICuE84/y1HYQ62NYAdtjrLcXaz0YupdkBMP
J/qIhz/f6azKDS/L1f6T4wRO+vtP5zW1Crk/3/pDCbKVLaqWj+b75dl8AUJjvsuN
1aLkoWIkiKaZcRSwEBzHpfHbS2g8C/Jw2K4wyBr8MXGA1gu9MK28DIRp8eGIRfGz
W9ynz158QZocCWIhLRIkwyFFEORfc2KnULPPzmGk95Wit6LnthuLGhMAaf3s/quU
cbxYDqywWCIZJLZbvXnBOI3T2BVcH3flR81/k5Reg1AKb6TCBuNkMJAysaajYCgD
MMIoIHhLVbUO+8yJHeVIXtAjm6uoy7aee6RLsl2egPEjyB6KHDys2/gkYXdx2jva
a8Pz//3YbFoWCCDIuP4tVKI6O0z8qN5/WaziI5Mg5GnYuFpFJzuGrBYAnkmvd4jS
1yvMGKgia1zb4oezRvyqtjSc/vpzSc2o674cnNon4p4BMmTOA/+NUzas5/rOYJLA
dll9sKgdexVRxgB/wETN5LxS/Qe/9XsuhWcgSk4FIOui6WCXF+pmTApRvied+K8u
mxld3wX6da+aYYkvBcV5jfM44zStHOvEMuVyMVJDuW3QoSv/5ph6cDunzo4NQE9b
3qxkcP+EoXoM+sFgfr3gswsltf/rpiyclYfL+hkXqIFWrf7YKli1i4PjDzEYYHvY
tkrDoviX74RgEUY7xTKjqESzmYqjndUZa+XCJBDcheX7H5cMxESITSIpkh9JYU+E
sQfbRovh93oPqS0S7bhsG1gDH9r/VzUfvaR+6nXXWR0YTv3Gl8AmTUy6FcjurguA
zHzzTW21OxBr5IkEJ/3g+RFnJNczIzLGAprFx9vNtpKTyDnHfFtZqyjhOEq99BcD
joDTHOJjIrIja1/NsBUoIpAsKw53CGWv7zXs2INcwn1GDXD0EFgl0qW2w2EbSK7K
6NqXSKjlIZFkIfE64zIvVQRRm98WiNIJzycWfPq1falb6UJY3lUl5/++wJYSYvH5
jfpIMhf1LueRz7Tx+YdRro0A9LywCBqS+xkWweherSsRnodrf5awZQ0bmC4wacqE
86db4s6tEIxDcKgWHopNXujMn54st0X5I2PzAf8ak2l4/USUIZgEUa5BZma4pCrj
rFZ0qNxNOxZbzlKPZRYaJnfmNsjXNUN7DNhgpBSLcpoa++IQqNx1HvEsoh/Dcftf
hWq7hf8aemYuECDEGPeDYPfkDP+IM45VQFmZrZOqKnu6v0Oy3TdGkNbKVXD1Pfa1
N7zv1n2P2X+samepKJ1mkHd9L+6jqa6nmYR3mSnMx48PAH2vk4UcmgBUxUsKzdZf
ICEjzYyp2U59vyEVo1I0hzGqr9LDgnb6Dnrv2V6hncedd2gzsKwItSlV6QLlxiUA
xhQMwY5Fa6h1beTxnTZcTBBh2/u5fArD1KJmryBlHuQiRx9RlFnbGag6Bh+yfHYi
VgDGV/uRd52c7+vEGEV+89nSVdRaUFC3MxwcuI2pV2sivjQ4Kix47NR9/YEw/nSL
ZRikMVifToF3ayFe5bhcX4wVHMeRSAnbchlWATEnbRRy81SLS0azr9wZG/apcsAJ
9dicLsyxD9xzcPPhUMDZwm64BaxqGP8MvCiG7O1uNOd2KoqaEqkozNIV1s0xaZ5u
hDyd5bToRPhkDEuFT3paBAUuNe9cUzoQ6jphKEq2QctA1G0feMXVd2kseQH/8hv8
mdh+/kr2SSxU4OOM8QLFQn6r1ZRC7wZaD+zjIiKpeLHHKgwI632Bbgoo65H1OKJp
C3Kp2GZ+fv3r8/T87i6rFSNQhLDmioy4lvVUHk3eIcvRp3mc/BtVXRomYfXa0LUd
yfs568eC91S4hF/8YV+63XfnOxAqNB1/z4AFo1vH1YGEsblnnYJmBBWlmsi0tA6/
9q5OHGSy1hxjdM93aLJReFJROCvrKNMYLNlM+20An/4Ek/OSfebNWCBj/gBRf6e2
BnYT8TGPX1uxQK+i2HNAWXeBW+bgOZArY5hRE+YWWFzd5OJbs/1EAA+VAYr6Plb4
v1DeABrkl9X/KvtMNhv2HI9RYzkDJp1jO//+Kpjp97hDFiBLJFkh5/9cUCWBM9F2
Tlur68zuPayqMWbeZYGCt1iIsxmNpxamDVjDiYZQMvtznj9V7ekIBEK2B9eo4dIO
+fdHd4ED60DSRByNqj769+vxMI2Wp72iLKXkLH7m/rQJhQv++N8Mhp50urPkDic9
O91WtGst7b8nGIksgeYdBbD59S1k0VPXbpMPPFPW7rv2wuxojk4Mj+P2jbAk1VfV
iwilSR6yIsWTGk/BI3LTZ5QxoIn7EedRChfxtjXQF20DcUEogsJ0w+Y306IM33H7
cQim/LCqHbckg5HdoecGCBeDGoKx9+jnYYCfZ6M8zKp+czEVhK6S2d1o0g2JpccY
9NPJQZu4WhthJ7L48whWioTsDGpCWjPlfVmKKU9Hsl9khrfau6rqvvvRfl9w/3f0
jnYLTUiBfFaqcdkVGRQGn8+CDGLT92IHIbnLg6V36UL6dpVwV36Uk2achTHoLrl4
0IVWVw6JMUu5rXQBSZbzsAIAHc3177NpESXpc+BRm9m915uj9RVfm+n2qVaKnUI0
3kq3O9vMRj4hd/ceXqIM0KARuh352mCTGWSQOuhZQBUu0NELQ6qazTTzGtYEC3/M
ynEryjJlw7qUNxWFeA7USK3zlDWzSD2cUi9ZUAYU50etMCqdm9B9HgD3t43OhNSc
IYApXUy10IEmURZoSLrLWPPUipEy/Fc40IIHw5HVfFFiigfWxi6rKDKfGz4J6d6L
R5roQFRHExHRM1BBHteMzvA62QPh0DgZ+dRuPojP8reWsk7LBg4bJ77Rx5I/4yOG
+LRWilmjbdbFgHAhwH6oCImNQTNeQ8jhL6GvRCotREetfzmvyhFBt1+UNdTEUCJr
IkRWXLwZpeyvKb1n0SQByALxi5ekf7qwukA1y7CBwOMAZOAaJhY4Db9RoBJuxMla
I1TTV7Hmozsm17k6Q8BIqq5FQZAgN3EN1lNaTZYKo8Ro0X+eBs3mhmo99GZirv4h
wxUhgg1ObDEfHV30Gp2JhADTN4+X1cPmHLmNJvXX0hDZisNTV3nHO3L7gm/qtwMN
0ap2F1PdM9fZSB+phiebijVbbS8mONKw5pwBiJj5WNz5VDsEwCiE8Z+4TWSQnfYf
N/ypgJLqtM7LQj1VjkjXhNKFDj76Y6fMXjhbXY3KFD3Kmaac2OmjXUTYZ53fnD11
efhauvimfUKeizoteHIemzZQLXPVwPtz5pMgGpFPptNSTrZM4YyM7Zod2u+C7IFZ
NsgH6fWOTt1CwzScYPy7L/YCm+LYDZY5TxuSgKEScbgbxxCNCzT7bv3kFy9Z0A3K
5EtoGs9HxoMRRoM1zHZgmb+nbl+awSlmsEXU+d8heRHumlN621ABnW0hPBAIhTvm
PXu28nbNWLCym2Fai89EeIZgeVfxUg9JH1TgkIPxEfm32Kv5hUS7/N11WKZtBoKA
zWOydOmLG8uXt5xmzIw9SDf4REVA5B4C8nZmYJWXKaaY50qYSbvZcjXf2NfiKa+D
FkSIJtHnwYdVZkSNhqc8ACGdtKo4iBs07OOLP8jAVePKoQWaaVB8we7ferpjp1C5
FJ2OQnemeVbHcx/np5dOkkEf82iKBmy0DnKYh02VgDP9VJoehBji10rMNWQDuky+
JXL8Lsb+CIQBghFomy2Vm0iuPTXicyQA5qnPhS83QZYiMAdvpDfONlUUBZiXWIQK
eabF5Eahjy4hrHED0uRqdp7yPVHqBHz48vzuaouckNj5n/O2G0ptzd7ATMURT6cg
OnDoFjRwqVVqzLefGuwKXMvwUOeJ9X6dOMUB2ZB8/fLFebbVK02odiZJLg4tAv5b
dXjBCdYPO8Xx/Sg/lR+XDgazbYL+IwSWp5AYtiKWSMqtZEDOCuJOox88g7J1l1p4
HZhn0lePTjem9G85YWhRdewIqXjU5L9iOYqiH9Ix5lBWFtu6A5P9100XvdVDpsI3
Sw78Or6N54UgThq8pcnQbuCcwqGGxDeXGhX++q3ltq1Q4HmFBKcaPxkCu6qCqFGy
ETWqy9TcVcHlWuykhqHOKqBGkoy7oLmLSv2IfbRrQWGiT6MMWmaqfAPH5bBYhkqV
A2zCiPqrkrgTRLD/eq4ppLUF4c2J2/E+FPAUTXHzTI8yySnIU3ZT/ICjhoJj69Na
xEUjTaz5e3L7N5pnvIeGsLP/enTgwuaC6mqKvjJ54anA0mN/+8bq5geBjMQPAwA+
6j+D0DR9L9lJvedPIzMWm8bhq65Renl4vCidfHUJ49n3Klo5R1lE5wdHerHJSwb+
9WO+JvPV6WZb/GOkiUpcEG4Vkmb+cec1QDcww1L5Bz/tJiK79+3Plj3LOrs/WVTo
TaFE7EYQkf+/gAHmbt9PAzqEZ3CRBk69sPXRV8nG+EOR7/Di9wIWBynacrVqeK4L
vNqiiqZn7O8S6f6xlGtxJ2w4j4RBBmuKzmCFMHvfTg1PxYuuOeBj36nGSJ3LL4F+
9doLGQIfGqpSDfX6g26/7U+GoUrrlsV/FIco1Avd0Xz2SVPB8LKUoEWrBRldsCkq
Hce/IitKLBLtA4tG9g6XJqs9kqhrCNS9+2WqapFcmZnCzMINjSNWCHCkVM22+V7+
T2YPDcO8sfm6CSma6YEDRmzFy36U8rmgFEaWXadhlV4/35QYnghrqu3+MgWfEa24
v3dLAO5gwaRnX3lY7LR4vYXtQKrZXvSDi5ooVrUQNJzvhCtrvbYT+Y5xi5Ck5Rly
Nfz878Agro7c80VfAIRy9f7JD+Ttk8dQMo+UKPABWOnu2W05YA0CEHWyz3Qe5bWJ
EMqeCltgal+qZ6l/Xb+SBvcI2fsgZpTN/jDA6PcR2y/7Q1zk6kq9GNfuEEWYe1+X
VwYRakd/6gxOulNf5ZmfS/F8FKDT0HZ9ydmuLMKpf2byHR7jrz4O6f9AoL8Z+SIc
laab4vR9JjUMJWbRCrTAZML0tPeGaSVxieXaftIOybkVAhuqtKZHktFKNESu+Kc2
f5NkeGtYq2C9KjD667eipsqH6RTubZ6/RMNryPykOEf03oEtt0PGUndskW2ePDQw
W8UuNR5IU08cFyjipTSYmbW9f9/lgr0Ckxc5R9xnW+Tp6nOArgfjLzpjDPJJHAI3
oQ/cinrZxwzaqmQ7KizPsXZuVF8PnxfrEOaJBJcwkB83KdM1pytBDpWxvAi9fVrC
i8ZmNiAO2rcOGIQih3aNCQ5Cyr/mVooD6cESwdefXi09joI/QJFW9nvmSJMbeqD8
xTASlz/FuU28v7IxEmn8na8/0SK4p1HiioBe7B5vBU1V6daI/dO2hlObK4OpkaF2
+G/jnDGPAynVfkLjYXazgGyf/RGp+wZDzjb1IuTR+2pi+778gfooYHFJNRHt81Q9
RSVIcPuGD+fsLmJOz3Gg7dBrGS1EYQFC5fNaQQU8zGr0zlJF3N9+lpQGujGRDKvZ
2PjWYYfu7IJi1/1n/d60BFen2ooc56aavxEU9PXIDJ6BeSD/Nvvk8oEy4wCu/EMe
BfJ82dUAhz+5lmF5xewv32Il2StiRoEGy5WAQjhFtoEf7qtc8g6qjOKJvGwPMdLy
SQW05ceLKLZRQWA2qUE7yuVazJ00ENaqxmY/xfe2tcGs+wvkP5jaYOtC97/nA+mr
Epq14LK2Yv/+f/GdDjYu5j2EygyoyHlP8AC3CXaOXWi4wnRJU1z8op4bsBtkDs1Y
eqChsbH5xXwdep+rtdbza8Dox0C1BGr5kcTgMlDgGQuiAlfl22psGlZo2XIZqrqm
MqUR4+p/Fchi28IeMvb4lwejkn+LmiOl/wg4KNBjGB0LdZuNMnt9NWHsmBAywOm1
fxr23w/T/wm7mX9irpw5LyNGiTMFwAKvLj4Qqb4NasDcG5VayaRG1k29mmcgcXlK
dgB5UJpsUr7KMwPYRXg3aRICIq7UXA1o5Q78zO/YssZnx1Kqdkh2AT+gR0e+Ey+4
WHNpIIuG/DCPN4HcPi8OJW1oO/8d2DHBihufMgMwxnw9K/wp627m8cYSoaVWRWLQ
7DSGOjSot/zPrJIvffknIvzq5daKbbGAhxTISkIWa913Qm8cXef+NW6uZxGwDuEp
xyw2KcagosdQzo5fdd5aHWk0Mpu69iOI4/KepgYk7cKt/dEn89yXRoSJM34UV2l3
79nBkMV3k2HWxGD04VvVX9jMuJy80CnykLepRP+Ati0tUHlibpdnm4oa+4CbW1Vy
kHwdd9+BLAPSJx8W56DC58ETVQT90KDbYMOuwpmP+h7wqvUmg7cyrdqvhON0kKub
kEpJCugWUy2WeN0xQ6LrfD5H7+La7NgTIcqDNP+nEpoPup0VHuNtBKnlbkc1+5PL
/1jSuGD35ISCImlTP9e0qCem8ZcmYL8YLtPowdjHmHJScb1hxVFQuG0EH92jeahD
1idEkA1R4PZhP3jy08qUL8L+XkqA2LHksoEuYmMCNhVirKobpK2LYW7/7HZcwhE8
f8N/Xsf3KUu/Ii7NZUqEx0kn8Rj5BVc4zOeMipjt/JN5AC7Iv6lx6HDlVVFID8As
tulgMF1QtjYtdQMTD52sYuCSuH2DcCZK/1lougtUOKILFGptWGJbup1aK4rwoUlo
PdLoZ5vh9tltkPUzGvnOlZTVe55GkPuahGL2WzHA1CK/TPwlIxyUL8txitzwOnxW
SrIeLqLDUUedv1iVqI40bHxPs4RKBEmKtavvewkGea61OmYeZbgqOH5T0ookgl3j
UccK9dXkiKUOttG+T7lKJ8SbBjErydnZKjjS+M/R/UuKUlZg3sxBQq7DjC4fH74r
ek/qK14Q0eANTUHJ7J8GrBqwNNurwVV7eQwVQ1lTY2UxgZRpY3mZyz5ptzuTJFYp
BWZh+ZDHO2GMJnQlVGhYPtXQGdraQ984XyV+mgv1TPqlk6Gv/Jr+I5KQ4/Y3FmcS
Z503kFtseNOJ5hIKIk45FQu+sS4UFWT+KjkIVHHjj4BAIfmfM7W60Dn//xBreM0a
HkZUTVe+7KeTE/TtxVcOvL7CNEbi0V2PC8yEYkcPu4DJ1ETGnKDQKsE2OxaPzRT5
HYH6fWQTP41nFwR6wJAkL3rTveQvHPKvUg9BK/mD952PE3M/Z8Ml7RboacKqMnTa
grg+6zlKvh342DEtr2/wN8iAJuolmraOAwwFf6xFprLCNZLCO+FKh5VQQ5VCUkcm
Spj2dbnX7/yz1i2DSPh9m9/Fe0vuUYbdB8KNDvgMW7MY6Aub1mWYkMpIKCyEJAg2
VstmUaufNrBzV5GV7hWCLYMPdfyNL14zAHjbI7JFnemdymjRCbUdUi+/G1P4pcbO
dQCXZq/E5aAmKFJNwmBr61Al6EGRd6Yxj6t1pS3ecDvBjt4U67EpUAfO0Tu+P9rN
Rh4Dinho9R7DEieuFpfOgGtyJ7Skmtk3MZsdn4UBDp5ke00KPe51RkSULqKdZ2nu
emLIXB1QYOg7zGzVUN94AeqAam4MICZScWsgbbxqlI3/K3HtUBfXWGp+fKEQVBOQ
D0HJb12AZk8MkuIdMa9xw9zW8Chtd5eWL0Dv/NGyFtChuQsHTYwfMN7368nEBMpv
/fdDHQag7JSJkESi6s41anJ+VGW5L/0FPRwCiBn2bnv1XKXLMP9wrooDA4OdQIA6
FVyrYhzIaorJGGSgw2ZPr5KqsVXzltTA62hnYkOF69Dw/iJitasAgQ4rgB0VnAYz
4HvU/AKDbl8t8meBz5GNC5qodWV9V5Tzsadlab7KoxfCM8HfQewDvtfaek+HOzSB
qYFMW51zpeBxTQoZiyWXXjTVNDdYPGVU2BYLS4Z7YlSO2pFb9nhg4nOFSz6abjKh
VaKeoWIl6ndAiFVkqHmT12iDeM9OesalCP7QRn5Mdplqv0mFOgmC1YZUhZMaWjVB
kfA054xnRTBL/Eygef+6knV9MMBZPFCGwJuoUkQbTZWX91v0QGf9BXsJXA5B32TP
BItyfs2rG8XX+I8lOjwB9qbA0/K1SFO3CjHxPB4xSgDVFHhLMgvgmeHWzXF0xhk5
A8Rg6opaPB6OlYKLNN7oJxtZXd0nC6h8toS5bTeRHq9bNEhUNlOsndjEnVzGRSvv
A7TphEiNc+iwRDqsyPkn8GyxY2KdvZYTU7ScIRQnNH+Gf+jywBcFuh5XSWllWCDH
vVfPRJ5j2aNQsjnhY94d3LnGxLdLtNLGnz9aYJ4ETVf4qJ7eRK6MjF/nYnjJ/U36
8nbB2aosiDA8weswsLpognLaphHWL5+ywuGDgRPjZV+AcVcZfZdezNQzjJHYL3BF
z63RnCb3m83o/K3uMmcKZ+pBF4+pCMSoC4FgsgDIx2nRIhErRu0bXhjpYtOBNJ9r
FcwhI9Ig1Qo01lVhLyeiEJ8jICxg6bYDJYOhvn79UYrCHg9W01jVN5LkqwLSs8Hx
7G32oAk0EssaLqmHSDtWdFOpRzbhhLna/jhSXROt8ajk2+ki/ViWAOKKMFfn2ZNJ
T6TyY+DTtLA4Pg/4JZ2LehGNUdis/Hwa3b6uF9ZWHxr7csl+iqWahfGZ6siec/to
tnQtgkQOdYbOC6VOabz876DxZSNkJ+otgpELHrJOYEoto+OEn7ossX5USaDdcr5T
bq29BpOHrtDbIOPE9iGe4F/+arWy8K91KXmTQGHBIGT2C4tvA4e5fWfk4ib45Kta
ebbYP35hJFOBRxZyQJXwiroxanaUk5NYkQzaQVFJmdOyx+1PIcFnbHEVMX09WxdT
yp/g/7XWJv+rcuXTdfPxoFefSzdYTqarervfFBu4LvjnpT09XcpTtxb3HJ9Zdspc
t0RWtb007M78atWPUEOrKVDf1rDvmEubC1UUrFedRAHl+Wb4psrd8IbM388c37ff
NOuNMgeikp9APWCDG25QWvDxbhtejMp2WK8CoWLk/jKLi1Dh+loHM0Fxav+wE1ug
pfdCDXkTMkXb/gsQ3f1uUoaDTM34npujVsbblKFXy+EOYWdPL8h7jOYCUK3UczM3
ShkYi4UP8a4J+IR8aer10kW7QyCt+c1YSDIOKucSJQp/6g59dw58IlpUCvqL+7qb
5qUVHPC0t6UHLjYDiE3Yi+RdJPXL9ZuUs9hLovIIx9edkkX578zR5kQdn0Ia4Jgr
da1gX7wwEIm+rtXey/8Aje+m23mA4JGZdfC4VQnZQ75QxkWpV2GdtGNzrAqOJAmX
hNphgEn7CVJgMP8InjvjjigJO+r25am0Lva20it/HMUauwXhH7wyoY3REW/JcMEG
MvJvv6ZZVv4lwwbwqPxohv260EHc/m9s0oJGl6bmj42+hJKkUHZHwEiFbKayzZ3M
YehNBPhsp7fSONQmTMsogxAvDYXEj1k8NLUscSW7FIdVZuXMekXanisqWkZARg7g
Tr7/5D9Sd0Euzp2/C1o1IrFX3NZOQYLWi/Hwcd+7Lc8R5aEP2Hb4r0U68sytAmaq
ML3BfMX1H7Q44edUq+t5jvh3rYvygirhmKS0gULfgUaO5wrlLxoQ/2OITiDF8Q/k
O6uqJJ2Ci9LC9+rf0BhFO+zb43J1G/JhGCbC1irfh6ChBlyqOpDnHq+bGtAKma4x
My1GFRJ18M5TBm3ml2YDhpBRKFg3rma/D1234lqvZL91nzYccG3/lZ2DSG2a/Wev
Q8PyHc/XkVK8gecKeTgJttmpYJPuY73NLDvfjJ+2PZ+mZ6cuI9XaFgNxD0RG8QOr
QRHrMOM43nOsxJld4bLc/8LB758IoqvEolZJaqYuvUBiyYZnQfZgnEuJyn/J78ey
PLix/jdU7hK7dHs0VIujWFIIYfpmHnm0Rx+FdX9N+MF8cGYxdU+FqTxR4R8/kL/t
Q4CZR0qNFXy6uYmqfDYn5seQWETDjX8RcnyQjtSbhceMttEbaK1ZdVZZMAeD4mP3
zIr0Mj1oOAw5mTnw0bKoWyCNCO1Jwo2QcXzrVbkmmjFgjv8/4IZ+ZMQCbQdTCqUY
b6VUPm2U4ehXgUIuFsfhtb8oWute9ndiXqOMbesZdfRP5MEfjdycwUsALlRoqn75
u86cMnQtvjio+C2L8QcflkxeKHMzxkdrrEvwgR3LUCXdU3aQ+w//tCXPwrhI+TjF
MOYNtktAPH8RCO7kULkRYitcMEVv125oF99IvCn2Cq28/BVmRv/kwHZw047HEAfv
/rDlUe+B1i7txTBdPQRSJUaKpK5AukGy+QQKBO/PFL/PU6muFeGoUdzNWwfXnfp2
Yc6Ru9OFcL3QkIOIXVR/DdvepRtc+3Zh6GkLeFqbBazMEEB/iz1UW1BTVPjmIDNN
YlYuIJ4ytQABa60dTwSzHmBkESV4iP9eg9hEZ+baQJLRT3PuDZvoHrzPoqEmEWUn
e489U/3se957oDGJk1wmzCAWrQJV0Ih4ss+1TgwNGpXcgyiqLSGEC7qkXhou7q5g
+9s4EABhRtHjNCojYV3CgqN06/YAVtN8dJl8e2NwYS7DRlSdgCjShPp1HkyrxjZM
ccCjX2qst5EZcKGqn2RWVn31p1tpGZzNAhWMVMqq/AGVu2JuUK97BdUh0ohBR93f
T1GDbMXzOLhpWG6rXUlCY06iav8vktISroEEettSyQCJSkxPgIylL5vYsUfaICLx
RPR7+ZWRWOVdzY3Z1qhoM8wXsEV/YyzojDFo2E9k+Bzemco3MCXQq9vOqrC63/K4
0Xx7lphU05ayiIJHd6ntZO0jR8wj90lXSt1BEI3qW3KMT7PDOGst22+K97e0r4XG
GLogOpIEfv+XcRJL67smotMntfGuY/mr4BzAu/FWQi9UZnvnKFzdNTQM4fcBZz+H
MuuuiFhwkHeCx7yx8bQbPRWg+JnYN+SGA9AT12MK8kYi2mL3Skyd/LTk2iLRZiFK
RR3nh6SvRXJjy4cGq8b3kK/Oti/Gk6bhM1ZqqHvrEtXuopeO0G4kLvk5uOYUf1y4
S5qtP6VuDwTKO9mdYHLTOwAyqVv0pH0bEXRnFzvyj1+XfN1wz+yIARIZ+c7IhGqt
QzKSEDI0mJq2nuyAWzTQ0mokzK+UtGIX1DJzCavtHvx4nrwBT63vdPZmEqHy9eJd
sC8rF+FoxX31VZ2qnTXRD834f2aJ/OR1bjL8rjYudwTGDW7jB867GORRTtpIXVmL
bPM32CFfqfSBMMVfgFtMfXtIUpMFzw7eKUE6a2gvlTzrxFeBmT4z7pCaKHmXZ2Vn
+u78uih0ew6LoLVcbxq0jzarPkExnYhyrCElYRMAc5ZKLNiK1fbkDrqWuHV2wkm3
YtKD6uNv7QIDmkkdvEnwnM5jyikjDCYW38ukpwby14FEOBBLR6lpayWu1HqqjE1O
GQ9fUy3yzkwdc/aGDaDSzznXwN3HE7PzhUEFwiAV7bz5DJWINoma+qJGk9M+N4qE
B19SkeF6sghbLZSt2evK8BCFCMHP672r0GZMpi5B2HUeMnF/ttcT7Dopi8RBEala
BCXLAuhdafvAHWEps9VclKtYHvUfLlnc0vT5vOprlThMd5lLI1mF+p0bnjrptDbD
dE58JuyMgePRBxoG9tkQy0H54IjMm0VvtHbYLv7xL/BFKiChI3YjTSajA4+w0BYl
Rbh9Km5/VdtIWKlyAv9vtX+k/65mCtamW+XPgP4qz8ejvGAPMkKHG1Z7Mk0Gv2Xe
cvnNj5v6irZVGhDLBj3TTPs5yFFi8ykJ3ZH/pC7jV3krIq4vl8F6dS9VILFyXMBR
/D4OAnoNI9JagZD/6x0fSg7ce0cvB75vlM+lS3XA53db2Rs8pFt6TKkQqI+Pztbr
/8AWSOLx6p1eqdbzmT2rywHsbbaSXC3V1v+LVPI9X3olaBX3M7KYPslApDA6EaGH
xFc7ZstRLeg3AvatB5+Ou5b2MnN01dK2Q7woXaj5FvqSl9WLZyqBx0wGAMlwsn65
2+TATAhJf58dRHMIwSzEKMB9+4eLT+LuUzGRz87BIwSgcGiltqhELFXzQcnia4hi
OsBuUPFNqnqvZLqrBd6dGiyhgXZxnjKX0/Pj/5Pjz9NZxmyrYcFe0reome1VR8aO
eRbUoXXE6b44Ht8Gwv9KNX5MSs3PrIUblUhUODHejK6A0pnFfg8mj3B2NZ9bOwDa
nP2B39uBj0ARNnzmwViuxDhFaSGqfFgb3ZTpohlUb1RfGyiKJR3jBowH1pvn6yI7
HCUqGSBbHp400YW1hXN2VlFvBsYmd7Nr7UhEiJdsXYVDunikqUxVKluryDPeJT8I
eUAuDzyjH2xstutysigobDZwVe4eq1vRJzhP7P0E8y6mzpLZPk6nrl0X67ATzX8b
hhmUB0joqtW3ZFMIpQcpp7N5Rs58T4iV0M4IMmSxj/lPyZyhjiNYCIPbZSVM/U0h
751GvvK80uOFimGY3bjC0OQEEC4NQDFXGumekSnNwp40j+oz7omtTbxDxqhw05zm
fJcBSGZynS8KaPpfUjYJJRhdh2us+t5lfxpoWoVP160T51GEw9pKIBFoOBgeDB5G
N9iMI0JvIGE0v8njH2uSfU5Uzc/EJsiwMqUf94zzZlrGFPnlcmUDjGD8M81Xq+ja
XpOvDCJRu85ZiM3jFM/kCquWn8f/fVCmGTLf0BtXGv7JEBQJr0Fj2q12DIjiwzxT
GCIE099JuKK82rqP7twi3DJxWpwKHc3ldkhFXoJSmcKU6zsXr9FisrWaHvNyQcIb
Fuy7Xrnqq0cRK47ZT2iAApcR87xDatCH35gUTn+u/2iIVace71Lp0VgctS9c3Tv3
9twtwWUTiZo+9YRQbceYJDPCoTXkGF6f7lMuNJgVR5Eehe8RPAA7Y2tQjKYdZRw7
dGu+RS1BuIKyTuKsUQcakJeZqPZI6cP8gOy+h+anLlGQZglz6Etf15msgXf2A0qm
+2bzj5qwJTTH9iVY/dRTcKjhG540Vz1Jz3AbrI99nEXtpRlANOaMc3HZtwhT+cuN
/QmYgf/QhzynXxtLMw0BBy7xUEW3kcCBKm6FPPvqb7BlvqUOqz7zuf22Ikr6acEJ
SkxJdNMO8OGR4Ns4cXIL9bTCbS7dWq5Okso+2VoW7roSVTxC7VIE3wRaO/352feK
BAqTgPtYUQ+R2Wse+4DzM5xPSrBl0Il6TxARZ6nv/yeqTBqfQWwvzga75kU3rRv6
0lID4E8H5cug91R8pAzQaAGFvFTDhLtqw5IQBTLV14msJr5h+7AT82E2W8sSB1am
Sk4++0Q1gE1XAmVnqzlhcOdqb1LOePZ/fBCvH8PAC8QTjxoit/lBgyAC5BXU2Vqu
wPYZ5lawBrYpXEUtEmLY7baNao5NFR5D717uISMNvEo+Mf2qDlLl0A4rKSMYn5zh
glFtevv2tpxd4Zh13kv4NH7dCxfBn0IxmloP/FqkXnqT2IbBToBwiaEV9Xqk/Vlu
kVU2KyZOg12IPmXLE0OMh87+nPXWdMBlch1+iU8igIpAeRv5z9Q3FQaIhkXlhQX9
ZCZepmGaZCAMsFJ2t4kqlrvqTKXVYSvQBM4j3Cm2FBXI92h3p7OUlyicNLJwV0oz
iJLVBn0kfyPJ8POMw9648JfDY+2mz0Gil6e3pz9f5rdsR15tFNgwcVj+7dWpLz0A
JktcHCWUPCW9HZgOzbLvH/veOtvZtmcAvZ9ilFOFQeonTCJdSik0Yg8//0UX9oGN
1i6W7SuJg3a94EC7TbT1prLIRogJB0LgNvA3rh81zB0znJZ+enaog48+KVPYpfx/
SVYlYtco5Pt3PDr/m+w6N6OXFdoxHgrrJjy4cYyBd7zh5IjOlu+oB4jKts/RyI5Q
Otozhs5HzBt5NtECz59/ft9JlHrYUwLU7u6QZ6u5ALSq/AL7InOuRNb2M0OP+BMP
zbTSmiEeGPa/EjjQu8JOGBkQ/3gFDEHhtTLDUf7cFMVoCJh+BdH54SmRebEHwIfO
BZQ9ak1futiDBpCO+OkUNDoVx91G1vDoiJsSFvhA1t2VvIQdjlTRyIW4uOTq8kJr
78hWRaRWNAQM8rYY1QTnMXxsT/gLNnFVkJ9vDPG2dBJVj7BoYSbueAeDlqvsOhDa
OCvEpwbouOz0P0CLfH53c9wbvTXPsT0GYoghVd2Lvul2yau2yOi6cajqzR43VKcf
aScwImCDsiS80S8PPCF0jr0G2xMdo8YSryoGroG13ij9pi65+qjezDex+chPaILs
hhGGhm+fxNkV9yauuTZHluZYvU1rrpUHHNDqofgcVp/HhMwyvjEVfFt71t+T+evE
tmo2ivNbbm1QiSNP7daW3xOm9qOe33YB6bWFVAnKtAZmJgpATvgMzX7FBePWtTu7
xU53g6ZPnfLeSiuJuD2vV2hVheA2wqtcr3+oTxzt+fCgzuUCTPr+MNs7odmOpNB9
VpCRLdDgd2BY5rDPQI5ZmSd0xAvNQO1rewblcF7+Rvc+Zyf8jXy+2ccm38FNnhr4
MhInBoNXoqvBRaTFBqhrvcXuv+KE0FaSDFMU+Te1X1DlhyVfYmIib+LKJsKzi0LW
xc3au9dvqc9kmRTbDcNVKRlme+6T2lfiLHnn8pMw62+lfO6w8fDCd5hX24PzrGc+
BQIfNa0J5UPT65g7zTr55N7ir4j90nZjewbHPi7bO9pYTxe9C5D7A/PfKlF5DiUs
HpDgTPA1MeVNZcZwJzm4LrSvQSxFI24UUxP4U3C0cgWXHldhLjPWe2bpzS/e1KSn
6jgJOBhcb3yiGErV5hRMUPulIYGucMU5P5bb6n86gsY3PNF+1beAPusLSL6AlFC5
P9oxjFuB4RjzV4SbY2siF1H9MY5tK6pcAdi2Pqo7QXKIxxlhwGy4IM8vqhNNj6ra
ZASk9opzaPYwfHhXJvmUKrPijgEwYK48MCMKnD30lEkMY7inoJ0YNRNFltnUebTq
K+NntFFFxGO48q1q1KLtzeEUNOdTN10xItLce+PPZYOonE9e1Nn1ulMt9FJnmwRa
RN9gsVXZrmxnFp591pMHWVp7M6sL82K7wzqTRkZDPoqa6DJZHH3eusBzDYll0uQs
DrJteeG5SpnD6dpI8UbsPASf2JGB+AdgMCPsd4iFo7roD48LpMMEsySp04m70Uao
lage3Amw9ZMjv1GB2a0yoqfGPfYvAX9ImRbILc0KMfXre2JZCZ7R0owGT+0Z5owS
EyapVrMn+JEZtudS6VrY+0EqAXsaeuRgffo9sVmQjtt7rNpLp2zNC49Z9pNE3GGD
dGHMwJooU2XRK5DPiy+XzUadKdtvykM+f9pzej+IKfYsMe1r9Bv/zAnggEEK1MDX
hCUzwjkK90j5IO6ow7PpvzqfhOWgROw7xXgCD1jK39hY18Ip/1R19hmjwj5N0OUF
QHO++82D52PThVbxklRA91YqslqyE+/CSE8+MC3LnUrm5zxOwuk+Dg4kpTG3SCuN
OwlxAAdbepepsSr2v9tE52WBnjZMV5ziR2g3AKggOOXZij46gpvdDKVV3EstDVHy
OlSPHMnYkXn3cUgfXgUUQG7/ZaRgjGAH2jDco77klh2MJdvMx1/xNnGUdFvLBs7J
MNirm8qicLTt+XQqOy5qL68R76X9OdRQFHINcN4tmRiOe7wVjAio6LK4BMl84OSA
zKzADNOSvhGG3mYRxtMQMrFYSNHXCsiDMrUOchY5hiua7s3iBC79HWyZe3B/DewJ
Uuo7XR0jaR5vsA0Tq7YFmmt6SByTD4et3UffX73uoInqLLRbcEnZ3r4vrN+MasOd
/W2BPuGBMOgiDPVuW0oKA3SN9lGH87o2LszN9Led8YAWirMtc1LjYYO5pTvzJFqI
XhVtyBHb+8o4BndbRb516UkavEKxbtmSu3MW6kD+/N54d75EGNrfXmsy6+3iDJLg
bfW2JCCIHa9JOjzd3PQU2x9VM94oY98DYlcS1jt3smJ4A0KDs1coRACqnzS0YnRl
chZWYTcipGdOFsVhQZRlhl39q71nzu1S+xOakzeFtaDugUMamW2WNP/UOzohKuAv
UOAXKyKuX2bU2/p+ERceqc/BllVbbjvzwl3gl7y1Dj65OQrlVsz+E5fsWv6+/ZtV
mJdz5W3r0u+XX6ECoHvHFVfe40yfAuk4okT0hiiDje5HccQg5NmKTvv5M/Ppatmx
l8ON+Xj/q7ruAuWawHC9YzxpRH5+UYZ0MOmPwwCS24a5z6mFLoR+3kzM1MpINV1n
YkEGVoaS0M3LrNWzhHLt7YeYXsbR+WXZdcXvvxPXQt9JV5HuWMFCNZ6BT5cm9A6F
rtMG4jhLZSmIDNztESCS1QOaVokUZyLtEDSi+4XvrlXdXnyUviEe0ddqZKFB7tkg
0XbveHA0dky1MHTuVytFPauR4JSg/9SKlrNbU73+NIm3Zis+WldPMzjQA/+8HFyG
dOGVk/tkraqDd6gnzJXwVJYULTCcgDIOJ2MgGl4HJxNu93j3OEWZyYlbdCaw4RWn
YwxKJS3tIMwsCWp/YnDSne58zF9QiV2JCB5No4NNBCTH5IjS4UCGXnrL89EKxrX/
bJYM4Njw+/xmd9esd8h++PpCtP9XGTN0pQH8NO/GVN/tYUwDiNAefp0q36gZv+4P
LGeAjVepwgpbD+zmiKnUos924Op9naCB9a8HWErRsvhANuZhb9cEaSxWfDfqXa9f
OvdJgKoCibRV6FLT/CjIOQkzzjlDf0n71spBk2VQHPYipSjewTVlmn+WyKHKIV3R
W4QEzYPB3NmLiIbDfs7czzECKpC/FVfJlE5009tcPTlLzvVsskImtNKR0P+x63sq
U9r/LOXWGCLXgpj3zIQpZXuHWlMaQMHDdggFowqkKK9zfqMwvuMkIi2kuxw2POWf
7LlOhZAS2EabgJ4qbMBCQWfTKqOH/6nJkL+SnZPjkqUahBFyd9XsXA9wn5sFaPPj
xjKoWl95jYD+H3vzRnoh1sMnmnLM7Mu8PX1UYWs/i5/vWHZXiLbGhKjzzXwYAJaQ
i+1UcFnoP9qgLF44l4lBYE/OBB5CnSrvq45nX+oyTlFDKEphNUvjJS2QoHSrLBNY
Ef/wcyp2PJxs/IomLiGYktbX2FVMzOft0tZrfMzAkdckG2pf5JE+c8SYT+XvLpUY
dUmguAfq5waGHMA4US/cuPyWmZ4duy2LYY0C9+wwgjcjOP/06l+vL5iEStyHCvLD
ZwVUr2snn/x3U+r678c0UvwmokJWYMaz3cKausoxmn2yI+pOXL0SwIt/kApdc294
rvyB3WOdLEH7GP1fkzP4Jx6CXLsGIcFlP3iB2+BxdeU7+FhKLqxQwWyaw/Fk1nm6
FxHGIVlQI6pYfDmdJ8Jcdy1ovlTt/Hx/+OWsjr5TiGYwgAdtiBFn9H9jzLBxGPxp
kntjmvpTjx3ORBkmdFGd5x156Vatu2zIBTomdVRuf56cxIx/W9w6JQaiYxkO4vyn
FpmoUIZNa0NIIvTR7duZ5DtCGO54XkUwHjdN7vn+NlFfvk0zav8JbtnePzaiNJC+
LJ9HMbxiwwNFy2rrIsPmsZmYdDgpTkk0eyHa4XodTWWcGxzAozrlP+DyED08IhC1
+XLMPD2emA1ZO+90QZxZsQNXxFVBt2nyA4MrHCToyE1Spi527MYnbJC1yVnBh5gn
TvCvfweLz2iTav6wj+nET2EM1cIzKL7TZT1YQFtJ1vVHp4N+QuN+7iIQoohOpq1o
DU5dauSM7BmHDAPoD44g5i8WQ9xdivpJGuxxxI3JDRUOtyTd9sUME/9dGfAKpT6p
jjxZDqiwwgPcbyG0w+gANpFMUCQZGdFjyDBSnbr3WkiioJFFvZMYMcj4NoUfJKmZ
vO8a4Een8VBdg7uXJtw9LJ0u0YYgcPsB+W5W2AR7ZFh/RI7QbisPoa5sWKr0QdgB
0kW/eRhMLlMix0S4hVpcXhPSCFb2uUaM26nuWNsMpuPZW5gmWEmDvpvA+e/kmbjc
zZ7oiHAxU8x5OaCXIYq5WDti8kZq4uaOz9yclm40+IYc99IYMTwC4lWhQDUwQlJ5
K9wU8LaAOwkG91c0T57Zn7GitmRIg5x///TYvgGTPL5SRLrTVx+2VLXYVFKwu9EK
leudy5upQQKJoQhQ1QUKpuOfl7HFgUriOdE+7fE9V9oxtzMHAbI6GFDWcxR0O3gk
lq2Wwocr9RwrLsWErmUqhtxepgYbAFY8Qr++A1e+D0muO2xGCMrhw2IwnDFIK5zV
JZO6nniMO2aOofxo4aU88U4pnV/Wt9I7FcVW4KCyvxhNzXZyKMZoXeQq4i66mOhg
CBkw8GbdRV1UjWCckrjS866094/+eSmy2sg+WDRYOW7f+4n0QTfPcYAo9nmzoedH
qZmjElQSEgSPIyAZ7ShbAAO5PkzemBGa8hRwy7wpKYNbyEOIYDZHVNHAkpznlvC9
MNszB8pTwGDU2huzuOl+0e2wZJSKgXQkY+WIleUuqcDGyDab9n0rz0j9oFel/4Z0
rB1vxMsAQ3kvuRmDT3IFoizK2HVydyXnlIHc+96F6pNzYUqImcwN13zEj8UmusIJ
1tjkeOSTHXs49s7TTTN7dttxkRNQEXNVuPKy5Tn+JN3KbbGfYSxdO37Bj4xmc2Lp
mb4JGPr85ILF2G/PmrjaO3kwRQ6g+X4jTeAH1eKed6rB3+yrnETrV9De5ek/vYet
ZG95+I2Az1B7rMBEFPZBWqxQsaFp8XHR77JtXTa1a0FXqmU3t/1xjY88XSF2hgZx
2oH2FcTTBkWaf9cQqRDi8oj37suEbLqt67gaK5H65TeDHvje/7R2SFbnOpl0Uo0e
Rn7lhvlHaAk0nQY1hyh1i66GBjQ0eSXXkFEAfIcfu3KoXF5MNIgT++FsK1msD4YV
batWeHa+Y+BAIYVnVy+nf3aQxy3EQ7KJ+5zwEKmn1vYDIhvRqWMKnTKpGf8N8QAb
q6FtvbpbuIm2DHU9SksnZK/WXMZ+Z19A3qKO5wtyYnM/XXkW8rd4J9jNYTzJCx7w
MNX6O8B/iTUCkpOhgnUSeNZGBIHrkomnwccTFRG4n50F/XZl3AFaKHSu2fhSD9l1
sk22U1lLhcES4bVWlkYlOOErtkgcurFBGIcLT0F1SR32AY59wPR33kQV21nr/7XG
PZ7NIu1LH3wI34Nso3JShoupy0jxtH55QfAJFtLsla/a2bh2WY0nv9aruW2OmSD4
HngqR3VahWMF6tCEiO0wlQPtsSc2QmTRfD72d0iaIbEOYpMpBZ6S47NpJMtdLkfu
nX65Q78xZlo6wavDKrHZW3eoBSN1eH9tfwC8CmHk6b5MpHRiT1wPhdBogWznWcX1
DEcUioUWlhsPMhkxL/TxHmsRtBwHrdFP4zenCZXb7tYaMsu8hFdofhXoXbo7MAwv
HgypuJEyJgkunaTDT1T3cozkVUu1pcvFN14JjvYmahR7jat4isDEIXzDyevfa2cx
FFAmRQX8wbob8nuO+ks93QUz/thnRNECfPVZGOXvc9OTWL1Z8XucC3Zk/Zt2Dd6K
KslK944K/C+Et7SBOsQJ9oBXVKauMAFfzB5uL0GxsQhPaK7kad/wSDQUbV84W/ae
CoJ3e/g2fV7Jp2dHcVxTbV7/+BE76i72nh6vXSHJaKx1MHpu4LdEfWUmLplPpL+H
ID6rEgf9GcQ6coYSgpvJzQ4hYghw5ia+pmVS9vapkhsHnEO+Sbep2/RobZ3D69Nh
8PJ+W2oQAlD6DCYVU1vj7G7wctbvLQjPsDqipy/qRHBNixA96y8JI3ZPZcnNlrOJ
fl5DC4B/AD3xT5Gkt+Es/lwMHZsZ5RQxsRW0CLwEgplJjQ8G0gIAvBEHOSOKaUhu
XDKLbYtUUCnhLIJw3H6tWMERsYn4h5zOp4j2bxl8zBpuOBVsWC4XhCVvR1Hpr72n
OsHxLSCmiStVaaQcDeZXoDdKLn5lhbDwjYnhSUDlL5IAw+W4Ozz0KHpkC3KTeF4M
HTYFYJodW3ZPSP78ovzY21dQ5UtvPuwxt3x561IuDW+SwGXjM+RbIStDhh2J0M49
dCVJgnwxO/rH6RJZa+7lezS6TgkRvptGA5oTBHcF+vtC4HmYCoUsHBIs2bbeGi8V
x2T7dpPj7t4DB52MYEGH6HOd5qYq4mRiCPyPMCLUgqkSoMOin7Gg6/ss70kGjxwq
DxLgI2SFwvBXczWTYIJV6mXyu+h8Oaxom94EBhuaWgGYcRH7xcJE0XPdALEHqNWh
hdHhLZPaHqEzZt3vNWc7KR/GNdIbTc+0lY+9ClA+Va0965q3MB8IhZC8sgOtqI8q
c0tOehuV6zm89BXTNsJ2ICljp0iNuRiga7MjIUH0V2UtkigAmDZiOEM3irez9XPU
5Znh3wRzeaV1KWpHe3X+ZlITCR2fvkaH1eAnBqj+cmM081UQpUpUMAZCknAYDDA6
8d2rVM6XjgjK/jn2GJUQbW/R61hw9AZ+M6itGk2bV9Hq0G2Msv04y3cL687nqNKV
qnpduGGUmP+LJJpBzFfEzp9eXBPpL6zvYMeji2LbXP7XbNVGv6HjOE17PPEHyWxA
7wXvFSwdWGdf2LDaFQIJfoMLWFn44KpRT3ftj9f25OAX+/bS+Oz/H8Yxvp91Tzwm
Du3OQdE166cMk6OXYLhjRHqQOBF7Otr16UIo5oQWuDYFTcAcUWfoKkoFNdmqkFQd
+xvY5IPbMjADpr3aqxpjb1lRMqC0HDP+1+JFXsU7yyx0jhHLCe59/QcX/oDh3ZVU
Q7iKwTOIJ8RpWrHMc/ujs3Mq8QS0sIeBFTI/O2CuJ97mN+J0SvqrmX0tfqg+MIxo
9o1gzHcrKw6tWhwUXELJRdyRSq7G+gA5EQNi68PDSjcoD+c8SOLQ63FxbyNiQMSJ
6fQEW8xQhm8ynCX9SLmHwr6qd2QoLafvC5i2xqfYL60Edhu0Dd0Yw95h4myU5xYN
kM4G1cS3Q0BNU4ErJsMxffU6JOuecvc4SpaLa4aniZ9E52UMgcv9dpsVY8nZyM3x
HAM4B6PEWZ5X9dT6iX0H4UtGxkZZngQW+zDO584Qm+qs2BE0ZEE17iWnYCSTwIHZ
UsiRNM85Ybe3TsvpLHxhauAfkrOUpuPILrzA7YEypX9NYgBFKOebFy7+3GjfHwKD
RbTaxJ0uMAlZdD+KVGybzrS4PVUTvTmaZIhLeOQuUMIbpTQy9P41ITtVWHWNWozc
/ufCBGiKHDUJH1fjh/hm9niqzPgWeENIKiMIL3DeyhhJmGAg8D0ulr1g4wjae7tb
dv2hgHrAFsEEEz7ebrpXXT4PDplk9OZKa+jUdbySGkcmsBFpEy6XZQ36mZVsxckT
P/s9jp8tnkKfz44MG8pMv+UFxahTN3XhmnrtVzSskpv02jvDQub99iLa4RFvQjsy
xO8++U0TCgY9YWKIppUxdaJJ1Xy6hHyvL+klwzFu/+Ef6n+DjcCu2iY2bbUyuzh8
Os9+1Y+xZyq5cGH3xZSc+Rh+IHEytGFFLEW7i8oF1yBAV28PSZEC8zcZE7UTST1f
WqX1ZhnQiP2dKKsBsYnK/tw3DyG1k1tRnXSFaZWYogcNEQ95NAIL1DU9vclduSPl
MgRml7jngTf5fmVGsGYN1cHCEuOatrnkyNcpEHPUbPkUA7o3rdavRW1n02saJ314
K/s31b2kCzRNzILZmQyS7TlVbpEJwJYy+PQGgwDuBQKa/nweMB4ihlrJsTGYFulj
/mhNrKiWKYJ7t98gCcrjYRlL3dTtP+XsxTVztMnjZ8pHwkGzzoz4kjvp03lr6XU2
wL+9t6iG2BOTSScbhIpKmRAXATOMIo+qf10Xx2WPVnNwGjS4O0t2mhNi6rItk9zp
xLXCsBGdZQ3PtiUOvYefW8uhoFgUwfDliVRcqHBt8UbQFgIh5krjQjRbiaJ/b34K
xIkVW7cLX+I0wNkb95eryAkLrkbx6dQ16fNElCKm38bPzWxLQDg7JnjZRkg0g06z
3jHSjM/emuIYaz8+KiT165g/ZcsemxfHCkOET+lCos7DmxrVC7uM97hZpOh4N8o5
4YIckMyIMRnMbFTHCe1LZhI+XVOSIwsFLW2k0dDoaCH8iUW7LQubbsSGpbXXfc82
5L4nkfkOE24/8txabH56fO9x9bLvopxA5g+DPFLWv2mhR2i3+Rp+Vcuehp5DtJzt
Z5CxBRn6ju+3Be6cr60cVXJbbdgnsVElOmNN9e1FRPNrhv0HAbDWkFNay6ugG5iS
aA+/t2q+vZgXLg27hlwcGxPv/4QP7vUVysGyXB72qMvHr42rhq+0pV61GnJYD7l4
rU935ouVIammx+izCwC1Ge2X/CSzLLyAHfoxaMArIAzmjyDupT1sjXYm0RcFovFL
yrXbsptoSIvAD/tWB6u90uZH0wMBPMYdKUIPR6/Of/SR3HmxvlxBsQz5++bWx/Iy
bVg+R5jxH7UdtbBAzF4B9/g6Bul4tOcNK/uahJ4/sQz48OMlBm5RcaSS1BwuaXQ/
r3ZVMyzZAWZ20qIbXcHdQvptloYHZRX84Vj+D8NZQL1l0lUyq+wbrRG5qIeBp2pf
BfTiZ+W7enC3SgWLXikKcDggyvFShkbjoGPW9DXI44O8UXu6A9NX1pSdtBkwOBl1
CxlfwLpxhUvv5aS8e38c1RphCnxNSMe3D9jXxb8az+TQaWxqURG6ZQomByqS8xef
pWL6ECMkGBRWTMmTAiMXgonGQWgqPwEeUUoeIlKX2yaQwyeGxEP1y+MCSv2P132H
YVE1yNQP8f7L6oXBHEMpT19PSEDKsPxp+Yelezst8lwPJEahuQ9W0v03yjVpQw6F
D3FC0CPa2GuF6PjYalzVAEMoYm8whYh6+wcLwQqtO3ltKcZ8MuLf9I9xcNZGmBwi
nEU3ozAdCI/Ws2rbD82EM8Rkp5uberc3b4YjWgpmbQrILt1JxjEwSuXYC3xiGEhL
nwX9v98Kz054zA1qTbnpMXzscavi8jh5OhhNdtn1sIzATogNQ3JcGqFmjDAuwqmU
0up1xBJVEyRaHdZqvD19UQqM3mwkYUv+IqVCqip3CWLz1Uk4LDCZTFVXVsPzTsab
vUgKN6aUBCk530/l3GkYSfBYnJN4lassh5M0UOMInvNxSKC1DEhN+BMJDimKJpIs
0O8iOCFLSAOuxfqjd3Jjp7CerrkHx6nG3cwsQbybpDmLCVtmDOuDyp098jctGhds
9RQfm6BmVVSk6fsZ7jrPsDsvc4jXa91NZ+UfHvDUlPj0+ZJvXv4NdC6i9YOWD4jx
RIRh/NdRQF5T9lPMAZQmivJsenmzR1sjzR58h+0rJF/daOKwLQzg0lGqL9g5D9ie
rMuDcU64bbgdqI7VbS1E9u5qdlkxjyph0LVS6aUMYY1KHWWVHMBpwcbEHSNdEx+A
VWP5Ongs8oRN+CupTNZ4Yhazg+UWote4JIHPMjHZ8y3FrsqMBtxh09tV874zTQK4
fJxS7zLOc/M67Q6UPBePOpJMM3gNrsrkGCFCRuGsWr3uQRM6014MYYdkJwUkJHG0
06gSwfvG/x/A3aBYBjMUCCUTkTXbO+2JzszxgGq42HFn74qD+5dIa72/PlwVE81v
PYGW+ETWLjtnlCO/5PFtRIW/7biuAiENjsvme4m4KEJljOuA5fEsVIItxcAaksXd
zibmfzH0aIGog8BRwBzM2HOvro2gatb4UTSsFsTOSEPxjNYlbM6j9a8UeKJKnNKq
RfzGEuNamlfrJyAn9oCsRMlh2rqTaGSbyW2v09BanBoghQOYaOlG0Dk1trZ5snLH
b5OsVNZrYhKEkIwPPsn3zf5oBGmKwMPmzbrHSNGxJoN2dvvFu2b0eeh/vOT5AtO3
J8/Z+fPVkky5oeXX6UoMQgllpv0EPgSvvGdudG+6NpR+8JooZcRAXcVuDpAKA/df
gqfikyZ4d4AHIEu5+Qd2nswzi+sk30QHNfHFqG5b1tuT2VYbatRJMIWglQa8jnBd
rI3Hflq7pLSd6Ljn1k3JzFOBIbubgg1y1ULKhDzTXT/6SahNwCsdj0skUD1hX1mv
WrBOEhNSyD6UdNWO7yz2MJHivFWgFPqBv4hoQ7iqk+Y/we0GkEBPjGwG0SolNGcR
uO3ffaf/m4hdEU0sWo5stROgwG4tVjNtl8DoymIcyH1rDj6YALvwK58WkYWelYgD
aE6qhHSITxdTFxS9p+kKarq5x2400orAnJ5R3AiGfdbaBmlKifwxZ2jJB1fatibF
am5uK0LFHwMYhwgQy8WDz9uun6+LSQ8vIE0D/LMEBdZ7uQOxwCYUjvMbJNk7rlFd
GuC5IhXB13S5uVQb7X/IjtI+LQNfeMtj6bT0RL4vdBzjVP9nkyYKuihGzlYpe29r
i9+EPrmSPGkt5S8vtvaIndpZm3iZPBzqMHds5d4hcATmWbia1YHBmRo25ygaLfoI
GNp+Gtusseor0tWjYtonL0o4YsfUnYU8HAHjOpc/6/67ft45u+58860YTPiF0QUa
NBPNdGTz156A2OXhQpRBiTiqaxCVwwwNMiFLrqteyLhAJm14CMeuBpD5wVHlkXX1
UYqxIS71l1VgB0aJ5O1lEen7HncMEJGx4cuU9B5UJW592Zl16hLsZz9bDJjg3un2
X4ufzUACIiSJ6uSlO4zthkdgD90yvRMu2xoOmRCX504aC4R9aCRqk6HCmSOAP6Ho
LD9Rpd3p3O4rqx+OKj0AaLmgMS4qQ9aATCz1+6tKWmO+7GB6+s52aR2mpQEEJo5q
5YrCRh4eTVodysTD+FjwvLW6kOmtgK0S5tMq6KQJps9iJx1IgGdDxnDgzcNbMj9A
DOLJQ/skNOgdaILFX0f80xWUTUYVh2960Zq09grWUOQySRCS+HMt9I8pGy1J1vRU
v1t1B/HF37F5i5VuWz222OvpBUYzW3ARMQxA8pUJ8cnbZIye7KjuynClbJlAMkTf
e40IVhstA2iwsKeUGydMv2TNe0anRGHaBgiULk4nnAgvZ+rIwTY4a5RXG/vdqN71
XVb0RN08ERQDG3QJdf6iE2UeYmn6pMBIxiT6Wtoi5atYYzAVVjyHGaSzXV0K7e9P
T0aPfM9oQOlGvLZNiyLa0WYAVN9BC09FGzCEfvSinxLxJW3aOpDEWGhyAEtATNWn
p6x/xAKFS0Kl0QsC+xs3BrX88xJviZON/S1jhsOuN4aLHrrATn1UI8W4jLirH2n1
KBqW6TkaA3XHIYa62/EZhAKvONzCBZ8mATkzXk24sDtQiAv6cpbWuA5KgIwsdyse
NNDWeTKLK/97mRFM1EdtdctsDkiJymBNNxhSqVokovc0JsWBVAMUEYHIOcfZ4cOd
YcY626eGmlFxKItpoHG9b2+zZkUM6l82Y0QSmeqzEJ0ROVtv4d2fIpL0CWUOcVkq
pk0ylnfwRIZLMxRqlOtAmojNIEBTCUFNk+1bjBuIbJiFB8K1Q530ufg19eERjb38
JA5MH3nnoKVPspWNHwabGRXll6RFqAb3BHT8JMlQi6LqZLHT7ivAyrFIP2h3hnFu
Rzzk4RrPyMbe5xVvK6gKAqzaaIhfiAZo70JB3LqxewZQD6DRuk/Wk/DF4s0WwCG1
9oFLa7gBcetrRveCE6bK6eXKkil+c5kYE7V6Vg+VZwoklYJGiEW4p3GD7qsT72li
jnWJzf5+/3FbbuEpFROuIb9IgUPw/zxS95QuH3Uv1Vwj00w3xU8zUYhBzRDKw9wY
1uTMWxzG3HsQIJkjqpPAfKQFZLlueHBwX9C4405i9I0pywjBpYlQKNEfJtGUbxBB
GY30dPJF76z2GDDoOaEzV3YILKFFHr9B0QqeljBHVY7Na3ElekicaY+oY70gAui6
YmA9cqJAYMWKk0e5n1IcqAS3EU09eFdoFW7zqZ087dQf01Quc8ehgPCZNVOnmXtI
F9wfDVYGvNvykaov/sdGmqHWUAZlm6IJ7GeM/Cy+D659Q1B/2BnjuQey1ChVTUwq
8yaTKkgiLcNfhYQg6XQht3BZ0/NPP9GklDyJpCUqIKsAsKJtQODKQ3xOFYDmDIFC
kYvf/5D83wDFiR+sbL4mKOkMSbxnGZ8zZkpgO8sF/yCGrXS8XqbusipuQ84Zqsm6
j2jclupTsgOk5ucNcCx4CLqO0yeGOXIGESSqjS+vi8DGVA7sqoFVvoIyWgyqMTlw
ZsOzWRlbiJs6JAcgs4eI8jkq4/jOh+OzOk9tToyOooKj4UxYQq75jvRwRX5SRZIF
UPby9Xn6iBCyBFL2wf4detCXZe9IFFXI3i4XxtWj6g+CoPgtJ8hJ2VPzoU2SwOKQ
LxcKvp2Fxdc0KVA1RDLE0HsUPA+E93hhFtVxRJLJ286/O6rWa83d4zpXT6i4CY7p
1Aqnu9BXzy/6xrK+2gvM5kXgaLCn9dTdOb9y2Ku8OgS9HuVFE1fnb4vFy1uIjibW
Zykf880UQKiHcDqhPZ87PVwR4N//fvY+VN2TUVzmxyJ0VU6RvAvprUYNShLWBKcZ
BV0IBWK1kSOGyi99wc/cBRShFR8KCn2qoITtet3wVBpTju0OhIou6WmC4I7llBw/
a+0/b97f49YZwLFvG1ldSwDJMKxz4gDGlRTnZHp9XGbPYLfYE9BzcgLFkBt3Wx2/
IGdiy3e/RYxtrTLqlJPS4iY7iVGp1F3VoOPMBY0cAPud1fRonrRsxhHvb427KnX7
DOkm76miQuoqZQ8WxWqcSuVqf0TiWONIOh53HFJ2NnU2+N8KLdZpbeJt4026FRVI
Cg1htamGMOoazTczFry+VtwHKbtxSgoWr4Wfzz9MX/KJWfxZFCXwFvRfYZ+TRNW+
3B9QNoFDJV/HSXCNfi5L+3Z9sqDoVKDooCGNDjjouVn28P4/H186/1jC0OzNC+EV
9y3YixQ2M5Ev1GBu9Ae6n6SzLJlw5WUpq9US+jrZlmhcIdKx00a/OD6GVbo7OiGo
pa2HbCbqXViI5k+uCZOEla2jOzQkQwxyQcoK1DmklS5vtl5TJCJxyRSfXaBvy80i
P+xPhx8pGxRxUkZrLdEUMwbpNCD7lJ/f8EXLRVAQVNS15ng6hivrb6RKKpI2g5wg
NgO8j1Zhv19gmWfB8lSXQ1y8YR3XN5GlIsKKiLM3Jv3ALa1L7G6mzfL7cSUQW9Jz
+mTwXuKeo6Dijseo1x+9WsH8L9Vqh1YmWn+o2ZzbNy218vacBYhyKZUYQ6AtbvRK
hD4VVkAilm11dil0oyzxyCbnan7wTvUuY0Jc0w8HxH/r2aLbj5Ze7GBQpF6e9vJQ
Am2Gmlyg1lvPf6SNQWO3Qwelt7W8t0ehZZr8vpw/KrursS7jP1RUtDYUfX/BnJ9I
pGGIYragS1bd24NeLOBR8An01xNcA5o34CqCKdg/Tap7d775WOlLsTYVuJKRT/6C
SUncvIZcVS4ZwzIZJWVyHHLVThMPsOCfzyDPJL++yO3b+tRA8U2VroaSBmDvgKVv
iqU/QlOwqwM0RhOpJqYNTKKa8GagXxsBgKr7s1G0Z3nKA9pSAiVRlx5fT/i3CGIH
BLkH7mxsV1uHbwlwgCIzXIk/gMqCnVtzogYheKDIUVuNUTFdD6bt8KhC2xDG7ZNA
xYf0hJrN6ldUz0WwfeaHp++OjdZXRESzIdN/SQ/FUddoU4slYRu9iOn19hFW5++6
jnvpjc43z0jXHPXmYJx+OqLz4byLtSbgIrW8USqDYFI4G/zkPyE8B+y5hstCiOQG
uPF+rIwWzHosT/PExL7UvAwk2Euj4VS0yiEbrz8XK6A5JC9YyJoZgAeLDiAM6DZf
aajfsvX1+nJKuj5srgnMpk6PhmRBWBWNF4qb4iEFVQwSRNi2ntcO0fVwBvT7vctW
AgxVlEKikIwXQgE8WsRcqkScinkVvI8rtY0lyg530T/npat5tphjeEhGNOD/myIo
rdcWpDK7ueXglcEMxVZZss6tioLrite4+FexpPajQfNp2IYv343lxPHoqfKpUUfN
LsJ+UmXoCTC7th86WKceYfk3mYnKttokzwVkr8f5uBnQTLFwcQcD7euzcGk0fCbE
yWmghBh9fZZgR56d5Bw0QlMgUb/oqynWIy9G9jylcoaPQXC6mdO0x/Na4dz3WWYP
IEkfnhGXivA7ohS4elsoFzH/NX2NeQDBUv5/4hZKftiJ5E/ngQJkUX9gAE6bEKis
iyNLjP6tGV4Txo7n+Bl3JQuc7uJ+AuwCT43uKF+J12N5riXl3QYoS0qLgxk6vPpT
4RtPNsGdW/xeS7SbGuxdZaW1wo9IkZkxg3SfNMf/Bq1qdQ5BlbePKwrCdzU0PD5s
2zpXJzlz8K8EOEy2RogEA/ZwOvXoz3qX7XL04p5yp19vMzOjjYs9IMGI9cacmfuR
JD7khrmrnDZj/aAA26iIYc6qhavHVG451diMjUfCNIGMKIkMHB9nJhKvzvBFlmAg
fIPKj0IW4EgThZfFQfzDvC9cPwIMNBRaIu9vkZa39VvLTZGTy7giu6rp4merIMET
qpS0KGTqE2EVIGnCrA70G/jopDDEbFgNeQz06A7ztGeUvlR7BmqK2Kq9Ub++RjGX
IUehmGLSu+GEbvt8eSJIBguemurXlfNrx1WdYaGDEABD55y5hs/+79EbtaiZJRmb
i+l6N8rAvAMRG6XIT1+kPCvbXja5zKWRG7IIWcFdacC+ws3xaXgdxMn07/sin7v0
Zi0tW9pkFpPKa9J7kQPyWSHAAINp+E7isW2fyvmc4nujFJiKH833jykGXAWFo/cX
Ud2W/LvLYhfalvYL1RrpZoPWT0LA0wh0lYm8Dm/KXtVE7akMJd3jenvhQtneKMwB
iBNd+n3w/y/3oxbGUhpdDhLnPNdqNHHhcB9XX4Ws6T54VtaQn0vwNJoyI6D9LDkl
5Zd+DfvbA6GmtbqwT4OfXgA3l3DIfR/UTEzTl7S5U+3Bf+dUnyTv3KXe+eyN01Cc
sXQTPysTZwb5M853Nva6ss6GlqckX3pE2E83RySi+eDJE/ONJtmWx8toQeLr6cHk
mviGNNZd/rn07ynywadXGoq4lE+Pfrxs9Nn3I9S67N6eUKpl9C9hCv7LBFNh4Y7R
pqBAQut22LIGN/apzzdyAweujWUY5n+rvxVscVIl+e/RTnN68HW1YObuwELa/Gec
iubtnxnYuTfWWiPAULM0bWEerVPQTixU38LyTTqyjUhmcKy0gea45qP3kD/zF1hu
XboPjpKCU2/SD65YHfZKBqLUW5xnuj/ozR/iRSM6QjJA5xSzaNl/RqNPm8HS+Cfg
H+FvkaThENEPWslk96Da3gfdFQ9ikMRD9JegkK1o5czkmnZ30nScDj6MybqizE4k
PYZEHo6oddPssiIr9XAQtgy0bI1rga1GV5i5NlbGw92syHlYhv8wyJIxquUIUYWd
LaSHBMM0SeVAp06vZFqd4/Fdwsv+loYpQlmK6pURIcQUt53dxsC1Fj0pB/8nqobg
C3/9wGu4ffWKHOFUm4AdLbux7rjqhHkFDlDrunaSnSOnZ0DPIV9iKVhdqs9FBTtv
NkANXZGrzNH+Vgz7Y3OZ5l1/Hr2BKISS+S4rLkoCwK9T56hwnPQVtY66eEsSbiY/
gMP96SGRRJSFE7L5YDzWMe5r/HGgpu8tZ0NYVyT+L4KP/Xm8Swzejz1lqoc3akZr
GmjnjiUIcYxuW9g/hZxZ7VQSvR5c4Pmuwh34eEJa4apwUskIwOlTUs+umHfll/HH
FjDtWri8fr12pm2JQtLDyVBN57IEaQ7SOkZRKXpDs3xbQ8X/FKcbaI1WDOpZxzSG
wkL2wygzTs2uLrapzg0qqljM68nmHLkxXKongL0QiGRxxBaJSo8aUABKLG8yHu+T
DK15nvJyJ0KZ5Y7/qb9B+5YsQ18sjxJlJdzt1hlzDlMfHxW4M77I1GHNbAlK3NGe
4jth9QfBecMb9XSYe3QfjQoNdkjcWeUkXXbjmp6qc+6dZhfHgAIQ42M7lFZcyfAp
aocHedUXJq6YOGJ3L6QiyU88FQwbFN4QU6RHm8YyBJvhrax8d9HA2exvXrw/l2I5
29KGqfv9mOPeF9an5q5mza5Nu7vxpeZvso8AYjRH83T0QQU76ZecTIpR0MFTUF3g
6I2HTC6js+HpitRAykBBeYdlyw+rKtIFKlfKrfO1YbAe9HPB4W1emKkCUp+nKb3Y
DL7ePMqQzeNF/xk9+7BZ5D1EF49946nSyYit5Mh/pmSQFawlGiDz7AFJeNkywYns
dRgLvYGvi5T0iKSnJVF9HXgS9yqvPxLeM4xUpQf/BYf37exXokPVKJfyD10Ze9fj
EtTDZ1llQkPt/U0NCC5oyifcRYYpvDf4Wl6LL85vZ3vDeR0K8zCkHWzTlK+iwE38
/XCM43drhcAmSy1V5bbqKz7SHKTA/xji3AZser29BmwGEzg93qphi9csi5DWu3gF
Ip0hGZWOeIlFFgYf9ACToQnJmhzKXGRVgCDk8xfOf2jDi0M2hu4SJ/ObZB9cHbPe
njPfsIg8kJvU8L5JnoHixu7UtpQAjbw5dFsyHirRDZrIYWzNvLV9n36kDxxqbQgc
I1z0SfOwspJqeizcdlldaT2yuNgTp4QR0rFV1lFMwxD1T0vifVFFy9XThqVq6/Fg
O1CdolZOm3X7x/AGuL9f8zAto3616S7gEXnlTa+8DGkkHNDpTGHfam20ewLjAmCr
OLRa8xsPh5yhFODiNpq5sytImq75+EKNTFjpWmDI3q3DtmNQ3ikVs+nGohUbYwh5
n8flNF44QK5YdXCOCopRuNxpTPLpbMx+TGsKvLcYigJnZPEW5gpFIEUHqlrkIt8u
gBKBTQ7WZGQ7e5gikaUmgjVxq2Br9pyiO26D6NGMM6rW+BAe/5wCEriP1EILP3r2
WRwhRMYF7TSkE1xFYvivYw00sUoXHWvbm01ULUaUbxsVZpuXOGB2gcJ+9HFfiwuV
iaGYweaQgefaSaYbCw2jtJe2NL8Jl7MBTv8/+cpVEuNaE0+qgHRArJ8L0vQUO4lo
D5DRvEejUiVDGxsBh8UqwEKVWns7lJiZPXP/sBbKLxdnhyej+DpDFozTLyYgZ1lF
MUXs4GNp/uBnuIX26OXUSQbAf4Z5SeG/6J89P6tn2MT722RS6y5tR8ccn+dQ7ADT
VOcgRaGxP1dQVi57j3PLGHW4ba1x8zMMOokpaotykr2eTMb5asomkKj1bH8WRqrw
/HHQCgZ2Ja7enTbxDEGq/mJnxm6JGuyG/1VMBN9lXQ4CTt+XS4DYQFCZb1ZKWOfj
YeYX4u9fCdx+r6ijf1ffhPSVHWBrHravLUNscCguHR8NFAb2kNAkHhnx2HS443cp
WKbaJ/9Hmnx3PRsLK+jG0lJHVwU+r3Z48JY/fxyjSd3DU9tLOwdi3cxBBLG3+GOw
ow4A5AYRDmllZe3Nghy2CgtPi90dVenz5gOGLf70DWOsSGYaMPj4dVZQzppjWZii
yDmFT00mt4WHqBdoKdYiQIZC2+yGPmQUgBkUcb4mvtDUCYTZI0DDujB8wNFoNM9D
cfwn0nUuIeKWXJ5o04NxzSQ7L2R+gTJdgohdyfwq3OBLTcjev42QA2eeDsEMLHpr
Xs6OAA4wW87Izy4+PaViWZiQSTs69y16yKl/jCwFhyPzGTalrpI2Ic76wT+NLZh0
v23eAkjorAIWYHlFqcIt+8Bjs4EaBqUORl1qKKmx/9449xJBoW4mllg21FA9rSBY
YKE5FNVLAdD6epJp1VgqZIy+QGY9I+W/meELfWLkMtw8KgpImwkVR0d2PbrOxIuM
Zya2Jne4RKcQe2kp+Vgvf039mKsDqrfZs+Pq3RgxX2pvuAEX527gIJmRSFdlomo3
j6YCVu9COhI1UzKCzdj5rnMtTnKBsEttl1deqNWuzzhGacDLiJSttYssC2aSq/rb
xeiwm+EEYj1lGexrVCPx1xhFEfHPxt9APHyzY0nV0/afa2K837lOWZ9nXoaAGUfK
9F5yHiCU5wgLMCdRclvHALRUkhfzuRF1zC0HxkBR0onS/ZJSBiQ+pOn5reMyY0qH
T2ZQr0tLtM0upBOjUYKAYvZoW2HRzJhsy5zIMGwgyNjO49Fr93NVKMLLS1KEhLfy
9vYvhIxqdwbSV9SfBEWHSdqDsFVOfbtqsFJ1B5dRKynz0NJW6b+BEe7MoYXvhZmq
JtVBkSWjynoRub8/VRS0vFTP+XvcGU0hyWpktf2+G7B0/KBr+MczCj1qG4LY+HE6
w9PA1fx1XlE68HUrL919wyCRlhuUBrqXUaGpcf9VLEKJ0Sv5XNqNZM9Yi60xd9s5
XM7GqxG3DEIObBC3cAMO9istnE8+9sHMZrTHlP+8oyiTd/lBswZI7VpBL5O0n46k
kzfLZJDy8Qa8p+NwIhHL9sgAl2hyzJ9kmkUa9mXwhVatQ5fBLCFcKHT8pIC9XWY9
CfObieZgvmDbFdobKSNL5uc2N7LTqBrVa5gyt/xAwpOgLj8OIai3TmN+FzVm7GuM
G7bb6T9M1Ba5zvC6WXrmS9SoeOOoo0rHz/vMrsfBjX5gvFl4Ce+AhuBCatQUTehg
TXITEh2lVqkrGoqIiBk2L7bftcMyUMx56BCNEj8iy0r7nhgKf/0G1uTE9zZXecMu
ZG0pjGe8zjKkbnJTZpIPn9nqXC8jk0qykH04f5nW5q9s5KEqfMCyY/Q/2sY0iTpg
3IAFIFt+lTMEqbeFG0fTAUJeL3wr13o1aHmi+62GuYKmHe+O8Bh3En33VC2DggLY
EIS2idotRjqA5Hwme3R1+JDgF0cDTbOPmC6mwVA1y0cjRw56goqQmfuHAK0+j1sd
BMVBelPPSyEqBHsMqHURMkNepeYWBM7fNKJSVasd7m0lOl4qOHbT2FqjeyMVjxuH
ujE750alpmrWHtqpmWiN9+0MjNLY/bHcF2j7mC1dI4m9BUy5QuSpG64m7sdyr5eA
fpQDq21GIy6cIRN5ERotXWKgloO2edTcTj7TIGjp2AskNifFFQut2ep8OPRhtIVL
4l8e71LsFqx+mc1ZkxPt3OqFNLye1qNgxMEqD6kZfrlYp3pqwhMnWXtPenAvjoEr
kzL9fZ/o2b1j3xIwlYwBKwIonwF+RluegqQT4QPvKd9BazumyViTrgrl1agEcYOY
jUwhWD2T1Htvpl80ZQ1Dt2kj5c1k2r0wrq6ie1dvq4SB663HqfMd8KlLppT0xiuE
Cyp0MQUx4z8cPb/KEExZhnl7SYPe7xDlh9HyjzHxbbYhGtqB2ULVhe5tdngYD7cv
IPyUYV29p2PHGROinbM5n+I3ykAp7ye25H+m5wuvxGvlHCtghqwkyLUnY52p5lbG
oAe1yqmlfk15W7AGLy2rpkAiwSm0hf0AHRsVWP/VoRMgO/qZdTW1Bd0YisCYBm38
VMFCUBueb4N/p88z+5OjkyYUx+pZqxV7FIqJ6BVvfZlH8kv38SJDCPJxD+oD2RCh
xgSs3vs/sAGMQOBS1BqwYqJqQT8DJmjTvBgyZyVTeN8RE4spnnKMh/m8ebAG36o8
6fc9xynsChDYE0Gd6AQLjV032V91okua16wIa6cP22bZ9U3JrAQaQ4oxPKwn41+7
FXpBjeW1xb65xRK6YN/GvwbGQHLxQkYwZUfzqmpJXqNCOKcmkTtIQIHMhywlalRa
/sm99GNlroKX+riAqf9MeA/keHh+wOYmafBJaRoqLQu0+gwxlIqb47qOl+dmiLkE
Hav9RkgsCa8BWBjtlep4Bd4QLrpi5o0JzpnwdKx8xXLXqTIgSU03Eb2UIJTqCBrN
VbIw4GZE0oqv9Aa0YsN9KI4o8Z7J+qEfkwz9Dff8I5pDMYx3I3MpXnaZH0YPYOQQ
NOBGI/2agf6cTSiDCFEzbgiFiyaP2Uw2t07X5yQfYAEVYFvffBsjNSnKt4/qnPlo
IrXhUu4+gKLcg71QgrhQMHSAs0PdRKhqqKsUO+vWHw/8bxfpRQenZuPDwnV+qomo
5R44vijj0dH7ccIQUxh7dyDnULAmxt9SdXZbbSM7sJn09X3LyBhAKN5zn1vJageP
P7fLwfWjSQEapRwnKAaDqnH3aHUQZw5neB4jDlpi0gOVvYlgmVJk75LB3b1B7z0S
1UhdTWRUy06+vlOZURoXBk+hMtLFXYiU0X+9hde0mZXcifZQyosk5IcFuLfX9hr4
OT7+RUe+b2EPzCjlvPyM8fQGlqh2Vr/aNqxGAkOvUXpGv72pkcbAa7+/5b12cEis
1XchBte/QIbgWh7JJSx7R+zkcf5QMmBtvWiAjdDrV7W2BBhhulOwu77Uz5k51b6y
WUAe9nAeEbnQns1Ee2cGuukVASQRkzDnwUbIO2TnsQJk020zLhUPDPa6NG+lRENS
kU2sG1z99P+XBSjKd9B1kNMX/1J0C1FiYyU8EtomPq5gy4gd0x7F4oVl2Rmv+got
+P/Rl3cX8chQUMJaumQGTyXeRdDlKByR7U0JKrytqWTn8r9ObGdVkZ2ImtXuIzYI
zs97UAroD3quvpWvg2oV4h3auBbcVvpdxBZGWofANogLGfbdyuWwTP602Z1Bor7d
ws82tdElTMHO2oNI44kE4WfM9RTPTK6vz3N5qswrfKk4sFCDzKaz26CUoM1YFkmF
i3r47Vn+R1ibcN623WEJMNLXHnkIDAIxjCGXuQfLxC2na2pyWDz1dLGAHziARCFq
EOs3sjB+CsAA1zEZ7LOmau2JM+svEBVfXHt0TuyYfKpyQiebD4YE4NHylwuUxG5W
Ld2ExQ3P99J9beTWBQ8Q1hU51mkoQ7jftbo6XE9xoubVUisX3a54tO0LjZAkhMn3
EHAv/UWKCbChbVwiKo0mca/WHbi1tMU1RjJSenxvoTwAhIliEHr1+LRjnJvUeUf2
0mafJCai6sgYQqPZTMfR6Z8lcQqiiiyUPfjtaIfGk4Z7o/ZwNBdzCYatV3wMbGQN
/JcCX30xPxg1uzCFza+gMHKtaVXXc+dYaRo05s0A3CH/GkodTlQ8QeSreGgQDTqW
9PXspoi5Zljei6quDc3YQyZTYoccF6BW6SgUtcH0WPcDWM90ZFnNsJPbiFerXwT7
kgAga9rzsM+K8IPGU8+rdZe8ldl4jCgdcpTVAGnnD8Y5tPdZvMLRv3xZAb5AUyhm
Z9DuBRyT7ngJNwP3N8gXxZfdJWpryNgwnV9h8nnqXK8CGW1C7+NrNYxTNC8+ElSl
jlpzICvGcedMa6Tqg1f8zN3kKod2XaicajNI6t1dJuL30ucESOAieaBMEHVvniBZ
/4iW0HfGj0YPA/OAVlD38MyHsz3PA3Myc/pk+e8gHTt6gYbHPR4o2VCKwKxwgjPE
GgzLUnCHFvS6aDh57rka1Qitxe0dh90icSIwEHx8afxxsnRonhNH88QFEdBvks8/
wjYLHfV4quzxcmZPZAnxSz4C5xJVRjRhzWpD2rTTm+sClYW6JsQUMG9Tv52WuCw8
GkY0FoQkfFfDGN7BvhOqP7w6fdnOHQa4pbaw/BDO72vn6+U4AUxQZ/VB5Esn0VDT
/GxliLXJIBbIBmW2ImX4PaitlmfK8Wl0rb0Flk2lQ/mGk0Lg340xR2eM9kGXdF8W
Gt5Nj6PcKbplLT5h3ubEl6V0MFn3+U1Z2yKG2CqpF363rPsXfv36u+CXuuMa2SZ7
HYHoQWWwfWceDSTueTm3b8PB/gP+BZda/z21zBMV/tRVSlSIGT3lZW8sX5mc1mfu
s544E0H2tTT1FRoSp84xGA+TABEPB15JpCcIxx8E2SUdSk2HhntEQfOA4MK9ZBpB
Ni8m831eSER/fIPXoyC10t45YhWaN6529x9FxJcj6l5OaIiY5J7y1O6x9ZJ4whmz
dmMFZxtWuYnHsE5hCdC4MblLIw84pUkKzHebnVUP/400uU9M2rnuYNuHJV87inyj
iFPsrPiYi97XbDWsFWecgv6Y3x8tlSEh2b4YgROtpW1PNraQMh4JQ5jK4aDBTpPC
kJsvpwc++ZUf3uMOkzSTO3dJmP4XWHrcPEwWhgjdkD5aK+gfuE3qgjLcTQBQjvj3
A5yPeqoeDul0P5FLDQJl/KPBPHXq4d2Ysj4jRt10LtwVwnGd/5tbIrUYW/N/ZIxx
rw0vqsueQp74ySUCklsZVUqaPnaUqOd2aDLzuvLU0NoWV/eZcVNydVj3zZwL943y
Sn36kM5TcYmMwZDdnweMnMh0jllSVv6e4lYGSMFQBHij9nRY1dUi5ORpcpxZG/WM
G6X+BMwwJTTCyrVblPORgAN3T3mmJvZ/AG0ZN+MVfZwBXq3+F+TzNJMmaxmOAjmz
teZvKWAx3vNEe2M+QdaY9YbmL3112rpxa4ySMEegUhdKKGVG/z2RnospgV59/ch1
sjdTN9JRl8b+OBYz2hWZC0XZMp5p0YAe1ODy+9p//jt/DdbK9hwHA1pi1/VCXTWy
0wYKUOx+sHHsH8q4ZdrFMxeeEMXGMd3XS51mmh8j8PxpEHKqjoDRIioHCKilEm91
SosAf7KK1DtMD+CXpovvBwQKtGSZmmvRaCEylD6g1AfYAPa2Q0Y1gzzaV8L6Zb5n
3yeO7vOJs9PNnxr5wngTuHfZu+fhhzyM55mKY0xiCGtBpxHHMi7NDULjtVI2l0CO
KmPhP0F9jDKFIa2Tl6nLK4Mpc8YLkNuRgujomvXps0a3EweA7zeeqGgZFJU9rk5x
XG0fawOkAyFP/B+CzyrdS/v5AIq8KIz5+e9csR6ZvUC9C784RoTULMkF4+OEmG6P
hMnPNXWCW5q8fjh+s2LtCk368ioA0yrnA+5gSlJaF7OPel7ah3z2+vQxHEAWA1R6
l1RWxfFnP40XqnkhS0VAfD5RKJBNgtGhOpWGVkwcumvpbWbowX88x8SdGLKXrI0t
sT+LDy8l3wlZuiu2gyWPp4n8uDOqx8mTVQ0dtUAn4bI0EkIy0eohScpAfmXTgXjX
EgpeOuTkbRbIHtSxUgcxzj7eLZUGLZ6g+tle4ZD4IsDvCgB7/i+fwXUeBcmtGYzg
bXxPM3V2BcYIQWP1XzY2jnf/y8IbilV+8lsKjyFabVxiyNWj4HrIGWLY5JXs1SWt
3nqGGH2AGObzBeAM2qeVvszr0p3qdw4HxqsZVmqN0Ruhd7qP8BeefB/KoEJ4plUY
a6JCel1k3Y6ltDzTI/D6Zz4Rxb0nUIxQ6GQoW/IjqSZvMly5dOlhWW7k8dWYJnHi
3UD5zewRf2QyqJrEDa6HNWIVHw/7EXLZXK5hfjgWr8ouTmAp1Y2yOu5LqlJ4piDo
9ExEZjU7j3SsZiO62C+05UKgVoy27/P+CewfzaONgHEAFysgURuOzO4Xq8z6RPnS
uC1gasTBkrMQmxq0E0kEwNaHBaXMprZAoRwUOltpCEkERpdHttJE7nYPTkr4Nx52
z07YqCGM2YMWqHdVn0fXWfGs2mHP/9d8ZiD4w5HvGeKSAL00N6PkNTiWkypF6ogn
j0KNrOZJLvA1gOsD5A14KkGSwPbkDmc/x+ojY01IYUTrxGKqJQa3iezM+AVAKQK8
vE/qAzu2M7pfacfCh2z5vqeMlWuR1UGJJSmTuSf0FEpMWVjLbi3usEgOa5/QTyfP
E2Q3Ag26AC3VawZ/LtcyHTr5NwNlbCMHTd3zX1jQHxKqXU8FtCLj95wcAdCW01GM
Ak0OgDazF46i2pz6g0/eIkoUk9R/Q9Cb4G7dQj2NzSm3+971QQScDeRYdQ0VY76p
dzKPc7+w7tCbvAqDAfG/L7nrbbHyUn7hZeAYqe9BP4Ow60hZmS37QEs7FB1kPu5c
kxSOgJesRNwYBazjMoDkFioGjuFDC2TY1qoyo71K+L+AZ+FYNcRgpzvP692iiaaJ
drsX2Ks6VqiV1pEW/l5e3zqlcCCpwUIJHhqAjFjW2JB9fqmr4b0DuKWaKG5skYxx
5ZGLhz4G1R1S5g1O606FRUGxaHqchQHEz/0VFxE7OgAFFpBJMo4J3XOayAacY7u/
EMd9Khb7IOFeRxYq2HxuOZXaCR59Al7POPe3eYlFIgu+vi5/4SERhUA1PtPU7J6m
ap5Ps+AXzSAVIVDjDCifPo6TaKnQiusZ2DSsDJVbiv5Wn8aD1Tj75iG3L+HY0lZs
RXAKxRNOrmDv6G7VPj2TO/FCS5AOxwWk/B8y9FvMLGKo2aowPWVPWQE2JhwOJM3f
y06+c/KXMmLI56+BZOO/rH269ntTZDvzhmO8B87u10GkXyUUUDDv2KlZJsIM/afA
Bu/4Q3qqgoAlAaP0k5eb1CIgmTwmhSej95sHlkPxh+Fuf0nuUT35eHBGcnI1aOd/
G0HmFm4Jhr5GQfkgXXlc36unYPka2DkRrMZpE8sJ3KhaZQ1EgAYYds6qQiFG5myp
Hb1mZRsl/iSMM/0WkoDX1yvmkAlvoqKGOoRL5jjxELinv3RRMwXc8WzeB7KKYnFi
r6FMEq/Brwh5GvxqiemzPTHTPoDW8ETe4gO9x8pPomtRf3XZxVe7K32mqkSiZgYE
rlwWRAJORX6SUZTUfjn8icCxawUATCUBrjFdc2KF/SqVaxp2ZvPcubxygQwFiL5R
ejJs8oKU6lTQZH1O3E0FLHclS79vRgNHidT0uK/Bmtca1ksem83UBQpLmccOYLD8
lXICekye9Vi5GH7ypiObEMkKiTy/9eN7OXSbyFLtMZo0IE0epzQ1nHoHGs0qRyHS
ukKs4ghqaAg4Mwk7K4VodxPFFcVdX38MLG5p04TVLAm6BOwFIR6JM6SuInYwj2sm
rYJG4MJ5vdxl0kX67eIjDAGsNDA/wzSopfCZ+Qn1PAUceTtZuBllZarUVjtxKot5
+VpGXoLEZjSgNnlUBwUlnUzGhJOj459naZyOH3GcEbYVAKGJCafS/tsN5aXEJ8z+
t18qlb05MU7DbXdLeg/uGQjG8giXDQyZvhRcrFtuRJV8TDLYZRqqXWWJvrFKPXlh
tVJHtKMYjfXRMzNn594wh5UhXv2TADUIj8yeGOe+/dI3/pASLJlJbOGDeNj8XjsX
M1uAw8fDCNXY1UbfU0pZxeDovrN9jzJKsMyhcKFWdo5FG/FFzqUW/DRRNqfwxXtE
jhNKusJlntKorL7RlNWhC8AFgMn7RQlXrv7w0WhLTJbEYoD70UAS/9SEuJBhbjEW
QQf9QOpqCY7zDN85QeBy9fAUu5fWXNciRNdKYWfHzipWMWpTSjPnqZ1jK+nQN6Q7
SwlywuOOuEwTCY4rq0XzdMNfxArdABvw8j+WOFhJd9+hBnIbcllqr3yO8mRkShi5
iu6qNB1U/bt/3belOt3x/+6aKpR8A3SHasK79Y32GTIe9NYRLFOX7lNrFcv6L0jJ
2Qdu/FxUJ8AINnMZOK9xWBB0KBlUAO/hPTT2AP10kodUi7rTZrogvOJNIN1O+Khu
PWHGgWd6Z7+HkUcOU/ZzMaGEuOTFU4boRlx/25+n+ID8poxDSyXyqijzBUDS80yW
Dv1hOGBarH41dILX4La+ApdvhuUsKQe0Yi3K8j4q3Cfqsl9/C/P2ij18Bnzm4Ryx
CakqvxTzSXtqza6kwDODmRxf+8OiBn43zo2YmriFG9I5ZU6tzn6nnU6tPkpcqhJv
FJpehKN+z4x5BQmGjNR2VncoYmQqBPEkjCvQMuGV26KgbOX5T0esDysYL6Fflitt
s+qJyyslMCJHekvnXCw/+BTZLHErBwMV6VHHL4pQV5zpOgxtzTDfyJLWty9gEYkU
5dgVR7ugHqg+FWszZEh0gawy70aSxfce7ssGogTWz1azE/EGjlbfl8B1vn7gQQHT
n56EbLSGlolYoeEj+Eu6zaJGf2XKR9zne1SYKbVsVPtS9cd+Y7MkyE7gonkNq68R
tOIz6orUf6HiIsuraPckjPTZsezjnNub6vUl3c4ZY3MS/iQx8FAI5Y8CIDFDIv3o
oYAh1D3/jzATi21XAGnbhz37Uj9qODwbCcMdmZLL7KjnLMS6WF+pSJTRcKrH/Oe6
LFl5yqNcnlJomB4qbvoJDI0qYRHz7T6G99BmZdydcMszyvvZZtGEyW/63aXI8zBm
NbW4hTzjbLDjdTGOvqxfQnxJ+hNa56B5KNJ9HL3fX9mpUZWINV4iMDEWPCg2TAF5
eKewVhWPRt/BwPFRUAFCoTn3k9nP+8uzcyvIXpYV2itHanpE5yQ2MfILjTmcQl+W
o3AZuMqeu5XwSiWrIYdYZIE96Y0wdDrKbTa+kduo9x/+gDKlwCivAGJWcWMFdbG9
bYFITkiEgvS7tug5plyR0ULhfOaonnoa61CZmDE1UcGmyBffhbbweStVBHSFr9L6
D6HBSFF+IJnzdtYXBLbKnkTh3aJ4xTP4m7X95WJsd+Vfj1toz2J+sRKUKsrsN7LL
gO/Tuo3OlgRinckQDPBNWKI31+2VSl6Fr0iDKj+jdV5MHM00okTutYh2hs/cBDVu
BnWtmE394vNP8qn4wdLufqJVFqKkGnYBp8Kq9k5AsYK9pQvhU1AVc8bp9WCsdRMb
2U4XV8p6OBGqAwY5wImj59EYJg7EE/9K3SxVOn6gv9UmHdyXzXh5Ci0XwwJ+KPf+
cMy8RZsnm+CB0BdN1p/mLTjm+F0IIcygiL3kDcZ3OQ1ej1bgYwniTjg75HMG3lQb
uBZ3HUJ3oisCmeo8MRpHfTcd3RhJjfg64uQZ+ElLeFRrx6Q/yxO/tinZ/jVm9ecn
6AwMsHyNEuiGR30iWBbLPOFlQTxbgpruqSs0ZReXU9SWR590aXDiaRCZwBCDE2VD
Uemb5hmViASFHgI2o7+QzIvOh44lSlYSeNURqHr58HC6aIxKdZQUEZweeBkPkN/q
IdpoVjDyiSgLo1peA6t7RMOttAvTdAXfuTyJ3ohjoE3k3xf1qP6nRzGwlL4OXY3W
j3l6xUI6qp02pcjd62UcVqFu5hZ1KUUmG14c9wMKI5MjwDQMGpgdN1osXbmt1rwT
V+xBrma8cSFow9yKF0zCsw+PJW5iolS+aGj9VWf+E1P9QhP1vkoXvDR+k2usVVuY
id+lVgRxiX9icyh5MvQvLMudZPnDafBW7F3MclrolLjiA3FLZmXl3awKA9INleSe
Xkqi7CWT6EXge43hU760Iwxs43JKnbYqp1rYV4YspSvZHGAUIVDelxO6ydXUpN2a
ud9cLUUNaIwqF2ZeCxeO941IC5+H6l8aiL+oDONFHgR768bQ7GVdCr3BkwyzKJ7d
qC5Ni++VvpYEWw7l5idEiCuQMiau1aS6Z5FWuOXSWwOTe5mJPIrTwbk5fD9ri8bL
s6IvTdn/PsU5XRpv+JsuSV+X13PZfPhtPf4kTfW3DWbmyno/ofVs+uLbw7tyRMfE
koZ/GHQ9vNrvKUzkJf0pOkQ/hkaYIxLZlbAFT7CSCMR93IEete2MjVJeht7kT897
TEdbn0VxIJ9pTcM92d2jMlRjCzbKJ2JexBBnFaqSb03P6O0QPoQtdBsxxu5nStok
nEj9oOXIXYURdQ/rtw0pYoB135rvyeYIPrwVuPnHqn+ZaISKkeMgQpiBjzBqGz72
7YaXOXCK455C/47jqHA3377f+YjTGFULizro178D5FCpJQAjx2uehZWFYBTMI0O1
R/9wg1N/xTgVTdRZDkvf6CCpUzDY5XyK0dqjcgQLv8cL9Tzfoe69rWd2haznmzfA
2cE0wK2EAGlnDOFczxN38Ab2GK5Ny8Bj10ZFqIEHpZQyS9mfP88uSbkC0CBGoVRS
vZn+WVozILbVjG76YzVQ9PueoB4cFlb720Z7iJ3Hg73QEwpNBJpqFT7KRQ7rpzEp
1Pk5VANDq5hILzNayPQH6j49BzOWpL5bSPRawGaztX/rcECOqTmgd5OIEEOmKN7z
dNNaGj/A/heethpVLnXkiskhuuTk6cHnYHUVvb9wlHN86yl5ut9ycA/1zrNeZFgo
InZMYX275MxUYT+I5NsC4dhY5BcloprFbu5hoDH6Ws8bZUhd6efYlNW1moASMR8C
b0bZ3P7e62YEFjSv/kiGgn8xR8fTpXcl2/K2x8wP+LolT17RsQdekH62pMqxLU3l
TInYD3S/Wd66sqS6I6h/LTmqrdI2qztRHFsAV0KSMyMOwHNtIINMSI3Gsn/YbcXq
osOK5bAV8f1N7sa0fc1IbDc00Ei14ApHHCQaDMefkw/tGsfMoWXG/k6rbLeWNCey
Ri9DiVf+KCH9ZOKTADaXaSfvop8oc0rhw3wH4UFEyjdRq1qS7zr1Vnxhc5nU5CRW
LDjJstpTa72VSEGe/8RoAyPYlPr3CWBYR5l+MWhEBsiqhzbgh1PL2BUbxeZGsB/O
Vp6k3FFNOBdKRGzcmTVZlmO/S20MgzCkrTtsR93e5aDYDtoGtNvxWFp+kmus7hJ6
ffyvrTLwbSob29Z1ufG/I8wiyWFmwtcm8ANQEw54eOqx3rLBXPN/N/w0OyznpY2Y
1DVYHNX9LEkf7STqNpzRNvA2JIa4MrZ9sTc6NUntuK3qMLqB9PfXHrSltnHO84+5
egFpsSZgwkrDdr80kVYnQJ3sJ9+WYz2Mkui18RDBNOQPxPIFrjIiB+IP2XSKEXYB
0Kd1fivNqOItyJQlSeiCP8I/ccU0QInKrIo8gHIUEs95zPDhYSTaePmH3iiL7TBg
Q4ydy6Ug61es4JxLsbynek7TSl3MrCdvDJ7Iinf7VAiV9InbV7V8r501A0Kc7ZX2
pKvLpkF7uYX1uU/OFvgrrsTm8r6PUDTdTREVA/O/9qgG1+Q3Nj2MylzfO3wWm6WM
jhUtuE5F7sFpgm45x5guFhAsW/xE+ZqK9tVXEwr62RYsLRNB01j76Bgol+1DYChi
vVOphp7hglhIg7lCeex+41YkGZONAUvwmVta8ZL/3r0sbA5DSX4sSZRiWTSxFmeF
EW38/LOFffS94Y8lQM4Mxo9i8+eDB/SzJ0umsH6jCOR9n/eXuA1BL8KiPaWDGybl
zlO1dmUZkG8gT7kKzVKfPRtZdperq1YdWmkKKixiY8QdSGUkU2M0najnKY95dnyF
zZJDM86nJMcqUDSzBYo8Z8oWkKGThQNTnyb1b/uc7/MDITcUzMHjzbOCjj1q4vSb
ZevgE6RXYYCntdrzJVXoLOBeISLItSovlknsEspauGtoHSo5O//rj8QRv87wr1vy
KxesGlwJwObow5r44YZcHImQb8dqSlc3U0hWfBIHAnFh1hMzoec/j+DCpUxWbJ0x
jgqnGDIrQ+kRuiDn3+JRp1WtCgEyga0qNUBVbS9WEWqe4E3R12lX2ZlHZZusrIw8
8EUOMws1NLpgKCRc3+Yg82uRFrSgF+HDx3lGnF/DABPdJaC9aFs4oulRyyiOuqc9
R6v4yZYGNiOtiohxgY7xGWe76Pu7FLTzqk/Jp5sgAYym5EeMijID6ggO7myCg1tM
h8C3MeXfxQeetq8j4h3JAyK2jyUxuAAgIJ1JLouEirT/b606zT2olglvRyYBKY/J
zR0cSwnNRlFUkig0ow1PTXxGYOKVSvPa0YkA9BegN821WcB/zDIO6KNCkcG6aBkg
YezwCIXA8UMFcE3g2aQDZ6FZ1l+g8U2TCd0+q5KNbW+OHe8ohi2EuLAwoLyATTI1
WZDnrYcRgxMfstV7dJ7YD8k+9+7YdsgfBL+6a5hhmYW7I6c1zu3ZSzMpG6R/LraH
Mwi1GsZMQLT4suA2HeidUb8MJZStJgrE1kQRga4QrzO/d4aBTamrYSRjW+kebOd5
3lxXp/JmBLq1WbTp0DSvlhxdn5f4FuDVB/lOdhu7MQx0qzf7uOEE+LQQ8mEqZj8w
k4sWPlmpuwaO1xIcv545y/ZZ1UnfdsNcl4YUcmQmVV9ORzVbgdnjqz6IzCEOXUXH
jf8t/2u0/d2HIoJckavxYc5wUSfw6YCWxNzns1GWbMAMuXzGbft3LsNUGfPA44rQ
YWu1hFbEMB8wdwF/7HBYBerYQkC2oWxP/CWY4sYchKA/zIset0G3qQGszjJIA8TM
HmGbvWsSNgdG2s2CfIgBjA2of3XDisvlmrpYdscGmNwqkihs8LyfEpnamEIZqUXO
M5ptPqq8dmHEpr4u6fDfNsnoelx1FBu4yOLkkQoKnjO+m0oexeSsF2WViu2F3Xl7
agodpT++Y1VnuLUlTUJnvOKgfGdgCG9tnj0Ts2WKz6TGapsV5eb+ruSkcBLEyg0y
b7sHrlpf1l459YOVBN4GkEvqarVTqLgreQZ4BakgO1BVcPOUN7fSqm6b9U1gmgwz
+Bx8jUba7dbvakzfVOfM//8B1s9K5QES0f2aUABXwrOQWu7fhOQ8Cikjh7LJUzCE
YplbLeJ1xxJhcOfoWIkwqfPo1dw4cNFBcvnOclajOsBgwIu2p1ek9xXPSQZpHJtF
6HzJuYTfUL/NFRq8bPliKkGIkt6GmCfyO+46xpFNxPsePVnciEHq5j+6CyyL0FfR
tZ62FQonYw8QPb+3cEJ6i8KruW6YIHqkHU3OWJj/UoqdlfwbgaNS/Tkpkeh/6LZK
PZbAfGvul1adcw7PQX4o4cm/Wl7X770PWs4bSqZxZZdY+qW9mQU/Nc9D9wGa4aoz
GRZT6oKwiSrV4nZUuonJeHsXgNaQ8Y+9R3kmpd4uJn2gk35lHEPEHRfNyadAdway
MQEgLNhnjLKZszkq46tt1MhjQB6mUN/lYX6P+Vt/5kw4j2SfF9wxZB6wllmallv6
TEKNWD1Eu7G7hXFcjzEiRg3p2HtweAblTgm0lidd7cnuxcP5BoOG5Lp2Gc2AAGNX
CsYqo1eXZavdLZCPQdGWXX2mQLLElQQ6KqWenrtemk0eZ7vYJD6zILMjLaqZ+aw8
jDCMO8rUCnEv8X+UxPZb4apbd+BEl1lnaDbVDAVZ7rD3uo9IsNP1jta6ejZuP1AV
xE9RCzws6ToauFdimauOzHWkkuacwFGO3KPyIDXGkJsByboE/HeYt2XwrWdrTRuD
FHPFZnFwRuDI0kMU5kRM1N7Ne+dKfQi9v/ZdqVyqGG+cuPg6V2xEAleLn0tevPvN
z2IrHQG5JaY+FCCBISFESQ3tOl4PcKe2sjwbazh3m4s9Z+PCC9+0A1fQvWEIihQV
I43S7sGp4T0yFiWTUGuCBIwts047Xk2TzbZ2hqB4ilfeGlv+GzYavCXkZb4+gPAr
2lVNh9r0cffsDRzOGEv+M2oxWmJuCJ0CFujqeHIPB5xuU3/AhZaaB0CVD6/qtZ0D
ZvDm1rpnItHVItkGmAmfZMSMnEXp1oUlr+i7b3SGFmvURzb1Hq5MnQLZl7uewmRH
BJ+KLQvuv54HXdFVBLwClqffQ48sUsk3Ta1It2WJ3uTW8mtCQf4GhxJGvd6sm383
QtfB4foABEpecCxLQVRfDmWuh7VxAMM31xV4wARE7H5G4GTlzG2okX9auAFfIBb6
Vuer/L8VgM+CmCMREQud/Nnql0ZzlcbBfyTVyujcQPKAKzzXorQFikL3uM5gye2w
4/enqxnaZwSd04V7hKbMvSOsGNRLv3PtenxPSFvfxSpP6QuG+qdhxS34LoStaRFq
ma3mhEf7NOCszICgz+O7UrH7wexYIxt//ySeHp21ALjUjMdCRZKxPnf7+4iDKC50
6s9wQOKXZYuvEQa9j4wi6mTx8vtKviEcvk8JLmFEI/NC3gtBOfJQpCuBkK2479ZU
aL4IjR7Gxr9aOBim1sKp+DSIIacORoVKERpc5wWR94S6hLWYfzYIqSXL8G0h2kge
1CFdiZHza8zH1l7vjR6Sgh12fHi42ctaFqustuIXUl6fGO/qMY+DAqs0xJLdudcF
T9FDceSdiejGLuDzOLL9hNXIVJildUDvuYp7n4fXLReJbTSOPVycv3G064C+6yxF
ZAJxZmJgB7KOmSAAUUfjhBF5vL1WQ17M5tfVkvHcqmf1IRI7xCEN7CjDZj0UocRo
zYuWZtMfkhHZf760vi/wn5ueZkJmwMbaEUEbDoCelOYzxcE+Aj7UACEWCrVYDUP5
L5RpDafbGoOTWwzdakqqJzJRSMTtN6Y7vL5y+GyWx/0LjZLS/sUc+uKJITNRKATC
7L9d33bx2vr927t4KXs/pveTbMhsxPcFdijhyZjqEw9cFzHbmHaN9RISZPVppyVx
Zky4kf76A5ikeRhM+erJ/FhD4t/tEpLUoQHIjFEreDrv67Pyx0dBHTMjD45UzKYv
NXTOgpLTsYyEWacZj8akKia517ZtGmxNjk10499fAozFEDpo1JoorQO394HJIcP9
dJgMZLhkgBG9doDCaH+LbfBqzShfjnbrnVt1zhUaC0ENCegn++RDB5oBASYShw7k
+HjglDaFQkAskVRGaorywleOGFdk9FHwcAPJwSyQS5+yeb4LAFec5wxsfwKmKJFV
axDW47Mm/INKYn/TlrRDktWp56d+Vcn6T8iJh4Q1xsWhQ+0LYSNcvWz/CFCj7AHE
KR2efiIBNR2ai2k4Zyk2xcWqcBtDN4++J5oBfPpeV4Sg3MQoTmNiXt+HE8pnaVl5
G+IJqPbAbt5pBCU3KvY9LMiRz1qN48R1Shh12GptnrRpmazCbIiJHTLIAGgFEWZF
vMZf6zbnfNnN/ezrEITryjM3CS4oeGip7TfFDhtYlPl6KAF81qV9opgQphG8GI34
0GD4cCU6hqab47vZ+8OKNMbx78T9EH6BqdS3NS30TaVknzl32L/oi+eAQ9oxTg1+
h/tJ3y39e/zbqIaFvwEhBF0kOqkATYaiw9WvKVtndXVmEcPs9hUwGaRTq0lJ0l97
SkJsVYTN+LOHV/+VkHGVrb8tpRjCECwhgzHgwIsPqOj26DGPPspCoFIZs2KA9xGg
yxiKVuTSSO7gfFlHvh9KP0HKidKlQMYf9w2adrsWjZu1h3A/ywsb2y5noRxkavat
GuYYoJqbF9OSSyaH3RgOGm/iAXHVcg32JQ98XYnQoUDSUrCR2y1qxdrgAq9SEKkt
i58VpOKZk9q3+4fwsTpgA5Pv7fXe7dkckinU6934Zln3AfMXV//qB0t7Dv2iFqv8
zfUeuFibJoh00pc8l4H409bczalLWop1Af4AkQXmlmWilJK+9yXy9G1TAf2ffxyb
UeXYB8AxI6Nxid6QqH/IXlIafTPpqR+9TEzfsHd1dlfU5YLj0hpdIfUyPKVrhCuK
1g9BeON+227cwmooH4WZaW3041X8jfF05ANdAOZuQllBORpm7GIV+1qeJFVrZR+K
DrzZ1qoMSNz3tDNDhjSc4XXvT1K5MO2ELAocPWtnJ1ifisKXV12EjrWuQxEbPvbA
QPHkNqGcVUOUEWWFfy5BqfLPNdw4qEOaOI9P88oBb5j8I37VXWjwmDUfVk7N6t1y
vOrx+JSA3VtuBfhAOOioPDH2FtnF4FF7a5HBmodEscKXyMbBcdk09P1qMYgSUljy
Rj8hiLU7aqhplToqsA3uhCUeFhNtJz8iB5CUlAjPzBmz/Vk3ZOStMXCRn95w4W4f
LTAnxkPI1RGl0LooP8BtOn3/U/iUfF+/UM1mzvL+TvAvKyXpL3+MHTH/GWGnJCsa
Gg9Hz44FUcnWzz+KQIuJqa6Tygt8xiEUQj2DdzVzN6niVgu/xVCcAu3io34MMaWe
7SDiZ08kzzcJaaN9W3Fxca899b+AfUpYcuzx+vYSr3ShLaXoWRobq2YKKL0OiCoe
ud/BErGmLyOPevvKqwT7It2V6is3x7m2PjiYIc55E1ISDqAjAAkmMF1Zp6ZFVgx2
MeJEnY+lQE31OOwEWG8Q04obtuwp26ALND9mnkWPq/qo4KLTZLTb8N9TJ3xkMOdv
9l/WDvWpbIEaj8tkvdBto2GJtBjj/RpCcxn7yUMrAWuIpLX9Vr2QefuiUQceDSqp
xFSIA0+huzeLRcTHE4HyolHZl6lciM26gira5JFvOScHRboO7VtxOBFHZCllsf8s
cMnQZyUyZvTIth0HaorewLTuCnXCC1YO4CHTdD2JiL8nPTFQT1oLMjXlnSWt0hNz
TNMtPxIj6ttzF26/A6vsFesyOiiv7dzj4Wb5w9JzjC4qkv1OEN2S/Wgyfo7msfH8
o5yA+ePxwI6W84m/Kx8Y12dK6LXqSrvwUWDLV/PX672A8FtBw0OhauMkSSz/Fg/K
uhiEMf7GY5VqjhVAGP1Slwjf2xwq7Zj98DhdTX/0VyUyDzlsIb+UEXVNfo6dvQSJ
y8WdFnXjaAjqUUINShAhCaFE1+Q68CDKXktfcFd6LZ8VmVz2rNc3nPrZVeDmKyhc
U5QlQe77l8J6qo3yKAdz4Hj1oj7OiZ2Y9QvqItmhIZJpRqTScTAynjrgml0JkRnW
ENn14tqvlrPR9+eCf4tHtYPqv0FATQ8w7E+eTEWj3xWdZBpRaC0qJtaExWuNtop/
tFNSyMaM5V8FW6OAwUWcNQ2iyZ0Q4aGpxU+5uJbjeiH3deJu+fv/dszZHwJJqUuN
ThG+K7unD4WlftD7yTBvT4HX+XwC3iWR+5Yoh3fQKFcro3Ww1oB50tg5BA5lvrpw
KUWgYCpigFUp2UL6AiVqpyRc49Ri0Gj77thtMbH2Rys8cnKC0UOjVIrVc60kFttj
WR1413DPYeCvvmtAu9zVuD5oRac4M5XEHGlBNybDMwNVKOiW8MZK1GEefLpyqmvM
O1bokF9cbCiTVJGkssQdbfJ/z5nGN61YKtx3l4YbpvbAlPsbGTChvZ6bnV9V9z2A
BqUSOaj3rtrvwGLKT0zL7bAfrzQ+dT9aATBdP8O0dr1BrsTpg+r5ORSpJTngow1H
RpxzdriUgt71h4zVMe4CRqCo/gjf2BJUQ7mi+8a7K1lEKQqwBwshX2HByKPQUcEM
TWih1mJ40LqBn9sTCShhOzhQWl7koKgz3y0wTJlqz0P476gzHOrYlQicB8xqSaje
+gu56nYZTegj8Wd34uLzB7JQJKyKUph6jQHUKl4m7megqB+3rBfR0TziTJ/RptL5
P+vigiIOG6xD+r03cmZRg6dHsIjqqfiwsG0GIC1V7OyDVbxxHp5Nux8x0qJPu6yC
Jd72igvdGLfKIvKX3Y1recw1gPprY81YDVBa3NVnaRqYWL+oo/iphk3aufQQgvNz
UoZ39TUgHGSSmgwofkzFaOCMq5KnOO9ZtJ9BT0U+MpvLbiFWSk1lPYMTqmSDlvHj
Ui/97w3depDICsQamvLFubYBWjHpxODfBNxjaZpKY+0PWmFvaj3glN+1e6YKwljI
jx0IwUVZfNFq0F66agLBfm5+GU8rISHv3GmYoBlMHEhmWamWKhI2v4kMqBxMXHuU
IwloHbI00s61bNfoMZWHUvrEhOhIgg/QQEiC3N9vBAzsApa+5zCasZIugZ16KOwW
K7+lZunM1865InvYBAv2QcpfUQn3YpC7sG0oW/SzCIsR6Vyk8bwCHueB+R9MwYJO
t+6JulAQ1+jXF65yNnItgc3KdOD5ZzbL194d4JVmYU0aJtjpa5vSpEFtRQNkMi1K
I6ivaFbkH/j0BKFi66d9B1uWjDkoyYFUn9augd1HZnkjShcwE/K56OJNCy5oRuzg
/zzpAjFjujl1HAQgiarwGzRS23kobv83bSyz2H8wpKnmHrJBxN0b6NpHGSwu7f1a
JcpAHPqs3qLIn5ezxp3VABjyD1BbPH5EK1gKYhR6MYN66j5V8/fY7Efn3m5eww0L
+VVbe0jE0JuW2O2llLz677gtKQWe70l2XijYRjpOmZYJGg7gIg7JuQidZsQF+fhD
ovuBT2JjdzQG+tBVt6FLwLc7WmNTz5sK59x5DM0lHBqO9uUX2x3+UHYMW6CdX4LG
9Y2zsFdBOZryUprK0vD61gsh9hn82ASK5Qoi7OsZm+gQSsVbKYT6gbzl0skbVH2h
BFQ28BLBBdHu+z58tYXLNBEZ3tYUzK2wWYkLaTBvKQp5cH7oATXFvI8OgsY+AJRf
a7R5WqN5UtfYg2BhI0GLl2IWa0/uwoAZcBzdc5VSco95QfH9jGMuXc0OOWVgYdmA
QWpaEjY5a7spw43Mec5CKqAyQfdGmDKqyDX45fugpx7zkNkCWVJaLCp9XzZm8RcM
rZbBaJ9EoCLL9k4En3WrultQ5+2r491Mcb+z6suZ10gRk1VL3VobrjvTi+REPQR0
MQ5IcQnaEpZKuszyyknCGNmhQzFrqsro0K6QgB0bRYAvZHu2rQWz3Q4nplegv0HL
j1t5tkXJNOlvCKuKbFEyipvhYoVTtamocRf4Q+xs7f5JcWNpTtL4IG7tEBgb50sk
WfGHs+kU0W3OflGAnjXHLlsSKKLs83vULENWQUUI3B+Ix9rfynEaUSyCrQSKmBiG
rMi4cav1mOyWaiSLD7amOYnIc+uP8ez9ic5lpzFQxMQkR2rQjw2UlLl9wDehcV/t
0FAMKku6hd78+9BEaEKUrpi7DcYKCHNWnQZiCh8sqGS7vo2qHCTf/v2Ais8Y6MdB
JEpNaN0F/f4JrI7rCDTCRbD8PjH3vYfj8e9eO47xU8nxp30FN2uN0RvE/CQ+dxeB
4mYSSnyRL24qOLwlIwJO1KeqIzS50c6U3A9/GKdmiGBQpaRtF+dEjF0Sen9wU9w1
Cf2LJomTtErPrL89WTmBvQUZTpviCPBBthQz3RZwQ9rsALn9dIdfO/+uM2gRcf+0
DlwLO6YI3v8FuMzL5OyVH+QgjstQyDIMY+Ci7L5ZEm+juZjRIgOdSz65J5AtCwFy
l8am7gdkxjbrh5BE8aa9GWcuL8ZXO51bRdLxUPRdyXbJhxZRPqCiW1onouKcuAcb
qYnNBH0If+IaflYHc7Gr1MAF6EZzPk7U94ljV7alR/R4iYBmPS7PaWcwxVjVL1eR
w0E7ZPV6eWnEEp2xb//9G1FwmucIydLjc/TERicx/F17XF7FMv0+MbvakOPbxfNg
BScQzxNKles3UYRk8DrKTWAGd5JO3PWRtCDVWqdOYwhT8Oaw9q9xo0yxG2rUT1nM
blnCCKBiMV/Zt1SONmnLj6bNU99WDhbIjG+DCoyGVQi7ABFZuNiC9SkBu32BiHjX
NHqdygWHGEotLvvBNy2IrTVGcYYC9XjYgxd4MpS8ikzajhtIzqKOZU9vfrb3KCmE
SlzSWqtuvT91YBxnlsIpVOskPOSmw+WeHRJxe/AG6+tAnvmOqy1YvkiT9n2yYgB9
/ClPSzCzh4tTFbdtPg7VS/J6ANu19k1jK5ztFejp9MLCXrbq+w4Eg/WZcf53mWTG
Mt0l02Yg2IxJQqqfKLIy0x8Tv410T7SKudjFr8oAFii9n5kzXJvLCakYUSZjIhoI
CvYINjt5EYDcaPY3dhpbpXF3DfQFZZBXowkHp1bDQUH+UQW+rVBqJmWCRhra1Pzm
yIU6Bgj+QX4SojlngBtu5fe0dIccunrxskTVaz1atEhi9Ec51Y0G7NSObyS3BAgN
4q8YHcJGe1k7axVVykMPqLKBK+ZVOuKQFoGa5tdeJNb7PBNa3lH+i0ImSlX9NH7m
YF2xbEQeD3utEf/6vznh/f7A8oyZoa75eDnbFG5vrWjiaT6z/9G8UHO/9biQ96nK
xjqmdskMcQSSj4FSROeGmvGD91BpAueQR0e8Y9+RrlzmoQ+ua9rY0omEgTSMeTUl
w9sGt7c+DdLR4cP0NbRRZQxJ4n5uzfwKLz+AifK/J4zb/1Jn5ifqNeoksIsHEIci
6rJ71TPeBVGlPVVhGkzjydtbWb1vzxWBKbY2rbV4GmN1A04oc6w0w6Q1nZM0Tu4z
40aYgP26/Z/cVefgQprgRwY5KBLkPq5Q5iprQHzu0Dh3Cj8D124mNgyIWXT5gpiZ
WFjezSViRw64f1dzmYAatU3S9lQTCvoMmE4nAMd1Yps3i0XZ7YCw13Bcw3ka61NY
E9RPaGotuObtA5l6s65LQQkLf3M5+wZRebF606cleg5aYYt8g93OTXhnzahSfQ2A
Ro0XtzAX7+weWHsaYbhPXBWYrxvZJZcESwD3iy4OUlkJZyHadqoQmrnioSzyvuXZ
5BuM7hozUAlPv3VKg4IcaBKXeVRVFw54uqHu0tdxOIkRlcXu8yXbb8IDj8RDFkwP
8efygVBbS8l/sfmTDnV1/fnx+pNf9Z7aZ8x1zw7orX426z2fRRyHYEdjl0WSXnOW
EDm49ZN3iC4+N4Sql6Wlhl+XK9UJeVEz24piz09Bg6R81dbehXho78hKdVEqBhdh
dZkd/LQUeWxF+fqpKhe9bRfmE0X5m+/BJTGDEyOAe0LhMobX6iP2YBhbfjMVs5bC
xx5RHd/0Dh/Vr9/W4U1pEzUxSby3nAaG3um93CIRCj0EXofvVtOirPjB6wU5sBvq
DblC8NJqFKpIOng2T3UPgQMMjZ+l46vlnLmD1kYViPESVXHMYaMp+jnjOq8l6QgX
LY40HCnLXHvIKf04Y1Jles5w1k2lPppfsDyXewWWfBCFSGlkM8LjNBAsdHKQp/g2
HevrKv3gL5e3Wk0v2bJOGaVjG59IdGJI6kRwOfNEV0ktPdigg0LnrviJdMJHNTCp
HHQ+XYKcfC56Y2nqAeqjJd0K9RpkrVn4FENQfDxKeCgwQGxz45gr6RnWaBVOPXlb
+1A6ET4rP65vKnUBbkNRn3ndBfZi+038h2dtrmIrb4JTLel4SVeJ+uYKL2mazv6e
V00iNWjX24leT4VTnkPdFFNyArV/d+712eY2h+kM4kbiiUeEuha7rWu2WUU2/75I
d8ALlU5hNxbNBLd1qVo+FurgV057vTWcf0WIEJWcaa1k+cMVJklqzLgXeNJmf6hV
yqRHzs928KhsnBcmJzRCdQYhfaQOZgBqxmNX7RVt3yp5aSJ+0jjkGkOCQ1vq95fA
I7Kga8HaQ9qHJSrIgVibxPLOd0BdtLhH+w97F64OUlRJ7bd8H2+m/GZDUHoDwflT
EkAK89SqXvIgGJx1hckbK5eackhIR7XvxLm2Dctr6QaiElYvO9MJHRG8vZgBqvYS
N+1CIbilc5Esh5xwEjr4WWILCvQo9tX8MPd7/b2Z4MfUya4LK1JmlU8Tv4dNMWTC
/rkFrGDHA0p9gtjjBywmv74YnukwpvL8vu4+mKMlNO0Kx/bNIXOvv+C4OeQDl0EH
mgOjB8+aDvSSoDHvkqadg4v67fkg7hHB918TiCg5ifP28toiM4kzB5zg50fEY3sz
OjHoh1vWsHBUnWZ44wgluxRSHSSqjFrv6IZzvkN9+h98c//SP2am9e59+hjIBr30
62+lEfdJwOWltNPwGnC+6QNZb/p6fr+152lQX6w++3U7BlI4N/LLo4hi69yBh1MY
/AWVQT0ziwqalGpqck1/pFKUYx0IuTD+JyzatX6yDXb/ohAK+Mv5p1ruNoHfl0sX
NpQTZqfQl2xg+cALrdaAmDayyQziNtuAsH+D1LBQQtcokkaEsiHbcV/YBN6lsAVA
ffsxf76AMSi2HDqMuHAKmWfMNMIBtdPS75zKrljUY+DVNm0j+dYg3vKwVZN8q+80
veolhCAwidW4yJ+eEtPXZyPY+/nqCKQV8SFrQAhASbZ+lrqAY+pXwLDUy3+CkpUi
nkMunNPtf+P74wT7xL2j9vg0PEDukRHYbe6de7B4oguDByazuAm0qtZVEubTZiim
znqAk7SNoDIFj8NNhdACdG029WML8rTHb2QMcHWBinhCP8c/v2kGH4OGPppyQdL4
zURWcq8eWwlJzx0rAA3HAKRLiM9Reto4NWg9OIfUEuKcVLUxqc6TSrwfRnArEPqr
DUjowd6nzxXFhAoMdcFu5I+5ucDno7Zqf6V81sA9GI1jK3lofS39KazeFzwynxnP
XaM3D1oNzTp1eP3UF6rlKuHzdXqU8APOfYmP1S9z87FCzD7DBRMk6OfNOgQk0bN5
/7QfCfvBG6XC3qS2TTXhnMjpdnuha0X2wkhVngnOfIhxJwqGlChIigCYNGzwCYHy
F6DKUorsl3PH5qcPAKKl+HWfH/ntS1AxZR8cJQoviNL1yevi0W34U9NoOY4nInX9
j0qfr/yKykeI4hy0/868yXfHchdIt6o9nXBL0O9/nNvcn9EvaS90YycLoq8LQMWa
uajcNIrnPvwO+eXfCxuZ/RAZAPVeFuXLkeP4iXsE35H0LU41AMM+8ckzi4XJc8HZ
nyfY/5TprCIGE1vNegecyHRtIpHD+76EZkGyXhORLy8DnTssmzgUg+RXQNE1NhcF
e5XrWQz3G5BfupOz+4pOGn13siCsD34kiynVjbcLYiK4qNcHCGr6oHFUK3tGX8hU
no0RW/+Toakf3ZAHQMzywoekX++MEqIxy1GuI0c+QZO8RPlcpnq3uH/Xl6pKbM35
3w9vM+KyW45GGraDti+NnUqNx2Aj+LvXqEfEo30Rxsonr/nOlgLT9pDqmtmqK2y0
Ln7qHtgmpn5ROSd1DP/r/eoV0OfLAV5fw16dI5riAS8owMDq2IBxqJsr/VQiGcqS
gQCgTnxF7wRqk853bZg1X6ShNE77j9A3xogeYpZpbjk1KB08aF9LwTNFod0wWqaI
AdfQh4256bdaJCl4kD7RZ60qmP8xiB3ndqxk8xeGQRPKx1ioZ9wpbNwmvFNRJ/Uk
SA9HTXQU5xFauO4XVbn8P+4lNCgfK/Ln0ullQTzqfNOjFsAJBRknoQUK2zUODcfC
TGOZ7fnMlVR7CQ+11e4ODQLIbQ29aeSLEzxZOwjA6tJayK2QGyf3EmHR8L39Ysql
Tupb6P2zEv2mWAzc2879W8fWLTgFcJnY45EEm1kKT1332MOVo4esbnMS0wR4ShGV
ucv8X4Svw7uDYBkvBORawuHXPvBbYHRLEOEZMUFxu0NP3gYeHh311TAWNQf6LXB2
GMVVRZ/kQf1BSPSJwp6wzjO+ytd1EUCguIC112ccTZEOii9FZH2Ead1kUTLGXmQp
U82NqXfutJGMdYs9QJTASttRkUE67ZwO3iD6XNrfDySUBzcyzNyWJ8wc0A7hzuLE
rT7bttbp9h+mEoVcNfQoOSEUJRJR+ajqhCq45IU6Mr/tOXDsbehJa1MvLccu2/wC
xtyYgGbGz42pKju4AMROz3xRx+cITh/uvi+MZuYjtnPVVF3pV35rMh6DqxRCXOw5
X8UEFtD94rW8T4eT8meZKw3EhHZcCmXydb4CUnHRjbAzfGv6TTH86LsVQuB8Ccqj
WU2G7XcC8dAoZ/s1UKsJP7jsdsOhZD0R+choGUktFkN1GcdbcdhcrvuJ8qUuRbJA
clyOvy/5SwfnFvW+OBUyBzqI5I0buDNIsUe/APA4NMWO34weZVUeQ+CIukE5wcIk
NDwk1Csmr7ejYNBQtqUwLOZ+GYI3zItoLXy1bni56IlUcGwl8YvZu7Cd3siaZegu
DvJxmpKwUqs2GuLxT27d/XovPSgtq0XI29uGCbh7bvK1TRqaVNU+GzrxnLUH0HEX
Sx62sydNHIIT1q6T4XF4VbD5rj5eHq2Uwe0x3mFcwXyiJpe9Md/Gnw93FWlXR4zh
YTgGyCgUBSvJORfn9PrNXNTP3x/2zc3JbzRmmf48qoFSRs0fvwC++g7iN9KmQ7pu
qg9PhnJYidQuTKCldoMMZayVCo7FmXEhWF38LAmTYAgtd4tImqvt6XMoO06DJIw/
/T3XQoJ2dh/7B+k0KSbRHt8oHaCgbuvrh4AQ/nZt1rBcDEGdr2/NAEOv6wNG/Scb
tkdUbWwQf5Sk1C83Gx2dEQV8OAz9PVjuebhtdTJJH4cGstIYP8CNV2SThjpjXoi0
ubiiTvnqSsv5u3FUSfvIFtLBAO7T343bwwVIlnRxbscKo0LIe2ANMbiak3O+7gPg
Y7IVAZWcFi9wQ+Cbllew24JKfx4XEgPNAaGCuMtcgB0Pfx7fkORiI81PDaqm0jAU
xGwKoLonpMbYAf/MLMSCsGJF08HmeiMnwKZp1lhJIqprEwKd0YeoWJC6hGOZ3cH6
3MCfqVA5Zn+G8d4tXKNkZHIXkf1WhdZhBCBVmHT2O7Lpj7ZKJJZo9rGp81Cvs3xi
77uwLbeZQpVHoSbP7XbJ9U+9F54fm58H5Z0tyoyDV66khrB4x6M1kQXCn+mzNPjT
bRDB4mUdLBYM3erdU3BEBjUajOEAIjy4VoUiXhKQEvRkQm4ejCG9nN6HAAwx+j8l
aVgp0VDFAWLpVkmwHdWyDQnsvR8ZPL1FglxiRYF1rdfR95PgqKAKyOmqDyO4Admt
Dp0PXjmXELYxGdi4eG57x2qCQKGwZAImRefXUro1Vdrq4lvLO5CoACOCQz/V+RrE
+4nuyuFqqiw5j14SQ1syo4uYWNYZZ4Bmne21O1IYla2jK7PHc79hsAXqhAn/0ONx
KQlkQiOrEumr8MR0Gw+Hxf1QW8guqM7LuDE0pKoAU91zLACuWTamoTHr76TSgjO3
KkVhug7VL1CU2kelXCMFiJ/Nl/Qu84t7FW89N3O2OucESkuSAo8bUQ0AXuXliQNz
pJ/YqdDNsQxDJK/ngDz/rxRAwA0Y0JWFC4E6DAqhgOgQnZbF48oQ2YW/ThsDbhaQ
mMXA2J7Zjy9R3iGH53Cs97IsZbpF5XujFJoljKUmZpK+eEuR0CKz0FkkLk7a1E2Z
kYAnwK1gOpkYHE4lCvtTPLOa0ZBSXmf5wGXYKTfvSh1qiR+7yBRw1kFsKy4fKKrT
UVAscl0bmKaqbdjs7rPP3AxWnN0gzR2184+b/ROSbysjltcGiRzvJB/tzAEl0uin
pa6UqVNcQ5R/7zjRGJKQ7EXeILE2yoESUG2njfVFsCm1C6wjeLB3pwyITmFBQNFe
RNXckOd5ctSic/y7jAtsj9SLZ7yl+wdYXorucmsB5mKjs1h2SiF9Q5YYpTtNAbVe
iq8+lNkCrcUvf/T0PosgWR4/+ufBPwExDfAmbRiVzmbg6hpbbTKgELgvHNVhCPsw
h4ajTMaOO4sK7wMF5y9av1v1HXrOXVC4+/laON8HfCMV5TRNd4C5YxIQeRyZhh7H
KzFBLBMZz3MKQLFZgEDNAWz5YEHR32jvnpswc+ZYnGh8Rq5ajn25+3zIiB/AnoOW
2mnp4Ssr+cZaBLQSvBvP8Hdi+FkPNhr4WozoFhQpfnN4w4mndc3r9YQl7vfmhsfu
Qs8yv0BlEPBQp/rtFAmX6l538L823PHk8PX7qNfQEeZKti5KO6xQ6nzq+TNMoXkz
iyGtlC2kpC+uwQqYfdVDcnvrALb/rKEEiLDnqWhRBS/7yMlaApdXF/MRfd6iMFSt
xCictWQABNMFYnjqFCHMzR2HjWoUaXkwQFSd3XKgE/iNIHLNuGxanL7DaXlxGrsz
LrVzDXs7JVtPdYE1prX62ykikkl6FTSsBUEj2ZGTDfspcPag1GTkKKM/WnGP2O/W
m1CquqCjzkSKAvjChEWgJgLulmP4EzRGstqToDPl/dXFzDVh17D/Mnb+D+6umj0T
lfRsSovq8pK1gXBkS914dVpQckLsejptn73Sg9ZW3GUtREM7c7+YdF2pfpZiRiyu
/GwyyCmbAg3LvFHE3FKi7rgQ15+iG2vcZLcsVDg7peLTvi/1wxh6gyxiDdT4CmQr
DXGSnitIFhy6obk+6FBWAHco4nXtroBvg5XSqR+rCqkK+WufuYaTFuheHzda95Od
smtFxJ/mgMRwl+4FetjW50gJppIJ8n0qxOQV1kgyE5v3OVPS1CkdK1Dc8bqxQtLX
ydJ5j3Jh4a/AhcOJaKVdCPPYD4Cuezmk7bX3VFRc6OGAf+PFno3sYwSCBxb9eZo9
eatGAwyliywOwSeCB3zvUQ8j3c6p4KroeuZ0j4TQXOhouocNhw8AkbDCqhSCai9u
Or8NJ1ho8NET767cvZ2VPW2Q72wHNZeIsvVLAlrqV8QnzYHxjy68oxaTTPPlYYxg
FjRVXDtAE/QKkoBGy4l8wMAZWJk00qCoPi/ITqJTPOmfTec5S7HUrRsgim7Xo0vi
Jj3lJR9CbXpPvOqTP3XIhwpLWobZ6Gwxi2dB3IwjTqk3sPUFkdnK2usEKtI41vuv
yDkiqWZrsgkdpJs4H7cz9l+chYkw251CI0XI+JUJ38/Erw7yPIQCDVAB1OGxaK4H
7QeXAmuSIBYOK89wrCzZqrJzqdzndwdnNwwIDezHEuEZOtcLZseWs3i1ivEIxCL0
k6T5CbY+7fwzNFM91S9mhDlHVMvojdi1b8O3OJohgJFRtcuCVzUaQ4/riDrIb/Hg
Pj2F8btrDe7fAHyH8W7AfzOQz64lLN8qefXkXOzLnM7a11X7vOdGEw/9htpVZGgA
PV7ccez3+LehInEii3T/Jb6Ogh4wJh0Y6RYx3ilGW8IPKmglgtj9LcEXXiQ1z7dn
9jeSnPhS7XK9HjCjij6q01p3XyUOUlqBsUPMikS4+UDM5vdkqjGn7tK4YEfDMzn7
Keb1gYzIEXDbCazrkeexAg6k6hjBfurb3bZ32+816lSrAvm9eQNIYuUAWAwzb559
ZTJi74gjHvUVgut8US1YAlZpmEIEI6kNk/a6ORYIYO0xCo8+K9Rt2XXkeZ4qymQi
kPBqkzFI5b2LENfgwVGqMhSMcAK3Fdzl0oV9m+mvY53+Zn73WSkh+tEcQi7wPZqb
2oVPoEf8bU0LVaRv41eOPFLgvTGjVC9Ukdpsr7JNx1PK0yk4TD+w5CL7ZVeK3Xba
XhQcMuS4ghnynHv4gf0gLqCP6B3JcZVQaYdnvoTD3dlGBhIoWRL7w+0Bf+TDFsy1
DvZDZ2OC8u/uFu4nrqHUFoP046xTSF/A1vWz0S2XHTvDF3h3ULa8TfqIOzqQWzZP
PgQCTZDlA6KQZj6ezLm7a5F7wkyaipm02NETlBwmyUCkpDSJBg+UJqOqzgHtBCd6
YWuHrYRbmyydtEdlV2pZVxqfnwXXNw0T3KIpSu2x9JQ/rLOrMpUfXs4g057YaxdU
8G9rT0fEI1qkA9YZwK90RyHGUGe5IdmIHfsN3ns7h3PT1pRnS1xmLGzEnawFd5zS
4TVIljgVuMllwQ1zUXzy44JuCobE4q/N1MhShSuQGHb3vfnAv78u2ePMARPQfbt4
hykZFL+DSBdWM9GTedeI8PXaVQnOEc8EOqaIKlcwQihBk1sL0TUv8c9AblgLz2PP
pLi8AC1YtJvjcDHrz4ITRWTv4Z4ukBZC9IXdpxA1SNhbGRqIYsFuOHdSED+jO4GP
6ioPByjh88DGsGTmzRdJpEbt7FZLL10tYJK7IXcAaBxjjnbbwKjNPXrqQ7BlsNyQ
EE1r0sFrAGquYka+RZBVaC3js5uvUgqGSfy5awk8FKOQRGWXZC4vtk2laz9pE42A
hTHQN1WP88uczHLoL3Yr9Jhpcw2zS0fwvFQeSVnL+dx0uEJxv83uQeSfhhWZ0CBX
0Nl3GdvBaZhT4l2QIvFFd54ZaeWiHPiwCA5R/bjUykojN87wcbKvZlT7pq3N0dEt
gjjSDn2EmRQb3LL9nnTCzNFCwIRH5d56HDlsxpVywSmLIBAz3TUBG3i2JAG6VpIb
uL3ErzFWVPxFelyKD8iu3TrH0PXPv0tCnDo6MnQf8Ydn+J4HFmzdTa6Hb5QUS46D
hNFTO2UqTDhBj3hM8Dc1heb5zvskWmUfikYTyN5T/UghAqHOmk4HGD0sdfmjmC2H
nbc8fYXLIAi0NqSv6jbpLfXpxWLY9+niBtl2OMXKcLMQ4K94CHLY6/7AI7eWcpuZ
tckibHRLaFkJVjOon6qo05KmhmfeN+btYL+B4IhduJnf5WQ+vDuu6O/xrDxJL0gO
H+5drpckqJkfQGHSlogAauZP0oGyRuuUohyM0QFOIK8UHuSOhVg4zem2IlIgg67G
4qFLQKJQzRvuQZHFsAlq2enlkgJZ/Qfe4njq24V4Ab+5Km8q+zxl33gzv1Y9289T
z6oj2gd8gQU47EypU0fNQRgMx5z0KjvmthRvWegeWZODWK2cmzZrcqCxMa+Hg94j
wtgoxfN1QHW9xUz6/30rp9xswXePG7a0un/Q60HHimZdmYQmuE3YEgoZAL/LABQD
eByuP0t1vnXzPz/vBqj+DZU8KKbcmFAPueiaWrOUS/iUrnjA0ZqUd6mz8V/4W+x0
DQGy73WTDHJqq88WtUnaDOTleUW59XsZPGswyRqBpm8QVvOQOhz2YmykulOUz+6O
B5CAVbbQuS0mM8D4Gq+EBWpH7T6VYcITlFLslmWDGZh2wW2rkG5kEgAitan6CGUZ
EXqKGFBWLH/BHf/y1hM3LakUid8dz4WnmOOEWm2v66PUKEyDnXXIMxQaveSHNYvZ
AoAq5bed/ueb1BbCpwQzSOryBWJZXdOaS/QUI0pZsSetyZfKuvgYZ9p6bEtELzZM
p7i6Exc2Q4EdUEJGRgCF8TGSy/9PEGxiXHys9gI2cTB29o1bE3fPar4DTq6n20eI
Q+W65TfUuekmuyLfBzUb4W7f5F1n2yZFwQSLJ49cwDpD1/d/hT+mNWriGEwMMttI
YK8QeO0R43sI7LAzrB7QCSmoVrlTyef8hqDMzffy7oSwnDAJQu1AWVhpK5jFPes3
jO4rJ3cscBXnxrSsk86VSod5ZzB0CcrRM7ALkq8fYiOjndOVVLnX6bi5FerFOUtt
uO5rClzNQBZQjYInpQeO/g9LzqwzeUURiqvoARGFUgMeDY+9lNMivlyEyBAQ0KNf
JjOayQqMFx3onoQV3luajTZ+kMo0N4IyR3P8kVpceiCr8JKsweEnQAg8vsFsMrKP
MwHzf1gNIKLXLJHDiyG66Iu8Y8CmOh5vnAy0oYgHNGNKv6VhuUdnS/5z0UEErFPJ
oR8+UAkkLZ3UX0gKdLsEp1aNwKRDAiIovEsJaSkwyfdVrA9w92C+UggmcSJ6Kl4g
LmnuW7OjP3Ea9EXV/tay4wP/DZpBkjgBzYB3SJFitcIISfJxT8smfazc+j2shmUj
KckdvAns4WiYB5Ch2NRS3Grav1nSpAT88EAy9FIMo0LNglaP9NS7OtUJIeEGlh64
4WcxvTq0IpTCsoeq2FiJe3ckg56dlF7F4/GiHmmG7HEL9UzIp4go/54c9jGh3T9X
z5FfQ/gjafEq0Hf/NIoBVlCS/oc0PQXmE4T2HCfZsKYL79oR56h/H3x6khvK6wEn
RVsFmyeNO/MRHRIfRuEbrcazwBeuAak1pMUiEjKP0gXoBz+8ML62Qcp90D83c99T
jo1yx2rJNFKR6HCAsjTWYhaAQQmMwlsHGT/3Wf88yNmyBisaF5LhzvHwiKEyXwMZ
zUVb5j7qiqK8syMzo/AIT11q/bVPU6s8/vp0LUIokKBN/WC53BxttkmZt+no4SpL
e/fEACOMv9WGtpZEUATSeqRZR4h8yz8uSuSmXn7DdZmJCZRfGHeit35ynh1TfvWI
I6l7S5maARVCVgnofQfjXLSSk+1BdafkDdrMeOuy3qrgQb02qiNoGDs+mfIEwjRN
kF64pCUtVwnaxDuD3kVbaqNr4kb03AJN89RI5POZyufv7BnsDTAzDAmXt9ieo7gQ
JoRTRXuVAwMKh/JqHmGkOF864VKK08TmmNPwyi6NI0Roq7vZ9UQvl6uamLLVO/kn
V/mIfDDV2bQCIHyZkglS1U9vimSchAegmWjQl19vZW012Sixf3Uhq11vafnBbqkh
NEjVW7dec0Y27CdRzyuRhZLeiL+8v9FdP72klXUOUXt8D1cs5MRdlvwW+ybivhEJ
0559FQU8NoO7zlqukFEfrFyHjEoPIqd0mVnnboJ7aWFMjmZETsD78J23d/kWX3i4
nlLmfOuzGWNSFIfj+6OdeYZ+DtxVP5RYUlpAwvhnQIBy+x8fn10/ekT/QIgglMCl
CkuW1OqQMj3GONr9mahjKAaPzTR/OHj648ax9Lk1Uf3Jk8ZzE+gDFrzWtpn1krT+
VCt0MhmIA9puTSHfcvj2a7J1Tirl8XB6a7JILvSnK79++RGlPmSQAdIGNtUosQWZ
6WqrtnM1ySzht1MlNGb96TdPSKkiVPvZTpwvJyJABprhcyUqNh46eQ0f/vYIgTvM
fW3V5pN27XgtvLUemR1kKU5alMsTWMKI9DF7lNwG/W4kFGNXsJVWYKcfwGcbwQh/
FSVqqENs+vYBVJc29HJMvp97/W3OWJJLvsDQbLQML22JicymK+ov8WtDPp7/7xSV
hg9m3I6WFcBVPuJ2MrIYV9UCOxph3554dsGftekwb5OY/lBU5cnb3WqYm7RX9Fgn
KmdIbX2XDXqs22LVnST4ZcYq/CpphHiYSxZViTboCldIE0Fi037M9Rm/32tCtm0D
adnSbHPdW0bw9AkLaBokf3ApxwktnSIQa7sYJ1+4yjLwLb8s+yam3NpoGbpsYKRu
cQbLVmWq4kzfmXn0m2Psuo9tHHMjaZ83HBKs4BAKs39TZoLKaywNeqpk22VihpqR
K3jy2CRDtDL4vaVOl8xrwYKXlm4TpmMicDoktDyJvrXJURIvwpZD5XCbJ2dn8a3D
FvyrqcvmSBLaxGzlAJ/hoiBygTzDnY6ZNISQzVpCweo+T87Z5gsZQA86SVSWq9S8
Fsmbw2LMUK1Ki7be6Xzdsj5Kvf6Xy6083Lg1GQvw2HzQiO59brXF/tr6/eFHZJcW
S5QzGFpbxg3qCxt9ELHOvmcTv1fQi4y8+YhFVA0hn/whyM+l6wZw1fF8GqURS2q3
FfVTaTLTTC6w5APYV4QLEJ2uW8MrcY+ye45IhlEXqcbVQTcQr2ZaVBdNTSYSQS4e
V7JVdalddkQ0N8qQ2mA+9fR1+E4okXWUgxZvecjFE9LDVSkf/dOAFGQ20WloxuAC
CcoPv6kdSsEPZjVa9w/PJtcEjwwWulVpz2/SI3h9nB4jcg1R6nAzdvRs8T9yYClM
vSkFekOg2aVbPl71w2EymMVaG58XO7n3QC89tHVExgUPQU7aGf195zHNyI1Nlkhe
PsD7PlPirxE2fBEs1Et1+L202AjY2T2QJ/Cwks9Gmi2D/pM9y+l8lWfpJqijmOeR
l3iRK2ywDkZ5Mx7VS5qo8BIo5q1DAFJkor1qjMTEb6DSFZjaG1xM4P4dXpnRCWSI
xJvOY9AWRoPhIXrrc5s/BnoHrf0gGH65mAOGtfQTNQeOgG4ZNMffwIY+KB0RrCdQ
lashiJLc3flp5qENrksO4mLzWeBS3GwjY1oKj+HjS4EZoBBKqxQKZ2f9w59hh16j
r6Zc3qqnmKgRAiqgQ3KalcCZQ/W3PzVUQbjtpdjV/MipgtKQui1+F7hy/EoyJ3x4
b0YaVc7aM6qYnGcmV2nTmBYdYPrPZynvROhToaeNU6ZKPvTPBrQ/aiNioSS5/6pZ
YICVkv4Q7qN2rkJPX+9qOHTPdpUAdHQaxXFu8iWyVfZZxhCmbNGkFhlHiVustR+H
+vTVAPJpyfgWTG1R80jzrn/kpaKp69aM7119bZn0WjSaZwGQDf5X1c01l4/ZxhpC
62mov7HQowl0xf9YXP+EaGFxmMixOR55WwOX2gkQZDvUH9nfrLFxEGR3fWtYjmM3
gHGnLVyPhuGV7OVq1BhiA7xjgLE+77Xw6qxe4W0OAjkGZgAJC5ckdvKPxxpN+oE5
dPIY5iK0xAOzgh0m5kfFkyPDEpcoo9tWiw0MiYeZb6XKIttGShx2iDbhDQi760yN
ZOGCBS3GHe43wd3aEcPHv5zfFo3j347CbuncSy5Wc49T1/67ktSG4Ms4rW5WD+vc
7N0AXJqifRK3MkQ3Fz4387zmJ3ForGk5HdtiR9q5YRwMhxz4dRHtdMkf+OJVsCH6
4AFjN8bEtXO9FaAlKeP8RSJnVUDeyu4JXnrQyyHVVQbAfvn8bt/W0m4t4rZrzK+G
816jyBt2b/sKvHEm1hjFuPo3cBaS708XGpz3M2XgPvWbdLvpJo3m/im7HvRCBDF+
14jeWQ2bESsw5BsmRgSHP+G9As2I4yQ2nIo936YcVWe/Ht6BMAuRhLRBWtGEGFo9
0/EAbJhsFtzoaIpogpPjdR199I5pumdYxSE9kbeTe4Jn1oifjD0vukl4nF7xlZeK
WEvN8o01gypJjRSr7UbC9jP/sYuPr1/SLngXJlMtRwKJ3RmxaQucf/gtxpigT7DQ
AsbtOOnaEU1Tc0O2ASh8Z1X9HR7PLeMLDNkZPlO5aAzfENKo5CIlo/S0hL7w045C
36p1JsGZxTkGt/vVONwacM8Ed8Mk7ZUUrRZOY8mibNgXLwumKlWKQeY0dRWjKP9r
pZfLHnzW2SIZ/2E067A+1VbOn0HN6oE+qb0YuBjAdSx8Zx6YxqNR7+deugC/Zfxc
rli6cTMyxayxC/w2kg/aO/z6BwbIdr8Rmtbnjs7eo1fSWB3WX2EUVWM/HhlPPyZU
oYSDHL+4p+N7C1xkzHRVFadnsglly9L3ogjVUHkSSmw9I0l0JupPR0asGySUmU0z
H5YlH/fG9r92+erSu7lm1cd7olR7+cM+gAWOW4GsAtYFnN90Td29PlA6MTm29YG1
UzJvGrzcmcMbrAuCqnihXflnV3gvJcOET7ZH4xHuUQzxS/yuWpubOkj9o1wzQhuO
TS7jKxAEoymdcyjO5YyQlnwj7G/mzZeeXmobIwiZTnatJYf10rDDoFbQSOC7fHSZ
nZ7lXOQMzX3cUNTKiziuZipAIoMHS2SH9R6yBnFNnS5T/tadk2wkbMnONh54Rpz4
AyD2Q0jKa5iNMKs4boUaXXsNFMmiZr50tmXRWwmc/V8bjKKdqJ9nn0VyyyV8rdUO
HkRnBmCfXiG4yA9OV6EM/l0fB24LE0WmYBNcDRSD8R6FBOrlKx7AWtzPhZktNSPJ
BSj+z/k3+X7pPDTP5IBjFwXZzxeeA0CWXXx3cj/hDFp5LowzYf1XSxOz5oQNJYTL
lGM6aIiLAxq0uE3APMevSrizQUB4BT/Db3oRUYkzqmeCrXa4P1Dq8XoF5oEgDrd5
wYMxmsp5x3Bj98XFo6v3ZfOy1CcV+KsjRLaMCXaWVLsJiS0kgcNpoDD8Rwcdep0Y
mm2QB/dBpJippuQuud8jXUtXHHb7m2yhmp3HHc9PgQt4LZ8PQgUqclW28Ir0+Uyq
eww2HIu0tOpbwGLLab0Sch7ZaKQF3OlaxLoUeRUkIiqvSjHoo85mAOAhu0mxiPcn
urzkrzD8n8tpDwrrDeigsfaJ28EYeb/yMvodrAZZ/R1zCyjdi0qCeXCbA6Lj6xba
zswCzzw3yICyNmmD7B0iVkmdVB4r48IWnVE2PWq8mPwluCYlnwsJAwq7ytuBy0/U
EhS5r2oKjsiMl+5bI8HMp/xvG8+bWiVcTZn9sRORVNlEqDZ6hbZGUC+l3q6ZAIBr
rfs359NsvErUodWf8U316thlozL0406STaOTgAJA8iBZtu/r/XU3AKs6wm5NkNqp
/sYF3Cd95f0mdsnZ1AWoPPrQOo1xeZy9X1ABJOD2thXQVE+XG71FFBDVW7YpojsC
zi3jN0+a8Vf7tt8/r5MPhAde5nNVbNL2stBIgL8vRe0LLOkSVJQJKVcA2/n8ayEe
tb/iMlgI/bMY5OHbBvUzFSNsIZs01QfblC68GIU6ChRUbzQEvspxVfeZjoZsW/Ef
AZMAiBkitVbYpMBQOb9nNO5itqr9sBwHMvUcPPD2s7Pv1MCfO+34ZbV8OI9xshQx
WKfp175UXxDqLRH00WQeP9UShrl9Jx6ob3PvHV4Cy9LnWEYRh+CnTiYW6nYrq40Z
ssT+FFljao+WLjjpk8MP0Jx0LmKiYvs+didvvpVMoKYrd9aB3MIQNYLNXJecwCav
UTWI/noyKrsVtHMLsP37YtuauCFG2HlfwD36dNUv0vVgGUk77pM4At0uWOsl8OkB
vFaDyWuQtk4n8m/lf1I8E6CBr8tbRea5NkdPxoPQSlGaCmpHqj3VqCYF3Lueq2V2
k2AzAXdtJkbnIlZX1WGysLJ6JNQFLbXpgQ9OUQImLjvDWWBqQCjsLDYmKHaD2dUe
96h8lwUEEJaPpNkpQLutP/FqSHj0RFvH34cyDe202cJTqz3JxsyeIypAVgTM0jw0
r9upaEG2KJQQ+hjQBhuJGynLBNTsuK4GRbNliGQD9/igPGOPWB5LfyMySYpNENYM
WpU15Nj5nWwyO5X4Ox1BTCdX6rMlRZJKqNiyxal9CQoxwnvMPjkQuvg57E3NSzZK
Ocpw+pGtAeNOFFkMRCzXy0ynbrQRCH/JZn3U9PKsDw7vjA51MRrkDbjhwKMdbo2R
K8Ax6JTUOXExO06gwcBlGN7V7N59xevVftXsFtIIBhGwaJjWOyWjbw8XvRv8RmLC
v9PE4K6UohzS3DKrxh957GAmea4xpUiaKKMxPsC1lwEjDiGZK9So7AoSdltMLvlw
13tWQs1fT0PlX2qDmT/S+zcbfNt2rW/6ShARipL5+y/szDADw0aSgdFcDuzC9Zae
hxSrkGF1wV8J/2T0oDo6GZTTV6VbWHkKprUNXZcMP4WyvY0f0GA237653bWHS0RI
Nb1p/crRzOuZDLQNni1z3EGiE0vN8KEqOXD+54nc2oYsEB6wcw79ryvQguoiNnu5
uX6fIlRh7Q5X8/J5J5XKhFfikFqSix2Lxfnw/ftHgdGRBd7ht3G9MVCCXQoV9UZ2
AnOmLPNS/uAxYSf1qlFumMu6o79kUavtYjAMPVQMamkt7Kc6x4gSMOSxoC75UIxP
Hys6mhsl+9Y4FDCiGpuivxApAv/+lz5sW0kAGMGZRhF2j0kuXImo/wt7R8iq7cRV
v0/nlr0OWV52ozKXQmQaCAGYsqch1S+IcStnuTCU6NLwzSTppdnxUoS9YLITLlic
hwd0nq7v5weIU510OqtrlauhwQV0r15BSrDVo40Qm1xfRJQ0T4BRfYziQBEJWCIO
1xcyeWaxDmkMY1bxAQq4YH4eMD71T30NFhH63ugz0PAuyTS8YjlpCVI6oUpdEmP6
gU4GRU6ef7rsusD8+anVipPzvCVxl3TjrGCHtyk70kCX+3Aa1SlZ7YhNsMRmjON2
X5298m6yRwNJoTdaMOqP/lFSt/2Ki8q7Dh3B6poqev/+ZKtUbhjvN127YebnFkwS
EPjBMhcXD4P9bfydTUs37Pfuxjlpcx8C1jbm3yE1TIWY7/vqY7pol+mGy0LDXflI
KuKCP35YC7yo3oXzKaqNAbbyD7B60oN62CBgRkd0HQRwFY3z+jsChWdxZTqcy244
lPXkYRC6Uck17GWc+xi+RyEUA+idkV73qnseYUWoJrESn6Ph5qzBGKZqee8wKMjf
1INQ+c5PkC+bGzIKs/jb8Q/9z9jf9fjOycdvQJT1pcLyn+7C66Kw6WoMbLoRTjP5
YcHpJHeD6spw4O4Kf+WSsaypG3fk0+GTwtSwARWQsyx3+eRBo/EEesoybQ5EUzui
i3XwfYe7AMhAZdXn/c98X2eoZyTsvHjAtmzT1ETvJuNrB+r+27EEipyQh09T/GKb
lkXsdiW3NqK4ueBUaJQuWl2rDuBF9erGJ2TavKI6YWj2gI9jWhY6LmSVFU69maeU
tOyu4HEtjao+z/0uXkEK3QfNdWZ9iY1l1QbYMKuLxEDGivhaJ4GK4f5aYZ+Hel7Y
1Qj4DZLYI7XU35NwcoMI7Y0F+NCYnyXUG/OO31NWlvVY66B9dqwEf6dq1bLsOYku
NZ+b5ujZkBsngWp+d/KurGEIHy5Cin1L/7Y+VhR2UyDOT3e1rXIVC/pEaHrIDZUY
azIhULsduWZ5ll2T4HRmZD5F+dGIiRvXm7+58kjCn9X+V30b2tZ5wrHYaSgwaSMm
3IkbMVJNtlZdkSxaYzLqQ7BnMEvPfRJZQTtTViHey4LZfPiXZcGaYzrFouqe2bxI
qg1q//mEQ6GMvQVIt108+4+5GHrEiko7nkPSw3t6kGhCltpl03WDI9dXjHkJ2Rms
8lQkIey0Q5Vagixr9IfvgLnKnHJ9n86a0OvXxcPGXA98yTn85zCrnjI63FpaNEF7
3cbxhL0bkcFxe5+vK0Y6qkO2czR1KKsj26IPTbvX5yhIxHzSVwPO0imkESpgNjWt
AxvhkjYmcYzmbMtXqzbZ1vilEf1xvKwLNIBFpC4F5uCe7aUF/HClxPSWQfa113aK
OgBMbhKZfirs4u9CKCVOe1gGBNMEHvCy02BXEkdzyCC/CBdRGQRFfFN/YgNUYH4s
0jYf820M3jj8/XAD6tqB9ek9ktpIExlyBeLTKirzlDQ94nbYkOQH20l4QD0tlSiK
OA5+ollQyNFQ5xBw4udlBJNI3qvxC5a4gcpFpZaKDVc1HD9JN88+Y6fnOkO7ZDrW
qJpGeR6OVh+rS1WgZgNMwWDlHttVILzo+64fwJxHTyFJCQyGFc3h7HOPIv+Toctu
vvFjplSp50hLD5mK620jIFDGeYKTyARpjOIsEtumEOeDsAJhL84Orl/DslNyEonU
E0kGCJpgj9aQYJSqMu/XteGpAmAOpMEspSqH19KGTqzyAadfNzfg23nWPBtbXKHv
wUoOvArgzFUoZ9wt0a37BiO27JtPff6NBSHxOJuFb04QZSdx0e/XZZXRNdda3Xuy
/xVK3PSZXrUEInUUOUeRi8xSEh5b2UlfJFiy9Cep1BAS8TFx5g28WVUn2XfkTFoo
8gyc4Nj5v2Yb6+D64sWjdRBxlM19hKWdFzrpqdqEAbuAn16bcjEmOVdTVW72p45+
XoiPia76ANP8BpdPa7j+zlDEKmBxjxLYfcVMV+VWP4YJfmgg+QSGx1Z57YO03r3Q
YWXf4OnMFN0czev4U86vEkMYEsm/hD1FU5WzjXTYdBm1Lu/iEEfgk3Ze+6bim+Dc
ciW7UtN7ZMYq5VyuuZz/0uDQohSbBBi/36ZkXjEPG0OBQ7rAbYhNb130aGDFJKPY
Og9oSIgjOwQyndSKrC83Oy3CTAbBTrdaftF9lerWQUDGMrMMS03mjyqSgNNGofc9
gerjuYTwADT6MbzCxEtb/X6tAvbSTlNeF4WI7q1tNDTMDi2k9hQvWZ1LXBRMoeu9
Kvf7KFA/LhrZKTlIn6ndBtKOzj38rycGjqGGwiJNAVY4jdY2DVEwr+hZ8LYAimOr
2CA4j5GX4zUDiKGzY7QPn2xSbmWCrZ25kftKsl0leXb3S+kWaZiVpkGXJZ3UQvmb
bbKtIVY3qGC4Y47dPsXqkBbPa8aI+NgzFWZEFMyZDMyti9iYzNuaJK94GDyMZRTQ
NgAu4IbhWgGPVxjpCVjUGIad9RJqjGNECK1ZA1RLLnQReIIeUNQZSkVpLq79YEYY
oKwtku/WLs9kYY+qniI3kM/0tCF889uZCQ4svuacRNLOJj30o5hPDGaf52h3C7Hx
PZBc/TKIzJXT8Ben02HydGGdzPqc4vkNnntF1v3CyCjcvYWzICTij7s46CIdhRFN
3PhEV1RxE74T3Ic3G7yOdiBJnwZd3E29tgzf5gjv7ZijPuGrZdZdK/KuAfdk2iwZ
B18BAYe+xAUc2c9iWqE/wepQWipdeDAE+PApkF7u3ZrCjnKH+r9ZcVHLemZhiUtb
nqDXm9e28FqM7YAPf4yymjWmxQWIV5dbnYl9MfOG2dVFL4Mij4L2/sS/qqt+Wdh0
/st1Slj5FoVOnHsQ7GGMQtWoicguyTGB65hUeBigPJe3hGmEWEn324VJFhk2nYSH
C+8Ldp1oXlnGc0/V4yh2pw/Nr5R7FoY8drl7ErCZYbUD/7rxsXyOKQ/N5mlGCvlm
XH6JcwnYbF8aleGyD31LeRatH3d0co5kpizrUog5oc20IRmZh8F6P5/mJfaubgwa
TJxK7aIU3BN4dBtxtuskMYNjefdBmAsjMKyhTHRHM9nMyTNqG3zyCio6hVLJ8VtX
Vv4b2LW1rrF1Cs7Gi4viuOUUuvVsv5fQtOT4zCcECH5TQxPhF6+nzCRt46EyQGb5
RKUHom/isY/IRoC1OcC7jr0zAJpDo66ag8Gsv0h5IsB04j7m1jGNnrqT+WxUWBpq
UUp17lx9lZUEXuNPd2Xh9FnJ8HIWiWDVmB4afLBX/Cpj18l/c9tQ6wu+35k2nbvE
aFfrU3GsGqFHybbBclkXvFWeeTqnATmzrMGkNDjjtAVML6H3G8iJJy8bOkVNP5ei
Fn+X4q8xKyWSbAw7hcAzBp35xH1B2wdpPHqBNXdN2j6wsV7ZwV+3MK1+F+utajcP
uuQeQ9etQZZcLLEq0/BsaxORIdTTLgq8KyNs/ZBeXW8pgotLwUToReZ6+b46I5U4
x7tICj/zfFpjSbhI3CQQokT2w09JJl0S4iO4A+bvPzQBYAwOWKGvye0b7MuNeLrO
sH15T1UBRubHTL3I70SUAZcF9sheqdcht0XhkLxxWp4vRfIc4L4ruH5+cL6Gr48q
14byS8nIokL+nwlPIZXABB0eeWSe/3khAvg01/YCLyThxTHhy5COMq7H6v+y41AW
01Gtf92ReKwYh3wpvUI5bH22KQ56+rODqXW3GVPnTbVrZG2mc5IXGjLdfIZg1Ds7
rVOUjiaFbK0Cjkl+7q5FEcpv/m8+AsE9+SVdhT/HAzeE2VosQhqrtXgSXwfDpyfJ
e0gTzWBCVGPo/06j3EH+r2oIxs2O2kQ3EwwDr9yKhaSXzjdimciQ+VRBglf3LQqg
/V9DtfyDGXjhUPjraVhW4KFGDuN4FWdCWI0s0MKc1Wftc6aJQcqvpuwvrjuZuA0F
CRWZQqfETe914/ParfMBzXrn+eUBoKDqAvJmgDlJbCyDL3UAufLz9gWZ6O9oe49I
QkdeBOzvYACEX0ojuLH1euOUGY8jR7HAD6ygt2io0TNRF5YnEkmBhUlI1p/hBKkt
DE2FvY7UXzcNAbs+/+atMj0IfzWLr0if6h+sdINxVDdn8iJRljkja7GE/vc9TtZ3
Ameg0mSmOvzY6GLQSRqT2Ausdwatz8unYXABUOPNtnCm7eh2LsFXMyOLux9rL/jR
K9PoUUuvEVvx07iKaN/K+H2uL7RXCJxdriYkO1OgLqX/gpSsF2C8nj9quHFhqQRE
1hwnSZ6EhuQeK3TUg2KHVBw/GKpq1mJtxL5EDsg1On6/BdvcGuib/lNBMynbx/Qx
ZbMG1ve6VTKQ2f+0EzZM2gcBvDdKmsi2LzyBIjXoQzywK5NzRqaEL1adCyB9vGbQ
igiHQFz0jV2rPJm7QMuxMKWlWGCTDfXeztfgi2RkAboMrNkcYtDu4hY66PfxR3Va
HBVne913rXOzYn+/QxKuX+djW0x68BqDWyZa9P/7lMQA5HDoEIuJGS3lyYpN+PLW
0mCeEICRFnUEvaKs28ZyJRHCBSBP6GS/4uBdSI8mdZMR0SXf4afyFYxnri/vQkdJ
gzN0v7HjmdFUp9b9E5w9myJQ+nycGjXGMq1pHElNAERF+XsRBpWWBbLU2FO4/52I
PdtRuL6V9HvHV4n5Fhkes5mq9qdUQ2Xl70TTrQa529SDlDWDhDrR70x1YQKC2/4o
27NXkpDFbN8cCr3XJ0T/nnhMrTdw2zz6XliJsrlpUVehmiVPSkkKtK7fAbVl004C
UKFvgPCtCJHuB0YC1HGH9ZYhqulPp9I8+TubkqfyFt9o1lU5IwqVWLcjOhyTKKAh
oSvEsMydCoeX80urAS/ssFTM251Vr2JFzywhYC2Q2w/oSeNhB0/VXg4Gkv0EQCjo
0UBAq2/d5EeRuGtCikQlAqTvSFR8lWg+B4XZp+ioz6LogkFHiFI+sYD4heGpDv2N
VG5f4lt6VoGF3ESuD5N/BUJAqUc9UNhZCPlTFVkwoO7T0Y3R3C0yFoSKiuHBxPcs
AM+AKv4zA1+np/bKX9EHuGhcHzSt8Cw1bFVte0Z29gBqmGWtN0Z8RXyQkW85ucHj
UTx5C1dRN9a6K3pnMi1amavKs/NoykODyE8JFa40KhlDpE76vapbDK6h7QZUWySI
A++QHiS2RF89bVK+ScOQSl2jEMQwa076iVqv5Kcwlhc5wqYJp9rVE7I/s+roiO2b
xJgS19DVixarotrp1+Ahg0ihRlzUNCeT9MK3IeIZDvYfxe/lt0PAKC3iOlcd4rjw
4vloDgveRTp+RszSDNHU9wh1lsXEweTQrm3ZM5jVrg7hqFMOEeOn7F4bALV8JkVm
hhBQlO30L2fj2s0sFqPJwa+zFlbbJxWV11GHazTLSqP4QcaYrPe5xrK91Znyj5fg
YLoOMCkZpq+cCdnuCOMDNvAOG0ow8slSItEWEAePazws+wULNcBHRQZn9RMo+hPc
nZrcBEc3Qx4EszHgtumvWFz5sJnbS4kUCYDhJuUCwPXWpok/A6j5iS9Vd463g04T
uxjIrMgHHftu0bbAHXTO00tfZbn8Hw3xnGHesC3/v656w2SAhRsb7RcgVWRbHurp
LkVLC6nB9GIeV2qxIx11muWeZz9nuYcK+ujpN4d8wdBtVU4NGea/M7BP8JeZP9dn
1fM8GFKua9DEsSmqGm6IwszMM3m5YxLOU6jbimVxKF5B+ueF04me5Stt4gavDLmX
7Zcu9iHDW0kjjggTSuNHkR+5Yt8UKDobEHSnzSCEFGVQjPliL+Bl78rOhjJU4Gcz
/AUp1IgXPugEDHmS1+sWOowk5oaZ9mMDQshn3yokWK9ar/HoxhpFWqEYJ78z8ui3
K+miu3kmptjRxecNg0iHlSduR3lTaBF0ulaPsKYVHnFx51MersHrTj0p60JwgIK0
z5tlEH72j1OU4MYZVb/jfK+WhNU98dRLod/O8uX6XJFdSjxr7jyFlgY8x/nMCeMO
LkdfsgBGtMoJi66n8mSsqngp8H32w7FJhHdyEgxNBpq+1SPJsB+QqzaCwJFlcbGD
P5fXUzO8CdLKfN6J51lmV0Npkm5p7ZQkCB/AspeCYr/B9Kyty3K/dSfzHu0iZcca
rbxC8DXeeMAOBNf4yM5bY4Zs8ybjTnmx1spa4t1T1OhsnSOYMr3quIXKEz6HM1sk
Tet8bsyM9K4TAbGNPsI6+wsalmbH98FrdWsuCTcSRD2CrQQ61DTwqYQEvSr0wzW4
u3jdWYXxzae3SPDqtsVaf8ARJigR2ZTIYVKVy4Y3s2+E5M2/PTV2HCw3F1jQugbk
ObDf9HFIZyLnYxeyJdnQSjrqBjHIrLHS7fCtg54JAoseJpOqzgoABcmpTmtJGoob
uWNoGE6/V5u2WuFgBBEWz5IcIgcPOLdGqzqoIB1fTEpd5JbPuDsChSoRbR5RMSm4
plBx4NjTv4U8+zNqMwbG12YCjBbaLXxTOBWVoV35PLgFU2yhZXRmV9YM/sPACRXA
iaV0Gzl6rMl3qh71/uvc8USvQM23gGVsck9Dli6lsurKvGmxo9+i4L8hYe+JxuOL
l9aBUkAg4SJQN0RhsEla/XsucFkNz0MZOPcI0CtomfR95UpBLBV8gwpfIddkmfRk
v5nEU5buGEx0nrS06g9QnohaCfuXUCqjmFdbNCFwWlUTRtEjz2j22G3Y29FxO4oy
ty9pL5PM0NRKSYcdBQRBsicKp7s6EZeyzQLw87AjzazzYpdrZ0K2IQcxOrb/m20X
8FaDzRdsmhNPipg+q+i+XoJcN0c/JhT/Ky37eNPkaL6uKbci698DNq8IDgxlTOHO
XHq+g3R41ZhRLgHKgmuDItIaufX5LXG6T4SlWz3nDHOQnSoxcCA7nGkyBYACFKq1
XE3K54xWPVOAjh5D/A7+jdasYfR8g/lMw9vdQjRd+RE+FN40uKii2QCdcUmfhqph
FaMHMTH68s9bbJldh/bbTOM96cZobpeNgDCBSDKZo1DZ0OHTWvud3+fEfJBeq4Nu
/MRDVlvIB243REBmYcj6D2wHqhaEpfm4jlojqL9EUHoGxoghY0oDs//5UFIYktXR
HsEsm06T8/sKZVKveMjmGWNtn+lMxG9v8v2L5gkSvHAwNkjMFyJXzan8xWziYMFx
4+N24nK/u8uTjrTSBuEKqxjJKEqR35Q/zjnbjjasM8Ys/GHXRFMqJqeChNq2Ho0/
CxQLp4fN+hK0fQjzF91/z4Gn6arTVu7WFyLGrheC5w/5LMnml0SQpJHORP5Wey6o
1lBI7UJk//PQrDpHKAOX5AO/tJcTIRDf9pdn0UcmIau6iQyuBLqPv0tXvAN7nDwu
/lS+irBMJ7g6p/SFHFNVx+FwZlfqqCSefK+srESLNZZa7NSFvi8ZssG2NSKq4fOZ
osOftpf2Qe9PzsHmJfaH3agKpMhZuejfzOywWPPJH6l4cAP2Nb95AxwAwT1eH9mM
JAnCKLNRX6+gXbAK0qk79zdWxfBVgTW3LzcdVmFiWDmf3YABO75NLYeGTCT8Ir34
SWhz6Yd3GLD3hp8wskpITV03oX/GjD7t2Nx5n7Ry+CBuInWqWrPTpfYSYwIsNOW8
eR7XwOBcISENNE3Ib5DeFluP0Dmy0r3h2BssNgLq640ZEkiSsDyNg0lCqU6YHxJb
yEaZnZzft3WWpY/M+tBXfaMtJ4HalF4bfov4s2RzldXOPhZfDWkqjiSxJOrCMtop
bFMmXkGGLHedCrze+HfIF4KEMJJcICROUu1r9CLn4EuR/8miWiab+v9xGowo+phB
Y4+J8aCzahukSYIXYjyJtusIzDCE+QpBe8jbgPAlp3EKOy4nYrVWbLhQabjjlhDm
X2d9esrw5om1r5PDidAEgNipdpdan/rFMRNW95qZUYGolNiAK7ndXWREbshX3y51
2uydAyTYXOZacH5PIGik0AKQBWIFSxGieoSAX9tZ7DpU4mUwXxQF8fg/sKm6pp5J
X1w6Fv7KMnwoi+DOp3KU33qUtIkgKygMhzA1kVra0RtEsTYk0cG0Upj0xAGRTe60
MfmcItGjJv/cUzH83j02boLQHsNGbRCm8tkfdpVAlnQnDaQlu+E/4quxV+9ePoxp
qpmcw+lYGTzSA0GRvw2ZjBZZ0aTyDlwLGJUKA4VR3K/6P+raIhRt1u/kYQDpxjZ7
AoxxnhAtUAd/o9wOv7Nvc9UlBb7VhhASSmH574eJUBA2ye2UxIOKwhxo5A1X9suf
mriiMR+Wg0+TrTnHIpXrM2mXuLAOEnVhtUOpU+ak6zjh5nRqaf2dYurto2mXYNU0
mJNMHoXvASARBSzXf6lFz6CfwFq7COcNiFxE5Vj7pTuT+nzbBRhH0IXbVEf7Gc1W
ipaDAMJa20tdcqpmPg84Xlu4SkuzPkOdcu9bqeJjFxn+hb0alu2KZqZ3m/ZRtwYD
VoDeXCwVRDJCIZdHzfdtdIQfhHcl4AGqnA5gUzCNAo19iji7oVH2ycBI9OgIbmVR
dU5+ml9KCwOY0BwIIqNLZWpGipECpsNx/kXwdGj9quhCtHes2xMqhmfETSzcP0s9
4UTQw4NYlVz/MJKy6zUmGfdqs/ardYMUJpfrGyvi0wE9gRZJPhFx/00xuwLG0vXq
owmI7+yqB0I5jVOqxPaZ5jbBbR0j8A3ubJY040bv2Cq4fBxdkzftgiFXbhe4Vdsd
KzRKGzSQsvwzhUiVqhoHqWFByWbvF0M7i8biE0stQ6c/kYyjAKP633HnKQuQFGBy
JpBDnj7WjUVMwF4BCGhSFTwXOBpLVKKwb1bo0WVmRpoYU9HHmRXN8f2NQ0MLMCh+
megYdyuR8dub1jFTiKqri2cAvPLJR5ghdAqH/Pi02PNWtIzVRS6mUs0hqgZU3S/9
AZV9jj7MTgrnJj7zWRsK/+ATFz11xeeb/hs4cUqrMXx1/vu0phFwfC9t23LWtrd+
xhA+yl8aQo/UCPTY/Wu71//kglkhxyeceoEJsdlKYyJ6mC/JO69qUTLBouNIYQBG
qB6XrSyC1+T5NJrs+JILw1qhGWFjrZnDcuaSjxe78C8t9PQCF3DyMqLad7Ng/yCH
IUg/11o9hLo9Xp4d3UEImGM40AvtlQH4I2LMv2P9o0JO6Bx6oIhQ87SddBZABYhp
QOfu2lHlwSU56yFygyG+bZ6PbFi4PDJgtzpBXL8fu7vnsVDiLhpTMYMF82pKt39t
5t6adueUAHI6V4ujevW0vleiwH2Ho6YU6WFxLVJYDgcrUNs3aREwSyEQL+sUMG2N
DUJWS4+iWdnMCzvc5+lS1HRRQ2JhLabI3M7IKBGVD7s+0Skhb1ipWTQEDxn8yoCs
4B8SbHxUqLShQgRAMldcghqUbjZNDuLMSLFVp+f/KYPhfIGeloqT/YZDMqTPh+O9
MrZpf78bRsopUvTjjpwHNm/oBeJlY9j47X5ZWTJvshTJyGjGAV6BK+Jzf+xyAfra
tgI+OyBEKbg2Ep+nEQBoTaXHblJpm5XBC6v3bliE6os5DTI82nWONdmVFvQ8Pg8A
7v+uUseMVJrAd0glfWNSpivVzZ+lDpwDGKDQHrfWmm1gICooCWT/3znhwpLoHTex
VLnGrs2uUtr7NK5VJb5lR/oYRLa5C3r7iNonFTDHKfyrTQQev6i12w+0mnzc3E7a
QHcxGMwyy6gTqTUf2tpOH4DWNsUu8f38wzFxJOh4k51a1y1c+56Qy6uwW5kpBh2V
x5TfiqhrT2JAvbUeI7ERWwg8pvii890G4DrGiI6oXE5q+OKTDhwDwURgxglj8N+Y
n95yZFX9ljHBdgRAIOEDbkb9gPMO3PuDx2nrSDi4Qel1o8NpvXynNlS5po59iRE8
ZhhKDsx3PRsUgtKblA+tKL8gtHPJxV4+N1R67wJqSmKKrVZ0h+PbziK5us3Tyy1+
K0Y4p4FYAtVMwPpjJ5ygNXrLR9XceFopOfo8gc2f8v75PC+ynwS6y+QvKBfS3kbf
8Vg9O4qknDCfpGEuDlWt+Wsfcyzd/6I5W7uEePsLAsr/Db8jOlodfTkAxJmIm5nT
DZfBqh80KVnn4mpoOfmx9LPR066YboNhC2PFRN5i7934rLgagNTivOWKXUHYwmOd
deG03EPFfaPQ/19mXBRMfbhrh4KZOl3DitEVPWzZUcMAstcthe82xIOmP90MGBdt
8O5qAgS4KzwKTHIL869qgFCqEle5pTTG2qomjBMWu6j/VfTIAPGadsM41fdDGd8R
z5yWx6skzaitAjZxUp9Onz8VLq5MjsAkv9PRIOwMfXyxaKT7ZozQ096bhSYr/fnR
zFZk7ebXDJ4UjSOUC/4+8VZCv5wYvJ5sqDcWy82lKbVQugBQphuhnskAS2bGf7rv
RNiEtCyRrB3QfNErjoz+xCfdUiskaAatPaVh8og3qKqopJwqgzGLYXAePUk2jf5z
6tkmNG26wEiDgrFhOnR5Xp19tzE3HkZ9AwMYvEBDv4QpAreIuBat8N3PY8Gx6yJo
DKMz7bmj/khywxYgSiGoSjQ/r+/5am1txPzuvWQ8aQMUKJVmtJCHYSs8FYG2ciIz
rbS9iPsL/EkQEfEcnWwemzi9QhtarGlSvEEoMJDdYig1yN4SRPvVMbG7K4m07NMw
oVxX6FMBWSeOWM2cbZ6jLx0JaZ+0zq2i6V0H+J1oAZXyuKs8GIdDLNgoBwLfVbvF
yFG1HseTl+vE/tyfTz5xcDXFhMg2GQlnTT/sGWtryr/UJwiOazS9XexxBdSF2AQa
mL1L8H51f5GqnBy2UlU5x+Wg1tyIOxJt7Y21tpgBW13lIM0HCJxMIJ1MC/jfawJz
8UBAIYV48WT/Layc/I+ygikL2/iliUW8rL2WJS/bD38TLSoEuJwCnkAmd+PjVOH9
xqVlB2UadP1RouJCFFO86OJFk0eeYl+WoORJxdC8eKMxYb0wjvp5wEQQ2XWD+J46
0jXtj9+3OLUNpnEODLrB9IjC8RfsP1qYKRGWZyhFvHFCaQifs5pKDNoWLoDuQWdq
VcENKA2ys0LVEDXSFewrhzMgUV+70EXnMc/n8IoWsGwNTdJyKBUcILkzq5s8EDpG
2fnpA9Aq1Z3kBroJ3JoN2atYX+holFSpLvobiIKWmJCUwMD1aPdQi9E4w4Feh9wk
GGyasXgBZ710kBvQGKnMA7619zA9RbBakuorph1ji6SET483o0w9IUZ1hew4NvRw
HT3cI4z/0l2fyzkIoRZDPv0MlQM9n1OnsJn9nKXPzsw00PpXMUSy9qyi+mzP+5/g
5yYDF1+gl1Qf2g9IIjaOIKt5TQqUxY7w7CU6c1DWGPyNY6zf5wn9O4N7Y8QPMUib
YZFfmLuhnf274q6bdJTT6I4vF53jateFqiOzKVrDqMD9zD/ZJaNDmM8LbHby1rkO
Gy99DbJANxKHW7Z7W7/KgqPIAmSrEZw+4Ws/dvqLOkRoahxfhlo7vJ2FgKKJW+uv
mRMQItPTKTr4cLvB2ya4gA+UsqA9nPCt1JRDS/1QIzjvlayUvz7rzTbLa2SRk4SQ
qAEAtqJMDUtnlWer6ZBnADKobbk8UWuadrCEE6v7fZsnL7ZxEQ5tBGuwV8wlKB2W
hhBpYjoqxp19EGCkENfO/XuUjA/ioGgETQFwJixveDPmwVKrH4U2YRmqNRkFZ8ir
16hoOuyraDx9w8TBG1XKD9D0FCqceWRHNHG2hkEhKSGrIEWe0LyyUTrZBLH1pImC
QIa7GV/n2HrgceEf2faQMRcGmOhxx3GUZqtISnQzFQkpj+9nDawPDrHWzMaDBBE/
5h0DFpgUIzcxXuwgvDlYXOLYv0ZP40tp31v0awmNSberZfdjpCfpgIeu9WIHFoQM
36FeVu/CHzqcQsF13fRpR/zO3K9gxwafLn7RoYp5Vz2Oifziu1AqX6gsnR6G3pye
wj078I7Z1GOPya4kqBKok2g0Bznu//GJIj90RyRjWYaFDFOWpSsAyYKSQ5DaCyY1
09c8Qrhpro0okO3uX0f8IrQZ2hFqGvhN30NOjY9feImRsiEntO+JOZxN+BvvOiHb
UO4KztNvhkdxxr+sHaoUwawRMtzh1Q+F03MbzYGFDsvrHrMWt1oY6SEiG8Pc/SfG
zNK7e/6bqtQ59askK2LG+QoRHzFViGHlWonDXyvPRVwHwdVw0fbqfzFLy8MHgu5L
YZhwoI58ytlm0jYTBn4hXEXr3DZeII2XscU02f+1bNYs03ALT3K+eeRIq3TjBPqD
BRQ6WWG9pdxNViZ9BxSKltnL4jK0lTGyCxjzjuKlmujz/5trC5lKp44FHieL7Xa6
XXVzSTL/Objf3Z81NwEiP9cjo9EEu7+1nfdw/tu7pZPCPeLQgKP3eyRCUzZe4Q5y
chMjCzOaEYM5d7/VR6FLeOujkm1YbDILIS2B6kcny/hxOJJ5fMRuc9CUbjRV/Rr/
5PMVnbvNun7o3uzNgNV/fJmjifvUvien6Bfrt/tCJX04g5Jyb+Vi4OozPsmo32ll
GuUST4Auled3ExoBboWcZj+/nN4EZiyPuxf86dOf41hTF7rLohwykbcceI2BRMfJ
tt3h83+OJi73GYnF9YOKtrqScrNW+I957y4HVNMZaWthh8WamkipMIaGdtvo9VH2
1r6pVjlk60qzgTRYnHdWVy2y2qty9hefTPo97GKlf8P2NZMCQDAFzQODLxSNePeE
J2DlG6cogrdD3UNzbZzIUPyV/oP7RKOfR5P58w2/GrkCvspLQzrEpkjGV8msLGnZ
QvdrayuETxPLXBYvN4ixPFsBVxDVkr45EkQ1+XX7GcRX1VCItoWzxZsEFASL3Y7D
4k7SF4oMbAmriM1210FnLzwCvoC/lLc78g3Jz+COKhvEEXbw54MhpZMdUodyVv2s
bhDa4lwKt8EBBcaqMc9qBg0jUtzfKBuql+0kaSIotaMbJ6g1OVQoHaPQHolV9O32
jf2Cz+tDXsLoyJB1/reXmQfSGC9+q2ZJPGtsT0mzaWH1hPiRzaNaBs1dIPlb06wH
w2XlK9Om+R2HZ3dfOykw2ZzCxnzBb0McPjrDG4z1vH6L4prtjfUm1BQVcRvItpK9
le5LywUMQ0CEAULgIP0uYxhFq0ZY+xQ1y8Ioy1FFYxOGcc8HtyIchFArZB6Ye7h7
cgMEn148l98x50YmpUjwRCbjTD8UrKk9oWbzyRR/De+eNml9+DmnaihqnBT+KEtI
aGNUQV6fuqCC7+gQus7M3JdvGhSxmIJxomN6n5L9zMeCIdj9q0aVQwumxdC+oMco
z5v3zdT8JzflyJ63BSHpWpzrb9GE3sJ102xKC+Y2r+zDXHoS8pwHyD1XfkN3dZ5u
5k3bSYvacMux0pbedOtMjLxqDagM73UjTgw9izvajVheQYLSm0veMOyzX9CVo0/Z
SJTe7W+WaFtxQsslmRDRmmnV8ylky44QCRQaMy353ZN3WxqKC77X6jn/qKeG6nFi
sRmOQ/KVKK7WjmPDWNFvJyZ5OwFnbt4aSxbZcbA+gm9/NjbQc0TgsOGoGtr4WAnF
POqxN/QHS7H2n9dVI4KSv9OXNb342Hp3lC5F7B+mNnlByWcgCuSPc4keOYdzU5lD
MPSCEyqywI2ntDNAC8pZxvQ3RhR77B43hxaZJXEe/mSGFuSfKdEgUurcwy9Ab5Uj
eL5SRXM/noaEK7giY5tc5fTUwcXMQ1gju5qAf/dzE+pLWSTAoiVCTLcv5NZQ4iVD
vbk1cfffHje7wGX7Jn+ukzJ7FIZEyxUP9D7pugUakBDlatEzCNOanNEiMSQYYu4l
ut52ykorI/CrUMN2ngqbcxiPzA/tpkEYnoXx1vbwwzjIY7D5DGavmEuSumfEJKvW
39y3nRyrwNCHgl2KbGyYMyC8eAEnxn42ZkvZ+WxIVymC6LR1xVPiZZFH6k3hXW8A
r8jcUml6KJyqNwKaFNetAxDfgw1xXe1ZykQKrQS7Go/QSHRnmGCfxZFm0vW4ojTv
STMU5C6wOGQd6qUqzu7qUMaR/T0FsYfALMQitrbe1y4wtODAru21FZxgcmXElwny
z+BOi+ElaoTTFeYVZmGxJ2N2TV6a+6yLZIKmXz85i/TzThfzLY5NgHmG61WoqdKh
UARy6Fp6/ce/WoKWD6zG7CPwPqF96UUcz3drHkM6zJNLtR8NTjTom0Vcx5GzaLif
gT/zYGBM58FFEKqYm/F7+6qfgeI1a4cjANvX4mxsrjV7t9td+k94YmWqdQx0MGlt
VHfFzEelkp59bta0XuAZdhtmrBSiHebKWSLFI8PVviDvxhfIfI03tTZwh+NDFMbu
jO1e1IvsDambThz3EALENWkslRLMlTjV2kNm2MtwkblT5wlQDP4UVBlRlXoskBy6
nCukfrtkC6FWFdFNB4cdoe86FcDMK00qBEQ5ZptMXDUbnDpfDDpjzgaNRMPETv64
kkfBWhC73nbjb70YXQn+DWfzoRR5O5iBeIkbjeqB4QSHxXS88KjOSLFU7nll+t4+
93Fe8nxgSQXxxvRnT3CwqX5GG3I1r93AMI8/0Y9lmOJcejk/+WDd1v4xJsgYD68V
JmFUHO0ajtgMsBe2l1bkL1DXO8bym+vMkJGIpN/btoPQLJExGeVtFfpZrfAn/eY2
pCjMsLAsu/hezjDL1b09Rntw7Jw+OeerlZdmd+gBA7+V8Vy6s/4MYXxNKoLJhcgw
80OJSfQjuepZsQ4nRM0mFtHNJetMemoIf07d8aN6HwyF223iiy/geGsMBidpkdK0
+u0pHidND2y4v0gCdEXJdLwtA/bBoDILqwG0vS8y516BLyOgmLVYYSo4SrlsVY6E
HK4bjdd5Uu9X9NiKT/8osHlHJWI/hX9mVVw5Qy5jOSMyilFLW7c5nU9Yu0RLqYmV
MXmurfYvrSvkRwwJQe99M0WxfhhMX0bmZ1jtEFMXtEFw7hMx//sy+L6HKduySn0y
TcCEo6UL8ihOOYKlQ4oX8f98Zfr2pHbsl5/eBpG96PdFFQGTybuuX56Ho8fPmPUQ
R9yK+e+t8vLA3C7IoUvzLVxO3w3tFxz+kGmswOm61F3o0LL7FV363CzlHnb2GIr3
WizDtWLVWUJgbvuNywQQsYYBMfExifpNue2fAOX4LtoqKAKvmpuYPou/TzMR+kp2
uJ7ez9mxeRKBBCVq1rmZH3qk/u7XGJtvHxNJQvkHEhFdoR0VsPNO39ZxDngiHMx2
lit+4fHsldqSrwquakLp/DNlZIERzv9KoMUK/Q9ZzOI7jcXHBjSZJsubIgJGlf5u
FERxxOKuGPruHn/8g1hReEgm5MefAqNPa0A1HexSPsd6X0vCym2PL8PdCr7gVG6E
GrdORNntpQZAqVjtKK4DSliP8X83asnFqHdcg9xwwDqyr6Vhc840D/4nYF19r01a
/OOTI26mkzthWdBKjHjYpZ0Hza8CO2d2MXDIKuZ1Q/bfUl8Dwj8lCq4U8AyJDcz5
20acKlr8vAWVEEabio2w+Rcixc+UuFoQS5RoHOg5tPfCKjj9A5VNWq6dsE44OX7z
5VW873wCjLtCEylcr3Y9tqHUdckDVrdfd0MkNkZGfvWq7bwLy8HL6Hht6dJ4/BtP
5JuXp+TF6rCOEg1LguP15yG/KyW7RphK5IkvluPm8fxtGFEeLOFrY9664E33ET6N
mqyJVDPWFY6YAKnMa14Eu1hY7eyGKD4eeMIaBbgKw90ncwveXxzfUkxJhHSXpJDG
FcNm832pb2DjldUIKCAMQpKpB7T+goJlRQMRoBAafKHlodMkRJV/onpqCnk80h1v
VL64E4hb2O7VShzGzranGcijI5baqMGrn8ruPjXa+MK2OZHLYzcIIbhJkDptfwYr
4bLmnmK+teFQoYee0X9P4ZQKNm07e2nd9jbBQKBkPNyRWbR548QSmDMAWsrIbPVr
sP9jqhaj+CE0/g6t8OrI86QHv8IFQ0cBs5qZGGMGYiyCsABUgtFXp28a8R2KUVhx
2AgdpuB2QfJWF9Cbr2qxnTv6btwd5A+uA3rZUmYJ+ghD655i4Q38SjsNR/hij9p3
j/Q4EW0apk/QoUTRMWTQRo2hrayrU/Cps137QcnbH3IhjEvnoa1mJ5CDFLk/jRsl
AQx/ME5ehiAv4LT4lCbK81Urs348ArkFtufj0WxY0a5XAnuQwR/uprOVdKdHDonE
0O3Csj8YqIlrIqf7n6ZPADQYzBlq8j2r/hOYcaH9FQc9HBezqF7esIS6NRU+e70p
fWFF2HgIqkO6hq2z5qLyGkrjL47kCOuS7KCNjMTS9s7WZBEVJjMDcu6Ko65TpDz+
ufpEedLkyZZOGB5kuCPhWGETJueXQ84L0cj3Ppv8BDq7atgkP+vb3lm7mvcyt859
/PO7TRbBQ6/bheFPhxW+Fe8vPuT7UoTsA6Q8U/2Bm9XLmaBMap67GODDdwna/stH
3ZonyJ2PLKqHO1Lp+ea69XkKijbM5pWOFLAKacgGupUj0b2sUT1EZKMsYjkKSWsL
t6QJ5bwKOE1540EKrxd0IFYSEroMB3uMX43jUwi499HCbEUvOqC4r7iIRywic6Kt
RODDI8s9CNuC/zzxcyLC3K79gAEvT1CuWTg9UE2jXgnybCtCFo7QBYrl0JrVbah8
Zzxjn26xU9g1k4/4N1gu3LsgDd1d4u3RmkQS1/qy11JH4blg542OwMUeStS/hlHV
Jwn0YN7pNek5lE3K6ASREg6cmOqeg9UhwJLUuM+PGDKComn3m62GUU9G+w6na1yC
hytYXz37fMIqGTxKdwA5btRyJvuhdpJYU7TbrGFVCsx1SEtA5UAq+DCAEjtIQQwt
Qr9+GQ+fhq1SK/jWr4UF/qaks0hVaSca2kE3IUXBOGzs+Q1tZmRdZ3KyrefPqrHk
al5yVrFHV/R1DETrIIvERYJvDXVlnZJs5EKVaEwlhJVDbRlgl+36fbkJb20FGoyw
ASk5QXTp9aY69dSKvnygP30exzkf7PR+u13+MYrzzPq0mVP/5nrWKUhfYT+gBp2L
bflDxWYRHP71LiiwhHNq9oxKvVjfmHpVbQEXEYSrkIm02qfYXF//WBpDS5qoSCIm
dNf6w+ZVWSUPc0YPAVihvKBdBfaYEFFtAIceV4+Dl8qr/sTu6VWw+LcRebslOjn2
50tik9PN8xHnIDrGluvv02zEtrrzuRVhkcud0vdVGDlcfQ/hj22MEnCA5uNo6Q/B
MOi33UZSqaO+I2PXOoJHBH5107DPQnan2Tg5xDsYX1oNQwG03Q9uXhirZP3W9nyG
Rrl3Uh9LbLic5J8Vz0LAm3BqzkULAUfWlK7g3DV3p6XlKs+LSqjJOLQCUp1z2v5I
8YHui0FOmXQHCkDxiru/9IEeFDD1H6rlMs3VnHSmqbEL/BqbJ0FDA5H0XH0Di24H
HYBIoaoIgE8uT4to4g0RHVW9zh0WbnatMgA+8JHSyhSW65HCnTMsodpYSSbEwNlr
Q7iJCueUQ+rlGi12YtxUr8HDpCaZesOFHeNcfWXLnPBcyxi58zCvlZqQVdlaxNb4
czEjP7LLMSwAqVs2fkhVvptcuInCMcmTgQxVO+mucy16B2dShaJkjGIaL5wA9S01
ZeJEEO8n7B5yEn7IlzsqUOuJOxw4BTdsOflMQg2hr0URb9qvqQKQ2NwEzeqHbvFA
UoCI4ytsc/7YZ7S22Ro0MTxwlvPrcYJHWQ7DbtvEvaRbvK2bKG8FB+ID6oCZjegR
YNDkbsyldD3xP/D4gArcvG9Kq8EkGmTXHmjkxpe3FesmTRD/pcW0KrYvk58FVUaq
u+rfgzCI/Nm39K9ZzsFVm5emEkiCYo75U3YDfrZ4ybinuauNQAhNCZqlqVHxiQPY
I9wAieJpdsIHV5ROMPWWMBfDKRjrZpD4xzNfF5NVUNSOoIks4vKU5YIXukk0tIY8
Q7ovv25h6XrYauzStZvv+K30Hj1GZ97Lk1aYs3nwanX58c144BrOnIEPeD/hYhI+
z+2cxetfdE99Erdib+P4nGsdZ/OfnbjyZMSXlcVFYtoJNvYUybnU2v4/oFySWBCB
c5pmSarLNYtOyMbEr4K+JhYVDNPvm64/1Moa2H66oRk2y4ScE+vTr1TeNfPq1akj
nZb8Eh7qP9veIPkg/PCHLhbI/FQ292SlnZ0CHZf5EUxUWfdhdU6VVx+1m0kCvKU0
yXdjlC+w/1Nqkr4bJH3d3hKg7IKe3faatpDJSndy++VEnZbj+4700tOuJ5095iZZ
fyc2pTX6o2o8lmkOjWbERGYh57aKofgltpXmVP+a4mZPbmMy3qNpGxqc3bA0hzUj
p1S0ryDcQe4wL8lG/arKXyfuLsmTTrnnAzLFN0DHOXOInToMGIesPtcI1XDNG5YJ
j9tEuq1SxLe6b0j9KH0C/lvg3tDLUgsprLxVv49odB4ihgZyuHI6RWYNaxXaYK1E
pXlyf4geUmZGTa79xruXNHrhlz/1SNGIjo3ssbS3CkdJJb2vZY3+9yDf1dTdbsJ4
qRbHJKrzJIJlCFZkDlTE1NucOQavlvpY0M9h4OGuu7WApVAeZAueFJGd+8Ebx+Tz
P7b/448ujSvcIhgoZecEMdem4BHbemJZkroJYJxVqEiKX7B4nwOv0DwICJLdPw+h
ab8NURAo3NVTmCyfkpNyk4E8J1kzwnBDl0NDcw6YRW+4VUj3aFmjSm1g5JYAqec9
kark4AgUbze+kbH1obbLa/sW2qzhKZ3QmGTiEd540UeqjUAKzPNmUmuXK880aZl+
LE/kx5DEQcZlaS7HYTxRCX175m3Lz6DtwAXFTfcHmDmngVm93aBpCt5LOU7OjM6r
kp0dio7VpFBWEUQNPDG2tpLVNkAoggwFe3nxdGT7SqlmdXFKgwkAVRPP4CxRFXft
zYO5u0alW7Bk7yn6czt4wuiN1jeoRzFTEnqb6nRoSuqYI1THBV9NhDOIAs1makaZ
Irl5W01i0O1uqF0JPF6Bi3z+vXdsGXNzkuM9DqztC8F3glnN0nxpRXJvgRQhDDJm
b/YSQIUzSw5HJresFSUSebKWFOdVbEyBj1XIh6wwVBeE1B3m4LltJRXsQ1kiO/9r
uWOAGaWf5F1Rha14vN1iFMfpS4s8rhA6GnckbuDhW9G2iM5iRxNw5UE9KJ2xP8Cv
u7YJl1vppZNUHt1Kq5bdoBs0IalgLDCNSAdiOcukBANH0Nxydi9bW8QlvBRplEpE
9s2vFKeWhY8vngnQVyUzs+AcX+2I7VJkcs4Um4f9e7OiK/u0/zJkMfkB3wZHUetQ
kMUiUmCVYm4pXzaLkVOJbuNJ7xfAWenNxaHfWhkw5dXmIURNA6SC3vbbO+Zs5jZT
u43a/DDlVWRA1mwPGI48QZX8b18bV6dgngDuyeTqXI8Hn45zX9HxpJ3VLTeGVhyf
oN68jtrCUW/i1Bv96ygw4PePVxAEoTnxfkI1ihd6KRSAWxOciZSyACrkOq3TPf/s
Dm9qBIW816rLXry3hZw/41ita4/NCyiL8z1Niv1nFBJd3ZKvrAzcvuUwn6rpsBkn
bifofwfEytN9y59ehz/Pbgd5C4yYtgpusYSyyZ8aIt323QkeHZ8ILaj0q/OPB1ya
++pUexNXYx76yYu7sudv+KlOxvlNYxdNMtGf479KnM51Qnq95txSccBw5GwerEAt
AodV+fKPjrotc9CwnsW25nX6Jv8KH4kLaZLPyAV+8AGpwKjTKLiHrVtg1NlDPCEt
0RZbESSmO+r4Exop+sgEvu1zCsjd+r8+bSlrkbUuitFo0tIky3dsBGpFkSZBSTGg
JwylUOA6tKv+gCV2C+Puf168emF0vrxvpdit6QtVQy9JbfABbClfb7pJ4ne9M3fn
PLQdt8JUwKnE1FVUQDkBVhHS6BrZqZzvpqhiGw/cN0Cf2OHznXYsFrMiRS1M7Pfo
AnrN9ACSgLx9xziUtMW8xEnHOMomRJ82rTsdWC2YCc6YuzJwHaBgQI0AKj8jTtqd
erD/ur701D7awyt08PZ5F8Cf4mwwafpwiGGyA2ws9b7BS3YVKWKecU8t8tx7u0F7
H9UCVj1SGs1M31q4yiUB9oHiml0QWwhiodaiBiRnAVauQ2bte1Tk+xziVyZKAyGr
rnO4Pj7bVp1zi4Cc1Yoj63hPhbVIovmnNf7pVyTbpuyQYiGHbdEmz+NS6VWTKEho
upVHfNhDz+1oNuwp/ihlySuy5MhB+eAcw40iuAZ3FKQT2eMOXximaGfyFBDfqZqr
KhGkfMp2yVpQUNqM58vK5VfLOElVsjofdKY/BUJopAmFxzqfYzyT95BefAQRfAkM
sSEGVaHnzYc+boVD05MfslGAYHYzXLDj4vKQfVCTiKdfAdDvZHM0zWMJ1eeHVoSX
sPWcl9ab1YU0Av9DDT2UH1G/SRn+rG6WNBzulOMgTN8U7fcDA/vioSeyfGxNGVkg
e0Gx+CTv4i5naPpcuKUtadYG7VnEvWVW7zCK0LmH4ECI95vmEYlckNWZEeNGmOpw
4eLTtoRkG1x7xrPHb06O2MKfqs0dKkmHFhLzVPJ8NTRZFTB6t8Gaa06mWusxrwFI
jgbRMIDZ/f7evwha4Tb3A9NZV8bA4Q+Y0MM+pz2kar1dggEvXeJH9xu2rpKJqQWa
pzMyV3mNapK8qGVjk0/rupoE9UrP1p1Z56Fz9YYAP3OukeueMA1u7AdpPnD0xu/H
fdOcnhYchgvi9Y8uLaogKm3OZYzOBpTET8JU40EMwS6xrpLRHtibDlUUd8Ob2uGA
YTuX9T6PHvw9D7va2hMlYPeN4T78oY+O3BRbQ9deFPENW1vCj4wHsTr7lzaf072c
nsp3HDqNJY7Q14s/Be+UFzR9gRWaBnk4FIyAdxeWQVCLoji817ZQDNSgrjgQ6f8v
Im9aCzVfiwBfX5uGcGoF5PxAgIAJ8QHubeKA4v8CHtqtkvaQSvSL2RqmEVm7jk/c
T7n6etlkbmUhYNWiJAQoSur5OUq+NkiiQnFdA/LzLPaXuDHcvvfw0vdEk/7AipTL
/7ZAwYePjGw31zszenUgwrKz6Ijo43jI09Ocz+faRo4MIPPy85mC9lGFF7s1g9N7
7cfE47osVsjOvtVPqR/GfW4vIEEuBKv2TRfc35YZ6KcmwRAzUJzNzDpqquqcagEj
T0qgjmu0Rp4QFkCNsvUkVlKtkdvnCZPdTQ7TJb7NHSirP9WJGpAWIgU2iu0fR20z
R80jhiO1NtxiYdzIg0BTgrdIsS2MzwlfWRWWeG2frlU9sMnO4eXA/tcsyg3q4BlA
JDNhnPgDmrg7eKE41/e013GhGB4V3lCuA5ibLD/aHyoLnWoXcC/Y29hldIUdd8L8
zL9s60hdcgZJIT0UYc5mkSAOE8EOpUJDWGBfA18p36oDMNEjX6QbmqvckAQIaRaX
uvPjNuoFIVhFYgwmy7kDodvs77/oFaUONikL4DRpd2+6pb9gTJcde2PcwVBaHRCT
4D4BY8HU5chM1L2iO9WKnLUIgmcKEhS82RFpDEtVzzhFaX4kN29nNzF1seYSbmGP
64bPExZpJRQgVd8NEkDK3TttWlt/mGdF248OLrhjyUW0z15CeaA2erZqaxKSeO+f
Ohy2+nDEVXGRoUGv6VDqzutnWE38UOEgZL8T0R897D6O+MVhMK+6+HNCMLwBURzc
VCJEDcVXtxDQ+CV8iYu71FUPPF1cUBr3/2rqwAmpXPCCD3t2tcVYq7tln9znAJ5g
puAa34V8d8Y8p72lLvYtQPLzVlsb0BafPCrNnWMfKfz62Eh1kZk5Q3Wf4Whabfy6
fduvcGA64j+0RtpvuTOMgkx4aXp/UbA1kevP1+gQWDJh+ogKyAoSXR7ABUrVDLPE
JIE6q33NbyX9WmfjVxOl0eISVK8TRzmCZJAG6SldGGSvJ29Oy3x3WT9Bhf4io6g9
9HFyzMVqk0gbQhpClWzYSoqPX8eYmyOb+cflb7/PL8HvbPbpZSon3lCBlc4hLGCA
2tmJFIZKVhjSxdvylmRv2P2C6wWF+gAMUH8iHikcSDlsHKtjzJL9s4QKq7vSnXko
3xdbWZgwcVnT98JCT38IocNFgsvvabXx3yhM96gDYA829T+2CZ2BbVAm0aWF3iKg
8/r+wWRUco+mqp8xUjA6wGiRqRw9Kd+kqV+tvS470hUKrWCtSBxcD1vYK+E6Fbyj
+qdWjaR/pi0Xj/mkoToQP/a7K7YQimqr+HoYienhy8XpD6CPmVpUiIAlJA2VYgu3
uj8bwN9/nLuiqPsKC4fHkv5DsS0ip612yzjekytDwVh0AUH7OEIrXleEm7d62J1l
qA7OYN92S+kVfqnuDpAhBgdZ3rK+zuGQwAl/BxCGP4q3wJ8f6444IlnWhxYHvfaJ
3vHhgjIPdKy5ZzmpksvtSOlmYlNeDpTG8FZhY2BOFxA7xUT11ezqqYm6q4ZZx05Z
4mxTOGs4TRkR5l820V7STH6MV7rk+tG/uCvRL1MVhs2rfFqAYFce0f2HzBr1YIGT
GirBHAWXxyZNPqyfUP8KYcELilnAeGLid0qEkYjnQm8pvIvcYALJla2k25bVP5/m
jPRQ9u2ZS2prfn8ucXEzb72pMRz78tTT+pgcSxuSoU5w0wpYNJA+AJWh/jPZHm4s
JdSwyae2QpeJYDEVaVyARLr7L093E8P6j7diBJ/nVvv62fXAe3qfGROzhkGUEapr
B3AoI5biYDlVKqmb8M2NfGXI2bpZJ0FjlMUdJiCiFUUNJVtA9XvkEsjsQWhhrUrp
Jf3qXoIP66KuDbloV1sXJzGRFk1uPmYTjG14dN9QjtTS6QQ19cE2sDv+9yR4FXtx
h2KQhRPXluHBaJtbqenzVw/2dDnO2FyJ0/xi706TdiqaViFPzfYJ0dlWwvPRtKu9
Lk82efZKCgnawZNyPWwrDDTz9tODF+jDUvKqAWB241iUIFcxPOyJO35Gv+suCuFG
ywH3PjCA7JeNoM1LSdkcQupYjjYSvNyFNwO2KEMnIuR2mOJ7HVQtrSKNjW3XrioL
sufGf/URbqooAqAjeCKq/u9T3uCTfppqmhQgjvMLKe/Zi7BzAYs073N3VnjVZqis
bJ1ChgI485+RiC6ijZGXGdY1rPwvdsmEOr2vqgSSe3u2/SGNFbY1pPsdqw4kB+9J
Jzb0e2Uk8WmrvI/+2saian7q4S10mzHUyM6n+txug4SxjLF6YmzCbQe/2/a1cKo4
rIWWEeZM8l+ZFGCX1aPzT096615Rz8lAB0cNuSNLxii74NR/qMF2kcSJAh2ow+nA
ZBqCEzGXGy1/I5iqzpBMgvGDSW+FuxWbnwPWP2bA1sfto6YYFvgzU6BgCYgyh7+K
g/R36gzuEn+ivWgMDkJMOTj6z5DBB6BYj4P92WOJVuVWIyGdcJchLJYlpXg6+Wjv
uk2GHt+LwbphfmPCFpDiEcV3YCkB/nj7Nw2nIaJ7HPoiMnnqdHfjLiP+CZj8OyLZ
BRc4DSfv3mLYr7NcUrcMYco4djbod1kwRI7tYRXj4UNp5w5sO2xCQ6AHwvFPpevx
CLweBVzE5Zcx+4WjlnKQbP+iIV4HnZHDsIjP3jFOQUj/3UxLBEwlel4Momq3DYZ4
D+uqWiqP8mAIpp8SItSP8LKu+na2LsH5oBEp63AWDsk49TVKRF1LDApK67prSaIn
MGvL4NYHPPVYcC/kcfRrakDFGIkmvSBC/BJQDoDv39/OtdPkHHDq7jDPt1XygPzf
whpt5MgXTziVYHVx/a5dQVl2q/GUhRT99PdHQoRAZkxZ7K5H62ce0PwaNz7rIT4g
Cbu6yceRHBJht4IzPUGU/kjlFtghWUk/yIfpISTK9tCK4tT9BOibtvI74TeCdB5b
3viW+rLsc2uklXCwpQS3vrMX1VWb/AEp0/sljPQT5VPv0UCLzZRN0zNrbYPHjP0E
Z5oipQLo4fbqZgtQP55XJZn0KKAuI8O3ZxvkM/wul3pB9deCRgl4O5pY4gZ26zcZ
Js/pHwTnKKT2OZMLEBMm4IUeSifXxUIPFkkFhHbSOpNeJ7THKAifA7OKV19M8FfH
/m3KYvt6A8rkF9CCLXAwAzFexnRca6ti93S3deSuUiiSahwVypVfTt7pQvO1+3X9
9Q/99Bd+nyszJ/a8UyvkeRb5/joDfDP0ozIfSUhXjo24VyX/LTNKU1TqBCHLOmef
gCULjFyLY+42+hL2rbftXulP7MvP+8e84ZVlNJoU/7j0EWyZCLv+Ty8HXqocoF0Q
iZXqis5Jrc0f8a7d+7tMt1ho/ykf/EQO+Uosfe0ouG0egE5uulsB+EC8njr0vc9Y
I4vlNFguOItib/jZwkcRFPnMI8OhuzNUE98ZruF0A3pLNWOQ8FltCT9+3ON21fGy
UhqUpR8h3EUJTmhKfci/MlSR9anSI5MimOS3jjaiPO4Dj2YfmzMZg0dfd8P3cedy
YBNALbUPvP6sjBfsoXliDrHkfuGBX0nxfSAHp5Zmcl8IrsCuFTPwvnayrckiztLH
mbGm3rQ2Il66mZdtzZZTGscEPArSyvUbhfyda/MjP0lZVyobTYJODlz1U6hItYZ5
3F1ekw+Bora4cE6UjcR4ay2KmKj+6KKp1irW2S2zHLYi39uPjmXuk1N+DYqJpi4G
a1Vp1rgArewf6lILRretMVKSv5tSS7XKivR+j8iMmfiZkAGws4yu1VzsrhB6pO4V
TaDWWAFF+pTwB1FH8aDE1h/mjOf+H7W6jmyh7Ec9Vg5quYh6vtZ7S2zk/rhbEirA
nqASvKHu0CRnWljk55Dd4P9+Xnk0vCS5oZvcFupOqLtHNPEndX1fbh7aQlXQKRsX
dhnKR2/+uXA6dCwH2B42ZYX/mRAkCWXRTmNAzv34kbv61860m0TA3rF0358oJRl0
jsf1ObxdDPgrRTDT6P4L8DtrYzR9luN5Gfe3Jn7BUi71Qc8cuFUY63vhHC0FF30m
zYY2yh677AbymEOTs6B1aEVTRQXXfIpTvve7gnh7Hs4qZOmZ5hjTA8QtjTufSRnX
+m7PjKyDb67i4wCq7fjg3R5fxgyDPfg2n3cV/6uI65IMaX6Sch3rCJZdRzjFwZfc
2vCzLLi3943x5SWRjoUEioZ/chJiUPnb0mX8tdz5exTtrb95C555aIU2qFLHkEXn
xp7nehPZSrJO8szQ7cUhngpmM4P1DOIK996ltNnjdxU/j/dtcp7GrH9NAPYM7Knm
whb1y9KYNmOumJ7U66CIIe8/YgDdrvQGaSK5qtMeYG94H4AD2E7Ls2aIOGXMIW+n
dTP60qaUWbwCNZHNTYt7fXShZkDEsaY3PzOYKSlbqB2oW9CXxABX9xN0gjTEkD6a
9kNebc+Kwcdv2GdV/wNavOFBZA1NkbDtMqmk5MIVQ6TRwO1JoINEVCQfWG0R0ur6
SFt2v4VA8g/KkjJayStAgHgGUKxXejmhU7MYUVCIsn3UFEfZ/2oHWrAa2+SIDDqX
hnIxNxIxanFWtFElM9GI2yehuBraRw/lVbRo7Bc8QI26tSth5muNfQb59prhs/BP
6SzYHDwKOcf5XGHNMWavh5XXn1qXt9OzQaCTq2pj5kVeHFoHVM/kmVpycaHfMaMH
dABGvtNoqAwd7VntuxaDMMoJFDKx1l1itdg9QSwu4ttn/4BjFfPA3ChtktXR6kCx
W07kdQHBFIk4xLQW8vubt5x8h0CsqThboLoX7OE0u1Ur+hr+lpc5A52bVUvK3uYK
uboyY+oT0ZP/HYzR/LCFv5SVWyNYa1DgXAcX3T6ih20VtOY6sO7zoG1dKx2yB8VJ
4JVzi/3u5G3hK6XMGr/fnWejRUUyl08lRPivS530X8KJ2P989hwmCsyg6AbS+wLj
IQBUC9f0pj53eODK0fCZRXcXv+u4Kta5chJWb1ojVgJrLX5l4iwiliWFczqO3EQr
xcPdrW34KatCWNFWz2a0Cq+A+IEvwOp5VZI/2o3HoJ69OL7CGzwDq4TMKaBVaUwy
YBXU6fGf5W8rQQFi/A8n76onQC6Y5ET6uFLS8gwXa5DYvtSa4JLMOV/gGpjzd58x
EQm1VuIZZ2Tp2cYjhnm0MkrD0ONP1uiT06pMJyPBgfjowVrxeKIE29LR/a72oJbd
NxiKkD+Db1L5x4rnriTPMK3jHwp95O6XZQwK4FGIZgHOY7PWgjwHE+G4VCAg+vy1
GL3enFJG2/UD+8NmvSGw4EqqzEN+XgNAX9S2aktOjrLifPh6D01K38b0c4T5T+IO
fo+9BmBMmzvj1CYhatBoHnruDFipHvLZnkQoyzwKGs0Kh9QQ2gQS59C99jtLi9l3
opMiK+tcYI8Tck6YqEhYSTnXGv44ATQzzJM9OYtMRnNW7SDBJXZpB6Ha5EhkcfDt
pglyBfUEdnNFHNROymlrSi8KOpd57SFc3qZXqx6TH0UzLxlIXJYUj2YTw+asLLzJ
g1llWCOn9DsflYK1injICQJcYDUAts3C32fEULjEDv8Jt8y2pvoNESMjHC9uMlbZ
0fkGzOqtf/u1klog8Depxb9ED8hLM60KohxRljFk6qTh1IN4+AsoJ4moeaiXlbIf
dcANWc9/6x/7C2t8dyr81ySbKGXlCjzcA1slVKyvYrcb1Hlgdf2fxHFafJBtxn43
K6eCpmPGqFYGI73CLDbFW4PZq1JULwafB0LWLj87DbcezyQMSYhKIIbO+XpSoC74
N71Nu6Zm6z4GYmRPr7hY/vOHMzhmrU8PpgPKSK1GABlFyXMzLi4+tGlt9cwbVkKg
UV/zlgI9baqcaIzSgsPk0Gf1TMmjhST3BYOyMR2i8wdP4y5+/RbkULEb3u/x7AhP
ScIDvR4KYD7dU0NfbzjcM7/M2FRaGxOM9+V1xEP5uFumXnzEci7AGw6GDLsmnWxc
Ox2ykhbgHjdd/9jHe5cP4Niv5roBiWhCYDu96WTWt2g6sy5a4rFEiSbC/AuVc5JM
yh6hXjTUyrXBPWA5ajLSx4VqlRf03veSV1WnXb8+Tu3hlIL5/3KD2s8ViaAj+fR4
yraygJKaFs8BxP7ChjF83qdLPWfhIrIKqv0AQnHd+ddSHCmEAIXLgxD7EsmnVZN8
F954uTAEpCX1yqV+07oB4S5l7w+D+DIn/FoVzzQMZf0H9/A6aTV5Z+SQDWrYnPA2
zn49Ay31NpQiMOBiW+laNWpEdAZWgloVX5zuh/FXnIYwfYaxs5zEHiCp5tNnlsO+
OuJVDaWYd3Z8ViKbaVMAhNlrGDSvdiUM6qnNEDdE23b/+nxMt9hSi2/eDklyN5RH
UDJO3WMk+VHCl8ndkDPIfcmHH2Rv9XN5jhTN61P21HPfaBMNIuQDlUH4jLNw+d9E
3UX9MDeMbXg4kxiMICQgCHJHTCkrd+C13lX52kYceo/51JhxApmGTVasRAtMyWjv
wiofHRGgYiWlfUS3ZVsJ1TmnC4DjgvauCUluwNmCc0cCWQRV2LjoyFUsJpfCWXqz
FZiy04UrWHfJQ2Y+E0H0PGHqBmASGzxcFXECLBSawEtKR2cXD9NlRSYnjeknE4ny
iGPvCZP/AyjRzopn7Z24ncxogA4pCn5u7ijy4yH/9lATrJ3SWULwz2nCgA59AVUy
56JqQtD6Jrry73K9Y6jK1swXTKy+3c+wv8hfmjXvXypQWu7dUJQPTF5LG4fMU5hX
79J1QSZPhN9XY6ZAOjKlb9WgtAPBTBmBFInm5xw0mCaTZIJOv7NEEh+W1E4zLtKY
1XCMMRxXh/vjFvs9kgSfKaGOJ5GNQflODLYiYAf6RdMfrvx3dLTpa3KQ5QdK7mrZ
JJ91t/6oSq4TUjn5AXmFU2VjLlOasISthbo6CeLSGrjImNTed6F35jWOYHbY7m+Y
uLl3A4cBGEk6GpO3BNGAMswMP6eDtBB0KnlJI8I8bOugiAxsb6mJ66D0cVJ1trnn
5ECLUe1AOZZ2nxqNAy/DzHl/u4rjowgfdX4QUWRKCEuLlqniZbiaN4t4Hj+0tlBU
YDSI08SlpgO31ZPOx0zxM7GC6aqFEA75Sl/pgcH4fR4M2x/x6RvnlgxrOiAb5Sck
5x0cx30pNAaetCiZjE1tQnEq3NpEf5dZXdrHTkQWrJp69sFFVWiCSf3eGO7v8mHm
pmippzctUYPtZOrWN3f5poJl6B+ZhXood34eHvdPb0hQmYZM64OSqWjMnMnOIjln
eSTJraJpgu2HSlvJ99fJPDa6vyS/I/WkVDtipJWTZj3T655N2ok6VNtQ5wOy5IbR
VGUAA2aOWLFQEoaefdPLqQfST4Du6IXhnYh8NE8WEGuYdu9u2TlN32QYdSFFmt8C
XSlejFFQmenpTTw1LgGj+5ppas+lv3uDhIDNGw7dv+gNagf6dHuk19rK0dURgE87
0/K2uvODTs6atLqAwUpqR4ycl7Qr4Qpj01bR9sdCNUcGynTV0kWinnVgjiA/W3WY
nuOmQxEyGkLhm+rkKvTm/3qFlaLO5nvgbs7cpV2ag/Yr3EST9KefGvl2MXZVkN0F
OwnxdViMv2chSGwNog+QPrmkJgtefUMFetAb5+y36jnW2EljlN3F+z6ccQtP4km9
nmWUzj9+lXXvoee131b8rMYSuQgZyR5xeG/IFKASwsz0mFHFr50Jknp0VPMXyJFo
x05ykZ1duyN+xcJGCniAhsBECHwZomSoMn88bydt9DxyQ888eZlk4CIvrgaouSip
YJ4rJKej0r4/1rlhhQiuIadZQdVuXUzoMMGcJmD0iKHH2TvHDDEYRLH6tjFB1A4a
CYKjV7R9jcrMNcMb/Q/dsWtBdmvKzw4U05OasPEj++I6WBACXvLa1jkAAaFZPD5w
TqRwd4BaVKsS0rUC5iojkbr8WUfr0aWJDO7xuKbN4SZQ9I0f2qZyHnm+ZfhBNxo0
37QfUfWLj4gyu/bCHvdluBwigRiGxZHqaj/ubT15gb1gXn/sOc3qYPU8n8WBXZwy
lpiU3uy4+xSzO2yU4Bl4aTAm1L0Wl8CejAj3DOZzvUcLDHIc3Z5otnXMjoIw1i5T
Ijjvku6LGK3s648/5kykRbMbsDKitp3NREpxCdvJQLEVmkLN9mb3AfY6Fsuquo9g
hPznQ1MEbm2Nt6exfp8txuHfBkMgc7skJqJbwtM+LIplr63PCGqBv+Nje6UbisYY
UPj6pdOYfrC40kUO3uDYq8rEG2bFARErfihLeeHch/6a0w1NtcExukubuwS0ZQUi
kMAGaExj2xVUCHPLX8+3dzA0Le65/V1+sph+U54OqgI91e0lzaglQMkmkI468Q0R
34g+cdCq+2Hk1ml8IqqW2IImiEkaKOJw8c0PQ5CAjTEBTucJ4LbvtZpTc4+4Le+L
8Oia3EZCosq7DhO19Zh3B7K0OtArqy7ryJKYNH3j4d5g+o3SYrbcyp1ZQq/pUpmH
FPEUg8cZTnGbzxAke52hXGA23WYqK/jzdxM25UQT+O/4Xuj8Dr8PP1ew5xiuNGBp
nQtZA+3N0d400OlIYG+58fv+CFpbMIC0ydHFOKDwgWhxZAyAIgkpIt0hBX/CLCWx
lD9Jw/0GIbmeDAeocV4KaL6hkRyhbM8k76ikW3HU+NpoalINNwVB+fo2ikYFuouF
F1+n5RyKlGzj7bsEOvyKqHYk6pA0jW8iBZuaLrT1JodULJFAiATvYIz3K8leLgKz
FMpYQWzjLAwAP0UDQ/pjj0yKJot7GgLoD/g6U+Em76GIP7zr7QvbOIamZU0Y2Z+3
DvkeU+3PHHNsTvjfSnj4u/V2iUK2Ra8cNaoa7k4orzseNvInsRIHW0a4Ztm51gZ+
s+n2pjBJZYVpTau0XH9UZUb5yWzBLfmyndSMV/I4A7/4qLFnXs43f8VpvmpmdS2y
WpxdSHG009pAkdvEQfjbYQScDXcWZX2mL53U0zM5CSSKPElp8bkugb9zvBhGlgGa
PK2vrbUWnJHmDxR1c3874A5SJcmrJ4+i+BtTBeaURjEmKHwVmHeA9s9zKXEVqv1j
BcsBfm7cqMxm0vBOLFKpicXqN3RgXYoRFdJyH9ru4qNz5cgLwCe2323bgRtp/o9h
WAtI9fobi6VqWHY1dGqa+niNbK7N8C4/v/qBV3XH136kTSU7nghpzeGWYF8DtHWa
tCO1iIXp7G9frPCSBzeow03UMEE9YgH2yQXSJGqt4helC3sYuv8nf5wiZ85Yln6w
dlplkOzNPlb0tCtC30ewjJRnY7vyzcr8TwNFXPFEBD/SXZLqGuTZfL434ES7IZai
hnG7/PT/MLLAVYp5kgJxntRe281wR+o9ID8/4U/Sf+lW+nmSNEya/BlhjSmjA861
rxyB9puNJF6ckjHstdTNKKymWsDZmlUhXPy2pA1OsxE6g3ZotfryI15HqI2klMfN
l7u+8Sg4ZHpgRhq68BTThSCmulTsTpO0JJvuTuJTDkZ8bZ+T+9MP4RRwoKK2oCi6
tpYkyTPHaNfrP8XPmrfjChdqziKvBKx3KBLGASPfX2ueX9FkG53U7qN07hVuPRpJ
B0/Xxm1nkGNXuPXGbdhKFcTtEb7sQdCSgAW6ybTiiZWgukioXlpHKQQ8A8aAuUlr
qkTvp0wBKMVq/bXn+uE5ei3HIaj0S6/V8n8uu3/tkMEORIv2Kcwv3KkQQjA/MWc0
LkKPqN5gm4MxlMDBpx4rrC0/7JneZuiEIOSS6MTftaSxV0GgiKK/F8EROr8pYqYS
6B6Vu2dQ9IoMJ8QfgFAP7WdPMI4CPVXwrL0uNjwUN8WILEE+Nj9QyojrdsZj9pjW
jDdGTnhzvAfcACFWrfNhNoiFK9+wueZwSKyDzynYGjPqlTaXTkV9Ny3GmZWjRRC4
fRTb3iPKqLnp6z6HFGdqX5R9YS2p/Dk5ECYzjEjqGMQffYVLJ/yW1Y4lS0X6FXAs
He2QAiGhuZPueOKNqLXIRuNXGnRf5KtLPRYdsTPsIJuiZuNstT6ztM3sFWXbkiIi
HgNWI8LbL/0ZL2D3mTalX6EU/WU49cAF9ziOMDGK8dnMD84wfXr+c7TWX1j0qNxX
2LIba9NPOCS4YC8HJ+NSSCJFse19CTo3369lWzaj5zjpsy3k4bxRlHyIoQLAY27T
MHZS2ndF8NphsscD9chrbJzypltnwfC44H8nW5MbraoswE4/+lWrDj56fRoNMhOe
RWICKlZ2Rny9gg9gZuZo+4IftZAGOWE2JDRnkOl6Dg6LhBGeptbBItQ6B+uMew8D
++gcsHkWP2AuFfOukgI8HLSTQm+AnG/qdcyCuaVWJrb6SAuKo/8y3cSxis0T6zx/
3IlF7iLtQ9hylBhBj5NnOr34wdkwCgE1AZOZV10Qaj416kwHUvMrDtFJDXtv//Z8
IhzGwnSAVszRfDMnvSImsgC/W4nIaXPWcq2evWwI/SLoXKbVmc49aJAvf+CgRO6n
qd9Id5srHoQ4WYd/IBlSvYDl95NOWx5NeLB1bFDXiojXwcKeLcd4Fxl/GJ2lfDCm
wr8GojMVnuIgEZUuNGQEhxl2FeSfoHwkXokTUXt9pX4DxzuMNPCfRCICSizCQCNL
zxSzesaQYjy+pYeEFrSUpOfliOv6yf662CmfeDfj0CEuebKmR+uj08MjF3IazU8R
BYbakAwaA6kCrBUuIJhIp3RH+M54r6T5/L7jNxI8pidp/m9tJF9yAEJ2KCyzp70W
UbSL+vxKoQK0bIgattSg0B92st4QFJOOb7e48hc4XeWAyUMWefvj+CHk7RvY1SHM
OUTz3+Tp1eEYuS6cjXkQo+Fslgxgsuqq8Li6YvOOlXpH0eUEOs4qNUX8HOr4s0+T
/pYwdu//r/9NMLh5JqerT0m3LyapgjV73eo8A5535dUIcmexLZg4az5Ffx+6/4KX
FshieMb4afY5n0AFbyAfPpM/gzi7Iy7Rl1Wfel0nguQrgaEt/VJGlYCcAiqz4tu3
dYbQbHmSNplEJCVICOdHimMU459UlK94HiQGU2QgCZqoY+l9fvVABxLh2gwUjEul
UDx1H6/V4cM5wPcA/gN8IScCiS6wUezyIK5UkeXBm7RGuUQ/s5d2cqB5EAhf0wYv
aCCnepaF0b7LSkWowYnY29DnwhHt66ID+C3Me6lebTYcRIDR8Dfj5s5NTc2zz06d
d7pQzzdxLqFMDQ9vluRbyMnXiVZvhPs3iUSZkyh1ZYTihNj1KPIobqNZBdOROV6T
NYzNd3jORL0IJCO1Hf/mNo5CnieD0HBuljks/QdIhqVWjG5JtFayRT4+YG3Q+9Ph
QVdT/obZilnztoImoH4uYkFy/YEg9exJn41PtPdEi5Wnn51TqBzxSxGfl+RfrNVI
RjgAq9USZejA0eJ+F2OuiZi8/EnLRg6B6vTIi/amdJO7MshArpPavWI5tcdS8teS
YGi4htd57tboyHsTKGEmzc14Jn9UVmBe59+ldGRzIH45BDZ9wLue1gUeYU5w1i/U
pcyZlfhHB3IeZ0MUDxawxQejnj6A9vVl+4kEXGC6Kh6Ih3RbdXedHC5UDlEOxmH5
adE2wkuEZsjjmxaNeOAlN+WPNu0PIqQBoFgVZbopHak1kDYP6nrRboiFwaD6C9cS
/bK4aJhWW74rjbspMVpSyTHbe/UatoUvIN5UFbRfImIPaRTgDlUoleQVAB/+g88F
oJCRXWvOAk01plYjlrISasGpWSAWhJKQuJ2tURYC66RKMDx5x20ieF8KUqVLJinZ
mBgTf15sq8aLjomBy4Scn5P/NtnJHf7zF2EuH3mflApYoqJhvtTXeIEtur1TRw8K
eYGgyDnzHISVIHB/ebSnzKQXyyLRx/RG0iEpMDkGrtvSEmGMWdug0jfDXgYf2FxE
7290Rshrxh5D8Zv3LGA5PV/CeoRemNOEfIov+877A/h/1x4y5WfilYWE+kU72mlY
K81mQiuhph7O3ZmoWgrzpdRkISq0QuvyvD0DZoGTBE3a6Vb5CCMcB61pq9W+JGKw
sGslFzry2yMFHiOzOSY7ScrN+h0xYsisbcNTsir83qoNE7aYB8TS9fMqqzzZdFRT
Ud/U4pBY+yLTs5andxWoQWzOMv1FrQIvkhNkpKteeZPGBccaxByKRbtO3cmmffjb
5KWH10S3h7WP+XVvMARbZUUMdKWmTkp2itXbdRbT6G0py2W8NpquqcMuVC6eaXCW
02Lau9S3NjzcoYMTXOgMGnbbCGcUL3Prd9/yhboUOrRMx8soZi4DMqjlE6xyk3pQ
o1mW2+TQvuFOGViNzVebbW+A6rfbCrxh+PPEcucfE6PDE8F6xK8+JJ70RikRil0o
Ziptrwkio7RAIxNY4SraEg6DLw9xqX5gZbwSjoToggfDaVl/PaHQJlpwCikcxAk9
XWNcuCxXh2YeFY67ehzU1M68iy0fW0RPcJtR6kHlg4d8qI0Ru1fxhK7APtdkuEhj
Ll/P3lfjOZ8aTTHsgATmch6WfRpBxZUeTqgF9vD10zGXMF5DnHFg3Xzip2NpCubw
BVa5wRQ4AfjwPgV3umPROnyALnZOGdebxghZXtsnFnCBrlDNFb1qOhU4Qp02ju1x
BQcm996vfgsEEzh1jMyPm5QoZ3nACtYcrzGYx7qndMGDiV58xbymCiSkiQRoK0XB
FgrM5ZqnNSO8jHJm2POSpd/Q/JTdCu0XzGenbpJpDYwQuDhokggobaNurxRAGtY4
TGPJFxtmWo74QHWkNuqHTXGUTjsiApIvdFKw59mF+3YUH38keTKYcg3WzYi4E4fa
S7ib/MQJ/h7G7axTg9cpAQCL6un/gTNY4j7jHk46kpx5TUxz5wfBar0x74yDPnGB
S9E0pJI+sJyxpBBjdTRgdWMttx9F76sklaTwffTysIh5GVflGWImswR1DE7kBEBI
8G2MAywQ60JAs6nOkIyU2O9sYEY+FsST0wKTrgPOHBTp+sPHiSIwPuV9es74GN6Q
3kpcRt1sBUB8SsaqeeCnzNv0kn6mzzQsGbMwte5Y4eWc/1RKKJQ+8EsvwDfwKtwI
aXXrt1i8kx1+91XmToPJVq/zzyo9WGwhEhtanpJug7uaPLANywMFsDX+h/WnU598
UxdoaJ34peGFXQM4gUPS8iubylnXzM719qT3TQE2ZPD6NUuA7h7BqdFFDl3caJid
i2m7mxn1kQxxg8uWFliqmvUfFjtJVRBYS5rdGij9vsqSkUjRipamw/qfuWwHLqh3
TPUHBi/DLwd8lE8B+nRZXUjDOWJ7OGhgrTGaljTkgI6FMoavSGctnZKOsUGB8rN+
xuaRLukgneP+JcX8BONznQ3vDuYow2WCcy8w9Vr1LrCnwaMYh6jHa7c8VtvZeBmq
yyzN1tm6Pwv7NSLBb/u9d+WT04lfuLQ71WquMocw8lchVCfzNpiVSRJrGAYk/tEw
NPzgucbDnQ3u7sMiLVEcrNPEhoor+ArJ/iLpXwqV1T0+roIDV740RBOM2VoERgdB
d8TmAJG0kPZ34+UWdwN4vzHOm72zwzALSUn5wwfHH3gNOpcpjP+QPnBP9341gpWT
64adCshy0eSjIeP6nwnfmQ+KfZierb9WRqXrOOaGqTKMrRWchZDXf31HD2DQY61u
/igq8YMivDT4/mbT/JQioVmH62W1q3EIJkmX9WaVcHyXfJkuZKauvy4w24kr3q8Z
WDaRNWQHxPJldZuJXOA64W6fF237Hfeu12tNUFrpaz2oz59F78+ZGQ23QtWzGGcT
1Ypt5R9aZmw5CGTaHRCPhv+g6kLgmV3oNnaecibY893o1kRKPakyBFBPES9uUcV8
GtbYBBPaLFgT/qV4hiZdu5cvnqQO4FxmNPexvDELBlxKi4ni1D85rWRbuPaaBCz1
aAhNp82cm80BK0PLRvT/Q2VR66zg5MjWueBzNaipAJfUGCgNMzuZwSsE2uKvGtXB
RumKfc78hz4tM4otc5CMPU3C4iHkuoPcvbbt7JtBMoozR20Vxj3h3aeOZIZVRsPr
M7uUoG+MUwfW7zZbUcpr4V+qor0Qm+nmRSNAkJl7FbXTqLo2tRB/r0DIHAwxiDKZ
u/LsYbueJ02yxiAFLLQbRdY0o5Ebs+5lFOTH0r6H0bhPAU7TbTtcfIdXJ0k4ZWO9
1TnET0krWEp7QOY5wiumALlpAJmcyBRDXWPL6WQ9coBCd9Cfcxrv5CINhRSjBruj
WOkDZ6r7acQyf36iwK+MT50AJRs1HW6u13RL2B8Z3HAIL2/iyHD8Y1u3ZU9n7Ke4
pG22AdBWr8pcLOUc5y7Aya0mNi7UxKu/NrN7qQVkLKkIWfV8RvHiP91ilsgNCRtR
H78qJgsgSM5ki2sxigxVKGKC76mu9Ez9trew7s32GYieAZ4zyIczNIL+Lc2OF75u
VefEKc9k/691bVlT1L7SBsfX4qDQlosklNpr1oHefaOvfN4rOWetPwUXKrGEPSUo
1sjEIvBejAAAODPPUEULa4xTGhrmZEVurwueefE7BWO6mEs5lwLa57mYQtUwNgjd
HRgueGGlu3hnNagZjKIk/z7DKB9Zc6uwY1nlvUh5PPsTNYQLxVU/oUmTrnq2jOdQ
cjMPWZyPMoyBKNZNFQy6N/bAFkF/Fv8dSFl8INx8+qfazS3h8IcmayiKD04rEdOB
c+A6gysdE6BIgqnY1X79qddpwmCU7PUuq2fjH3dZcyH1auhfcj0Uum0OSxgwHCOp
Z+PiVI+RsT1AA9LLDBadFBP5BgtSiVkycz4kQyazrc9kD2nCOmA4rAhwRVags2uj
XQKqoMYwOu4eYJSsByUsIhChUpbAwFOnm7WDS1HsBw7qw0VTAZWqK6u9LtjcynEk
SzI9QAxv47Jhu6O31LhxiUUNhXU1LP3hS/iVHyGgfNUbOhnUdIdh7WB36j1h/fcb
xnrij4noByZsM5lJNj6m9APAzITC58PGxzBW22ceAXlcHDLa3mq2qOJYAOVgMXcl
UX+uT0XVABHD+SqJ5Sl76bnAZHBLc6FLOsITuJZcc85pWHl7V1FTf/VsmsWxThBF
XaVV99w08G6yRDjQM4hJtvvhos+xIgKFdaOqu0v5xbcLZM/JpSNBbuG12drD6hu/
kPcn0kk8CIi+6NUnRQn3CE3vGTzKfG70gz9NMCuplHTOpdZb+gLQpPh2VyVcNl9e
LRH4c9T5oHUYgRmjLoo+WxxEGliI1KjobXlEQx2VnbjXbeHzq0RPjBSzQMroHdRU
6C8JrmrFQCF7M6yFqzow2gjGvvyk5AqkvIZ52HjY95IG4CK3iuEfrY0vK3v+2HsT
biziAe4aInDKwvHkXCF7aVQ6NQzMiNF91W3RjjjTH8o0DqYHghcDrwx1oqAr4NC1
N3AR5LrQugBCOeo9qIQz0GoB9LeUmeIDTLYw/C2639aoyA4jJ4Bcj5lEo4e7/Zip
+Sx1ChLNY2uBPxT/hzmNP7R14As57D+dshbx+QaKjr8NdscsWRML40Qp45W8bGEf
t/zUXxCgaszKrztfB9r9SXOzxNscAp7aSlgLsxj5pVVJ17YcbfOt4WOPdIM5GbYc
JfMS6jmCVuKtq8SKFCSWY6QwtfYCNhrBApxIzHh0TBHUFcyzEB+QkHW7JgULTX1U
1Z6c5CTvOAB357zQoeOdnP9ynvBlW6/ewQnhJK76D5yJdhfxHANc8b/nRwy4zkAo
ep5pEEuysXWYvunrFwoKnn1L8JQi1K9/zNM7NMmRc9jzmeCo2oc6m5HgN4r0dFoT
fIBasK53WhLpj682lpXQAB+OxGQwm5yGmTuFQK5gZ1cjw6tyEol+60os07/zQa9p
6WGssBe3yFKiBlBDX+JGabbxaR1CHJ1WibYsyJ5UDogKZkOhwd2uPOycEedESw/G
tsn6cyg7BzEOTJ2GW27aHCSUeB+ruUUwzSmkQAvJNU5XQOSrvaDnrud97RsNec7g
qIMFB8VCKlQ/bDbtO6sQJpF6Xmzw7qKl3xf7xTp1bK7sUoorixY0CnCoufUZTP6A
l1H04dd8i0K/qyI4ZaedPJMNB9zar+/wsIxPJvI1QFwbxfMVWViXZzdwippWZPyk
uj/iTebrf7Y4Fb4hzXYiCbfIP+VevKfnONVauWexNgRV+yASb1gitWoFwl5ctk6i
UrI/vrTL7CQ2yXhWVuqPABWimQglUTYuYZ/DlBxKlWAlDLw+OyFYCgXfrfy/Juje
dM/30tDZhDe+Higj00Rk84zkfVGN9F/cDRV7W4AxN6cvRGdiqyU3F5l782sw8gxm
3pEerqeq9QQG2NNcbzCYic1DNCqs/7IVc3g9SHGQ9JOPbdVOkId/Qm4McFx8Oy2t
IK11MbCRZGfD55sF+/lk2jp6HNmW8J7UVdDsl49eGcwBnKSbE3WVqiA/wwLPXCJq
CJzRB9/uai70N1bdmgMRPKF8zoBYbghvztN+cVMraCMVasCU8xko7iOt6IxLJPHq
Qt+81kmy3VdlX6A/uWfmPuTpQZhChEWlhWfM/luoWqTSsyUBqQDweCuSZad494tu
pa/C0UYZCJHwc7CwxOqF5ttnYjTlBhvdlBgdAcxQHArnSjDivzIBr7Lclh7eyPIQ
tAeEfd1l3k/DQKY1kGdaBruQnjVk6/6cXZ1DoC9ECUkc+MisAIQgxQqj59Fe5Twa
o9VfrU77isfSpggdFkaMtdF5N9Wo3fm/FUkJvliAi83Sgm/XUFE6Pge4avCMUoaO
XPGDUu4ulee/68ZgEwTpp66H3lxtqqGSTcQZ97T9C/mfsFpd91fCCepPVRqI5sCk
u3hdS991SERzTQ4tErh4VIOg6W4XhVnO6WDSzUBO+90tHRV/PJHizFliKE7Wq6x7
b5kLw9VRmampw/NVRS33mUfe1jeyzWscwqatfz/JlAGRaV6osVSoMU89SNjzxPGN
4RLwI3rI4cWG2xPtCIJkwKL4xr8PvWjZjWrtniqLaQYrANzOQjh5ipClTqAlWzV/
1FsV8VtDhOq1pRCibc565YeDMINsRfKLnp08nMsgUi2u3HweBkpybJM4HIk8/PXZ
M622wFkjqQ8a5KIRk2cP/FPTJhUi8dBP7wQlToEJ4P5Ru0VOk7vbgDcsRrDUisFJ
a9byUdVCjCDP5/eyWKtpQikkCeYEEaMgzM5IZWU85z6XZN3lYUcGyuI5gNrqlWvp
tnjNxMIpuflS7cFQghbrVprpaFEIsLItiVprsN2Q7lhcxW9Hrh6fM4iZQzA3bmqb
kIRMZxIuf+rzY+xVGY7JM9wctivpubNhMazRvUFgaXOC8qA10hbgAW4rdh/G5RNg
E7XkX3A9A2cwENXNfGftdybrblvtK5W157na7q9TgQQ1smJ0Oawh8rp+eQDk702t
nUYm+fp4pjR7QNkMVta63B1l2OZEqcoILWdWe1/vg9u5CUPx7XtDzAk3bnrTM23w
4MmOLE9Jr+rhLp5A/G7wYp+VSVNc2Bb/cZE/WQwI4k0qjID/5sU/69w47ssafdYr
Ul0NSgc15EMnQm7mCHm2bV+5I8IxMRCzaGm+Qz3zsCQJIB2hprLvg/XmjUNyRuY3
aYrCqjWWcWhlH7fq6XY75rqSGch7J6q5LGrMd1X+SrfR9g7XBbXumaewyX9bSC05
elB9+KFm6rPQ7Z3XK3p+Qe5tY/dkBRd8s/wJdB9uBOpA+ijsFuwjvuhTjEZBlMoq
yLfNAYL6cEdoLYVX61uJs7UG+yyoYAbrmXWrw6npa7kUvVRVSJx54qsLgWwQqY0C
9BVBDA+gA8zcvo60ece5vI8yxPHXlRnAluVyR9Rbu4VFANzSFVXHsWCUWX/kQHO7
ssbNy6YQnkGriVp9xNJCKwDKcQzruAacOvhNEV7RfAKI5vXAxu0Kz+pC8KxQn5SM
Ej1gnf8CZHmNVYY6CHNF+4/gkxQ2mBSwmSfJXswL3F9JlnufnrodP6TCtoUswHUi
YAuywjLd6CN5iZJsoUXym1n+jBhD/GXbRv2OTebHRMq9Py1nCm5BB3BNilvi4IMk
a69uNTv40pyb65Ql3CLZCail/QhZJusUb7K67pvd9RmIdYaEteKLiMvC3Ylc6pgd
yQK/pRe3y1hBukcJw12+OXHRaGix2miAueFXzqXp2Tt1ZkIrb58H8nGfzYuN6wrg
ZakbRiZqQUpyESu2DGqcj70Q5U93dZJ31XNow5aYk551lJUX3WbnKuCBFNCpcJVH
Ij2JDVGACclcpPvD/7nAU/jCWSltbpLfn0wJ6emZuShAtjDqGXTpP+W/stWPHkV5
DYQ4178RAZ9rsL2WbSuVlEWHnzom5DFmBB7ib1j+RooW0TlxIQXPeJt5nhYoiWKH
ANSHxJeYUfIe3H1BTvseqhLjKxB94DZoJMmTOiOfDsaKDbBJ87mqrbyLpoh/wW77
agoOgs8fqa9nQNJ2yYFdhxnUCIlVuV0AbQtOnK79YqA8+wdBjimsm516KNjw+aWE
KA/x/X6ZlHie5gU3QlQ83yHStYnFpvyTOi7oTVQQj+Tim1dDffYUpFWkj7j+tpal
FpErwVzD0EyZhYbntx6XCv1DSd/wg5uZr1Fy1obO3x1L2mORx5khI+sPdA/Cd/Z7
PmpIG91hw5ht0hXrY0dGvSr3QzMcuiZdHDIo1UwMbQHnrN/Uw+YhYbza+OOFJgOq
BSUCIle8/SS5GwyTErgeOh/rGupwi6sH78W3faPL3b2d6BYwpmui/RYwu6vsNzO4
v2J1GUAmjcdFx+5IRTnH59shRt12eAqn9/A677Qb5NbHsATlov2BDPL78z00hzUO
c46N8pZiko5UhLNF7EErS0Srd254IhZBV0bf+7oBiUclHyZB5XUHhHt3FHg0xOYT
q8x5WUUHvj23hKUmlgoYMZoIxBDZJnPRjLeBfpnR8CgpOD5+7eN9kyTmHNxyiGuS
+sNA3f6V5NIrqRPjpTAuVRltlRiyKbqiCd5WTK5fEawCVM5Xyv0xdS0eQS6UuIXo
Au1Wav1JATpriX8AMWWh8WK91fJwyNjwXw7hEPpRAbvd+ZpCtRaIgx634LGX37Hx
zwJd4HVZkLDPfP3/mCYFI9u2ie7qBw81r6noFA3o+axmLQxvUG3BdXCqBnEETM06
qnTDJF7vNYinCctaXTIHFlKXTAaXyWYqmWy4WHWi8tUQufNru2ssOqkowsZZf9bF
JaagJRVkPCK9r5epsSUQo2OaxJQexpKYqz7hYYxNivErfMFy0UV2SleezPca8HaM
KG2BeM8uTgPg5xw056ZQk26SdWbd9n2QfGlBGjVLy0nk1PEHG9jJvDSvV2x+LF5e
UocAuR9ldfCkxaYqi3ni5bo2k0R/3MMTKN9VIO4Xr/XLbVfAmA1SFg+GZ+Khq/IZ
/7mVD14hxWczhjpDX4U/oucIqfXnn4hMektMObM7LBFuj/hisDIl4LD2rKnSYipA
iZcriY9N3dtQEhXeQHouZb0a7VU2oUFeQLSOgZOTQ9u+bQ4HDgHdBKDAW/8EenAG
IxoJXDTXpNRSsDzA/pdi9nGGtAE2ag7amBaM2dcm+BTWOr2Z3f5EhjaHFKer+PGf
UxiahtOelDODxOpmg/G0BAnNz6mw/0B7LwGZwyEjE+gOXHWgIpwPCGT1x6XWsb6G
MbeeZYm4EK1xUKzOvy/UUgbdilDhmYhLbWKycrQS5u6gMiylMa68cg0zEewZ2u5c
q45s4B/iLr5RArZBrw9d3bE1kLzvoeyJntMzmktU5aX9wMq65TntxW+4GO++d83B
/BsuiXaHwZ0U9EElOyYclJduOlzaBdV8R7fANKxdvzHa0Plfp2SZ0XiBWPk+qwJx
OUANL+y6SZ9Tn1APd6CLKd4/PTJYay0htgHoKWvlgGojdglEw4bFHZDMSFm/0B9Q
vmeOZNdSGukLeJGV6TBmqA5ZdYoRfWdJbFskf1p60uAM1aKwCfD0KIDi3H6slFCh
5UES7tMehp/efx8POABpqSthcOTffJG4cQVQLH5VL1O01IrC6SUBcAQEkLYKx9Qo
FgYDwG2Uqn/oPm7WJZxjtI9SPYu7etjYVsffxvSYobE649OhzeunFbZO5s3ZWWGT
xdpIkgeaUrb07jDkfsnUHtok0tymDdyEdTZZ28MsvZDhThcCW0om+bfy+xQ6ovEw
9+67lCGvWA35iSU/71zWfjwITLYhlxkkVenpmCMfvQwYcWvzqUkxkMGBcji+Ijpv
t64VFizRTAUbQyEmB1eVFLCt1kptQ1Jj+sAS+apTzVa7LdXwjh0aKifqEFSBG7BB
G4+2YE5Kyp3dVG5Z89n4VXNXcCgssCK+qzQD9wIF9z7XMpWrTSO5i65Oe/uEWonM
ar8jDNgsLpI1q4FYn32Q96kBhBElH0rqV+GzKPy7z3pb+YuhFLNuoXvbmPjlUMHV
+TBZHkpbbAMKT9PCGJcnpFiwRFB4D88yIaRx6U+ybtI4C6ouRkxicPLSMSk2HaWd
3qIcbO4aDAjJVGY0P0j8eCOprynv79PdPD45+1yGaKYsnbfRaGsUkWMqAkjCTPQA
zeAdfQ+wE4ukMyvp469DfzVNnI0ekn4sC2X5REdYceZVzbBtE+631iuZwZWC48Ac
RUI2eZKPSoVpVSHzkR6XULiOgaudMl8dAPx2bM7BHQoN2/6VYMvZNqTTx7vatGyc
GktTLEnyaolTpRPbXLY+3zVbpasJCNGUFGTJ/kfHbtCu/9tK7+T6O1O8U0s7efRr
JvD3QXCy/JJEY8/Sq7xxY7S1jVb6sdyZZjTBZtmTH27QdFDcmZblqPZu/WMH5OZL
0GlCAQBIuxlBdaK5e2oc32RxsetAoIzkRA47EcCJqxVAtsXKvRnM11ZrcgcMTS1l
8uCs1oEOwwZ6SfitJj/853DhEFYx2GlyYIBDub+tZyiBVnXn1x60QklBPHuGls2M
CcYrVCNoL8U4WU4+LoxdLm+9hh4qy2ixaX+1QxkDK9bOuB6XBkKi6QsZqpBo+zkk
3mLSetfedhQtu9ooZUL+Msc4ILgamBUh1us5gsvFOC6Dbj7xtGveziZBhGEyi2ja
yAgpxfgTnJFD1GIVk7gQx3CMH8mAqbFf5tYAnJrkxmins5HQLwTC0zGcg7HHqqqC
X4yu6wNaTvSo+4v04Cl5THsNWHDfjlkkQgG+ZMnh0yToi9a5gM9TKFCBEao1wmF9
FRHRa1smR6ha852Xll1gpKAKN6KpKKEu0WnlpYHA9+kYlkTB6Pz3ihWTMHCV21vI
nxaiY/zabmTtPLa6lY7+2qAdqXXaz30xOMdrbmiKF5AJpOV7/jJSzKA7tn3SS/fi
nrJiJwT+U3Bd3zo/2dgJGDobKD7r0XiEOt1UlXmjb1dsVZLin2G8zB7wJTT8GKJm
K0TCVP7bh07junLfj9qCkSqM/1QfSZyez6ZeolrhPSD3WIjB87XsP2TbkfX45jPZ
Wzj45oR7VJBr5hXeUXAhPFDggvm6Qf9VjDrYEtWlj9+jK3zNuDqukX/h0qljM7ZA
LHDKpWRS3mKpV7U+R2rrC02aEquKFWZlIlnR+rm05zRfGkf86xXN7X+fOmdCdIyv
mWilvT3mi6eJy2DDG1Ozc+bZJdY4DvULPavPBDeGUhdT6VrGrdgwGy5F+m4jTviO
5UqdDXxxVPS4w5t45cL0uk6NW5BA6s7QoyLUENM40jfJovCxzf2ALQpAzKqGNFKL
pM1CjxAl3zbfAlOPHgUp+d1vQB/oi28+L/gMps/3rj8To2PsFAcp0WN4oxAlPwvl
NGF/K7UedMGSknXauQkbzl9Fn9WuQJ4BdIM7bFSy/MPYgX3OsUR7QbuYEAboLwUj
LJFWiYfPeOuE245Dmq9Eq/7ye+EsCyxo+UCLezXdLNoXjBlu6FbFYTY+54XdthV/
5fXKbWV6XZv4TQJ7qk3EWV2XeetY9bnuBWqsF2BCXkh1s79uqnXgfo/cAeZlD8+p
BOZe8/rRao1TAuOvu1tUdF/NgVukVOf42pnC7NCE9VWCqnffDpRKyuvau7UXmVxC
gP5c/iRlr++GMTBDw60jEwdooNVQJwgvLWQihrUWMiFz6OcVx0ER0e0dLmKfGxBp
kBZS0BSk8QLz7j+4eB8LHEVp6buV7tl5EWhREyvMcYp83Ao0ksUPjEnpOTitudhG
cgq24oZ6GWQBnUwHVYNnwn2Elqh42cM90GHwEC/qteLbxAvnCI2zParb355Nwk37
jzSqrU9fXlislVKa8J6jUL9SC4nf1UfjmlY2TPkTyjfVQMBd0s8cSFgRZVj3qp/6
xoYtpARm9qlnPQIb0cpUNbO5b5IUFPoC7w7FIKu6fhGOc5j+7VcEmztgmtFBujwP
pXmx5val0mpBVUL6E8aI+2c/tqI3VRTqv3x50rivb5aWqqqGm1AfrNv7Zw6Iq/8p
1lbQlOHr4zuo4I74HESBkdSoMw60ciHR5Vv+EQfkg01iaPTyWMIfbEYPwiXn7azb
MYOEF4o/A6obXsx3GvhAf+uqlGXwWqrbdIgoBE950KlPvh2bCh76i7eorFRGk6Xy
Cu5GVmEY1AdWdVt0Pxj5iS7ljLcCVwxAxEM+wnQv4CdAsH79xoV554xZDOM2s2N4
J5U2MXIBH3Pbzmr48DU9c4rr62V5kqqVEZ+r925p3oggMkMCQ6kTuPEiCc+GZUXw
p1vp8b1uAB84X+2zjTLeJzpCmwy20m+myJBAKI8i3wTf1F5D4TQmx13z679XO3N+
ZdKKa0O32uwJ4OzN2jerGL6bI5T3U2lsTw7B776C74XAfaKyMSE2uE5BklwWPcqd
rEHiSqF/ti1KshJjbcCl+psgqpIQgCXlti4hO7WoO7ho0c37rbVNZvSWvIkyTSgl
qz2NkMF0GdH9CXT9WbHFGWcv3VaF4Pu36iAxw+OqGNf2YKrkkI+/L1OwGkUUYb0o
lwfCbtObqkCGd5m6YDY22Q5uPPq4do3ZadQRQelbFSBLRdjYB90MuNeeGEDb9fY+
d5MIxyy2rp0NgyOrkYfxfa3igffpmBZbhKiM0ddN03GSg7RE74uZ8uGWXX/r4GHv
yIux4ImhxGG8e8vvmVZ6I12xv/wtbQkm1gGvS3DxaVpq99XbvrbswjvmucOLn6TQ
9qHv579a4HT2IVjS6Z/KR62HKrBuWaQXgRBXoVMIdx8zao//WFYQ+zJ+oghLk9u2
aYHJyNbFkp+OB16tadxZmDpjxegGfGQ+FIN+/vfVAAOEcHerPrSFHv4c+PLsw/YI
bQhg2rWjNw69bI3P0zAha8fFkPFP8BJX4idXrqwcB5xFfpPwF9Tb9Hn/q7UTys5d
xw2fD+0C3vErNghiWuXcAHFou/Hajmsax+wqumwjR/wscitnnRkGhKdo9Vl9duU0
uUmGLyz8DCVhY05Ptz9VMNrUdQEAblqbOBbA8RfX0S2wkQNHDqDtdy9trjn0EtCo
ADYu2l6urMXKqiZMejgYu96o4WsFJqoDxfX9JW+/4hoL/vRgoAYnC7Ity3AtZ+A1
odCs3Bdh17L35QVH2oBipWWH3EgZgHUKkPgyxDlyMgUn2JpeDO4LJdzciUTwmbpU
Tf3yRMoTJfXv+D48WOO4aPOqUBrr5MCkK+XkccDmLQlm2IMWDV5O+PNs150vmJbI
MpCY//5d8O9m9WfcyHhj2gKkwDcI3/9dWmIS8Jhwpp9xaX6Rn8rMRsRbKZoxlWLY
NYtxmj+aqM+d35Bbz2UUq9vHDJYhx+YsEyySAT+EhjedI4p6reF7rOhOgE4pfBn4
I3GSHCLFQBLz8tHGu8fENbSwO5pVtuyMNNtI+n2EoEYu1CVExCzk2HGBaJQmf714
UVjcmtmrGUED3k+AW0wpNNUdvcguv6konnA7E60pe815JbVGgcGat6/v3rzeUlWp
+Lbc4prEUjtuHikWXYpr5G6FJSv/PXX4Ef1jOx7Do7MP5y4/JSeO231vOGYZ/4j9
JvXArj1Nqdz2HVuBy1pLlnNcX8dofzE8GAXCrOo44ObsOEbRZDcPVevXrcCJ/gxw
+bZ6purSFd5hqokdJnxzfUXiqJDRyzXKSdwcNmg2vDjOsc9N8Veu0xYc2ixYgT6y
uGYX0byjsygGFN91tPZl9mBzx6JpWwXOIyx3ogjKNglclzRCVjCddFnLjnFml8Vu
OgZzUVDVC0PZQfuMBukP+oL2H7oyyTTFOdHCRWSlPCJQKI5afqRBvJBzpkKsp2tc
OTZyKSdzABcFp8cU/aqA3eArBQgT9nOus12lUmlZUy1TtRWPiuylF39DBePIuXBy
GDrZiUGWkoJFRjKyh1xTdy+dmWC7yAvXsUWc0x5mQY4lQHlgfljHZ8+Lu9A7lXwU
q/HfIqC3uwM9xD9Y2GHU0L9q+b3DBuNDbo9NazRGNVgzO9C9msKSyJlW+72DgQXv
mjdpipUp0jRFj8/ibFSX8rCrDjfenvb4s7528dUMcpLQheIsfQH5XXwyJ600++Fb
3ximG3ppJKVo2EwoflYGpQiI1wAWry7Wvc48cy9XEJ8sGHIOQzySE3P52hO/jJa/
AJV7DF2yAyzLIZ3+J+LACHsaYBu41/RWyMSIdlvPNKZWoDkPsX3npiWFUcnCQT61
CWLrclEUAz3X9OtCXkV0Lib65oK74pOa8d6wuQoFhfkzIxAXEigYC7axcHwAw8c7
0BCJ7HplQq6arspwVBdtouS+h1+cbHUKXeMctUKQc9k0jEOaNH18lh3EZdx663rN
AM7O0jlzyBBRNOX8/MsfX8cGnxw6QIAITsbGvdHKXWaZ38VXxo18VkBHYLgdldSc
hu05L0fpIkmVnsQR13WKIqYIrUHNPxZvxuB/w5/MXIZbxuEwf/flodsXaXZ6ZcDI
22n7VqXcUMZpI8bVtjpcorwmB6tZHdm0LVX/8zvzNUAthawwHum6UYvQ+Xar++fN
8K/DFHD+3YkclGAtHIxD6RKvmKlwiF56KnvMX+KZJ0OLNZz2iU+Yc7idlQ3Pc7Xp
U7WAfyfD3yPJ3yBPGxSgcWHDVuWGEpZSQqGZIQZAuPTM4RS0MxXoEXdUavn8FRSP
gVRnFTNro1RK+AIsss9a50MFOd5+W5IK6mJ9IJQ1v3hhJHgrYAu1yzI8eVcO1TSh
VaoHYRyIANmBQxWOpnQdKEiwOk6DE3eeYD9BhsoRr51LC0dV5nOK6hPkiWpoxeBg
n8XxRMsfqgZFKFAvAHjyqiADeOU1oIzPzgPJ/OpkCU1yz5/5f1HS1v91D24gpXzG
5hVxL40jjs/GcwIgsi9Wb/FpeCDWjctNWBrNlL6InfeYddQWoOoSERynzujhZvpF
Ly1CTB3wdhj6n6eLpavbYemuTtIYoNBde4kLwxgAvaNi8cot3wU2l0GyOLH58gKH
yrZNlizp8NsTHja4Q7cTTa6NKaAk57aFHVpiEJDfRlvK5npQpj5H8JvXWwXUpEOG
wtI8IF2ReLEXsIVHzqPN7OFZJzCQCxERqliYs/z7m0XehMXWSCzJUflFPfzxYyqn
24ccvcatpw9C8ljf5oizAOmQ4kFPhUstcQBvBuW0MWXxDMIDt8l5w+nkuI3NsVCO
B3W/Jvfd3sWp6R7AeI8PrktENpiWry+iKrpzHUs2VjzHsU6Nt9H44G4s/9xp/lOq
TdzlQbVd6yzR/PDYO0RA3Ce5Cat5r9y7UByuGpufiYPZrLPoEAksrnxZNhIJSAmS
nLEbix72+m5yVN/RoF7o4s9MjCBYa2yLAErW8Jr0GM2OZolpTPEtrDzOWl1hdgBw
rUl0JtTe/adjrn26qIVgfuhOTClHTZVbzsTQcdwA6GKyE2+/rfpVVs0y7acrmCix
YZzwukxtOg13c8JGL4A/MK1y8hTQOIpX8xQJe8v1wZBYzlBq4vmaofIjiuJf+4Kq
2zD4G5PDHq0kxoXHhLRE85YaG7dW43fujNb8wcVHtj1wIrTg6duYF1OlUQ+lCFBU
Q2uvzr4/GNNA5NTYvU9l1zfZZqhfqUR4RIzxQP/aA+OZH1BUcIL+RB2oMdCNxYNQ
Md3RA2fTuoRjlf0g5j0KW/qFXHOFw+D/opQ+5sD3zvI+oMmwwTkQc0HsmF1BQpop
825HCqOvcD5suT3Oo4xjKbsAvaPd9NY1M2kU5UEktS06piNJhLBF67fCzkTK2n4G
MkoBMdxIRbzMnhvRQY19bW/vkVyAGDFOww2FOWGn1drjlIgVnws06As0AFWOX4H6
UriDnvHHe1PxoPwUXPgIzv6VIDCSHBDb+JBjgqDj9nRhP91jPW8oHEiUM6S1e5kq
0oETzV0TckM/hhSaDNej3pUWMO9SKgA1k8yngyeWSjnW9q74h/4OnMh4DoH0FxiQ
fJSfBnMhG1feoQRDsllrabAqdCIQdNyKfE4/eI2rC11OCEBetObk+j61WZf3ELmx
Os2TEWHxitTFF3uTCqq1xTWnbA8PsBhFkDZkvxXTtfAnIq6PicEhYdtEdUOnc9tm
m8SV+teTEyxX6uDiGpgWLoINlUaB70Q6n7016TzMXMUwXO0HZBWw8Tcbz9wa1qS2
S+2dyShSnESwVRvJ2gb0h1S7jHx6L88lHM+WntroKmr7M/tnAszwLRuICDzOVecq
AUx3ywKoHGW7kIISVSLG/uVNon8xOFzU93YMAkPu4SbqiHVtiAIZ1y1YaQyUHLza
P42OajcQrPJfpjkoqAoiPDs0uWe19pZvilBL9gVGfKf43dPDHWbOnzIUGZLr3xzG
X2XPLWy02RKzTUhpT01JYLmoRuWhP5yj197/4SALF1n7fFiN06K1MZZ/Z2bRyGFY
ytY/HtpPmW240szR3CLGbfF9aMxrWcqoK+h/qXgOoALz+X2rF/8JtoTHsIqRZGLf
Moaa3VEyVO6ehPo730bCv/WQZyZLqAGQT90Xxn+uDa7fUiCeiWBAbrYCVLui6V+D
IDQZ0YR7Rwxz8TSBFUbNZ9n3ert9BdYNoF9gunNpLzQIkmEzMeMqxoDxdBW6wopI
tBXfFMXDURmvVFffgtRuIdC9AaR3oHvAWbeo1lYA4stiQg1TK5uW/QhIgDzVc5Lr
ePj9GekrrXLUdeQdlAXDgwMu+RypZ9IijFmJ8CvyTf4hB0UxV82XusiHQyBzyyZj
r1FG+NrOoLhx3ikCw6eiVo6wj9N05Aa25545sUzEEJTPcKPUnI2sA7etGUezwYkE
NEUaszJmIzo3RYeoiRiIv7hL3J6PLhhPPVOImDBQhG2jvIbvsIvJ0Os157KbswEm
fdeoR5msns+g4spgFclWLGhSy9mtkQXDM1Ksi52YHXYiGvTE3q1bkvy3MW6sPX7A
1rGdErTCS2t/UnnkM5xWlXTCl0wYQniA3H+YkyKn3geGVpaen8vrrslKIaGEty6z
Ey4JY9EGp/NcPTXS1TSn49jFz/94TV/Cx5XpncY70go3st1QDiTf24mBcvGu5qW3
MfLC43W7LfjnHBMTLv9IX5t9VQXVtkNKZTez9o9grmBjppNjnrKpgelJzwSGRUEd
BI7S5+NuAgOnzTB4RJdIG4qJq0ohjsjz5VFShwDMxCWqXjK3Ed7OB0va2gobi5h/
iT49zjTdu07tqBi1l+OiNQgrbuE37/+0PmFyP+6aMAg2HbCe41VrhiD5BGYea+Qn
1mRnGda9OrtW2QVq+k2/Nk17LO+gyeZO58OB33KSxNKMyD9KqhDsmpAc0aydZ56n
pZ+EbcpWVNxTWPi9qUTLGhl+Gt7ksf04I8gG3SKY9URU2SEwgJPaDsR39mVydB+S
FQl9TBCCR0yLipCqjQJn7vRE+Uije1VsILI2bLdnI7H7/Bxs3fJS9VUs2nli0GY0
msqIQeVcEj4VE6SwmgkulwtuiAMXCpeMzg/KON87nT8L+jckT1DPbQcPbNrO2RNC
ifjezK+0dkSlNWC5Qnx5qoWpCE79JwwGiqvAZQKFfqxUVFifu5K7HXxkHcNjBZK6
gKrWbd5NbOR0ZWuwT+h9JLqFUFQaviMbacYPY4E59aStX54UIKpYSZdqugu9mgXl
uTTU3hn+ZDA/6LmVTJNRFQFvCtjWADBxGsewmB/RyQoAzBB4R1qYKtn9/ZAzQ788
DM53a/ZJ8ACOeXBv51qiFQ9jOIuqn/oMjyHf+th/clluWQfHB51wbIzlCj6gKOdW
q+iObjWdUddmk73gaEk0e24M/NXIbvLZLmpDiN5TUU4ubn/uZ/xVekL+GfVm3CDx
JwmlK+g5yGwnntAP9ukK8NakXN6fezgxPSzCYeWMjaqS+4XAS42vzcZxtVgJwYIZ
/hbEFgOu6SdB4HprGyBiu1++M/ZwLm6HmLdXFHjUqxsmdAyIFxnqB+C4mPKAJVi4
lUGD1HVqJDtMI3E/UTwZDB6dXtJwdmArK2bsNxtiZftRZ603kKAiI1S/t48aznqT
F/rkP2w4UXevmrzFGwbgToigtluGgxgZLWGHKFB06LubvgSceQDbzOYKa6P4G3HN
A6EIrA7JnGCkcctPQhQhmv38htbyTBngUV3ZFufUja4WFPg0C/r9ZLMYG+RO39mz
YjD7Xfkf38/xaA1TwS/bGAhiMzHgdlXPybNZD4ljchNTU+6AAW2oJTXWqBQ5BDk9
Sd1G9P7KAt4LwmT4sFPkR38YhUK+lU09LJhf6UgDvFRbNf5Lds1VuBhOn+jwrHkR
mpH1bU7BkZHjlg32GORLD1x4Ds0FbME6d4yjHoJDYo9q/MfJ9BoKsb3w0PB39XXn
3LsBBodzCNAafmFICt4FmJLy68/3ztGpFTouVOTQUeVEvBeQEiVYr47Jeebdg0dq
XozrjMATQlfjfX76560qKzS/IQzHqpPhaMWWJHVeUcLTaEXEjuMUq1+/TXjP3xA4
3b3hvWSl6qwsxS92ovmn+USvxo6J6e7vXXago/NhD8nMiLLUxMKOvPn8G4QZ1jml
ddSeWMkKl09102j7XeF+6fKc8lDqi0mBgwX6zECzJU7/wXt5fZCff+0u8qKdPLFA
Hl8zchzHfVw+ZbkfLDlI7JPaTSD+DX9MIw/5bKKHsMbb6A4skluq8GTQ0iGMDjWE
GICHkt0k3/k6Pn+mP2vYDMbaZka8EldH3ZlaT1ri/5hfQ+Dad/jqMSgersClG+Yd
gulkPOEZrm44drYIeWKPDV1BmfUnevJFzbAEtlwAUjaHy6ut5/uoVwnrVHtA2GWw
CGVGQH1o4Zje3vMoMK+Btn3nWOz80h47W2i/LgFURf6kwndOQT12ZuIziwFSqjAx
Q8vw+wFvTHUz5q3O9PV73JimP9G9nto+Swe7CoAkLdVi3FjrrlVb+PtFXdpSZ568
zJAK2SfRKSKyCBGnPSMWvunmjmcMPxkODqJaawR/1lp1iABNb3mOKgeAGVqlOS0R
6NxIbJVEvEjF9mqvSFVDY5xYW5aUCCl2PT8YHDIJedAF7ddO06p+KbYqOVLlcgyc
aja/UordT90PD+DjmQRZ2uNV+oNXvEvO9uDNUp9/qyFcPPzhumriTwYRH/ydDD9V
Hgr/WPdFcLcGoNfuJxhIMmEe9PKAE+gheKJC4RTMmxntMGGs4ZZ9FmyqyJkRAOoi
h5mDkQhGXeydmVpVL5AThjzkWfwvUgHSwcHSDwEbUUyWvEuB3LCpNrzDmW7n5Pb6
QCTMgTY/qF7Ix/YAxqaowKlDC7gbMxUU8yl52hksU+UYrXF+dylhepitUS/LNGfg
9o2AaXxffCHxmwVryttUJhMCTCAuW1FRgdjVmvX71vbW1/5pQTqMlGGiVNqBy48g
7881nwc6YGokJJDh1jpIKL/0GI0qkOMHVIbYTghyIeBC3hHQ35MQQDDLF9VVsY9Q
bzIYFlv/X5LnR+RETlfCjXBt3Bw6gkpO7IsuZ7uLmPpTQeN8OmWlMsIQStfp7Epl
zU5XkVCOa7HDY6YBcdGAJhMT7jqGQIcGJuVgF00URwxqMVNlub13oxC0UXMqYo+r
63rWpwXALPzyVe4wZEFufQZFo/UmQ+HZy5XdNpBynJCqsWoy5gUhl2u024oh5579
wWNhEjxemozceff8d3YdlhcYL5uVAUNRXp34wM4jswkwRyrsQIozAhV8LWd2JiMj
tBAW3NM2jNEG2N37eb0xZL4jtC0tfBqmtJNFibIRW5grt8AETz05A2Zgt6YCAJ6C
+IO3RvjD36RveZXiTSp+4jN0rWBFBHgKL/A9VugqEfD/u5EW1lBajhFY/7gwJSAQ
m1u0ATMpBvActnSuqCNzWhqNNQC+OHD96Xpc+P/vMRqX8iZLX7RhPzV1jiZUHTGp
4xQPJ89lxfPTJvLgikdSw7ipe379EHuGJMZDtZZtgShYMzo2dqa2xN/9duHZ7Hmd
Vjxwj4xXJI35bb8b0sQOSEsINTLJP8vpMnQDGDM6Lc7XF+q1cBScZ5g5EzDLZfRx
ar3OhVg6LjuXOrMHNk+DE4xLcoLMXBsRveC40c7uAcFIAR5VGBrAQoBwhWvzogkS
/7MzWUhgq5oumjBeYwqVia9PWhhEyORkQo4+Yg1y0nJHoYYNMaqurR6IUzB5LQJ3
lrGUZa2qOMI/nPZl/k1YqZNIQ5wcux7nbPqt7kyuAf9eN35ONfK7VkNOyvmEbeLu
KjEqp3yqjLspqTb7pLuDFsJet0qYmM72eOgNza+FvZsaBkkhCm2rFZ9AU+E+rKCk
iqa4U68HuuCb3UegpUe+VM7IzisxptgIuW+AaLeCYN+KGJvjxmlq7csxlppeLaep
5ft1AAIk5SrhuF3BY15l+MbXTbhRh3Ft1rS4hYi3VfvYuxGmS2bdgsRI1sSyuF59
bx5g5XpC/fOU7KxE9GfHrdsa2qXca0miB3DJMuitlJkDUMmVwDeR9QnR3hWZiqQG
MwSwzdg3ZXtAAyex1db7Y5+J58MshoDddDbax1ScMJjT6Uw6ISJqIwG+jv1AMSHO
wDVVYOxlGNItLvDIORfqDg/klMsH6w9jrnwGSS/aqOU4LjMe1Q4uewyu/1qqtf+v
zzcdceYhBlw3qNKAcnxugqKIab2fOBl0E/M9LxqLo4QIszTv/hlkXp+NhUJ+ASg7
5JPVwMhD5nSC2v9nHq/1x42GWfqeNmxZ1DmoNH54NOKpyvXml4L3upVLUCKfHkaN
NP9+ZSro5smfpqRkDpJRwKGOOnd2UZbBvQLfT4LhddSgMvFe84SIYxzxYIkgLPNv
5rLd9S/m8wzK9/Eiro7/UZzhkJ9YkRi8c4GyPZ/DmNwihmH0p3K/sS6Uq2+y0E+E
0RVhtDxVI64qcOo+j8N1uCEHPXNPHjOpoAYCqrSfyguiawb3uX5Toc9oFRS1jJ+D
XF7vuIyrxgr8jZ9EAs8JbQ/TxIaL0f+t+Wsxw0G6xmgBM90qw3z+273wmqHusg+B
RQAVzPA/BhPgkThasCGVoEdxu0VfG2Awe5Xg2lUmkjUxHjuemVaRXtdbKIPAiAy2
nt4wuHkaqi1isagX9rI1hEY4DJ3JrYDgxoJySqBUJl0SzEnUTEpiOe00Pm0zw58A
0Hp4HSjDHXJ6mTDeN9VWAPSqJGrzjJUkub2EqdvNcgadW2+4FQsCfnR0+tbzFUE7
aqIKjiNUeyzavmWl74vKkB0xju/MBPvPZk0ziBCql1Q2HREkWPKyo3BLj4NKUiK0
Qc5u+o8W8x0iRpUamZzesjSRgV7t/3RP3CSPWZrKrriWAmwZ1zulfOTh9MJEo+OQ
R0cePCEVfz29mFUWdCYVocNv2XAwDJfWmZwtzPkOOTfNCinbuUozRURDOIPfm/FH
5uUPWYfwSzOKKUz/QYie03XhGV4gpGkLnFkUd9xhrxUXE99rvq383Tb5OoRxI/OM
pJtlrmhZAQzPXj3kK+L8VXGtJXL+kzjJ57LEyXdjzH5rJ1stRQ25dkn5uRWpzg8U
TVf/B1+JS3lnwR5xc3Vq2Jk4NfqHZVJYJsJV8EsswsvcXL31XIfVUlqdnCHuwGDF
ZiRNsPx+DkAtP6Yvnyh3ZwZpNeu10Hm/798tqxP4GkwCEZu2oB+RdJR0FTW1noaZ
BIYSecFYrLPU1lOPk99uPHQ8U/9uDh+1Fvg5sJr8rmUpeSAq/WHbGgDy61XpLzoS
2sqPhGProMnRRKnk0ujS80ei4ccAb7DdrxvdNj69qCp31dReYrPMiVwSZQ9e2+zk
M6L5Wu3MOIHhp2gLKwjbja1GQHTex31kbS03A5MyjUiKJjmnBJXMbJ3vdXDDtKo4
BrsMolSLIdbqdNvDrEsf3mAIvh+WyvmT1kZwvyEEYbEWIU9Y2x28op5vkLEiTisT
RCFNQiIYYVzeV7iHyLmEcziTuBwsnE5rXnybGBIhIC31EHgVoOcLEtVFaqT8Z4B5
MTSaBBIHBMSxlnNPWNG2hxT5VGBJOeGCQTa2ZNceofns6w67XYZn0mVvr6eyjF9i
DV/OnGy+2YFECXmyApSP+cKl9ky4zfmXwne/Zhz1i3Mkz3eiecNzniR4Tu29MjLy
2ZZiELlCqxzW7N9GYFst1qMJAy/ev4VuG56yls+RBjE2EQn9sf/0uBBtYERXaGIl
84apEqXBYVH7Mkl/jLaS33zwbXEVnAfU0V6WzFk2bpJiCvp6beHXRt+h9Cqu85+i
lrxKgzQAQKkg9C5V5CNL2lRYXRkJ5BZqa5zLndOcQITscfyXpIQWGE0nxOimK4nL
cAQT1TsWjwiAl2l82Ompgv13l+t6mJYgKUsD++aHXzbdwEd3lPXSa11iBaFXx9Xf
AP6zuF/ZzLnov15FIL+RKFMMQP7OqN4hZOg6dmND0+IBQQqEIvgfa9UKwFAaafjM
AdmBZsmwX7AyrI1+Si0GA8OIwz0gtf+1CfIK4FWSv9qjYd0UTQHALfzl2dwxKw+n
CaJy5+pi9PNLTbhqv2Z9qay5aBP6Y/K+8ciTw1q18455zfwgtbIKihurJtA+C7D8
nZMg2aZyGc0ejJV8+Jjhu5HmWhW7u+jGv2a3j42YpcUke1k4AKGEmOeU9c0w+gvR
NgpdL8axwRn8BoawDGrMfUI7gPV9N9l5lty6LieHLBnDafvkpZyKOs228j5csuZn
y6fKtAZqJ0Q3dGPzNtCCQt0Xp1Hg04AiY1VwPA0aR94gSj55o2k5wJy2BCIOXmcI
DtgqKjRzzhSj1RtwOkfElxNZMhfRZdBX84CgY8GLelrU5Puug1G9+80/KpZApCdV
3dx1YgwOGcCpo9m15+WBxXI0BYWrlYJZkMxhCtYXptJNiyJi+rYGzxVaRIV67UU7
RVzTUH020LJh7uUVidpZn6pb9uCeu/mb6RFp5Xj710QSJpAXE++ECovS8tSUyMqI
6tf24xX0RVBXRDn7f/oDvnri/WCU85yfIi79f/8RWI2NuIcQ23g7Covp0UgpRYmK
aSslFxQrjdrPc83Gpyc6yQVgnsIwW6lbfL8awpyJVo5BaK+86PfSuSz8XrjWupi3
chTb/NvGODZVfGrbRHn2EtPJioKqBwAYTdfMUZupLCTLh3jnWehPqgR9zZM4y97R
gKMFVGfTBcauYG50uw6YXB6ktrd6h7V/sC/auDHH7XQlbWUOdtwuKFCmnW3Fbg/a
51WwoR/uZiUmqPucThhcIHdVQZcsdJIHqWzJCmH+8BqTilQ76I1l9eCByHlQTDz8
1CCHvVzZINrOf1LZz5tZSnVzj5s9yRs+nePT3KoM2FNAnRh1ST1tT0xhn8OaR/dv
4CudDXYWMQ6htyFzdQ5PpQM8Z5bcxxjizNtb4HHPmAL1o9+9ieix9CHLAI9xoZVZ
YyW8EOEZIFLuSp7mcIu6sFz+sbj4ckJojBK+nBfkqECyGdJx/BT/SVz5bCqp9bDJ
mdatQGYYYeYBau3ZhRA7YrsfA3HLbUE9e71o9Fxbaz8mqv3YlkT1+5+dUAFGSZj2
9GpfhqrlJXc7vwvh4JWykDoigWW7KZlmzYK/3gYXagGVDEKpnHM6IGplsNBb8qrC
//VIa172/xWCMP/NsEuUIk476t0nCgdCyU94ncr2Rlsgg0N7OowosxDHY0Saqyht
NP6RLoLFRYYg+a7KgRYus8Vsbl8fJndfScbpMcmQmU6XX8sJodjunPOE5Oya+LaN
nHD4RFESb4o3p5PInBD8rZWRj89/X7AQJaKFf6EYGGrUltB52e9VEUS3X4noSGv3
rvORS/JTE6oxiQYViKFu04SLUl/E8I3j1nasAUJNz2s4NZjQ2UlTdCMfxtzp0uJo
1Yf82dcFl4ASWOxwfpM+rkxFtYEuHxeCoYSHEm4hioH7dUsmVz5z9715azNReWHy
JE8c+7wbzRHtWCL3TM78ajSdz5f+COCqHI7d21RDov1iGOYzN6EaDPgbqgFibURk
S8agt+swkg2lvBa4Nn1V6K6x5m6g3Zcsw99TmGZrsDZvu/0t/YlKTuwx9LeZIy78
DfG6bIm3O4mW7BeWfGVouTxkJLRSUG6vhApKt5SmecnqWl6oWmS6+uTlUEdsOUmk
58aqAq2gcXu/tyjQTsJXMheoLx4pKKq9Y4CR7q+HGasl1PjS83wroVp6hI2j70Vc
N+UaMh5B1wPGDgoC7OnY+T1Pqt4MyFfYun0iM0r1ZaygmZNxpPYZaQ54emwERWIi
NWzOnlOJewSquJbzMjSo57IkQWvRvrip6uQPaNFvP0gdKRY9MVg7dKhi6pKsNQUu
ELF6MSyrANASBCkbSeXA7BZLxoDuVVnENGgSzEJUOQqU23V0VpWrHDqFjLWhxXdH
B6JqSxxIKpagRzx7BviNDcrTohilzNRiaA9s6ZQmGKvEkDpbH6IqWy/yqLPAHSmo
7MZ16RmuJmA7rD1MaOs6bg5wRsLwP9AQZnqTh/GigDoF+g2Si/lMA5bdaiATRg0v
DbfXpfMs2WrEiAavGL1lZQhPLYlXw0T+zPH5IlgmpxDEnQ601kXZZrXtOoajT8Ik
i0wZDicCSlENThzjPYUDxqvrIXJ3f40JdwIu9sHZg49VT7X9FEcta28gqXSLZQ2Y
vF2PPaq8qUc+vysi72qGPnFyFJ2U8OuIH175sf/Hfy+vAS+qQmmrNN/DWHTyrIbx
WwxUK5Nb3fZbagT2TVW6rULBY57+7jQeGPDKKcu7K8l+y1bO22WSsRuI2j6tB9zj
U4T9Zeu0IMwpQTjSMFcoXCGH4Pb/5MbFb/z4j3d8ug+EP+EHm3i8/aeS5os3qwNR
bnGjJFZfjBdlYh1rzmyR9/QxmDQXL8cO1nhy/zgn369llATKRHy48o5KRFU53SXX
K6SP2kKTM6gOFV9W3SjIkGeZhSYpwcnoPO/xFachIEnVHFQERXEhwekTmkDBOVHy
3JR4+tddmfX/EMgQVnkirxvS1l5aEZHftBlx6O+pRfNvQvdHwXskPbGbSjqmE9pE
SMdO994yDqtyo+C+4taMJ6jNdRlQZSVj9GB095vd6/RpVYBeS/qzV/t3cyUfmDxE
AG4wzfA1ce1NKFqekgkF9Iq07F6bfqvVRBdnU8QNGEJH/YaKRZRs4rK6uOAHxUGH
gmwCAXmmhnUxmfpRGWQNX5CfP3KV+qM7gGHEpcIvq9e+0OQKPj1OZ5cJj+QNUc5H
SSfCUYAUj611m1rWlkkoL/IYsWvMZVyy0rIr1C03THbnjRV8FVyYPOvfKPGdsul8
PjHhDWnuXPytYMe4i9d39LhVWVML1EnzOvvtD3EUcoLCoKOD+yYVKAHVOlzXEGlG
FqSYCeMcDVkA/c/4tyof5NJqVFlcBbcOm8E9xjP7Lw4HY98sAFrnHcmZxbeK63Yo
VbXAHy8hxvH/ZTq/3cmxJc4ytGXFXQLDy4GeVl5/xUm6KkbQ25Tr0tbtzvKVy3sh
EQfZl/kltHr6cf6PeWuXKXH6pj3WT9PRcuXnW/wINyngICZldIBd3iotRHR9VB2c
gvUvRHAyxY5yOG2FACgejbeMbt6GQoKLcKUlRZv7sQwQuHdo/ZW7vP+Yb2fHldRK
7ZqcIAq1SWPPVtaiS5kolTxmXP6NOL+jaZyZL4S6reXu/6Qlr6HPogkmsuuwHso9
h9Z+rDDstm8ztAL97VJSIkKPRizAAE0LlEXQ8aQWzCTcBT6F/tNOXkYDC7yyiXGl
jQI6jQWBcGuEa4jd9/lYKk9vWakO0kHTjobmIteZ7DYqXsgMJkqF/f11YWqY1r0j
gpsd62NsNtKIKP9+NVZAj/dilaEz0glpGs1HU5G3QA/ivBLU/sFQKxyFhxGPLUUr
0S47MSdhpp9hbe6L0riOB6ErLBLlZwq9NG+SBZPoPLRGJweBebqKpc713tVi4JMn
+q8fKNlNFsnDVOJWDVOa2tp3tEZc5w7VKpXuI74ilnvfVGJ1Fx9iAXY1PgGxydYz
3JsnOkEf+HkNDCX4IzrIHd8b34uw4xLshqSGDyW/xyB+D29GvROzGbxXG4RRkBPp
R4hAY72ec6ExtMETrVsbvjrUcFWVoNsFPkUpvcOMybf63NM/WdTYWZPpcgzzP4yG
Kh9fF4USweLCkJGnYR6GpySfzSkdPpR7yRs2bEEYeXpU9AJ5H+llpSzkaWJtfOyP
Yj2Os/3NgT8p4ZBiwi5hZJV+3RdnWvGXRBwgx88YySeIwLavBsyblnpGk1m422tk
LEW3GNGatsS407+aA3i3swQ4Oked7/DaTwU6nS8wNDylKypqJWQqM2Nw+ryTPCAY
E2YPGOMoPceSlFykJOPynyQJczDIH12v9ncjIMvr5uZUBsZrwd6YrdJPGJ707Yjp
xHOCXUz3lzpTOyR2k5EonGleeD/BXr/LQoK0ViyHhduxZD9zUx/faJOGSXLc++Du
pw5oxlgz3v7kqGrFfVVs8c45c1gDhVt0zHx9TVnIO/ie0omc/dnjKpgRHvsYCDmv
OM1DQp1iYz8/7WaM5trxfRFzrRCesoi8ZRyI8BY8dcRsrtvyyGfeYvBUfZDmr1zJ
+SFy9cdScqfJeaWAxzvWVt+xAUY55P1gGC+LI2o6GlT8FLEu5rmAq0vu6Fpw890k
Ve1/JSz9atPX3j5HQ7nDOpgqjM9LcIvw8NWsMXarwDf/+WiXTsMcSriwhvCZh4Hw
yOvdhpxET3pP4Mnav03eARPPT3FljNI4SW4B6ie3tMVvMICi8rgiK7zKd0zXCc4f
qq4F1W2Qff39DLx8fKBGnXg6CbV22HxN3ni8KKtBEfXwGEwgN5r7h94Fg9FexCOc
v8/XA0OJuCnIwcUoXXMUvJvyABWRXGmJNWUQdp0+j7qGQqAiVUhR2D8Wv5RTvcw1
euunn/vyfzCnk0BsR0TXxo8Bnl4K2RjKGKt0m/wCAFX3UUKPbEBiKvKHw1lDgcc3
E+rvWec3VJvCNsgH9y+6kMnlTQLjf3sL2O2vZNaEpWslCjGXNYKmUD/5W+7aJZm0
bFLG/07UDagv+HtB6aSERIQJ0dD11/5WJz0XDGsS4I2lFioP3cbJ8b3ul52TfoxT
eqGU1QmiAcqX2c5g2ne5ZlcI8c17SRUgFkP32mzZvPKDhhB1sYNZiPdV0hjF/QOa
uFc3sJoKBskEPFfOj2VrzHNOY0cEvRNANNOnnnVEkLw3RA/zPFWTOwWKdoSZ7T5j
4ir22u6sLebh60ZXVwLlkNUKf6+c9JBRhGY13wrbbQcicFzWOns4xB/rWb5Jtip+
vPBLeWmyVD9O491Jy7JbEQPVICn8tnzDfUjWGGiKfdRT2qNm2bf2xC8PamO6cTFy
xHwNFrJJEKegGLS2+Su4ql+03Crlcex2fyjgwsCawGuidvilDIkr2GcepgEBn8ur
BaTRt+yHnjYFq3g4/Aic5vmNZhONz+nhyWfQJXSmFot9Bj+IkVZma8JN+TV+OzTz
HcNG2E7435cd+tySjlMMCd4VTJiFI0ckZkGCw9stSNIntzr/EbN07QwAu5TZyr0G
FawMZhYshBCNjhXJV+PzFY980zJ44WzDbFalhvWiEEClrOvHulyI/p5u5zq0X7gs
/xkzpQx4HxMYhLGrRuuWMlv8UfJLuelN3eCrZjvdNR8iuJed4wzbapNubHoSutU3
fOWOTc3JYGJMrutRP+GA4KHbL3yO8okqtu9Axyz4h40RK+gJRZaEvBTUN13lDbFr
XUJ2g8K26wLzcY434ukULRB/GKJGhU6zrBYH6LRQoR6HaAVjcRi0Li/P9phqLvio
O1LfrPWqfREryfGfmfr2R6tmeY1KklakymjB63OWoAr153yDUJdMdP6iJMiL6j0h
1aP2vA/f6OLzD8+Wn/vKpNhSzTnEQxWODoEF3cSPstH7gprONRwNk2HQLrPDrsNK
rf5v05J8jsb1sJN+V2unu21miccGn+T4C5Xg7NBXwhxjYBKeMyl59K97HCiAtaOY
+hHwGTcWn9z3vdnWBQtB1b8ixIvDEqm610oTo2aF0RNexfr18PSojhkkgn1ST71U
E1iKRJhkCwZSS1DwOpmdNTpa7sD7mkjd+BMLUhNJtFwQMqw4OgTQodM9MYM/YQRf
AiIEz98Vx5HrdMv5nZOXHrLzWCJoS21rUnVTEd3kXjo0XXOCf9dfXsr1wSfFiXsS
OPLPUFf2GOlwrzAS9jHsVQaVb7pvrHlCrqpHBaFPXNMemcx+Gvk8U151xJYaDCwj
FDeZ4Nbzh1yTOg3yYOrT5BsCfO5AFiF8qCgGGY7epDotIp3Djys4eoEl++h1nDNl
vdESaNeBXKPfueEm4wTeGGTN63I8DVlUjqVesSOBLPR0iDDH/rFViJKIIpNBlVyp
PmUDZWbO1QU2aqoJsgEdMLOgAkpveQ2/GWC+/fkOQ3zXk4bKcBGY2Rxdo5fUt6ir
7T6R/qh4PUJp0kT4N2b3d5mXQukuEpn39jQ9Okc0x+3d1N3SqAqMnBWK0bfsLQz8
o6NtIPQhTzqYxx0ycKguGZfH5ZCCmwK61i1Rv97IAgK0dLqlEpI6Rn1D7VDhHB+4
QNizwPguu6zf5JEWqdNnIVtavl32bRzDV+4snunwLeJFmgQ8jhMEhupbDJ5voSlU
pjfFYr0pa/U37zFsWa3p0pSxtRxPUa/NoH4Q+evO3Jdqc8oeu+IqhVEatJVTPmIz
AdDwYeGo9oSkuFT1C2KxUjFjUbaUpnCSu7lJc2y14MqFcKCjzbZBndLO9FITdjFj
wo02eAKdApYco0lJspRn/1QNsffn+cAhNxTPk0SswZXeoGPAlqyUDxM34lBcyuZX
dS00ZbhpCybDVc5M1wSxD8R5NZb8rpO5znD6MrcAXh7iFjohzrWt1kTGXXldcYZs
WCM9MVzhzTQFC+ym6WcG2b3pdvkNYVthMVnPB/Hrt3VJZbRtjxZ6VmqQy6K5Ysk8
TsXyik2SWV+5zEYSFoKu457dYK+NW7/AArQp0SUhgvMvgMiUZjwL+wyF3jTCyAM/
936myMiJT7TOGDNtDNyKk9FjVSLd9KGnEr3gfQsXwTeUk1ZZkEcX0x2JuxhDnC5o
sr6fAHsdyYV3L9wsCM03o9xv+kr56lq4oxyL9M8BLhL3vW77GPyzgna/QZ2/bwgf
nDZJ52BL164PxSvlPY0NNZUlxSX35HzRHcoIa+3k7EOTTmpdkqRdoU+fzln+tAJa
OzrAfUtyJEmJ3h6I76fO5vaMp1WxifZ2VHPpz2W1c2WS38JeQTJ89VZMxihYOzFz
yC+tle0pHTT/Zybo60wBhXyla29Q4qq/qX4WhM3Y9kLaZHeNNoT918RgD1GIsXQs
tf6WWVmX/gZuPAdpfbI909myvgrSXXJyWGhQwUykycTXPvAT0EW/7CqZAyB6hxt3
7NpcBgSv6Df04xy+YLvs3reK5gQ6O1h9tsw6wxB1+SBpREtuUB4LOO1yZ/Nywprj
3+1Kv2D/zELPm0tlB3ZU5qU4oB0OaLPzD36nx9HJVcXFC7TLOxMdM8hVfIXWjzyk
fY0+N/u6p3c6pBXiimDj0hz7CMqpQYuQqWAnmmDUWmNHrdtHE+p5wpWM8yglgKRO
VCpLpVmb4mXLJoBvT4DUzYGBc4/dIJ7PLQPWTvlb3tH32x/KHWY7OScM9kR167I4
PSvhNldzgD3PKF6jUVybCc2a72I8lk+WJGUrERDo/I06w5l6GqIhLNov1YZzxeRU
fYMVHuXSoO31MHXtyvKp31v83qDF4JbP6m06Ur60JaFxi5wFVw6eVeonCRVXuunC
N+g3E8AHxY7au9+QvGhWmec+YpjK//XSMBSgPb2+8ogE4mCREWmpDDaZpCwSvDiA
2aCC5O3LqgoaY52zynAdW1v9Hfd2cHJa3MYSUwknf67PT/eM0GXboQdFvpana77X
U4a4DocOMW463TJ94wJ79jgkdvyM3MXtF1ZC0HkiOW3u4I9FC2zElmrBM5fMpKNN
f+1QVVlW4/Iu6GRZsJCdYgelW3K6opZM6P7PE1oNrb3Ed4I0KdPWoMSpUOx1xVkc
M2vqQb9/XvE/SQEUtchFIrUyw8WEyRqWj3LW8AwXQWzn0nlcy0IMfVMnBOpYmAmR
96hFW/69sHxfRvJLJcedwxGJSw07DFjw+mLhi6F01XcAY5ewtboIcebBXoTh6l7G
TMB4Ah2P/NkBuAJ+dxYoi/A17WS3ptQDwXFR8HvQX9E7lDJGzo7ovP3iETpSLhk7
POQMXvpoCE68GgxC3pDf+0z7w4E8stuj6GXlHdY+ENpUtNyFb1ichPdZ168+NFQ8
mdYcXU1y932a2J306TUlN5EY9j5FovOxldiQom0sJjE7B8jr33Yk+utvBJqGa0W+
DJHzJAouSH4NwdL0qDOgRSUNncmsVhzL27bvQC1h3XZ+861gO2fVqH72rS3RObV3
pLuDqftw0c8tjplWHsk0BAqPaXK/AnTx6mJhzS7T+a20qFX/dE9XeTTsANA4uy8O
zIf56bwsED6XAb5PcjyNP51LSSu11pgF5V0EFwIlKTDVwghr2Lv1aqg0cSDe7nsP
4Sh65FpqBCiTSytvMLQ074m7hLq5llzchG6A2EilmNHJNiE4E4MNn4B6oaxihD4c
lV3NSVOqGKlWCg4oFcL839Tio4LSEzulxAwUbNmOpaqnrm6z10zDcjSSyY+dmsgX
zQ6dr7ZfSv7LA6WjLLw/Q7UWp1YDryz1ExRiVJi9quzREhlh8WU85BzYiyj1B9ia
vg4SBeNn+Yf2/0Q30X7ErnUgemdiSdC+nSEaLuD4yQbuN9dFbT3RBpQVqUqwnQZm
9xTW+Vdgv7hjl+ZuVDzAwRGqubD9olnzLBptrp42W6FgKMNJn/qrUNufbNZg2WqA
XnkCaUIxpfQttFnLxNbrcy8kt8hKgrT485sr49PqQ2pCCK/6PHznH1AnB5zcocUo
IXfTSogYtVpTnFmloN36mniQQjrswiK3WgQhTsDFPCMkEvu2d1/wRd20CghVWOTv
gww6IE/e4i1P4kpk8hh+BNJokoe8S6Sw25H1+Srb0L1LylzpMiZ3Z8hl37rVxMc7
8HzWTm7tvK7m4Fhywp5qF9rluUI57vCjy8x4V9YZOP65p2S1ycpY1uPJgbjnhPyC
m5j62W45jU7LLKZ8Le31wocdYgnaBAEJoSDiYh9sK43AyremraRtKPeUc9Zb6SzR
KIlD50LFk4N6XgjsNs/pDouzDmvLIiGsiKvIWSbllNp4AMK08EgnnzsafhUKvgrf
KkJ1aWkV5C1aVlOdW6r4iigUisapY/HN6JHqR/uD4pkUe/APw2VvunoSv89aH9qU
0OyaHQrIDsBr2+179K3ZPJR/Q0NtojjKahzS4rcxP0uYU4g83Meact36WbiBstEn
4/tadrFUdEMVjxLa0Np3qIDyguovid50hKpvgLTnQSHvEcT80U2vpzdSXtVv/QDQ
RVN9rAzNZdW3eIRE5RUIQRBlW1W6JK6gzQ+ZhBt3j0UEyyfcoJZ29OuXr84UIZsu
2XSK27/F2TT0f29AkTfyojdtdiuu6NkKqUg5pSp3xdQzAtRFioOd+wk+aqBDs6Ue
wfpQGHd7/GVYvIOM9H+WyI6aL6jrY5rPYDGMy9XMaQ410wi6vu9/7+Uj2+D+hmG0
YSWaPr85EHdaR9fb8+PqBIpxZUZaVUTmVm7NmC9CMxFY3W+yq7IimH4RMdysdHn2
OxKqkueEcv5m0zO0M6OZPqQ4AM8PfPQPv3Y3uf6MxRZgOEZUy/RDCwmRIQ3F3HQt
NK4UwDbn09RgjlNwBwyfDzX2ad4+EWPq5Ct6nbuXHZ/p2iH4NLpxUi+dfkEa6lTx
5NB2eDDkJzkZK+FhPYqb69S1jdrYtqGD8D0zejujcks4YagfnJBrT3Z6hPdh/3F4
ukoFDnn0bIxwhIXEVZIJK/DGL8DxUOaiH0FEwWyku03GY8zHBEd5vHRyi62Xby+J
zUKf/SkLv/gNuIRa7x4PLRNLfo09/lJ7uAuwZsoCF+uC7IEjK5zit7+hxw/XP68k
f5kd0Mem15tHq6VLTM9/jyEqp/NAMkvEWzQVIQN8tn7Yl/21kei810iVIfLg2ynZ
teH/Gg8LmU6UtmqVbq/RCLPF04IlhwhR3Lv3juE5UeW/g8WTnu2FVyjzqa+G1DDH
ftdIgIxF2pMnICMj0M26edXMQY20AM2WEJ3LhrqiLqeuJ8+P+Xc1pbmSToOHFS6s
VZrf7RsfESS1NTjF7sqSNmTi+NnVnRJBLt6wak9v3V2AZu9NpQWhf/rhq0Itrhyr
ir8MZRLWEq8jZncGCZsiCfkmPZzhhrE+LOL24TIbm5EeGy/D7jM5796o+SnrxVtb
xxkqFodOM1E6NHuamhpril7PhBlK7glTkfE57LasJQCmlVmDxkmAzjej6kqR6Ogz
PZ4OqTwn3ycBLo1fCL4tZ1DrRQNK3pTZjqqD1vb7YbQxa4pRNn92v/cmpax5wRkQ
NyyHE39K32ObACiQk7BC5c52bBlHH6peLdB2iMIPV9bACOfWez7VjeKeuJN8ZmlG
4m104CZ3M9Dgk5+klE988xNh2QdQvp6EdADYBOkm2xTdvzcb8H4Q34QqxdfPaQ2Y
I15p8OPPdwtgumU7AcGekVuwauHQ/xnIrCVu+5BEMu/l/QxatbKAtlnwbn2nWzbC
JX2MhmgRw3gF/78F7aYtq1rkd3uDRfkUj4yfy4dF0gdOARKHHAzaHbZcT0BMT3Er
FZRQxQvuRhppq174RkyqtDcIJdGO+3sOoG1OLCaNBsS9vcvQswU+/NHMhjybQcCq
TXD6Za8jA3HmLv/PEOUT35Kc61dENuI+xChLEl4hyFGYl9Xknu+yd2DJK6DtkgvK
ZRHX4ouSJ8QLVvI9xirbChe/t5ov8WMz956tQsvws06vCXAktaEn78jJyXRGCWjF
A/+/W4xFBxyt1eyfKMFNZIh+0/xt6s4d2ZOn37qEhKo9N2yvqkaLbG0SHDk4mDi4
zndctglcNZACaKpSziwZc03swEHljO6lGSmcLuQ8Qu1izAPS1DSkqOg56ltXkb1b
5cMscfbT6BlMTx9mPuKUyoxvfERWrP9Tc8ktLLubfTl2rS+vKEfvtj0cgh9Y3Bnw
Ewlq4hu5spQOqRgtoKRlk+ebNyVXVAgjMwEv1m0VFF+M/srn00SONaRAF5aJx8Sn
hEcI2pgmO7C9vLyMSfBO4+ugxOLNShBf8au3HqgSGEUNTVsoOevPTpkft7yN5csV
TNev+mwj6SLpFKQjUsMYtRf6j9o2eW5Amk/WrWDWrokOqXc9tiT9OaaAcu2fR3a6
RLRtONqsGyiIvLyFQoqVr8twzlf92rc+1zMNKZNhI0DajSvCkOpRcUuzUPcoF/bQ
6VYgAzVXdtxGc8wnhCx01eHuGp8N2ZOJaMaBVVz8JjzAuN34OKbUJ+FtyjFOPLRP
eyCPjSm+/Dq7DFJI5sB1nloRncP2KQyKKFtDv2JMswnPoxiVu2pqjmszjmf8V1GO
zwhcmgPzFqTM55ooun2zIomV45WZHEJipw21aEcspP0ZDbdm08ocmwCdGf5mfWb/
x/pwzyROXWAF2ulGSoT15EXyP1LAFIrxMogkq/Zls94jjezNF4GWFV9/vxeS5P1e
7qCu3T0+vKSLEe++MMsAh7RbRq3sIMrySB6N+6Gvngr0X3SYRm6S6FfBlp6MA+Yz
4zBReT9KWMtiKwcbmuhe3pJSir+CSaYZ4D67ckKBFnrAk9hoQw7C0pesITPQwVQp
mLX/mmyGM5P0b8hfzC/Uq3rNm/ZFTiX92TAHrIGoo8tm8QWBmpwBaLc8gyB6+rwn
NaCF2V9TjuhI/hpkuxUHDwkcXOObOs9hNRSUUVjlYiDBwYbZKnFyFP9nIk2GqusN
pHRwaAYPV2R7Oc0ffBIcepEWrKdANI98bs0qCLWsJGpCWDpigFiTIg/kf5uF10/A
OYVTNRLFj+pTnUj/XmKisuaBsbIwsbSw/qBECdNzQ7v+MG6dB2McVlCKMSOHrmr4
Sg31Rtu1JswIY5pFsxqviV4glSSNFKnp6ndq9iqTw0qG7RhnHvHonKc7FV+AtkiS
I4XOJFV6qNnZxgaEldLCVcktvYOJT7HikekUztVCK+fByvkX9aYBihJ7edCWX75g
+11gMlDqUwyJujExNFkudcfCiKHyrXCFXzgKmcJgdLkMeTqbN0kVlN1RdVdLLzxl
q1zi5st6UBjwMZZzVo2Xbj8SFbk4QKMx3UY3xqjn5/y/iV2XVSY5zwZtd6cRQHhn
yXJ4YKbUoqG625O/sM4uxnndmgE4WV4C3r53vE4Jaq7Zx4M2k4z7wWDATFqWkviz
RugQ29k5/+Pw6/rCzUM4oyS8cikpHHspqL7BClqZr7BjIHcUQfAMr5GoJfCr+gBP
CUbX+OmvjQxpUdrGadLW+hwFjB0MZ2G6G48KXe6A7AAL/qGGMvA3lIyui+ckTCFe
vJUWcGrh6dvoj76DND5A8yRi+bxq2a2oeJc+xxJDC1B2m82qVbpM/QITNqDbvl2B
6Bm0XUTTpLt7HfEUUms0CkhcZPrPkRAyCRJ0qR8hbT9KA+LgjHl7jlmkRc9dtPSN
mSOLqgHOxEvEY/YsEKlYUs23R7nqlqQXIuwtOhwo0D4kiZxt0HZkdqCyC+t8l8wX
mpvb7QwK7j+ix7hsSdcdrztQ2Xo+AVS1CA1VHf7qoWq0xlflr2+Pe4f1L26WYYSL
WSzrSmmz42JQCuD5tttl+BbRVM82ggIZuovY3pqh3xrB7gqgGaAVo6e/xR7iWY0A
xeVuva0GiWUOOLgk6ODkAfGLfQGzOmKIQ7XRgkE2oVoBofkDtYpnW2hRJ4zpkkJ/
FIXbBMs9SgwTMRppn72WoEUikOkub14KzvqpCIo2ab0tLeNs375kESunauewCoK5
xCuKTYW9k3elafHilEg82plP9fDXB1l4WY0AGEll3qGGS7WKZVdNuglK1+CNX35x
6urBQiq4UxxE6QuABRG8d5S7zbLPLupDqQcgDt+thdGtK7Fq7rSo4gfX7covWMpD
F45BjY1+Rk8zLmDhSfQv08Q/B24theAB87CJQFW9eNziJcr2auljCJUv9Go+89b6
OX8QSarV8Rdgd+g2VnnyJlEtVvu+OTgGDYmrPkFhtJdfgrFq4De5J9ZR5rw1X8X2
Ydgbu8qo+k3oONQhijj7WHVwt3MA1/NgQmgqAHDxaz2M0DNjHBnus54f2++D1cKG
p8ZY6sMJFNjLHke7ezpOr3yBSj5hWDlxgswW+87Do2rVVKqNUU2F8B9Y+0Jxdvrl
e6veL3b0yeBAe4VHS+ZOAYxtlLayBKk7hCEregV/pSDpNUY+ZaBnNt2XDQo1kBMK
tM2N7BOKZK5UjaF8CoY4O+pPnSpb2UIE7WlTNTOvZF5qPiMdc5d/WJsSEH/EKVVZ
fADxxv8QCb6Vt4ezC8o90GigDItXh0pNBYOl18nRWpPzGSmv7lrt1xLMh8AtpGXu
ux00sFwf+rUmYpS2Z2/OmU6pgT6kXQAOHQTR7l9pYvXiLVn7g16tHTJ+4RXvXhfS
lgVzwP8dRo78ihd/X+BFfdPWV+mQWtmXMP51ygmr+k/boEsMfcTU0XAQsQ3pkMar
vTzsfI0F4hK/gCzjgM7MBuDp4ybGQ7opqPeZsKK+8YSFJDLxf2tV2nP9oAyMmgAC
H6EP3GCv/M0APJ4rAxLBatSODk6QW59ytBYC09bxpjemzEmBkivBbUlGBEVfXbkM
4hdZma7QdKHBow6WM+Z5K4gH7164IHj9fCQzj6I1TgoMGtviESZYTeUXbil8qNEB
XmAoGuZ1FxgE0eWWthQyxBH1u8oLCrN9iZLJ1+XmeF1kwXeM123IwAy8bgBsrzdh
cqslG1zO2FETFXhJVarykhDbuv9soD+9CdUeNRVbBgiISjcC59JyWjdYHs8y1P/k
wLiww2JohivW7/u0rgJegAQd7E5VpobkQsZIwgYrkzjShzm6H1T26uPS423flQOC
MQ6sj7KJpTEy7yjQDphNzj4liPLo2pksANxxxWANTTHB9zR2GQTFZsptU1qj5J7A
7Pv4gMNOayHe+jZl3TLxrpQuqb5wK6XxsO86lwQKdn0RX35SLxxcLNjzklaI2wq3
mP5bN1Vv+cwgt5N/sOu7CUjygQb/hocA6imu0z48He2riL1aOhOHTP27RmstcRCa
kYFa1lzlu52oU5H+sjcOvH4K5zLTEvfOkMBgrUFMDkmTU0HA4OW/wBUHslHvewwb
saEGTNfDzjVZ4J2b7OQsKKRt+yXtEa9UodKsaz9KUoc6HZFRqYEXhcIZOKowC7Vj
Xbvigk3yTl3swzH4faqs+12PzDJRKVyA77CX4Zzi8EDnxEonU6PxRh8qxxcwHnME
Djp5VRcG+uXy3aehaQ1Mr5kRXdIQRY0VHzDf6qO1OztxEwRLpSigZ1I5iy9p3opG
yAlpMK9l+uE4gSxZjtq8Mo5BCCxts97Or9XEXP/Jr4w820a6XB4sZJi4fUELDyR2
NTWRHazZnGEuh5Bx7b9AG0lh1p8p+ayAg+ZD7zMWW9sa2cMBRfTkEzaHt4oATPV/
Sfc7iWmkWTP5bxQwKPQVCkOD2mLOxCc161xk8lzq8roVglWoLG1EsBMy1e35DAa3
Jei0BhLVNeJCR1u17Ib6CuiJPiw8AmZhiRwbRefICCHyGpdUvp53hWqMxxUX6l+5
cLiVawmvjCHJq1Er/E2lcT8v1eOoa59TOLIb4A0OSMAYe3Eo4RQ0m2P3ZRvyDpL+
uD9l6KUMslDaq0Y6BKPNOxZcNctVWIjC5Xt7Hdgvd4jUJTciA6QBU+df0J9ZOzHr
sjbPH9So5E/eIyAQZSWG5FNIu0WsWOlEqypSjdHwinVX7kqe2nscoOMDW5PshHFg
fKUqB/Zx51/zEk5P8IMGU+pN+hxKfp0rd9LoaZWkvsrBcAjuToZYKpOUaX1yhuT/
Ya0s6EdY8S/tOIcqCqDtJMJAHr1wd0AhzH97OFqtVPLnISiIl/eivuF/GhjYrq3L
x5xrrcIysGZcNruZeyFdM7MUm1RpHTH8AKjBn1A/AoSd3iyhDdgk4eA4FpiiG2lV
5ssHoo9A4vEcSDSlsVom4NwujB2krNa1nHpRBzaggXwpqibgEyUDwqFri7VUdSQc
UJr97MwArPqtDw45QTSp/UYni9fN/DiG9fNLl9044xMGqGn2nhDw4rC5yOvxaPw4
vaUNdENsjmBvS6EBbj+1zXzeThzflm5ktwGqXZAzs4WiwnKuq1mDZER9TVyxAvpW
AW6EuNGLksvlMx6xZz49zLi4U5JwVslPlUyQzkZH7BZF75AEwxZd+aVJ9UZn00h4
NhPbNDLRv/qTn3zyeaG8C3Q4HqmHY0x/wLODL9AWeE0jfyaQpXATfxAx+AV65YTh
QHV7oOnv719G36dWGPZSeFA7uesx6QG9tIKm8zIlQ62HgyUEWFyAevQ1kmT3AVfE
Ny7dmei4LEa/ewEGg1+jiY8xjE9rjzrVTkm9uNNm5wzuiwRiyr29Fad4HKnWDxcg
FZaPO4CjHpms8onfewJP2r3jbVIlvtNib8dga4Ine/6itNyc6ozWGWQhQpnjZMti
F3HZmtNT5ZxnOJFa0xDujY1yJR+BgpVrPYGRBezktrT6ZTlpVrag29Qikk3Gfg5O
1yxa+G2HGfa8RESccMosCR7Jw1Ru6ReIJ0KhM+rrnTCgY2t6T7/yIX3Ad+f2nXxa
9QnVkz125yJRkBRQvAYrGjHYpig2Fd5XWvdPLVCNB7tOJPIYFjVWtmzsL/1+6nua
qwoMGpxg9W7vKYgfuXz7oggBEJcwvvG0HnIhigFmotGBLdKC+EW4Fz1GrHWF2QiP
zBm//mznZ0HVztrRH+0VY+LpRLdJqp8J/LLySMYRKrT8jG8F+SKNhs7vZdIu8I+h
37HhRoY3DTLfxrCW4NdxE5q39BIcpEqzfj1bECeYetlOi+9Y3RqpYZllsJArFWCE
oN8JxKg/y37IKRKBRrgcYKoV25nm8pL6M2qAnPss4SH26899a8ySHe+sW7Q7eHAn
Q/uEqMusWJ4lq7ubeGpaVNZJYPA1tt8vATK8v+iTtDFFsTN531nVMQlbjyPlhbHp
x36nrtzpRasFjKVSd+PRP7rafg3GS7bmmnU5+R5NveBw2L6eXevuc85HuFmKE7SA
3uEDzBe+7xxE74PdTwcfIVO85EC6Dcw2ixZcBYxmbPLeJhhotEeMU0nf0Glt3H2X
kfFgGEaRx8Zkb8j9yDPsTGqQ7uObpY84eGylRRJOu/HGhYK5JGe2glT4g8eOhSp8
JRv+JzVNONtQ9vyA1oxSF0nTi5OFVG7/Pu5qymSJGcivEFK3uv96A5bFzHSGJhVx
epIUaDRjLjr8W65vJ5/8DxS2wqqonidMJpKieZGnP1pH/h7nelafa2zQmke5WTsL
ScwBCSeOGRpvWGzvpG2zOcmqX8JTm5QzrxnduqViqdwToE1IYSXy0uMUiIUvYlki
AH2QE4eeeO0nO500J+OvUlS4EX/b64N3cr2i+eSK4Xm1ijqHGuIfZQsiEqyuSvqO
LL3s0BNoT8EEP0salrCFj4pK3JjX0Wa8i2QG2JIX2sMj+/VL63vzXf7dGbGFth+K
bkCQ19J1BM3niad2xPCit2T2Wbtz1BrosDpykBXewc6UBlL0lqjpuk7PUBokFjof
EU/zgyDAxOTZTK1Yb83tLYwBdb3ZPA2sbDg+llDq+WVGhm/ieZ8Zjcl2CqKAW7d5
CkFkrSFCWzXmi13AU4qaQ7WWjMfdwpucxV3014nuebvGC6pfA8p5nypmkIhocFW/
r8aO6TWg0ByPUbz7u31z00j2OqXdtwrMJjMR0zquONO6DIn69164d7gA0MmKqM3N
eT1KCbk9RloY7RlH2vN3Wj5v/5FzmPeL3rmg+6aIwpDjijdH4GW09qHqj7ZH7GO5
U9tcNiHL0xFYR+Qxk1L9CgPSZPL0d0sa7fmJ0yicF1NpCa+q93eAlpTT0iEG1rgN
db8/xQZv/lrQkcPRjb3oPbT28yQMh6Cyseeu+Kbu/C/zwzqJmxjaH/MFlJ9bCuqV
Mvi4LaPy2nS97td6W+P0JL04wgTVVtPsMgOr6ZsYORqs1r4v22A6wR1OtFSeMmr8
F89sFaxWcMiqK2i10lJ2oNq9aqQiLZT/58+psDE4xvOGCWRO6vSha7JMIOLj7jfL
Bkr5yq2/sHlzCSsE2A/V1cflDyx53dKoMlnhDE/YXBH0LUAFB4wPcql7/i1dLYOG
t4AD5L+PIY5d8PpPpDSG4fRkDWaDO1LjuN6xSDbt5UH6VAU+XqA8k90KYY3EF9L5
BNggTgi/P3HlzzZ/8j7Hfk0wI5HOBk+YD2fBppu+zTGo1kJVj6FbIgjUoaDkMZjR
R3xafj4mllXBJ0XTDb88goK/Y8eFKo+plW1o+DOfYgwFBbm7QO1Z+bOY5E4EkSzA
UTbI2HRCyYi/kUW0eO4rhPsx/+3Cah9PvJ9YWzOXzcWgjHt0Vb8mknc6Z++qOpQ5
wvifaeYQpKYNi7lFyc4YrskNY0NTE4+hd+LhrBy6A00xLpxcJ5jxFDRBl4xT9ABW
rhiEYZWrqxnFzl7xhCnT6ZwpAkDpOcs3ISqYTOAMgZfxI0OpohD3uneTXIpMEO/p
y017ao5SX089Fk+rtpmApNUmwpFj868s6c74zZ4FjsMMNxt7c5hXT8zY/sD7kQ20
N0zS13frXiUr0YEd10TzeW+0pu/F91Nz6keecAj/6ztFpGpWkeTmOmcJp9u8b5XU
1FQBEksjsjHny4lT5eBbzytyk+mozb19Naz9RmJF8Wh36E2y1b5O/TaRnDbieKns
pU3ZjjfCSd8vw+rR8UhphuON7V831yHM/R6dYooESiL/1kX/5I/i5GMAljKAaBvO
+4sFH0qPbX4jC/KtSOO4sk1hxiTx5HoN9ux6NkfjswQlssrDQQQe1iiJi9mVJRfT
gAv6X47oGAJzOYg3HoSsPmjufwsEoe5ID1i79WJkzwVQBQSZjM7sRQLVrg6L47em
U9vD2HYqBhi7GwWTvELKNV1mi+niXpmUtr0S4qnGvMzivAIUiaEKgJpJ04/Vp6DB
H3N29G4XjZpUJh36pAQE3/v1VIeDkodprTpV1ezyr5KSpDMZL8ogYvKjzg2shEC0
98URhCcfAWEzWCGUv3gmtf7LTok5yUySd1ExGnvy9a0BqrfrSjhsp060hiCGn4yE
D5MvTUhl7Dnz2JI41AQ6ap28RYUp2gASbg61dFc3R8Zz22aqM9M+ZsolFGrY2SHr
0wZPuDZtq5CtU+8lOz73/irVlqxRR2QBwONFGeMAMpKsJjR8lzaiji6qiOFQAbQV
yXp31uKw84ZQuFocmVxrs7DTRa9PJTYUK1fyuK96p7nmr56QY7WbxZ6gBHn2iYV5
7faMiMHBvdPcWSitrCNaco8whWdYAuMDRBdT2lZaHVZB4JyzjSLnGDW6jKebne/c
s4R7VL9GB+5Tia+PL7YimyzbZbYLWOyX7ESHH66yzHvzNoyZREmkoAGx39PZI8ob
i37gFa8gjgAP8pw0wOX31ehkDzcNvvCXdsGLiZ9kxhTB9BuUuPXA3UCmkwId42lo
h8BSPfEH9GlWeq2z2yBVVLNlxqLGhdu6/MojhTRq+6VBClkFlm60R3fUJ4n97o0z
eCRX00oFjn8Wo16zNuJDDchmofDcU0TDs94ww8T1auak7AeNqZSkAyPxXxW+jHkj
B7D8Njy5cx1WWb8RXi6iJGXr13ajj8h854x1rwvTfXSzUUjrxw2+MopGSP8igFyy
ilwy+9VzVgllj1XZbB3hrpchU0Pys73AK48G9rciIFEWwgi2DvDGuV4KNnuFGfOE
L8/LHB5m35otNwa3S1HVKRU2VIOK9Ad2m7hrSYVHdlq9Jm0/0JqT7Ic1BiSGxIYj
TQDnMuYlG1GhjKmd8o1hTVTZGTOu4f1RKD5hmHVofv5GeNGAMnvtkuMCK1SA9UmV
SrbMdTRwXe2Mul2ytunXsEXyyxF+VbIh4p3mqnkRtgzDVLq2LtQmakoAZpfW2r2g
QdGosKtZbYWnKb5/bYzbvqP81KdVgSZy4hRygMCy5iOf3Tr6ci2COYVCPLHz8EVY
VZCJU/bTdYe/g6wdBhe748M2LD3Lj0JXoHFFhILueODy+PLahuUKlFSu5oXJDdFN
mftehJouwJ3h3u0ALL8t2KoJKv6xibW+7pLtohDG4rVNcuedD+ZoBVtR92UVVocG
t0DuQVg3BHyXeDa/R5FlKnoCp0vvTXVyQcbbQ22d3f+QL8/hOO7c4H4HDm8xUXCQ
g9PtStfSdFBdP99hZ3cU+rnlCuANqiaJwA13NsnoFjjjzyurOXwSObezrYLWpys5
jDZjTgdUIZ92ZtuwE+VqnjPirb69p+rH1GoZSqVZnz7TAgWSj5E9oVEEFmv5AoQA
YI+eji9SxVEj9N6YVD3FPKhDGgIHDtFBmsksexr1iYwlrdV5oQpo1KWGXRlooYX9
cRK/fnHO1DDGDCkI1Z0vJU4csTvpqCio2m3lrmtEHA7bv25bOThBXza6tfPlvIki
rowIv5WrlSstfJmzqbd0KMPChVEKV0yGZj7pa+4TMcc8FuuZ2DxFJaZD8ivbH1An
TfwG2URN8vpZucorOo/qC1iQAOumeoSEyLHhbZjJGYvXfkiLaGrbZKpdwJtQCY14
hUG49O35NfOSqiMhTCTosCal72Kly+zxFWja2rYLWSl23EpV8/MA7MBEn9SeQ+zd
pyq6vBhKwBh+N1wRLvHk9qAfzE11sbgjsjB+43usev7dfgLNnS1s0uFX/Oa52UPU
QfmBroGGYQ8KQt0id0RGuwy4x6tqcSQHd6QMSfjtSX8D9uSApDaE87PGzSz5dVyO
rRHwfGaZRbbPzU/1P/ocdL8dgEsRF0kYn8tey8ljZhQWPjBWgPt0RQ0nLIdP8Coa
Pgs/L3J+E3YM1Cke4wjdnz47D0GOQhaIoyDrYv4Qv3YW9ApiLAYTB+ELNhSEO2hf
5gMlUBugdyAqQfv0KvT5dwOCZtpn0wTc3zlB1SyKRQ3gbpPRnKOR2LrLh/13Inmd
vweGHamfs/PEo7iK+/5urmq/+V3y8nDcbBrx6GDR7IXuUR0Q1f6Rys2TkdUbhXFK
5gqpXn9q8gb++j0HSJCReiV7LyLY2IjN1tpnDmcvYNm0Qn7fhJCGXvpPMlwbxL2G
BHB+P/tYwFNkSYIpSh2jFfMIlgRTABy7207XgxG9H3cy0QFIP6h0eCHiDRxpNQU5
TIEjmO+gjbDCWp6rhMmFFtNe0bhKSqW09hKsutN5fCYbpaPQrfJWsSofSlsFPTKT
f+gBOsZwrFhhksEf8WuoLnXUkWp2URbk1M5ExftG4s/bkcvBtYU/lcbObwoqdkNo
GTHCss8FmxOTwa2olcRqSI8g2oSGYqXdwKmioBgKTOdP0JwFWYhJXjM81BXvyH3I
BV+HkSUdhw/4pqwUsq9xC8VGS/LZ0cUK8dBifDTiDr1zo9BrPESzHGZjaAEPbUiB
2JzZPeG5Wo7Ob3ZREN8xaTzQXoqzc1POHQoL2DPamwlJjgjSixsqNciR80aeTR9j
29O4rtLcWWpOjg1G9Tkl043LeVqDKsJTVUskZC2lpqZiJv55DUD8Gy9seZg9Kl7F
bz7d8B/4iRqPdXqlGnqVIxROMedME10pJaCQJrSu4/HmtLIKmTKVg3BgMu+DzLCC
fUGR4+y3ft7GMneQUeHYTNZSJaybpJLi8SPCKA06hBH0lEtAnJwPybgYLuNqkZGJ
SVh1ErEGAmv5qlPKVpxf97XTqNbpd/j4WkqCrwl4at3W4htENTWvK0CvpVA97w90
IUi/PoeBn8EMVKV9w1whgaglK6WexNApx9szHV/UaRTlWcRH0wfvp/dXF8Wu/LLS
vhuEEiWIwfu5ISm1YTbrIeVtbtGiehrQIOvY3SsQ+L59UVJhkE9XRm1Rj866vVZ2
3GhP+0atJkD6eV9ZvgWNGkngbojqPtKxUtz0f4/grqWsNobrR33IxSJYZfYRmteg
dMmj2pUn3ikK05aaxf18Ne6sNYm9TkPNcOcP95gfPsmnTaeq/1Vcx9u1UlHhfbR6
UnFId3ozhFrFTnPrYvkh5BkWUQgxFtswlil6XTHPXGgCImiOxr7mMjL88QZKhrX3
3gPqIVAq2IWYymCdR4hP7ruaPibuqIueq7aV/0G647Khy1mf6fsXvNhLva1KHiSv
1GN1wkA/V80SS2DpJdURwPIenpoG7CpPWdIm4QOZkHWvFxXY3h2whxfnH8NVG1E3
qsVaODXkSRMu9u0ARlQ3GZ4ocKh6SyxK7kmjJKtMswyoknfNifL/m4bFPA8wXOPa
8BMSF9kp5Le3ciiSjlDQop7IDRwVIWiXgvyi8RILnJTPBz/Wa7CcYwMtyAxUbHRs
+xE4TEYespmWCjHGQoEIVXTpetw+MdnRzVYNK51eLqlJcT0vE/n9d3gS7FNOFCya
3luHJpaCP3+2NLH0GJ4ySPWEkKPkwIUV9zoR/D2CcYC58pIh3vaFsCE4X/8CgdWO
Jh5qTG+gpol2RdCDRzP5Tq8Jb3EZYPVjb70AkzmAXduftiu6JQU+FYdolXnl54gt
G2J7JDnf1KTuTjiO/lrbN0SLU7YtVjNc8Q1db8IE9luUi108fV6oCSjTgbnuUQzV
u8iCTX68RuzNdXK8kdQaEYXXNLY61lEyOE2Kzxy+2k2suEAvomK7xYz3uaz4z/9l
reBA+JcmvNMeuYmFLgRCoGIg8/OSaXPmyvgHFQIwUHpmsWB1Kiop4fN3jOxf1F/n
6RsEtsLmbmNiV6bAjbunssSptJC3gpzCFrGTsvQ1dmpEiGQEXmY107xcltQ+lcGw
YlWHQv/muNwC2p+nIEf8QTLD5xrvszQHfeB7H371ISo5dcw7uVhOXiI5Qz2fMICl
Yhq/yRT3QkmuDqkK8KlODhQyfze/meTojFjP2+34Rh9jUyfMWVCD1QN+6QuF2div
ZluFyVNo3fqGI1K0a+9QZSqoRo5/te6mLbtzG1lleubkTns0gG5YMZ2jXGa52PsN
XZ9PJslTFJSdPpHN9uW480Imk+MXHJHBEnMvSY4z7F0eBgd/gMabVJpfxcp1ar4r
DgVJfaFWe+I9HCqK9+qQXFJDqJxSzP/VD2DxQa0/++hvnIhiQDuBuORLx6EQ5ZKD
25AtB49MAO0to2W5S99oS5iDbeasYqba47ShbyTVcjPx8HAg/Uo4BVtrDOYgiGks
KVzeoGVvPO17jsmP7HHrPQGeXvyVHf9cRqVeMzqfaz7iu6KX1cb9kfDJ82KUWJLk
3yK6uKLeQ4DGzVu1Dhdv6Rmq50w207/Vvtq36NsdOWdQ37C7QlA2EC2sjyvvc4og
aYdzyziZM7J8T1KRnvNVKUhyQlAiqAFQwX9FTTK8jeXGt3+e9e+lWy4yxFUlluwo
d78rVGIxUgEwduR49Z7eiktiBtbENCTJQvVwU1QixHTxkAeZ7bmbfUpTYtZFpDQh
Dhj2HZGO7Zv7qUOtjsLyovY/1gwkHyBDdnFyI8Ln56rKvLLT56pc3/3WMNSjLHqH
5RmAhL2GEjJRyNViv3egb4uBIA/w/j/K/xakYSronwrYnU3QLPP5EeotQ5HN7jSM
vPd9ylh+KqB55LJqOVK+U93K55EAacj2c5+6Hp1uWcGcFPCJDHlWUZv0hT6oyK5N
A4crh+TioQiVAYn/ffGySzsWl/jgBwuz6mxmuLumSPeQcpfoI1OtFtm4pm1mdc6e
JuDRF9koavTZpzYfMmVzALUFvQOfCgYQDWJ6LU0jMZCz02ms5PnystYAjhXcRsMq
fMzzsOy4SaK2/NcLeFv+us6fC2O5V1sGdojeYFwYO1mrHiH5d52/76olLwnS1V9f
VsopnLjpZa6rVXX+HRYuG7Gytn2NqDt1zDapQYQoSr7rNoyar+7YazlbffZfyUUa
e9eJefSXHquFmtOdFqnHXc0gXk5riKCAQYcsmfiYYkm7RfXfF7+7kEWY/JcLWbnd
+LboXYAn5XzCEpwMTI0FqlPEGh1GXplwPX0DLXeWv0d0enDYkG2RBicMnmbEDGjs
RUzh5Dss4apC/kWeutXMQQ5cHNN47y8Jz6cj4UWQLnvMN79wBf0wlswsp7GqmqGo
JJWZ6OOVRr9Wa6xgmAemH3Rxz2cxRsp6tjInJtISUItwy19HeoRfCB9Dj3VLy3xj
oKi0TOyMdc0kFwHN76/PG+gKKUTUHVlyx4FWvukDHWnh6O2HTXzTcNI9YqgL4oF8
zNvgXKMfU568jhVXVNAaK+NFT/fvOs4ZKP3hFKLnXWs/xT6C3UOmucCpaWpSRCwm
SgUK9udZ2xcem3Eesg3Gb/FMfAmd0WM9udHTgsDgvBXX/Dh5m2uWqtftpaPD4ZqC
FHmfzo31pkrut8ewlZaKcXZ+PUjZypvnLThPVY8ZHCUcCWuMJe2vzlq/ewgASfB0
ZWdhf011IJypKOvfrGdWrUFyIpFGV9NpzNbzolQz1sfoFb5jexFfiH6t+sMfxl5y
AYhmyBMS33i2EjHmp9rXQi5OQo2xvVYPtwubxUHifeacs3jdA3ASJG9ttzLk7Mte
XBiqRFWerFGTBzDLaEwbAcYO/HDxUhxDWf5A4ckxC6zaxHEJGJNezP1oWfaZr2uL
yrExlXCq0pPqytk40oVSNMcNBAHMio3H36WRFZQcGQCq3peyt4y5CFcvnf4p7E8p
ME8JsPGNyLqh3p8o4TpBzZCt26Fw0iVH8DX3w7CExShc8RvUQiFOKQyLqd1oq7Fm
SktgHSzklz9g0kZwDDznwBN5KDZS/dI/Ag/AhlbYSGrnvK95Br72wUJF0K4lXFsh
CWElOHW9H2YWLdVvpnlfwodH1/ckPbPl+8LeoQKbCZnQy71PUqe+O8iOOV8cusfC
15iGDhSW4bENkS8tT40qfrT30aSx6WoMSf/IGNMBLby4izpfri9e1LkESHy5VygH
h2SLF8Wp+pOCkzSf6X7MARu4tNSF0pajDxbY1NxUA7OiR2lHhjpnqY0hOP3R57zh
cGKTceHOV+Gi5+als7PCkYbizy8k2ANDD9xwoGz4l0PwhfUyZp3FDb0QLsbHd6ub
SWJOBt17gLHXmSEhkZmaQtgesk/ZVfxjXUCe7MRfa0nrf8SHW1rpZrP9MuRSgfuL
GiLbzjS08iUI8atY/CSalfy68jHaqr+zXrFvkoP1ILBaC/xKVmUsZ/pr2pDthtA6
+1e4VwzL3pSs4PraRCmIid3I5U/pDKr2OFGUi5Pvt5fE5qFga33a/0s+AuUdYFmR
2I8PxSRbPDGvozl7e30g2dxdaObg/aVT2gAFHR+uk64W+KxCww1ct+DyPbukW4DV
2mxCqGEjMVdzsreLp9DspP6pVghUpga1mcZPWBd/06EHxj6VkW6+RxpTYTmQkQOb
UCpLkJUzsFl1JTdnKOyfODjAa3Q7kkdx4rmXmtMZzPdLrWQ2dj2zYgsFqomqG3en
YpQBo+KUG8wa+eQRVqwwvf9mAcv9M+Jae96Yk3grerDl9heK4A+N30fmatmRRos9
UX95QYRPisEeqc1oIB8/0mCo+ZywssOFZTkx5wbiiq35hCWfXswHCg2BSrzUWFax
qOdUf1ePToxjPhgJcN597X8nLD70V0aB8SjTY4KJLOYN0G3+jGzrp58IJawsCy1i
QmJV0zg6jkMiJap/B10ycbP2hi64YI2LyX1pY0mgippY6yjayfMmOLFnbJGJLnAX
XA9PcHEUp937ugbChB9qffJgVeVs1Ju7yHPSMx0J57846VNWXt5Uqgel9VXR7V3r
RbjEw5CXQRJPaSoKmkP3tjjam6xZpvAIJdxmYCR80phfEVs0I67avHBPs1iTciK1
gxT6R1fAs5n+EQ9yXVCVkHt8250qQWnXGjRardJWZSxV59vKkHNEfmjlmBO0S8nX
mBc1nzYcP70TQc8Rnj+Gp1ip0Hjcqf3vZLRrXo9pdoY1ylDAP0SfrnZ9Cq+QBfdq
H2FFOSG7ee8+WHxHxRNT3qNXN2YSRkJD8yy9oW7Ij5HF3CmwZfE+n8l4aBMqYfS2
SdgXDxGzwTbR0luMv6viu3VAo+ksK69qwXrEv6XrAKGgg5KBYU7lao/c2jh7HyC5
8yDJXvIOlIz5moBqc6376X0TMxvDtHbqJhVJM4gIa334Ml+jIZojvD1R2YJXHKTr
xYHL6JaRTwFH+sf5VuHMc+lEIMcOnFcv+GAeOTezkGfB222wkiip1WHGl8buQhty
ggnn9cr2RCGv0tAogQlbixkI9G481+fGAJSsFcUDQ1fPoFH1vSRhYXaE9ou50ojP
OH+G+EaTPtsSkoHgETavEuIrzCK3fbza4T93DIvS40oFJW72P+r6gKzAV7YspjJe
lcT2uJAvCzB5LnwmB8nepyA2AbKSmQW0BGrR/khISt+o0LUotljd3WaGu2RP2Zt0
4N1PAijGzSnPiLQAbqV1lJfZnxziPE4BLzC7AQ+ILCX8EuMijM5ZJj4hS5yeOWvG
zlRM8I3ChjdC/5xQ5VPOJsCbcmv+7HRyJW7jCSEQl3qL8ox0RK2sQ2VDAvtMKfUn
zaIqHeI9RonR6jSgHTrP5atpDF+d1SabBePo+CPa3xZQ6mSNnD2el0TvIe14kNaN
a7iydCftkP3xfLZIB2WHHhswzZvPyOe8Pz5QnmYvLL935q3ICw2HloD/YUupD0gS
+Uza96kd6HE5cRjpDLQffRgOKFNtFFBdWkH4gfj6S9cEUsQyY7a7rs+Vn+wTfO7u
ETCLWUVb+9LwlIKijKClrkbLQDSOlt6cIiSIgfH4lJ21k7iD7XmhhHeV9KPT8K3j
zf1pBRo72S5UswMDHEBHAmyNLtERCAbSA6iFJXwP+mO1TorywniIzzHWkb5cjoC4
WRQSkkK7XAn0hV8Qqq237IZ+6E0Y/O2qioMR5ZqldeTjrvPNi4xB48PLRJiVXP/U
b1rMBw66xAE9ANdMws1xFQF2NcMiD04zZeeCU5LsufQJ9OaiyF1EVwU+S1aoyKR+
T7mTA9GU49T+chStM1QkvGdvBnBIOaw7jdWTntQWDUuyIlwGELIQ7prOzXxh2gXb
ftNTbtMYsaIQVSupMgdFoA4ulOXbCE+yiQbnvu1HB9/HiXqgLDzhxbzXWX4p+w5f
OiPPXwgSCSX6f+ghbMQmZaODFnQQv8SCDJy5dp+2AflMSuI6IvyEO0tHNnGbOfT9
VD3FHqwTpyeQO2p7tKYnIrEqFFeL3kJ9lNVh5L+yb3rwRFK1BNa592Lr3tYIrt/8
OQJgCrp/dtOiPX80Co4s7pqdZAMCGzouA32tRTg2bW19WVkdxuIdUUyda2iv3khu
Va5ut+v5A3FHzpI6mzY+ozcm/JwbiBGDhGgGr9S9koTyE3eMsf0a4nc3XWtjKZIh
vxH2hCj66vksjJBM6tid4HzA2TSw67H8oYHTrvD/DySDlYLL0l6QmpiOEO661TRS
55hcp00/pMbvjQeEH7it3558V+IlykrC6fOfsVcZqgM+jUvHR252SX9e3lf5hliw
wPe5tV7y0bADGxQ77vzyrNkG29fPgLlugYAXumRpBQFHLljwAyHmsusB9/AKSZIx
HLPIIuHRB+nS6nYS48QbGF7uqiVkWHg62i/so1ftmoajNU//kpAAPPVTFGhyOTaQ
tc7W4+vqx7KivrGO8kTeSPDr+MSVRD5PsG2U9GaoXZNH9OeLFwuhBq15T/mevbmd
IK01jKSY2lNGSoovdHoUZqzH04qcmzepG1S+wQAA8fpFZ+czoi/9L08dZuL196D6
K0r6w5hfgnq4JuQc8xsHRngKpJ0aMHBL0SmcTj6YQGPZqKKLmPPGcn4harm8CXns
Qlwq1Xqnc1x/todUy5Tp6qL4NrJ1Jo7gaOexOCduP85l4E5mqnBIXBGivQJyeKQ8
SyCZ5hAQRLrfx1uuRHrv+xC8pNMJqeVTgkVfWFbYDXbck0qzCydxQBPZDRwYcj3j
HKa7oU6+q8bF63eQKttPR5QlWWjeToAxDhzRrxVaj6c+vOb4B3Gw0IGsQjNhoiZ8
/17mf2SzarVn6/zMLSi8BZ8yxbLq5nZ6QnGcKeXUdxq3CAh3yeYflAXuae5cNcIr
ssn4BQZN9kTP/1ceEz92N6XpQMGvEV2vGjoGU4jLf1FsnsBQV9CBcj786dsE2+7y
WFNX2CUXuEiKHopz/0UwOcdRSmsJiq3G1O6jJSSAKIpkAdsJeMY/y1qy6NpqaJHs
4fyioqOCkCSHC5vDB+S2d4fPkDrH9Pd200inK28PS20r5tkxdEvv4tRBvoc3lmCr
hQBTWjEgvCUeQBbRS7qbL+eFdDRfkORJ8C0ctTBEZukQsqWVa79Scc/Y/JtC5H88
ngxK7ax/QI46fbDCTGkdT4en3FtMglqhAkdB7NPSR9rlK0/bjIGGpGTVnmp+MmED
zR1KDQJeglfhJnTiNvDlpSpH2EgKnuUNxp0Aym9QeQmEiEfZDsXCTdWStqxdn9iy
ZBmv1P7qZQxw54HwgbfhE6mJNF654vA4ZRR4kAS8LCZEfaKCm3gf6sFxirJA2nMN
QgtwPDG+G547wDEeoJ4QzPuh3FYrKuWftqefr3auEgSRrgCs4tn+iwgJ2tS9x69g
FYf33YK9/cma22Fc15Tk0WPz2HQ+IzkFWdDRqQpcQCboLlg/ADfP083jYN46hGfS
Dh+luGeYgkfclOYdwEgnB6uAcJ67d9qj0swpPglJTNPsvodcNFJo9bVj01NyksqM
EvTgi37GVUzesD4DvJsWyyj0NiKHn84Bm8A7Ay/q88jTyPgMQK8/yvbHT7ekxn1S
PKuPROfWfqOlb2La1n+vDmEecyvMbmxJvNRA7mtaGzsc6TYMMviAHgSdGnO4QUDW
VTGFtxw50EkCyp6zEyZq/pLv5//md9mR9XDbciE6ZAUf0F5elFmrAiQVEbcMC96D
YRzuiuRXmIFInBp+XNt85R9N1myjUiyjbajidkJS1SUlENXVsqwgwhbw0qM68DlT
I+I31kfkZWsSGjDI8fmYhcLtoOPbPhlmivGKTbEA49TYBYx98+tll3DAGmn12txX
iVY6erNri+Jmt2qXew9I2ZoIxv+oMdLp3/hHkDF2LXoxv8aa7l4CWmbdW3aaFrfn
mCM0jvlj7JVJrCBoaQ9gtnetu0PufZ1uSGMakvZqfzo8sseSACg/Pe5HAsOirFzV
u+Tgpyea71trenRtfSYHpa9YvUP/fPzkRxDs6tORsE1bOYTXkNLD9QrGmdgz6KCp
gStirTF5Ki5I/FJIQzEVgqXW6KargnPIpB2uVMYFn40fKyiQlQz7COaMlsWUAUZS
4sSjseQt2jGOAMICp3cRZysfp+01IfNVd+cmFVNltPHuauxibxKFYgjWceQ8dwqS
EGsHTpKdMg67KnwASJW56rvyleV/kXpRJ2AJ6j9bkyLKNkyD1a1Kvf2wZJsWSxsO
GgN8vkK52gAy/CalD1+vfQw2EYEMG0Q9CEH7IIabwtaV0lfhMHBxAxr2sjRoa/w8
qBmRbenRATfTFDDimdaEwjdVB1pYR5u+rShJ3/jJx1lIF1RONcNlPlnhK22GoExz
htqWKL4RKhEa9woWTKLuDht5d35b4DjBTTtQnlMG54KQLmAhLlWY5zBx95K3GtPv
bgygCo0JT8zMCUX5ekd8Bl3W5gZENlRIacKd32i3hzWZ+zmJNkJV7sgyubMIgdR6
MxHQackb56WsG4MT9YioruY/fL4EjvGf3F20Jc3ySGYDRhFxtXWq7XnYEI3Y/GdP
De2cjmd3zdQgeHfGQ0IFKoeNbBwI1WLZp/KX0/YRmgoYs5ocU2AynjbmwBcMf75q
ysmo9bdWCvxfjv2rgRSXEtDGFyXrzyXS6C4yXGTGt9GW0IdCP7KB/FSOlmUZ44V2
4OStedSFORZQ4KEqa4jdF54KcREU4PqqhYZE8m2/5Hh9bLlGAVF9L6YXp/6TFgaF
q6DaOYCF48D72yL1ohB+AWazo6FF2e2nVRkGJzJ+CFBZKv+fToAIWGJQAluncbvz
1YwXtgBcqw22tmCRLVdnZ9GldTTnHHSmjFCaadsrqHJ0+Dx7AFTrXA3ydS3siIlz
pa+XCWPRPzn0MtlXzLXOU5JaiPdIGy+mQa5f378SgwZxYs4pHy1FbkFY4zRfXC1K
/yObbLzAORRARIPCdOVzGZz2odCrna5tzGDZIiwqmCBhNACLdKBkpueN1UrM568Z
ThNZAHB1pkJ5MYsf23DsDboUjB0Hc3XUehVb/NYkw4U53ahRaHxISaU9G4iOHZeC
up0bABa4kJJpsKf0ID9VzA79MHxkG89CAY87xDxZmqYZ8b6MdQNH90bOYiQY2bK5
wScdnJ7gAy9H0EO6UkiqATuVxzLYkPBrqDqoKNx+sZhjBwV8t33FWaTxlTV5Xgej
yZlGPoRESlfY1bFdLdiOvnV/aPROWbLuYyAJifzWqd/9gRpkk37tDwH3H10tkSaU
q6oWpCxvzq5vihBrcGcAR3546APxcrPwGrit03IVFYwVXn0c0S5YMaImHih2qc4F
E2hG290U+zaFnW3G4+2N6NHvfBAr9NXKQGXNhKB/OvxGRvOb57koDoCSAO1YaIZx
7M9TSZvbYJazX3W/CV/PAauBf51TTYHq1QUd4rIJ/gE8RdASN7BIo0bdi58XcAfh
olRI5BqTMECfbPSUFa/+7aKQen0qPeQDDjsl2kovCS2ZQ1cS1/EJsjZHa66+VpJO
8wW3wtpw/zbAhS6uJUUXLQq+9Iq7wvZ3Uh9c21WgTutRGxZIWK3WEJXivtuHjMWN
pOleN/luYuU+FsfDDBUVQlb/vb9G7GVmeycet4m2DgLAU7Q5Rnswt8CY1E5TIXyP
lZ1BtiXzhad3bLN4WaVcYIKtwi0WR/26UdUmbmF4xhCSxA0xrYIpqkzipLv7JT1a
T8Y4dNYQMZKaX8XBiZtU3QRsCv+Gvb3lZug0FYLBjlZi73br/DjV8XR7C70kJfhc
frkDed9fa6S9iwNXowzD+KibarCtW535K6OXkX/omaRFezMUtZrNw8WFf8Q7ZJvx
9NsscQCVy8Kl2BczwbptjAXHw2lzuS20QrKzMX7HF2dRTkzn02FelrqgHeu+JDcz
F+TpqSlUrO7wfPp3GR97b6V0ImPQr1S0TfvnFef4T3Fn/Y+8FVwNo6oiwGoiEigY
bbKeviEw3clXQHtQTDzycsldyyTLEX/A9D1tmAnc48us9ARCWsKDnDfpRqfsGOEC
DF76nanOSv3n8vqImJiadRTdFkmYbJWAD9Ku+QSIQUdtFlw+uaPvC2eVq/JQBGwC
V2kWuJ+DxQ1S+BL10KSDOHBPODSh7N/YC7KJEpY0sbz6CLv4k2xxRkwImXSKcPiA
HwSEo1L1xAAhoOBc+7KSld0y3fuQfFlHDWKnHBIPaMis3TK2SAebMCOw4Ryla6Gf
F7a/jIbFGP2iqhMW627ddzov1xm5VqY1WpXIofAicRL4sVHuIhOi4r6DHG3t3sXJ
KN3jqIfiNRVskmFd4dbJcJju/UlCYSG+XIOLcM+QojqEeHvJT52lFhbSgN2+foyU
IOCnxtrkpZ5FfSTGXXlW/gmSEMKyawQOQJvEYhJB4J3kV5rYIz7B26eW6VllEBeJ
VidaUh44WWahXSxCv2R6L13lsCZ4k4VrW7MQwVQXYstsENQiZ48m/1YHmovHSfW4
15Pb+YW/ecF7x4Q4ZEmM2W9iUb54GJhR9VtrASBM0nSJkuFiSkLLkiUjr9BqtRXq
uof+913loqbhm+j5Xpek22UkCpm7/BmS0cHXps81On/UHqlZ/LS4gePbHQQCgLh7
6PsJwmCLWB7Fuxo77dD9bxx6FpXI6OrSd/gIEQEyDhoRJZ2Pulu0CAp9cjXKpjeR
rdmTbHZTkeXBkYhZubExO5wIaww84EzFUOKG+7djQ2hsMv7q9ezpFfAHp058yZVJ
6xqzxFxz9feIuu8KCCFoEldrvAIB2j8gzYuKNgKh3QhCpqPEiDSdV/YSTjKQkj7/
MicLtLJEkAe069VNU0eNRLRp3T3B+iNx7btckkt0i9rLP26UUKvx56ST/SOavTeq
ADNKuQzreKif7nCOcyxnNP2utOlYOUrQ+TT32JmRHxDhLMIIIjwkK8KgooMTvspd
6a2i5RlrsiNgSEqmRsxE/nSPVQuJb7dYCUUycpvvt36pHq4XEJo764ShI5Y5SDuh
BBVLZ+gEkJCr+X7TfJYE3SUwhT0dpbGAplWcxdVXrVvAEk4NIMoqz6OOGczPxvqL
WUiKB0iZ3RM37KHVjkEfcBEOgF1Ucx6efVoTbmMu4Z7zC9NHL4+WL5alEEqx0+FT
bokRhkIVKdNbACmyHMqeKoONH6zEuKHF3QUMRxDLNbnjrVUlGuoADC/JCOONKjNT
4y07niuo7zkXJXGyjegb965yBrpq+ZPuEwNew82ioTPWolAh27vwD6LR6P6Z3kkL
G2u7XFiTbD+6ImCy6eEveTGiIGdEccOub1ID+7qi1cC6mh4HfSOVCQUx0wSYBnYm
lRvYjUN+9LIvYJ5FgXVfMFYs/fKQndjoFBg16yEbXWxQk8pY48qyhS1RUgWojOJy
J0Yi1mN7BNpGC/084ZDEUOywxGVcE4HrjT1YK1sf11StTYFDb46/rSxFHCNAQK74
cfh8pED/bTsoYlhjoxVKoJSzpzV/Ra6flytmzV3JCFqZx7/2SxgYD+EYsnMz7wG3
cMmLvDR8t5mpydDYxYHwuYZkacdo6xQtSKPEBovlnql/ipZ2CJaAaEOonEDqb7aH
L5cT1mt4XBJH5ojwWf3G0xZU3gq64RUNRVupVlY4gq4dChAZp6e9WgkRE3QNRYVC
94Y68DHqJZ8XBn9xBAuS0nJ17oxaxQwGlAjHRxZmez0KDDXsyNS9EnOkT0OUIOC0
QPxDqfD64NHwPU0EA60cUKjAIl60BnoNjr006Q9DhDpktDWR92uwiyd9o2AjSiCB
ykmj2F02Rj5nOA/hrlI7opUmsLQE5/mgz2pHVI+iNn5HQQGnm9jHZu7ZNkeVaU/s
Nwfge/NVNEFzOro0xtJURjNjpgNuY3hS9OhHfqc7NlqgaTZcbfmacKXPHdmTtTWK
RdNkmCNNXcsJtxrYhxGPeenEfsXNZ5ixPLlw4YP2enFNy1GEyKMEFJGjmNknvqxQ
y68HdTnPrn2+ESD1puy3OFG59cTggJYgSbbeupq5ICmYVRIrxDdYP7vvt7tCd3/E
TyRKSqpksusNbg2cSNS0gMn2LDZLHTTzvknbwmO0bgij8Y6+oMFenkhNIbMCS7ah
jd8X0vXyHwTByGbmgXOGltVE+s86n9m0BjM89cDkZVHVFal0IF0ZyGM4ItHCY/0s
G4aj7cg331W8rGUle2cc4dOPft6xj7jHvDgPwaWyrKwy3ge7PxRWPsFQTE4IKO/O
J3yJwTzVbJbnuFe0d0HGWELl/bYW8Rg9rdtTlBSRlXJ9+T/V/wMEWQqHS2aqoaTY
9V3zWODhEctbUeq4nVo0X4pKScjF5b3v19w3bmNriGXHGa2PIDkRQhqauZsshVUg
0iX35cetFdgu+37aLHhK4qeo0n8qa+TmcLtK2++yQrLVm3PMFbDFZ7ass6yx29mO
+Hl4Tv4g37nOk+9GYNGEFoxBsleHWTboFjutkl/47tvhcE7x/Vl364usQcTVPqzN
GJXkbzHGLyaZ0FtBixZ8UiJENgGu6PvytE0nUoNgXHx71cOrcdQPK+e3mp0heoVJ
8E1/qzmyhNsdNv2k+CVFN5ZKcXryt/SSI63gLHwZlCe491B/MeujXTmtvZfw/3Z8
ou+5hj9sbez2pXj2VKp5h6Lt507kqqFcF5C73iSnADSYt4KIZDjEFthPwhkm5p3A
iaPrGNnXFfNzWZ5ERwp2DdP3o+lTDd0FLdjczJc7Uh5CIlLpSjSYKp4f3AdzViaS
/Hvrw0xf7Ljy2uVp3llHJ0BofiYXu1b5z7jCXR7a31OZOsgMDs5+B9jVix4eeLPm
pAkgde/WcOMROiVtSI5k9PCnJSAsuVzjVwmto0e2+HN5ja6LljzrYcQlPTXRFut4
iuGF9FGSkDtMCI6QGiNGbyFXdt4NwFxZK5OXSlwzHCszvCIJBpXPc0laOkrseg9x
Lbs5j/0dDOGA5A6LTaU+xkA3oqeWYTVKFfh5REgMAMql+AhaQgYCIIuIo1Ggs5W3
WKunNQG6yGx8C2QWzL0+OAmIQeDIDleP4HF5EPoN1s8AYJzu+kIFD588NYGvHyqu
j2AdGpIoBBWN9Koh1pG/yn2WUaG3DqZAjlciDPpa7c1RyZvnjbHrIi55+tl8BVRs
fwJxBt1q8FuZsltqq2OQFKnuQj8ql3NkExmofI6oZ6vrA+eiUr/cCPisNUQcfeqn
6l3iVBskGZcD+ygSGhrRSbANwGMepMSb8XIfrCa1V5SoLNp+hGQxJa9upeu7FkNK
+YTRgwMKdv7rNHr72jIZ6EUiiq0nTU52C6oXybzwHNtaI5LUE6axMeFK9nGBbfGu
25VEGYSedELtysWFUjm7uhBR6USJ96rYgfS8XkcKrOjhmgDqLnO7jAkAz+pAL+k9
gRz8i9R87z3uMJGOGcg2VUgd21kQ6+gYdWScal3GyiNp0sGhOIeogL/fo6QqTNnR
Hvf7VyX/ZNnIysa+ZfpFRvfBgSAU6G/1IOvEPVl2PjBh9PHRgszrNtEv7zM6XYvZ
EtI8Rw5h81e0cOYNun5Ef0+uH+biN+Qj4yKis4zxyFyu51mnoyW71gtsh3WT54cm
c0oNUMfQpgsLUDBQRd1fOXjIf8OU1umJ7oQzHCQ1UKo0nNfTBjRN4MZr1qrtDy1r
JIAIGiBe6gExetUors/d4UT6wq1HV9kg9QBnxH6QeKVxHCYJv41TAY1u1GGBaUlO
M+79LPNnciyQmx7o4HgSu97aqju6JK0Jpxwu5Btk/IjSVzCDSHxnEvk2ECovbt7T
0tC+Xs7AFpwe1W0xihsxeI10v977ulj1MmdmogKRkRdvPEgYYExLrYN8PO0tUEdS
l1FsJ/ElAXNdbkRniPUgHuVzA8hmlhPNvf4aWuW0ewbqh2debPM5jtfrXtJVoBA0
ponxTI0eDIvyMT9q8IsbpvGJ2ObzYzkktSKUsZoviV2qPODV3Wlq3AzbN/YjrQTH
TxTG2Tie+rBI/or//L9Vtz4sSqtOGZTEtkpjnPZRYrDWd9z0FXtncpowgwhnmdCj
Tiiu21Hn21x9RpW7NePrsSmstySr/l0ud0mnqdwCcToC0o9AXxnihwnCUls1ueDR
u0mvDpYp9eSmeWCkD/ApurVVuGjoNToANrKI/b4Dt3sGNv6tp9tommSv8XLsCnVP
Q0UBZIKALgJniIj0ttuORZr8dhVjRqzsdyZr81yJfV8IRDeoRUBJgKBbwFEfJeT0
JYA5PTS6u/PcBXVnFlYZRZ1Cm4wvHCMqJdBOh/pnkzAYe+QuGLQs3myr1WlfFb0F
UnsfEvaZhaVPE+LAsVQfYPyZnrKCikjVK/qXEX36yFDVHdrtGgpVcOClkNYPJCP6
7mHi+5F0EbY1U40+4tuLi28ClGGHVt3DYTid9mVLqJWHeW3LkN9VLr52xnXracGi
tASBTK5WVxkTG2aHslZCJojFaLw/ttYJICgZ8//37oUy1ykm2kws7WwVzqBoN2vp
UsD+oad1Rb3VUiFlXI4GzY6izmb07XjXVsWP5uEKvLFXZYA4QF+M4myDsXy9iRBJ
Z/2Cpq9pZqL/CQodXL9qish80NnPXLcAFW8ZXCwjjiSjsGRLp07IRv21roae4mDa
T8dWdq+RbKxPIhOiR2SwiXegTfhSDUPxm3IhvuqQrNQYj8eiddFumkHiQwE0yk+L
OfegtN53SZgM/TVB2x1/g6kXB0zMwpth/rfnRhcfr8Hdt8nPmuO5ch/orzpYLT4z
yT6adTRtBEJZwai0loNjGzMvdD4hlvh/84x/wpCBFjwBqbx/sWM0TNBJZdLYM2YI
c9VWue2hsfRvHIwSrkngtMXruu4eDMSGxCUYwlb1N7xy22f+63srlk7YhJrQTYpG
B9VHhankJri0n8yZAfrcJPMrj+AIR+P3/Q7fmkuYy5SAE3byDpLh5FYdnzVDliIv
MwyKe9XkQffn2vWsO3sfSYpIGMcvYp1eMOGt5ve8SJw9FctZOLaLXfn0IcFuOY2q
LqDKIJTKlCrnPScb8iOEZTFrZ420BwxVXdlQMe51nyberzciIfV+bMWinOqCyuEZ
4o3V2IGQ7otQUlVxULSZGeQPKpToi7ucuGEc9Xl6f1tc15CPNLMZOHFeYoW1YKry
rJdbg3jfKLTc2DnYsCy/p9FH60m4H/NRUgWVX1z/37xCsDymA1rsDtzCzOAEe2Xv
0r5fL3tHgcj2QFAuu4zJmurF/+XpDoIzLrS+U+Gig/5jRHKEVrWUpKDLsLkt0krK
A/J6lWyJ+sIxpFrUluz5r+4px9qjvfPAxytm2XPa77u/G8Leh+dFN0nXKTZUfUld
v/MeTEUpjQogmZ6M95nc+zjasnDQ2s8rasLxkujeLcOTP0847+DYY9HtUcZvMquI
rqoumVhMqmppHKR4iX261tujmAuIl3wQ4+MxX3Eo7M0naVHnn+DHnnXyu75Za2ny
GBJASP32tTgO1Mh002n6keId9HKcKfEJKOFKIULwrjDwmsNdasXgpv4DTJgL+KqZ
cQQuWp+dn+iZ351FCZkD4pOERsvFsmCR0JhQ3zvZFWdrOxQ/D/6ugEoopQT7WSf0
JfKXRZkhLnJwMpQIOdS5dD8ZpK0PYw6wy/o9uxto2IQb3AaJxN7lfJlIMIylVXM2
p5rkaM5IGuwxsIazZ/MTp6aQ+pFkiubCYYkrAWzlG6j7OTKod+IosGCHIuQPQFvZ
AREUkooStZWIhR0AbxHuAms58MJYFcAQGzqYxfuN9a9iCDumPTp6FZfu3bjRhqRY
F+q7aoS3LJBB2HNmTbZv1iPvCR3FtMBeilDiacbnjGzDvorY/cqUuDLeEHX/JBk6
W16O6FhXIlQagSuD89ihTO5E9NBltNUYcw0v6EfmS4j91doFs17NY3bCkBi3FQIZ
YVJXhwoMLfFbU0R9GdoE6K4IJeUrhvkd3sk+FXJif/RlGoZzojrW+FlFeC6/97I1
rCpHhr/n59hIqURxDv7hRietXI0TXab6uFfa34JMke8Yn5trYBeJldwHoP6a2Z/Q
iuuaiW5G9i7mkPBd17+OtTO+zudFQfXmB5BN3WZNQUlsXhI/YSodZxvNuPhwO7Pa
J45EqeeKjDLFIhKEB+rwJkMlhMiwYAoQGTo8M3iQfyi6QHqfE6x2hPLFlTfiRQBk
7C7d45H5ubffVMyQ+3+LMEISq5zsDiTXPvp1twHuzdfndDrgVd5wSbRY93/40ePq
cFIS0hKKa1EC36NwCXH4J3l2wyJRy2u3lekPuwOu51dVMKsq3Y+cGWYqkz0mSQjz
YJMMxWIUktYyScLw97eJtG0zCZOw2sEbQaqUXo9eJQ+sGHt3I4WUtzQYp8Na8xDT
B5BQS5ItQMcyyOBhdlBUS1O7gzLn+C4PfVeYpTJ9ovX4Vnxr4vHvYoaq1IRTe+rO
SdKUO8LrbZSzn4PP4mzsWKQ9RnqKJEnJ0F298wqKY9UxxVHc2evhtQjaYMbD2nsz
W3faN+it6Yfoz4M1C0R8fM35oyWQMhsFYbbqpzsCHK4X1uXsrmSKIl31O5ujguTW
ym6I2LLxaZmPsabQ9m0xkej9c0E6zBTwoeO/1s9vkNPerTbsWR7sNVpSvpCJixCy
xTw0LjxyS9njQqVm+E23zy0GU+YhI/BHaJ4cYUJXMvCOvh86D0ZsFjpci3TyOqWn
k62v02hd9HFyg7busGnXFjsCxN9xNH/EGfamoCuKLAsjhNOqs+rQDm8su9VhLvqS
T29TfZdyZo4bzq/nD5jOt6yL2NWVMYQ0A4eI2JpLBJPSOhu2Vxmdao+DvSrbGWrq
QGqmfBNEy9MJ600/Sm9xxe7Vty1KLDaU+f3KGBM9nYhKlHK25LX5/8ymoDiOjgrn
FTGhPAgNvENa3VP1NU+D02CC75G3Ts72a01GptPEait2kY4qmB6hQOkYcVjUY0ya
WuWvU8lQVr2IGmpAGCN1A+uFogYYBfXoKG1yE4cPJQ2kCbidSh6S8qn0YIHTTEHc
4ulSqAR5bWMRI3rCoH4ihFufRS+qvPKmFseIjofzQl2P4A9dXnoBrzVxzMQXt8Ln
qMkCdYXycsCiwii0XpRIcC2a2TG0KgXXWptknrmjMSr4BRy64U7wi5dzMrEpMMjj
L8F8UlfDILYq8syZi7vR/T6fu/bTQ2VQ5Vu3sTHvD82UJAF4cFW2pWoVEn//i7pJ
8QdgP+bWjgIYMfIORBPEZUqSppJ6+db0RDS8g7sG5J1oXoyW8buVw/un4Zd+yYqL
8+4jivJjQ++k+xF20lCrUGQh9Yf4LL4oTD1a4GnvOaHV1tu1Cd4U678swpkU+dkK
xFSNfw4j+lRiSzGaarCzXWN9HCpxaWzPjRNQgsK1C0mAHYW8miR6sxpHcQAvdHLI
8rkrzY/khrShmlaJ6u/7mbldRIZA8/4d+cwMRxiy5GX7jTccxdMT04t1Jn8gI+Pv
RO87FL+DCbHER1eQLiSFUJ3ckC3i9SfRnfG3sZ25gmXPgwRN8m3ginbpUX/cAer/
KLKahsWKl2FrCRr5jmP8k36jNZwC6mk/wG4ZtD9hc3JsGwQGwCdK5e4rIyBMJ24N
0J97J5ThXw3TNORykaQTazrLP6lRXDdRM/cBcL/U5ZkFFRmNYevnQVDvO3Z2kG3Y
FkWtWtbjJprBJSNmAPGwhasKv3HGm2SWbm4TmmDDea4sSIDMjaqTI73oo9KGSdDP
Vh3c+dRQBjaYr/yNtrQnGauyKr4DNgLsaJKzYxRR03wRwjmjkQhNxjKYy2SREZ12
RR7ERXLdWdQ7m5vwWqIShQJZ58Ea0oD9xGp/JzvyZCN+5JpnDMryy2lKl0v7/jEX
gnFR/ttZOCxFxkPtMWR0gz8Pjbwxd4vVJzLdGz/xDhVOW4kXCPvYE/c3RTXq2Hil
D9af8S9g1xrQ35eZnAcAOn3whRVAIDY4/JjnU+5wmjd+w/N9wXUjxSdYoxJESwfQ
35ZwOGCT5y1ie1RGt9vkgB7oqNzlMs0Yr0XIRLxbDJZ+FlP9teqDjKkKPQAWfcFi
Q5JiDK61eMZjz3inRvyTWxN3C8l6gTMPZ67i+Fih9TmrnqcDzK9b+7PgPcL4yja3
QAlgE5S3E6AhX+fx3ACBcuXI49coOKdD7WnzSA8WYu2Ocl9kUIQkiNNpwzdc189T
TAyQNqEEEOuQjS0FofzqSMrHkinJus1ZBM5V60Gzs1RY45CyfwXwiVEzOyRfX+r4
QLHiA6t2VFKHOegnwlBUS8n6EF1dfRTfSrRUcUlJ6LgUsakAl8UMVmLmoApZ/7ti
nlRPiz3rzXFi93i99RFYDOI3v252odFtn1sKZnJiPfSbLD5XbDQ5jTDL5bqrcUrN
ogSgoTfyFRpOLUfN8oEH6Nt5L7uzzeKApEzzIatRyDzM5RpMvSMk/HDCCM7xpSMV
4UY9+tTPN72uuIWBdDhzvdIrUlcbApYmzp37eeRsiyJ+YP/WzN3ihNDHuCWSQwur
NtE5j1kydgzwNn17Ws5Uj4sKSL3lDoU/IlH454EmwngNtiUrdERDw2VTEZsSuj5d
Vfeu0XzJSZiKmZJOO871SIK35Tg3lySzhUWeBo4PEzUwHhcB+zONhzj49amwV0JP
hulICOTM/Wg7pIzZ1N5vR064a8Jqlpq3GAp+m5i6xYrJt01IhXUiAzAAh0zBXXYE
WkLJFToZdFLCiSVkI+jiXnuCQ1Q99gnx44N0OevfdxjXkFVhneOUTrjKFPBMZ3XF
9fUJD3c7VWQpdIIcjcZE29jlFnou582Et9yLs4d8EG5BrosPxJdgUtVavDX98sZZ
WDbZboB4z8roSDZFTvbgZQsRDnM2jka23UbNp0Xc6eg9wYaKnTOc4YlkLNog6ahi
jWnDXW8J7e9qzAl4wA/rTxbVI6QrnkK8tND8Rbbt3fTZlRPQ0usOF+OlJO8Gw8Jq
sf0i+B9wmqFpv+QnkGwFwp1OQMNaI5tBZEGbVhnuWOTrxzGVFuCugKdXyw0u7FXv
0KYU54At8zfNPlTHYFi6kXeU5tYWNY+uvLjs4y73fnfTMOJ51vVL7shblk+SjvIf
TGFtZ8M6xTeLSvubMYRgVKakLit3AK5gRZT2DprVBYMxjkzR4JVOrFxpWP1NbVK5
k/iq0hjPWtWk9C3CuNfpVsBLJ2Gqc8f2y59yHiUGVI1T3AiJRFi7Ql2aYL54pQvQ
oMMNwAW+tZ3m7WeTeySPCZzBx/5usrb+cWzz4j/tySP3rJ5O2v52ecsslUsIQcn6
m3vEmDkrt6ig6S+/zyCkXtwE14pxfTqm32tXeskPEGve1oUK59C9zm7bTZ+wJ49F
fq+SyYphUqprBeUohcHA/1HVeBaCdtLuCro4gGGSrtLEuTh9iFoMpNRHJ+uUYHyt
UU77p5uwSgg0izsqmZnZWHVvW3itApDBFmWfy9ohoNabHKoy7MyNyMJ7KqF1ZLBm
zjB384xyvKlP5cF04keXwiIpnC9sT40fYy0LhogKA+7Ns9CVpVRbTMSyCUsx2utK
rOpUpyi+0KCqRtvLfx5d/7Qc0BssGm43CO/zI0aqvxbQZaQ1mTvhsMrW3Gh4Iggj
ao1g+BNjvqVT1yVWCgoc8q428BTxLBJv18/XUJGM4NRXtQsuCmeYmqvGE5xwlTOz
n5a9ADO12H/bTJIOXQEAYqNAoC/1eQrcdVKy1RkprMv6Nr9hU8RJH6lERXqFTbWB
gRRWR0e6Kb1yocg2TYKciWDiEGxgX+mXeTBHOrx5Ca872dRfgOC/jTBQb1uDcI3K
cbjIeDTBB/SUCf+XoYBIl/vI5QcIBD0zv0t53tapYMHSpmjhUb2g3YkFdR7EQgjy
vN0n/n3t4CNZALmJn/siqwCRAgpM1f19HM14l51w69+4oKheVgAi47De9zXIRf42
pPHeEaELfHAVCbDjdm10hMc5zRQDyEd9Hu1N5MfkA9NbYmqXOX8NKE7TSXPvvLnR
u46G3s0fWNfLCvlKtKRBIRM6SQDeotDYy2HBplxNct7YYhyrbgXJodgYrn6ilQAn
XLrmJIEAsfAjzSkn6qqtlthgqLclgBMn0CmeAdCP9d528ItSj2lNldz5cjFzlR7Q
shganWezf+vssbAy2q7SAaXJx6n29WsS0lCJkAEk6TN97mfVinngZfAHYDTLqZLy
26tQshrZaIZH8e5du4q9zFatK5i/EuDK/eZEZnLDwkMISbAo2SXLImRwr94OIdft
0l2C7U2pXcXmEq4T2ocnXqYPKDBdiE53GOC53exYyJaFNr2d+Nz491l4Ydt0X74C
iGxPS7jm4iQvCyAREDtvD3lCIPfnwnSLz7/KZUPaTgJQYsk0kN4LTmxZDytHSVSM
gd3ZiEgPwZb2mvwDuyG0zaPBms7vuUaDKA92uCZz5Zvv0UAWrzHX/hTHvILLc26L
ml+AoJPMDCXUsMTEaJ4z2oq/CUr3ux418zyXfRVtoB4zaSoNubiYNYXnZVaJLpYU
oGdfbuUzU5S79HZ9t4UKp7pCyf5QchzIPofcBy8WYxy1/GNYmvTpg4jU3Jgim8/n
gaJzXllBM6MwIt8DW0qf7XZn//ufpHWbbJwcjsMC36X4a5IDKMJ1YPi0zKw0uymC
w4+w1jrZynKZ9uU0Yd7VwBxvPLm/uI0J31SfC34JArkfMNAIWIGioGACMf4jtpt3
hH1R53mGVq1dvakvq1cpc/p3cO2Y3gb1PeKdig0m1HdAZGZXKt7MC83gTYDeUsJ3
gKms5uZ5CMhu9shlkLY6g+qk5xnu5rHBdkgm2B4TkolEp0QGq/e/OypqInpGD/3W
6KYZlzElD8XWFpk1Q7pBO6rx13fuUhcCXuEz3NT4I2f3er4PcA5KrHb6uFnx9K+b
3XR0V4DJkJp6Go9YGXvBilZGUuQYXs7MsCYbvy7Iit1knwpZWlCipQyO2n6fnzNN
HIWDzXSHtY6mhPsQjibNNOdILYAfGmNGuK1SeXdKxAZrepSOLRlotJESWtt82fUD
7lqCGq8UXoYaIAtAR6ru8rXW+tXkvwfToDTpKaCOMsOAmb4ybLL92uCtWm/KBd8k
EgRGrjfcTD5KwyMHcWN66I4rOdfzx/SXhQwaYeXdmJD3MLfj3ZiPMpo2W9vBSTB8
t0LVZN5LW7XL8vpEznw3fvkMMTmDZIiRtRzXSjUlBNzULXfSFrMy0rxLkOXKGgJ/
k81Cy4Z2/hbINlhw8GcXIv0Tt/YOmMUzuSqavysAYB1kwsyhLYVsNP5/snqCzNKv
Ym+zktAKn0DKIgbUFdZaQuGkkuq8KtFNDjfcFY3k/hCLvBft78nxm/FFcdS/ucx6
hKIyCPo22wIHbtxjycFJoo61qu1TdFyOiARS8sENM0QvJ0LNDaWbl0ALdnPM2TOq
Av6DheR83KlZH+u4QlRXJQUBF+D3rM5N9eqZw39G2sbHJpmqem4Wq4OdzeVjflsR
Ty7jP6/VEUs4/6+ZzdZ8Xu70JiZEsvlgZZdSH8+GLWcyD93adinIsTOSl8lOdd+o
COZnvodqbKJFmnPeH09uwvGvic5KOq16T08H1oqirm2LXxuhUOXYeWib+gmlTEyq
Vi6YDYMKmJb3kPBownGASR5+A9fid5pYuOr+PB9nih5QvSwIVubJvQTkyKnY/DSi
NjqFPTId+T5V1g90mwAYqtY5kkag33LEnxMaC0oFi2LTMyvJcBX+MlqcJKIv074D
e7px8O+GwhPQZZavlUmitQzRnrNBqSRBn/nW49sgFkkrnyEC3brq4zr+s62sIEgZ
Wo7vitZJAdzsOCuS4HokUhzYaJnuJe5aoD07ps1p+NNZXlkKbdYzniLvv2hCQPlr
exaxSKL52ijlkBjYIHOCYzQNOUtfspV4tb3YNrntlO1aDV3melSN8GVpg/nuss+v
gTrNBIqenNP+7qR0r3vYdcdARdk8W7lh/bygaJ8szukcQfX7md2OLx6ci7FC7dBx
vPJ10ykQD7dcNhWdDX0jA6ei68AKzxAjY3N+zCExqXtuFf5jAfOSXPmR2CM6+hec
RqyWxwhcxs7Ec2lt1tx64j+BdcTmf+OViG1qVBlpWQJTPHBIt0BacqeungBr6lrx
J99v5MCAV4+PNqkfN6XE3ShzsHqOuT/pmBSlKfOYpeJLj5qxndehkh19CPynrgcr
u0JJcft+llo0MAYiMcOnUM2LvKRvxjHm5rxH/f0whekZF38aWMi8g11/XfeDvmUa
2i1yQZngAZ+9wdfRnIzIEyua4RazPk0sCpZYBjhFLTfvDtdxQbRlfp+nN3eCns5D
tS9pcZlY/rC0wTvOE1bf5YRBDu28CEIKrpJ8popjiFduaC+jIBQ2DG/9COLFw4le
rx53BRZyWcrFiGLsrRDPHmRdAqX8cDzgSQ2K1aCi/aumpsOHJxpLml5mSzP8cuQs
jnVUvnkUkoAQ9suriYSyZao0qJSBWSbN8vh40+0szrpFoElnU7oYnm3ifU7kC/A3
tPxLVhlUgMXtE84fP0IR2UarBEHKimIh2oiDIzMSAgC/Q3FrI+HoB3zfCIFNc7pz
e6QZvVpvnPddxpDoxLGU3O09l1bAHDIpsWk0lyK+lYi6YGm3WrFblPryiJmunlKv
KOJxwiKucoUSxReCAq+L6HXmO98WpBAq4yNuoUhs4xww4IZdg4Edoam4/zs9roQR
4GtZfQM2jyYj8eiJ0d+I8YlsIBMQj/KP6BvC2FKCNbBdfATOfgUVHpqIS0ucVIeJ
2HtDmYNOjCIlfw2k03mFdvWR4o2tpbJ/EzM/vzN4PJYnVqNxNFE7g8ABKhXYJJul
allM9HFDO/K17iAMMe62Mvll7BN3N9A4ThpgxP7ZCNp5KwhHV+vktDjMepYrl7S2
Bbs6fai31zZ45fpUVoHv0i5vJ6BLeLMqiWxzsL3dXl8EumHe0E5J0cVTE4X1EbxR
iiXJ7Ib/D1f3TMqRfgIr9Bivhsf2UiQUu1o7qsFfvZwO4aukAoWPun40VTvUENyD
tIQXtaPwbVW9/wnR6yp3+RN743225gYuS35PnbpMBjORteCvkV1KNyy3pXsnYJH9
WMXJrWpfnQzh1Bb2UhFWw+EcU3Wd3muDzfjzvn8cTONT3Khr2f5ukulvhJEa5hQw
/FSnGNpawnXRvV4YjJEbrW3NL/GWAnRCZ+hUzul49GkTagNOBRsidroRhKFBcta+
k1HavsGA7VkR4KwYHLZzHZKdp8zXpncLbPiX2Mkee+CbUD3oT3D7aqZx7Mo2hJ6N
lc1cYgtJPWfvFcIqKyRrWmT0p+7uOE9TlPKAxiESo2eS1saTCwU4K7ZECy8wL/UM
Za63L7WVKpsxDiw18nvaRiNY2IpgSkgZGywucRclROsXDo8mS3AQb78mMV2ixnSO
ocJsO4GYXllfbPxbo7EW89hPP7sHZhTLbFHMNC/af6jlWdslTn5Gw9lM/ZUsUqjJ
p6zW5dzC0Mr1Z/Cx7YSYlhJsrq9trect9qGCW823HjPFxzIdgnk0/dOXjeUepggr
LRI/XngclGDjZF+PhpxI9d98Bi6sIS0QcV0e3jyAPyCnwY33SiN1IZHPFAecUQB5
vz1XY0mI7UoCvlXmTofvB/5nEIOiS2IfP8f+9KjQ3z5rt7JeyIUE3YehTK6yAwLD
+Xxsu9icn7bTPPRaEU3y8K2wMKmiKceCfM6DHJXGuZA5PbMBcu6dyxtt1cCpPdbf
TWFXPFD9kP6NaMcSjnys7QEndyrjSFptQVNC296dkecwWUn4w5FeJF80+K00L80Y
9Mp/XSGT+uJEYFU3eANporWhVKWYIQmrR5EvcuhcBujXu+oE2LTMEuZJ+4Fid+LR
V+zY6Z7fKWJy1DeXdTA7H9SJvm1ZhAF+vFf2QXhw1poTxQpmyYtE/RB8puJQYPJr
ErrTIiY9xCuC+kjIsA6rYrnmyNsERgGozQ4TmDS343RsqgQssWlRhURJ9xUIG1DJ
vtmF0nx/wZNrXqTnH/nDC7qTLFaKZfIiqCuQ/dKdLGnmefn9kdRC2m3uj4oF6VlX
6NHvio1IE1bCRBlsgd4GrsS052GfHu2hVYUmGDOI+NwGYffYt2PWvS5go8bJdMpv
VFAUamD5JS9iZf4tbPju2t1gy5H4U4BS1aID1vaS6v8OMhw/UGP+qVJWPWvG0rkR
99YxGmOsv+o+gal/324kkWTmYHa2wZP1ce4lBelexMcEyHk1EwTH8Dhuy05iTg4M
5UhmFQBLTfbJgFoKl6DJp54kahH1HglOsnmdz/Fbn7AFLUcn3i116Uqxe72hmFzf
MaYs7Iw8Nq3tgPdZU20C6SPpJcCElXV1q19PtXNA2aihgrlqiD8CEKOUHbuvnlhB
ApVA9k+UUKwZrJAW48KdDatCXqaYHOqRybz0kp2eY02mC+Yp2DS0Ix9VpEzNbNDB
UR7hgE27WNOiUV+dTGZ6lvPtnO8ZQY9OBK21ZAvrXHWxGU95StmGSgH5gcPHotsn
aUsw/83MGr4yaUv1JnnIO6aB7d+s+vUTjBBW3T6LzxhXfg+BTjW72qzGL9rtBnNP
Bu+xPsjWyad8kbxnMrJ0wLmiBzv6yK/KkP31HCRmuGm/khQ5jt7nWMwk/fm8wewp
9w6VJ+dRDOv7H9MvCtYenRp9jiuhk3t90sims9bRH/6QoVsCpJHKkEJoDa0jR5G9
yPIJfiEuGs6i5ccDKjc9/f1NsqFNeOm0zM5p7zTXsFdl8kPxBJLJgU1+HcjMNRUm
zZCrgqVah9RPk5cKJO5l3nOx11piIt6A9zA1MyqnqN1z0egjpzwBZnDD4zmYNDlE
ThD1IU2jQbfuM37wVPH/B0x5z5qmZOK3R7ZTFjQMYsQHsmc7Dw/eqgrFhDR3nJ50
sNAEpDzGbB9cHg5mSl5MCckSN2xuhN3Wj4rKVPYHat8dlyr54wRt+n/lJGxeSrR+
ricdOJfrplNsF6LJkZ/AKZ+rTQKoU7GaL0KXRbx1pJ5hDV1ugHZQaPwFfn4pmpzf
zeRlnoE91U4DCIedGbSrLAB8t53l/0PLJYrPtnRvzpl16tnq3lszntKurXIC/dIA
cyWI4DDLTri8OWKghpw5yAABbcvbigs5v2k7KHzYSp52OSp+49JPS1HbCuxWLouN
Gr/OzbL8JFv6ClN6CYxOXDEI6bUloP4Gka237DGuESwhiqP4d3mN0T6Hiun93YnB
L1Y4eij8Lhdx/MwUFJXCajNhIndTvGk5chEqxpsoGGrDLiC1xTPv5n5Bg0MIxlyC
WEFsBPKUaBdJB58V6Ol0nOQxG8oXmyPAgZH07KuyEHmRgP2LmWTlRseH2wUAb+0S
emJsFYHH/XipLG0RtUFpiuIOMyApdxIWO1sW5Hcv+MQPuR8fInYCTsM68v0GqbEj
u2FLOFtqCH3LYjf1263ABR7HWodaQDuN8l45zF1/We+3MoVG3QvqZ2dl6HrtbP6U
EunQMOCA6JT/Lk65qIpkV9Hxx87R5F4g/o2w8brf+hTKVKt3W18I/PmkgAMHyfUv
JWGI1ZTodMpn09OhtR8bxoNRQ1Al+QO52CPjyq6JD77c2geYXjl319bSso9Ew8U0
9G1z3VdV/3xjRXxUS9WRyssTfMGqh9BWjo2y5K0eZHN5zuUICvbt6QWV7EVrpxfA
V7vgZJ2llosCHNbGS3kdIngIupvqfflIGsY1TPNVnIpJmpG9w7l61jN49tqXGBOD
YF9TNXgGRnuEWMrYzevkEJiEWY0faYtk1n87ydxCKhF+SpuDggEQlMcwm8PrqFbp
x2izMTo2gkFrUYKkrTj2/qIDW0GtLXhwWkYFIYwVeW7RMtt/6w/u3MxEUINSUZ3i
z84YUAHcMnNBm4mGN2K6wepIIE/vKlYjRzewTkySYfJnK9iMlxiyjUIuvSqvGMDP
R1HMUAMcb1DJRIGqP0K37JA+LYfPMHmQ6Je65DZJJttGoz+ynCm2naqz9J5VMx5z
dgREN4KFXLnPvH4wREAKrfOtQqjMg7hIKxz7lkxiiYFUyXZDq7DIQzE97t5oeZTZ
qAMrngy7mkrzbyczN+lEEM/4gFdeDHU+GahOniEx/V5RSZ9chwY11/lMdk97JcSU
YwTanK8P2xDrFTRHDWLOfcsJt12n6dlUNFMSaDnQI65DNrP4+vqhbJs3G9wzn/aH
7BiHj5wZHwEQmqbQ+hnkIiRvUK1soH29pSsRBMLFU+gKb98XQwHlzSdZF7xZcpXl
zvE0V+tpmEZau0weZknk8LaQxGCQK+WomGggYjemGAZAl4SddL+nrub82fbpINCM
sjNkmDeYWbOflQocn5oQ37oKTGcSM3wJ4e8iOD6b8fku9I49MUBY17d0NNXOXHx4
UNCTOUeVYC+w7tcS/MZkO28j19tDA5RAaj6SbB6x4Vc275fLLpGJWyyXFyCMlMzh
m04KMWVnR8V0VVhvwdZopL7r/JMDQPPbBtzJOvj6Tq7gTJWC4VP4mU/kDoHSek9T
lxO5gaePS88Oh7hIL/cFhD5peJW7xLlYOodTfzm7sivb1mlZ5D3zi5ka7uewBexk
Fi4ZVJZYfK5wVLjvJxDhlGKUmr7v8PsPBQrd7CVigZdyNPR3DHwnc812uqa8ZGY+
XiDOQOhLKGhc+4dsg/K21+wECmUFoGmbY0pS6gSEc+29KsyadWxJP0prOhk1O2ZU
5rg2ueRee6VFl6pTDJBwTTK9H0EHhy3TtMzvj3SZ+64q3xfh3uNz/3WGmVogJwT4
4F6qvEQOcqVDnV6EpRVrv1qEGUMLF13SwaaoMagYxXbw2jNGU8X1Kyz3fDyZPdTm
97u14D1h+kJp39YgtsBngoxscteWW1JCt+kaMMCLbZewepnr2nvYMuz9FNAvJStu
NycJA9j9oF9KR9E7cxUFHHXSdls3Mye9925p5VDqiwPDoCo1sfJIfqHN85LoBvKI
E5tUnWNLhxfYF3XvovYIHmMKUiEf69WbFfwrqAb91XPbL8jCk0Pi2n1e5m51xVzc
bv3REKFcwCBYIyISffUqYbpCjdEhxY1cekfKeY9LJa+H8F0+lGh2CHAfczM9C2Cj
C16elum/G7WpzZXiOHWika81B49ZaYFtLuC9wBMExQUCLKIaHPJGxaV73hiqqGPs
HoktAfTvUcy1jfjTUA6nip52WHPpgS3o6d0kgBq5r5JQMWDc84ER171ZTvtcl29i
EZTksc+KDwfXoVQXrbpn9MaB3Y/ylLXZU0kzooiK0SIyOofkpnq8iDCqVdu6lAIq
zCVG41jU/glaJZCynV/OHYkXzsEinKxHrkF6SNXTnF0CATbn+zH5TkUSJTAvzGEK
YQvGZ3xZAp66qcpESalBon67qu5lTXPIsXoq8hYeo0s5PA5uIzxkny2pjQEGtHIj
S29i+HWSXXSrRlZkACKCNPVRc4MNT5t2Av2VEzuLlWBrVg6O0XH14YSRfve6LLef
PQdOY6Z0DhkZC7MC/Pg7H2UTQxC4msYekezSDU72O8+9EQeead7RJ3ECgc0B5r4U
r2YRHXplHJdgmPlv+84CQcVN0xUG2V+fsSade5H6QcUQPfl884EaQ0o5gBrtEaec
Gs2KXbdmmTnEOqKnUtGMugnc3wkVdl0lFXRpRtYa3fIvaLMnDH9MsYOQtQ3a6M3b
ArMD3W0AGzcKI2vrNto9o3oUOV9eF8Yba32qud6OKi/cevp9ED3U0Q3iNJA1t007
BmFtUybznZ0W4wNwNSHHd8UkUkRFAX9FkHB4497r1WAHWZ2NbStyjJG2PiK7AddO
DeWEZQ8qB+735FbQv/OADDOh74V8pK5MLkCt/Rl5XdVZoUKSMxtXudRO/pyi9NJ0
cfXfrfWk8pG26ZMtX999S2RWCErwvgsfXePg+siDvwYO7gAdOPTkNP9zNUbxnOrh
xwMyP2CdDWWwc5cqRMNfH1abv/fWAP/hSPdXGe5qHLglSARhVZiMoGwdGioISTkt
ssQGOsAlxRV6gEVZcO6XyfUhLre3txQudbZv5mTN1LCqTmOqhPfO8+fe3XeWR5tj
YB6vv9NuJXxkz++jYgJQo1iI4XNmAf0YueMaFX17V0wJuoknc5c7SWwQnV869gfX
9g96onFkEe7cgbpwJnLVTSQPEawCzbGxOKyaRSP7/HZs/AOgOa+5F5+DcP4viyO6
iXv1fVgX50fcfU9oYmMQOK0cccQRnUW9arx/pChj0lqRwozManM//i66p7/v9GAR
klcrNv2l/rSCmUw0qu1kUeIcLwCJA9MzNtDKrwWpZu5G6sg443q5uiYkJprgLFzw
CawrAWCMCHEKstgjbRo+mHK+rdYbuf2m4STy7TTT5pzQnFs+iaqllY4jWDKocWvJ
ESx2OyXVkzwf8RhoN528idcCffvobISKtjbsnzyoRDLoOB2MEUN4pdNkt5VWT/2U
Or2gFh6dEe1Xx6o7ZFGtuDT60LCtBTPEK2Ps90XX7gBZBzHwZoBKHmGOkdkA0Bil
DiTna3xVOUJFPR/IoGxXBpAU/vLXTxGHOpebwcqm2xzhU1hvfTCVO8HFY7US2O5t
vSwCbM4aZ3793kQE0HaMEU9bhoAnSJC2b2hWy7S/NEYpV1HloOwPU9GprKJrPbLU
8EZnS5aXioV7UQNAtg6HOOV25gSryPDs3YbWrJNxyjTJ+YIr6EkIgoAt00LS7P3I
Z6gFBDO6or/vf2/isx9PCT3XhNULp59HBVDTybkJWwkriFtppHAwO73e6D0t8D3Z
k8kcN3/ENEAWhFm5FFcv/vHaQHRupQxOwS7BoJQtaoP0Zzy8MtbrFIosVP0MH315
xpdEoyPfafl4QY5QLZCbCxWjLmVGE3idfTyn4VXNqXoHZTMEsiTuXePgzUGVotlN
r12D+eGn+iZpNVU95I/tz3t3PyWY0sDwVctt7Hwl9snegCYcnwD9ddoddqB/1/Mj
SGVrfeV80TkLb18TksoxwSLasA6iNwYbh/q0ptxxMnrFZAX4y8l9AYtk5Dy1fnEh
EG7/MW4sZ35o4rrzfV/kGm+iq51QIFSaPD52VAx4BoD0yQqkT69QVxi7I4LGO0Gx
XpcHsnIL5dyNwXvX5dZeQ81L+fBGsmTTC51gu02sFK/r+LgyHVHVddZM7jjQWXVu
6AO8EVnCvF/mzOnVzmyrRyn1G2QcTbxk62/guxK7A+/7oAT3IDFU2gBGLfmlSoQJ
901roGxR1ipLBaa3d8sNeGn2ogMsNkgnAVqwIbTLFNNj66Mgaq8DhQW87HtLVK2N
ySkBnPS6ocD53tFtnlbtByTCmAVlO7RCQEd4y2iMuqsTEHGpfmPznafMzgcpk6Uh
ypffFuGl+Z9+FIlpfq34e+DeTxdB4uYgfnr+/d7Uc0FOnMHxCQ1EgE5GKmmFX3U3
xXsSbUht+0c16hyqeLNDRPWAaJr9MP8AVp+LStXU3NX/ITsCtHTHmFjA5AMjdB+I
HNcGvvFlOSLQB27Rnf9AcO8FSyinD8wB3DKV6cBE7yDZZIaumxopnOpOMyH1uUfS
drsZBCsAuY7MGmJWKE3XAEdWZiR4/PiVlJwBKyIeHWjE4pcqcqQBdDGiUDJRKjFr
RUTg/g8k+U0+R3QkoeiDJt/omWytHUDA9jB55gd96SBXCCEnkpAbI6ltsjo/I4AF
x4yzuwTeXtGwJxPKvTUL7Dz3lXZyO+UuEWLDjaQIrFLdrUBE+RoPZUpbDspaiGeA
hu0KxLdbMfnyTihbgFfsyUW1eVfNBoNGdL6JE7v3+sWf77yFM3MwRIJLsi1Qe+4U
ThtIvcLjdkwyY07uqy6IL5PBClAedtPjHRBD9PnqcZ4VqEzDi08buytdaZC4ZUc1
w163oMHbKGnIDhMFzRSKleLWCvEq47Xtpz3qBMWKLX5B8YAdRAcP7lhSEhKE1JEo
CBept+5d/rpVIVF7OET6UgyR36YsqHvN08RttlmazwtkgHqHNfNPEySwqVwZfddY
pZSXffrTarX/9Uc14El+7XJWS31T8IvJ2MYNHLsSDLce4a6tVX5c1eUOeN855b1P
K7J/2lje0golTvmM47Iph4IMOx/6e0RI5dIl582aAF4tpXpwiV9BV3mNM3KbxGw9
0hcNdKuoOcisVnwCRqQKGOYoyJt452jXm/LtA3bLEjT+1xv2u4RbyIw/WqaT9+S2
i7QuG4ZjLlkAIzNMpL7nx2YxqieOVUuFKb3OVvo9gJxetV7P8EZF78t6TUCgc8eh
h51ZqMmzxpqwdSfYIVKxlO0CjikZX9yBcXZVUODp1UqtrUPcxupAAl3n8vZIB4Qw
vFmCxl7PNVFh696/kXvAL1ZtBj24jQa3UqhjvLBdpe9S9xTIewqPkJYps4i8Zn+4
zwhViLsB5hseDQwv+sz6lzkcJ2EH4h+Qn6uamW16doKYgr7SaHXaU3HPj1ZcoI8c
NlSI2ffqmwn93dPau9rIljJfcML+MWvN9FqEbF+eLOsygss+r4315DXZQ9TfeRie
UvApoztvkw9KJqfwbvwkPOHwYpVJzihGda53vOM1hny8E+0OnqLzYGsfhIgPhLj3
354J5ZX5xD/dlisEE81q5wRuSxyYzde3P22owBRQn2qOt5DPMA5yh54rKJW3Kdcr
wVlKQhrIRFP+NTWiZ/AMo1j6quOtjgYjS7XuZkfaYvJyo1hu/+0s89m4iSTgWtge
4rFQIcfUH2Swophim9cshyOxvyTrhzBjr1MYsq6g3tg+OTaq5lROQJ1XK3RXjlpq
7KmGAzceZK6Q7rApB8Vu48Os71v8BNPaIIHRzN+HI7hvdARfBABD8KrVH+MtijWq
8ea4zDYpaDj0YCNnhV+IjhVr/XusxAFpDegXe8EXMa9x9GtoATi0n3pIOlMdfKsk
1hyvz13QA7yBUlEjPIw9EUgbDeJRaSDX/2GUB7pSsv43MfpMjCYclm2xQ0UudcLI
6SweZYd4DhyPYpVCE2rQ80TS8Vj4t0enFx945Rhc/9qOi2A74CmcvcaTWmDEUWMr
kre1be3WU73HdDVDCEnQ6YtRGPAtaROnuuZyF3UurQTJJn1jDnt22LKiVl65P1ou
5xj2ivANQbZbFaQw7MmDloftIum6kHU7tuF+xTutLFhXp9yFUbJFLC4frlR7riDm
UWCDUzUteDnI9f6/Ujsgn3k6CkOdKTAZYWvN3yFuskZwgbyVNsqmbHEPIiahFh2O
4e2bCwmFC4BZ66lxKNQj6wONLfCFdoU3L9tC4HxVWjRDodIbC0hp2KRJxa1xO8qQ
AiaYB2j+3f0U3YoIkb4ImfKQTbwSbb0PD5o+T1i6s0rvac4v6uzcIZ4JCNHCXopO
JurXWpiEfZUgcSwJkEQWg+mIQm7V44x8YHwCTUfwhVoyVwrGwVFK52cJge6r9L8h
ZnHz0ypERaAMz6xGBoXAe09HgLT/qBDGskSuoL5CPsfhWZbZF5ktyJvQsHYV6EkZ
35ANMdhMYZgShYfG0R0PMHoHQEntwEYRGkgerfkdXICOOisxI2IXb7rMljWYA3oZ
dGccCCxOqNLREYsdn+mXdijhwEzYCL47ft8HxPMaQ8I57jodqJ9lwjx9mFA/lIsu
k+7nnKe9jZikmH8SYCBZWtW284ySqVxYkM7VwP9lzvWe7vOnt2+EPmCYgHrTBAve
DEmnIm5cuedKe2mc1GAPDUSdKkkTB/iLNgBKkRLMZwyqI3fksOVkj5Q9bkSdAIUw
G6ImlxGdIA7V1DsuAhJHP8k1QB4ITXIvUWVQPgc6kD14xucgk34/JFB5Sc9fBmca
a1emYBI7JVGckXN/QlQfYOZxiRJQmQ2J2FWfNG6ahEryGQRI0AWv8n9OBwZZW19/
ez8ZIPmRum/byqiybU1m8TcglYhPhn/6vn9XYT1wBTzXC9JNJEjHUv3JVrWOpZ+g
zREkB4kShHdQg4nxWy2Ws4OEHOGv6s7AwCvRdbBKh4oI6yEqQDDjpuWlcCgbFiTD
oRqxi7ksV4rLkZ4b/jPYOvTYRUCMDEhpbLx0umRDn9t7kcUwVjyQzsDuK0c/TpYM
gAjqJXEECh/G1q5alr+FMS9UB638c6P8chHr5mIkBp2ZbmRLzYKVkqgB9UvA+a7m
azKi/6OxSY19GBD1ZUCxfS1zArchFOkkvdFuKXwNfYFaokm453//YAzNMC5mnnG4
9E4JK/Wj/BTXKajOyBPY1uJlOEANqdWbFNkSLSwx0JiQ7S6AnGHTO64e3ut4UyPW
EVzjMEGslhAXEOV5HgGnP3iTynqenyRUV3MLsuj/db3yu6IZ6YBj8islJCTK0R74
SHjKYOg0XLMzzbPgHFKXa3+S+ucj+7BobBBkVp3QcGiVv14pkTFRnrnP44MYwR+n
0stmlQR3S2nMq5lHnOdKkvPNJtOsfGn+NjmqT+h2UPUWsgLJkkAUAUelIDjlOz2y
XDEop61kWl2FRknpUb6ZTB8PSyHByD46GRhbIDjkzNVECVcofef8COfFr24L5p3N
nGW1pRqeeI1ymTbP6NgizhVsegFdr22sAbYTNPXPdzYOW6fKyWfs229Mhnh7w25A
tHHU+xTEO4COKF8mPH7oocGVxZOJfkUh8jU6In6SoWoCBWhO21PvsYzBjSgdcOLO
M/2SweEBFaGJHpDjn5EzNlZwvYviG1dOy61CcWvzBaSEUzfZwr4ZtF8HAoWgpiPV
CSpS0xFjn1zOF7aqN6SnyO0P42lkVyRAKe9Htb/LukxmR9Sck/uJd6YTeZAcgJp+
g+ZCdf/u7i3s9GCoG5fEk/UVUUkojtBwQHRLiGVVDFGsdWus0d9TcixxwxyxrogM
A5Pl8lmjfHq2dALy2RnbB4EB7juS1GaHHSQ6i3Zno6MgdEBoG6e8430yMPGuFZZK
3UlYg5DAh7bVJZ6a7oCqb6nsljfzR+EMa8B3tIO/gJrMLuLA2o495zHi+6U1e+9D
CKLA5y4AgiXI5q6Ln6gVIWIYn09wO3eSxNR34d+MDLlbGRVA4EqfvtqmF8EyYJ1a
0IGkVjTCJSBNQvoLEe2zzhOcfDciSsoJTqlfJGqVVt7QeoO5jYXQQGjpN15hl0U3
ZUb+GoqtZsXJFq9yTfSkMzI0FtdCjDIVuKQ0xD6N64/u6C+7koaJCRsOCC+J/mc2
oEjtATLcWGzHBKOJJOraIMhTsgvKupX+TlB10FNEdmSsGcj2wa7gi5Sj81SZwBCz
m4qeVrKa4GaNymMBezp/AGNYVmC3e7ftIHECg+wrhdJ7o9RKmKmRUGzLb1M04Gp0
oewsYHST5/vx/8HMHOIitfyRn0pxJlnST+L2OUoehNAmju7qzgfuIq9abb381FPQ
YidD2IuRPeOO39pQzh4XGOrujY5wgQyMF62qi/AsS54NicTWR+BSbko47m9w50H9
nR/sffiReFSdgW3NxaBhvaA6f/kAlO6CDM4yH1FY9SmyNRcOPJipEo5dwxGAua9W
VWCZHfKlZW5Y1jI5OTaZTpt6RucDDlniTyEr19KThYrp5uHNWspFpeMFqmn7MT9C
0V4XcUrXRRFwh8hs/va7gHCwAqe7UJPpkS9ctm3eaaZxcgMez6d3xFuZkEgm+uwY
3ZkzRVyo0bhLBTHHObHtAUSdb5g8jjPz4lSLblZ/QS9yU7chorg3uMMvPoQKcCLl
Em4SrCsQnOTFLCDlpTYjW4SdWi5hs82pc5rSF4b5ltHHv3N7e4zTf/UBTQ6SU3a5
ZwF8iQOrCvPZSZ+CNctMm/NtH+l7v5fsL/ALAGN7All+Ksj4ulPnW81CVR1D8EHN
IJ78zCAWx+3+MPiyqEqpzQA5rC4+u6fnox4UtT2QR6XwFqSmsGcgpxctDnmautYt
Zi/cRcWRLaQOwM3h7ukYIBP4pGAypNJCUlPNtIZNeUd6LtNP3ivWeJKkgJvjKH6q
/UBIx4CLQHmLw4VqlPFxOPVQFi2M0M/4CyoTq9/s/BeItay1pLd4rXNJ/jDqNgxn
9sV25KIws17UOykY02QIuvnp9n47HDOHssGhDqhZ8SwABe4yYBFpL7FjfbJ3bQyp
CCOf+L9QDQA3vEa+dAYfkUhxab3KJYIYjV6wPp+egOe376LgE6bNROIg4p3S1w/E
9Eh1m/nQTr/fTwz5DoFXXZ1M2C6HgRYkaXSP4ZWJ3w/JMoNt9ohVpB0uMJYs5wHs
fVTECuVs7RUdnPtfIXmth/e7lvjyKAn60/pWMuoEGNVrAzFCZ/wfUzdM9KlFf5ze
WPZIaK/UpvFHtDDoisT4huzE5ZiZuFGHGQSvwNX+uDbZDWotBR/gf/F4Uzf9metf
xtdsZrGbNoblZqQr9k/C1PdJv5AfQDt0KVjg/645ias86R8BCgCWFuQUCwvbDhxt
Uaq70S410FEkk5btIv9R9z/qaHoOPIhPofpenoZaFK2SASvPojmFy9Fvky0PVZEs
R/RzuMcrNpw3ZqZP7iK+9uAlu3y4XYJ2VIa1K+IIbFPrzzJGtms1R4hJHY1AGGrC
ggbXlK7ICas+ZvT7SHVIWCASHBrLXmTVD97VsWaC2O7fMTRnsT56UaLQZ3FgRGji
etjVnslWVRlUJm7+OhBMHvwBwHR6usnGD342Gky3kjgcwMIPdKTeDve58O850e/K
+EePaF7xNU97wx8LpmIFW2LtKIAbcWERBDLcG7VWbRHUmiPrldNDq9sBeWaFBokC
nmjJ+zhwzsaV59yvw5q2KrxesIH/XoWwx9jWTwbgEHDve5rTiF7Sj5ne73uA79FG
PcXqhiLP5lg8U8LTi2O6I9Dj3AL+/No8ru5X8Y/bFS6y2jz6lk6tJq8KHnduZkc9
VtWpDM4c/q9OQiPYRUihhm40HONh3YD+4ujcNYxNtPr2X45fsRv4smFkq69SkuHK
5qgm025elb7KvdVAbcresDsw/GLjIPfJvENnjSHuuKgpBO8QkXABS335kU2bzSxK
bhBdo8mLoImumZdx7Igwuw0WzqsFx8feup4WWdtnCI6Lg8lbkBaZfxHNYtMmLbz6
TCRMcn/AgXZYAvY04o4WF5KIH9Rony84t4vyZetclIJ/tYwbBktMmPjyHL5TCIbP
K5f95XwlIFTOHLJ0dwh1HcoTb6CKQ7njHX/Duyy7yAvQLbyxL+lbO7fwKB14xMy0
1yDMt9bYoU8PInGcg2I0WfmlFPRcq10eiV/UQN1fb66QkaGY+ByurUThGITWIEOO
AnVRVecArrDcCyGaCHxBs+WQ6h1a7qdUeXBt4YdGfIgQ+4UvWz/pAISHLkpLaTzn
0p81iE7S/kVimrfNEIkuUtyafC5KAjFiQH65S93a+dbaf28XAUcNe1wTor51Qt00
2od1YICnhXwgVMk6W21DXjon7qpC4dO/077F5/pHYaHvhHUWRe/EG3SW95MRA3IZ
plMlLeRvXvlP0CJSoO7rcCdY11tISTfXMX3uWlgAEO7AS88lJuaQCiD+1Z45cZUD
LNze9OtObPTa9/iNNsRaO48KRwgvb4/0neTJH7Ez8jB0xvfnVPucHkIe/WQdpFta
tszm2du0BTFcNrgCkuAuY4marpWHuo2xyOqZTfkWhGEN3hKmWPQfduF24tdaNKVk
0CvQczazVT4mfPYNTj50mwrvAayh3xORFp4SGHod8H3vfujygmKSjjr1zAsNca+z
WkOj5Xz/X3RidzXveXekoT9NkhXVingtCVJt74/NZZv8PpsettrGIXMFhdkPjnAd
NQbvXkc2NV6eME2ZuDY6SyeNgCietPg2eSI0y3U79UVjTtAjKtyM28xN8o3d4LvD
cNY2w8bhGw1TmTainaL3XEnalE/8b6JXg5S8/TmBDPAq+63nfvRDGs3G7y8dxoYF
1mPMJAy3VggTFgRBAvaNjUfSz3e7Sq42WAvMUMeq0fFISRk3SDlrvoRrbC+XRUGw
3jvius29+3MasUBnspov6Q+FTyyNYMlc0SV4F+cvsWczAYv5q093upQWy9LfxA3b
gvWvZNChPqHrrmz3Nc4il1C4QgirKRpgdjI0H+tHraN0kj+cTna1QNlQPZPLwE5v
mx8y9MF5CqS1fmtWURRzpmoFyvo0C1+P4p//qQNNsdi3HD8yLe/uMQVim3H3bQ2E
AEDGL6lB2C4pg+3GXdd1feB6GhdhvHZrRM2wM4NRgAym0Wtn8PV9eaOT6mkQuGol
SIplnDO+KeabJvjaCtM5mciTP4NPfn8e1UTPGgcBR0ByCWIaxOD4ClP5DbC5V8Ol
3/2jJqeiAT+mt2crfgJA/Gh3qDhofIMznedrvuXpxcK0iulpxbiuMMGfS8iZ9q8d
SB+9GlkNo78ozV0/pQ1+EwUA886/6OOfplSPodHca6oKlkbRxvXbQHl/fsig+FN3
5SmO66Ez/zKiOTEaPyyJPQEuZst5CMqEuMbnI8J4ALZz4emsZLVfJgHjHzXYrWvG
wXQppN2vpv+VImxExtvDLHYgMoA/usg88kO7fQGBNpQPYKzN8f9j/V/aNTeFbL3B
K9PzUjdbEMkSyYS0nh4whv7KPX8ZS8CVfAxcqLeTISos5Fs1tBc2t9317O6GZ3lU
/wbJmETemj1ZHpSERmaNoQBe6l8z55gEGBfWaVVXH0bjuKrlyT8FAdHIVvSDnQdj
R897v42poO1wrS7cyFq2k+k3OKfnFmPUWMgcQopTXA3Hjjjs3eGAB+fzSSjyAz4Z
GqSFvbbqCtcHMymNHmTxhp+UI/KThRXYvALBuwD+t7RnunyCspJXTjaAqhhbNZjZ
qcUtrMxlrhCdbjvB7kkhh5D6i9yVErlkCxP9I+mkNgX130BMyeF4yqX/Ft8ld1tW
0J6TmGInodhhoVooBkrk1nzXljowov01K/9abW1RJg0SACiVLrvbjcf+jx6Q7k6U
myMYiHXyBFvm41Yr6M/N2jEMK9aywMcRt66B4ZzlYYUwUseQGF7W1ZBgQFdmls61
pd2Sgmp2d3Ih504X4SS6VN25nE88imZkABHPP5XbJLFzWOrZAUReA8b4600C/HOF
QnfdyQ3DDNuIAkPqE1q5R+S8i1oSQcfKt9zhAsmJm+EqObX0WgDatuPAYpT/sd39
GtwyppIbUOQVMFwD8B7urpv4iAptH5ynKOrqcQMygPDPePcwyDYkLlJenZgsNk/U
DFA9BLbz+aT2f3Rn3pwv95nNZMEQriZj4Ha8rJt47ASzYC4zQv5+ubtq8ZW/ZKf0
wyP9BRl5mnR/FNjEt+x2viCAoMhVA/uyQIK0fUof8jCSbQi5ZGvTzrJ5AjVNorsF
Sb/0mHHCeumJLQjcZqKJdsvuVh6T6AROIds6XVBmX1MgYHbzehoabqmUQdLHySQx
B4SpZsezmtZdGgkIIsYO05vvseeTVZxa/j1nKkmzIoT3Z0HFBqdJHuKuPmTBa4HZ
2UuoGdvLWHTAXYGWa3Dn//6+vDr0q4AJl5mPZYHBbt8k0Nz1KueB+Cg1wVyXxcfD
FbmwxVIBt54kYQMHokcZnDHDJAedqkzt3rEZODPYmM9Pogi0FSIiWZRPhVvXurny
RB71eTjK3E5EZY4fdMzbGsWjvuLQDo2Q7pOWmMsGpj4EViHS1bKARwQcdGrvtnoW
8qxA7vY0Y+e+O9rbhdAUU7ITq/9CqByKAVNJfX0bs0GW+vdJQNfGuru8GFHQw3CF
Jzv9JYDN1RjWmeAdjU43ksYt4rI+otsRhNJn7Tzsq5r9GjwEeiJ5Z70nDM5A3c2h
mvRHIxXytIKTyqQfWR33qSavFC/BMladK1CM5YOKN7xQgw78YhMbjFDdFSnhKqfa
k3nQfh6VoUDvFTeB/yjxdSP9164dsSpF6FBGQOJymBZMhlNg/NRhzVF2C9Mbs5Sg
WO+3PGqPNpOho7JcBO7kN500f18mIyuhPRCtbkzgQzGjHzgoGRFJK5+Qfvr2EH2o
L85mE6aVg1DM5LMMO9sF9nPYChovf6OTn6e3OA8LDGpVz3uzg2/MKpVocyp0rBdd
/c6roUKg99o1MrT+nQDJSUiDqtq2UXnkPy2BOQdLg7hzQS2mp56LW7MnfEsgpbbP
QDpOVwvEWTP0A5STTlBCfzSwN0J7i5Vx/ntrad4ZosBnCnukC9lX+SByjF1esVNV
JGvXqEMftSFpWWL9s4HRBBf5gXQoy8PgjpZtA3eIWS/X2qNUTA6kI34/QkVXbkDn
Apsm/O4QYsWrwt7NEpPhAg9HJ3keL7ZXsfEBIUivXTMbocTbk1JX2bs5xpcSILyj
zkS0mrG2gpQolCfWTAY5nWEaebijiuNO5CI2TJgP+2gDUsqAPCbeXX9lXaNlRmj3
/UkZ529WoGGeBnqGoj0Z1pNPSxX+Uxv03v0TOK/TaBZusfzpu8PtF3vXlq04leZA
Txawt6OPyNcGoVFh1oi1RDtpw/kQt+vaBM3s4IiPzQ3kw9dcHpfy/xd9LJBym70P
oLG9tpIGNJnFFyBdvtlVfkSNJfa3UynDfSTTKqoZzmBuhtxu9grUGrAvXkW3Ns3i
LKDpA3l5OLmy6ougXHbpxxjduBJ/IxwLZXHM3lKIE/NpW5KWyQlvdurMMzI2NaJy
ybSwOT1R63iSr/czzRLqp2WxiZgo5zYVvAQD0BILuNPRHKf1jFcBvR74oE5WRj7c
M8TPutt3RtR3Ity8QjdbTj8J1EUXVLYk648fWtKCM0gQLsZOH/6UnTVS6zKIbyWI
vjD6qEzv529U/SfvizvDxfEvc72do2odXjlc9P0/DJIzGzEkH9f7HN0GW5srqfh4
cRJo7dUJ8rK419dOUNA9fZFEq/YB+XyA4bJ1HDLCM+jN0GjzFTEwlLpzbkg8aAe3
lc1bM0N4B8jajcS2ptx4FnEzKEDg61cD3uvOOhbdGYVm+AYXgZbV17bRKxwVK5Wd
kguBOy0b8ZLZABHWi7Rrtgf7L0CADDq7Mg+qfAdfN+9BO+DRldPyJy+hfqu9tGAB
SY4H0o35cL0OzmPQJf3Ue9clAB6O/vQWMsFuT+hWTi2g5QBa+YetwfP+Gu4i5c73
0UkR3IrzcnElxXyw1+7Kfkv809YoXN02LfW1NHC86cIZkB72DSgMoj52qxpDkR82
uGqZfOX9O/t347fuVAKUxgPHMHjjPcXCagI6sHnw+3fANV9UlySyR5E23xq3rL3W
Y6xo/89znf/UyONHliGSXhuDWiH+AfujtjyGAmEajeqSpo3FbOyMgBBt8ONuq4r6
+usrPyjfa75vzrap5FPBzasEh3dtbl11s/tbksZDaY0cIrELgVZe4tQHbXJKiy2b
hKiMNG72fc1mL5jagxkeicz9AfRONb1EcLo70Xgl4BDc6EmNQrolsC9PMs4gSZ9A
ThGwZdOV+ebgd6kl0wAgkv8l0dInhO7iVq7l5yRG4zlAIC+Ht0zrmgU2//iP81fp
LCgfj9YNkHfWVAmk6mrMpPbqrcSrD2yt5U62dHoCbkVl+Tzn14jaLLlgewcQPxnl
799gR0UhjyuPjcja0ITnWjRni/H+tkagViCWYXC7pcgnXgxY5Alx029Jgy4phkvf
Ag9UYHNCmX0ScO8pklITE3zoU0MOlBhZEWD7+Ac+k4HtPmLknBQBJQ/Ke8tiyjpn
7lzMKUXwSpMaVOg+3JcU0SeR6pmXukCUNDslBf1yjjXF0wcw1jI7iFMYtZIe7H0b
oV5nbcR0xd70vTeQ1HAlkqvA1D6565vZzbt2Tk1DlPfU2Yl/dXgVPktCgkaZLIYc
fqjvdCAvPPN5FowHhQujy3VvUSxwUZRS90JODNfoJsmqE/WGg0suKXM0qvIK45BO
tyNZuumHrIhMcjbU+IxYtqIS2jCKGzMAPfXGpluX5AKsuYNnVpEaPOMraTUNnbW0
C5ikt9YzZKKGe1nrN2hMetcc5M1aPfj3WApAjlnKZhcFGwoEkdtdEuEusj8lwRII
Rt46e684QK2+EZw80hFkyJ1m/bqkLyEdLDmS34pbiT3RXFJ92x9dqXKuy7Ymm/81
Yg4PsWuHHDN/oFNCwImqLQYYy9uIufJRh69bV8RbbfpeBOnUzFus8IlOdie/rzsr
HBekbgjp29Z/toaVhyofilTrreKJHxvCgAanMzH+tUXZFDrZN+I2ABLaLHJeREM8
/m1jEQW402jazWBvMr3pOTS79+cq3Ah3FMj53HiKB2dxWZiw/iRnGuv7kdDOpAmc
yZfXqnhFeE/VFM3bGwPLzeQ0WX5VMz0j5YF30ZiDmhrcGAGL8Xj4KuL+uhHqJ2EG
MRvMTNhgGg44VWF+zANtSkRZS5OBk4En+fJgVkady/YWG5QTtHV9/PPpxOApBh6U
JOtc6qf9JlJeZmiK4LXvxrUBfHmejznR5CRMoFiR0EhhWHwQgGcDMsVrjFg+kCoN
C3C/knDOxNnSNp0Z4kv8PcOhscsg8xLlDKivRIk1ngR4P0UBAWgLP8uDAHab+OUG
DT3CuqZVZCt39img82bNEHh+7PFKUMCWO5r2JrkJpU/WQx18cxIAvdsWR0GmXcGd
zhy776wKJtf2KQoalW5ieSyOoozgRHWBBwdfurtr8ClEyituD6XEhVAsu2X1JP0G
OR5RKtb+vH4Rtpr2r3pHMePUp6A7AqaN5TYMq/or+TM8Gux0TMKMtyh6qklWsyRM
EF9jJFS7C906QEN7WVTgtz2Xe3jLR47CAZMr4yFwmhmo7kaQjEY+i7GXg/Cs62rp
t+w8t7xKbZ92zI2LnA0tk3Xd7WKn8X7MqpmOXuCR8X4QxEhpn4BUIWuCqdDeHfAt
YtVdnHNNif1QVAPkw0gxPcV6mEfSvVG1/LxWRb9cIMvoIkSWznLkXibI0LDce3tz
+Whu+ZBQDTMK/wZSjcd5aUsCCp3rrNaffrV6GkcyRcT/vlW21pYISvg7HVsQGVbZ
SeVl/q0piJ219/Pw/U2OdDeWA3PZJN+JzswRsQSNjOLTbQBsaFcC9uTVHK6AWcUV
ygkZ/EeHPHSxMxb6ZvZLPZjSHKQL0hSTsFGotASabqR+ExhFp0mqO2FVUzXryC3X
bb9ObHyH+ZOHWs4w5N+Zqea6vJkV4btBFtx0ppghjlpMU0a+ZH7yfiWaKVknzHA8
TiLPc+W0may4WEp5SKGdKhyMosJXACnkY/e4l395tLcayC9wFqNdaKgWIPANUvZm
he67SPRTUWqHaDPkoehjRH9s1tFz4uh8ujaXQP5oe/o2lJr/11ONgaeJRtcSmNGQ
vLKnN7UgR1EjjR47tA3Uytyr4iQRXPcg+ifdMVGTaPm9r3YOxxlJLtNYL1s3Vskp
Vs7YeLcPOhVpOPcTdouR4ayHWHQU3UcXfeE2RfgkpSRPOyG9fz/77749JC/qAdhI
nXJ5cN4/VEZDvNlyAwgpYPYn8XD9KTOLpaBDvOTC0ZDpAUzxvNT/BYJlumVdEsij
7pKo/Uc39HApg2DWbDotR9ZX/I1/0KffUoa+fDtAlK38psat4Yo98TwE2P+Py85S
wMkaLome5aHWruIIAHdyJ11m42Icqxvv9YuHbt4kqOVwAXw/rXIbjxDh2kvjyPH9
gR3wM15UM7xUb413R1O/b/WKqCqS1jqoXutDlKgmOCkLCndBuWnFd/n/W4MznZ3c
0u7bDznutXSSNAUeFDnsAcGSmrQB1EDXzk35Kvb+8LG/KMuIC5+8buDaYjUWeg9X
q8UtugLrKBjlVEcHCOj3lgcjD/Ui4+D5g3QbXWTgHQluRDEUQwXYr3DJkb6FCRrh
WYGwchTcwAdFn99PaDaG8xIPeTo9nSdN66n1gtmASP3wJd0c2/sP6bLxVJMK2v7W
T77uKFuM0NjJnWPD784fueLutPHqyZARcZWGK1In+TplAvHGM/XhtXHtk9VLWW4B
NCz0Uzrv0ISJK198iSxcahaeNZgVOueaFQGhpsNrDUw5efxw3UjMWez3qipVxD0D
wwQQJWXWDQTHQg1Vt7noGdO2DO/w9TakQUqreJO4xSjpUohK0h6JmubVnXv0+Mon
cdueHBgP311vhgQtpNQY/6BeyDHl/PtwH4yJgMBWhM5Nv+kUqlPsNReVO5iu8ttp
YJZuYALfUqX8CYJOiJMEe6OZwHXgJJ91IgO9Y1WLp3WIpica+JJAzwb/BuqW5dSC
g7XJqDUZ3QdhA4ZrnQsDz6T37DSxpFtIQ7wAigTaxWED56J5yJKq+nAMPYaFHaO5
+29kxJhpIMwaIqqAAny/QmTCqZNykzpWQCQCeUpxTn/4awEROD9MTOx8ZxmI3gsB
jMg3hrr92rPUTdE/AdyNil/qz/mytl6nSgubNauGVshWW+yabGfsnbKAnIktmCor
9F+3OYzOCZnCxtR2i1jhvkS7V2d1tlEqr50sUHhBmxgh4UIL3MmtsymH9eLPyaNe
nirPyrSl579LWE3dttIMPgdiwkwvCJIPAWDwpdn5pVcsEqAVuZnWYGOuUp4q3tRA
+MLzB6PGRO1s1ZQA44ycN+dbHipf62tVh+SiAvEb0NA/MYc/SLHpi6o3g9tqn0OH
6qENqaTcjt8mxKRednbsro8LIu2fdTEcmv8pxckHnlyZFm5KsulnQ3SRiXvmEq49
J+7RAKTDzS3j1xwtdOe+YRIrc+3XIiImwHfZhVpMImTQ+ooVYEQJgMTHsVs5+sn3
5eKEuheNVLI1i590YXIkCjlo0NZGLbicPoY42XQeWFbtI7E2BVcorHN1MRWIcOTw
WqG4akfnMJ8BlllpfcFg70g6EF/3CuadHkTaCSaCggzGxD75Hyr0JnZwoJ0lVV2I
XcoU0prkWiqhGOouk3/hXW+NIcdX8lfKynG5CP7F/yMKtdJHCAS5ribusJg8ujRW
Sn5W5pd2MZdmBWrG9MhugdBO1lRvlc01Y1y22XuSxhKmpWCPrAYH1flHoAlnH3nl
T+IoRdD8RTFAxUqjDrbRAOpit/F/l9yuzu/haX6Gsu0wd4LN2vWrViELJAg60PlK
pvK62OFMHqF1E5KryZZiHQ6plDKRRP9GPH8wJxZtuQfmaZ4Gb0u2qrrpcxkWYmON
fDx/Yqnns9KraQOp1fgYFLGE7N2jq2A2qW3iyplD8Jl4EEtfM433ywsQ7DgIe/3N
tDF5KGPJmuEnOmwm1VQ3Ax7O+mIeIgBuXhsjvgcZcJ2AGmox/7d1YB3eoNZIaYOT
lyCgYDUb9V4eSgE090X3Q3SWBjfxau0adj7eQSjizSqzI+pHzoa2Gja3YA7LvHEF
7vKw0Bqz6P22IQGe7+Lim4s/js7nhLNLhGrFHxbxbQCzCqj2d6ot516f8jDTXXOj
SrLFknVofslccrcj7o9ofKjDbN3Lwm5N7cLHH8z7JjF7BsGUM5GjkSLEOHnDD9JZ
vZwpMh1SuzTH67l9PHYj7vSK8z/Kos26qTXrYIv6rFd+a53t08wtXM5Mn/DtWQPh
D24jaeJoUfgfNhRCormS9UHyoYM6Jjk9sBbmy/Qzzu/5aKc6r8oKQz76kcddQm4l
ZWsO1lrMc+vq1j1yW3EnROvrFZDD+kt4G5mq/g2lwypOy1UOxMbZJK+IPpr8lfUA
TCdTQwTMMCy1VJxfuBAkL29rfPwYAuDVDv7UaTqHw70VfljXFfsZh3cKESCchnu9
bQj+5q+vTGUU4dZUi3OmF6jG2AbDycqynTGY/rwGHQgZp/bzWjJoSWS6s+yIXrAz
Y1l3tD0t1NIBEtpWxht3kXeIe+X1opQiRVZy6zNqAGrfKW7rG4bhjP1i9Ninderv
8DcVitPvxdytFcRIcxsLjcN0b5+QU2RBJxHg2ilBTeBaj7DH0BXZTPcVUdR5tLOq
oVzt09fsKTmcAXb+OPdcUO9PxfSo3sSZgUKZxTJ/8dP3B3rid1DgPXVEK8vhPC2S
weK0YOgzdP170esmE5b4SrMX76lGisl1KiFOJM3Mv9Hurik3hmOwoAw4jWEgmxxc
hYXlesGZFsoc4GWmUh4FphF6ogoGQ6FOLA0p5Sv/37plS4gyCWQ5oixFqTMAQ5QU
NwGDLtfp5w247lFjuBFDn0kf423DS0wfMF9RAIU0Oho4TGSlyBnpfAIb5qPZpGx5
mJQG1o21kuGXYdfxL/KiBZgZIttLHd2KsjmaxLtwDDEoTsEuvGRtcdk9oF6csP8T
rRFS0b0hzrZYdlXEq9bNaHX12TYPv0XV8K8NV2DauKdo30Vtn6TzznQoi45QiWcD
NqlXwBjL+DCi0p6wk6XinVjO+5LqNmieDnCg+mNS4us8SFKdR/O8NRgzvtdFmEQh
tIAFoxYqaP0dEAchBUhKznjgnwHXUHAuVpt9Mn0P7fgPjoYo0povrgrRENkSG06d
IMP/UMykPKsHRAd7ss/sGdlfqqfcDDyXnzNWLYu3y5GQCZNylL8akdEQrOA3ReUW
VPfMckfUFOF0AUSQrH2SiMRgXBHEuEYTIId/4o0cWmLCYXwEfzR0CIBfFDkuzAh6
Eo6e1i1KYGF045BZZPXu2KU1DG2v86nOFp23ZyEIiQlfGrdYpJUaLSgMubwJ9bVt
TsJInRPBQhw3gdNT4IkXYRIcEU+vksZRwcMGj275rM8VBGSwW07zuTstoe+D2Uaa
QRioZ04gzkXf25hDOOW5myMAl+8zs0jkNAUV4p1CDTZFlf/dMkhFyVwTCkcMNnGU
9HX8ujr25k2tgR4NtG9j9yoCKTed4BTXYzaEZDIFEYjO+nRj6iO4jAestsEIPJen
qpnMHYMC+Q7I/xdx9DVAZqlSF4tZpmZxD3sdgAzEf4ua8sZYf/Azv93roQZ21OPL
lkHfY8vCZin/nx1WMXYAbQX0Kfd1XCFsCEnpuuKZIgNKD9t3N/EUyv5nYilHP3kR
XhhTlHxIoMsvnSG8wiY49/PaKyJO4i3Exef8wtTtVPAePQQePpMtFa388pFQX+Nk
JE3wG98lCjuipRv3FWuMfqpdM5MuGJhuAlbKX6Fobd4FqIV/8y4GIJWsDkw1pD8z
NEeSR0iSjb9JMCoVechcIF/ZwQamyqHrLDGWoH1krxG4Gflet0QpC5zICr+9rqpN
EU2r400UbfLQZkfAIqlqVpVsQM3Z3hk+L53h/t0qQ/jJTCQUtvFduODbvWseIWQZ
2P1zm+vG+5R9IDsnEL19tYJZpcuNn4g1Sa19Q0n8XOvgxjWsWke4KMYl0cSUimnj
1lLWWDd/Vy3NEFrcxReqShQJPNXRVRdegm0j52zqliVj+c9+l95rM/Jvzit4duO2
vYfCOfKulcrv888Hfa+3LTUYHS627oUBtjnZ4XnYVpXIWFf0QSi3VFMA4OzBOx9k
dnA7gtIbRH7vn/HTncAZP26QgkPYxcUfjcpaPPBE/w7kGqj+Vs+4bBfhKjQYaIgc
YyxIb7fszVImX41haFdOIpR6P8KtBMACCXzVPcKH/Z87PQgU2j1yyDk/YxUPG22T
b4oxly8ZqHGhBIGPwqFeWZCDegi8Pt1/bgteqIlYiMpJq50goOMqSBXiVXcMAeRl
paxkxWnPcYClq75QoMTUpso+WI5bKUl+ML2KO1oZLkXoIaIIxZLC+aWTOSOrSPzH
uk1c4T2ngWGu2f6LVYSKCRXMQ1tHR5uXUpjEaZ4bTPpCT8ReFwnl6L43dP5IJBW7
D29g6nVwAKvE1k+zbVCT2XCgJAjQj/RvAcl5TT+6cND3wnuJX7TIvVx8etUHRMFi
HJmazGQrTkXciFyYVQK98MIu6N7qiwI1wkAnQ3Q5bi3NH5HSHXWuH1bhM8gkWQgu
gAde54HCqG7YTgqxXSQmd3N7+26nZ4vyDQNXnc2Ix6MaGxL2JE+T4TPaKOwmpWdr
0kWA1BA7McyCuVvXQHo8FNeEBZi5nfatLkk00/KfrwhcF8OVMLz2qzLAE27qObJt
QzoxE7VLrgUXgW1jTpDi0bKTQLXoEuowWMof0uAOxE2PSR/ijVFuvvzf+7MNpJib
cFeY6o7awDvZrDN2myimmuo025r+jJQNf03ttsSeUcWknaYqmx+6WQ4hYUAgf3rP
iucOrSzrT9XFb6+OTj3qghITo+OOC61dTYDpAzgGWxBND8TrUj5/3Tro4gTocXA2
Cqu0EPNsjKSuVTQRZH4ULOuYoWf/x0EtlG5Z/8I0Ehhc2gDCMhWSRLPs9xWXGuRG
6lpQl0poNJaC4eJ5TRNUdiuE/aSakLzX/Dz0DKUbtYZK7k9GcIWXu0hRdJeSS9Qc
cKRwLlT5KKhU89yBRJs7QKj93I4klh5On3RKeX5C0bYViu1UvGitdfFwsVsYlCOZ
3CbP8p7Bg8Lb+67y6AdBnrcQsxCcPMMGUzds0OXJzeMtx/oIIBSa4PyKgN+ijWx7
mmL/+Pjos2f8CGixG/IYXNt43olWKnGXb8ggFvgf9kqauAs90ad+99GD6F11Tv9Z
ByNYYABffwmgGhDvsIDeu72rHCOm+S4rlfS4PNkf9ucAbgXQrEu3In/FSTsC3ScQ
RVleMuoyOg0cmjVBhaiEMHTRfkbkJJcP+SWp8Zs472rPudHl6jLyDgZ3D5Jl24fh
d5WetyXlkaBXfVk/J5dEwn78/G+gYYHw2t55O/MU9WjlKgwuJPt+86+aUJl7s43E
L0zDBuH3oz6dJxtC23+1QndDg9iJgSyxrAelS7/aF75JwpafWDocIyiZObX+yu2f
Xjb1nWkqztTejtXNNUjioiBYI+wKbcSa9RW2xZ4oXhQ1GTcT3eKvE2qiiecjm3mM
K8D3ifHd+vz2jPz1TowRHG5NSVSOJzyPUCu+qXEsC0iFbWX63r3zeS+U/ZNpxT7V
vVwfcB7hTSuFQJZcqhA52kUkClVqNxLdGsQuUt1BWYbWdLitFudAGxYJPxqvZ8sy
c/6B8iXhNpjimMEf4pOdgXCbHjhz6DJKD2Kv/RdjoDgMEjfOc+CpcygrE+OU5FCf
fY+gm8Vv5xYpJ4aA6Bbd7ms4l3HOtXmHY63iGgIudcMm/oByqwoG3EI7Y5Xx9nDn
4NVzPWezD5D9ok6YJsEDy1VLqv14FC8kQnjR8HmD03akQL9OeiyW6yL4ZREyfUpA
2YBmTdi+wQMoWzfxAg0Dh/Jv6s9qQnfIry5RhcyTBvlOMpznMxcfK5peVR/3O8mY
G+bB+jNxiXDG/36MPyfcy2U6gPeqL+A0LkAvtfT0qDhpZ5EWcelITJ87QsyNQlKV
3GJi7JbQFXwKWyjInatfSqwfjdp7DwqmUacUSkiLXjOat5qHVn15EqPFjgi3PYuN
0ItTgLyFx/s/pTTSNsehccLRVY6/Qdh+HZTSEVkM2QUvl7gLR5FMcQW3SadzEmB5
ABJC9S0KTUm4IE4/IzgYZJ4XWtHTB4n7dnB0WV2QscaYya2KNe9aoajlEM9TFMID
i3auU9DcCx0DeaplAo6N3KGxokk7FhbxnZszbbgXPD9V+nexmFhrgR120eVLoFUX
DLOXCq69YuK4SSf59DzvkDd9IDB7jYqQnux4Swvb/w/s5lJbSkRS89UBkmYtbZha
HsCwAfaumhjSzIWW13mMN8vPXfqxD9Vmapm9HZjPKcCQwC/IxkBjGGCOYMUdgsRa
zOcNecmbLJlbC4Tu/MUuREaIYefc8F7VGoORKLwqH9s0YcA+Bm4ygGEHDR3cJCVk
ZDnDN7kggEFKmLkqlREFDTHeAU5Ov/lRAdgJLCU9JzfhLgo9aZjbMs06uG3/OP1d
ojgNiBOXyVyLK1EqbLMCvC54pXyNDhcRrZWOyNunFE6SL4U7rs6e1w6SI+YrAlKz
rE3aIP7jxvZs+u1oBWX0DQtuSk13oV4ioOWDDWTJLy54+PjwOHXNycTByprDnTFw
XXV50bIzneDZNG5RHTBNQviFyhYnUhYhcG34v59DFmJsfZ351u1xTtKsjqT25e0x
tmkShcuVi1Jmr9fOWHs1Lfxw2+gfzuI+c0/lV0JT72HjY3U2v3gyxMiiskFTUZlf
ocDcBOwh+QpyBsUbI7C/T6OKeJRFsiyBrt3H95deL7vVAzGaDKpG4gFAJvLLPIX8
m7a/MMDWXGFlJP2gGRA/VF2a3tLpUteAFxNxRoFjF+Dix8nQNhEoqlWyHl0aX6AV
j8QnAeijsZtp/fmQ8yG/2j0VqUeppyoGOiXxmxbMbsfaUZmb9fWLDz62E6ksXoO4
rpU2NtZyp6xzvh4PhhGV8iaOCt4gDUXw+F3PVCQLdiAFC97q7SJPBQXlceErKAPy
ApveeOx0uWyHp5LUCznkhPjwHIgJ7GBUSNNR2a9EuoqtdLjAAcqj54WdBRV3FSlS
fYPuMrdgwvSORanGTj9O4msDlvZlNDRL14nZKzi+ATp05uDXtwNtRoG3LCUhPUIR
togMdtdHGJEjbksO6w5ilg3x2ORT2Md5dAZJVvIGEPSwB69jPTrfiVjvmUE645B9
pn1WebcR4ySi0kZLR/xFQB+5Tw8jERDxhzgcsOUd/YrrbO9Lm96V27acsUxGcML2
64ZpKHd9Sp5fqKXFdUf2PCyTM3Vi3Q+MrnjhuuqcaWuY5doOGme93zogJ/fprTYL
hHmKAPDJ2xg+XzH9PBOWW5W6YiL8411lyxm9oTXq6e2WXIHeMwegn0xIoyiWYTEw
4QlVDAh9TAawnPZRxXbD5BM5+m/gQFTqBLSpcNcuj2WhGIlo68+SIboEAHcannEa
rXG9UybHfZsOi0K7DldNZIeCYr+l0m1vBYrIlhAjBk1gyl4gylbuSBh8taLrqVmX
6p4hUtTp6ZdupYRIunz3nGKaPG+kxs/zBErZlY3VFFQiq00ut5cdAgtvvphBPC54
zBPbD41dG1U+g/FDYRCpuYi3BewCpjdfO5RaNHs6VPOaO1aDa6fGuLFX28YICNHf
VSZiYMjlw19ndw3ZvQpOTBX6vv0rNbZeDLnPa22qsE0GkvQrWi7R7CxPasJHP5gw
z8uZex+icAI1kBb/ET+pbFr8DYPYQsYUSOCNQcRqXwhy+9qTBMR6oV7t1FPLvWCQ
/prygA/U1j60LIRkSgOaxpbJif071L5ik356X8fNUO0mL+6bn5ggWXNl2vBRPzU5
TnG4Wm7cq1cQt6bEeXiP/m42vAsL8daAgX5XN9iTo8kHOQV+Nuw8wlB0L8PB0N3f
9hdMJad6eTzRrjWBGcFaZvEVwQT/85iwcHMkzRelWibF7Yiz9nBvv7BwnVhf1HWH
g0pymvaUB7Wl6W0WQg2+19jdOkTU5wvhSmqlxyt+ybIY8Jq8kWeVqpk1MHLstRL6
TOE+AXQ+kIRcjOjQ38QkWGM/JBAcnI38HG5a5vNulw9q6SpTxbbuoRThR0GQNvSd
hngWG0jmYBL0IHwDXpG0Joj1d63SMO265v9cwi0ONdW4uRH3+Lzx5xHszUps609h
AXW/zoCdCVdxIpzxEKM3wotpyuHn3axPgzjl59kxVkJzrh9dVOXAC9KmlNoCQ/bt
D90jdBPQgnJF2DeOlu7SRu6iCZgn2rNpzFCCrX7hLAOAgOnbaCH9Em+pwOZHv6tV
ZHhYg5DRRCUQnAt953X5M5UXoS3W2tEvxNgMZu1lQsaSrvuFTM7dPtba7/Nabn8L
58RKiUakSS0nPo1bzHJnBIYu5BAKbN/mDgeowfhqXf4WfmtIJmA7ipmH8E9sCoC9
nT0ts0mretCHfVeUKb5+Vu9rrD4pEXFhZeMiLEPP/eW3mMjd2n22aCPxAaXc00Rh
C6J/QCdcn86XRMj5J2Uf7F4bdogpKDVphIjs/XJcOZsalTU5QP9++pNnoXEvrkdc
pdwTryKAyJTB+AmD+eHhQHtsIRCNPwE0o2OB2ijTn6EpdB1v3MuHvYpzORip9pjG
x+AI51BTd8S0Pm2BPdE6B3kmS3evHBgznKbmYY4X1t6tPhdpr6bcCd1O7MIFDpAF
OhD+hcFG7187/mdP0oACMNlLJsDqclk/t2YFUcj3e6fKaaoyipxGz5LJ9zC8JO8P
9OKLv3Xw+jFG9XAQ4fHdt1oJFlbUpjJvcvxpnADX1VyLO+kDLWMrtIFFB670nMxz
Gxw08BT4XYNgqocyeDw4DesQUBPC1fgYPJuGumUZQcRm2HuLXJmQKduEenBhGJIw
4kkh3XU/YC0YSj7cSQVEkKPA2VZ1pDx146UasTJosBXVgbUixjWTl9ZUmrN5o5FD
pdcaXr5ZRR1B3/AhAGqBNU8TwmJX+x0zymQ/w+tP05dUMxhYs1zcx3+AU5ElpS7N
rJCEHEpjzQ+jPGo592R1oyVNN92xF2/mwMBSi3xhEvVLmzFyBVNI88y2zjyM+Hjf
aP1gA6PNpv+7t56OEjRKZoI+8k1+1XU6f+V0j0ekIh+udRANGBBdkYoZP7n9Eguk
k9EHJY02ELMbEYRilIMNXri6bf/wwYX8YKSvK3QfIE1HdwWf9uBrjaRm9GusAQE2
WHYwXNjZt1ph5SJHAwixU07l7aAQoFiclD2Us67LRwn6xiUC9LSbcUYj1QA7JYSH
5lF50rtDgw/hW8LjiqO9aG4vgF5IqiSA/eobWAXtiBpk/BUhbUzn73QQfZ2WnCEv
mUQC6yPtuTa2SGCs+C1RYuIQ83WaCXfz+79fnKej1pLH8hmJMNfkjeWUPbf4v18K
F2h5FMTyXEN8gx9DkOqBK83v9S+U6CLhy6QSFSarX6EoZIw3Qt50osmX5UkEFou/
eYffBzLiSjZjmcEcAIfrcwAkcelx7nMIYcHSzJ6fakKWSzG1uz3MIqgJylcIreP5
a0friMjrF2d8IaUcRV00Kl29GJZSZyIdQ/DugxHEDIi04Kw/NObCBpcZCA4PeX+V
+co13VKsiL0g6Hf4b0w0Ae77csE0XDu2LTHHejCNnQEdqWr+yqDAJ9E6Y+k003yE
Yc9hzSqRS16G1GjMHnHBbh7YYKvMDlal3pKsVfd3SmnU4Tak5PsiTXKIe77hMUQQ
buDw20scEfcQOE4L0OnIrL5u1zNpFlp9GLupYtfTCnvlZQb4uBp+Uix4OBeHdEdb
TNqbi42l4DhLRT7lgEwWEUBaBTh8QSt3IFva72LzQ++Ig+Q16+B1jpA99E8eLddr
8p62PG2ffMaiXAtyO7pT/t5i633G2z7LCd25uJuwF8DuVYN1i8Ilul/zE02MyyJe
paJIFzXCvzmimrpI8cNuQ3C8advunNFuJ625lM/eFNAiAmPa5fPi4B+/1v3N7TV7
df4Wl2zAJf2S04r/1+2oQcN1WM6JkbSjU7L6WiiTNKtMgDcrxQXOAfaOvumSTzdM
iKNeKqrwJrxFKdPqi+e4Xda8Rvk+wD0of13+8p9XQEaIt1S3BKI4s9S1CvAU7zYh
Npt3XkZy48uSAyRdIUSloUSrR/1VSmv3kg/psXve+bXWAGvWhrTUrBdm9rKoBRb3
n7yhpQyyN5FtmnCIoRgx0wvkwjmwyb7acg1o5mIHEeHaGMnf9Xj7jEi+IHNtEtgh
vkTKIq0PsAapVEobrAkjfrVZOzZd/IdGNRagojycvNY/oWfDniZ2Z/HkD7kD8rrg
aSlWqG7VHbjQQYOAO1CLk8DVjRWB3pzJEDqtfkkdAPSRBSMVOygCVebRJfzxa10d
kKY48Mzv0olcXK76+ijSSs5cB+s9OA7AM77fUunHmMLGXzJ4ul8dJng7PzsM/Sv+
rMirTGm23HN12EFqQF8ID14wLTSOeLvG2xIp0PoWx5Hl6vVbRU1yrdm5LYixbNKu
68+JTmYgMgE0k3ZrwD6FRkirrSY4UThqjt/OQcHz/N8tb7e0Az6YPMz8AeMWjKjw
NQSTTOrv1p0gWzg7CiJptUZUznVDrwhoxSgAwdWS2BXeFnbT9MN1izvMNt213upS
udnoylPqlDVdB4BYTsAMbBQlYjHdjiL0OuKx2Anptm5Jr+so6cf5iNxuOxc7uvIA
wdSwlrrqS7LyjCiz8dtuo66K5Zzmjw9Ouew16FCSjCFnbM1SDi2YKQn2OJnleI2B
BPmf7TZEc51iETgtyx06L3/pe6Xt75dJGr93Md9gHQFbgW9DwbcRw6oP1xqyY2+6
l6LHkDHPsPFcn1FQfyXUW93wVUqy/ceoISsE8QF0IxeVJCUdNqfctie2U0uzbVEZ
6wcmK43j7C1wU3SkSLsrzn98u0osl4JnabtYgdy6pCBVzbkcmyHAQxdpi8CVM2Wv
XFKF4NoOf+ITdTj/QlLDjFP/vZvmKJrUCeaJtvOVrSd10WG+Z6utXnxM4c0v3tI4
A6puUAIsJHv48My66Hnecz1mw8yN1l007Vjhui+SOK65kPQnO3uO9LQOy0p+dBak
4gBZpzKdqSyB/HGSIqYcmYfSMm5Zqwos450O9Ppz/qS0z3GHymXd8W6fFN6JFf3G
mJdU6ozXj3tvYlo7IMrUl5tmA6zec/kOG+ZlHTmov3sM+Z9CX8PumUaDf8RNTp7+
i4zKU7LspJmFMWyCqSmkdEegwIOciLe38tZ2KAOokcfqdNbF7PmM0+DRasazKv2f
11m7AhW3/v/P7f3+OqrcUPNzuvPz4HgV/KLNRnWLceSgo0p1gVMcaL7KA4UneLXw
2pUyNUXtIsrqjKSiM8d9BvKe7aFxMCvp+cD01eqamRyntQSi2hNfMNdIM72j3TQb
3LaIcnfsNqtsfZdgNSDkGsDFYx4ZyEEJoxBvfVJPmJrZErKWFjZnSJ2J7SwFb5DA
UpGGv/gqK+/W8ysI62vabYP2HK3/nxIV3Ce6UUO+90DN9kpQUl94oaYqI8OYzvOe
KyZCofd/0bwvpE8Ss2dNhElwtYpPCxui0qinhh+am+GwaBimybrQ9tjU/S2Zq9zp
t6C3oDyMmIu+jsGOdRbZJ9QF84ERGDHjU50vu2kZo949BS7Kox2xVixq6DZFB/T2
C/okxCvVQ+dm6Bt3e+6HttmhqrGDI0dwpN1Sm62G/V5hwQWvrytVAXYr/sOs8FtX
QcXXwcyo/ACo2UDtHqCUbIxRVXwquuTXg0PkGYPUPmiTsbHzG2H1XVOeJ18itFj6
X5cjvkx5hFHgvSb/vjquH2ibdEDqflCHtRKuyXKKtbPofCLRYSDQiHxz3bcwC/mz
bL/ks9W7ptnDxoU0XO09Y9OVi3M74WW05U2m3W6MUlCYbSQ62vDZzruqam3T3zEo
ExGDKvP7dV1WH6M/qz3AF6mNb7CpXdwWN/J/0O5MztPKkzk1wjVjJMlpJJ5EOBd/
H2cuqbxabpjMPGzAnPykYPJAEOBeI/klIGZdcWb2uYiKcg8nGyTO10fvFe4YQ7vS
mOqNPy0W2ETXCyBVdMGbx4yuf2uYUKRm59nQAX7N+qQ0nTj1P9QSGqtkhwZn2jLU
m8nCsqvH38kRlmTH/zq8jdLAPx1V5XFMZiazL6bB14Qq+w/SBow9nAJqSPs2Ii1k
BXLIAxxH7bswIukbp7jd3CBnvNGLAol+DqGJfqqiH7yQe8QIR5vUNSHGZBimaLYY
i0rK+nCVYn6yXdzaUOz68ejkOt42+VDmZrLDabhCsmeF2eDnQ/lcSxnLjoKHtygT
4ZWwZoWJlgpNt7vADYvqiZzuuSYAIqN7YTrhDItlIGe4TwmdEUg2G3rpT4cakgcJ
ko+rdPKjIPRVnGyrdsG/+4E5pAHmQB5aIKF7gyFrqGQvgiOcddOFiNWv2R39+dQW
sN9V9Ba3hexFY3uy+IVK0/vczlhq3rztWhAyvyhqCWwdmk4VBvjD40B9m9lTNpSk
qmxYLhnHLK4eWEfcGym2MgcYqDDqiGucDnK2VApWd7FYaJKUd//o0midxiPQuR0b
o9gyu682t6fLnA6gBAkhJ2Rnj9YtIkvFERM3v5qEKp/ehZ+GxkzlMt7AzWkJ251H
jnH0t6iHiKYNZn2x13mWmjsQs30Bn8WdZKfeoDB0JK4KaASd0I1Vp+JWZ+NcjSLa
dELmI2+MY8u7ghG//imL2dmMZMVRJzoDZy5jBdiZdFJd7g+91IC1ofEOVYiDJN88
CQn0NeH6qr0h+IyrRR4D0GpwV7d6N23XlX53L1Uaah9DJMY+eEsMfju4KvTxT+dR
pBKOTnuErNHdXJQwGArKTZ1wz1mmrF+gTNywJLAPAwELNLh1+Gj2fneIJhcocuna
3cXtuF8LtYr5i1tg9sxcUA2CoZG6R5WPpcXiEOdekUUGUJdjsQ/kgSmPtr/EQtdV
VuLw56752kMMx795E7PRmbrfSlGkbCdWA51OUhR+j6YW0mOSZK8vKtfjy8ohoDkG
vFbF4j4fx9DyVL+xWhHTgAHk1Yb3loiVJ6Yx8pO1udKBL5/ebCUjpAVbfOaVUjcN
7n/fG5N82kDBDN+Us85IjAGgOo72hDX/WJufg9v5XFXqLBtpQb+meZhaa2thCMeY
Mpv40RLa/jGNaElG4IpYVH8CPdaxMQ2suhC4LQ93e6JMoHaQngRl7NiSO42Tjabz
6SWJL6Zyu3048kGHInEbZbuuyxSybN+wbAn/QvEXFlDoYUDvQ1s8rC5dgnBq5fRW
Lu/rNbQ1xMBnUugL8Gc+QpzwE4huvniVTKpFzt8BkWgvL+bRJFw5ZPcO+m0oiJ5K
kcYTUpXccVa0tW+UDgYN4aGx+KR+bEw+1RbRoHaErE1W/lB7LL3bBXlU6Nc6xd6C
Z6OQx8a8Q7LF6y0YTDvWLvkXoaQu8RxKiGaus5T156yg7xlwilt45iTLDgR8aIIi
9RvtarKXuyDfh7U4DKSfUiq1yJvF6FHnI0q40J+huLU44438mNTbK7oRcpFpGZTK
19QRQ4yMTwp154r1ZsU/djHqTwnUCx8VdbcxjSRXSCX8HH6FtaMLZ5Yvw2skaCV0
5UDV7d5WNMzsqO7RSUDYEMqODTHWi0z//0oahG0qeA/7xSvr3fJjQSYjYhw01S5X
WwuxTIP0J+WcezDPmuL8uujIu6cUyzJWWYJSlqay+gUbguGMTvb8W773vIS20pov
4k9yooixQG4T21jqEBqtFUIsvNGVUVNcgx9fGerOo1N1UQQIP+Fw/Fek2HNN3Bu5
5Q2iz1Ecwj4eQQ7KCXsGi/VHrffnz+9pwwXGhmb4nh3fKGBjBmKfWo0II2mm8m5F
x6iwX4XsOy+eNmSyaz9NnWRVKQJnw0nTgWTXI93LIi/bLw7l0go2trWCqwhvvdHU
IqoRy8OWpF02pU86nWXZvUq7bIOOEQdKRFr52PNUYvqM7RjnVhtD9yBTngrIH+y2
uJZznfaxJEfCsqo01+Qk6GMQFsQx9bjQm6WxDgXeLS8mkNBKs3huc+dliW+iJstN
77uVO/BmU980MdSoF1q3hxBWYoAd0fxUL2km3z1yYforbmqX6fi6Cw0f+fp46uXd
0+Szsj6tgM3HASj3QbkdgZNJD7y5gSakramLmX+iybWK9T/qy9CbdnZ1DMzMgP2/
zrao4D/QylqVQT1dnH53jPKeKkFX0eWkFpuv38tvywIlRZOZ3bbvlnqNUtjvOL4q
kFMV4O/IMkTak3raMl9jUscfuQvAPpqdx2xLDE8Sjt+sfYCapS16vSPIEnvFSDkX
tkmtF2lVEu1WOBoemshbCNeJ/Z1ooWH/FPWDFll670WBhF5ZXJQFLZyAef9eKuod
Qi6PnppIscxjhQghGNgFnkmm3vpg5Ua5vgSCXkBz+DQZmPzb20UodbF1KeVr4aQZ
GhjGFcIL1Xn4AUacJF+3VQ1cIJfThvocaX/Mf62M3szdAuvPlG7cwrcLOFjFPgh9
02Ozqoyf6rlDLQ6S57ZQAn2oEjVGMKkvbWcnM7ZPCLN6x+zs9uWd0UROGAyttG7m
J94zc/UJkrX7DTbjR7VP763MVpjabYTy1wcX+2USJ0jAKxesDZfvn/s5BEr+N3d6
kd3Da798MigJsh4Y3oSM0wepOilwirlnU/LtLgim+8zrj1ZBxGMM0L6Av4OqzCAq
L2g/51NOZP+0bchtAzkk9Bj9I0gITCZrmfLQU/fGJUfhgT6h9RgIVkjlCkHZ9rgd
tSFdkjDkEeVP4pfTrMFU1SrRs8EBMETWlzMHCaClQBhcB++fXQNbT9PMhEibX4xC
SeYSgTfYHSHYW489m2ZUbzACFKKIQ0lis/RoZItuIqNVbOkmc2JdnHpov1VoYuPV
FPPW91OyIwLyltKccwFvCLhEoRRXd/3hx8DtWKZQ+33DYTLE5kMYGYuFtNDKqyAW
4pkpvaN4wt/pCekXA8t4xbUNIyY0XcJNh1scoET3CulcI3j0MXcPi5bSnow85OiK
eHP8498mma7yt2F4cF0leVI4n08pd31jlYvHkp7+mrE0aCBsANr6xLbZqL9KjQt5
alCSHVjmKc8WCZLe/C5gest1zcR0phRaBVbgfk4jXH12Ud47dhVu8MZ9djPzGdLE
rwc92TEt+OhHyJaX7vDOWd4p8t8xqBUlZHNam14GsoqMTDLY8PbfaxQZYr/fv6IU
LCSOcd5uou6iU9qLQE3nErpXfnTpVnRrs1l2pSyKVxPfnvSSlO15VT4pJWOwxn3q
+CYQNE5aeuavDIHbZiZqMGmgvxduMSrsvsyHI4Qiaonx74bsyHH4Ag1Dnx0ICaeO
5T19M6vXLZNxuuFVFokcKfPJwdZZMwgLZ7ABQIv7dkiiNj95sD7n3za87xHDYR0P
dXK/VqdHcN/sIIgASD4yYyPkaMEd1DPUEOOAazmAu40x4ew9fAvhDW0O+hZ6k3bp
pZcCcbQA8GG7ry7bOldVaMBjfctL5qGYWDhENOzexutS/rnSJgBoZjrUQ0b9Em3r
ZUYevDyd/jdNyVu3gwek1KlpcP6s3/BjAKf5Ax4SXdFqIknREp7HG18wSde6kdwv
jYokKsFpC1GeUqQr5zfPEMsrqLCg1/R1gnddVkjf4UNxDxBPNMEdaku1W/9jccXV
ML3U4kK8+xqcpjD3dFYudxvfJuK5885LZyF5LHp8YwiwYFuyfcvGmy9zcYKQ3tM2
Dyqi6K/uc7MqSM+4bdhH+ghumw6BFopZt2StWDFIGBiIuj/r04I3OHpwl8SKd9I6
rXzw1KWZWB7P5KC5o8hs0bU9z/OENR+QxGxTr2uSQLl8wVjUpTid6W+c2J3JD8oF
GZ7hYmpjqlpSU2HtXH8MFYMU7z2rmR3jB/LOmKkETlDKgCbs05tQKLCloeleRSDj
DBE2nikK/BO0UmBoFle3hJAyF7kHPHY0KYbmFKFzFvLHMTZ+o7dknaeHl9kFYw6X
rp7/lna9dDnH8A6upbopzqQQIpkfodG8zpbxZ4MwACKx57nMY0dqfVTZZLg2NdMl
7jWRoWuYU5mAJLVMwbvZnCUpLlg9HNBo5eSHPGfdKDSe/BgelIoyM+5EH3YsmvFM
Ai0wmFiwc7kUS/zxba3OacWHM93ZIfTATVeGx+2+TRmVX631S0DNkjiHvzYpr3g6
+PIor9n77IWyACUQZAy8vBVFM+nU8K6nZJlAj9o8EGe8prNKDa6H7iii2gQWh9Iz
XLlPDlpXRFrtkOHP9LriLbBd9snOKeW4pWKKTfaQd8ID2wQzNwc+J0F4TMsKyGOT
aCcUO4rXwZPGKWeFOZObYDCliO9cUAKUSQB4wHyNdd4PzxQfmDu1UAb/R5fNL5Z9
ueja2QfmLFUSJcGbdD1NC+EMflpHKF1Tt4jNEJf74smqnVpyF8Y1jmQYlXkxxxTE
zNxHkZjxNpmKngQjazaRk/7U2kS05mb1Hqukl5bP9y0tEf7AfYw1IM6+t/6HHArJ
G+IeSR41VliYF0Jm+s0hHDRhGOJ6i1o1nUQHtiT4S59u2+GxaPkGLS1OouAyzytK
1bJSh9kRXg/6IgQ0FUSuaFQv6UEZa2XzGdG9LorOhJ65WUoKEt9JTCdvsfK/i4Ms
h8pNGYXgTJ2DPBBX64s8Q7NLG9xFiblOXp6GYxHqgTDWik0GhL+jUQjNaQ8S6A2+
7jvsYil4OUOgGTdlPLKf/9nbg+cne+iwPdrKE775t4L+ErEWK/L6FZXe5oVHr64F
vlCaUvI2Ta5DOajkZJghagtTyE2Gashigvc+K/SdZlAqxjwgXo6wJi1fGbsQ6eow
os+X8ZC7urZFKDuDQ1m0eBBJX7ZtP+T0+7EfjnHA7btKLs5nIuwCKuoxoWPjT2aR
O8JOdWDMCt5t4IZ6HAmLKdQMw84vc7BPk6ZEwlDuSkRzxqRT976EgdOxU+UEPpRS
J4EYSZluDesSbvRHCoCGa9twB7q5EUBo7b0GkvZTiANIFAYna8SrGMlbXdmbz3rW
4uYrqK/TF3tkd9UjiTCny+jumqJXTpC9XVMVYC8Qx9pCJ7TuIne+CPOaSl/jjxW7
C6npCkBSv5R5Q4q2TNH9TAX3MzX6E1UZz6AxgQp8aJz2KvvGAAoMdEeytubmq0XJ
67N34TOS9XZ9D+WIsnArFCIBQl4cO1KWdpG6N7p+kEIvWFOwr2jIsh6VLsCZkdVJ
PhRfv16/T/+zBUmlUA1s63AFb7VCbg763C/Rbu8vA3MVCevDNz+VoA5ISNpKzqvA
TiPYjIdtrxLZo7n2moJe/bTLQlSGOK4aRi3asbN0v1Ju//NMulIDTQbsrjtdTX5j
zrYxG7Op1g0AV+pLu6CPI8z3ANv2zT1f8AtDY7eBrVe6zj6ZwN91caz7SAMDv9k9
orumVcIalLJxSvcM4Gug8ygDGVFCFNO0dBIcKVfvYuRS6icVQRztesvlEQfBZiYE
P3Lc1GbqepTYZm7B8yMVnLa6No78FnoIuPl2vgeiBQ+uNRWmbjXO/DtIbO708ce9
AoL7CuOvZMvouxP3qzpGehPN3CDrhHlPMMV5IgFJ9/oEo59syY7Sp6rg1oCxrU1b
rsrb4L35nwLKK9sSILiqGZLRLhQumEly3oSl+C6Z869Bd4H2dsJe6QzVe+Kcmer1
CV8pbpifOuW7MKjWASfQjAQQz1zt3IQk+o3AX1QKdiLnWyPrznGoTYFdzJCm/qmb
RHgda0SLWN2zWGsxhRN3qs2y7kKQ4YmbF5/kItZr9oY0MycnYqybxvzn7XhSxT39
O0Xl7Fm1wL5Ww8LA/pHs/N17T50is7Aw4VQSDTSxesBt4sBFSZ8IBgfN65jfk7Hh
ESmdSamw+zRqXstTO5E+iYkGeNw8lKYVE4Bkv6Kpkcw1emZ4kLGjs1zq9e+2I0cP
h0J1YfhyFdPvWpkwo+MG7KcvM1ZnzQGZnfPFMGUZGDbeOyGcuD9enF9ay7+ismUg
0m5wpioQDDkWTx0TUw+cFv/U02YTT9D1/duC/bves7igpOxwI4qZ8MscqHa0uOHE
ExJ76lmaow3txwAFgPiZsyzXk8Mz2CfxFU4dekhqbMQW0N35SsaUbPGxZs4rwGC+
sAbudlz0IBI6QsXRIrkDaGB92FlxMV0tYiTMRcnVJKJ7GjBzbMrLHGW76L1AEMmc
1DCLYF3EuSz+LznNj5JhUBDkuJZ/8VTZ3iTG2njrgP1Ctu07XtitYmHLsQbrdeHF
PpssCz+ZQP8jqTtjMtZjwp6a0vc2teRxeFYgwS8Sbz99lzYqXIebKSLrqVOT3DEt
VlzjaSirRSNAdSHBEzmWBKJJyWW9gbxrHqOlNGlVrdSW5TtxaWqasVIB2ko3gla1
NBGNU2aGA/RvEUBiyilRZxhqLsdcQK+XrcwKCpuZ03AKj1ongdDkzMkoRDVGYWfD
nK2rEzhaoJVdZsw5tBvEc5VZIXQj2kiqdZ/BVHiGFrutQv5WWcrDqMM3Uab7dHg0
jmtmsSls/JwbcoEZdS17sBeqGK5s7VPMUTFMTKlV/m1jt+1iWh3p/CFCq2z6OgOG
mxacS+z9K+zZdGlwO1zELeEx1fK5UNMaSGkILt25lxyOz6jZzFISjrkWpcHs/Sc+
sUUaib2b/vzYoVY0opqo09UHss53sCsDgtEJ3c51PeRBVhGRzgGqOYBb9QtE4HVY
78V8QAxec2IBwST1jQb1JWFSB+kww7OI3YRj57IccFQeci+VrhhCnC7NNC2gF7fq
LgvvR2EJhvt5sbsp8XbpKumjhEPF+cHLqsqJoeeJsQFt5P2XoTTLOxLMi10RAEbk
iP/lXdR+xbRjS2ipC6JCsh02/Whi6mMBe0qPidY4XrsPyK8sThdsx4j07LnVp84w
8pqNg8Bx/durasgLAZIYkRqITfZYVa+iF382aRcHPRtxD0fE1a3t070iRs2dbcyN
dVUfUPSdWNIeXF7WQbd3/5qgBiUOdkVgey+EPG+Otwm1sOZjZfg0mPA/nfzrmTh6
60sfcLi5qF7MGF0+x8VyOaYNoX+584lLS0FijqmNNaPTWQcxKgIU+tw2SCTbnrkP
tE+ydUzozpqxLIdD+uZrHLzXNZVWVNFyOjindjUSyjFJmDi/5JTuQL6vDkJ+8G6i
HJOMAXZhkBDSEdRNNL5H81/Y4FB6vpV1RKgbw+AuwFyidEgXwPue9pe4SaB4pUkD
1nRi0XHSmQ8Gf9RWuUrF45ybKsdb7U5vai/n22vjeF9PYZjpZ0QDDhQB7N1rVObC
4QQGeoqO4DY3aGyttnAa0sp+S93IVSKkA81ftQw317/Lt5YQS4CoMtDUYnQxZv//
UTtoLg+s/PJpHCzzDOXLwy65caz4slerH47HI8ALE0lYiU7sB3QR1GQM6lHhpyQ8
fG1jH+TiWe50/HPC8RkZU0vB0F7rVXpUQcCqY9ro5bHcDnn3TehGnoABHWxSdgjK
ryEIvl2g1SB9DeQkvcSTmmBJD/x9RVmiedmJyCPCvC36QQa5MD3j1m/FI9Y8acec
NGhg3kEsED70+Is85v53+Nn81FikuJKgUUuLvESwVR5/KzUmPdn2KVY5Qm7LHde5
n0Jf1tXFA5OwOSio5KjPIkRiA5hEm1DrxwfT/1oftJHvw6p6rpSQkZlhIej5sQEw
zEAAfkxZytXsuhQWMfRLl5m+HAMgWLdM6PkJiQAAaeoFqIuIVEAiYIKdWrAugLeM
XKm/wjRJ9IUNdAP3sGKmdecOl3YJqFizCT2lP6HaWnebIH6AAfQjMqy+UIJjuXwc
xZ3pSOsy5xbqS+YwWGuUSVhxDV4x7PxTGa0EkhQxfxfz36sJUmzkmnJIhndsFrP6
M4tLHSm6Er6ujqKejuXan3KUVoHOkToRq0drxt52LJ/SYSHMMTUjLl7Mp5zSLxea
FlPyBeD756e6K9ZwrqaO3CRu4Z8K7dDKUJgTD9IKhV8CXYvSZV32PA8/RNLZgFML
UO7cFB4ee/l2YPF9Jaye8r3HvBwc9Jj1WUUA0rA1U6iuMYtsf/2C97gmaNYit/Ex
NYW8Q38SfDiJ5JaFzwnpMoq8ZWy/5Mu43PAnJT2n0+5wmVF2ATGcLWDnnY4+MM8D
ZSTpP27Jt8ckGomqQfl2dCoH/g1ml4eeqFVFzLtpKzpSxyakTNFBDIgzs3P734VA
1SWI6b5kJfdfZkLNh3o3i1d5nj1MtQPzThyxjA4T/hl7/ptzB0a1EcxuKaMwRYit
NxT2TqitL/Wcg+vV4wKBbss/osWjrel93VOHUuJsh5j6uPQBhkgAXHSLILZBNjkB
6yhrtNRPb6ZNf67XNSruWnEqvHhMt9dkQ2Kwzm2IE5hRshuabZbqZFlVOTnrEw2b
sZ0nlmfrGDH/apgbAj1cvlsJrvcBmx0k+iy7IQ9nYuVcVxKktYYr3epZ1dCEkbV2
oo7NEVDqhu6R4sZmvmWb+9NEcnEONXKajuusgJJt+H5tG01a7QSw1S+tvbb1JEvz
L9UmL2Ri8DjwzY00eiaOzbMzup8XdPYLBakyfbZ8vjrKkBXiWblh0Txk7m6KsTbE
J9nCaEtybMygiwRG76pkwvzAe1EzZApTwCNddo7mNwzy4XiaS/Sjd2WbYAtsHHB7
bckdDWsfskl2qXbhWoomf5uNJVgkGIQ3/XncCxZmNxjY13ic+3ezdVCa89BUVfUc
D8i41lA8/X6sgEeuR94pSPBSRwGwRrVKdxUXDeFPSv04cMluXywhOb/jpMkqOvg3
PfYIB0R4h9v62+M36H5hjrvtFvDZTGiuplBb3Hbnf2HgUyeSc7XvSiJOmf1ztK/k
jmObhmd9BRtSp2hNGwclgna6vGqvZ6rIvj1Jz98sv5NKs1PQGuZLqpiAavkCF9Zk
GeUe7R0N8UCz3tfM2zxNsjRbXU4qzvKihKlomTNHVAnLLxPV2DgwXoTFa5nnvBLC
2EqQPACjADeLJtNXZqOc9TKOO2QiiIYUw3U+ZalHZsYPWj87mo2D8KFZ3m11X4R6
U/N7Bl1QW9qiAnDZgmiHDIWpZa4H4mS3iz9kZGmm8al2DlCA+4+c5yAPtuWkDIBn
Mv6a3Bwm02jK/eTa2VtthCN2LNq5RlHQULzq9pffqA+iqEQ86bbLIifPBQ8uuB5x
sr5d9L7ejGfO9BHVM3PQffBpOy4cvfgL38ZAnpvaWOA0hdOdubKKstvp76rO+f82
g7lhSNwBn+RYnoqRIzjOqbJO4HtSJdeQbwaK7l4Ecg0/ciA6b4Sy9U8b1Y1u/pqm
D8JiZzixtBCe+aomvj+DdZLL7q9mz/f+Jii1F4pCW1nhKLnWRF7boGR8YRXCKKGB
6mYfYceeQGk1//bSvPapF9uliZ75QWtKCMeLL+F74VTpPJE+VE68gjHvDSvZAiiq
7KUmoYbUZrmWk2E2yuTtqM82KMG6UaFUdx8Na8vD57nqG9gowm6aOxnrn/h8L+D0
24Bz2bawNJ6QbtuBuZfTKHwKdbEH0ADeyyk2aJt9obF02mZCwISqqBvC7llIttV0
VcZ9I3hYuQ5JfR2dugKQK76nLpJ5XKzjpHukAvRUBaD/rYoNaR2IVpwzuzDqysNz
0Xcq5aJoUuLWOa18pF48lSXcnNWxdG3S3DAQHX8WZx3WiZoMRbelTDeBq72jaZ4I
x/C2KakokRzv9le77BUuA3aH4XpJ+ujkzKM4h+sBJZuFFNTZb/Zjro5lVJvR4X74
WTFSjhC4F2qxgIuMHcbWYYTHoGnwuvJCI8QXvIbz8hhd88v8PqVg0T7UMDLhoyf4
i05YS6x9GmesciSmg4HSVDu735B30WRKz04qso0+zFsbvajg7ueyy48exY8+qS1N
eTsq5qmtedtElyYFrmxRPyv4BGpwhJeF5Fga6GuXJvaSYM27VTgUgJPKdA0n+6QB
e6NX+q28np97ANvr3uJhHi2lu2HOc52mkGYHarjUq8k7q7hSmqdd04eNHCu4knqZ
7s/0D2tiFTPvBtLedWVp7ZizWaMcG8yqkATxbx2twiw/MmTfuCx1k4G7xNZgYD/+
NBMpEhDYCvpAc14VvkUchi58NV0TcWa1/GGp7WBttnd4k+769iafSZPyxzNlTF5R
OH+4bXYlFe1DYstBWy98jRC1QNDgCQmH6ogIzq+akmTeRWMwrH8SL2XEYquBeQUJ
TbS2/2mMzp+IcpXFRIZztksdHo3xZ93F3beR71g3SU8jzL1kSHJ5pIVBqUQA+xJH
hPDuFxvW12Lk/uDw61i/HuPtqLr4HNIcoJyWiBD8Wrx76N42Nl/qjl5jsi2WRuh2
2QUjyBKefLwi9CpNobJ4zTokosGgeGBzNmATUJS3SZ/En1NSEk/Lx/8fqzWHDF0a
fvWYzmSmCpDKtyU9pBD6n0y7znkjmIdPAPmpMsc8O549Kj+CHv3F/pP6oMHjjBJc
DHp81fx/cRT8r6liW9nh7xrJTs0zl49+1i339jmmxmcCFFR6N15Qx3fRtEkp8ujU
SiElKRRZ40p+HoUh8qZOob9o2vDm8Ck6YndhepMwdrqfLWHB9asAFOwIAVwmfLjW
ozctYUJsknWTEPFxtGxGDv1NpEJUmc3TsMjbchU6tXEVGLlFNXYWxji4BzZUb8e1
HFN6fdIn8IWeMAmb1v/5QUZJF0t71zV7Z6wpg0nLEiBaoN4dZToNIwp7j6wADLdB
o/8DZZnb/eQ+hhcFO15zKvCz9dlt5H9qLiOBVpQlNLtAIYqIEcfZn/PyA9k+PR2Q
xt4PsljaPcEiiNw7e5T8IxS0DWKIMijzUD3wojfQRBpzE2+M2sBCLVAxvMD1sI/q
JvkpZRYMTmwhtTMhG1Mio7nAisw0gvn/JTzk5LJHRAiVuz1wj4LRnONo2nCaHZp5
zTUbNwiy4umlf6JGNUYL56pZYHKQq19BDk0NEFobyAoL+YFXoPUTjXnLQ7L0FgQc
x2xc7CVD07cWbelLU50lzp5Fs7KfhJiYDua01zyXLaVmYNxvgA6adyrx7PlC8l+M
f9hGxYEXVEF59GlOrZIgA7Qdj8XKuY9OPITHTDdg750dpq8uLkVYR7JEbPGo2IOq
g4TREqFBBru+ymNE6vAVx9ZIRisMIc+pPOcPmcVLBozuptCjlju0ixTAtguffU8T
QUSVEIWdh46S9XVRSnRDgY3J0Lt34Hm4qC8dI+KVXNxJYYGKj9ndVM5+kMnzVNUk
/PhkFg0CpZ19CUTsiQIhaqbdzgGuO/AINVezuJq69mhqVThFtEcmLojXBNahN9sV
5bvxF1yRWDa8J1KJpFIiTaYzJ+84SHo0XK0T58kkjlbD9JdXd6RHyuQSuOkjnGqt
kEHqS6FOKKGpy1/0CrelOmeNgqZ9ubnEmGvkPBSQTEmWHkhKpMNXAan7Gfabb3eW
UZT5vZbjuhwYeS99D3To22Xsr/o2l8MwScHnVx8Pu76mahaK0DQqiL2QbDCU0DNZ
4NeevwxKjIbKqdWRZqjfhHT/PFne5xesJsUOJ3hq0KfIjhYz1GihOAfZRCVnabBG
YtEg7Crhk6lNqd4vHxU2JK2//VGcZMO83Wpg0l1jzWGVyl8n8ocZe0LmylQZr51h
x/cjbVCjCbt7RCsOWMURTCYlCrAoI7Shwk0Idz+CjNf5OdX/rnJmPz6aGXqe0z/Y
yZ/CKpFLtBbx6OqYDsXlMgw7mtaimxFUqM/X5JDMxrhuOPFUUbcqvHGtRUJA/6dn
47WL67xSpG6eH6AsOoty2GSbzu7e5xZYTCRGBo1EzyKEZtwZE8glpw78FVBcqHAG
AeRq8de3JCa2cRnc4EnV+EMyhfIdGL4IqBKSrNcE9JYDQ6wJoA0iAYgKMeJjoVMo
wJpWbs5Z98iq79IbueHOGVh2kyHHiXrwnOf4zBT5R4PWxWYFr7c5oi+jFbg+yqXc
DJ7Hfg/kgBx1orVar0cWe8mCnAe+xvpHf/SFebS11v1aPADbFEfV7CYfa93WjxxX
RgaD9z2h+jqPPGeEK277bNEP4plD6DFuoHMB5lUBfUqbj60GW5JoaLVi0DHSFWrp
J/Ed7i+38coS9IhdHKa2ywBqgtgBsJx0Xna4YR88KDCFx8a85h+IwXxHveEjTKau
fW4HL7ZGRz4iiRJgXtAVWL+50SIcEJ9TYurFziIsZ2vqvGSh1OvFOhSy4qBhTG59
AY7hZsU+cK9O1dst1eozH3rwVuFD4yZy0OMssSFN7zUyQ83qZtufLkmr9NE2KMnu
7wbaYK0NUU45FLUFPy18fyPM7Z74WuMbIRXoOQPhk/K4m9xlJWK5gvpouSwtKlYP
/Gx5v5VPhGPigp9a3k3/445NrqF7wdx2APvhLjNhkELpDExfGDtLzmtVX9Zyf3gi
98vlFcAN5U3KWFRbMhn7a845y7btK05kkDEL8JMm+IWFgEmk9zSbGJl9RD3ropYq
ZwvSIi43MTNU4uI4V+HHFdazdyuEb7xYWWt1BBmhD8bleork4/6b1kGxGXuocnwf
KnrEuGzo48osEbAiuIj//kdwSfndEIhWTTTLnkZAbFf5h4EstAZwkvFu1rCxlLyI
wJXxFsCHZZci27UJJwOeubceMwE+S8lN6IL1T0aIqKyQAvoGyf5/sYAbJ6UcCRwk
uVVhyUSW6lqUf07lIMH+9d+hXpCMqMGsrn/o/Cibfull2l5iYPo19uzQUhDGYG+5
quWbgpiqVRh59RdY1xvhwBhLZJ8ybBcEIUPMTliySH6NpGxTab6glMcjKGRGxiXd
C0KkytnmiTBH8s58Om33qxsO+PX4xeMq1Y7kwqYhjc2lsooiyu60v+uLK9/l3cuy
W34WQ+xK5O0vAiY5F3II76gDe2faVWqWfYnCQWBe7UuyA7weiCuOe+Fr7yT+IntH
9z/nOdMv+z4SUOZzqfEnUhgua0aRpp5BJHj/ZmMbHIO+vR7PDfl/ySM6RiwB6B+g
+/D1rH9rKn8h6L1HkxyihCaVi6ZztKjguEZ6zWevUybrf3Lf5L+hzFQTa6+zHm12
14Rsysk3SFxLZaBofR/3KguWYhmDfGQ8kqtzakNimlvKPcpisNjeQyz6jrYcYlPJ
pxFRUusSlz3NdGThIxFj1H6WC+DRjyz4Y/5y8zw5hlsXeDBrraLxgIKUEifutJda
dbkiL/HG3tBPAJQA3bu4u5f3pWYEq7UEPRuZpjCsArw5vk9XXAhxLngSRKIX6052
EwTQBwJFJXlhV+d1zGXd/MbPLtlE8V2eGdduNjaHIy1AWCnFuODoOjteZIOWgh+0
PlkVsC6quukbg+9mQ5kZ9ptzBvtVzr5AjHNDosaK2FaD0MB5e0KIZg7c3c9TNsFu
zOKZHqxpXybDZwi35FPF0DEhjpNNf1I+fbEpAOA97AY28+6IHoYupJcXjnZ8drhM
1rX6/7IkiR9r6sQCptmf6qk6o+wGTd4bTPGikGJ4i3OB0cmA9Vka7sqH/TlYZF2b
i0BezrksVAl/9PDxPx/DSq+6jl8iLiuP6t1F7vWQk66QcSPcmv1e0sBg+euvOFOf
4MfVarzyOswVuu+7f/avqYskUmYnbJ3aIAEjlWUAQnbvB/DT53UacNjjKeo2g2w3
Ti8otig21pOnXIybjoIO7oPaeyNQWypZ0wMefiA4OVx2EXte+4mccXosbh+ipfe3
gzTCEKa9uZXkbJ/IoAG5JPktI5R2Ez/pHuvoZ7XOFY17UQykNsYNoTU73pIGadUp
ec99uDXt5Bh6LmPZb8eRfz1DdJ5U0pWobpPB3m9MOX/ObSLsGIUNPG1PG36FYVwN
IOX7JZRIP8TLMfW7znivJhc1RaBPzHpJA/SENrDWbIkyWKphU+15MwAULrpn0BHm
brKHLO7lwl26P0vXZjW4K7RyxnQU8ecvE8lWYtRrxymBhEicQAsV4K5yXweHeQ0r
ekljoIU3CFUJX3kYgRHqri4Vm+oXyWUFcoNqI5Js4/QFDIXJ0kHTRyPHpxP6KQ6A
c/h60b1uzZFs7pLJ63ZKlKwUw9m96sh8jeGiZ+nKQtBZ7wKvpim7nJBxnQgpvFwJ
i+o3iaAU5ztXfenLLJ2Z6OJJnzoiZvye6zuPPJCGA+TLSHDmuqKZryV56UoWS9Qx
R6Ktb0R+d7ytYOCWoajYBn08/KgAMkaUc3i4dhDzWiGsvhnE8LmbQb5DPtGqdDGS
x5tkn72k8C6CjE3NnR+FRW7omuUXFlnYMB2ZdovyJSAdttuP/HcGy28s4j9i5P73
+NE9PI60NM+uipOEE/El7UsXjjn2H0TBXVH9+YMwjAFWNiPeELfUN/y/35bKSDsl
rQH9ukomx+xn7Sue4u6lj1tEAw69ZOADckg2ZB2+1elRtuvUz9iE5y7CcXsGSuqt
pzR23s1fz64N2ZrkGjd9nJBXSoB3LjMe4oViUnlSsI3LaR1Kq9xVY8K3gXYnHNC2
L26yjXk0L8pNZRZem4T5mP4PhKquN4nhCrDD9ZQVwBFk6WGH9kNbrLkqYIt4bTeN
4KIzegcJcRSZdtgmerdXytfuu3LCXiUC2U61gYooo0jrakdtT3x7kNdNttut/LG0
MujZneaVNXi77SaYE2SRU+FABj95z4TgOpcU8mhslBMF2f0qllek+kO9wSv2ATWg
jQcFGXpl9hzlk1kVCkqSL6Ef3ws63tiLTyTMlQlNtT6o2Us2Hw6tkhmX0UFOk/uF
O7mQEd5v6Mwh6gr9qjKG9+1fbGbj9f+dzLNgULDYe5DoNMBiSCbrHr/yBrg3edaa
C9udBdVhJqfbwWnVrvoHEL6wlVaMGIyR4VurJt7Yorxwbzcyrqj0IwU8K7nADf6A
1VbePZ7QbOc0XacyLB9Sa6SK/Ze+ISK2SO9q4w4GqwAxRN0+LRW/WXGejgK9nmZr
m/xoUtS/RAewQxbLz6/SQcsBeZ1PffpUZVrcAv50Nm9GWPzBdobru4Dqnl+HLTqZ
RCME2kdEPbKFS6Wm+n5M8w+NWn2P/Kk7+7SMnGg2mczM4lsAPz2bLVkFadRYEZ/n
8aOQAb2f15eq9LdFTymjR72uy4bKpRVUWA2hqYNcwn6cFQOh2BM55EiPjeW+RtVI
aGW/CKzAHQQkE7BxWLmDLRoB+nwo4lSKDeqL+raLYqMHJGJjGmmEzz5FJ+J27D1i
WmeKgCJMwEUp4ZsqrA4PK2RruQxHqRbi+3rZg7ZdbH56LIbfenV0Bblp1qne14Qt
HM3ZOWEuMK5TU95tFdAsKGdY2mtYqFCj1iupx002HQ2kWUz1qqE2N8SZF29yBxF9
349ghpQKfsmCK2krsOmOXdF9xefRAmS3x6Ud1KQsq8IEyhcM85yRDmYQwNXknZSu
Ayw7cz08R5zdrpwEcQ+Wu8bkIUQzKCzH2ypeEDc2LRtp7kIAVGZz89nfHJYhdphi
ITKr7tdB+SMIP6/tO6E7slGuZ9aONfbQdONG/9aBtClRfvj94yB87RwWXKH7CsfK
qd/x6gEdwqa3iBlI3G1sHRSZCkeY0BWe8aPyDWoWKejEdEt4FsgkFHIup2ZDTCNU
M7vrPgTwHshZB1Op3WiBVOqWkykIBgPoejw28UV55bxc3wN0gJq0UYCIf7C0ld9z
LIU+52ehibTRVeyOPlskaBfvfDE/AZ1Gw8udDfWZ4qgplEukrP7OQ9IGKglV9G6s
S27FVhd8GsBRMIuvZTrk3dbGC9AqDlnbVfWrNH6KFcVoY+K6TSH1dkraVtMxS78W
POHCqwPRBxex9C2/4RG3ZGDv5TTwNYJv1B3Z/zLVLnaMPiUztaiEbImpeZPCaOOF
2V4SgsqsOhBJiRIFzSR0S/k/EbxvThzd2TDBmSgB31YKCzUABrTWCa8bFJsJlPWc
rk4WbayXAHlVOZF2tqRy9jEefoV1otR6JZsnLEH7uK02oyjzmfIuICk8EgHclZZQ
BYy8a71C6luZVtrS6QhFWnO28NEmT9SxcmeqlJ6W1b3xB6HTr9tHH/TO4fBfSsl6
niHT8rrCAUApD+/91LHHRaCOwsCPTz+TwCGPZqw/mgIUgjWhShfYk8sJigHmxGMJ
S5cIhHsts6Hr9x1E6KOlTDETWGHXNAPd0vuC/0xffW7m85RsRylO6TMct6SSipfJ
Q0d2abGyJqtjGG+OEdmUrLDv7oEhZ4EsfvYWzzxM9LNHlZDvoFqW1chkC1Uk6V1o
LOzQ5XVTxFPUEmi6O3Vg/6e+ZBrihWVHTEEnlyWnnAQOIKJDr9HQghm6eJsKQQtt
d1XQafSHuB79YVTM8VdSsJWjNl3aCAgHwLHsXbcPgDTlkLvFKiqkL+jUPInjJmE3
SSLnKfWHRBLjWauv5CveDIGJvanFfryPbRTJtuWkxC/q2exuEn/kPIbfxZyvWGss
Gf5OEsV3qfJ31bw42epzHO+fPXoVdS9eg88cSlvznOQKv91aZZ/v/4A8ZAJssBLM
AOJnSUEoKUsfRzdHw8ZxKrS9/34kjM1y5lEziqCpuhpS6TpWgtuReOlKMlO/7c2X
DQsm5LiSFrwI+7d+USzqx5aJLxZ8Tn+JttENR7yTEwnPivDS/H+GgQ2zhGYOd+Hk
zhNJ351NPoQHiCS5FRfKoN6ES9UPM080MLWLzX26QonsJFNyouZzg52cRGLyKojx
+qHKtV/+r6EP/1bun3J6ifBqxPxDArJpIyAvEzkZAvn9hp6dSZTJKni3KyNNKo6a
kXgQceAiVWxwuWTkDg815l6ysV0kgj8o4k/3GjhkkciV8AHdkfLQfi9u1HK8orrX
iKaWZgr60aL5vutC2ZQK8v8bHhfIhNA+A3H59wHBu8qZlHVwGcnbRiTBVE/H4Eld
22K8oY3IK4N8tOgQSIJOL9Q8GREBzqXK9II9eCfu49L0P+2jgs/nBzGcp/ujZtSx
UevqEBPvSNz+YIeZgdrZ599LN86ziJwNgBzAwI36VDGIRnUaOS+QBX2mopyK+OS4
27Uzp34Pr4RsVMd727cptZANyWy2YhqGsiUdr9rcK8BG61H0yXTQeFvyrrJYTOeh
xQQ77msPE/WpMEnkVfxsaKQuWXmGVkdZt1nHYHztcIZqoPK+ZW8L9HkW07xM7YTH
+FPKsb0ImHInwbfCm0GRX60s+FLqHgl9yRAbF8wUm01YGTA83lgwUCq+b3ryhSXy
7YsC2E9rR7RpT8zDL2KaftbpkCm1ok0DSDF/weonDYAFshEvUzhTUdLFVQlk1J08
5rfkUHMjzHH8V+Ynlz6TR498sTtrHXByvyVLk1My4HRryW4Wbj5FyVPJs9YJ52qQ
NfKUFzSmAF3ROjS/wYe3/UKcZ6LCgrsAUXaq2tJEwoVUC5BD5gSYfyGVRzK8Y0G6
ROVKp4VvSDiQM8MgrCfLW42cPIYg7kndT7M0g/wwYzQlS5DhV/aFA4dpYoGwC9no
nVg37t6B/s6KG3cTZ42Djv6DOul3HMza5VQ9M5MUxuPauJprfY1xi1whD0X2ykr4
JDo2GxRbX1ULpOnKgdXHOltzY3o96CXjxbu1ZMef8m+ipEGFh5WlfCjQSZs8GCmv
r2dmhwPtU8U7IcaXFU9M0F0gDk6Maje6MzcDNkdCZrUcdn+FSFL8MZWaZp5JODo5
E2lYsMgnJnPRG94gHQNQ+ng8GJyuEVtxUEXwk+pbsg/mzRpRKr6rrHDEspF8+ASl
t/fy7JpjPKTM+1duTG2ELgqXLYnsGuSyvX0KKmNukGx8S2cKoPPLWeJjBncf2CEe
ZsyvujfOP28/RdtPeKORebruhv7ByoJqglAi+6T15L4j3P39MXnO8UX9LY0sseNf
fQcNMpqvWTipytjiQh0HaCSz50Rhk2s0NT7r/bJV9hgNFwT1nM8uPnPc+fBagEMl
isTRv3zHMj+/hz5QaxNQo4SVaKRszZB/KCSeliR8aHgzOc3dvn8bXWAOTDiRbKka
DKXw4VZDRWMUjDimyl90o/1BJgRgywwgHycjmaaoIpR9w2ZJdpDu/rirHwYJb+Rr
02KLIJS1qf9evhV5gMU8kMT42BAcUpq7bpTuBi1kKgfUTbeBMbhj3jK3per8IyDr
EU0UzliZAqFTUCIdnmbzljfmRPHvrtFvyP6OPbsonNEww/z4+ryEYOCqAp7r7No8
NJk/1CKhWXi5PCqcYUpQMt+YJdUoWg3LDVve3Aw2NRZx1EnxhihMn6aUph9cqUeQ
EmsxhMCMVWo1KAdyJSaqB5UYDfo+NTuU2YuF2xRo1PogHVR4a0W8Ihav2/ZCbbG8
PHYoh7u7npYCGOzEMK78A3NLIob5OjTg/jpcwBB5inj2ByU3ySq5es4P2KdWgcQ8
5TqO/JIu/oct8jcClhvwFka5i/SPR13e8E8jucAt3XoVACnS6QFv6qIigfu4NW1O
Tx5a8krXbUCGt7b4mVnuuYiA4JTd7C+d5rX6T7C3bl47fqIh+4jklJV/ZSD1KbQ1
oEh8DnrOiubSa2/vZazHuA9Xa+9LePnSSIkS4qCVhi7AYFdgkpC4gcXlnwgnuO7t
xGF9m9dKSHe+nI3gDH+QE14etZRJGa6HxWJ7eseKFXmax70hbgcN9TGzw5OQHBDP
4haC4dLJngksUAZcQ5K7RyjBXubH7FdEocbu/fXXCYonGr/gQtSCXwuJOfOzC7Xm
GMGtaDrgcqzKzIqEfy9jjVLcN4C1uyv0sbYHmZ0a3gTtEbpNNfGzjeKldfDfktqu
HN0xFb1zHlEjAW0/TRCbWI9rmiSMQiHpQd57Kj/mFHKV50MkiWEive/Z+Rcx6eCr
HxQcQKjNuotclrKUbtx5BdatE6alE2MQ/W0fI/oxIzskNLRyKAMT39Zr8k6Ydil+
VuUiGkDoNeUgup2AtjXS6eInR5/7eQIK9fR3HPc35a9H5+El1evC4ZXJcqqHF2kD
Os74Yhg2zQ4RgnALZ8xkJKNlfrpmWkhasaW/DBK0zZeQJGk7mirm+B/XDoI0T/ka
B2tgeqUgXEUuGoJdalVW5Dyy9UdyrixaM6gLQqsWc+BBd9daTNTDILseWDGKUY7W
Juqfh/zvPn8zCisXzwPqsqrKGbFDhYd9V495S0D/NA7qtZXWvYNpkiTeo5zZPl/G
HhyZZ5MDIAGbBMXsExkgD3OrHK81PhTEUfnyyHexqj57+299rsiDDaOcmsLGYSoA
QXQak+a/zlMpGhn9IZr3Et5GTg01z+HyHJgmXdPh9F3vuGOWpK1XEJFh4CVxkkju
R2ppWLz2mDscbCdao7IlL1Urx6qtthX6RBdCERzPdE3PXBUkzl75Ie52Jm62OAYu
1prA4zljF2/cT4ONCmbMVpAA5YnjZYZNv0TKLm6iSqmM8MdKs21wlCwlZ3Zs9EYb
IBnUIQX+xzO1iZ9hFpAHZ8Qw5nTyuqhjdmJGuSlNxRJ1xynOmQNJuWctIqFast8P
uLNMZ61WLIQOTsoahUevx9hvSleZlWuiKH1q7dKdqrHWukRY+qUVGdLb+0+e2OGI
MIrLfPH/eSUiLp32NkZ+oEU3S1R1RxLBNE3lrBQ3r53GZsaycaaT/1a+85BNQTXx
uaHffjNxL6Am+2SgtMssuud94SYcTYNNPD6Bxgrcha/emSHyrGWgqoxLsmOs+i6g
QltxgDTRAnJTjwxwIHXXwhAekXtRJJGtiNSrGNNz2X12v3yu+o0AG2zhAX4L3Tma
aXJTtuyf4UaSRBuRDRT4gozfnSMiXts2kRGriE5TkKmaHzZbTyw7xoGD5ldVxt83
9IDvfoibpGhrjc0mGb2DaywkNnbGFqYlqR0wS/S1GAdLJUrhwudj5g9KtS+n4mt2
K+kMHuIgTV57unw9JEAGn7nYta/8YW+TfMbj+50+9LV5OqvPiTfTiDFkrJ2Kteu5
8tcp+qEau+RdY+0Bo04LEOIWng9j0jXH7otmLSrS/whRkhrty1Hc77yU+KuulbrM
lfCjHfJ6iV8R/Kyl3n1V/rUeAqPVZ0QGbyFlcTuATJ9NwwHcvOdR7yaiqCaiUuzL
AtxmJfEai0DlH6la2Aa+PSLBKA7MLvWS7gqGxjWdHw8Tx4OP53IJ8L61gdsZr35j
iDF04P0s03kErGXrdK6mVdtCyR2o8L/qtUf+kVFaADxX8YkETlDNS7+eL+zZgRSc
Fj3E/oJDV0Y5YGqnwkOKsjDD6pUETa1GRZv2PJiibKhbrp3agIsYQaOhs+z/LMgI
x8qRGl1Z/O9Kla5qumf4StbkKM/gMxhjA4QI9RCEe2uPgz+iA5gvxxrSuit+U0Go
Q5Q4NNoqI/sGPSxH92iKChfhEd0ecqKzCpCP1/hdH8R42l27adkcjBTKfijkC5Hp
FqmUuLIlAAOh2xWR6lZG0MgsSfnzsFSmj0uEJEvgdGj3IEMUUgdWorcSCddu4XhF
fH8L/z8As0KuW+4lFOxFUrn+J7q5dfJ0Qcn0FpCffr7rS2+QkzDXl9ke/i+oz/QQ
4+MQpJRmfWbbXVeqvt1+NFlYPvo8DeZ+L4PZDwnbb93XHm8mGuD0bGctWNSZW7q7
rjwcQmCWWgXoBJCG5WHH1tP1I2tgoFLNcFTOXbOrQCXVlhitbiEZv4nrxGEsjYVm
hzGawz1WVO8gW39bUXdSMlmza/QYRHNplXFTxg6iCRTjyYrAQd5KC0xMyDfhrBGR
R8ZlRFeR28M/Z+ZWdFELPUc4RBouSobc7SE1b4OSDvv81lQYp81GK/WIh+EhB5Gt
oSnBhoY/mS2qOU7FiTOx2prTx7PD2HsIXJKjFqzQaR2S7udjnU1Bu1CRjhtl5yM6
+cudGcc4ri2C+jszA5CksUmmjqXUjdY57LnXdbRYa9KUpdy5Nw+NKVa0/9YJjCZo
5qpjpKNaWcXILGVL28qTbNaI8Abs+7akyWox5VddueLS1cgU4w/XbEVEF1CyOwIF
AOHyj7XFOOEUe3m80Ge//uLZMlBEkz5jAvyzj04BigVZjoJOOeRdJ9S6anu8Ua40
xTKmvOUTY5efJh2DJHN4NUUjvq+5zFBy60HCxO9u1SKAW7jZkqVS8h3nZuch9tZV
vF4xmptyy8YklZYPXC0DT7ZSwC3UfUlBbU556VBAnRZ0/OW02I+EuR75PPHdJL3g
yfxW2z964qQtzGFt/OXhhpmPrwlb20iMldiSFsfYhnMvRUMHUj1JZ4Vtd7X9aTA2
hX1V9wwJaD90olK/IbZinoVjE17T+EgROgSWxgb7Q+jeiVkewCdQ7tXzRSbzEz5w
GMIfvVggvZ2Y6Fc7ohNxO1Wgcy+/WfWo/4hgnePsxlZdsRXyPyqGfEi1iJhOvLVl
ZxbuKd7F5FtZvWCPkqymaZNk2gqXCqTLMSx1lhyEPUlglapk7fRFvAxwE0xHQBoV
gZo8awTJ4jXq3w7c6fjS70LIWbf6ximoTfi9FX4kGe27kP/86OtIgG4cdd+t4QaC
Mn0VGJR0NTtrHhj9RLD6bcGzvfVJIKRR+rB43NK6Gg5PwO8366nh+adllf7CcM9k
Gs4h99WCiOlf6kPG+dXZRnspcvxJnkZ6XihsS8YEDSDT5Griwp30NAnpl0FVGe93
vsW4eCGnHMVgeZ0r5KTQeNoxci5bHxk7TAXlcLSjge8CYS9sAFKnAGjDhZZWswow
m5rVqbF2gVdm3be8o2Ic4gOoWuhxjX2NJNJv334kxJekYW7eu5ky6VQS0QetjOiH
kFdb567paTkRPFEPzx9J6XrlOU04sNCI52hve5AAf3FEMGW2mvi0BGbSfo0kcbVB
gexea9oX06Jy/52y8kOZ9gptAQBlpibI2wv9mT8DrwMvrqjp/7eGp5w9lo9sU3EJ
tIIX5xfUWFxtx8o5myLlODPWsGravPbzRYK6xIVkvsvFNMzozhHQRU4TCOYg1/OW
Wq7/1D1MWdFBEJxqO0NwAkLFbadQuQpgG6we0eOQD+7peLy3XBBrrkl+bZZTPnc4
ovXxHZ7SENInkohNH7OPHMIJQbySwDX1Ot0qFepzrOFtPt0rPYWxj8lcG0EMIkCB
eEfrkMnZnnyPAw+Sl3YCn3K26mfoC9Kc6pofZQJA2xl/IlcQm6jlfoGFxMbyWsQD
T4P0DY0cane33+QCdCqQXEjMuz6/5jpr8vxyH8LT20dsAIgRuP/Q/fzlmWWe9Dji
gv+oszlgF8Y7z4+fhzqujUCz8qvnO2alAo4zmzQTiqJWPA+y3hnHOSluZlRsy0t2
GgWcpAxas9SkxbjyICZJcTKtMr0NjqIMyrasnHNvxCO8oYh0VQ9z4tQjoPnalPaZ
AFhLnKfeTilv38PSPZZmkIO8uDmIT/jPMCN461km4MUTLC4KqNpnUSbQpjsqhX10
mhAeV+H9CkO/VJIC8n5Ndo2J4Re3fPzx+dV1s9u2lHfPHUQbbJ0huMc7lv8oed+W
j+w2l44HFNE0qEezmN/PiUfKIh/debRIGRoIR5CV4FDDNdvoBad5h99ReLtu6qVK
2hIHUCRENdxwDsrk/wbtDdYDL7PKYioO7xB0QhlBtrbu9BHrBfAtYIyZufTqCtPQ
pDuFh2jgGq4KUz14S4OVVa02CO112DXkmAPTJFtZz+9peoqyw/YIPeK9X+wyabFl
ALofuEFRG4fz1M1tdOkXlCuGj7rjQyfgHyw7I5Geett/cfdZRKwS1oPwmdnITwQQ
417EE5buxHqe4QZJNq96NhoJzZlsO3cvKCB/0ZQ9RQxJhxEBARnHte09YSYq7NBQ
ObmVdvjR+NJSbRWv1CRrXVzRCnfpkQ0dmEWAZuBibKU9IPiBtO0AxiuvIHPyvGMp
4eJcu+XxhVfx1Q4dDJjg5ssAX/8U1OBUwXuaGo4oGPfa15YQLgRBYREW4oLWDD9m
eNwiwFWfX5dwFpLZCg+UjOsK07QbaP6wcfQG/0CJ8Rx3fMkdRdsZisioj8+BVsLr
BwQ0tH8DUd8TgSWc5F2GTE088dS23F+0RhnEsuxHuo/x9+nEGu0aHA51qkXodlWe
DmtTieCCGokWsnPfebWsKG//+MBao6WBYWCtjz0m04DOWl91jzBFvempmh1TKCuz
bEfMTRFAhYYahE8nVciTP/6bqs9V4B6uv77S0Z/NP8aoa0r3rXFQbZJy+79xiiuZ
Pm7EgdzNPNsEvP3b0prsMnk0mMAulj3V/DVUogcUubKEXI4kVG7eYp18826GNoit
DVxMgRTsVh9DRUKYw/Y/NRVKKy5KcfGGRLyuLSFHZZrGPbuSUcjJ5ZOlBhsI/MAl
jjNyOBAla8qO1aWdJySmjXPgQtkjPlw5FihPj3Lz7BwHaErLDh6O3GECk9/xZgwX
XKWJD4m44+KxWcFzj3usoJojJf95MJhleVyLnhOKoXmzVSYcOuHF18DdOG0rADRn
7faTDjPvmr60QOXQPXNgF0bn0uJuctRlxkhcEW/8hRhcQB9rqOOyhF+MCTWN72Ir
88XrVw2HdwY7dfFuBsZRScptuLvfPhjJP731GG9vJ2uPsVz3CNLSNJBuitnGe9tr
rrC5OTM0CZPCn74Sz9WD5X/EIzLOQtBq5t+wvhNRysBT9z0XQWi27M3GCYXuH4WJ
OGfSNpFrqDr2SWbkoWzovU/bUElOrjrfU3I64gz0kUWSwbovkW2Mkn92qacr67f2
P1DgFZiHhcczwpnjDthlMaqiprJi20y2Aargyu8wEfzJSBXwwUuTxNs6+1ixhF6n
nrUG28NuKAblNRd0YFV5fItI2vIVyGzzmTdFjt4NDzIX2AQZJhQhrOfJ60s1KGJb
6ygYDH4tlUu7PZv4z7ZhTdh5I8JMhSBmmgyhM5mXfGlSt/3aGZt6pkVQJL6qoB4z
FtDc0adBkHM0hEq0h7ClFp2A6Cnk4PQmmrLTaLGkyLwRrjMe75LWGxTYSgCjahZx
1o6S0gOAWz+HtVpeJmJkrQxm5ePLo0GG1Cjsgu1/DZqlIuD0qlVJ71kz/ddhuloG
OG+FMdL++/4Zphhu7Lam+QuJsfqVX/6klx8lvsKIqwboezzYMwOCjMi1LRIgwp/s
QbWzhoajWshXzP3COrN9WZ/5P9u3xmVK6pwQqPKLpA7/hqYn/x3qRwENSqUGS8Oc
xk1cBjwlSCn5RVQ5QCJiGAUs5vAZFwHk5zTnpIXoEnnpNJoUNxj2+w5xx+19xicE
qoqxsLA7AeFn5wUfSHA/jocQX2BnGpjZn5+/RwH3cg66XEl/ey0aLcxg6a7DK/VR
ln0A9gkmix1T+oB0xOcJ99NO6r7kxjcgaKtd4KWXaLCDOlN5lfOKnFPc5FtPYJL6
SYMcqblkorlBxHDsmLMEZqsVjtOlGA+hHqi+M+LzqSg1hqVx8RtSu7E5JXpd5oFF
IAKAes0yOeNIMPWJHtaQe8ux6IXeE2HCj7BbrdfSx3IwNRHODCgXDcNJINNTbOFC
DcYKCyNbvVilk7xYLVTZ6pcEeLBTOC4kFHOzCaN+bn1NREsqt5wmoGWtjjeArlU1
Cwn+zGvn8P3bu5a/PzyrghHixTUZI5v2+T2UUqvNwmY+HCA56tH86eiP8pa4yqzt
UZGo9QOaW2+JYlpxiNkiLH+TZ106buDui5vijvHX7xGBuBB3u/z196bgnn9kzSZ3
Zqxt+rFkWDPmrBMPiC9abdMazIJTc7LcOmor0k9i4ZgRmAk4xuqbklfsbCUxRScu
+woRHxr/NW0G3sKiYvMi9sqK7jJ1HsS6qI5KVUfDCmAx3NpL6YNsow1LnneBkHVc
DgTdpGHX2pXBbhQlWNwKAkxfzL2M0OQjInpQKMM38poz8Ii+ygqW+ns3a/BiYU3y
X/tOtudKNldiIaaG4Qlw88jrXD7of9UelH50QrmhjGg4u/KIEJdUYzddMeDukihG
ZgeBcqpnAd+haq5R1EucIDvD5j7qpjZzUlkTRN+e7K0bIGZ2kHhHLNsPu2sGYzST
swOxUivNaNigVhY9k/x0UULP/PIPmqak42/BbrdKowJL7Bcy6hGbMmEodg6cz0TG
RVINbvnVbcmY5/PHmOzEhrn7ddO9PKL0rcpGSWZICA5fypXE/Q/zRYE8AweOh+kQ
0kFq+x7bwbgSVa8P3hJgTJswdp86TQI0wYYvS6FKiwKh0/A9y6frQNzlasbcj0W6
AzPO3Sw0emecX+k9YqwpvdfKFqtoSlyarQ+24EVwuJMWa4I9+Sa8fOC2kGRgxiis
uRb2iRWv+zSSmAcEOMb31vkurI7RrxBKkkkziTd2NFW/DzoC9xWOP2W2P95tTV4y
WL90rmWIvxaRXtpePJKKfjJgx//AjiqHb0n148b8XA0QOX7GFS13AxFmsWwmRRIO
tFtiX5oe+dEqtkTHw9wAU6642dHn5wVm1C0yXgsOyBCdQDsWSeC01WkFsyTy05Ie
U8hFBdDUEpxIqHsYIPWjftw2+1SOKKasxu1uxfIcvKVv9WMI08TeYUwlO/Ao5E2w
11hYedq2dsWZmMRlMZaE6s+jRU4ec8fTKXuMxWTA4Sy2UdFaxgSR5YmvArO9bBY2
miigrNsQFffoxOx/4q6GyOqrd6UtjtoEhDvfgPcT4/aybM4TKOK5R45mrhiY70KT
1ItDoTDMYNTzRS7TSQv3JuPLtpeBE9pnYI8qWx/PF1lQCIbZXnB4jgV/SWMRamTh
ccDdZi3sz3nTkvUGvpngVj4OFfywfDbok5hfEpIP4WB3lfVj1YRQKpj+sKw/wBRa
PSPRwzZMSbeOMCf5oAiVogE5yeIxTXK8kShuiwVzlfW4TB1mcq80c8QqyHiR2fu+
ug631OkWR418Y9kAgAf3fK9ypaPedZ6nKLICw4x+JVFKlRoUpIyvAegWO6I1unfS
2dU2nvb9TCU/xOUQzBQFUaMUlaULvOSaqrYXunOWxny22zeEKk6htPbte2QPXTHJ
i/nH26PCKoDfxIM4bSwqQ70779NQQSrFcm/6D1X5UIJ+4ln4hIvPIH2BCygP4ffj
d+P2d8TfSUjXSs2uf24NLaB1aNTeC4KrcI/59c8cqmeoHxQqF0hUnrbyWh1SL3OB
1dg8N+1mJORGpLmHCuZRksNT5ZG+MLACBhb/ZkAn6hX7j2Top2M9l2tLRSGIZtzL
ODcbMIRsEoGWDnF8ITfHf/zDaAR6yU1iY/rA73rF+t57Vz+4kVncsR/LEDXHEV87
i/jTOLd3/JflrZSLnVVdkUfqP/p17/fvT7hC5QrISSfSmbN3vraVebJu+3yQ6GF+
dqxAItLASqCMllXYXvU/c/tbVqWB7rpIqVt5gzVFTAQU5SNLV4ET4Bw6jLQ5i+JQ
lPPOBSV3y+v8UaiAoSg1hzJWN5joN+VyIDLh5nImSkws4uL53xlwDsbBokKYhdvM
czMPmgdYmHNGkNwsDBTRHTlo3MzN7VHiZM62Wn/X6nCIKS63Nyaw5xXDAo7UiqoZ
x6vw/8gvVBUkAe09CR+qmRqYl9QIIvgASiR5rXoXS8a/Wwu+gR1FLMh9I1fB0/YY
AdqGQdQKO89N35nvhftuJCKAt+XnZ6AvrH9mJU0L0C6pQ4m448SiDi8f6pyUYcYg
GvBvUmp8FTHsUU+ULpWj83TlAuI66NiqhtjCtKbReHxN6z9hXtcwjDv8kWzpfEDO
Oj22DuiWxqYDVjIfaKuA1B1GfZxihMLOuZ7TROEZZZ/3YpheBK/O14fo/SU4V6wZ
FQV6NdgMCOLOO3TPvwFt76Qa8WIo6AquKtQcWf0omRMmRklwYqJv1f1l8iLWNOAf
nDG6H2qOMgp5RBl3dfjwYTPgo0LKXmCMPVErGBc651H9rA4XOqA+6dHjo9IOkGU5
zVIEZ0uly0iuALinIzAxaYP7DmZnqVjAUDh1w+0iPiks/oBNiCc0jihn8nQmyyy7
1lW6Rb021A2K5mW1WxeVawHHyIzHO+91YQgZhFiy1RGZM7XopW4Ak3rd3fRwzjgb
YXDWuOamUlPTRH1uekuqfn/REw0mtHYI3gbBfH09d7Z3AAZinj8BJcoEOuRPz5ZB
AtB3ICSH8OJH1LLP3rHv2+o6BAcvagfAhSm0tp8UGAkRYwesbZTqDWrfnmwVKpbh
A92LLW93FFc9A5tFH3vABPecbOB3HOCLBn2tqxYilFRWC0Nm+qhV5bES02s0lIvN
5WncY0if/qXBEN5PC3JD7G5gn+2fWpQIeh6yJR2H7LbYl6DBq9j6hsHOszlFOaHw
dzTchO+PFCbX0ZggOrmYZ5OnFbKc+ZNC03+qwfWnO6HbvphUeiMq0r4mElm+k7Iv
EN1L/czw7ldfToSPAina3AreO1hLI5Gil1cg/9TjGWb1Sno6s8ViK9waJetq4iNA
QyVhN0vL1m6FzXfgVG5GIV+oWtBsZySDTGc+s1bxhaE8qM1PzoNZeI92ZorovZaF
a5B3RHrh2vitwt92/ymZAnK08AYMOxAf94gNuLy1KDWFx6UOjSMSMeqLdg4f/PGs
RGqFW//KvpaOCTMbsPm2iMSdpsuVB55WRHj8pQkvv+wAD0R/hIYUL7ase1mDlkfv
ClCv5EGdH3tGuDRekhOrn/YNhOfV62Kyp2pOTZLowR6HwHnVkRFp/rQAVTzAm3Ev
krbxk8wXjbREL0MSnNjuUGj8sXFvF0kRoW/PCLEqO8y/yfFZ8kwxzkV0ECR3nTn6
PmdX6L04Rdyki5+OPbZJROeyKcqcRDJGL6ETvFbu2s1vboxi158CPTnE8sQxXCHE
eiYaxn0OKTXYBJ7GMARU0EuYz6FYxOn/ZTGMaKEwFGz8E053LV+YCeE1xAgTyuAW
xusgvKTfF+OfdHq0iYLMPk1AcxIKdGgQVnC7xmBTpeWxI/M5d2XdlYuWgwKBy794
GDZVH53oZ2qzvxVykRTo7N/0g5HEWbCuCFXPcZcbTCskgpNNNcLKN0lddbbHwrje
HMyh5mus8f7v5JdYVGhBeEhSJaxna0X7Y6OnLtjseT2FstN3kwUPDusKDln7WXx4
UeArSiF4OKm31yvwghoa9baV+owKPtP/5LgVIV0tZLnpBSFy8qW9UOjjUzyqVZiK
XT2eErfalqbXRReneF/boLrxWNsPXFmaZDVnphRvqdNxHR6h/bbvH+We0H2ZkTMh
MEmmuGxuaIp66Xvv+qvyGxcbTuCGMcd6ky04EytR6fSHuNrOV0J1kv6C+C5NoXGU
BH0nNKpEcYqL1jwgfuXeTjSvAvYmHtjWgXpq6/EitlRIZZPZJs8/blNXSoR4pcFe
nQ7N/D3XPIbbl806P5mweFzc6fS75XwSo6+gJ0oXG48jrtj7x+GcV6yeTxPZyUET
UV780V0NJCkgmwL4UjeT32EJu95djn0GIJqjxIye4B4zOTIFTXqwejFfmbAZK8CK
XXmmYs5kBlGSo+rpgrwDbb8izwq2/O3YHffcKJOR0+Lb/waI33Yob2CpzauVx0T4
HoWSr2W1qhxyVTPDcXiO6MLVwpebnoix7oQfmHKVX+wfMj6/Edwudvbtc0RvJrZ4
sw8XklNJQUJix0caZd037RaK2pG9bLs1WmgtKAMFK647dt+n1nCiiZAKDY3ZGbto
nCIcT2BvEi8q9sXqnqnEPr8l/M22nUMRd6uGAR2Z9sGTb+k3kElNL8yfrlqiTq57
NeC0ExLME8pLE+CQcG8c5+R97VKByQ4I5t3LYCZV3uzG5BDxesZFFpsK53Shq75n
bLQRGR4575XHUEocMqQ94JY56NYFiW03pz8THUofCzqgrlivRNFenV/dN2NjxP+U
6urosW64Ws0z1ivOXuyjL9K4T26uvjVwvo7Fq42UCQfiCo7v1VNzIiSgMONzldlV
YLWxctYhNxc1w2eJN8eoKCwDK/fPlwCGddjqS0LLSrI1REWVKHETbHHktH94lC9u
rO4fKXNniLAqAVX1Xb1De9CP6T1ZOQfaN0NYxxO6uTLSSy9c7tI2HXe5jyBtg5NU
q79nSBXT69rpnQU+4npIE4h+SErBwv8T4Sz8sGB7xNo1RTxADl2cb8FvFgCvV6G5
KaVfp2vkPTOQQ4UaUJPfAo/zIrTgsm19wWpxxX+k/CxaVTgi1ERJRRSbvV7DeD+o
sGgJq/MwdIpwezFaQS4MmiSGZx6ZnsVFdx4ttxDcu6+QkHeZ0hPyYVi68C/eZIAJ
gNx6N7wONzWalqMXIAA+6IQ9nx1kgkWNos5d7ia8NhTuU8cU+k8yOepxlk2n+sIa
YVH16ZgQzpJ4gjgF8lGtLk4M+NbIHPZsp2AguN8VjKt7oFClrYopcS7Yqz6DdvLR
7HeEUOP6tu3WjI8ix5TX3Doid8a3TqSX4mSMs/QaQLFq/9ubz2CuETXD/mEAJ4Cy
4ID2oSDcs4jDNhwXjvSy8jv+nBszROniw+/olhSmUlUVAfqH3zsUDiRYERftaX69
1cinze5wMq+kH1cQjsHEnOQqtd1d5GqG1VHVXmimTUSBXbX79PD9RnejcMBOBh6u
al/mUr+TAZVA2htXykx5TGR8yuDv+gFMj8ckv2ekV/FfC1jcJFjcngHTYCTGQ7yL
tmm8eKO5nvCP33xQQFBKjJ9JgNfrKH4A2hYId8NghVJIU4NJdIXjPEiK5PB0CYmu
8z1yRnFC5klmWUkZQoC/BFcoz+LQe+nqUObgeYs5CcrPofpIeZ17c05CRxwdkcim
C+p/Kyvz8mTt6cn0Asv5j5JWKSh96pdd4H/g77WveA3fhcf4rmvjjYLKhriiobIZ
QMTyJRo9yTvHMVuMfXr9qVmgOnWqD92FP8wAz4YmnZzEn9lLPWVJxMX3iV5vlmMy
4RGkeq9+HaKr9qXlIAXd+rS9nxYiEwGRg3zvpp0Dl9dZvOmar24znr19t1neJ4C7
csCqUu4wXvIoRJFuMMyp5Yzh+3Yh5fqu/5ZmSBnYvVvet9wcGoq/uFtH3scsP5yy
3Y+zAI/9Glsfj3jef/4N+vw5BGuVVqtSBOJH9jta9yeotNP+Vt0xEGK8Qh5M2OOO
K7DU6bwPlPkXky9LYSw3B7DJLMOPqVJzuKWphe66cKcjPkRWeJs8h6UQtZTj2tSc
BtCZsf2dfDK1gn5OCQ4fM9vPzF0pAapKbc6pq4KvRuouvedjMoYPIXsIDAHdOlVZ
t7HMjkQOZn0iixrxUaQN0cfNbwsMPLH67rZDddXutbRpta6jDYriLZCm42lpaDwx
BWLs45a8R5NOlzDhXRgqrlQySTSTt7ldEeH3doXa22J8MA+ioCKw5sb8/l7OkjYX
eJC4qKvK2umIOfdbqejKro6V/wLAt95lB8x8WVzTPkwmHjn+Af0PujuOXkckj9cj
y7OtKREmpRggp/dWFiLF41v+G6ksFpDz2gNb4uHclKJalJxR0I1fBivxYOoVxkUJ
qvRww7EAS3siQUwr3hwGB20Vm5qsWfBIxIRzJKDYcomda3QxgeUxGqCCHn88u5pn
Lnm26b29dI8kaI31+GogHB6xh9cVfMNYdabX3MHTVaEPg+CgY1ChOjJ/PzHbM/X8
6wltcZKi9BAtwheZZ4vCw9ZNI4LW6lVmJMmnZwf898DRHh/9nQvzas5OJckw64Te
69QzXig0WNfzfCbJQrERc/SQ4SZxojCoI9Zzc1ECUY5luU/+DR3J58EfTW5OS8Qo
1itCaq6iFFnEnZPCVqC/B09yZTO0nHA5U5PKIs+7frAvgxHw15/LagvIf61MNHec
CCQE/EQp5YYXInAg8ErHYXXxwiWFZ2qGWZKSzpqIEBCYExoUrzsj9jBcZZfpxwgt
iiVm9kXa+scIAg7gWFIgW1JMoCHqNrvqZARYrJDvVjI+LjQ+d8ZcqVMPJ/NfSZEr
LrfFeqFlOwmgHzbVQbNIWwd36d9byJLWK5L5l1EpCyqsppZRE+z5xI2h4JZVMeIH
aKxC/xRs7PbJ53zf9knDsZ5Pq7R77E1CoqbuguVxvuMFH/O4CLR/BK9Wl6Htnhdc
8zvIEXEnu+RzRQL1Abv6C3kHp3sxNnnSZm98MJe4I0GyUamQNF9lprGiYab9qpBM
OOVI6NtWx0P/q7FrYj70w6N5o1XOM0SCFCEZn7xU0KZsXzueIohUsCdcp5k4lUWR
M3AaIOQZ0rvXwRBLChbYN3Jh7OHftRzyc+qww6BSzZCXWmoLloUo/xEPH5aNr4t4
UjT/ro78aIZQle6UpACFRTzOv3lSpDdYw6G/AMTIJnBwctX/grEGb/2x+/+vcOEp
RyGRr3F8y45/ezBl1507m0zTNMMdQpv//jnxgOVc6FMrm6rpJVW8MN6Lx4M1wfXk
uCypY4RwPpwwAqnwdTWO7m9oyMBCJVCYrQ0LH/UJyRC79JBZsBrDDN3pkJtmFuUm
NzJo8Den3Gvh6C5+oGjVEr4x/VX0SSEWQwLITJXduB3BdHQde/FsB/VWPzYYaHER
LQqjoUE36OO08LJj2joP9Dj52TLGTNHwsDSg2vHfl/Y4jER4mH5Fv+GObX9iZgrx
kjmpl6vr//H6sZ/lk0cOodYhWH7EFr3nB1KjAd0ol3o6sb39PqC0vHGmlLv9poPv
Gf5lAOG16ljxf2V87YV+Q1Cfd5hTM+ujdLldo7EA8N/1MH4bIBuSf9GkAHb3wh+8
klqONPwZdAMXRrrrpCP+epWOhJEGvHEQ6asjbRnYWKFA6MvgQqMEsOzARue6PCWT
SG8qsJjNXQfiIwdeJs5voZfX0go4YtJHpZ0txfYKKrwBXeUENUJwNKIYVIfP6g70
d7wHRZSGRTE1qi08oKNEN0o+dGS7wqgdbzDjyjQKkblzCcuKGM/yf6bSgWwefcXC
80Xwn27BpVuWSuamBfH5dIPRAShKrKiGKXPkcLy8rdUZicYZb+NY+8uVu1H/32GF
B6cQndBQfwM4i0RcbCvgKdS1F1qrOuN+IF0u6PREB64ovoQtTP4IPrV3PrSZBus7
ubnZD3Ko1u4py/VhG1rXeMTmcxh11Dg12D/fLD6CpAzkZqDLagXr1zosLILL74a+
zVSl7ce1xcamxbkFaKcnH7mpfHLN39RhjlpPb6PnIGRXgDPi/U2TPXRCkOuev61b
jpStx32YBY8iKLJ4cHC2diZQOI1iyP8PPzuzCIzQV9yGipgjEBQ4bWswtoDg5CA/
dhpRgKIx9Vce//2B2xJpwp/KDWbxNR5hdOBxTQirbcZdXX1SlDpsk70nE+AO87UA
d4Ab3BwGm/8BNguWBKZgAgox8bXucOYMhHTI7hrOfNtflUYl9HJY8CY4BMAlKSG6
54wAgwyTsrns4UIG7NdPaFFrEOwwpb4YUexcaDdwcnni6+R1NNXft2ejPohY8+v8
GB9k4vaDe7H4jmxsAGof99u0t5fPSFJ1gEGxirVyeKyAzU7XbP+VaLGiG0s4/Z7r
BdIGE+zm3XkR2ooFfwUmnzswirPu1052P/ad7oBmMLj91SD4DRbtN/zgwgE3AdnO
WLeSRvZnGPZcnCIzPrGFE109/frgO80v4AWAE+TxDwvAvk9jE1O4hviWFIdrnxPx
KN881b70ZYTjwkoi6TGLMgx/7aiasqI/tL2zISgpu0zr73nSL4Hj6awjvU33WHRT
alM5pC0WejF675atR4LqLthWFSW0cD3L7wO7aAarjSMoNPlTWx7OUHDOQ2Qd2kaT
sGjjgsx0ksczxe/rZ8Tvoj7gu7/gHOD8ErusJic/RluDdB1dAMkJydRhUjZ6lfXh
Qu/l1ac0AKkpLAvf+KI5mx8vyARowpO47wOhp9bH+V698bQyIxT0tRWC5pa60q7b
sCJbvGPBY4LvVqxbFJNW4K9H7MrgOu6ddDgpAS8DF/A/fkSaKsCkVW0d3pqXk3HN
moFSk4JdY5B7QowYHXLoj1UAR57HPKJKRjeB+FZjU+J6QhKz7/+wXWTbvh5VjtL5
/fDs7nvVdu6CYxxCqkvDW5S5t6nsoDeRipr6NZcdq44Vgs0ENZeaj3yz9gbYZ0rG
neMlJOLYmbxsLcxECwolko160KFHlz2TiTQ1I78aHcPxMiiWJiyetV9UE7+OEdBh
nAaMrCTmmX0qcCkmqR091IRn2ZupPiSKnipijywnvvJXny2mIXhDtBzxs41QiBbN
6vY5dEu3G/WvmT6oiXumgNE8sWL/niD8INukxxB7Bx5BCAgjHdT4bmwTiFtlZXhm
u5fumdys/YdahZFgJNYpbxDGFvxRJ35AmG6SV8ytYwYM7SecmyNZgsonh0pIBXH+
/JitEvxR1syhKvqfBv5dypc91Cc9lsaUmjRqthYNmqMpbejRZgng4hWMCdPk1FIR
wrecFbLLaaRpK4cHj+AzZ8QmIpBKxTvxtNZNxmjUnvW+W0HdC1SgIeyn8/8lplQa
bM1GxvqtA3/zMjEOL0pfkOvz03IxqI6ZFiZqJZoSgIQsCa8eDMncGDgb1Q3a7kMe
SJYY2uooTpPZVAgGjdnKlwhpZqklx81dp2IuHQddr8pG91CS4uwH0Sr6DNKiI0FQ
MVh5npFfH8GJMpdxMfMEn7injPFMfShA9zBeipo4HYoVZWK6GKf3THAOUi0h7YGA
r6Gd8dmHRi9eZB84JCSo3YT1PYjuPD3ipqU/48caXLiLYcp7pKxydVNiVhmRqQe9
yOMrCLpLoT8QVPfbV0Nl49te8h0T1IrVWTmWIzCjRwZyjBXcpjLfeFcUHEUuxGVY
EclD6XR88Ed5BfmIEjl02oUVsgFTkBaKLZgFd06ivDtCdseJbH64uGBk7xAlwd2r
QwpFqugJ19iOlUvqT59dhZLTAp2V5OZtVtOVizJEYsFKS02e2he2KK/UJWXMjcUD
ggqcGa4GV221tfsEjt4Tg3G5YdDF0smr8x8QD7aB+GQBx6mmxnWuHYGtI2XGak7/
HDDzEdcLrqYCAkI8SIc9n3ZbndyLfJmmMVmGfZLowNNHLh2L8K936A2k1voA8kif
R6jFP/AKs8qW0a02CHQOfbsxa+H+R+u5haXJFatoxUJcY7RRuYNzKt2WTxtma4L0
ev/m7mRpWIRh4A/FmVzQLCfvqif2e3z1ztp+tHFl2zFjhxx/YDHNrCo1qJ+I+9Yn
Lkkrdo0oULNcIG06TjHtVtvmXi3IHvutqxgDOgY2OcqNXGbbd2xny38+e3CbiBVv
xITdJgU3tGXz5uVUJ8GyvpmqbTM0mf9XdNbNSHHvg27NVz1qJl1YcAiUItu8KNqW
lGKoa4QZTK/GPcanJqoICXr/BnVbh2yuEukn9tzUlgJSnGSozRd7cnJp8+QGDLdC
nVa67FoxhaVsqIIFryuxOOlj2f7LW5aKVR7nB7KdgC8i3m9vrJ3pP8ENhBsWbnWd
0paLKqpSPpXnMZgMIb2jKwRMSLQAeKvBZhQ0oaVIFAG9uGhNhoJXAGSMPsps3LEe
k52SELo6GaI7gS7+aHf+z3R4AIbKSaNVhGX82oQP9e2TeiQoJiT1XXE+OcHjQeA4
fP82WhLkVKTJCdsY0OWkH+TACg7TFWAQ8yajYSvFRIy4V70H/8T7mFf94tfEIkSD
rmbMgBA6q1W8j8IQXbVmka9eASGDzn9LIHPVgW6TuH1c8R3MYP3cAGBe+B786rOu
ZTqLNCizVGeBUd5v0yhqiJKzsJZWI+RO7nt64ByKu0Yeqr/xMb07t7UljAm+UYop
pVj59xu2frYFYJlSHY88RskGWLEA1OQFLV76BcfwRoPdxjpPrA/JU7uwsmDY6aOo
q7eFJpK3/67d5a6oOOn+uGLkRc4tpPCfNnebRuIp9C7BYX12VZK+xE2W+IWqbMAE
kX7TZliYs1NLVG8LqvdY5oviUmiw6iKSkVDpyIL5JE5Kx+kHdOz5rG9Wu8801kYc
mV6RrQ2CLhjT2+Mjrn6cUY9A0d1frHAFMej1uwmEQF9j68VwY3Vdh4wYoqXCu9kK
UkZswTDqE1ZAYhSDkRcHRAyx8YJ7gSO2BNHQV3JHWHK7j/5oEWwkQgBbdq9iEhAd
3zsD3Kr7/sJUc8Yje/v2LFtDW6//s/vhDyXzVQzDZkG1rN2L3rMgZkxknTljniMw
eSAW/rYlpvZQdtvjEc9yVIBhQMtqfZ4IKxY2qpWYIMOb82dfuSZ4tylOCDgLXIs5
HLCbGic4yjcAhtpLl0YNQb2vcBWNR2yHq3M6LwcP0izYfCsmPZceL49Ag0sMeUij
zBiGj2kT93wgV9BEyQkJgjXWBk6DPa1dkAkVYgU7DNuz5pMWPJk2M6wFgFZ6hRu3
LhlfeWAOe9fr/275Mc4CgXuOyzVUkb9MUf28SToLDp3PdD6hqQIH3B5PYwkqy2HC
kAWyWgJmgGhy2mHAds4IzUwm+1G3fHd6S2Io6S4M33WaPNGymdTijoCivjFG82Cu
QGiDtd1HfIgrYO9HZ99GGIom7wYfIlXoI8KVIA7CtcTU5PJP5V9oGPHd7wrKjDSG
gt3x4e6q6iiPDGLHqjHD6XeG+j2btHaYEg4X1i4CBGjGq1qsF71Sz7UeU18/vOK9
BcqEct1/P+Nfeq+CfUH2ebdfHMWvK6zUEF14IYHVRtw4bCeuMmfMqfTUIumDF08V
zLeyH48WvrSW8LvBoa4UxBRtP8w1P2jo815JJZeDEvRIpcREWocRsud6DyGtDB3q
XekZkY6of5kwi2+B89TXu6baPsuDVzFoYDKDj283PtWhP7lXgpWFpNxcdEcEfLgY
V1RKK0jETjwFRrUzKv07O8fhV7dW5uzNcqL0uYQom+b6B8N+cnvsEaRbV/bYwbPr
eNwWzkJ30SF08H09/SBYyhQctJ02qIQwF1BgKXLUgUF8OHIlrsF3N5BxdMiP0nE9
Rsrsb0NsNKLj2+xDKqP8yQFvbmimIUK6YljotlbQ8ddrzlmxPtuBRBRurwC22XO3
v5ycVkjEskshkGIYgPUTcIQDhhoe0YDV9iI+48LgJb7w1VQASATgdncyT6ICi38g
VSPjpshGU4+K1k1mGXjK6vqUdB7OpqJ3QUYpNQJBw2nBGVoFEchAPNcRYCL5s5Vd
ZuWvNOt8ez1qWkAsCvjtMQnlOMddSPeV/GzdSm1H2edZoQQYv6rYP07RUjWU4loW
vUQRYjqL9YldTx/1+fIJr+TdUwXZke6on8clGkYk56P0fiihwvPDZQh7hcWjH9T1
4sdYCiQoTtvqWkVkHI/iA8bE5GVndSB8WlEdq2g9AY0Nf8zKAf5VQfB6d/2e/Tx3
Rcmj2Di8RiwiJDOz695rBjg/AVkXYO3gTyfC9YDqpDamSwv0DcOIS1A/WtKIu7y4
riQ72HJYT9G8ymtAKgt9AZyMMuMBfVX0dnIHcjjqg4s8r/47BlSUudcUAtkffOES
RgMXiJtfJmaRBq27TRKTP4nubSQ1Y19dOZpJZykGTGCZ+CLIw4z/VQnFZLK4snPz
33fJ7jmEsTXpJzr1TPpRdmemhsRGDfrPe1SG0HGJi/ghcttnJmCrH5sUCg+FmeQq
Xg7HfbmEKYLQvxTV+AeXBP+W4l89qfQx0LzAt//XHWYhH7r3hICxXTixmQwpUnoR
Oy1A+IXfvKygFaaRe6/bYZYCguvv0HJDYdvV8Kmsq9uzqzxyeBDCFfJP27fO9fDC
Zp+J+6IRLJ9IxIRSjzrkPsAH56MbHJVw5mhruaXMuYVtbIHc8Xs5g1sej3t6oaUU
q+gM6fYTcJhBirK8LtlZjOTLKacYQ04Hd61R8evoiOIjPxc6iReAgZ/9DdJkbKTx
Vd0TcNp+rTeo1k/MkDdUQcZRWwJe6Hq3P8wc/1B/Ay8jYMr9JSH7j7/rsf4n/NN/
hMYBmhYGiem3dbMTFnydRBnzeW5l9m6Aj0BBH4TeqH39FVwooYRKNwQx6k2KItkA
10Jpli35x6cPmkDPf8peaJuDlyXCc8XgeyL4EhrT+zTtUhkJrOtLrZ0Q56eE+Efo
6/03xmhoIRj4cR1UR+tuGDT+/p5gZ8P3nj1ObNhTKosapD+7unj2R6z4s0v/93PO
oA+EMUxQpWUW9McIVuyOnSmCI+3EQwA/FXsbVu3p8v/PiCsi/Tmszl30VM/BBJq9
yxrA73d47YsqVml+ptXx+2VFD/VPC6VNlIwNJ8J+WERCDEUW62WTnZ7h4xzHYqpN
b6lip6xYQBRyRHCxckfy3GlZG5lh5eD0solz8YRWkrLs7bn0b+z1Ynth5j7XfvJh
UFiXv+aGZ4JCT0CJ6LX112cxSqL3OHyk3GhMEL2omnDCJnjv4PIOPf5gX0AsfNZn
/onShDJpppx4P+gjMTyJJAjY/k0X7hk6UOh6LPNcSuppdgl6Ohh+IBA73BtJ9HSI
xoycSCOAW98jxXusrS2RKPs7Eg8/7wRmP/ch8SS2aGrXS7s94qtCPoXL50SYw+V3
RafQc58gug7lO0JI6FhPHsAjYaTQomzDWepsWu+BIhPZtVc5oIFEQqVqW2xya90A
0R1HGOoUBJY8LhPW8Y/SHmnU6cTNDDK69kiguPnoY6kEXwudq3gk+yk5kLCOJvMl
/4sfvh24s6O8v29gT01VmYxeyUuPid6w6sqhEj6zCRfk4lcFJwI3tQqp8vJBBgcD
rgd7duuw0/Q0fEB2Bg3RGMbh4dWveyPqWUuL98Dqb8EyPK0/PujNsNS/TPpCJGbg
QU02dD3khtU39YGwHxtrqj9blEnWveAdM68Rx457Dbnq+qEANpC4qmVNSqy7oM/6
ZV4gdG4GndxfZ0mfGmortXa6b7dG2lEOnITo0rbSVyGV98x27NhedZZi0Kc3sh6/
2Qf3HJWTYWfoht9nDlu2CwWfBWCoMkflvlFwyHot79V3xwyN9M1yt7P/kFvgjjgM
rxaqGG91qO3T9ktAT/koBdkztsVeqQoWYIrqribV+AIT0bzmR+gONohnIapJ18Ry
B/bY+TGddqaj2rsQCOm/V5/ohy/0miI6CjXxvWkDQH+pUnvJArIWWHLJFOJNB9Zb
s6+xIxWGzb6p8S4XrN0A7kXocpNqCkwmMLPo4MRUR0o6wwjFdS0EOgDI7Slt/Ap9
t7SqTskOs2qdy97M4u4wVbtCNzsCPpal0ttm9ezkEmkY0xBq2/rvCW2araaFw0Eo
B8rYmMYYMLPORkd0Tp4hsYnj1j7Xr/l6UAahzFUr5+slxj2Js1XiXtrC8UsUDT4p
zcYYlefUxJQUsjydUET6yCs51IfN1xVEcOkM4P8V7RhF94H2o3tuN09sxvfLuUVN
mLs/ij2j27+q5taCkMM8pbVGzR+U9aIybEXePZ+dDkktPB+ZR9k/tm0nBWGiL4ob
fi0EfmQBOMrR3M3E2N49GodiYN21w/3JmVbBeKdxdDoV9fyD5krJNQUsa6y8jvbt
dg3fHt88zZBZnhG1cwFUhQX7HIWHOHSx2xYVcMs8607yQQ/VvxnB3zwf1hHp+6v/
RzqBj5vG6DP/BNe0XzKKUQdexINAStikAU10TobCqXPdAwuw2wSwlJ7zeM+cMXEM
8KuzzUPTis/ZH3MyZIIjnd8SM+yUqojIN+fToLuc2lGtOpy48g+W4kK21aq1pZZN
tK+hKLfKTwf5ukLuceqLlGqPmvhE64fH3dUcMBPZlY1q5V59bV4cNPQKHo1C1Vms
eHK0sjdl/zTxkIhRr2A1w+I83Lk9DxI5FaBjybY1rZQIswMAKvD9h0mTJtobQWII
j75uL/vgOHmTkTyA9ousBnlil6CsVGlixd34RvPFhkcGpBaTiAtd9cH0iv9rumrJ
fzzd75DA60WWjmpjGh8UCOzvg0GrUzd7zLuBrtawnD4tWjfW+pRTkYIJm4QOO8fi
wgFZZ5skRprb+cSdY5v7yMSbegVNL44SABJbc8piQJE6ZLJ1+uP7Bnwq0RL4wYEv
1xYI2gt3HexPlbL/4FrqkyjVUgzTLpBB5ZURiBlZHhke3ed/jHi1cqrc5okxBkO9
GUegGwJrlRDARyA+7uAdhp2ssBSE5fp+86PsHjFrKege1RfLEPsBGiGIshj/exPe
1cH22FPfg2tach8LzzyYi9HYCdcNC/ogYVh+N+IPNtQJ/6IzEdP1elCwSzQE2xn6
BvuqeknRygIqvQbwxb3zENc/EO+6YFiMSoxZXradxPj/8dT1mFCB3Kc+WE9HRadT
hjPSfTRk5SakS8EAN0Vcjo1lDsrwhzlIXCWmXRsmTeWTWv2U59pCXhxIxq/HmdrZ
6IudHhIACBLetJeo8XC1qAVGDb7rmCSgQKQc9pQxKOiHQBZsKEMrNl0e5qtGMPiF
KFecT1QUVVofyHam4UKJ1CuUgy4EmIsCwVmZdVEU+SlVeuQ4b7f3YDT/bNamp0ns
V9NY/SIEwps+1ltpIpFUeIcMQ+nj2Iq3KGlh3OYPGS0eRv4PODXKNrQrPTrUJWUw
zaaEBTGSn2v7UhaaYEVj6HvRBVC0RcoSvS9Q9SSTIuJbBNk/8VCdiBX+dAPmeZMt
fcuzgwThcxilynfT4sfzRxbblzHJ7A51lKWTlAkaupkXSxzzss4objhrW4dGPp+g
TgQhmTaPy0hiuArou76j4qNXCbf6gITQR8JRd3XaGkFUkiMu5MRrfghd3v8rEREq
WDRHQ5MiWMDpekEIpZATRYfvV9vYVjLPkE64TZgHtCGo1BUB1z+pxnkH8b4QMvgi
IzWVP9y05FNkjQzae7uSX0SqFObMyT2bKs7/PlLjuSnaHKBX/jd0U/wy6NHBzOWp
Z7Xj3qDWbko+Q0W3ahj2Bkkx7N1sB0o6fINGJ/3r07RR8a9VUW5eK9MBMW6laZAE
/NZO9NHRCt6tevZpB9c6/3CExNR5r0XI++nwJ0D194h2mbm/zCnPZ44jJ43Sq2V2
VhxRw2xwLZsaWYo1yfxehpXzfuQwIxQ8fQNzNxBj8D3iSTJFC7I/CuVGN+Wk6jzk
E8JV2nt3GOpF6inANJhkXvVTjcG1jRbIiIzLpg0CZbNd/LdmMHYHcoyxYOIHP/BO
e9Ebke2jUI0lK+PR7Twgdc36zGsNZ6r4ydTQ6m1+aJDFaom/eFAawhTRZYQ6YlRu
vt5DN37iW6oyQNSgsfuaGCoiFbNeKfzPUQG6Kg/0u7myoFOoAF6WbZxxBNdKDrbO
jYweqOr/pBKARNxSUbp+3WZf0wTslzig+6A42Utb1r7fUAzRt5e3/grjr3/wkrzw
EgYT8tLXa2TxLV9de/asyKnhL3bYbVzaEpzjPkl/7CwurA09wHaXytQCxQDLnB7h
wyy1xI4mg/tVsH2DERJLMV+pTvkAprBch3HrkaziZrwwGuGHA9/z+hhqJBOs97Ae
ubddO1xE3R115E3Gb/e2JGvv5fdbz7EsWj8FptQ4M90jZvIha9JOGQj79dDzkcO+
0/ctUmDD46mxqdr9neqWZWLoluM7XKw/+uN99xaOMPSEC3c3sHp1rzRnXcM7AVqp
BxGaTbW/NGr5AX58pRFD+NJxm7DpWp1R1V8OmwQII/PpJIaE4I5aaYo6RGO17gTf
TpymaPBBG1mKQ6eAFbOwwArzUVNaVj1ZLubQSD1eqS8ldEmE6hY9/IirJLfu/Y12
XL8TNcn+9HoSD5nUGuSCyEAR+M5Tkoqe+B0ussT5Pz4RuZaQvLSZr7QASlTzEhq0
oMWT/MjLe8zCGQ+3eTDkNMFCeNbeYeN1ChUgY/v1+nj+Rzg2Fy9VyvKzboFur50M
oEpauTt+BzA6SYsjVb65Z/+lPoez5asxo8w/JqeN9CHCOG+e7CVT0ytmlCVlNhav
4B3P3ncUoBi14RqSecuTztuIfXvLLG1MOXU+u853DFZ69eYLZZ7WW/8UpQzSx/PU
EtsrzEmrUT5LBzmAnQa0h4BdNRI5hT3gkxvX7Q0COJSbi3UXSp8rScWdoyrCgdJi
Zh4BuOCiDLDKm592fa633C1f7ULYLqz1Sw4RAEbx4+U+W14cZfDzqyO6Aty51RFx
wr+D1vDWiRdHbI/Lg7kjqYvt0Mmx1xMaEY1PFutLhlTFa2pvem4ALWud7Em3IYvF
ZXnbrA2n5p5zOsqpmMINQdocXDzAXKwPgF0jpeRa6bANTKeiXNnBYXHfwvcvyYzt
acScNo/A1JFepZ7mApZ7uMelP7IL9H+QyAr0np1kswovuGI6/jlvHXtIFm8fMSV2
3Efo8wvDofHxwreRH17VDH6Dt0HWcnN24Cx1wE7/5w1WUtNn4kpuDkLfWD62ug+1
SW7yH6ch37rwm9/SJlby12rgioEm/FxicKPM2d/frc7rCrzKEKJj7UpmjkY2DE4c
Q5PZ8oQo/dQ2nziFiNXfIuGAFBJ0reY9+IEx4KziMLJnITxQtrKuowg/VE8TztyB
FxWVrqApuG1aefE77ROUzeMqvFlRrp4UJj8FBCvO9ZLbuxeRRBW2sicbLgcWls0O
sGiD99gZWRUWt8obTYzzGHB5AMvTPgpqKKo0RiL2yvGFYXPd6/s+WIUjgVnH/Pbk
i4aYSIPDEwvGagvkahF0yYW1+PRHFr0W1JDZdrFKO2+kUxA5g6HcTTWJRxA1vw08
2S2wfSDh+zhtyiYKxLvshhlNIgld33Yb+hxdxVpTHgKEYenB4CHJan4SKJhUw16R
SEdam7qqGEckgfhCNvjfSuxKATE/4cMNHELpOyU4hrzlIZbrizZub198Lf/cvP3l
OtRWEAx+T8w8pNNG7Py+i0H84YkP6MyksUdatPOInCuYnkJnk5DffGmy9LMGV/CN
6vpk4z9UDOZ6WPQlstK5P19XKgn+tfCJpFneKa0qEyslOzY6rLbaAiYh7vLqKysN
5suJAl5Ch3PmUidqVlLc1iNaWoWq1dDCf2S5hsTcfclZ2N9GCcGM2aoi404weN2H
d54muDAQM/TxH8/l5atd1b8YHNzZBqGPHtkR72kWfHuoIcpYfrQ1r8k90/MLJYfY
+8WFdIXzpLvn7fnC5LARxY5srF286g3pMa1UORzhNR+EOxQ1vCnQHV8w3+Oa9h1k
g72YFBCc35UsBOkyNxJnzZDTK22ZGACo/vKHmB0K5hNxp0KzCn2ath4BfCJzbJtH
430CTPfw//z8/xHtq595X4kedcNes9Q76i3qIsN3zaG3QMgm3ykVBw0YwMF16Bbw
cet4M8gA9VC6PkGiWqP4ChxT61wu34+nQHmcScaW8EnzvzuEJg6KgrdQlwoNd3Pd
4MUMpbhR2KVVCg43+0Y/+Q15RV3kiT0Avv+r6S2T8Hr9qoEgdKPL9QpT0A9Yq6Fo
C03upxSIR/Qso/gtD1V1QzaQE+7vOxakQTG1mfGg8IFAyuaZklEoDIn/XchlJE55
p6ueBkVsSAaFL3vq4oG0t1v+iCdettE+ex49l2QAubCrym7pZQ+Daop9EKQAf0HM
hLCKeYR02YOIDmaGkeOoilHgZizXiKqSZDhVCo24oqXOWhlSZ7h5MGKfJ408zNZW
QMe4OE2lCU6aXC9AHrieOl2DzDhwCVEI2qcByuH+JJjhGyldFLx1hLXNpLCAqQUP
SCAk4D9njgurAm0z3c7uCMf81fvxLkZMSAGGi5kU2SxWpXlW3FynFwbAdesuYFYe
g9L+NJs6/cwDpWnaZ4YFNUiADwCfV6zsUv/2QAi93LCu2RPQaFDsK8ajh1h2XH74
DCDabTaOlJhNt6QQhZ8Nh/1+Q5NVsuPSCYmnCUdxoDLUSziQTWs6OKxxL7kygQ0+
bk/VBzvQ/KyrE/tw4Nc8VUz0i7rCGIOjvIOeRojQv6eX67kqvJX+BjvnLW1EAlCI
makXSDqdXofeGLbPwEtjtr2rqvbc7BDl2pLVYgLFRox92vnhbYlIUGL3ERDiK9La
TRD/SOKALEOdmgKttHYjnwaBJMeAo1eVn9v/es8LWj2owTGZSMmzuIKTvaOh0m/b
vqKSlUdSmqaQ+Ck1ZE5/PJsYWvlAxmWwoIVWdN81VVmo0pzgzH38gx1pU67VnMea
PvfeEPqeY6Qg9gjwFWs6AJqS9oK4qpGCZw/nitL3hxsJfz+bY4jiZeYSblrWnsdw
U4d5yfd1wy9OG/ikWp/LVxJ24BPqbZRhNooQgNrHJ/ADQO4JCXHjMnmusqyODjny
2rx9fc5nlDU+Mn713lUKyF7OQnhcXSy+eoo2u+7EqOYKAcKv7My9HUHkCQbEjoKn
CPkfRuJ9ItA1+W2tEBJNfVjKtB/vpfAnpkCU20skeMhrlqPJDVi47ljeibZUy+Bp
/QyR6TmMjwS67kiRS2Eca5PQUuahUnbUwcP0Mit2MzShOP6Uxv+elDccjePPuUS8
H3A7WR4JDN2+0bp6aDSc2rcs7+zPvGBkvDT6r2058EWMFBlZ0jtXYQLfRw+1AFkZ
UaOjPpl/HsgoOx+TAYugLgZFkU4Lw9XCsYQHk/ICLvWzBnWXDfW8us42NMbCw02y
R0pJzAbxO826AFDbBYjxpu/hlpyxn1AuguYkD9lqEeZ0JaWgLUUfDb9TzuOJh8Lv
GL65RDzWDN8k9jmKvnDu7/k5PRYN6C1SKgsHwmzaKn5r39O9wLZ+PoElJcrnZAvl
qfQcJpdkyENJJsQ7n0ejCbwktr3ti0Tnwxa/alk1eZjU80safH988LQP/HjWAvoO
XMinppJfTfwx4T4whyy9SIufPAVKVb3XF1ZaJXJdJ3VEknBVqEFKPXDDMAjTJXzI
78ngbiLxZdRPbtIbVMdQMw1eki+jzY2AvzCI9CWLuBSelXI7SvQG+3eB3iYRTt13
I1qvqmAOezhcm0IJx5v9qStXmdHWJXNA2nLf152NrYtYZUuJ0uDu6XxQM4q2gTPH
cU1UGsouB8CtYfM5SYvATEfNjE9QL5u/y+q5BUoFaMwWLEFgGl1aJG2VZ2F+sIPL
H45EaSlsMYfMdNTc8e0W3r5tEZXcRwBWgzdXWrrJgfoF4Ffo7Zmbt0ST7oREmdeV
B4Ng2ysWELBmbI2fumE3gfAQptb5mNpmY2tGOXZ4n0/UfZTKJCRc1JaX+1RHP2ee
Hn5EMK5g2LLXoFPlBlHLdtyY3zStyzHsnK+GLMhn2qTugnKST8UY5J8pfhtvifuZ
M9MyyIas7ROjmEOFAKHxGDTbD2zSWa7hx6SHbrb0iXxVUTxLUMfiDOJQlfpa1Jhq
ROzYsoDgtlm19FgETDW7QmfP8k8vkKLqiM3DzGE+oLS5PZZGWEyieB85BNaReJPT
NxFYuP24HQnPjWi088l9EmqrRA9TkbseTLIJeSkcmjSSnjWpwPYn9rr1R1v7aVf8
5xCc80evyt2ZQevdZmf3mziPRWZBAzH4AzCg5Bi/GnE+Nksgub3+oIRgZMu+30Q9
8E34sC4S3nF42G3lSHV+Lg6Od+oK3AESduqcGj6Zfs9aKkWVPFbKlDkEOjjc5+VY
eo2Hn3G9xFyIElWNikNBzOFAH+tia0Yv5xGtKt8lnEkV5WT61+v8asM8K8HcLJBX
jPiNHPT0o5WVUepeMuea+Cm+99Tw4LK+aeWhvlayIlZLDNPrgzuo/Oqdqa5Qljru
wSn1lP5wAWQ7rQChqKJXeCFLOEu/TBBpnSyTwmaDblOVm84pXf26peaZ6R+ej3y2
MUiToNhCalbBCamRPN9Sc196woAxiWpOUEXIE7D8VSm/y0TChwSBVNXAjzZ3WSMj
2QZ08fq+f2+d57JLJ8fdMBDmyqM263015JVunhwzV21azeNS/VSRj8vfNUSRVg0F
ZKwyabtUAPkEf14TCYYgXUxVoqa+1Gf2xFEerHNb/bVApJcxeqSUD40aGENWRmp+
vLe1kzgdjMMpay95YrcCeuDqbyc5K8yawJ36FsJRwHRuH/97xK8WG5FaTqffHt3e
0PREQ7sz6Lwsx1P8IU8aPplCHVioKFuXEG9OIrD74rhleINhlnyKCsucUWcsWACT
rH+kY7wlcq9f7EUZYG0xvMvFIjffUJkId24Lj+4uPUy9w2LRfX+5KqUMcXKz1sPH
hBk2Ysrfo3EeVqAuD8QLd+dCWkkwhE68CRJNzZEbiZfTp+8zCVcteg1OeI/IHwdH
G2YKHvh29eKBxGNcH9sqoMeKL/LmQQtkxeICw5mBKjOqaDH8N5D/074GT0k6TTiW
ga4B201/3CEJiX+24sseb86fRcf29NTA7heiWqmJqchCZNZzBLnwfN/PYv6i0wE1
qoBaaaACGSHHz8BUquJUj7Koznj2EPoal9aRMaG37gX93nDJj80DM11Iz5qZ+ycF
rlQepM79E/wCYyd1cgqFdHdhM6FlUgI+n0SGRgupdmegc1ECg1h5fdmCObZy/kY+
QlAMixcy/fftjn5dzeM2/350KlmaG7ADbmB6IPAeILFXSz7lHqo3Y2M+ui/M49u/
2lmWzcoD03MPR0Dk+i5K4f1JMfkVEtpaG7hcCFsVuHEbniOwbwXElf7ucQQ07oF3
2irDMZ5MICWyqAbNyxC+67GYwmHKugm1V16/vkMyE+b8k2mzlwgyj0htEXxKpBFa
xekbAeHEuHxfpaoqqhzf5q581JXGfNU5Fz+cW/06efltmbHSFBs0Vf0kzP1lhNfq
KEWo3d0+f4G53JB5tVWWGgalOxM5UpWk4XbX/iwOyl2T7D0YNHV0smjk3EzEp5Wo
F2ZT9PYLm52tvDEfZRZoupvsusfROZcEwVTn3FWVL9pVvCrRWJINCJzAHjfV8mEz
tjOe2RWJzD+fMwsgYq3w3LuuzaIE9LLYMcwop4ZeMilriFs6aFSynR6gSJ8yHGlA
VjgPBQeUvIrTbP0csFR4sO+Za9hapZIdoVzgMT3a27byjK3MX4EzrBr2BvivGvTQ
GXdYIK1C05FQDB6ydhei8hdQvb29zgBcm/8CtGxNSKWTr9bifWu4p2GY7iKOnhhE
41Z2I+8yEZ3xRQiUy/MDVKk6nBEqFRyUS3L4JKkpRJ9vTCfwJUHK+HKYV6QgG9nv
RmxvvBjJCzPQw+MzFsUzVWQLlLH9wYxEaHBtTPAbLM5H+SrR4xdRnJrxlvrkoIEh
xJnGyjF5KxMLBIjLO0mLJwq4jujPfrp9OWAH1HGNdM0L6fyINmzKXKYB0LP37m+V
1U4UbA2S9bQ1V+Ak69B87NEx71aOZN9b8ipeVYJ7uSPJ0Uij6ow4YhDgIL9wE4rB
sxdG6a15SiqC5ha/5+E3nlepzxuUC6aD0Oll/+XCftrMcOPbbfovNKxanTjkqLvl
wHe7qscJRb6zrI9E90bG7TCqDQCYYiHLTXgKKPlo+WNJE+Tk5vQ2r1izO9GRpS7A
fF3XYJEg6lA0ntxhtJfI53MxPE9k3y6mTziRgmHm7L1cIF/R7f2sO29Bo13UXizd
mpO3K0m9GNVH+8VNd2SOmU9eyhL7A+h+VRwje1Z5lqYmfbWqQsYo5ekKOVnC8Xat
8sW7mUAq4nZrM676K4ytBM1CXl3A4nYyGu7HMTa7KDnFXTpJ9NqMbbPk2XiknFIc
v7R7ecu524lw7LlGoUTa0/0L6BKpdWjZxGFeJBJYX0rRWUc+zR2H2F0ejiuldP27
8g/XJWXwSxQ0OpsUcWBWiW11DiVJoZlJBCy9OF3ozviqdLlKwhylXIdjBLBrlRa8
+p4ParficJXZop2ayT4sVaeToFrhe0JIWxHnLqQYjneESCFVKcMEgaKkYtB9yd5f
pZTDexVpzzwLcvJzMMSOBcnF3j3ky5ms9a7ms7+dsoAwb0s5rRAyBHYXTdgGfL0e
lbq9YH6agqOSkbATrm+k+lDhdMb3nSvEmCBRBsJEbf3bTtXc4zHArSHlcxTl3HZ8
2qIRIsK0btZcOyniM62yvbPlXdKz1TSydprRLtJWiN+opIl+emKGn+0u7SFcvo0G
QUdz+pyrP4vxynR9zuiCHjHYyvekzHzuaZ1LZBAk8f7WGYLtzb8erBxm8ziN6Ywh
njcYGLPfa96JYH4XN0oe2fAiqvvTCU1Tabs7vS7BanF+m0tyOzpD108OuQhDU3Pv
+XD9bALCPIraajrKjqmazUZHVk46jrahIcSKxnXY9nX+V+kWLw6WP4MGGBQRmXX+
JwSRIlqLz0UvSOIF4xWKzlKirLWbskIrAIzC8xAK+4xRIi91RN0Yu6Z/2s/VeBK0
WuHJhGKtPmP4m5UP+/rTo4/q2H1tnJfqifLV/KIUdSzxCOvGKapeirRDYRuVIW1+
euR/AvFO+OTbmhQsuMSUJEpoXZXPhWI6J3aLyGa+chQkf2RVYY8KX3FAifrnIYVM
xLj2zqv9q1pdEFQrOiGQ9R0+82foBMYD7c+D7odx0IklUYwsNPTRHot58rGpjA/G
IHjxmG2EPz1tase0J7WKBnTcDPJxnQOrkla1adyMSVmJsPzYNaAa9viBaXyRVxmM
50s8DGRhK8T3Kr3AtG1J9DBzdUuZ4MCDEj6DQjSiEkKZHupfPsq3yMFAa+vhzL4Z
LWeEAHU1p9JywvpnQWFUjcAm/zVEGln6tISTewxsiGxPzM1opRoihPmpszwi5N/W
DD5MRCuAlo0Fyz7Sjq2aS+UBs7jjEIWNvhA/qu8Zikz+sPdcFS2cx5CKtPbN80Kn
EJ5YuoedOixlgOke6MhLteNF5jAZ9+IBdyABMmhU5qVWWF08vXCy5UAfR6/8/3jK
MawwMsqAN2H89laKHXVmo5jty6FyojN8k+8Rjcg1FFJF28mlvqjDIDeWf8ZKFf/9
TLDVG+tOH1SIaye2MTaspF8egvEOEWeIQ1p0hpLBkVmSJiGH3Ai0MYN0K4p2AMBO
IVquXKKk7vVPeVE9m5Iay9QDVKH+HoNHCd7D5ppLjBa/RKgFU7/69d26zXfVRyvD
cE231rSkZj1L6KzcMHf3MjZFo74K4wVuW2moFKfi8ZqiUuR8tca0MZikGgyZRZhm
PBSBVs4HG47OsWWfCiann2UcDpOn8alenbXvbtOmuDLouJg5t++EJ5a8hHLGrffa
BjGfbqJnZlutkXIh+xGYhBJxDbEhs+8GCoOuHu4sKo9f1D3jykpLVSdUvIvWgF/G
9fzdPYy4+rnG/4EqRXA45IedWNSvXAat+zrwwlLpdbgtvwo9PUP5ccslCMfX32YB
p6DbX9euBOGagzHVQHWhX3lzj59lAImxNGq982lwzacaZ0rGS8O5ZF2Wgulul+Nb
G6eCimNsb7sDuBgKcwSNxu5bMOy7BEHR6bi6j2tmL4o5t2ANHChDGP9jsrzjsy6s
UpLiKS5kd5j8rV3vI69X7nxz8aopYsr/TrjQrgPFP/k76OmYDhZSmP6cVIsTSIrZ
QXiYdnFZLRnVo+O0L4RIHwjlCRDN9FAXyp6sP+KlOwnxffFikcfsBJEqRJJKDeBv
CxPorvNtxx/asOaPL7M18OWDs77xg//8yK3167iitjDXTc8DHgJivLHsfGkCkvCD
3iMZcCie3Qun/zxgt9WJgxGqeXt/ZXHw5Nq1buSks8QSDNdoDUSmutHXwvGucCvj
tvrRHZO/ArRqAmCjkZi/tiry9BzpvoOTSa/4MRZrjJEsLxyybUvUCOZcljsZi9DG
eEwuMu7gFr4vayS0d/adwbyTyz8BrnqSmt8vfv/Uc584Z+GdyCRjNY9nBIrApBhd
wlDZ/CcT2UYPPOCB8cKLgme16PgtlBp4UIUErkL0s8Vx6FE4ZsaQZfANyPkZb8Xa
J/H2+vG4SQw8GJJ+p1SNJKPyo2uo7v4DXbLHgSDq1UABXrwKaApLS2Ci/AK9SYk4
bc7hJkc59WycBvdPhyK6VhzC5xHtMO86kc5JJUypv99xPwqkQHN774egChwRDQx0
8FLJfwMfipGSL1VrT49wJ0TMEr8O/GzC6XBXv3vGhbKLP7HzpOgAox08g8H63feb
vyUcsdDlz40M5HwB6HzJsb1ngLjv/9CC6jEJj2oO+RgTiuUadHAI0rcrp6avDguZ
jYnTnLGDeJnks3wjWhmG+H85sa+TbLbXF2PdzQb/ZtoYzwx37ohsiie2UBmSfM2Y
qNBQVNKr3yHiTKB8yMpJDKG+bgu55FAdre19k5uKmzF/TlERg/v9iUU5hFgZo1VQ
3QXJShN0V+tiSZ+cHqQlq1ZdEiB4LtXM4htnVMTb5PaRVjKvcyesBczN02au7GGL
zR2XDQrah1vKbl918Xf8Lz8mlNQjPuuChzREA3lNJWJI39cV4kAsCcMTIv/mm2tb
vxHIchy6JuJHJ/0kNINEW+SrYA0PvR7P0uRYq22ZOEGrRFBn5LOf9CC3+QGN0jQv
1NXWzbHasxiGMqiYiK2HXjQJIHkY8feqneHD6RFuceNXGNeKkvcbRyTQyTXW7Bd7
g1LSvsI+JcZlfo7qYcFUf6FL/ZPoBfloy+DBQ48zNhFeGZjq6wN6KDnsUhf0fmzW
MaEPiqDFQt08RatCpxVOs371K5QrFI4xDceAV/u8yxbHWQuNC5GeJ71/X/ojhA8e
1Xxk0bONrie4+5DjcCGt/Hf3K3CrE0ZtNl/yOfeGrVaQYScB0v4LbffhwTxxuk41
4eHn+Xtt266lP+6nwdRjzhVPy2P5seeJMpKptnFnA1PoL99L09R3j79AK61yOw2X
9B1ysQHn8V7H/XJTZFVtIhq5fmF+67iGOBuSR3YRBpFlGoSa8Vl/JRld3k4jfD43
QHkX6ZfU/kiwwnZKu45xM5RC7tgTDmwnGdt3Irea4e9dSpl2oXjXuzOI2muUPxTT
FgNeN9rJPOudJl3AnoyawtRP9FPu/priC4docpNrB/+Br3IqZAbpZiJQg0DPHy9T
MdfBccW7cZWUDNNjGQEj3AOM9ODFQcydXTSsO+dReO3GU7ukPq7K10QmyxjJFV/x
qB1Gd6nJqOp+hadVnAjS9ccG1X1+/1KgNUr6kryqZ2gfUUw2nQvVGxKJ9OvCM/jW
u2Ut7om9rwAKsAT2bch/GjyoIW4wCSQCiEcUrJs4FOMDip6p5wy9QgxGIFcmHoPC
OAIKIoUODBDWw4kPHMrhWhxlJZ31x370Y7zKriYTDePTyLFGZXjuYjEJwfUdFBut
cyNfTjS4MuWowL0ydgb0McbpMESnsU1p2voHo9AkKgsJSsyQJeo/TGf0VVJ4m6z4
TlazUsggzl/6rMjvfhKqP1HcD1d30FnvwlRBvBTaIr5QYTKxjXaDmBhccrJ17aOF
u5e7gNLzS9BVDtVXq/ksyURqEg17K3XezWq5INXGVMgzM7IP4E8VpdFJPbpOmDQy
2W9IlYlAzKAburfNxyqq6bvCIA7aYmGtaE2YRCb88CO/3YHeCTqCmsEc70fGyGXo
CerIj9Zgp0xJ13TG6Acb3n7pmug29hqQzXJmCr4/gY26RTdQeoIXKwfE3F9nVFwV
8Pr+TCgp1WHhH3Bx+4PAG4pVQgVNppiCemgqGbw1jC3LDpvEf/xuan1KU6ujjHXA
ws5wKdZg4yi9m2lVj5cqmuFjmeSEpuA8zhTWtPYEpKyszwm1rx3AhpIu3eZTrXtu
gWEsgCy96kSrAiz/mCYwCsNRp0S81Cib0c/EL4kEnsqrquJeh5nVTL4Z4x8OwKBQ
nkF2i2LnDhwcsgAOZgkF7qpJiVZH2Pzh5Cef4KIapIiwXfziKiHPXH7r72zQfBM4
gLbhIb6exNgghhNqeX3b8OwK6ZDJAqEnxdFwUXEykpRZRAz5bS5SWYASwRCauJde
l3B9Cd8SnLrbhGpfIf3UMNsxeG/dOj4JOQr02r1R6afMsh0IPW6xKbTrw5a+14FC
rZXH4FaCFB5JzhXMZB5WZSNivgrlaD1Fvy7eIq3MEdhKhMdW7GbOOWg0S6I50cKr
WjXpvJUsW10gJos98UyiVTUhZATOODM60ldQViDuvQBEHE9qsVhmRl83p9Ye9Xko
/MDQ18jLW9RDijgD6Jahgmlp9MESJGZZ798TEzkXK8kGNRVxQ4IB277FfjJmP4cf
jGPCiqs4T7nzu57mlXDLuxD1QOJQpACQjeSlQ4bUaDaakweBLwxhYwJyCjMXSXd8
RVb7OxiTS+Ws6Iix2r7FLnGPtdRTZcY0hJhOIiGWLqteNHBK8QyfNy7SZJaUjGUK
o0LRgLgiThwaBj/aU5HyEY5an5jq6sYcFpYLmxTXOWjcWAClUMZ2tvCG76YdZfHF
v7JByvFnzBZKUViybt2hoz1u74ENdXORzcqXLX3uUzWrqRR0i7Vtt3OuK4DNsNQr
vQIBDEHV4mUVPHa4E2ascVS8xyW0zpD4WQxqJbXWdS1pNQostyzr7VXQr3hYyAhY
5MQhal5hxWsn3kUANNEbYKfsAQIubh2Zw1QslzXDp2cSWjsCWhLuFuXxkvtwOagj
N2l/SB8epBc0dRkrFmEYhzBncMyK9e995OSy1ykKJapgIUw4A1toY6hDJezmCeDw
VZD+KTtZ9BUKxfPrEUPu+o+MczrMZ/Q/9aVdKkkCuETuaQUGiV0RRQ3tJiTNCqjI
O2QoRUF2s/IEjoUTh2uOgXZtRiN/BBGj5C50UvOXAzj+3DaX0ozlORBjkppP97PF
wQac8n/IckV2YaUuJWl5fDimkmmJUIPSdOBXE50lu/wjRiedbxJmmxgrdv4C7+lz
vYoIQx+TJ523K815/EDlFEeCTfSHL5lc04v+tGT25iwhQ3ppKrrexIJzy3xHQy/s
OjNo3mJ4eNkSBJ0NeFrIYPK59ulHr3G8HMbYfLfQL3Gb7lEjL6temVfaxS0M+0Kx
g+8oy+ewKpwlH1q9PgohgmeaUNa7ymjjhPf8ApVvo2wSsGytuL6LzX076kpzIzn4
MLH9GdnHVK7o+ucXDw16UIJrDRHdunTO8lY7Yzq8AmQ9PFmnOaO1y+84pq0UQboK
mdjpJYdV1sjaTn/efdwN61xh3+6+Dd1sY5Ub7ygrWYjvXLkgTTN74zjejas3LdwV
Q0iOrqBRCrwHG1q/Sa8TsNHCaPIdR0OWbNC2vZs1CmlbMiHpoh527cXL4ZTRKGRn
MildkiOgEJxEQXbUhIbT33qMhBCi/MfnJPG5P7rQ/RGxMzqar0Xb+8/Hmgg/MvHs
v2RVX070AIzPXjeis03N2hF0eko9c6bTo7+pCkQc8wPF7DWfav+OdM/PltoNrdhU
y8BTHJkXqWwGH0FqAjhlbaIjvmCmhQ75hbZNV6JUycMSjKPJ9lbkx4R3gZ2IACHa
mGFo0Zgn0aDMan5uwt6/4MeT1vqkznvmdxyjYjMawxzYpXtAOPtT9rb4L3f53eH0
OiJQ7hC2Bw87p197J+KMXotvbvfaClwLPlyGbWGEgzq9WZNaotDawdfDclIm3pgX
WuFQsvdHsSNfSfGcdaNSUuzoxEk/Pi9rc4qXFCY2ZuiWEIGPPXt5L+gp+GhtvGLu
suNFJ0iQR09A/XUrYvr6jqBnp4I9IPdd6SyIqdpmDZ8EpT8sAJ0uuXew0LA64/ul
MsWFfqLP0Rxld12p9YNsby98Aie5UMQHx705THgqTDekd51OiJs6oIFD9L1MCqDp
O9rjDIjHKWc2xJbZBsdoencBVPSEHdPLdKKPwgE9pbcD+DTBzMddchZQgi3sd2cX
qokDgbGtCME9mxyH/nHv4lc/jD5jo6vAsQgfzB3IcZGEp1aOV9I/xNm/s0MCarhA
GFIvBScgO1UIyXyxG3AgB2rQzHXScFzk4SGLOefyGIXgp13BG7gDdfrt2RYKFx1d
BqlC2lBEeMfrQo5EBt6NRce75hS6zhDotzh8j+N7sJkjyU3p4YSe1xTbFg3DeWMA
vYxK9XwEE+9RCXXdPVeogKQQpcHkXCNm7NIrDhmWqCLuMgNDDB+7E+ownLFR7hbC
YAYqmSFkztqKWTKtVkF9EmcjK4HAZnWi9Pw/LEEa19gpOir9J1fd8XpR6sABDidf
A/df/96PN4ijqXwWtF9hROdWjvdMqh+VJCJFDQlS4KCz8ZytDyx7EbV2mnXmV7/O
9/MdsLUQofY6ul/bOTBOi67B+p2bJ69ofOwq4E0/quFSG8T6EippAVnYwcpC/TTj
FV3u59Zqv1NSap/8adwgM94MPgjZrg4bYBXOxlE8c/wiapvg4RAI2f2wSvvLsMbD
EpmZ5AD/sbSs+qYjK2B3oyLGZWyJIDSWwxOXg+6It0vuyi43ncEakY3UiMToY4iC
UcVT/SO0oKwcMEp6zv46lxT6bkH1xonfB+RBcN+Oj6v7PoKJRTsOWpb9mew13BIF
WWOEEkaN13tncAxKwgP/gRotK6ww2YfT2CT7B/KI3Dd/nmZDmUb8ehu/D9TXnSEZ
3OeHUq/so1y5sfuqr4ezF8HLu4TH6r2ODfj3fqAPrAGULKGBxtf8j9BTJ2dDaO12
qAeo0rfpRcv8ro8PqZh3m5FiO9A3Ve7jgY9kLPUXJYaAtzV8y6M9k3SWvhT1Vj85
cKYlJrduVHnPmf3iVbN4ZXc/eTVb6dOO/IeNuNqx2vzSaEQVf8KbydTic8nrnHyb
u77rKN0ZX8FNF7KLlxal+twc2Xq4DfxBFOjj49i8oiW/C7eIX9Vfnzezx1XrRsSv
r6LqhgfW6mlUlXsHMn0lwpAcwjoDI0QViNpqyPtkbgwcUPe2Wmb5Ao/psAqPrEhU
qXIeZ+krO7A3utxspW/rvdZVlj2PzWnuUt7YEnBF2LR0M76TzpkT5ave6aEUJ9oE
uW6457MJyTdeIxJVjnIpNx5SyUjtSntkLLJ2y4vaAjkM0TaDhbb11cD8j/O/0sPt
xkjHsXwCX03kEetFLxkG6YupwOr2rcxyTNnc9Uo9n7HnSGa0qDQJ8pN1CHWUpDmg
Eoe5IPPL8WWafx3gNU2eWpDfgz38CjqczoytSlNP7nHqWXbrLRbSFiphnWa7EzpT
hvZ2qZb3IhxQ0I3q2fnkxqCgs2pFxbaPoNYrGnSXC78kxcADZgHw7h/uyeRmUb1x
V0SJp/yFKxXtBsMgfx7SEDO0fqC50ryI/cMFjD3vVcDZ5IcQ6cFuIhpUKQP+fpLv
nLl0mQG1D7zUq9kBPKilneKDTMGMNxSTDbgehJQgdPYlMF//bZMjs3ixjEm0S0Yu
1cFwttDJIDzbtlrLTZonKHdcgmMEYzWAG927G2RPiW9a2fyFHhq5ikHiN+GWtAne
dVQ8L/kF99fOABJ4v4vlZyd2AZLiKMpN06uUQrixfBGUmmF8bClZIfY+CUrZ38Qg
+Gtuweqe6KmShxaac872P0WpfkqM2YlploEJ3ej8LZCzh31KvLVUGBJ1GnQ2T7oa
zGdKNEUrJ213wLTDPXzm4TMn0u+aX13C9vn5gXbg9hIES8pW5IwroV5sl+Jwecf6
Vrj7BZwzNf63jgNUcjIjPRewab9yX5F8uT0UayzoVErtIt4EOx3htpIVTtJxBbJ4
EbCGX24fMgX4pE80UyU4el+qw8UhZh4noB3iS0d1V1g4et82hrkVD90gc4cT6E4N
t8iUId5KAxrlylsBfv5rZE2gNeWhm4uPMcQTTB0+EoZZKvSdtbFug2Oqw3o4a/uq
cvHVLjMAKUapKpW3NckT22y5NKEfwLKOYM424Fzymm5gRTfFu4ptmufPItABSjqJ
hhdFyMjI9SFp69cMt1Dscb/DuOibYqVBotkWPWO7D/aiWKbJr2GnxqYY2LD2Ixp4
smFQJC82r62k8n+p9ZNgCCN8wpAQNPEEye4WSdXEGV/ilA0QF1OFPWDlKR7BIe1/
NoRBr0I7a5QyQbILo+piClkRkhnNWy7SRzKwi73zmyyZN6N8NO3z+Tx2ZFW/RZKM
SPQSyGx9yvxlQoqViDag11N4QZ1n5zlTVpkxTl4L5MefOAsgGRrKDxENGoO7Z9li
nbtxsnkGQI+IfhK3DAEjb3sEFPvUuY+J2hyQEGCrao416QnboB2bd1kaIQG2/2Z5
2uXNhAM1UOA5Fp6cbZFOh5Ki8ntfmdlqBbKYNFHNOGZ5rEb2lKTiSEF78L54GwT6
CLwRxVQXvXIS9wcKj2Q7Bz8fNAGPoOCvnrvRgO0Ra1OD89mjTzY9nr405SuEqCv4
/Al+MA2PZ3C5OemhJLhB0A83R9Be3KNf19ysnVmo4P3OyCeN2GOPB+AzOz8REA7+
S2GXDbdd5J450RHlB/+FU2ADURs5yyOxxU6KNptqnkppdWNVId17JEisTU+j6WBb
kzAKAM/RWtzO/GpvI/FM0C9pitBrHUex7NCiqpK6KZdTjADcwoxI9CjXGyQTfcaZ
ci9Iq4lNJTU5bureehH16FOC4Kv5045ukylmHJBjdYBlIiGENkYXOR94L0hCddfp
ixl670xaHW0IW7EXelL5TmoWp1zlZo1OLEqCiQMbn54+2oUCXZ+mqUcdn4uZB4kH
lxBWkf2TzCUahkinU5f1mqHTjB4yzdDcBpNGe7XX/rgqWR7YFUMLGErTRtxBKzDN
C3TKuQwS9iBy1EAXr2qxQ5KmNue1vdtTebk2p9jqT02fXA0RDJxLtHvzCHf6L2yQ
rOFy7obwxXiepj6Q9vaNf4Krwfc/c3u/D7IXhjuBaHmOIJPqj+YADYUmrClhJTTj
lvo+GSsOzQ1QsKuqpGlsuL6n2/qARfALhGj2UyKOL3x1K27ujMRf01+4/hQ6XHkX
+8PlSWI+EbJkYorDm1GgcqRU9jF2PcMxPhNZhk9M+8iXytw2LMMqdShDhqRJaXOd
eSqWY9XyvY0KYgBirh1Z9ThkN3oZym4crDxmLlpGgWN/I2eZsai3pnBbdtdkEuv6
fmaiJdswoZGapzuVCoBCz3vXB82u0n5zjdbzhExIUrHWNbomT1Mhjvsa9sHyBJRo
jGPzeGoLZ7PTYtTWQ+Dhz3YJNJ8+BOb9WkoMhVxGA7UtA/jwSL/IMK/ny/WgRuyh
I3lEi0/Gp/aHiHNHtEu3uVnI+0ey2dy1djTgFONAlRFJeaCkNNo/j5MDjFqv/Gov
3rlTkx21Zi4FH3mkuICCUM83KJRAirlwI2swQ42W3jr4kFsjXA1pO62w15/L5FCU
jq8v2r8vQvClReYLCatR0KGzmLIZ1f9yagYJHwXnCm/LScIiSoMMqVvNXLctmOZf
VhvvIH0CFJgKFsd2TEKpDnghPwMMfi4B+XxPZF4l6MFJpSeJIPcmWUEh2//KkGob
ikmna7HlnT7jd8t6NBeXF6SZEzyPQoT9e81xSQLl9VubCP+5UT0efeIkF1kxmPHK
TZ0TchL7V5VPxzD91Rk8KWykwsX13HuNS8MrKc1XgqPfvIyLdP1ZAqBGTLGkG7Lp
uWicuElf2Yw3gzJScCxmtu8L85EHC0oEiz/quyJQM4ydwZCa/owGRwAqeOd2ft4Z
OPyeVDmKYccvNnZ1cwQsUTigZkzr+xiL/91pe+GBPA9HkTE1cvC8DMsR6ACJ89dw
P2+3ysolrfTjEgOc4reFW6tL49wpWfSJ4OVWCPsVVVFQLdTdBU5BLW7HRTSaI/lX
dDYJGe7l/UCDStuK6ojXkfATH4EZ9bJwroHmivEOoZqElkahim2QsSDyDpy7n/d7
oEEHg7HL0uoVHebw1JqWl0GGX8c0z7jLYFW6zwNFS7BuOBaKLMoFtW69Ne1TWqz9
4H7qw5qgGleVkdcNxdrIqknHXYbuFlInwq7KxuKsAlGtRrVM1dH9CuEuZ8mlxmJH
irOR5J9w5V1lMzteNRsOGv2xk5LbVVLnt9VOEl/fB0v1neY1zhgP353i3SUKgMfY
2trreC5dEa7ouuLnhosHBY2ZuWtE4J4h/ab4Ar3c9a6yd84Gt5Vzd00RavrMQSTv
9tBqLpXnCY1FnDbz+1e4enWuN467iI68OE8wMyuXbtxe2MCF6C0Iak7QPqkFfyXi
a0N/5dqT7P++l0i1suNToLuafcWN4BnVRyeFe4t/LaejaVfaZM/vKqal3GQYu/iK
l+dLUrmdpFRXXTtSET4pa5WvBtP2dSMekEbKoNWFIVlu8MEUPCy7BP9bAyJoMi5o
vy0Xo9BI5OV1LNu8Fl34ngNX/7kRN058LeFyCs46frdPKb9ZHRhkjDK5MTLTmXCw
E9ibyk8q8I6x7BtgbXvwD6o1WRlhZcsMUDvdFB+Buph+Atw7yZ7YbpQwY5zEFkWi
i6LmSLkAQCm8Z419oQNnS5p/Dl8bsZod1yDqEzrShf320TO/V6foRaUb/PGavQHv
G5xPUhv8t9RfEzIRO4cKDdC86yh2Biz7nwy7mD+r15w/MFeFoG/iSpdXeR0FB6MA
bkULTfw97LpOUmJoH8EP0Wz5jUyQPZX380t6Y/SKoMp3Pn3SUS2gDtcqKD3yLNJX
GruyATaKYu+EmzfQJyPeYq4LzauGbTobnpu5hSYnN9HSrJePquOx3ovubVFNj8CB
/gnLJn03L11CTLHWfD1K5KWIq14csT2Fs0J2/6HauVtOK7wO2byOJPZFcEiNNyJe
L+rSn1MHJn8aLIqNzqRSuTzVmo50BH0SeBxJXBqBkw4pzX4WM2mTEkh2Xs/V6SVx
lRHHLHp/PtOv+V6gA3JLTcbQtTsmPPfVXgN1M9qwc9J0X7Wdg/p7O9KDV7g8FocK
s2wZj9SCjJPvB0DA+dRk8WVtVsPSGI/5Ha9f/ILDx1ckCHUzHR4J+UsYpiui31jP
SYPnFYT2ZoOIz/uEzNv6Y/fhuNU87No98ti5c5qz1IXtTwv+Ij3mEy/322546RkC
CleBQ55T+wW/aHxPd4RU+009XiOVvj7wd0RpBrOmwQtSkTYhxYYdZie3w8hQ2PRN
3zjMhuvQoCa2gg/jVPDVZi8c5Ekv41kJXZsqkkKMCVx1zkc1lAQe6qEKG9cTt+Xq
eiwoe+vydXpV8o2D45zeNPShM7bGxx1iI1XXRBUCD5YKavishuE4oLrcyCiarIJX
LJUJtnu0We1YRbsdW0YQtncQZiYYHeasoIa2i4V6GveubLJrOzHt7j9ZqdurhVTI
+0Oi/W2ki787+F+y3NO0+4LjuSNYa2EiHRHuY/VSag9emjVPUek2B4gWi1bNneZA
IEyWJeb8dCp+L09x97RfcKRM7eGbo7uk2e0r94HQwupykE8qx6EsXpH8e16PIBkk
V/rTNg9HMvKZQ7iW4dhdc3NVpYU+7Myk4JvLIw4PWLGfAk8eGygW1soTWNG6T22K
r+fNaLJpXOo2wmORQmsBMQZxLzvE4emz2De2TBwy/eDpu4avZCRo5+/oiJ2ziyu0
5BWpZC6uof3JlkhMAC6Kd46foP4M3Pg4GvPBayEQeso/KOVuyg4YT5pR21/zvRLT
bx4n1ekMJ380rdjoUO74muOETu2dl3gm+UXc98O31jm0hEFYcyNEzw5Sf7m+irhN
vy7TjVAlvvo19HvdEpPqHVn6JVvRoC3Q8UIrBUZEC/+ggNyvV8/KuDNkHz4xPHwy
99bU43VE0AoJTVk3xE0cjY2hObteQ7xwB9Hiqi2kLM+42EQwex46foy6Ffmf4h+/
KFkAS/A7+y0rXccBpsQn5+hAAfhgumw4Q1fchwKFXSApUfF+XGzCs2+rqpuu/rub
Nk4KHEtRmCrQ+p+jVNuYFLwx5TPrNas9j2RJw63Iy6ECuO2xZHYYgCUPLihhrwpj
ekndMnFl7OJS01RIWSXt2WrqFiVHOE7IB8cZdJjNCujl/ig7q4ZSXn20mKdfdVAX
8CqETbdofzlLcgGwvCWLeD/YKYbT6ojwwtQuUYw7dJdOB2VzLO2ZjK6DBHmtYYix
gZ4DqbUTR6rOXj0Vif6hc6nN3Acu0oom5HeyxppZ8fHpuJQh84vmPfUByWewfxb2
1hZkAifvTX98zMVCvSGi0EmezYJBzLpU6GIfISgJ0lRZOPjTuBKsO3wxce4BO31J
HyjqHv+ptaLAWMwUj2en4S4uSx3mW6udEDD0eGd5jcZFLgleahNvBYzS15D6KaJr
BMk52RAB1xB67LeZAfAftX9zzk+QS4uxOo/9KeYTJp/Om2s5coq9dRTHVnNtXRSX
NRuTp2aDdSLhRC/rZ0WmWEAY4hSS/2eFdJ0zBbI6k9vGV5hfkJFma9nDI88/l0yz
8UbU1PK8IW1ZmOBAhq16oerSDCFknOawe8g6nHIHthPOWPliYAGHoooRAXNIod2s
g44pqAnud14Afqn4qDbmLdZG+H3pNQLS6wV4j2SaPf1j59gJR+UdOBk+xU0wkgDs
YX34wX1mAawWzTtP9/GxYaCJhmG2SRvMfsmZoH5FZ53UnYW30HPPEEZTW0LuMlvq
+VXA9kpA3hK9PTqexrbGjokJQDyI/ZNs0SGd4fuV0+oA0haHWdmtKPacFmGSdoYk
MbEjfz2OWBaTys07VACDxsEpSuwBEjy90ZL307vfvKODJqxzXp8zetwQhsplESIk
SdSn+ahaz/fn94rX+yeAxnNGdeEpk0S388NzpsfvQYErJiyMQW6Imw+c6yTVWJm9
7kEiXP61Z/dfM3PP14Adj+BDHPhKJfTHOpIQhNLvHye9UvpDogARE3cKfx+Ql/Eh
2m7du5hwZJIjxTfs65/xjwWDsUm8VQCiW1nYr3vvfzBfL5c0N28V5gpoVQSWUyms
XqEd4rb10Phsyy4UF817/2xt/Sn1yWoKPmT4ZodMBagsTX+T1wsQcQg8zvhce2fh
vIs+NdYjD8+fTcJg3zv5gbuCsg71ffGHW0FCbxykqp2URzq3xtKhcIctAAYSGct2
2aFLh/YPIz0Jtn88jT2qUVdzHcshL9SN85u/Y3LHqZaoPTKJmVVfyiyzhE74W3c9
JGrTbar4RPW4plMfnYIg5p5ODzmL0u5uB7OkfE+2CLQw4/Thc9k5jNQ1tr6MVycq
gdkVYjrd0CU3Q0NwgiuGTs4dxVvkP0DTrb10Zpc/4aLad+P64PuS4t9JogaTU40d
Iv7y+fL42xmBGgzmWkNSH3KlIln6DOAbWSknuP4sHu9qG7oSr0dMJdL8jZKTqCu6
IsRyP+BxFXzm33Fkr0ms5urpaYcNHVzkrpu6JxEyuRhPusrT0/tr6Wat52o+fuez
zALq6Iqm2PsU2+XvhIlCrOCsjMfC+L8Zf1Ov0H83ScOvQBwh7+h9dk/51WwUjhuD
lqd/HI3zaWmc1Q+JI16YXPSFMJBmW8FPl+wKqq4UMtkdXuEV3G+Go4m/XJgYGgX2
xHxHYaXeVvL2IBDOjOJvAWdMiBGErgcL7z50/TbuLDuX/ttBu5xynSu3twj+5o4n
xXz+zrTXvZUmTuJF4iOL5NVfBnR2IYUDbnOu2puFWeNLL427C3b7GUK7ogVnuDbT
l5e8y4wuw1hEcTtpqtom/0mTUwqlVsaQAc7iGsrJGj7P2/gj8gkJ/4WKNP2CssXW
/Oq+YONY1Cu8vm5VygI6g4LWVZTlhUNpcChvqo6isjz8jRIYLRuGzOEHnUuQ0JhQ
a0yMtuBOS70WMbdm96YLziyel7IgQ7p3I9To8WqS4Owc0bmx4OAijXl+3q954E6I
Oo8nyUcVuFotev0HUYUyT0dTS82bHdCmv4l9HM/pQZzlpL74X81hjA7//uL+CcQ8
6CaaV5TiZinfI/OMYP9dp6oqRU3T1EzXzl8t6mJaOwxiTa0aLdF/jZP7bgaGXwLC
2LL3YoeGQDE1DojWc7WEcAszLyIGOm+BIrjdjIhMHRX1IaEIN7dfca6TrDeOtOFy
YHYsrltaysgkz+pkZ3k5VulWZIbfLPZSXvxnDCY4kEfcABCHZjuls2UWdmsxvMSi
XF4XTtc9EdzP7+0Sm8Y3MbY4lkCHFv/Sa2rMkOElCBtXCSq0KQiNxAzkeAxlTms/
bEGc74itlS0AX8/VmWkL3mfw56zUfNNz5LzOm/HqrsdNEHCYWqIwAavYEBDOpVks
UujzWoClpSonFcgTKqKkw+ep+YHfH2+myXsWYDAuJ60wIrIBxSJyCEu8EpgDbbWn
GCi9UHnH3/Kecg74LWtRaLbw0W8oDIiFKQf/EEEG+scBVAn07bc8Q5o/hGdlVvxT
m3Ar3W+96jJ4etNm4urwe54yi9YUcHFa+BJJLPT5YoAvipgs5Ny04Te8TJB9xvRz
oqMjxxu0oc0XSt6odkQ0/0C8xOkM6oAz3EMZMncGQHNYwEcZDq9padm02z2/tf88
K8f8DPvJDN9lNT2wzRxtngFoQp40qLQtsdiCjyrcg09WvXDBZC4Nx4BZ5VaFN5o3
rzMg7aQMF4KU2iPuZsgKBPyEoOKdn/eSZAIPWS6dEEbj4MT5kNeQL0jOkGDR6nKo
2fdPcpBURSn2N8pr7W6bCdAB9ScFoymO9ug2HrzR1/RNhHv89A+RhxIZv9py6/Nt
wfdy0FJWbDCPyzXP8Had27AmiAsDDag3BWr98Vi/2duCsxCMSuhSZW+LHKkFlYdc
FCe2KVm4i1fP87qgY1Gr/IKqib1GFtQSmYmMXE9T5dm0rm9R/XNoZkHV23t4ptnM
66Jfp4YsboV++nb0QNmuLIjAvxTgletYoJxu5NzFkrkW/zsH/ccAuiOHTuFO7j/Z
+lNSWk/byJ+9JTxV6kenkhdxp6OxzjMoua24gVa2ZLqBqPuNOh9JyaIDDARZga7l
h6RtlH+7OfseR9vjZibfVRwuGlez03XYeifX4wfeWyVNsk4pHZ35qj463jaE6bmT
5wjGsTKzP85/rEIiMUWPbIS4QuQnFLA9bYrg/zj6udP4c8FH39UJ/JnmnWgyfNX9
/BCCE3VpYIp9c+kkR0DtfcyX4/K5ZHjgFDdcp8ISzDzz2UBmWg/5h+91E7ngPKY8
Xcu7YDqGcPfwWIPdyQHkmi1kMNrSmD1uR7xDpbmPk9gzPvzNcAkuXS3bFBupD2cJ
+DM+So1dXZ5LnLZw8QSBbfiZtMURN5TXdGTiA36PTYKJeK0kWQlLv3KEqaFKFSE7
zC1LHCYDa1npSu1SWFyjB+1LeK7E3+vJLDMHjDOoaNKiUx8FltfRmV/jItYLZjY1
AMQDtEa+RH9YeYjXLYabXp/qdRrIjdVUEeTX8mhroKAPxA0JKwHOXSfetk1m8fTT
pwNmY7zHZ7cUvY/+BXjQF4Rrn//S2nV2yfleWernNhrHlEr9VRYWcf4qvRelF7V2
RVX74o5lu4o8I8QYyfwNFeotkNvG09/vMmKgQocCcMEyXuCRATnRwdTqAUaIOf4u
U9tQRv7mE/R1WCqr1P9vs6rThAX6VdjzvI8xnWf7DglZCjsPJTcA0kEdjEKv0gB8
m+Z2wHV/vv7rIVggSKenGS4e88L/bcoU9pkHc7K/0YuO9PcdYjY65hhu1bVXvFqV
cMdpdvD35SK7QorH0T3YvWrnG818CyRx/AljFrzRPrdi6xFAWwLQUzZ0cXyqT3bp
frFOf4y7+cSQjcfNOdW0kif/+uIdvKG2dtnFWvFHV2+25Xle2IdjRXdG23/AgVuk
jgsogMFkGBkgDTpSoocK+aBqBir4h1GNX2Gsg1ZjXY5YrPHTwsZf4wPuWEZO1OyI
5SBxiGxg6jJCqu+BHk+56CK86Une2pNy2g6QX/dEa1343sKIsqqMheDKuUyJPBZu
HvNwaEQ30gNtuNQPy/e4azpuOvs5Uwj1cKBqCKPbP8NK3fKO8M6qiKHLjSbKjaQz
4G8xDwB3aSr7fg3My9hQcQUY2aSqVBTWTfcIZf6pMIKzqPRU4JGK/hg0AFERd6b6
HU92IOzc4b2RY6dbZZLqQR7rarKwMyzxRDIsKr38Sl8qb4IWhqq49nTEJBYA10vM
ML4Tb8h80sMdMqFFNDsRfgXS13jnwjiI0y1rpCA3ueVsY/9S/Nd+ydm+8+wUkHT0
LUkV/7Tryaau/JgZJlqdKelOV0KUn31mu4s6bPONTqwo5QSRLlK4bO0dQxpa3rNT
TXBwboorsRKH8ICv65cGYiZ//3uoClO+YvMMiKDmy+kBw56BAqmCpQb3GI/HZT1I
eUpFy+guKIdEybTImMnTFEeyZsz2vGB2Z0Xw93zInxbLY4Ncmutqg4TbBihEDtcZ
H2AoZY8O4cB1LaExORe2zOSIOCJCh15bO2qvwS9bpXKLrnIqpaGrTjaokv5TX4Qg
EvquZR2ij44oNOtl6FVm1D/7g+uNzVwb66B0HBI9Xz+1GqgnKIWSFmKjV89OXWlz
PVPumvSSOIhUZ10m21Xz0CeNxfBwD57jhINRvPmMEuyLSiI+BbENOtpYGAi3LK3/
rxCoa43T0HY/Zt6CE+1n8zdrFvYbgj461W2XaFSGQUuS70mbbaTS+6PDMeiM6NEv
2lwc+u2UjTEkYwPMiDfd3/J3UiBHVNRskUCYDYH5atPVOLKIzYP9+vDreqmPeF43
AwkVUBmPStPZEFxG+xyM6f9H36Y5I+KjTlyWiFQixuIFiavaTKgAH7o1im90apvv
hy/EziqgxiR6iva6kLAOPAp8Tcr2yNhFhtHxwPk7kuopQ+UKwadsH+DXNy6tD9Ky
8SyVcg1PgpR2wcGkoQVHkf2AUX4xd+3I3H2HJdjSHsMB0MN7JUt6ih7iz4m2VMYt
PQ3nSiIRFwrAqDYZzGIq1qKHle4LfNJS9sSed+j4V3J8tRz2zoLvuiu/CjoBuhYZ
ry1WGiV+rY7AWXfkJKvvJLRsrffSZdwpUjKfCV4P1OjBqvvicjqZ7bL+tCnUtxQn
LI9PJM8vUajWZifCEyiwFRe2hwdpGquzIL9rIOYMlK+wh5VbCwppEjDvemZVWXyf
0KtdhPA0bpCmKgRSm7tsBwoaQH8fuvN2atjX17dd47So+jQWrGRpN3V1snCbFgLa
zAGkiQ4wODHlQvDIVU701DnwhjdUPt14IYnsCYOPsfRxg4kfi6nIw9NyxWqlB7mQ
K93/duFGBMLe+TkjgsYI0hVkHpiieWW94aE35Exi3E1kvZH3SkayNqflaxrz8AXx
p6t6bpUZju58XbpskAUmwTV2g4407oLLKqgH6BEwcjnAZdQ5hkC8ruNZRntaP+S/
CVbbXpIUyTZiQvfrUuwL1ZgbMBs9dhoL4ynJSSok4ELPNphNavqVFA4KxfZuTp7l
0O70A+Zcgoi8X5+ooA7bvfIM+vgiLmi7/kMAokyRVPacbeRteg0AGLp+FqGraxZJ
jXyKqBQiF7+TVjpb4ByMyd/aLW0XDmWVzuLR9n4Le84Oc7y5wJ+XKBD3qoaw004E
0jdUS6Of8Wm+KYQ7RVbuwuwXlDwygRbLb60RmmZ3m8CgVJjizEPy8x9jH855Tb3y
RtVvt9yRqI5sQocpD+O9g8w5Tg718RQNCDRokXwYVLu7tOL2d8jDLgLJafpj4r3E
F/ALD3DOKBLZ8T6B2j8uo3R45DlhUseEI1kAxJBQdpW03/a0Zd7Wa6bPcYvUiFR3
gjgd19421DF2l3S76C5/O1h/5/hhMm7RNAIrMhPzu5F2D8Al0p+vHzyhc9CzM9IO
EzgCyOEuTz6vEfO2lUTg9CfkYaMv7tfDnc7Da38VCjVQYAyxJ7Rod5nuBIIJHB8W
+VmyGuLMgRdjsEbOaP/MMpAHbSuHgT7SzlcL+cF16qBfUhe5oGowFyWO2Il1+tJK
cy+U/bA3drhotmfO/oRk2USEeJVvMmMFp4DHaP5el4WOkulm/nzcklmu7FKhHJdN
Z3RvTu3TJMI2EeE/FKVuUFAw9f05NmxMHLfHL/yQ+QiNeZgAoHOf9VGxKC2OqAA5
DcTNsecRmpbC55Q9X+kAe8mkKiaL6KB663mbDpXKz/Gbfc/uSqEL8TgBN4SVHuxM
wC6R1KQvN28lT2iqQFFKBwxIiTNyx+v8KTBFtW1o4KL86zjTFk6NDPR2Lj0p8nUs
7bz5jsVHkkuAz6mY1Mp5t3j4Tzmcc5BjkDo/weoNek0PF4C4/O20u2LeAwJEiMbB
oMrsI06Ki5IjDwx8p0mBFucr4fCR3xttrFi7DpAtPQ8ttbCy9lMcqZV1MKyOxuwt
AziW5ZCo0WMY8v0Rf/Ci6DAZrHi29sa6WWxwH0iOIp70+kcgdbnaoKh3mt2He8cP
Ar/+Lc0GpFl26gPSWBj6lJu0aYrNm2G9qmurdElK239nNnCTWVe9M/MuMOz4pm82
mzyIp+0hYRoqJ/u1IPr6D1XSsA7nuyBQbXdw67CwvG0Jbv5O2IQPf2D9qZtRXTPO
4dSekALDVZ7a/w8vZTnqXb0k47NvsgPkH2GI8i0slZ5V58g72UCe5MTuwUDJLGZL
HU49MMe4P3elY3WFpUFB7CXfDvdQYwDURqTl4Nk9qdYQcj6b7Dqw60UGnMwX5TS7
ecwGq9B1LPqwOgzWXEpxKno6mXzxbaEAx3oFtw/Y8GxEuSmcI+AaJHZJ0m//weKX
meFa/YNdUxvtx7vMNxGsEdUAitMRqO4J2guU6QNBt+pIYNTVSW/t++wqkonEehw5
OMhDCMpE9jaoIQqHJnwHnOOElJrBnS8RWTKLY/9xkDhs+5gXjUrxUVg6scyYv6GU
0Po/EICHmOqu4sqrKaB2jEdNthg7d68NuVAORSGvyELvNpXDxUUwbsXB7O1Ni1C0
i0Lo0+YlUSVxS0TLrr0ubYDm+VLLJhSUuMSSyJNZxIGgy+jS+TsxMTvzEROrRoUU
Jd+iiamNTkTkxCIcFG+BrI/rCxVPCpUqK89vp1Ts1ufYQRl2VN5/cLwNoh5KJRLT
RDL2HAgmh/Xjsvwx4oJtWXZhtN+CZ7/bZzi7GIcYPb2MOoUzY6b4afwl9pMbJjTy
HF19uGwwncuvQaEllWex+JCag/qyp2ynFbNvcN4+e4MVwjPhws3WVKp/IcDJJdRp
IZitOo78zTxYscFjkxZVfGGl5+XQxhtF/V1dgiXevtXWwYKvtk4JVw6zA/12VCzz
cEuurVQaOWaQfTxdOFQartRpIMVn/iHu6JX2Z5RLPqKh4lHKF5kjLv9snNNN7u+B
qfCSC3/3bmIQfgSbuDkDF0XGwvuXSrashscucdaqRUELs8FFvC/GogykeOrluRJ+
DM3zvtqYTkZ7m21/f8CE8cKORmGRgiSm8BIAR7DTdyhLxsAJg9OrN/+/nL19OV9e
lz8sftBwzZj/0Skyg/jjqo6ipB57flHIxLMlyVJWGLLzfxSftOWOzVVfdhGBW6LV
GKQZTd9elIaq58Hj/TSbkj1aTaHo4C7JOTDqwz9Vf316ewUKyyT8L/TqKpUoydbZ
b2feEcLnFb1kInpTIvVVfNCNFqTK7bp2DIfL+8/P1RfCTXhIvGXF53w0Nrc01JyL
qMVj/rfelDCfP3tlXYwVVhtXhk32r7pgmP/3tMJEtB5zNbV3Tp9H/19B+q6lQPUS
UizIYrh7rrutKiwMvaNbx5XVKaC04TW6MUNN2rZWe24eheVFz74Gex/Nb8rGXTz0
7Rya+DLJNb2fTGqECpKZzd8TxVF/7l1dHFNs+IqDX5DSqythz2sEPqv6nxHKcx4u
vxcZZqhpLc5hnjlopMfGf8yYIOWDgByGCb6KZ5JI9xqdpRHZHuG4e7ICkRGDYCcS
E2CD6Dyn3gLn9fiDp+Lic433QkmwI7oEWSELq1Ys1Jx98jDsD/vmNUlobtb0+7wI
7AMMZ5vn1LRA5YnC3fsFtJ1XMl0z2tiv28+kzqvjTaTgB0/sy4OK03hiHoQ8vNaF
JizoXofgY38RpmTMK8sWSd0N0DpU10f/TWAL5lIppE3dmYztQq59Z6Vc5FzWkuxM
Kj90nziFQo56qLhCDwB0lxqRgJw9717A5pDFKpCE6XAuEeapM0Adgdgi7dqZyMjL
agCIUrnVEe21OrrH0tMrQzPhCxPFhUeNx4F7pOEfR6VimfX2zWF8legCs/5TUTxu
NYgmrP7axkmYaFrLim/Vju0GPYEbvgnBCC97Si5eIoRibR0u3+LnZtn3oqxLK++g
VNax5kSjNdVxr3y5EkYp5OEWGq6G8RmrNm6bBf80mHjIhE+uJU/4QdMIw7FXehvA
/1CtQnH8v+AnLsbpcDCqq0vz4EP5kta/BvP7R23Ikf7wwk+MwtxeWRlxn4A59iM6
R9uek1GaHdYXQsjbeXqAX+BdYpo3Ug4544eFvUUr11Zyl4WxR0hpxkEIUqBfbHJL
P+9qPEHkRKh/MNqTCifWqtHSeqVe21gvv5YmoKEi0rI0lDf8DZmDiWk6D2+Ofh/S
Yduqv/N+nJo7oi/Jdcs186jCXdub8sVb6imz+KLhdV5Qd9b+qYpWFnlVnO5833Rk
tSJCqzVEWLUf9+jJmDIo6zYozIrgfGv8lFg1+N87MlzcVqn794LtIOm2EtE3Ffs1
U1UA4tlT20/oOGlHQy/qBSREN6/OSEWnxwBKE6os3dzn0YE5HUVHXjCEq6PPgkbT
D827Jk5LuWRCeVE7rS0x0BQtuZGGU9dpEzFpeQQ5Hl+3VzUCAkVlUHPgB8TV+VvM
2otAQ+WCpzE5eiZthJWjPR4Uwed2gUztC3s1TRtGQI7XlHpQe11bXCm43L3GGJnA
31eZnxtJ0cBictyPXEr7XkHKD9yskkV6vSUlvqoem/GcdvB/hPHzPwNu0/90EH3n
9Z4TiI+1h0cZ9xigYZeQYWgTYykhYZINx8bZDnUu/OZ2x1/DZ/oTnfaLIjz3cApC
hQTZ8GRHbr995JsOZwqkTV0wlA13LtwBNojzlBcu1ZwgV1TzSwAgCbWg9bS5oLUp
Eq8adiCsQzAG4Ua2Krq/WYyDXDQfH46RDHPKxECoDjg68EJn9cq5G7vOmvoYWSQv
hrDUD17Ixl3x/fPbTGW6+ufqrHJ0juqy+EVJLZdyGxeQT1yd9pFUG1Mk792ZVbhS
0fmkQwiJNUPyeUqJTt+p2R6j+6LkYWVeSfyT9EbaLOlmlG98ZUscWzuAIS9hzrSb
0jAR1lOl+NlGBxSRFv7Xfo9111wEAy01qgChgNcYTk7jL+sT+Bvx8RMwDBCpxwhY
SR24pI/W0tUp6HNLs3fXAkzZXIcoH0adNVuWJZZt97XICyIBclqd67pJUSQGmgLU
EKu5MXjL86igZvo3nFI8lcKqOzN6x0kbBfRE34t5su6s0iN3Ugh4HhQqzSXM+Yxs
mTJHN8GpUVCXuZCqIKkKcj2gf3i6aos+i329/FccQc91hughcVaM/aiQD3nxYQEj
Fcy79CGvZWVcrFNF/U+frSYV4Ou27Sg6ddRmb1x9yROXn/DoLTiKXdywA/y7ox88
UJLNEjXcYDcy1HVxHjC4VgrDl+BwZSjElRLV9w7SU07BWljO4R8HckGPSHJP4v0/
wEagFamJFgL7wdPXWmboqmDDyPCRQI+I1ee6ZwpaVoB+/3+6NG/XwPA9xk8ECFgc
LE3bampjx8FlAY3QbbKWAD+QYPMKZk0h3/a9aUqs20fv5nRTrsSCE1+53FXeW349
Zt+kuCg8C9QSO8kenApgwZL1LgUhGYHJv4+taCcKL84wJs3jZskN/REDu1ZM4k0h
twKOZBWUGpSIVN1elU6osIcjKf9SmTwxkxXOrxfqmJR2nHYgR4XxqVu4E7NMTT/S
2+om9KwFzFlpusG6DWKGJh+6AYOUN/KV4akXYy854Cn2JjELNYRtjGv2ztqN8mul
paahVSh2vrk6xKjAdqVoJ2fPH7g7lqs8lTnPCzNTiNrQ8+WGcQ5c1dyHcItRXnDS
TsPmomTuQn5LGtXjHCt69UNFGtCw42ptf1UCnzvB9G/GRHYlom1eeyCBUonE/0qc
zPIPp56fOCadW1Ry6pmGMC2M1OxD9ApfrYCaXDlf2N17sCQ3eKdZ5SUK6dfkMXzZ
br1nI104t28uj7R2iFHSJW8TzTIRzdDXzl0T1kUiwl+0Bt5yviTY2hB+EVj0c/gb
jXZfN+91jn8XXzSPzM7oixXLLYgExj8EJMS+peQzQw73FPfnEQ/9gl9iKOm9TG1L
aUgQUQhAzZY7knmPrcnaxzLPX2bziycKRc6goFlP8e+kyqpweOLZ9mYPBxK5TBoA
B3dkubFa13qa/u3LYKbhLeuroLKccyIM1GbhyB9uSeruOcnCl9J4Zatv7SgyHssR
Dg5NSSCmqVJQwzsr7r9qd+9S/OXnOGhamhzmLjTcjSmiiMTUw93RGynn5imdGAS6
yw5vxNwJcxa7F2l0SDWxd9XAYFY2zr2sul+mlhjI2KONIBS0Ddkq2vpOOyE4k92V
fzpqhIFOxOfkIb9QGAQDbt96TeEcAk4lg4v2XeH6ngXO/N4ZD9gyc5ezM97q59/+
mcOhTDeVFh7ozv+uKDsQnK4nRu6uIa1Q+qFNfQUU3z3DIRY/ue+CW+sAleDosvQH
iheg5ArMd34TzICpJWWUp+buAiRib96Jsukdi9v9WDW5MQX4QW4yjWrUqqrOiPK6
rQ4WJdqkRzljXWPsIy9ve7fUlQu2Hfgnhx1vP3aHJgeotGQlg97XRCAyYW+ZCATi
opVLXR+x1iooNSn6aLGbuBtcCHQN1+bdBxN1MyS9psiqc91hIR6RNX6oX8mrzCwV
k61TnFN4HRC6TaP6wIdjzvjIevCHvUGUH80aBDxnlgl+nDv6QuLVGjqQCn6N0oTb
s/fILxi9DZ25fszJbUdHpM9/OPjkOUvCe9pzv4UDAwRisAHQeRCkr3kcPOOaRAh5
Ne7DfvCIMyUMfjKhvJEeCLnYqJdECZ0XnZpmoMmLI4Cum5NJ2Rslr4n5OPU+vnYk
J/ceLo12AjFMyeWXp46U6cy+0IDYQ52SwM3XCaAef+0uGnp39pen3qMi0WJwc/Bp
HYcdOCmElvFwiIGjvCKinpOht7chC9tbV9hLIA4gwupo2UZGaOwyQqiNVnK1sTl+
zzGaLVWLaPRJdfZsikvOQFtrigPQCxKqVVowuxu/v0MB5imSGIKokUFmRmbfTOev
+lfO20XQvHzxSk1JMBGNkggj1CXex4H/bYlmp2erEfinHgININCF5HNvuVipLb1r
wFEKwzTuDRD1Tamz5tFXV+eyzLeygnDJw+o2vJgGxwVlKYr+z4XFU6Feyyb3UoQK
nAs6Br0b4jVZ4ZfuUNDjLRcLRJYpwNEif+2PcTJ5Kd4bDptu0rzBKcrx+Ivch6W3
H50hMWnnBPonPQeIdEGsIjApP6UjF+yWk6k2CpI4EIbGEdBl7+eUnxTeq4cPMpH7
HhqBij7CXZhP8AqhWtlqdZI2LA0nswre/L5OVb2TrUh5ldO5oDM48DswgglPrCeF
qnGACy1k19fleYYgp2j9TlC/LrCjkit1OWKuwm23XSOajyhURhJ2C45BUZ6xBgJ9
rONEv9qZbyd1/KINStTJUy/NlNLnNOJ+kI62+jE6R/Hs3gxt73OmnpxbqT9rji3x
E+1MGlicBFeT7PSwOESJ08vjNwX2N2K0dtV656PHbeTEXFJhhbd6rMrwI5rYWq/J
J/85dNY+69trchGRSeGjtm6uA3ZlJMhQJ3oTuvB0v6+A3ZpcGxsYlkv9oRoRuHcF
Mleu1kCoy7BY7fhHcp7h5+RdRwgMPJHTin7eCbASmh0G84MpuTY2G9w2Tp7fIQ2L
3DnY0jey1/Irz8chNdm72saGLSW95BubbyTBwgbIR7gzVuU8kfP8NG5BqX8yPuxe
bFTfKoVhhaahIodGm5YYfUAgIgmG3KehdPZiS+DoJNVGCHstG8Nk+kCfctdz5fZr
5pVrOnya3qS6AblpGGollsL+he4jJe6IKGQStx3UJivUsp2YOGvQILt3v9QkQutk
Kju6hlTCARcaWxkNx72nEOXNel26cbblfSkjfIdJZdqDDNSjcJO8x6UYq2tWUUu8
O//uJKpI/kWMP/nD5yQgTYh3dRqROZL+/QcNkl5YuAo9XNXxVKUyGrW68XTFB2Bi
KZ/IUVJWS+niXKajfiR1InwKkCbQUEpZnvSZoF5yuf18BWKpmoKaYwRZcwL2lEUL
MmKy1ocS+0bgQA6tLw6b3zxyQChld5uyamQ/RnI5RzchEmrFKdhcuWxftWDCTLK4
+h3CXGV4wZIbRV9hWxhxdTmQ4AR+KxzYqzzK+ex2bPZiYKFL0ZVsSADrptFtUGxK
IV7JOghJWhoFpyF5738Iqsggh2+0XOjmRRLF7x2k8r1PXkKkN5TtSQ6rs1iqUaMi
gFQrVquB6S0EAbKcnl23ktO9N4qNUIN4E0o8v41QRUfAScGLmsszyiEX4lJDEtfa
tWFUuVQfbfk8nOipprYLZPSH3Y01Q78NMpVRs59dU1vGkkaEeak0agb9ySrBle+E
0KQIqYhSdQHN+86q11yRJkiVZUe+ptFK8v5eAWwpy2DGCawFdWzoWgtaG3BwUqqa
YlnhxVikd1nQF1NcGlUWFXZmyGd6fjlG/Gq7+yNl7z6ZdzS8k7+yJ9yDh8mSwGWI
DgTzdwa8jeBEaYX7N+5h6uyjNt4EH4hqRbCVLkEKk3EXRei9Zc6MztdvLUqvErsv
r0kBMOE6Su/2fx004nKEnxe1r0dFD27xZO7uOlh9eXy8Hh2uFzblV3ltU8FGshfE
OhNA8uKfLO3IwIMac9C3XsrD4h398KCMhRTqIgI1kZTduB7Ppa45bZ8V65VwCFcO
bO9fPZK+L+xIRoQFE8abv7G5r/NKzRfEYyKOMZV+gZwfLy52xklo/2zuzU0n7sgn
E2uzOKmIDuw+uvaMR5LSmavDJcMme48nH4ym5D8mHE5E2DDDs5rLMOhAxDpyDTYm
4BBZdLNXYEhHezzwIbBZE2OKi68Et0+BTjmZCkXPtwU2xdqZZgOGr1rBmqaLDs/c
CNmluSooLPcDNSSOchYorTz8Co8/zmN9grFrumZ0PxcOKKBYZ1fl5+GB32t6HZUe
tbY5+xg8npkS4OIRBXf3SV1BLymqEAQOZ/Th+2yiRW0xAEAkrNH2Ys5rHA85jlIg
lPaY5BVE1+rd/aPYtf9k4BzqutIRDNAiCQDRJM3AXqKfhjTD6lNzqPzFww4tIK1g
rfN9VHfLbIKx6DFaflzK2apkQPPph28yR2JrLo5HVe0hIBy0Jd264ybs7xefzqyB
+GMz/HjKtTfSQUFcSlZoV0IuvIr8lJQiY/hvKNeb/dQSbd6UrkMQUFcCaUa5hliH
YolcCJhftG0XkEGzMqEWG/BSC24RStp90Nf4aseAGQqGYwPBvEBSI/cjczT3yG7U
JlTJE9MdvPsNaq7k5I3xW4X5jqIdkbeN1j87wesH5SLvsX1MtXlm9pBYv6UA6PCu
YKFJ1nFhHkhtfxNQBmSFnkYGSt/J/Cr19VSjyDhgOKqfwEz/u7vqCjdI5vLiStsr
TZXBkF91X6qu1cUvQAZqwoNeK8XYtGoiCELqLbxY2jOl54uwXCuzt5bbTRcPGcn4
usVg8qZ0pSaS0BDFkkesS1jZNB/UNB60+aIcwhEKyg79+7U8k1xWhVfNNCZO+DzB
uuPR5FVAzt8Bjb/cM12onq+wqWlP9D7jRfTsHqjeCTEKhGsoPtwMcRxVp2omyBMT
3nag/ECgFLS5RUrkwVfuqvEBqDF7yyDso0oCSknHGw3L90MoDC/sgDJLouOaaYPh
2oq2NMErMT5KzUBHQLC506EXSkBQuE2pXccEoSS8TWCbkFg1KoY5fL5SbtbsiG/2
S49ChMcy2zp4FIts5iLsnmOcB6b7KzXT2mKs5jMiDV/Ug205zhPBw3Qqbp2MwrHv
jfxp/MKRnAxCM20V5Eds84qcF2TFY1vFdekgC66Nxc8i0HtdzF1JFU5F6zP5pAsw
9TdqsIFerEKSLFjO7a4voHyuwl6TMqt3xaQN+Q/D+q7B8Tn8HquZrLndsWapN7b/
dsywPK3qsjcvzLpRtrNu8CF53QcE2/ciFTfy1BLWDSUewYLxT0m5xjUtztgBZUE4
eHgHC4sEqi5u6aMqKvbU9xDyZNUHwUaw7G30JTQ/FjHSR6ZnLGjPNeGxqsd494zC
MofPKcJo/ssPlr9MlPJ3bqZwTv3wpUhrjiU9PMVV2uoEBnC5st8VQNCsBG5WkQ26
tBHMjWDagst+5CStEcA04uNj9H4SapFp7J0tfKVkj1tPKmZDUMqjiaT504dZmCRq
Ztu605aGSAFHHBJkAAjoc0Y6gr0nUsS24DQ5MCtrbpTPtV4t6Qtf2/Fq5fca//bV
a4l10CROnQsglA5z+6HGrCkCTDGmIcqehb+l6RTN17qZOA59U43EAtUUfqyWMTkr
tWPtOZD3v4/msJ3V91XD2EVTfT+SUP9oErZLrwv4J8CJHDnAL9s1miTNSehRuEn1
C9yT764qMzBxATlgDg6xdWkQXikCqC20cg9dwZNn+piSr7+T671ibpLA/tD7rVi3
RoxEpkLed9ZuCXUpd4SR6vqf8r8w5z+xJBpiLRU32t//W+j9Y+umRGzRUlo7Y9la
jWax20X57WOebl+iFtGacNQt8qCkafmtfeNjyr+AqNlhQPgEOKIA5SRMmXQsE78J
hGFAeGTcf7abXqPomXr8llAvAmfERf7UuqkuBWPFvVcxxeQqc4rPkNw4lOXUoGhH
XNP7Jf7O85u6V66b8egUqIw0pYyO4EsPtUP99Oyhy81zkcnb3M/R6gyGkeYOhYYB
+3dkV0uS+wJVEU+9IQl4zsHKtDO6B/Xv6s41gjaRVvJVCM+IzEjYW/w1iJPfoU60
awnTu0i53ZGLyNGVy12EwXpdQQ/WP8DLMuvvPgRjxTwRnTHfpsZsCXWNNaZAxVaZ
zTUbe5E+QFfWTgDNB2nqkmJrIuv32VFn7Kt4SHMnRgmfVfUJzK0d1tjkR3wyudZy
fNn+lUebdK2QrkC2uDIyZu77hAAz/tn6U5WVzt3zdy1TfPpcrWB4zOIkMg8EZDB9
ZFbYfaYZhiPP1DxuyJH3qqx0s1U+OQn6ROPJyGjgPMlYjy4WY9moSmB9Sfd/TlXv
I5cxGGons70Ps3z9AlLJsvN1Fh97nX2RN2FF42iPusUIqnqd8/yfoJvcSCBot/2D
Ak6u7NNufDyltzytXVR8qz+ZCIj97M95XsBpnFvDN09bhhZ8PtEL5vLA9+SvVCqG
EBoxTCVVfjkdVzoYBZ+FVFpCgXb5+5jYRahuV/idV0widcHG54JS4KxpnsrWqsXl
1vz2NTZztfB/RQ5uafWVAck9Ibj2KFnfbHXtxKUtVflpjX4LPhbmFDIYOTdNmt8n
wn4EqgPatzcxEEjV+DfmISVZ6LHaAGtpYt038J7IcGIoq5LEQ72ljesXdoEAGs+d
pzHzrgBWo/sCy2qLG1j755VPzor1CzzjvonecvEIMIhxl80LGIzno/XB9gxSDcKF
jISzBQeoeQGGbYYELIenqeCJvm4eN85wkV1RHI4IAgYzTVkOBsWonMgKvNMFsU1Y
4O027Yb4jFtCNE4qcJDYaiXu5UjbZE2S6cqncEODPWwNtbh9YK9AgVf4HNQzdDju
yQpp6WA/RaWOpHdb7sPqF5YD2ZbAK8I4jbRfuutx5J09/pbMuK8i0X1xFlP4jmTq
dcOlpVYKyheISgsADOCqF4Ikb2GN7mGiJ0HvtLGbAzqX8T5nCa3r/2vj732pRX3S
VPZG8WTxfN7L7FLcQB4hqAHrNOrER0SXUwqUZdulTpu5LE/ARgiISP+jrpJuNyHO
wLLD3GedeHht5DMm7SEbUuT7XuBexkgGnNpbUEkAQwVp0pjs9i2hkhqUnUmRgkm0
zR+dIWD4SxHcKJR7dMXGJZe/dyqhmX2KjmS3sFqXf7yh4xibE6B0yKoAhPbWw9YW
MtPcC/N4FtNPOuS1bk2fi7sO9OwBZbUNTQTHfcSWsJMOV7/x79Lx/lEkvEYMTSi0
g5ha2fkXs9fieW1bVBOVWG+Qi9RmS57aFJ2dQmEtsvyy2sXucySndOgYLdUM5+Oo
CSI9A5q55xaea23Z66oXlFCeQNq36ofu/9k18kcX7S7ppbZM9HIeSj2fp/NPt9i7
Rg5xhoLN7Vq1uxjPwu2++24YPJD8xkFk9QR9w3rIfu/dqvVfJWkd92h1pKAGNV3V
irBNwtXo6WgJH4I1Ede6ryy/2RFcDfSgUaxAcsu0yygTcaheUect8qdrsXuj/ND+
fN8PHGAgRPpqQekAAcau7byzt7vf4hkCHkiM1LRlOZVmMMy5CUMfeFRnwZyWJ8eC
Ealt4eq9BGycrhs/WAaXuF+ECgkTN/pt1ht8kTGg+OKrT9g82ZKLaZJf+Bv3epwf
Q3QPmgFh5oJvyKo3zc3KXogUIkdVq3s9qtDKBnIWDGze1haZAM4Ynqj/I8BdAb8h
ahbVEaDuESe+IXB0dYwBOa6zN+pMjkzRtMK64Niuv6PsYHouWaL9GkakYFAoxJWi
w+MkNkjm8dzSGRaVsmqBnvBt7r37AJO+UPFscKK8HEec1zZKujEsrXiT046C5jSN
I8/SVND6y9OkQ7geeVdurZoLvxW5N6k+S8aJXNQO1ni0VVVl2GaTb7bnQbC7ALQs
lYxFn4hc4u7QzyfksMPGg7z/2vCY2Qj1e68swPKbbjEhbeJvONhb53BFOCeGQ7Ju
lZ/jFvcy5QwbdB5jxpP0jBwaHbQgct97ncP5GFLB+ujrM7VnzwLgeSsjFr+E+h7x
NQr2csGKI1/OmrJqWQWoAUExwyH5nHZm8VXw9ihMDA+fYCvr56h4IoMRlI7NzRnH
rr1rikrg69QvYuOdoQvfZD7TLzHUgFn56KTNsrvT/t+WJZDpFX30H/ZbN0W5Oh5m
ZFUX5kdbsj8XQ/L7IittMJVr8qhiBKoFxf0m8rLQjqTgWza99xAHgqT55k87+PqI
K2bQF0FpsqXnM6nLqtoORiNHKnLZUbQvDhy6OV8jLbja/G6+4IytLPhSGZOu1tal
XJvKU06HlDQjAI2fjvZM/JAbaAQ3mwWTqCqZGZJHX4vaUr5oXZfUnz9IwT4ZS9Gr
SELcZ209W88jaSZTWVDLR1RU+GpulLbRBMfoHx9poiOGCd9V+EZ3ByyvD685SiN2
r9hRKHTqkiW27CHRZP6wlvsFwJCa+PzuKwri6goXy6jaieMLs14Cu7DDi8NJnDzB
kS/1Y0M/z1PN4TRldmyscRrZvSgjJzCnoELpV6oM8yBMiAsb9Kh6gohCe5wt+IJ8
S4b1TidIyUWGlRtmAnGEO12nU1117KApfmSCB4akEkmXZTYUhQw2lY6DPgCX332Y
YacZAgGB8oz0TIQMMPRSXGUCPhw+3YWJeZkoZ0jSKcTCWxKlX0KLQq1g7iBLOy05
AHZmzqnut0JngnKpzh7jz9v8WrkPxH3UROVRf/H7GT/krCYnDQS3tWqoLHfO84UN
W1BFCddYMTV79L47rDRzul4Zs8XUACcSVhuKN4aAIa54o3O4kXEQwPKMEtwZUCHD
uA/9+Lm1hgHbswcv5qmbJQOu36u2EesoIri6gySZBZ7G3TjeMYmIA1Z+xpZEN//a
hnmY9ZejAXxDKB467pt4l+s0qMCrmop4NUlD+K93axZL91D7/UV7ddtd0I0dHqGt
B56nuHwXyeDH31fQaWiD0ebS2vWfv8fQGkTvBjLFSVhpFTxP8Y+x9t4jcztpr3xM
1BtrEnSCNM+i5ZUfbsjp5xbifj6dPACPHcl/Mw5stdOlIaqy4/X+JgV4fUnXansH
LADOcVP2pUXSgf/tCDm88cbiP1ZyIFc6hIViqS6nsqhzEx7dwWERyUfiC/s50kKR
AkqO4/fOPXDgo/xwJUZ7pck77vmCnns8tIpKPBIlBuOkw9ws/kfcAB5GV11zlKGZ
TcgwNPWiwfPLI32+k5/68zu9gll44MbnaoeVFw+EKt9Xtu7lrTrWEl6Jn+yQE6h0
uz9YL9JQ9N0RyfaXvwd98cXradfX6hGyxz8bw1j02ZCGXwBIKQON7rog12rZ2e7j
c8iwuL9HMzMt0z56qp/ASB/p/C0zd6eJh74lK3FMwQpNFl4Rge9Qm96D7tJ3YPLu
xeS2fjHMvoo/xGcXSSc71SDqww2WXbe6CTg1C9qnMDMfKWQv6aTxYtf7gze6KBK9
LnCLuOhBncKFEUNp3a+X6vQIVD9jnGQaUTkLTkC9CyTzooV6u6w9vF8Gfh0/Zd3C
f2106fdPYlMeADJXVPnumehSH+ZX/f2nriKWIy0At72L+O4uUlodUuUqQIbwhdKW
DjHqzIP9LLc4En4+1hzlQqCfkXUpP8OVWDzgJAqSOBHZ0/8m4hvN4qMLlcNQpC8G
zLPZN7xslZE6Jk/XCaDnBJz+9oaFmSNTK8Ck453IxzdCLwfWTZXvxX79k8J3bprz
8qG5YsrqtHjXgGGuDYtJkdSBxbL7ENJCep11tPLPV2XVcgJyTUB7pjSy1C4uo2Q2
tV26OHFEEKdNTP6cV3nHCiMSvz2c4avTJyMB5uOzWMuk1PMcFIkaB4LyGnkuvwvj
1uLx8ROkxdpvkXNFJr/gl5TqivfylehYlsoYiiaf/Eyvbhp8WuBZlByqHotEO2Z9
ScL74GHpMouQOLrPvRd2SWLCudBxzkmL2UBp6OWmtcmkWoxMWAI9iBokpyUvMH4Y
ZwrvsIG1KZt683wbrS78+9CFE34Fjohw38/H3KEmAFplBKA+K8xPWwITcHJ+zxJn
YQFTZs6Pd/fbAfRejVLyImutiZ3WdQk+/3TooB0DrouNHRE1QPUuwqDOfa8g5Csp
Q2iFN9YUxrc9diez6H1Yu5n1D9aY847b78ovdx0LAjMlHAI7hHk3NhM4DEG2aW2y
yMX6alRmiq8gQSszBomJ0twiKbQ9HueD5W5488tXFBpP/jkpViqkjEPL7HgYAJIO
B6bBo1ohuKWlJ9lnHs1dGnInprJfCg55hTNpKJumjjksKjNr0ClQxZ5wuzAbj3lN
KWXyjTmRSBUb2JetmyBVVN9uAF2WLICDTDq3bzr5xa1mrLLF3qEmc6Joc3XLop4w
16eDsIz73507anijvzvvp+XNBBUbmWBJznGaAKYzR1ijhSj9B/Akt+7Pais0KMRE
H3bxcADSfKOTzEQOc7Zx8j9XPguKpzXfO0mjZ4371hbEvRlHNCiDMTDngT6rxUcd
m9AsT4hJl6VsBPRylvEcEDY4P0q46l5H2u6RLvDrLwmMfKyCBQnhMa5hSk+Z1RJI
mi9Atu68DboUSSVNVGs/UEYCgFgKu/OGA693sU9DAfrg9es+/MYVQGeNzMYyOKmk
rn3X27cFmr3Ej7k4NuuySxPrraR8RSKWOB6Zc4DSg1cyJ+jF05N+AdC0dZJZiW3a
6/Stwd7/L1SL4BAK1TiqxG1Apyp8LXDA//nYZzND4DYIjzonaMPno9S2ITbsGlqZ
Yhn4bCbrJyTEZR3y1Tz4OO0OKYnuCJarRE+kRukXPdz+mqySER5JmPoy8H8HOhb5
UbrSKIfnGiutxFQql4HePWi5UZmqKRWJ10Tm6aa8QCVkCe4AEn9yHEINOBXmqGPI
1ffVLQKpHUiOhU1RIiC/SfgD1RJCBEbcKqFNPel+0w5qCefmff3iA6wd1JHNfnOb
qQJWghzOazx3mRU75mBzQOAoJK7WjvbU0friEgsVvlmV5v/fvCuhLFHmKK6+dqAC
wz+BqaMpOUZgb2gkJaUfwx7voO/kQWF8xq59vak8Z2YISDxHiJ2a2co3hz9Q/ZZO
8JGcQ/j1etdW97ODvj4igdHfNfu6QDPmSijWyZZ6gd2Mc4RDbS4cALIAxdFjEAyZ
/hlidvjqqLQpkthLLvgQ6JAzA9G9t08Er7irJAY5Hp2pWp6cADvLrUWDWZyIbk8s
IUvoMPrcH9i0sU21TN5dY3lfKiM2+9zsWBXN3pA9C6hsIUkwL0UD149zCBCER6Jq
JiZY5/yDScvxXLN3zH+4+KPmdBzLCGktoTP7lPs3s4+iGBJ0rszQUWIJLKwiyWgk
e7E/kJbAYBZeBS+cTy8WB8ak852j7a7XjGXvCVEOti4lNs4nLHQXOUeEBbm33zET
1QuW1roIoeS2YTA58LcMjaL1usNsCzutaBJuI/GApkcWIBmX9o+zS9M7KGXK6nlX
c3MYUC9jJwL2FTBBBvUdXuMB1WEwLZ4YXP+mn93CGX/L7pWIGZElUrU4jYNKepAf
nK4eq8Rkz3Ij7Jl3LO0j6WDOUoUnBTZa1T4ZtsEqL5J/IJ1gAfBh0fmEeyoBN8H0
BZmdFkKk5nGYQps7B+l4gXVKSNKLt3Pct3dAMV800aH581SDj2ESIsV8yFacPfDM
fXyLBMhlMg6w/X+7ryn5i73icWiT6cqF3U9vhRmVttsd5xrfQynLIrBH/Mo/XA4w
AwC+G28mZhY3e7QWSHiFaqyUqOghOunrIPAKZUVQ2pPTJxlhKqRsk57vd9gqNSIW
aZ8AGWXHMKj/+fpfxzUVvztt6aQmz/gts8NA9EUBwPsIfvCVyImgoFmV6oTeod8J
yLXZOWN4SFKlyT1vFLYLE14XWxnRpp25dm16IoSgzISz7zPIGphtfhB744Mfs0BU
yHZ3d8jdxwlWk3scvIh/zi4OQnPzlS+uGS3RweTXKVF4DpvncPfLsh0wOk0vUZt0
uM22a3evefTuGg/eaix87YiuUmqzyMzalrqggtwWtOomBH0O9n8BpUmTaWFl6lxj
7AmP8CxL7rAMLdGs0S0YXf6n6AS4x+rDgMuwk18okt13QLddahFJblV6XfEeMCiW
zggc0g5w/NWfgmb/chUyQBYR/mFdFw1+Plah4LqBV57JgEY1ikwgP+k+1St9Dbk1
7PDbaSNvWoMN4zCA4c0heKRsLSHW/VaQwbswqQh7ou1V5yvjdmOxgIooXB194mBc
TpO8BsPCnujzGyeELsJ/cdhfdL6ofQ7UmXPVK8d2IZ6NmWIcVH86BCbvnAzXBYw+
/3BlZ0y2I97vHuZsGl7/FAdrbh/bEsMFGxheav+2b9y908U2I3Gp8hu7hOrpHPOw
mcmngZMIcdWSs4GZQnz/Nh81F90ShgNzCPT7sgNdd9TNbVsMC1q3MqVYxVbXlc+K
MMzMvHHByDxSt77F0xh6VIUxIzYz7ogNFFYvo0QmI2EmBoiFxiLP/3j0CEUr/dkC
VDCRDvEijfQMhYCkzJVf3a+b1lWBb9/xyWw8GCMg1R9PBeOMWkSfn6u2XMNQ/I+/
D+sVc9f9kRVbzRgLkAE187Z9gpKxChJU4g/oS91WMzz2PdMUpCqFoKEGjSc0Rvfx
1sNt+rRHMrJTMqzIHlbDwXJCuthD5CyOilh+JcTPn7H5LGfHfVBFT3RshGlC+xm6
E9MmYC5Hhwudug62gZa8b++c7bh0w9VwVVDnxgE83cTdg+nad8ylF52g3CsBQRug
/brScIq1eGZWQc0n7TPoYybCCtG35E4nogaE6SrenOP+mWab3BlOU9rxZnrLlhg+
gPV2o014xGNw2HsDSFe3fQItPxt8ePqSeBwU8v9IzI0mOxlosqhQUe0eTgg7YXO9
i6YQT1UAEHn3qPO/uADBoDFqq+XNe2Jl5AYWZn5QEsPwvMWJGN921q+WNFKA2QtY
OJlAAzdOAG+3WkOKZTLpYNHBAqkhckakVRWJCShSsgwD9COwFpMtvN9bino+Vke3
wTMZ5fVvCbL6Y+UG6RbkU/We3rAVw/EXJqArr5rU27wH+eKL8hZXB6MLR5wMJJFv
a5jfZjmp1hnPnldzLNbWusmHXUIbMPudydVwPsJv8aGsiSAdZb8LfePe1lw6TlnM
DdYkRFPZuK3KmqN0EsdbWa2KpJzSgw4KjxL81dIq+uLr+LRV0r8j4YCdCKU0nfIq
R6LNkAyrUrahYpRU4ojzrptROsWchZ3QhzEZdsjr67ibFjErjAYMXuKikqeohRoA
UF6ctmrqunHXaUf1r8cm8mqAnuFY4iLzIfd+MLrmKyqSIJlqdaGybJFfku/f7+1X
gUUrtTViHGp74gbhRavM78CByWhXBs9PNHRm9f8aLJKWO58IHFNmVk6uvVCDhTWg
9fWSwToXi+81QGMuGV2SSJk0Z8/Y7jLAXKeHztfIFOOQAbZGBUsZocWMFKLcIQEX
BMsi/aHkzkLQtKz8LJ5yFCrE/j6CSb5jbzNK5n/lw3DxiqkBdSlJM/wnCGg7nGZb
s59hPqfmknQyDKbcDXaEHDB8M6JSE6cpzb1iDa8q3VPGJibigPx60DyNiSDdvzEj
wETu8Wve53kWt5YrdjvBz3YBtRWF1ZfFZpbnkA4hTdkZlyaDuEhH0vBAGvd9jlla
kpug4IRvl9VOTavf+xKWmeuN7ppMObMnuNH+9j/je8cWRxDy+um9eBruZ9fE0wK/
yRKPLPa3XUWnp+Jk++FV9TL9VJmdHtNonhnUZu5RfQGMFIp70ahO7sd5Dmi/O3p0
wXjDmMaFEdcjGnujvT+kpPDEct7IgUG9KOvlrx65gKu0tJATFFmfm3KjQu8dTNAs
eMUbajuOzK9TRM2smT5W2EpUNl6bLALBukQgX2eVzFquwl5anQrjVEA5LpFECyTy
vSifM9ZIyEjOGOYeIKJhRWywgGJHcw8bcNXsYGPEJ2qYBEG98GEQ2c1SAUsnMljr
IXeSC/2HZlyVUIqN7OnKqk7EOXYjHCSCJBQCh3dUL1iSPgE6hhwp9pv8ilYbWA8K
YKJnyF4vMJy1zlXHWrF0s/cJ+4jiKRduixzO+/VFaJLJKkH8jJ1CwrAMc0KdWT3w
gepMbNcJ6Wd02hPAkL7h1L3rOV7uTFl2H3ARQrVO24UwzggZfLOGBfFpNuOk6RFK
KK2M2SLJqiZSaHvHMup8A5ypybfdj8EDzgS1lanp4TS9gGjB+BZBHZfJgkbxr0mQ
4XS5J6/lJDRFEJNZwvX8NIbqFeKPcil2dRPU3eBom6oYwZaJ7C6m1HY+W+ZHfe1v
1pJkpRg0RvgLniLDAsVxiJl7D/0uAsAg/hfC479Q9mMJ2dZePJmHYZph01295ZNF
SdbxEZgL34JhZsMs3wHPIFEs8o0fdKvHCoERa9n/SQ55f0J7cHTooFVWfC3DjRmL
mJBPLNHjM3Q1CuOTq9EjFTZKL4f+GEtPcBvWgkOcvaX4RxGREOg59kG3wclPd2dd
E6go/xMOnc1qcWh/EU4gNFJ8gZ1tiaLqxp2WSxpx0njPQcCeAzjIx5yNuq02ZYaQ
9k3p+krrlbeUDcHgKWAsv+oNyWktsg8vWFq5exwcNEaNxr6hY7CVt1OhX8sqILcK
rp2k01JsyHYhP5Clzh0dY9MnvXQ1K7N1UQ5Xa/HOVUzdzUfJUff4C8X/s/t0pDwR
2cHo+CU1gs7usw1I2ZHy9g0HgPUPRsXPLX3ELj3ylPbflWWdV8l0Ws7vCcBDgU/T
9rgjDwXn/yC1LE9VLJIsDHfuDOedbWvq8ALc7MiLGYNNibiM/cvEJB6FLKiJlFzj
HSrWE+PS2GeMcr2tf0Ni0d0SO37OVEdnRgPgRfCQkkAKSiBpHskjDqHjqxuIT75U
I5wi4S5XHOpGJWL2LlcdRtq0+y14fxWJhMYVyfadnaAUSuU38YomsaCck+Le0NPm
1gW02W7jmZKAoTm/zq+egfYZEHtFszhOO+/geDexuEW1HGdEgXEebjoV0C/0qtcP
zJ2flayunb7PqJ7SZiGUaCoVxwY8KwFBysx/ryggP+7p+xYNlXLSGPPYMG9010Ef
kuQlf2bVDyaElWbXdjFVQR5OLs9bizXhN+4hwIo5DkCwKMPD1AYaTxt6x10PS6aL
JtGk0+xztDsuDERPhwELZCZGIsdh6iyVOsERX9k4/XVtoksBeFv8OMSSw9F6M7la
wZ/sClAgaxWnZlKPWIcVseOiNZQjkwnhqnJnk3+wjM/ykW2/Zi8/13+NMjtwQB51
AW9xPiKOMqzKG4pGjxKwXjQ7r0YyBCJNHu5AhSyxZD2ghIOXkyoEyM+Pd7Qy2oZM
bzGFtMZ8LXVWBcIMznO0qYHjo+PD1xWMGV2WcZKw4nyj8KgyUHT8ipMgGKiVLjRf
BUHIO6JmjheMTfAGJ8BMnGPB1ApaMcafywOw6BU0uALb3Zc/W1eyVVx1r7N/WAew
KLoHgEBy9dIqNei/261Gm7kgtZVJP2wCxk/a5Ul/qJtm6f2AWzWthcTIFfoLKrHa
i5Msbrx0pfkPaUN16/BkIEOfpoPuks7vwQC5kJe7R6gvCOCF9xO1ncsZYkH0pBMU
KRXqWvtUvfG0FukvVyLnQKtmOptT3Xxyz+dC9a7cbGdSao97EXwpEcuwgOawwqR3
AKVbKcGfaMLtdjao3qgbHYiHXF3lRNJVWFa2OxM4kkC0c+KD/g0tsYQAd26Zs3A4
oGVXEVwdtUO8PmtIaLH5QmC1+uyVUeF3VxbfeX9nmimgIoQiOrYQsmA8yqBylQvw
g1oTiJWzMtqjkcVs9UH8YNC9478r7RjW3UdrD5lr1a+fbi5PWEEUtMtap/PeOGGi
AMVPCKn6VtOgZ1n8NOrGBRKS4zZ+cXopnU9wfqHJ7essbm1H+SCB73gPCcyOU+F5
vqIAMVIXG+WVhMCBaifKtzoIMeIeOQSwyKFoCfT5gAwLfeHp0ntLVTUm/gqwHOkJ
vcAK03hBu9VQUcbdI52tN5ooDloqdbF8rYyzpX1sw9s0fySLPyO/v6bq1Kb/SW0I
ixNeMYgCegvk44lKGoSqaGFcGZk/7Jp3tGlkSp8ezZNme3/0qxEjVZinXebkGjF1
fWRG+++hm44yqJG1+pp6t52/fuaHJCPig7WsZ5qgUK+3Mw9VnObxAruin3Qcy4Hx
OT7QDqba6YiQPymO+mirSitVrBxZBsGPfSNY7Pop4fhfwsxq+xMspxjEQRLFD1GM
gOfdW8XlY7iPlhYTuaxDReBOlTLgEnPNmNCF4XRTE9cGIHblUURT/9gUaezgQVa6
hV/P6vOmyCe8V/WewksbSBBpvC7ux9SkA3Kn5jG3WkXTFTgB+8EM3qkZKn6hYNZU
rjfY8+GJeJlEpP4IUAYvLZzHq3wMK8RjOzKXESMPc9MiURsyLxlIKsfsvhnaljkd
I9T6+Cv66W23gPrw7zSQ+HbyXRJEmOyvvDdiGYYEhYwVLDokSVPliTGf2cBUoeIg
SCeQeatRuRLVl0Dofx7wh3Y1bKaP8ErggzbiV13sAExKRKwHtd4zKGcd2P1gWaVi
f9+anOt9PD+8xB5IKlqTUib6Ta5RdjHcWp3nd+aSqqIKxHapZ4helO0MyYNiJhQY
NeBM9JHQA4FGBhyf0esSzGMgMMrl9XMSs7EnyHvSjCF2F4c9V1EtE4aeniI/gU7r
DGnA8WzmIwwHiBM7JtcPZ3w0ZemfCpOEF5mkEL2ZkVdqw6rs/9I/UiqjIOCzmLHE
MG5/YGKGqRswUIozAB7NRUqMfy+yC8UBOzTS5dE2Ucd0C/6Y1FuMbjMGW2/Hd+UA
pGhJpsKzexr4CcbrHPcg/Jq17vQTAWy6sVTwN4Wn232Gbk+QwYU77U+8d6dZgr+6
4dYejhjPx9EXOL3yGR7PlbvErsIUEmtVsyBPIkOxsNDrIir6puPtXQsVMB4es4+r
f7UvjsB51/U1oHUcUuv5N6mJyVIdxCuR/ZtCfX9yYj7IbripR5j8QA/WEiAlqs83
ELLq+M/kgL1JVK/YzrRvNOTdUskob2EM3aFjqUE7zd5HtmdsOENC2semWNoI8L6/
cXa9CHC61Lq3FQ/c9cfs1S1/QNQF8AM4w33CpQHA6fb3qDKcvwcPj0+qoKoZ+7bE
SKEj9gV02inH91G/sTtS7HDt2b2t85Z7iJE022jTessJG0wGh5a/X0ZiyWqIncGN
WF5mg2eY/knUnjMoaIlEO7QYNTWCN8vpZL57IyTmvz3yY7J3PKkCT/4rHWVRwuUn
Siy2GVoRFptlXYNt/0dnunktMZgbwFXAusNQm3Yq/EA1DzViiuJgHnb61ktChhuz
OLICDJl2kmDxk4GuUvE9hlRHv2hEbgjbsnivbj3dRpMIKxIuDZvfnIdlfn74Qx0d
czsv5UEqvhGI+77+zASl2hcC71mDBdpFOvQWlR1NImc4TZJrYq0uibzKms8kam33
wFnNQSSngp3BqRXGzF3ROy00X6/D+fHovLZkSSUuEhYHLgffNGs4M1QY6Qn64IpE
K/RcLnkC9ZCr8dkhyNZZV/KR8El2E3b+lqGcw8uA8etg+5Gk4OY8R6a4JiNYjrqz
FrKEgAsmGL2hG7dUDFjagXSZ36081JNreGILFz67kDXy/YT5ZdfIpHE1q3EOuADb
JiqbDut9ocwlQYjekIVOd4YqyE3QL6n9H53VI3uPYlXRka3BMo/Jty1VrVFSTKT7
EmXymxyzl3RntsyJKuX9EhmRybcLRMaP6NEYm1oeqHYAD6Dgok3Ju2SRixHfsJeT
KArifTL7z6t6otNow/o3x7Y1CZFqJdBhfiMjrdOnWkqf4TiZMjaeFqlZHLnYnwJQ
o5TzkJ5ZYfMBIxRFAKZC6xbRzuO4MGUyRoZqVdjzMM0Pdumb3KfADA7v/G9VwFpx
Ur9H7mL2teBuw5812X5sC9WgzyGwS2qsfDORbNANeBtStgXfhYjTksAX1a+0TPnG
EEraGudB6J2I2kUqsXnsJhyUQrBBdBym5pSopyYUXzKHFowvQUUeWObjI/bUvtNe
UHds11yxSSWuLy4tUSRBJWLdfcRopDSDbt5PE0ie4SWyeVhU6HfvqjES6WNUD/Hs
G1rDKMgOZPpGs0ZDnHnlDO6qHR5zaI/4RyEQbZqqFlkZ/Q8A9idpobYYzwwGe3tL
XyMmaVu6aMYHzG3IUCHbleOuXXE9hFcdyfwpMuKcbspBzvHz5en1BhYqXKibiw7U
Tv+RkLgaE9FcRZtJ3hRl3YJOoLjB+goshk0hoz49b9UuSan6t+k48yaOTFTQXu6X
pwxZF1DUpohKCoFpcdYGiCf9Q1ZsNmSLglrwyZHSn579BJ62Q1JuJLksy3J//FJV
c0wj9F9hGoyOb6r0ybKb5QLvpmtUdfNjOGpUWBRESgFSz62XPL80YcnSgLNtVboQ
i+0sp0WyvouLjUpBY0t+LgfOs0QeaFU7M9p6K5DMVnHDVMOLQWbJkvcnQBruOOEF
8eXQUffn2ReRhjTypLsO3YrxmcZMWU2+j8VXtTVhpjEHXgK4FunNK1KDW3UDjNXL
8ApyNga7Sxze3Ay/QrPcIZoxQdH5H+Mhf/ub0aX+B+tG4Hquo6zMepPirRO5lXfF
r0Q6GiO6/d3mtete44AH6C8b4SuC2tIxr7QCzrbD6PntY2H3Mr+sRCBQlmGgacCG
4n31Bkre+EpJdIZsVWYr56iUULlyrHs2rKsDU/Lc8rxs5izEiWPnTwKJKCXsHXro
VkjL/vPBXhWEim2lYGIp2wCBmsCgJ1UkSCkEL+Mw5jXqu34SzMR25NzcRtP/oxRB
ePUTxyk9wJNsl95QrFP57UiJz+Gx/h7ouuIB3KyUIiU60Tlu3BmEYaOdji6PXKCU
JHxa+YutH1BToRMGWRvRyLmU6cZT87Hk/aqApm4so3GeHDqXl2PvDVhQL+Kt/Xt4
BByVXud17dgEIFG2W0yv1zRdBc/UWiC4RiZRoa8zAHHO2IkjGNDsOf0GKD4oOfQM
Cs2tGWQJwoTI0hyLAG0w2yL8s5ZjuLvzEStlK7c+P/tKbwMMSHTd3iewtb0xPZbD
lFywMg6oWWW5m7gxJ7bm9MagqT5/J6PUc2i5wxqFZvMEUPibLbUuiXCnFbnnuJ7c
z6AeDEFgzVT2lfAaSvnU2ZG4bW/bB4KFoJWViXANG5h8M/vt6RO64fy+JTu+99YC
b9Bbh+BaXp2P9LLk1ofLw/XRmVxznVnvPSs9dOecPfQW2FNPdTi1bWztqjS+8n5x
Qu94zXF6AqBRTtRu+gHvDUJoWKs0synLKJwnsau9AqskHiOutUFs/DGqXET7j9J2
TjtyyKQilcW7Gfgy2NuYxDIhsavpVKyZB12AsxtYbVWNEwqFX+o8z6n9lS1D8SGK
k2BoNEcKhm0DoIETNTpPvzUsA3gm/et0GEoBixsYcWd/qq+rZLDQSI4f8IwhENzl
NHWdzzAfb+2jfFEg9jieKCXH8WBnn1XbDdyRyTNpnHS5VspQu2EjM5e5fi+3F4Kh
nOSeclL52Wf52RMnam9Iwa6j6m4hD5XHk2WcJK1raEFSqd9omzBn/B9rTJAJB4HW
HeIeCVzBc5dsuGgeKuS0K/VuhWp3Qdx22ODELz2a0fLwgaAW/qtR3Zgjh5CNKEML
FM590lg8AmHGVnf7qQOTy01NxorZxcujGtQiXl74FOaijG8x37UVfGIMskq9aptU
j9IsdHOwtUwjBXsHt4K3+O1nZeArYYFQ3iX6U2bqYeTJpF8rTCE8OKlHWCtVY7eu
VxlsvgObT18rAO99rhfAmtS4fVFK6UmzCT3R5cR+lsKsc/FUnnuvDnSpSmrGy4Xy
EuEQt12tWwpB8NZSLef8dqM+f4DNKAdiQ+CR2abScIc/K9AHjdN2u+c1N22JNfn7
ecCgvlybMQuzq4pRZ+7CsKFEd449HdLY7zpGaPfCgiF8eI4cqzRZclp//gz7y77n
lXCVd07B698HaVWK7dgCU56U6LZcl7oWYdQK9LNIr0ZxgwvtRezKlh8QoHltcymy
EiwEvUsbb/tnkcPEOSjK5puGbynIvJFrxijzxrg8qZ0iyPmlkZXxXGCXQhB9AmYH
m+OeqZ6Bb5taSFGGdV6F8Xr3xh5kS+sJFuOJuvPhlPa/2xyixEOyNgJerE5neeDc
08jj+cn25qNSTAXzdOz8xxHGlDoUmLGE+ERXvw/vb0pmRcajdyRGHtJJRc3MfidO
HL7WjBhbc3UwXjFUwuFfDXtI/UGZ1IkfQMx+6sblCCoqsthSLKqP/gh8AY0NUWrm
RBSEKU5GLFZKVE4btxYqq2hl37JSM11/5t1js+vHHpUkmhqQRGdqJBCvjHfAfOeV
yAIogQfizwcx1Coi4F/YboX2HTDWkzmE8YjCUpD+9aTWfoaBI7LG5ffNCI1gsno2
dJy9STygH1V63o5ykP3xvUMPr5QACjW3f51S8dvio9hGzA6PMrLCyhtF2eBhUcLT
BJ4JO6yAqm6H4J4hFAsuiwUqZt41uphCuoS25m/FMbuQOwM4cJIFRXRku2NZ79cy
V/TXYMXv8mxLPG9wLtuDUCXRcv5KJchPzMMtyFljjz9+rr2YhGdBPrY1Tn3uv+oU
lh21FWpCyT/UgB/Cw+QTBlczcpIqO6eAm2Mww36Ua/n6Ud0BJFAThVn+goTWk5aw
SohpLjDyjO28yMlsq3CFnUFeJDc8hHuEtry0gQe0abF7i7sMaDYKqhmthUH2v3ho
seQ1dCZblVnd59JX97T68gy8UVp41xWijQV42MyEeezUCfm3vX6SOrb35hrS97zl
oqnrteLJ3g3HUGZmobecNMWtg/NAj0bBPYWi9dNjPKuSyqRWT1kz9sxb3h0C504F
7jqy+4E1M79MTvhYFMv2lskE92iQgq9O3n252ZkZ4kU1Q/vZvlz3LbkJ+B2iBa8V
NJGJjLvnMAQbxd4e/EQirJc8Gi1F06OhFd+ixNm/N1yG05ajlPz/gqhAv64U0hpP
7JgyFynp8ctF5ghI4qtY20qVQEEZYMSi6KNzHRNF5Vq9jg0HUHAHCXM7ZZGBXOms
fGJsw482AJycvoWWlM2bFwPxEhT2JwPueDigIHD+lZi74HeKHABzhflQygEmCyHv
lUJdVaVhzGqpd0qSopG3kfQ27VdIATULAEU4NRwjAl4KRa1D9skjDdKxpYclUbU5
m3A/G6DaE6dLB8yPvYXQ5TMo6lAPbh7P4bKjtoBr1bjr80lbKJpspAE7veb8CTes
YF0uTOL8aeJynjRCBw1SKHBj8UjzWuDHOx0bA4hWAcTO0y/aDv+iNpXvco6jfT/8
Pxy8zJBVLq7UuwnqvQOggRj7Lsq35JsKFTYIXy2Jt37T9yYkQeodA4OErA8AzofS
repGhXkp8ajLLhZ2SNVGU3txLW6ig5fKCyBEU+4Lz0IMWaakpbP4rNh3Ym5/9mAE
9trw48AzyhL/6idNqqqnLUTDiqx6DVV+5ru1x33aCJrXSdvP+T/1F8F9VCAiTXeL
uTaOvyjGXjTk2Ytv8uXl6QruCuMj8ggNaFAUaM1gAEc0Bqc1Nt8X0DdFOfpkpNiM
zQV851CYtpeNRMny3AcnJfGEfKKwC2sMxdeEIB0rcFo4uf2X2Lnl8k0bhk9abdDg
KxchE9+pEmHMRG8M2vsp0eaf4YZd7n7Crte1FOY2ZMRld+VPbogbDPSBAZcmZCGD
7zlKUKepXDh+Yov5jrVZq7G/e10StOtwjnz2DXJ9KBs+80v6jeZGB7+FZBMbU7mg
O+dijhSTXyBbQlIo1/iTsU4vFXjKtzIruix+3kiGK6YQTv1i+uE1sCbxYdqqsyzS
UCFgcQ+IXdvUh/8oCUibWE5huAkaObG+FWrZU1sVShmM2H37MgCvNoHJEYMlkFMK
IBUwE5/Pyum6B+jATeGL/4Z8LrO+uI3IVRVWBbG4EmXNnRAs5LNi9htw05HTszKw
mJjMlSjCGRziAmDvzqqqovc5tO49cRtrBpKKyX/nOUHFOSYFE0TbR94b7LJaOqQL
TzWPnW8LnmV62aKawZ4ayVLiQwRgLT7z4IC3nLYIHptT9YHEX35yv7FW6d7pj37f
cx+q9jwOfr3xXu/Bfcvp0u10G6LAqun/Yip9z6KgATxrXfFd7JWQNsdih46nxNOT
v2YlpZpHvc8BL+OFNsI8YIfxgkCKHVg5vvhGLUvW+mvVx48nFufmqtRvrwm1Frbi
eXX9/3zVXhwmWujmjuZ6Jz/BU5iSRsLgxuBAbzA8lpnQyIe79u71kX0zH73zawHo
jBDcv4V0tFSQpwf34qkgn9IoUjdJ1lpr8I0Jp929O+4SMh7q8IOVMeC86/tg+eLY
ghrfzuH5uTw/LrHdWk46ts8KC5asuP3VgcyPXgzAnUT0E00NW9jwnNP9TZQwDYO0
ecTtszkTaFHi+vA5WdxGEzxdkXt3tUiTxwg1ZYJFU+0X35cQDBvuJUUjwr9HbZ02
GCnrh8GyJxB1Q2OK/EXol5Nis/Tuu09w4ufvfhruJtsfVmDzqQvhE9kcI+uqwWaX
K+z/lub2C8Lb26X1bUfmMYHheCYl1PZBDLnaaf4+hYCDruteclGgpYm8H1nH3Xdk
h2kGlKp+MjcrUfrPxER3FrRijP/2yjVDAYULBN4GCJgSbyrpv3dVBoUFXUD2xtHS
6D/cycWH8m7ZKq6+kdvjhD5fEkfq8wgbUeRClNWvMVzhNXhjkrQYjEAy2ozOQx9h
75nRE40kZHtD5DM6CEfrCo5zUqYLPgUBFjlur+0SsWc7ztq3kDJRBGmGCUHX/K7f
tF5zuy9PQEsqQDRVoPNNYmzh2cW8p1OuVVu8vbSI9Eh5UHI7r50Il4kSC7S2SGhs
Jd0CCmph+7fJluSOw941zYQDR8KkZ617FPxiHUk5YYY+DRP8ApAb74UMyTvInEfc
2Z9CclZgLqSs80S3jT/OzVX7GnAiJOgYjzN6BebO+gCMXI+II7b2Y7TLev27oX0h
dgqgfgxS9m/bKcdJJVj3IHpykM9vl/fyBVIM/7+FYn100GYl//sdTIkKkWeIPB+s
lDycQTPFTt8OSRFQ+ZUmTk2HMpxLK4YaenyMvI5KF7zwKwtekZCICMZVw2VkFFLH
tjf7G2yGnjqCP9ALqXqwy3cH9rT5vgbMyuoJZMCbdZBQfJR6lZUuKN7U86WTUlvS
UCXAUjHTMyE7jKKjQyzYuKhBeLN1LjHcd6ucg4nF0wV7DZ/xutJSi4YWTCP2tDH1
YT1SXgEHv6y/V9RVdQTRgwnNKcsASQbNvXzO5x0wupdhXTe69lSvcmGkU/CWRRzI
SdyB4xBEtkcjgetR6paMW50zHiJB7A/amNznPUHThXMGPYu/AosOopo2YT5Lt1vL
ppIVx73U1MSqcUfMjie9yzC9c/gPmB0KlHc4+YlofNylKv5z6mfdRN1ao7ExwZjT
oBftXR06loXUZiByjIpESYmM3P520hjuycjcWRPVzPmJnF7+hPWRpFmuNZriAnJ8
UbOde7xIvJaBr0ZLBJYj7TS5TaA2Van9vPE+w9UxXLxd1s9uY9dQnd1XBjUp1lDz
HiGc83Ya5NUN9Ayaebq9lTO0NHJDS2JAz9OcUsZdShyARLHVCsNyShiPL0TM0Rmj
nLllJIdTt0M5gRMNDJFQKDfMdrvx0MmpQ/GlJ8eiUCExJHUcB9ogXz/31c6UlIOz
m225A1D+VtcBfFhxmYAHfywztBVaAm2vu455VaBCP1JDmHhsqdltzZ4hb8U2I6FP
dCuV6hPG3E9OLNKXKJH6NW2XHZE4dY9qGfz9V6gvZoVDLXEuy6z3S5L7cgBXYQYz
S10PrP652q7UCs+chyJymAh5dHACm1ksUQOw5xkRk4vvuXs731kWopf+xWMYrfwr
K3jzCKcd3PMGillC/6qVyYr/OxJVU+xLUhmYl+qteLkAsvGSldJ0Fe7skiehBFi6
LVChlLnChgZQNHx948nV3I+ZM4YO4NcLqxxq4YiiNgRMWG/nc1eDYk9+Wa2qqhDI
9Tk2kwhCw+lCvZ0wZzF0vJ4UQ8gy6Zb4ts5VQO51c8SGdpwkZfLBti2vFJ1zk3fJ
vMGQAICjjU4UZLQ018gaUT6Qx27AO6KcngrldQsEbPcqYgE+0rJ/Ag72izXDtmNx
yZQMTMTjBS24Y72e51S1UehP5GqVDIFb3oH3bfXf+zuFJKY5oGxuwODOQ3yGnVvn
9cQMZfcjLN4/elk/G8l+cfrQCtOsGPvLu+sd+zE6nDslL34yUbLYYCaLUyZHfWGj
PFR+RC9wwF4Y6HHH+OaitVgn9t22ym+HK7+VXqdcbMcxikLGwxul6j4PEligi9Ye
M1jAfQqHQfIW0mTTFr9w/XRRmYK1F/i85iJj+YqbZKNOHYV23qjBJRNGTMsY7XNB
A67nKxQSgfwoi7/z4arX9Ln/AFBj0afs1vqup5Zpwu4ItsXhzhIDzhjwnLSUlAah
f6dU35xJTO5uMGbpW1dJb1QfUkCC/+jQo+KS3G3JI2UWOo7v1L/CI6H5afMUg0vJ
Q/07Kwj3pH9AuDSjmvwrqqbcDeiGEcrRhkVg3gooPjn8NJDf+lr0xlbJ8fIa/XB/
41GSJJDEWh+fgXXDXwE2qS9/cc5zbiDIjMaTNdhP/CnaKwDnOM6MPbkgn4R/myBB
3GD9+EW9B+rfkuNZibirckEC+NWbN2km7MmbKbU3lLMpNh1y8GL/cFTRkgPEc8SO
aE11TS60iUGy4ZGJvoUFuuchuo0PANZekUIeTQU4Mkg3xvGpLRC4YUt243t/5NK1
iRBN8bzeJNc1ekUoxsNorXInHX+ul7YHd15ucDiv0CBu8e3lGdO+D2GdWHx5pvl/
dfvEpaD4q/U7in/+6lPi/4kIUIkhOSfEwJ7RglUKIgXexW46967HUH33N2La79wN
ysHRu5nn+r1XcmYaHNAfLpYyDVPB93RyfQ1dkMLgMjzP4bSjkofNOZIcG+Dvyi4s
fBd5Bdc09cgf5hqD7cj0ehgCvPY/TMCrb86fNBJWoxUUs5PWSFrzqr8kNsrX2RJz
B5rY5NAQuku3ni4dAPUzJ60XMgvdniZHXlGYatRs1HEVcYthJmKG95wRay9h8Un0
WB8Wg8DDDfCoxr7J5Sv5gqYosIFs00fzHL7FE8b3dKn3GgQxOUIww6F7bLexi8NS
5ksI6XPx4o5E2PA52vVFqx3yxaY93qvVm8o/bH1F/EO+MW/uCJrhFcSQPVs1a/Jn
FtMabkU/BInb6feOx0uvnfeW6hnxR+6sZG7dab8QVlJs7jHjeXuJ9sDs7A+oSpA/
lRMIMHEruoVyAKh1YDNmp5vtXWi7LkbZp6gVC1vNQLsVpCRSv/VraOeS8TZ3FWf/
anA1ikm3bn+MtmxaEBYHuO2TEqgh/tWhxGnxn6m/To+OY7HBwhdhY9+yEQgyEONP
+ez+na4roYt3eO+F3nlWkZQJ+UhFBHRy4nWcdQb+XwjtrlK2oYP4vceaXulNlGB8
QripoO+jpXXGz6+NvIOVi52/N3arprG9zQxQ9AOHs3+Vb0eyV5OiUg/0AkBQPtiu
2hO8pC0HhB49RVlgkEqgX4nGaq0K178azaKehsm3Oag0GBTp4BmtVt8nZq4oFfuE
M0WRZh6R495Wdp8UXihU3hdzbuupEoUi67Es2fr5rR52P6re2wJUBxaT9m8Vs4sb
vlTBagEweB+oLEMyOYIyyDaVyboJ6ktlwhxByKtIqZVdZbYdn4VjRqtzqEC6DOPl
BEA1/wLniUMB7oXDh+Hm7qFYr4Rm4DjVdwZ8LsZmSMMBEVzr5ETpCIc47Plh0hz2
VX6yzeS6uGbUzhMBZT5UOW5CxXoPBvhNJcD9+KaOthpYVQXVmLVUDTlJdxVFS/Sj
kicymTRT2GAJzZq7YrBb7rr22+p3pLemaw7erqJAw9nECb2l2UY2lRuCll5GAzE3
bX6Xzh3yX9cXIC5m+AG0M7ZIoEDGikfmSXO4C2QHI9hYOiHN4UbfoOnKEvKH3FfH
AbaxgYwaY0H+2c89MskLTnsd9uIbfvtwXuSm4D6yAIOiaOtA2YadT1ddRl5p9B4v
alpF4jF4NaknTdemqMSRLckBXrkw7KfwJ1ymZ3mc7t3iA6hWjch9LY8SkOsURNzJ
HHvjC1HOg5HZK4xfy955dxEroBmSnAXLKU57vGYw9ftOMLvc0FCmeNzMzWdqF5VM
XG/uakFpTmbzzg33NMHJdPGV9yxskcIq2tWDP2YOBTVfXUQRDGkFoySSWd4bbxaA
jKr+Zor6JGZ7bs12rCs/igJO78aaBr+es/P+kYkJr371x20PLgSSl1m+TKaQV4YW
T9eo4UjiEvwAPhaYzlHLuRtcJKhFJbgDKZPm2rvytqiJY4OxbQ/XaykQfZIvGGl3
aag8tpvzPinWzMqpKB2dsvae2CIqwhwK+YjUNJTFIlHOKnrQDU6YA2vnVkXaWLvN
WxXUnxzYihbknLZuwjVz2ufRoZH9+j2rCliiZGAPGVclIbiLGd7aZtL7fW7BQc51
OIrCXq4J881HwmS8TCDFeUqt4uN7rx0RphMfsbJPvXnoHm5+xWD2x8zN2dpOSU7w
agP4Rjd8uB4D7IgPgSygriL5Y6hcUgbu2mB+jXXXzm/tI2ZHakuC/nsXIvF8XUY1
k6eX/jvCmAQFDhKue+mR49JpAzMPYEfbkyiJc9HI+hYcNtBHQ9g8+Zc9+CQ2Yg4Z
ViRtvNZDL5KZVywoX21W0ydELeuMlogLzptbO+Mpp0eI13TgaONjGX3fh3LN2AiZ
IWUQ9e1+n91RP7bop9JhIl7KiVJh+8nCzR0E9vi7oBwhlzqR+2sRhh06MbItQoaO
A++ttCan39VVXec1hm5v/W5ZfBNf/OQ57gMmgRJ9AkEMQlI+HJB8FOMobTRWqiEl
nBegjj/ezYc38GtWkqxsbJvcH94dqu8RtwPibMEh9lpR6NQB7V9lckjijqtRxRMm
aGvSuPgRYeI+3M4mQc4drAShgBkx2s4byXcBIcPLIsFDBrka45qz+qlAKag3HQu/
TrWtCaGZ3TwhUZhH2YHM4ObPUtdc5CasjPXS7eRsTCfzNuzLXCReoeOti3qHogcj
iyeihuRY6ulIc9Q+9R92Cqtlp3jKFVHDI3XpFlYnbFjLLleDOSiEy1hJSks+yism
0NQeBuANZV1ZYYwTcaTdXp0yoOqzD9bWfSRfbavzgp3C0sG9EIrRNoIPPzmX51cU
s8cGL7ywkBdElG5TGD1bsbPbSHfEM+C9n29NNcK0HAzm3LfHMcGqKQVkbDhMThC1
0+layy7U4pJZ9A2cSW3vWb8q0T2BZKbuVQ1qBM8gz0yJjku8D0pjnsWkCwM61hZW
4vsTJ9TydewJXiR3DzR9hDJTMVt4FQGTB81oBejBxJnUtEHBqGIjw4KMVGbb4sWD
ASLCdpXG+LVYIuYWkIVhsyJO1b32XeD0UciiPycK8aTIAgWhw1KrjXFmxqSndl3B
VvT/tsdilvlPa237JpZd2i22604BPx1uMTzCfwBh0XM05ZTxdco+Rm9f0f2LMmgr
C+06A8QQBBcJI50mVhiPj630xCZxjeqsUrFN2ZEX+bVnMsLlGOlXTy2WNrTN8R1f
IJrsXyGGEWOhpb7NRbxCaeNwU8ZMDo7k++dCNISK6C/74rHmFYP5aLvuV3/oiaEs
U6giFKdTPMQoXUKUkAhc4l7argkw7BerlwBfxKAapGeDUgMpPU5NO5I135PDGEqc
9/yi1R4P/4PN6kVY2TgygHPE2X9N/oo8hA6CAqGOs+3DybvN9RpLImA2fn+I2TvH
sMEun1AT5fStvDqKENkMWcmqY5dcuxWh7Bu6v4uD/rG5UsZvbIWRdFSzpgwmtn6z
SiwtWfXJo1UpNkbZYQQMyuDzNOb2xhaAEyl8t5iEYT+jhGDEJ8i6zMaMYdT80Aiy
ZfztOrroN2OXuZLa02hlQRqzbf8CnVplxHe0vAr6Rwg1HoGgSc80qj5f5uhBGAw7
ZbKPTr5Vy5KPc4QoPavetuZ3ExUIh7Am+AopSI26pggCEmOWYGImAxunbH+ggp65
GgXcYiv6dP/w5/tgxHQ0Xm7QpDoUbT4eGli0+L2hA8AXmPYMAN9z7RV0WbyUs6qo
Ql0klQWGZXwSPiuRaafiEicsEmQwx1b1axHF/Lup7YJLOHqN/m2IyclHAkdpepUY
Zf2Wq8GUWK8D4TyKKNddYizJ2yv2xrQ/sr08hKrUHxIr/3lH7gNrW7yZ9X/dVd/w
NjPcoD5lxOuvp4MOJtWQ03q8la+v/Q+FUw8IZbs89/1f7ntfyOlX6ZXgV5BWPEtd
YFIdCmtelcEVQdb3ze7RZq3+6Hdt85f2Dy3Cdn46YVwa0gTVJHCCCP1u4HEIRu8Z
G5ouX1QHCCgC+H1YVibLJl7z8+D5xoC28W5bghf/uTrHk8NnDLA/KkTOOyzkq4/a
ObNz6NMe3um4U0lXJ+BxmE1IyEoeGJTaBD0MLXu1xQbedEBJHBqNQdpVwkfBAC54
rCjvAWJ8fyyR9juKHmUSn/2SzAXJoFcEaI1tMvEEpKv2hFoxYPYrP3gPvccNrXuY
JxWcWjXUvPF+WTITd2LJ/usw9nXEXj6ywQw2kzK1//4X4ypRMbnDjnkSSTCtsCbF
YcoCrtDhBFT+czvGB8fh8BnQlwt2ydHrXN29ImpH7KoocJCjZxH/noer4Qs/uE4d
TpPzJoCe+AO1aVMBWixbI10/kkP5WH1bFgkHcU7ENJIKvWIER7IzHYz3S0fX5Pih
JGS1/IPhLJHwOTSH7uF2PgP5jErDlv/ZyXVm2+XFF/lx9pJUKaY1RSeFYXTe4Xwy
DrYROsRz/z7WF5DkjBy4gPxLs8uRASD+/1FG8fl8erICs8CzOSFoDD9cegp5mA/C
QnKjmGd0rjKmE3M2Q9vtAMyZWvuxL14YcaNzAa5Z7AuvCpE0TU7cuoB7tVtCDr6a
kzTxKJ6FN0tmcP10fbngLVmRow2iom+kccx1jLotIA51dwU8Zei+VC769BNrgg5q
zyXU4XX7Ki6l0sQZKnsGi/KuF5uokaTjQ+Rh/NrKYqWzMYmv6o1Ow5fpOGNFcysb
JnkKo8rLEFGuLzpjltwgiSsPYGxc/0K3J4qQpDVOPJNYwv/U0GzHZN4R/52M7OAA
P7H5XnvCmZgO92q5+P9vbHLH47vMEuM5mrLwTuE2VCDiDN7UXC2Kew/2wEmCWWeJ
+uwMj8Bsd9MT04EQgJ3vfZKLsBmgaj0PvhVJfKxxq02GT5S8GrPpswPJV8jsOZz3
dwDkMUxIZZ59Y1xTIQG2XBflttmIFgpbs+gIjmgz4rZYmE5qs+vlD7/J6HhApljI
+BrdELPzombAUreKtBL17Sbg6/Dgm7KZONmy5QrPYLDcUS5hqaX9+wUdNKrXpKkI
k6vlvmQc+GjjQqD3mUEsk4vhnP+refXge3EJiujLhFqmz2b7geYSsz/SFqUG3OAC
iMRQlDHb36OOYeqwCqo7tt3+u4L8tB4ZuNC8jCLCO4KXl8vjyGwlL3cJ6lH0fRrz
4bxVRJuqQD8sGdrSoNrO8Eejl3tbb3ky2zpFijo7YObP+zPxu0HaSl9xL2K68AwY
juicQnJdN38ltSmhLU5YzSKu6O5z2s93Lw3zoOp7SeXRmI9FDHAL6xRpKyqv3GK6
9SN0Yqkleb0ja2C68+50fVhCMFO68SAIQNHbHd6C3ELtvjphRGiCYsrhpRFkZWpU
lcyS0+bcbK+SiMXRPUe6VB1mlAChPArBQaLfA0+IxdfoHGuXYNptR2FGkD25aDr6
zY0YZ0rc879HqEAnUIH/qj/yA+1iAQms8+9YGuOjFJDppUgkqKwmAmUW0h1en+UG
2eeycNb2PtBct8sGk4QIV5Dzxho93kNLtXyKKuqDjqdwt0r64hAdKgsL3fcXAAJ/
o+rDqE0ypdBbeWUy7gLs+8FDp7qYmsnDqiqTlKOwuyzpx9ColLKDUHYJ8JqjWLFi
MwUwg984MoqEGQvo7rxO7CHsb8e/M8es7yrBmFWICKHcwIzQT58htFOlD8U9lgt2
ityQWs4+5hZxOc1xtYnXLvmYWnEEypdcX62e/71mgo8ecmjisWvDG50uEHeJ0N8w
r+/i5tFeAR8orAVK5NmAxcgXqkTAKA4BxtFZ/3u2QitWyd6v6tVfS7K1B7LHWZBV
bMza+JZJOhoaCyKko3O/tMsZwL3wTFPGL9RoGEKZI6B1zV8jd6py1RzCE+Gts6Gr
r8ZPOAStxvH02iREvwn/SY/pLEFUTiQvcwSUrwF0Rt4rsxiEzz7dW4Qt912ecov3
djox2mUVrRNAYM7DHDwxI3wwOtxyymGb6aYLUqRgqLvGJx9W93GHDHe8McNIYDvB
8spq59uSLvPQLhoRDJZsHOFQF90qVS0i208XehzWhs4r8nMxD3VAbB1zbbxdOw1O
fM28vKx0WAiQ5fVvx2viZoGeTrb3VVee5cabJkRVb0lH07KbVqN9CcTM3OPWsERe
XuHvw60XxJZ0g7ggLLN38K05XGFhBtwOgBgdfU9pBnj6qowc/gmQ5MMnD//nwQB5
oxsOmGM59BobUs2ZIF4ZdHNKI75l5VpU5uac7rRzdaWxI0CC5OrdmQGt1XNE9odB
33g1KFIMxJJ6hIRGvedSgy/SA+QdUWvdeCTzXCZ8HKOYEl9PjGKgXT6WDVTXXtRT
DoHz1IktNY7IrCFWnoicdd9fnpHbxqDv5o3oNKpbtHABsdV5J72PTOnUClY7xJtj
Lum+rtAsmWeVbWhQG8830tLfnnv2S3CMIFXuJNspwrRYeyaPBBA3K0vikMnX18rX
nl1BPn343HK7MZJNZpADq3KV9k9FYVku4XgsRSICb3x2p5C5LiZgW7zR7jl4KhwL
weEhxvVaBnYldK7GPbaezAsAuW7qoujozl8nut5I2YGKvVzTSLJVA0A8xZcpRlzC
Cw6XeZeRL3XoqVPzfZLe9JAz4hFZ8/MpNLfghOgH+PNSvJsFq8HHtmdyJ5sjG1Y4
oTS0MoFBquJdGVL3GX1LbToXyuOLOpWgEFEzWzYCUJJAdFprZlGsF6i86/GSyjle
5YE6jCzbo6pWHYqEgUzPrP3gQcc22Ux+w4hxVO0FdxkbT8JVzAE06y2eclWdnCfw
R4xwxxxerHQ8tczuSrdHFwVOggMrZmS5JfP/w8WlepZJQW+B/WFgTDu7gAUF03o+
AzHRnxOkppX3TCKD4oJflRs+BlxbeCExkmYG8XY/ZZSXwAHgESLphttVLAMxMjfQ
18VpKiv4pbEUV6umswXAs4F0/2HzlGU8EseuErH7wdM3gBazFGWQz9w1wEqvH+Jh
fGX4yOFauQyjdUhteMRF7Q1nykjJnD7jT/s5iUjiz+uaozSWIxaz9balFEB33GMF
/PzxVsnBekdbethv3eyHvZIsu3CsF/tICTj9VINxYu8Hp+pEbo8BPNzssemWEg/3
Y+gcR8CPmyubCB5/P9PY5++L18E02ctEnbbm5z82bzUcGAOSWjHoSjf5mAnpRT/N
FCphRiEDJ0tVKznw0KdFSa5NIZuLCJobmEzTWroDebky7+JG5pye0l9PNfAkXAEB
gMl1d1nOG+CgLE5JjARdbteNA3Dp9JhMqobEhAiPLMjbSOOEnFIXrMwgDtsKC6ta
A4rAMDIw3zvKH93NHB5PyBcor33yKW3xbNnTL3Lmc6RepMX4FbX1yGXqVkyWKQBy
v9CyP66z3ZBMETEf7DQBq75LU7SD89CkOwKV7x5QCtjjr2zrySCseVAYmzjMrIL9
vXa+Qtb527DxgvEZSFJJh+rWl60KMHY74aw9/ebcwF/yljRGgFyxqMkfDdSez66t
3fvwMP8cD5YbC1ZU6fCVAVK2eKj15qts0rF2cXrX5eSp8criN6vvG64wMYozVw8z
MGWB4ae7p8wHTEla8GbcBJpHimi4HQNKnL+BCNfP13J0oDT3I5nhw9QR6cbufniL
b7tdOIarHtDFCh+dfnhJdzd838pNdLeiON3aKMzlwm/FgES54bPmAPV72zNGSVBW
+YPcbSkjGZ/2je3IEP62OgGooqrWSNdEBBuQGkQ/hTtJTH32geF07sWjDpoUKwRg
a3LVfCAt14VnMwtT9JF8zbHuEuqpNGp4xLzw6q84RbDtzpN1ui9apf9eAGUyvydz
Tf0r4Rsrpv15e4HRaOm8aGM88sh0d4oN9fqFjCW0eIJ7Lcfe2/Fu4F8dT7td71V5
WOcbEUeDfiWB9f3Zbi0qNCsG9Ir8blEMI5HyeeG9+cs+jkHjmqYx2tyv1DqE6Khu
1RM3EcLuLxTHoqhmueZpPr0JeO0X6IPMmT21semdemxngXTYI3AxqnuhfQhdTLVu
1ge/dMFDpg4z4GZvTYXPkBwXClOnq1iDBotY5B7jDbc7Zrqy0Av86bI+BSKfvOF6
k4P+Zo3i/fOZTIBYLA6WvCItmNe9TnJ6i4S6iDGVr0pMUufn7VgouM/LHOLuvuIX
jPZeFQPK73GpjYOPIeJb7n5uZW6guELnUQqq9dSt/Rz3kNKwUHCMsZgLJYJcbORW
V8+MlXeX9ZM/adE/+uVO44MDjkE8E58o0EXfWYF1WnWht8OKyk3Qg5OyrcjW1OiL
zcl1NfKlF0MpSpikK9xuTSsxMQoQmbzmpKT29Te8JPijjpOd1wE1/SA30THukBuc
JIGnO1/9R5bFeb+8xKrMBYaYDuVn/adZ/fzlejcepmt8rFG6ug/csR8lv2DcnK6z
HQZWEqt1gCXIaVogWyT3Iy5pU1+5mixc63yWDaNH3a6HhfpKF7KgBK0TKPcXA1I+
frYh+54kCxUt8Hxga/5zh4+1J1umHVzBs2b6Po9z4IiQVhie1PbLKJU5T+Gn8fpl
pfp2dpipcyDDv76dm/UjjIVSCkAnSDLCmunhzwV4/ElGRSWI021FVBPQw0KBhxl5
i/rReLA3nfpAiOkcaFGM2eZdrwpPppTDxwlE6nms3FB04/31bX7LTNrhrc77xYmz
HqQJ+6XG8k/uMFB89HfWD2JngNAtxUiJbPbwE3E7mAc0J6jVqcQKQbXoWVfvpc/9
bSVvAAVuDMBOQ8iKi93bX8mK7T9G1H+hy+2Zl5NHvYSrJfFrWEidjw5siv/hWZ3O
6caHpwoY04cqTBN/cBaYhsonrZzMkCBLY4kTd1urLRVor5+Jhg9l55fxlyOGtPov
rIQcbFxn0D0D6rIneemZ1cT5je/CPQLnbrkVpLUM+xRwswBPSga8BzpQf4l8yuxn
/HyetuOpK19Q8R0ykGLrN9Mrhvy1aWGzglwOvOhULCBjOtnA0Y1RKqXKrF7e2RXu
yRf2sD659DBMddiydIpWTj4DTYbcVA5xGt3Y+mGV2ARLVQitxujO7FCW1FHBCxjF
48fNCjjDp4wXMmcQOKXaDnqTtESKSkeQrCJ0RYx5FTc9knKhPd5AAw7g0Qcrz1YG
4+Ih5EOXMwZ2uFRER5ZLDf247j4ObqCAg6JiJqVgfUJ/ad5l+xjB198pxJ06b7cr
Zq5Mvu75+ZUw4BWRpDWldFJ7eRdP7k5YzeZJESB7c+PcYkSdNQio/01uizSf7XJA
auqWOKofXRJ7VA9szNGBuq0tIdMylPXUwNCK1KcesJg6NJqv7GqM9mFVHF3Xanby
0f6FY91f4fWrGtrbhooMO6loVJ7eh0gm/XWBEclnLlnuntnD9n3g1ZTML6QusBpn
cCwRrneWEGvr5uiACkw7BwUmTeJfyTBqPX9n/eXIaoL+kGr8JMXck/EeK9SV0dI9
flp8OPhgIgoMO+MHM+326Mw1RSpqAC+I3bzUIbhUD/0kQHiCu6RABAUCmHxgLUIQ
E3QXifEyJ18bClu7TjkFIJ/srEETdsJABnXZNg6W70MSCZLUtB367ZT8tKxr27/T
upg92jQsYv5GENtsqS+Nx5DgUvgtkBRna05NfiQC5ISxNVmDFyC6j9PUxeE4rdmq
/7aX6mUVNRrIFPbEkjzrom/FH71vRAj74W/5XyagJa5WMoh+VuhRiSy2qHrR8Jn6
8L2+7j1fKcI84MfKekBkTIIwy9+6Te/Odn7b5poCqY2tjPrgkAD2R3/qF5/IqBBG
83E5Q7xh9BKdnvN30vFT7iRQHQJFq5BkCGcWaJyicL/rjbG3Bn4FsFH5VywJDGmo
QPx2Fy+s0TWumWmqcv3eWTZ2N7HJ8dHmdxVNWhBIJnwGhJuERg3us4pRqaXdKcYP
iFMZhe+JMt97T4/GveJpoc0X6pB1y7A9k3fMs1pyOMzoUQJ5DiTAZxA9ACrU2ivB
lI1OLuCSSpA1j5LTCEwazVdzzWUK5D1GAGu0yl/+Eeb5obsEj5eTY4ys50amrsSC
9i/J4fuNEVrI5jAn4wxO1FOsooUdc1q7lNAJBD6nTUVIvOXIl1v5fjXCS3qwLokz
9YwkHeAd7V9Yw/j+SyxY8M5YaMEaqCBkrcNoS4Jjmlj2vjCS9M59UO4ZyqPAkqRf
ZAYcSGVOXDRQgR/hQByovx4oT1gW/swvt5RHJdZMs4SvbYj3soqxJ0l/GjBsMSIt
IOjI/y3S6sxR92EJ3BZocWx9xXbIJ4yJlkHt1dSMrSyNOdsmmNCxXgUQZocMRbzu
JMjPFH+jBYKArOM8+qDtWtsbvbPEeWDWGknbpREkYwDshk70eHEliar3gpxdkbVp
S+HWiar6TA7secvlCjK2Hr+6K5NRp9VWVgKwvcXGc9ansowwPAfIaZtDFT1tpxZY
GqOyE1+imUtWv6cCEjSq6HZ5EAtFJgmur0YZmvSdaeyrHkKtqXi6lqiduUGX1Ess
Hcqs9EhB31tCRNUaqrSf2k36vzUYZrip76dXOWEASQpojjeXgaN/x6rKYXcy+Pk/
FvcPqofUZMBiQywj2gj6PNf31S+ZCiyjdOzYn1xwYelXNWXLVWDVkEmc032QO+4J
WKVfNzDUPeyXo28pAEJfbpJh6vojDvNHA8yZPH6757tPqsPolhhMh6mTJhcM3mZC
zTk8UMSUhM6RK0Wa6uNE6d7svrs4ZV/HJ4QOhxXTPNeE6V0/4l+ETP0jsENEYjkB
Xm/FN00AcmNcR210pSMGxitvSy4Go4t6pobx1HMITL9MJ3pajGqdk57Ye8pIbpuP
Ma8bMDd5fRuce27+QbQdtwbf2ejC24SEicbHJ/LliqsIoIGikeliLDEDZReqmk61
5PWPfNGev3tWr6Wtmttlsb2h9HUVFpcbN8fabEryMMupbWvKjYnPYeGFlisU6twf
NuCvzbWAVRqsMAoVlKdhnetk6mVVWhanoKY11XcZmoxH5C61etDx3aZNBTks/ZEo
d3ThmuLBjvOahonUSRIIyhrU9vhuGFdNxXbz/XBPYRwpWnCkeGY4naLzVwuJMPX2
p1ijgk6ez3augTTI0FypU29RPQopUK+/NjFVgueMknbwXrQGVJA7tqfIvYAQFus+
D0aX8AYvQtPzrtVIj+ToZ7z31zTOXMyuOFjxH1/Rki/ffkTte5OzsQNUREfTzZwp
Ip5CJPBzRH9bRGMqQO22jtE3tWR3CuDJgDWXeckRKsZd2bnOu0OuyAFxhqF4srDx
/KZpK+H8dv52NwK2Ff4nlOGhAXtOQEdSjr8UL25l8OBNU7iCEa0M7fBhsRTTYe9J
InCJ7ZTWpujBdO5cbVVsIZOZ2ukp+p8HCFEIji94Kewk3Jo4w/59p8vtVrWaoweP
We8lu6ZoPzWp6lXK3KQ4rJnG0V9O+PzxFqA+jOv7pR3WGhZcfuEcCQ0a7BV8Mq3t
iXNjHmkYyeLI5Xn+0XKY9Sazxx5K/s8l0KzolCLpuyaVOK4U1GrLz+PRkGf9kAj5
OwzcFWQV6joeyAXupmHosZBjYNgG08RwpLNtgzlLDVGfOLUSpLFrNFo7I5HCcfUc
pU7Hmf2qBrvFAOyVgpgyIUcHETL/0ClqKS4VKA8A7+V4lOBzEEtMFLUfbboGUhcq
52DoZo/md22ERsHMlkhwAjzIOU7tpjoY2zmyiGHcfbSMuNBHgYNgWxq7QMG7/RrG
IAGesysopcjATX3NsYeBtNyrSUCSzzOYziJokb0INpoz/wrDRiXskHPOgBsIr0FL
Kfmdvl2B5HI6pk9pb5TT3G1M56BWYDorr7EtSbfi2nh+4W5LtnpBhb6gq/aQvF/M
M3Ki/iALoW0UGvxGPmSVYc/yozmmjLmHvQxDgs13i/eHjoKTjf1zC4BIMFLVH1zH
NJ1YkSedwlMSK5ILB5YD2p0htR7lh/NQAcJMzaHI7C1QUTzoEQLtR6GOCprPMM+p
ZfxKPMhY9XPImEPt0Sxm6kamhvMEHDTYSZeEeIeBZnwyn5t09c1QdP/rlROaud/C
D8CBn3vUDXeMd4Fb/REyy5Y2nO1WezNLaTxfhN5ZAHkw7qw75tTol21XFW3O3U2e
EWTEyEDWJ6P8F7spLhbu7yT/NiZehewzTK5g1gzFFTLkKjFJpAgq+yTGbDHAJI4m
5BSd295DMBevFr+ZAOv/gCTX+9x6xk5mJmXNT3muiJ/fGlEoCwwtsStn4vBtSdwO
rTcmr2nJPoH/qNbHJlikyel5dRuTmRvx9s15SnUMw2ntZAKOk8y7hZlpzzlJ+Jf7
RVIGgom/kkop2OdfLKZ692os1iP0STETkG8m++3I//mOTVtd5X7oLc2rU/cnjglY
UpZkxA7Ni/FATXIU+G5JOYdE52moYbWJZjs8tC08R2xlwCckscBkuJgBUnwjoHrD
wuApjftbmr/sVlqRs19CBNj+2IwNUXA//qFOJnFngiz1O1Eokz+4X45GIFuqMqHU
rlgZkpEohYHVZFSaUeLp2LLcKRY+rT8nG2rUjVD7Ot9yztzgaMD0Bz1qZqXcrbaF
ptPYfUHX0j7Winuu8j8MalCdwI7NEhZSOAv2W5Qv6h7sGH7Bv4Pqml+FdjdStDif
T1nnPcgDlTyLQY1oMetX1Cw8ZfXnuT3T5z1Mb1KxxxHYnjLtyFiT7Tiy3IhfUNTR
000Z9oZ+wWUzkTvtQdpXckSs88H3vtzPh9wxbGEd/KNOnsDJKEMgWfjztBYfsVku
JjjYBZEHrA/RfXB2498iREgkoQufV5drFsEEl+3D3y46G8NpsOeB5yeLWRic+aqN
MnkWNeoP/YNezmpys9WG7P6S0uMkgq780bntW6U2MDpcCecFeFPQVBzuQ+XXJN+N
9GZp3SWq25/NhnoNN+ddETvGyNvDVd94a4ZarFZ29ZidHOq32/SU9O4aMFw1UREx
3CMFwXwAWPT5oL6thUc89oK/6IkUr8ubZsvXU+S3NAzxRv+Sj8lNwQ/myLohXBnU
TDdlumeza9PJgHBnrDgW74QkY6sBMlz0fCUOvHp1/Uv6LHX7oF+rHitfCpdI7Gkv
7josMeWeZwmrDDmg0neydvwFbqREtoVr06efP6Cx5ljUsBkZ9yP5ttvl53HlQRGV
nWa2eBBxoyoLaHfc1v2x63ePDXZ+sBgjLENlHQbiglL9rMkWmVn1Wivme5qcJ/qg
axcHr+kcjEY89NuDuINO4FlZEsBClB1hs+UWQbfTAkHNQFeJSffA9zDbuISWvCYr
mYYPnVaD8S1Sstjxq7T9kzaWAfsnfc5zCriWLLAc9qlj8OI7dtCg0vz61lARvB1A
G/5Yj7tcUIS1vM+IUOMuYEDGNJg/CMG4NyVvNo2XYgcLx6g3QPIDERZpcfok1hfs
KGAFI8teULcsIockfnjVfh3lrXhN4xfCUYb9zMsr0mK8Laq45ZjC/QKKyGwYavcY
3XP5bYo6dloy8B/YTf+3bCg5+H1Z5vaZUoX+4EAbKOqESNS5xKsiJ4gFboEQvqX/
Hg8OhslKB9vfsLaEgRHk5Gx4hJN/2NfL4/fUW8e4ytahek5Vs7iuU5rKkPjeFQK/
XDXwi9Bc3FaQ6W5IpRzhsbL9sYX0+17X3D3nqi8Qnh0ZyPTnDtdM1zzdoz4RYRaI
5xDEd8BhXqjfR+O/MqqBdIp5DGENHS3JEv6lIiC97t9XE9ZVMGhYWUDapwsYdQ0g
omAwRDrgoyQVARo2q7dklOYnxjnGS7e9uaFwLvfIv9FT5lVg9CiyGbLr2cEZXOyf
87WRgsXB3iakEJG7SxDDyWx3LdbKKCLAvEMWd8uBawxdgnUb2NB11/Wj3PAvsiCk
5PDx+X76sZSEhQIh3uMLCtcizHfliZoyGwtMIZjZQ1s9CN70t2fUfRMP1Rc4G8oV
Afxi0aEmZOGR5Rie+NIQgzU51K8w+1jRKvpnTVnMsFNJxD7NG2WItfs+UIUFlRYP
AgC7ZQSwgBceHPk1mxjN17xPdjgRwNCOctZgJgUuALJVFEhsdNlIny8xOAxTD/qW
yZ/8cYVQmqByJepkVBGuJ1XyX4c5namCv8vETxb9LosKoE7EKHihld+QraozOTFr
mnX9vO6W1N8bv9mh0GTdYb6tJ9OUzWD18p/owICaKYED4+K+IJKF7zGD0AuRjLXX
thMEOkzSLroeKwu2/k0dItuFw96dvnFIB8KZmnTPPpdT1a44amAAQYc3p7cI6oOR
G8ZYY+a2YyDLT53L9Iy9aKieFJAJQNcje5wU2AhltPLbKcX3R1Wk3CQDEAjx1abu
9h4rCAa5zDqGRUYeqVBfaSxWS/qzKsAS3Q7DK2ghXEwzI5ZDkygNtBwdJCEfhOQf
RpqiAGphor4gThYzx3MptWEqZM3Sk19WceAFQyrXSfzNuYcbUcBm9MgK9o1GBp18
YuQSS41WGBlYGQvx0DKRQAgBZmpy1K+l+erOm4dc4AXAf2aXiSRXXumgsnt76Ls1
/kLyiFYfcPuScmJZXrtN/i5YDZitW4eM/93MXYc3vpBW7dn40jkktxm+YB1VpSpJ
o2Vy/P8dIRUMGVkB+X9VI3KdycB3YuRKCVT/70Ud3ehEW9SvqFy/FFcWpEf7xu1q
R6ivbMehIMkHZoxn59Z63FKhPHC3LRPpwz/iFC5nzslHGpgt6uczqA3J4ASG53Z0
A1tQE4k8TiXaAzTXXn62dqnUDziOSDBiUSFZNPftAhccZR4s0C8plAUs1jJGJ5qH
UpAkd51m1hXa1a18RbrCGLaANnZrBBbzUG6a1tvVgDTXHXVCenGtPnWcuEyEbBvN
uSwnCFCgQN1jAhlgMpOfOcKYFpy4Xne8WNvhLk0cwkHuXa2SOWBo9YyR7bYTNobK
WWbWPhL0aR2QaoiL5Z+cPfNPUdcfd4sXiitJJoBDRPorWIiz9P38i+OUfpAuAGo/
Yaqa1aTrE36s0LQaAX0/LiigcJM147Yahqmn0f/o21+r8QcXGKoEoEshlaW1n14d
FlHDTaoUZEZy7Br/CmgDSScVwcAseu/dWK8X3a38iFoXve4uv6AfKPDnpGC9z3lf
/7ivpT6jlXrTgrjKs3+5LWMljfo8GCy6O1yF/72mOxczWaM2SI+0XAU0XoBgDnGv
zqsQaP+DBHYdYOxg5Vkdz5vobWzGN+BpbRAF/W7UTTTkg19ecIqqbmw7DLDhTFQh
zrq1+AuZCElDRYYN/skuWS6G8IKcqjaPYCAgcAPOw47WXDx6uSVsb/aCPsDzJR9o
I+ctZ9nIWiF9TBiqoTRB7kP0yRAu+/GI+q5ngTiLVSriq73YvlVCVC4Tz3KfuhEA
yIvlRmqWO23iQxTSkFZcO6VezUlnmehlGHFitJ1nazT+9zLfj5wFqbJGWH6DlCVR
bSquAtl3S7XwiXLrMIk/L41rM6Z+THYWc3ABSkRR5qFiKrJxMj9m/luq2lAMZDn6
/qvM6yFw3xg/3v8rd/BIgX9t6+tlzX3165fAS/sIVQoWCgZfaac7fjYS2MhGB1T3
qlnRboY2XfnZn4MgD0fk+eE9ihT/Gvaz6dEKP8ttjm3gCX2FV02TKs7yOzqu1ZWP
h5lGdZtSN39qQRkm7edAjPsGblyt34NaPRcJBi+xL3Uo3MQUN89KOBTrx/kSPKyD
PIyNKkUprFI5ezzXfUCjLhvWXlIeOCviXtlwnvNa0RKpj/d0EkhKjZfpr+5KPGpt
CHXsVzv3W9aUBnG9OQSSdoO+2FpGmNXeFWwcdrCubXDGqljGxa+GsCMlUBjdFoTW
OFpxzprU8R55v9gejo0r1m21V7Vsu0tBdXwN2fGXdhCa1K6r5/zZQr4+3i6xKdQS
z/ahdOlojMTvpPtrfUKGC+xWmtALD0WCRTPvB8c0AQwRPe9aS5KcKGMrl0ycC3wD
0g1YDCEBYoVhghA+JQxX/Fe+wm9Uz1QezFTmpTE1XzLeHURwe3ZMTQf0vzaq5Eh+
x8q45se77sYCuBH/NtraSviRO4hNYh6b9tskjZbhL3GeHp3RMPqgcAB+UpH8cFAS
/TLMmIYjK06SEKWaG07q3uQ7XVY+V9Vjqr12KVm0X1GTFNueZANFtALGhJZqIgr+
XlskjXSniRDfW9iAC/BYOQYnXn7i15uSil7D85D86i1VXJX2Heuhoq0xtHOi5w2z
2g7blfF1+KSEpzW2NdeOOmcWd7vZteJ4bKw5fFgY2KPsc8gEicsiFHsf8xNQolR/
ygE8MwtUgXNjFxLqUZjNkqYaD9B1DCSl9dF7dncZWkyBBgYWc6aZjvTMkBY6as4N
THh8poiLC5vYj0b14DUAYjQs1/4aTmPBQ3+/wvlmayZNky49sU3q+7evlUKWHQ2L
jEbNdDjcY21a4wu+kumNIsddG2k5YeNurtBcfL7VgIEhaXaefb3rN99hvC7bFYgW
yKrVf3b7hN+dHiN7I98G11EIGn0oEUodYFVTKNY+kVBu9JKIJeefnW2gN7JJeeib
3R+x6T1Q89iMkqsjkOsnWiDBAwdqdUDn3hXsjAIwqv8eD0zyygrkEskmu5hvCD0+
qF61tQ43f32RlekZF09FtGBlAh7kqwP5uTextOssjtY/94pZNFY4DhtzgqlT0XeB
YEfvKG/YwgHK2FadMWFeTdc76f+TIrbmJhnPYd/nD/FyK8OQox4+Rb/sTRyVsCXr
UJK4GFSKq3Jn7+R9MiIU2Xjf9ADqGWVDRmW4qgXJi08XRq1IIDFkQSrDp5pM3m3V
SN/zBNw3il+sPaI0WS5Inz1FS5L+UmIAQfWIUt1MpHosjHNc5rGtvCZIvs3ZodF+
FkVi26yA7jLhdqDbLyZzx5PsivItFSo5vKNZMg/i+jO4hrRohKz09wqYi4TWpWfu
AY+kXUjJPohZ7w54kpMegM1wG/NDJtJ++zOitv+tT6O8nWdhdIXmvnY9nf/XLt6H
XSZPFc1aLFi798pjUY2GcD1uLNCDm1N673C6UFDMWLdZSWQdeTqOciGMTjrLm2Yv
EeZPvhu2najH/5lKuD1SsKbrlJ69mHVvVKP7X1MhwnGs+fdBD3hpSIF5V1XS+RTL
LZwRmdqeHcEh6HICdgz8awyrhv9vCFZsJbpibrQF0Sg4rwVNVnuemVgxeb72cUGa
pjs0Lv4BV7nRc2QToCksdwZjMgcP6oF82hroesPpzjdwkgQAoGVfBi44EpcOb9e/
P7ksYML+CqaBhIL1nt2PzQWQXmpqZG3td+SaTfLY658nlJv///m730L+W2qjH639
hIcn9dSByp8R6uavujTu/U6t+eWBrTHnT+1zsRjmf2rKIRr1btG/y36qFWLv86cR
fVCtBrDH3y/Hv1bq3Hm4KTd7sPvEPaBpmXXkqQTtFLPTMGsb3p3OxgVik+IBsfIc
X8KTZ2bo1H+o7+QCatE25v+ckjF5WEWaP3vSZFvxy+v3HlR4SAlHr3m/MRarDKkW
yHG/8AVbEJNHuZas111uqs2YyEhggyfyaNm8BT8lQ9BcN6PKwvuYKPhnBimt9/Fr
Jhd8EXQ8wCWxXplpoSyFcbFVMhd5XgOjMdWH4QtSoyWqaUrn5H0Xn9XRAhO+X4rx
/YjNW7BDVBPig9i93YK8UilNZI8COOkgdbLWQl7mIarFMusnocX0nzKy8gme32Fz
G6e0F6+a0EJfoVefjmnURsI2C+fIYnneu7+J/QPiL7Cp/p1tArN0SRTDblhqpWey
1U6j+AprTLEtLOclrzwF52DhbPyzMqc4pZSFieEYXzq0O1VlNKs1VFsCZNiHEW0E
8VM+/HQSTky+qvZC0LQyasHjuWXBLtpdCOQvsYrwTUfTFJEG1KQHES1llVaOuzo5
Jj+W3ljO18jYdrMK2jG+K4AGDByWwFHCK877/oLxsuFCq30KobEjeRa0Orja9ryu
KdfpACs3rj+0FYKRQd5R3KDHkH/4kkElz9UYG5dKMhENlEU7lBA/lSk3V5fcf7uo
D3DnKpuUFxjhIeNnpWngDQsSn/nbXvJAQiPl/sc7kvHpxPrc+hf+zdr6i84LIaNb
nPteHbKTdUJBUihBPA89gaywypatN98dgu9tkXWRfN4HpixxtuyYNTZD1Rk812WB
fA+wJfiwbPLOZyyGO8KpWJCZ/g6sbalIPLlsQ/rsRJMpcduaGQnsD0NsABZyr6UN
xMRFnVOmw0QHSG+76dfgFdre3Y145V9YTFLwdGMC4SLvVzRxwPuKOGCDyHXpAxo6
GwBCJo+30PMC+7PgKmYMnQwS1Fob0KaRXA8QpT1oOGBNwbYHiWJuNWZRs0xm64Z7
hCp14FMBBkUtlOYbb1A+r4hiBM6bpfrKkAm6W0k0qXus87MInKq2ZgdBEIz9qecb
7zhW95E8eJEm/NL+8hyqHJU3ae1r8N/NHhTxfl32X4BO3DyPnlx0yQ7ahoaRO0qv
P7Xrog4Xh91gBTqPsUdvJqJNkZYjR4FO1lzhRhUpbJQED5xu3CD8nVtInOMxFrxf
n1BLPcT2HDCXPZgPNpykLMTXIba3n1wiffvCWuTAcbuKtVSDln9XSv5jFwJPfKNe
pKF2T+00r3PnNa/MvbVoywxOM9kcR1w9xQUMXz9Z1uXfXZf0eh6WK+ay/c678FEl
X+S4rLjA2LxjV2VtP7IN8up/qXL7OkGTjlSnbfppKkXq9Wy5OR1qlAmSRgzgknoc
/ITquOQaidfSgqfBgCOLgm7M/jzghPMJZe4fynM40eNQ23c57W++glC+KE6vMdO4
Ty5y304NrpfCoX15cboON6shw5Ck4QzVFkmNCre1YnbDZ1ANLY0OlwX3T1QzrJSP
IiTY0ggoa9OC+PeIZAY/OGkgRQYnYAjd/kMoUQJLqd+a511wDLWAPOZMchs3768B
HAmcweZz2Q3e9Z/B7fpaIfFhuckE3JIRUZG7n3ZXCbKxX1SosrsP5FBjyVUELS+K
n50CARn3MXDPsPrWGx3QpsPhuT+XhrLqvIKd0MApSgWSghYOqAuIjQEHE+/Gq+YK
31n/CJT6Eee9rOP2EDB9+/2+ho7FZdMFlujB9D/yUyNGQAxVYJbUhnelBy/SvA3i
02pIO7wiY/GPMtVlc89jIs9v6t5/f8kS4Rgw1UtoAQgEbbqPKn6uI7akdf7TJEku
ChM92n50JnfYPfa7wYRMv6R2QMqnUV2J0p/tyoyawUifaleezmzOK3BQuocDWXAQ
6Sz75SndaBC/Wv6l6wBzhkOmmUA3//8/DJyaZ+TVIOMPQjinprGmkHRtamIP9K4Z
Diyo1oumnXJLPFrJ49GlXQ1z98qGnWj2wgoUKvO0Vs1vhA8yMDq13L9dif5e2ThE
B3NmJ77qHLbs7+MJxdCqp4vC5kq+fdj8XnEfsEBV6wi+MLR/X8I8DF1PMOnZFxV0
Yt31DbYUnIOGiVY9xVNXQCLV37Qeko6gFdn8bqMPV3UdwL/aqRN8bzfjmQQfiqt6
SLbr3mkmb6PUhGoxNe7BwrhDXQoZtOcR/Pid+6DphYLAxW5tXyvEY1dM0tYtHmK7
Vztn+Fv3Osi3gsgJg7dRb/t3DAy3S6UB26f9NguZyFBgh6KCetxVCQBYs4IVwwMP
h27Z1zB/0+vs5Dvb9wslB4+5dNf+4xHrxt0vSBJtcbD4Wwf2xPFLrDcEKtcNKA0t
U2EtFO3zRebSkeMuC27d4C9tc1bJZUpJue/Z2xx+O4HN3tXBXB36/qh7mXDlzJET
qo4ts0BktXCgg7gRTI0M/7/hgl9XsEazRfYJ0NESKgMC07nQMa/FL6p7Ofi+1FNK
0TXBDErP7l+3gAeYHGClnC7dCTV8vodBnzjJRLHo02tFBkWEDqi1XDLG0g6PWpbs
9nCCGUIPSKcAa691repidE2IXENwwklafiOjx+t14Uh9SLR7zYeeCBc/vpnOugx/
OdVwFpj9+F0At5VgRxaZqTpEPBwr638ZzeM7l1XEXfgZfYovOiGqhMPWm8+LeXAv
LACnkXS8cftiPrE9JP2684VwhQxKZ7NW30jmFTzMiUg0wI2BZWBTcx4I3DYsg9ij
9Pwuulf0+Jco7PuZooFqM5KYeroy08wdkNH5OkTgYktOdfTVOJ+F2sB37azbQXKA
3glggyOk37CRWDbqwT2epUZcaA/iCMCfUeg6ykzllVTAi5JnEz766d3CHsWqh8J1
Duh9s2b1lInv4BAB34/WvwTuGX4hE22MiaPZZEFSVOVXF6ZnOwhUAQrIdxvqUBgk
5gs0YdhCwGvYO5DfwvfLorHq5F6WqgEISbBJ29cbxoOgfimBh/STM7f+PNXVk4U+
1u0OrX2daVo5lLJ4thDlyV8dEdCsS3c9jhbSgfZAtE4VKeDcgY6/R7D6lTorJQ+g
JdVUUb9AVZLWMIhNnsNHZUsvFFCgxge4TyFz0cMSaWNa61kOECBbAyFRaHXbjqEd
67MMsiKMWbHZSSKq9eloqrbnvco39kjZShwxu3amJ+NBRochBw2IOqi6dR6bUoNu
TJ+Mw9aSPnsL7EIk2lRjUm4Iz0ZZMJ/apCjbSEIJUoqhbb5yPCCHWJVfJY3IEv2u
n2jF+NOT0cdZJoTa/ZuIjg/W3XAru1nEXSAnmyWGLml+tNmXOdlhwxJemKwT3t9m
grZeE+D0gJP5oz/FFIssqcqegAYkhtBdHP4arQiJIxfxTifw9DogM/3cMCKpegPK
JRczIhoUagbxb80C+F6lPRfn1tJ4ZzIeFcg3cYSoTmyxPMEqfdgjQGpP2MmzkSmi
MEcc98llDwzBRd63p2EqJilfhW6DIxQu2M8T3ispi+MFNg3/VlE3KRVY4hg++E2Z
sDASS2XQbs+RlcZxW6dctc3STa02bvkKN8ZpZHFDdwigNOC60FAEcAEvSsL6kHvs
CCTw5mh6oRjpQuD8zSPrO8YD+r4vZbt3dXodObR3pDwfXLJeB8uoSLzbwArTfXVZ
qsiaDkVjy0Rgqxow6tWCCgG5TTwOtpR4VIr5do4qR3rk+mfTRC5yzsOJUFhdRIj6
5TRYEv+6ObZp0If0Sdjefx4t7Eol4E9FhK+WsYgBln+KPoneC0XSwSHSt0uyF6Iy
Na3c3fG7IdEWEkVMBuMTpiu+9M3rmM1DuVMFIUNz2Bye9Eh+yXyi/OQ7vL+c08XK
Oj0Bb4Dv/RYWerGBBAMkzONefmkgv6/3Am9aVgTYaM3RyG8k0Nj6eux+pgb2Nkid
TNTiqoP0BHgXJAJF2UUKFP8E2RHmGBkjTjChJk64crCiCLRYV6TjSSZj0V8kvuLV
GbWTj6E4FkKJsOEZfl0/4VJ9rjQcRhi3RW7fRlTWFGxiKIfDuIR84v2qMpHu16g8
xDInmuY9LBm6OYHs77KWnlku57Hh5Ikol2ewRTZ0hT5eblXvRoPosvo0gFvn+Tg9
TDzoPgWwSDzVG2DC3fivpzcqWxrqrI38u2q7fXzpV3WTMtCmuGnkv6J3UOLnM96A
+Q/Lwj2Ap5G4r9Zr3tcwyMKEQK8xrQGMD64zqYbbcZ0wvHQFD3iIVB0LfrcMeuXb
0MlIzd8Ngimygy8tInJDlzYqdX45xiZI9snBFisnI1W9ezWBIfLnN9Vh9t48diSB
ycOL/9NaQCe4moVLXBl3uteNVSJISxs3utm5KeZgHucfDlSiRv+781AKk3sbznL5
M9hUia72YlaSqDhfPWLCvLdgCVmpIgWSK0OnQlL1/Ah7gNfplOn4uzhqX1IwtRB6
5Nc6GPs/NNXnOgMp3Kr+VvJZCFld1GtFfi2cQrxqrFU+bnTH/mMS6M/WKgYPssPL
pjGagFQyzMatdfKzhbLwL5esCLSYrROMV6zVI4gWDkZpcyH1wgCGHq7UF7fEP+Rn
zeKH2JQW85IsKfG7dnOavXWlUZ2MMyi75vuHXHeYB2XqWQx/vB90yWD/VS0273WH
X1KuCVIXdQgTqNHcOFWYeOaR4YXal2ZX4Aw6h32GBRsgjQwInWNH3cchYgrnI4Bc
ktYDQgPLsCb6JPwBZxt1DQZDg55z4ixJd9ljuLPDpBVD3zCwP3LwfXjONog/Ebov
e5VPyekeYpEoYl2zZYnSscfXUOv0f06d5ZPH7gjs7O9a30b/PdpInKSEPiWLYPBG
hNoVpHy7ztA0wemiaTNb6vghyYIJuyonDhQYjVCaD0fgyFe7gxuW8W9HP8oQk4cB
oEejvmPV4avYYd5t3kMShNeWBBo5BWWk6TBQ3aGaPobrfKUiUpbjRXh5Z7gsx8BW
6PachZhwtykDyUy0S0cJHDsB+OhNTQrEUJQZJvwqxOu6FmR5YlP1BDud1xNXspPN
EWU2pEVbwYpaoLgMj8XEyOLoCY/V46lqeOu24UwFx9zENODVSlcC2720UCPMtDuS
ulH7hJ2vnHymLpu78fptB1CwUcG3okWlBSIZKcb+ZgGyDpyVyO+giujNw55g+RV6
kjB9MwsOHCzEeN+F3G0DUEAnnSt2UE6B7158tbJoQTyHLGcOi4mqMv39405gLX12
2KCkbMil8VtWeHuDiamtUeVhN0+hqUyM8yZq1jFoZZF+iDqKPWWZ0+U0mzDbw9Pm
G7I3uRRxY/vwWPXQvtowv3U/+LmScQ6fgEgY1tnQFWvdlEZARhOO3bcKMiM5JCJ1
Yr5kRFO05YKQGDff3YAdps1DuWdsiS0vHOHPTMHvu2/b+4D01dLM0KiXuit2nK8E
Q4Z7Yi+efo/q936ess4KQrTkFkRDcmpiZWJ6xijcOr3jojNkYdAzUBTRdOkRsgkt
pcNaOYEa4N2FLiSFUrcgx6/SWGrQEA+vwk1iGAfC2bOBMdRJdm6SNMO3l8nutvxR
iaryMhlVRxvgfYcSLPCMCmoM35g+pFJudduw6KGQcBfzXmO0G0t0lALlpQV2s1br
/6fKqUE6VQECtx4tUprzYyWCzYJGAsLFabp2gS660M/+Hzcxuu3MeyxGrpG1mdxd
777WbuLihRjMXDZkdVO4fyi8aowPCxKFzCwAozT/qrUtlhdH4y2ww/tmcruReVZM
XK6xxqFKPHEuQDmt8zgb3EcDzV+WQB/Q3g0Mf+sj1/D3wIOElHOmNJ0RTCCZqKoY
002fihyAddEfvljHz3BSvCd4rzwC4LljDA/o7YKquobxvzTwXcTynQ1rMFL0UdVT
x15x0BLuwwctU5YXrffTtUTd7XnA4g/FQ3Ls0nAHOlOHN+CT1W1ruSKg1DCLJzjH
Jrx7ZVtEn/JbVOE2ynC+oo+csrYEjlSmzK9pVfkFbe4hrf5zvS/TwVN2U0Bawmyy
GqREyLOGBlGf2uKoOSfqxazLzDmKcX+HLLKNsXS8pArbhUE63YWf7YAeMR5V2J8a
9+LIZfLJIz/UbbUkbV39Ur2IyXyMwe5lnYtzl3k/16semDPdmBK1oTN3xwQH6EKw
2JxdFPBlhfLanRMW7Zj0JPVty3oWXkadfUnewSuM2ysvlfciLPyeXwMxA/jcVEoI
YEpDzBP2U1OtO4CqaG+wuaa5Cfx8VL9xRaR3pRO94Ii7afJuewokmrsWC2FHTcvf
zEuhimhzotsLhFHrS1YFT35BNf7qwgcpOEElDXaf6iaNAK+tuqTpGrUiHtqv3slK
jngyadSU3RXBfHTPw3JiH4N8oJXmmvpO1T7DcGNmPCM8ZjCPR8Jej8a2pWuw0Zin
HfIjD7AsuUVWDTTUbORQ7Gv18ls9i3tdCHnjbA+hboeULTtEjYJacri2cH0weUPB
+qQn/lLAWt9nU4KDeUrFurc+p0Uf0N8prClEpxYOQX7v8f6GhFQH0GoiXSoi9NhH
JY+H6hhvluO5KPPE6yQrHdg0N/EASK2o6hzoJhU4FTDxgtV7ZYkh7MBZSynp1Kii
1w4jexW7LScZMLf0iAZrmlyLEpfaDCOesm8+a0F7D74xg9Ta2beG+49D+0bfmnCv
Nk141UO5feiI+rp8Wznuz5vxJAVQyTsHYqViUXufwoZFD4QHmhHu67T9BxGuA/TN
aRv6WAJSzrTwx3M/d3YAD1X0ROBlM+REmFysGiS0N+f7F5eYdHZJLwH/ECK7/kk5
oBwL446IT1836SnZZyBtt2gcEJ0w6GFd3G/VN7KAUxmlBJ67Rr+LFgKyHDtJUyle
mUKXwiaUpRo55TnjofyoO0z1UvLW5SZWTY1kN0knaZbmaWuh3aZGgz+Rg+RBLRNB
bwjl2FRH/lmlxZWECOXSdVfQTqqB85/0f0eb50lXTQG2AyGwKCWB0ec/siJv3PKi
HhPo2TeVfuedqtUc9e/gUHo5vDTeRG9B4zjgnwfCoBhSW+Xh+CyWziac1GZeKFrd
Cxx1DWGD7SkJttLAKmfUz2BLTtkndBimb0FAWR66Hl5XJPA5X2Y+AccFLncvH1Nu
ICj55JVzIQR9ypXNHoyZZseUyMuZhltzuXrGMEylRZwXCs7BFau+d7ZuNPBx+fnn
bvdGI6J57pckRL3v9cwiEvGUYlc5g8AzaLD3hToRmKVr4v0IUD7uqfgJMp8npWt7
y+L416J/YQNDbQiX6T9keTq30Kra0J8uImzYl+iIs85F9aqvutsVK/WcUZ2z0ftS
xjTtDpS22t+JN3meGkIINQlQ0IxHGBoLVXlcoKOiyNS5WpQB4YjEk1ie7v8VHb6+
oakL5qegTVLBliBwMx1msw6NAI6spq6zvnHBOQRHr26C4Fa0kg42naNdCjBBGCs1
LIBJTDU78m0io0+JRqWOPoLPkDmC4gg5jhfi+Yyr/thNozEhCn2Eb4I7dQZpYAOp
yDfoqaLPz4UFcAmgZ9fLV2CGj9NzaoZqa7Mr+LDCDxTou/OzPrXpGm4XQMJPw2xV
yoAwnsswFGmh8g9D/A7m0Yq9fH8oVRQAXiQ5McJbD8mw4kN9coBExIj8d7NlqiYD
73qk59Zr8TvZrgCICG9qgtB8jawYpnhDUG6bgii4wUNJhtfuenrHHiCQ84SiM1fh
Lh1QQ4fyEczU5cP1DVs2QqLMLq425uY2IEaXzS8w6wQLS8b5/MDjV5grv5c+GcPW
Bx6al0BUNVmgjUKVPnFjTqdO7tezAx5bXpZi2fQwdw6enpOt9WHkeAlyrSxemJA7
XgLiHHBzCNDJzVG+CDDHWzFpDUfhhUkH5DjZf0EsrSI04f0LkRyH0Y8iS75Qib0I
WSrdVmDx6DWW+cyUlC1xDSE6LGwI/cT4VnA0a0Zvj5wkZeIX2AFiBeZWB9exzL+t
deXeOTz/YDBRYeEsksZ/zfCcOFI5yFvxLiLEa8qlm+0IziSWn+u005MBi+2J+MJL
h55gMK5KYLT4Axt9zjUa7hOxlTEtzySzMdZmCnQXFZHCiIJQ0cLH6JWZlxeV7hxC
Akqy7mC1Ipa9BHOyY+s4zKUw4iiJ1xnCgzq0LKSnXr0KmEripd2Rc9ahui4Ex8pc
JkYbJYv0XWodz+IYn/IfUJv6AlOuQd8O8Q+D2cGkyB5aHQMHC4Yf9Ff9GBvtP5Sb
dneNxBX9uf8UutNkDNyCRLlS2lZPdV4iYOW2dQ1Q/Ir/tf87aPMl8l5qiGeH/IJm
gRWrxlS/S2mrQb7R+Tam8hnhlwFzq3xbMZAnQz3N9i60MOhQ7Y13g7tZneQpZh/z
C18syez8bjsrLIZiK087c1JYduJXIMpyDoN0iDRnJrQm1227Oc9Y4J3aXJqqQCfZ
pN8jJZoVTfx7fQBnVccAtadQd1XrOjUMVQfJvZpxfCxfY6Vxp6Q1h/b4qlMaNi5T
IAsTXNcKGOseArksHlaq996t1+YkWmCa2AsijbRBvwZTz4c9BWjmqes/HmJxP2Wc
ddSrdBroAMY8hrcyusjmZEw3llHFw6w9w/EAhe6S+wrUjpcm+ERhf/jDWJzeA1L/
8GmWTvdtS7Z35XOyJcealefWLwmL3QkN8+f6IDddODd0kFHeYg/P6nmaxmMAbQ6I
J611QJbRzhmtzE3ayKZX5Yo9nch4X1LRPb5q+swZE9XX+YNOG6SOjUJN3SwCeQqm
2CSt4a/TP8imdl5SoXsJwpUIlNHhtYikAzIFrA3gjtx09w/A7s+Y7DKT/Bied7pa
hJ1RDQWPY34juTG1A8LcmRzMdyK7bGmF426OIlcObNXMtqcIBjhpLtEnI/36/es1
EIkC1nHAyXDgWGbDLs+Kwp4IioS/M+ypgbgVxL3Fvl5i5OzQmEoqct3IE46Rt8Mk
STqFCs+UK9+/Ng0Ccjq1KeHwReJnUKqFjZOzs5MHcnjBh+I4m6mz+jlw/I8t2O2I
ZcHz6GZpDKdAzXAx6E1alGDHPjrSo3A1sbNaBvb+hZc7OgjDxvUIi5tTM2CYlY9x
/omiuHMJ3V37KNJMVK5wZtpLTbX+ygBltwZQZK9ZsvuBRbPT6xVKGY0vMFOy/9Ap
31k0qh9lqjDKv4uFaEvqKfgs3f7JZt4wtp39gtZv/MLpQhdXGMlZbzpthKSLWfwv
OMxTR7WzpG8V3un39Ndl2Vg7koF8irDQWOQtHPTK/JkQuJ82OZyujyoVvCT5wRFp
tG6D9yUnAisy/luQFmWu8En4jildRQCcaIMMJEXC7Gu1LlO2Snknln1rIVS7QbbM
PBbfYH6tQQnQrY7dXpnh8uvoPm4CGmYuNHswwePg+xp/OZy520aogw9yJAchSDlP
BCjt0/rtYQ8kdDiF3AtBr9SaGyzlwGUDfsmh6R2GsgmHYEw+RLWqONUWYs03z0kr
fs83fR861NEkK9IValoAVhPulSkWTsmqAe1YEQGm+voNxYGLi549cjhiUxUOpnUZ
MI2wbT1ggknfF+RoCz3Qf7OwwJW7MXkJwVg8YtEvyLzwouZkyb3N5fUuL/VmBWzk
itkEaSYhEuAiFmOYsqqTPY326WX/MWArwEzobo28PrS7vdXusZVTiIMN0OODTTP6
u5jkRkEAcw1uhjZ67VFmANSvXA7cXlE3mMkqBj4AiAbBRZvEVehPFRarXgxMhr+B
KLt7Io6AFB7fEfkD49djLeJMrO5wpGZNDuiWN1IRMfztGj2NhguIWZShvvlJCou/
Qges/JLaVAL3GSrEgudi4OH+HoxXTHAGPEar4WuY7NHklE+gKCW5Zml+eWvCOBy+
jOPbW1eTjwbDdl5kcWdqe9hlSqoNNuPOl9yMTX/ZujnD/ECkioiH4Z1QrLjuZvW8
8LSCK/xGIoXZpI0xm79uBwdj3CDqN9YM6IzuW14gOhsLjTLv2HM92ut/w1T0PaR5
ZbdHbCh530X/tqQPC5ZoHZ2yeJokKM/l03sJND4gO8aSnyQcloEG2ZBC3arfmydQ
ZWcehdNfgoAJItC25K+dsLTN8w0sjD2iVg5LTB/frQAjZfhzf5Zx8gxqjKknLVwQ
Ghdk/I4yHIGISpn6FgvebvkKDZ1+s3cA1bJnj8ziV9HpX0kwzHnnBIHGALb8ajDo
BQ4unc+h/J72kbQqn0/TAOCK5drygVY1u0m3XeyHGE/sNZev009dZ/5/uP8WxkK7
7FZdIi49vbAc6xZIO/LI/ajhpXb8QH+mHZ+X13HQnCnhSjsiLO+ux0NRuu0hF4Eu
/9aTs4zCX22dWT/7IkF0w9i44KwOAMoA8D8LmTIzD/15ZBbhIdALxEqEAubw2atm
hs01L5ZYZJCnJB0pZONVJCD6EaXZJQ0WqFPOv2KrBfArUFMi8kw70PsrfBVe0rUp
5gfF+PWLJDi/w9k4E4WNfHSY7VGjwct3T+UdfhrxUvjjDvY+QydDdf6805RdKzHk
FbOa+2RQhpH7n835yIvLCUjvKQ0PfN1/8BrpbS8hEDZCtxyisstNwxKZ5sV9cxI6
31vT3tR60amscdPeTbQ7nXUvjmX76aL4aHGAiv7J/2d9xNRRY7qQIwsMvp/Lk3p6
SUj38Z6ODbQZlMR7G5MlxKJscRmgxmtTOCpulMo93IYvtAyfsBN7IW0+FHUykHV0
Yv0LLlbK8576mFBggLHtIMsdf5QkUZyndH8VBxxeA6io1jmxPt935Piyq7n6XKoS
wXy711OOgbQxAEXlN0XVcnCARwS5rhCv/NQLjVu+OPfacfHNFPXkRzlt8UOJDvFQ
H1bXcNi5641e+CqrRWeAMQ6VM/x+WRL2wJPy1cVx6vNEqZjTWTZ2rEDG4WKzT5G1
iMaUsMIs0H9DVU4hQGaGcZpRWp/2CTTpT4g9I4x4zusAMTxEIprYrL9MX+VNK0Fj
rd34PFuxBcSa+1v3Ry+6Ei8CMdE12sEXw3MQGMKZdjs4zdBVKeDK/fMhjfFFPclV
8A8gQNB1SFlHYLda+t/O6glOdy5hsTAJaIzkUUW5ug/PqPcfJ5J6IiFz2cwPxXpr
PcgTMa6fXk7oDtJqK8xE25jZUJDCbV6oQyya4WuZGJxvWstUCA3oOdjaoY1UT+6l
QQg7LuFfX854Ac7K/YFiPl/Fqg/95Ss1Y4eNhFGoBoEFx9cPWMFaq3/Cpc/1YnuI
n7lMreia2Uk9z4Wow7odqLTo23XzAJheYqbbw9PmMWcqXaeCSklHZtCclpIPtVJo
87SQLTcVYOGsAts67z7TQYMJWUYmKApvNglpyt5V0nzcZvL2ZJQRRFjX0Adk1rag
hFmu86PVXMrplrssdQ+4jbp/KkmfbFKH9JmrQMqU+yJiuyaSEeqmKeDPtWYLzxLM
w3VC+2CJanv9ttsRTeKu/XGFaw5D+yosC36PeHLt71AYszChmq+wjdUDBAchbDMT
wBP2YyEcEjJnGrM4CBCLerGMnWLhZMTUD/kBzoOxT5zJzrZsMBAzE0TvtQGhVxQt
WTH3KQoUL0sr10KW1J8E6EcP8Bt4toKYt+K4N3fwMvRzCS2ibXVpMCHktowqz+h0
aYHRoQvZLuvElC988mbNlvjvGvqK4kRC3n+I43QgFfAdxv1WOHhkHsVWxJZnXuky
bUGyO+ALmh3xOlCgJ5DF1ZTTiLR9D/fpqWtlKaksYIzIgZ+umyTBh3Sz3L5h4jgV
2Se5VcWADh6swkzGL5+QL7IwAP4CU8MSQ8zHgJ+H3rNuHKesYCal9XyBhT0o8+AI
ibgnp2pq1a3BtWg3f1QqCBGWzGN/IiMsTzlOto0HW5xEmnXTr1sHng1Nx1gNR0Jq
vZd6kaY0CMe0oaIVqfNvO/L9+CHamkz2O/D+EJ8sxQnc2CB+uC4McJavfHI0n36J
gANrK+RhfQf5Kmsd3JmBGzRf3/o4EtWob5jquWoASOmdaV/aMoDawpxYfOrJOE3d
SRLv9RTxjlmKn2sPiBmOj3ZAfuJDFyyx/ItWGeiX2qpsMcse3F3EIPtY0TrbHjtB
GmykwNuXmIcU/ABg/Ad36/KFiZvE3MkuWmIqQi2RBtS/CDlAgvkFcEC5bG+ZxDJH
x00F/y5cHgRAAXQFk4XsZJoqFNS7rPxJEj2kCSqIrcSpnsmpPvOkrfxIpEg9fWlH
fizJop9uKIyjOCpeig6e9Mh55qEp7ZBSThYuz7gPOY7iClOCeKG1zpc+QIOWD6y1
oR/S5Ho2gfuh3uwZqxT6Ort8oRdw86rIprDfYQGbwPrRlwYv2W7+tKHD6eU62Eb1
i8h7Eh5CwJUfMiJanQBk1da3Is/sBHjNmVld+G8D9aaElVVhAccorpK6UKcBjFQO
QlkhXbCmkVWrwVr7Vtkect2NWNxFct4PwlXML29+kmgUh5L50902FqWdqwkir8n2
wuBqEwAV04co9I/MlDx55kMuEb2Wfb7j9O0OrfIB/iNiH0D2iU16uyPW5Z97p0Xo
DdLt6igNMVWE6nHZnaWXH0tkDBBO67lpMRKjmcVLLfMc6/R7ZZVtSGjmRWKo7/2T
IP7Lm2T74PZ2qZU0tnsgBHzh12UNr7d8Zbi83GEx1Ims53CQBVovGLysB9vMG9St
mZ0B/jVwFjolWf4Iu2TUnCSuoAyK7o8D9gppcOikIBZigRwBJ2Vz+P0SQssfkjKw
B7KO86vuWo1Sd0Dd+1GGujUIPrX/tg81TBN6Ji9SIrwkbf/mZweqdhjVT4ecXbMd
dGDvIih3DPUJJu3UXNSOYg7oLYktM/NrmmyXQPFguPQHrEHJPXyvT1wcQSKjN8Mj
glYT+P23g5JDEq877iufp0iMFKlMDP+PHMnNmE5Y/tjust/CbF5qNePfM8T0vIOf
ZzAQTasdp65QFPbF2WcvhktDb14OejdAaOf4hdDEB/TeHlLOGtU/62tWvzhR4bB6
8MQGvlhTkXGfKu5py4x+vo2sVVKMDkcwkUpyzH+DGGAZ+E56ICgIv7Qktv5fxtBV
JbiwGbZEkZI+GUsbRw/uHaBc1PdDzAAHKxN/D5ugFlGRYdiYqImzvW5QyWx5fH7y
HJBJ1aUj9wqSss+7GxpbwXUXr7I1L8L0z4UQwjNdR7/MJVjtrfmXNAI1ZZAakwIR
FQl6xY6PxL/b+fwrwHMNoJDLRbJ8tti3KI88nP63iLxR2xFpdNJoWSLPmcBlcSsN
RZUIsTKoJx2LtQ3BLJQbEKoCMNnTpWE8WsCgnwI1lRrFYwjr7TtrTfbICmksEOCR
1SMBX8o4KqWYbMeafYxB3sm//01n4uw20xULuQaK6qc23mw5ZL0v073OfF5m8R+2
6xEkMtahrSwK4fCICX4KxH4jQpx5Ycn/3pjlOxb/FxhXgBPt8jx1GJYaiPyDT31D
owXecCypYQWOtC9gw8ZbOpgIYtdLURV35UXkBFfCQ2veLgRh3nvvrrEHCOFN7SWp
YMI//18PgdA+6aT4V3yKkApnifALV4dJjuzuqoEaZ4TpgOw94ijsvdEzOcUW7eYC
xsMtb6tVHGufR9Rm7/vuGn5ZkwDtKj4lFEu7YWxacfS+sDY3249xZSYZFQ5ZXx9F
U3l0UQvLUYm8ZwXWuV1YRhazYlXp7r6Rs2b+7OmDuXx4RRLEhmHM6a/9ajsyimX4
qz6fbtMlzejGgXc73w6GszH+qgdlWlWvROWhtuMu0CausfW1CJmaukLATEfSQP/I
NgaSC6/cvIDjSfbo9EjGC9w4+XQDJ09fFZIP71T9bSXE0l+OID7xy2H/PRb/Kf/m
7GIGsZs+Fc2nW2e78csuKMt0wqh+t+OjEdDHjFV8sxS9m4JpxEQZiF+PmKYl5QY8
lEMeZsD6lmvSYe7+LhYcHCjiL1ArgFzLRUTA2wQS8+mR3HOovCabnvf7cCKt0ktj
9KKKHf97lEgN0yKLMy/PXVYYonDySBgF+VuttVOXVOXyqc+7HF3aNEZIOYZ69YBX
B5JXtGEh/frzgZkK5c77ZgvkaM9/L4sinVe2QAlwcb9X1cCjpOdfUljj8k5Q7OID
YbFCBeqEY/BF7BYBkh4IOdFVzRcLD4cv6WMIvxMVOTFUtBrjudFSMQRfHslWVyPi
qtKS34DBNLw69r1mwpdrVcVvtaADL6weh+YPP3XH5NgBqlgbPCrVij+lFeVMMlly
9xaZPJVHYzKApYsjzJeomAZ+muMp7I3J/+AGZuOPR/GeLhxHxmldODz+S2bnO48f
vQQdfOvjGDhu2xXGr1MjzIbqF+jjkbMhMza0hJ5SkWq2oHf8vO5oST2Swp59Z4oy
sMtF1wsAc/q4UaRE/MhDPfChb7nPbIOR8s/S6B3iBt/5IyLPmekU5u88HzVgZ3Iz
CN/sEDgEq8hlLXW2RSGIWgM64O/Y5kF5OvPUNlt/mV77xzlo33zPZBZKxNDhGv9R
jIT++4AAnwYYdawyWaCo6XEDrZyceO9xSsG5KEPf0lZM4Yv552T7xd/9qCWTFxlt
C6c1j7PxG41vhz0tMIleLKGNgjU1Qg0fCTuNx1OjI3v3CqE/LYgwRQURQCu/pMYU
75WkC9Vmr0rMTmV1MIm/UiABvoPdkpemFvyXbkierCOYFWmme65qdc0/zejbZDc8
a6w+Dx8JJMWhmvYNerzSFb4Dd9Xq+2wSbG1G79rsRaLMHIzIbrBOOBCI89oeZTHe
GRajLeEi2Qr3d528n+nlVnaXI8FHZb/WZUSMvpowhMMq8WBwF4Tp/+ga2h1YdASu
zfpfV4vNAloQn90HlK/EaGB6r60mOaiX0OblI6uTfFCug3wcYD8hE7vf4wJJmcRU
RzbB9A0Vl9q3dkcgRJtbkZ7A8jQ+4plXfR+a/eaUV+Zs7UZOFCAxB9qvoqCreust
UlkAHd6uFD6isunLhAGLRRijFuOmGNlTsewSO65DVsvkwUd4xSA2Y3+zIPnt65Dn
MYRnPjQD+uLIgoKuohRXltp7lPeqnUDAj6QsMo0k64G5meM/h+oTXK3vBzgAoYQS
wGh1Iqyh5lv6sLb5HZUggzrEEX+2z1qdLUiEj7yuVZMNsUTGZ0vc12P02Hn/ae73
ngYhZ52biw5fgvW5Bn/Bhre4nd2BxVGEfFw7Xu4MgSf5Z5MfiPZcRLL+Fv/geQrq
2jamo491uI7LJC/FzAHzDTrq8agxFhxiZD7+MY17o6kxAnyIQmZdw8i1poHamwSK
KW93+bVEzbyCl4SbppGzpbNOhTKrEDfEEI2FeCNN6FVcXQIKFKWChBk6BZq38Y3y
Cxpct7pSIL5M5JGVX7jE9DT1pjOinRO4WMRkqg+d04rdiJggRv3jsqqccpZCmt1D
teZocaEQ8PkQL+KEVraBlc9SOtmtn0Ut3iiwQmTyv3uC4a9t/QTLI3apcsLeuv9X
qEZQUxXmxevqbKto5T06BANs+nVD/7v/weBwiZnidl+OcaB/5j00Lw+ok3lPbnNx
vyiadme3SLrD1CS1T9TWatwwldlthDEMQ/ZpVKAQKOTx09sYEM/JRZFJn1bSfAEc
3t6Vn2tlgzWKgJPc9f5tZPVIfMNp2YeOZlk7TPAXjewUn6Z7Ik9gRCxwYvULEACN
OpQoKBwbsUdFjUZmPGw5ZkFVaGXUhb6SKKKX6hbxnjwQLjOKCl5nrIRLgpNrnKdb
jHm132+ivLAQfuR0BgW+Lpj4HzXCQTIohsse/FHEJTX8j0Jmi2wpdEV3vAts1dLb
IWSljxQCRb0nEeW6bdLOALxnMM+JQYNEC6+rMHaaNZPGdS5wHhM+QVZ73mbLKTB3
XIRkYZlmV/+Q7OzFxq9G/FLQ2CfiBttsDWVSCVCtgc3Gknp/lJyKpyeMLIZcUalL
vpQzoESE84KWtl9x3uWE+TMdp7D+XaEfjgYhyt/B7D/jxoLSJyfB3fiNhhkl5vOU
n88LZuvBHcJdkY8jyHOZ2Eo4Gkb+XekjbMPc71bz/QIRSMcrVkIKSoPhJx7Ibcvy
nbJCLm5EfJAeoX7cJ6Zd31UBEXASa6hNeMuiZXt+A7tUMVoPT3/GwkJbOKLnDDdY
JAxL5Y0w70VGapcWfVKw38X6pboAzWrALRk78eXeWBQ/W2AitfeqbS1ZNfAQ8S4i
niHKwjoicW74aHBlWg4uRZztfGBOwbC8snnjhcGWL1hWl90Ou+0w2qvIhQu99I8Q
BJtpkAe+f0UgEAIHRQbGoS/4yIHUj34+BzhsIIA0LafZk8sBdYR5od8HEmtr0MMe
Zof1uHgC9szFofBHqilg+Vls4c0Nk3yT3p7mVi4sLks/5zY8sZmdrN1uLeVfOdsr
1I/a832FRKw2R4M/G44ht9DUWU6myjWol4ZqwrKE+IBbllR257NHqLG4fp69oW+r
oC5VERu3lqLKMbd8KTGMqL1SQiqXeUSuoDuXmRNlPPI4WMGFSXdr8WZPns/wRekc
kZ9NOn+U5HJu6qK9/6cFpBBXYXgnchfXKDTqZGP5drzDEt5GtGRl61paRrq4/53f
gf5U+aMJfMxXJnb/a/io675M+RIdIC8s5jAy8x+zWKpespsaRWnnQfrB6WSJ4Pkd
GM7vz8yueJNPeXj18NszdlpNdxfGxsxhbkOw3I1w4XLdE1WtY2PXb4OV0qKiHcAm
cswDk6hGxPE+r9cI5gUxOGQ6SyvhYf22DiCnmeI98klKau0fRZd4/Cfk43vZB6wu
ljQdb8zV7jytZL7e+1jjrnlxHQXtSDZg+tHJNFu9K6mP7Zi1RA4RMEx1w6wh0IYs
1DWC5QceSfCnUMtahCJxljFTXruAnlTrdettuOZ+9qjMMWhoZzXV33OrITzifAtM
9Tkx5fJh1qybID7PV+laNXcaUj6VIHWgvrYJRdX5kE/uttBlTjkjkGlkIcPNtexu
3A/NLXbLi9Ad8n6S4zCd/bjQG62+T5n3n+UX66lmoTZlyVcRs/R/1PMruLxDqwJj
50CywzvEoIcp3HLYCyx96RKBzA7oXYIBokg5JpG0BsjrNIW49YF81qZSNiw7VHqc
qv+BYzG92HW3WZCOfMCPQu6FCx/YU4X3c5k+ApG0ECvBTKZR04gKJ32O2aRXnL0z
/y9TTXVn0gOnZs9EV23X43pcBbvfac98b6B8gZp+IkoxoQSsGUzYnP3sCjgQqmZ7
ZyVtGKv8P8XCnVlqPbYjuDgyAmtRmHa3sdEbgFVZh9o4Cu62xajVwHC4xpQYwVKs
8MBjIvQnS267pa480QiBfohw9fims2Iw69jp3Ov/U2Gjf6qI6fE8dTuuVkhpJAih
XIq2EYHHEkeVPfolFU0j7pr600wbF4FQk/VYhsXvfbsHDFt2ShqIhgYBcMeapc88
w2i3PHcYyfzKXuwq2q7jKQgRpGCo3c8TsgLJ9Atxzct4MLCFvR3CM5HXptBC3vwt
BWMD5Yjq+9UXHqg8yyJkdECU72DZsaPYQxGyiU547spDh7E1D8Z73kd83LNLEC9N
SOx7+dP+1BZEZQ3p/9V/mRTYRA8Vm1EP8ZrfGt8Kj6QAYb9oo6qVpZW8jncawKwt
KlHV+vFMkCyciq5O/Q1IJffoWOxJqgAGF2me0PHqifWoQH9japrAVzZv4rklS+/r
BoSifsJM51zBMUP8huQ+jIyTRcty9k5pQKlhI6ru6NmkoZUWqOt1HlOig+Er2pas
seNhGoUgzCURIEG4728uvhfEVCxwlQzzaOmNuMXqEC5Au27JSNiZXP26T8jjH4qx
EmGOnP20YR0P/hkwa1WYFqHP6g2d+OTGvG5sJQoQPe2OBz90aXsZ5e8XhnkeqAb0
JFh5butmVM++u8pJnXr/8+Qw5ukB2113fUEOmzSknq8Ray3kfcVE2enlJiX+bFlr
8wqaTJiqsur4aEn21iD3RudxRGty9kYn0ncZaZXw1H9Zdo5nR/w0PVcIW8iGCoEH
G1p19PcRy6vH0CXspNE2jBziL9PZIdxTUIzQlDTTZ1OMXdCTUn9huOHqrKDXaxsO
+wAn5BpWC3iSOXwPlBFTqXlNaSUe3gY44POoQmahJFhpzidZeNVMQgBXD5AcZE3X
0xUxUKSCnxa38GfDHqRLmV+8APJjWGYcTj43EAy1DkrtVeI9z9LNPXX1OnPBgGW9
gg3SdxflHTam1zmLn3zdGQlC8iiQan/WKQL5WgpNN2RojSpwlkHwoeIJ5D6TE4FH
poWPZyo59Os97jic0LoCzEJJulNPzDgA7oMq+h5lwN1ywztZsp6hn6mIx9bXUyIS
mt4FW2/671in6C0wBWctB1ATMYnQE8sh65UMNv1tyLN/U/v67dmVALFegznkVNhJ
EBuP8tSMVqpNNTgCGueJIY2+WUo+vc5/2QKS58zMEJU/HPOFR81XCVkRgd+PuE5L
ddgk2B0Gb0ttRiW10XNJ76Crj6lG4TfO+CAgvynnBKl6hYd/abJ4aDE0jAQkCBvq
V6XjA+ASIvnzS/XIZ/zxf+2SzislVORadzuFxoo/T+FHeQgTDNoZK3D9LA4IRHNA
lNmgzaqf4GInLBNGqleSJB8MCrdx2HHOlrxLcLk9tGUkMaQsi4zX9dxOhJMf3dK4
m1HT2XW1eQ9Sg0FSXj3pwGsejPvzaFgFyU8dVIqiUT9h/Vl2y0tlD0FMNzzQdP7J
gduvFrrKMj3UyAioMJHovU0ge5BwkAOfRTEFDbrWPJdUx165Cw1zFQPP/OcN/QvY
6+Ag0uHSMvu4XKLTvC4DyADw9DWjcCmaWWh0RBS0r8QBX/4nvqKqu5zsoKGn8RsP
ODyNxyB1JcJ7iVh0iBr03gdJZzFVRzKXWVS4WNgOZ+DM6jSF9JwLTJ8Mn+ctCKpW
wN2TamfKq4VKv3eXjI+qbg2zd6a+XCmz0R7BZH5jXM6UTEbA4vJLScfgHWh7S4KW
S23Ex+kfpVNVbNjbaOp43kY5T4i/ZLXF3PhffzXSeqOZ+ItAVZBkgmSY1kOP9OLm
W61MF/TE6p56TB4Rz7yq/Gwhc0qEZjBR7C7uGnEjirc3tYJHLgXAdvKUZugvDZ5y
hzqNQm+xtaLe7xP4Ys+Bxl4IAtmkUQPcvHxAiX+LOq4+zfSFlum4w0G3OTbD+dNB
Qha3AOmg0vK2CERfqpY0qativ7PZ+7BV2dGUWibmfF+KrbOwol1oEzuSN+5u49ZX
96GoZOTCcVw28FJC+Ej/T4aIFyd+vbXM4/01dxKdl7LEUT3V7Fww6qMb7mvWwvJb
7FPSPFz3lnutfofqXcQYj7AsQDZoGf5l3DqXdgCoHGqYRopPwOyKvgNPtchXKXeZ
79riToEo98iS68/FzLWKWpmn4h4WgbQY+EEq4uSWUbOhLHEJtDQolqLXxSYuTH3o
O/aXeGGYDecIw2+8B9YcgG+CCQBKozSkdmMcq9uCnsvA0TsXiO8rkf2iRuYwUc6j
P4QsLmXjIZVRqJbJWFJ6+JgweNzTN19orxGT6/Rj62at9Ss90iUdFCMhQMx8If5x
tzWAlHC9KO7elYiRwlAuTUVPHcho5BIRZNrOSMXlrQJijIS+LhL/+jLFI0vR4Oni
TdU0UHMv/vb9v1stML7/cp30uFMN1UF6W347xvIpHlZ1IcxQg+a3eLrJXiU82EU6
mlkOjg4VNns/9WEqxaC3jguylb9LqhzNV3b6esa/tHKX40VhkrOtJ8cKCxyXA+bB
StOroi/cMeYZKvK5f8H1lLdLc7tmoiLtbD7FU0IDoiKysz7UYzmxjNMfXIXRc7se
rSQzodn2cyZzDc3TYpd/zIuFVo3fJ+OxsNkd4DPvJ/imZRQjTlrkM5kDkgXWUjA7
unQNFGTiXgNKJdm+SwlOqUO6ZF6sZP8pVkbwXHYbwsXzb9ivA7xAA3S9y/v+QH8k
8LxjMKsuYJ4L+fzvdzjXzUN3yHjhBq4ekHQRMzzRcy6VPqsn6qbGvi9BS1X3oQ7G
Kb/ro1pjJB7oMsQPPPhP9T3ixia8CsxOFswyBAheL+t0oTfwkQ4yPHhBOy3C//qq
aqaVjDPcU4aCZAMh6gSzponJaOsb01iTPt0ck++74Puwp2vVpyuSb08FQN9jkySy
hFmKZ6LvTKM4c9fsEsogLmOiqSZiS60vCFe0acsjLpCDuZIoSDOaJ571SmUE+Q/5
+EAbXkNucAIPOy0TCFVU2LBupw9oOvpac3F4QTbU1wh/Wv06ekDgnvcLdjAB4Nr9
oVuoQEpxgBRpoSI1jpYR5ABOsZkOG7eZng8ZRPhut4R7CQW7+H8lYIvJQpGlzyyj
e+/YjesemqAO0feNiHU3zn271++0fDa9cYAY1BJ/d5/grKCjgP8YI4bYglSCKgZT
gdQnY8pQQyistiWEldQ+eAP01OsUqRI6tEhnxR8skRpd+22Yiu/jVIpgrm/lfqXW
5gPgbnRcA5QSXBiV7ptZVEIYpj+1m3OAxhEP0D9Sn6H65iHR90CEpJJ82fvB9yz/
W2fwsjufiMXpgYCvrXCweGSUXcZEoNLeiYRFx8MTg8S2SFK7OwRJRKRPYE7ZfFGl
wGmwmo1qouNI6mUZ2aHNtZqWCHllMmbElgvF6uk5ZilT+OTF2wD7MAETKOWLwa+X
+Njg2pqgCdnCcLrgMrxbFh1GFEyxrRTkD2vSMBt7lGApnt060mU79f2Ui0gORf4v
Ilo6CukRJ82vunpXQ9BrJ03+ah8RMsOy4AaXbzwCl+r17fPAVQHtfAng/AnSKMjO
wimFzdFOQhe9L4eZOcZLVpI57l+8Xu6jsZ8RzLQBhhWf91K5peU/vstyFpX0EUg1
54ukKFD31Cdo4uTElwlb4HVbmv8b3ac5Z1XkxUyI15wf7weR2j60/n8+aOWaH16k
952UWZZrpCTJo7tJTeM2zERl/elyGwSMch3/b4ahr/fpcQN9gkIfTZuz3m1SjiOA
kcJFt5OhTpdmF2RBdVykuWdEiHxjOeUbqOzpTkGbAlIFI1xZoU/NmGe8fScFzbkI
T3KyktxHwqIMGW/yY4QNrzN2i0UqlRh1N5ODPekRaZwYQNe6euo7Vk7w7zwN3nRp
DLcmOyc/e14Nl2QITaKAIUgQ54R0IhY0HrZNxGLabtU/vOGXzJYQoJAa7jCWgZC/
ex21zIoQwEbykpfmNs2e0VkKUtuBpvhBVxf29lcsrg8txsuAZsqhY5tkCXHGazkF
tlGwOQT/j8pGPgh3L8AqsDleSX4vMWmurEdecqx1qXDUsJvoB/t3RdTTAeBoEjGH
LQXvwABoaNC9S5g/hmS7DYZLK1pvRQoA34GTySI4YamdubNvE3sx6QJdGHn3s+0s
qwokJ616NjiAfMQ25icpMYRI/h4r5XTCX5avrYLlfcH3yDpqnTOKfeF6XhoVm6NB
McV7LJpgKFVwqOjNl3GJL13xn+HIZBwJK0G6C//0RvOzNhMDFV2XuFVyM7S3g0MO
MSSYwXkuJZ5WEFTZ7b/aKu+nC5fR/o1nB0hpYCfNyg8z2jLhSXlhHUmi33r+zDU3
+Wxsfnf7KDh9/u6kJm0/MbZSQshdgLduZPfRC06AAVJ0B32iXsxgrp32VSlKcOy/
UwN/MCqlJa7ui/ZyxgbhFMv214p+NEWRCSTze3ns0uSgqve2HOnsmBQgX9UWAORg
kuDXARCtro3y1hrXxmyU+el41PGLn2+ZkfIAKM1Hmgd5yonjsHHMcHncNimJNAKh
tXg49mbIWkZXa6YIIc/463Uih1Ptsrg7BKjdsa1M1arTrCvvTpMqOxwA4PDJPRbF
QuEj8zX0rbX668h8MzSBd51mJ1SsXyuWVtKcZl0H1Sd3DY0RR4oBcH9fmZY0doFY
YFdWI+XLz7dfK44bLGr371OMQbmidFnBYR4xmb8l4sX3pR1nJf+xWQYzuHeze7W7
0/Vm4HDmHMVzurR32ne1yllb6ako/PAbjU7nHpCSutbu/omtjD4KqzGMrFEM85zH
le5wi6WqiQFdGW6zKPhOMfn3Wkux0Rk1LNWXJNzXlhn+u04nIIvyiL2A6ywYVLPj
SwRIRdZjprMQeBlOZvMPSpOgLW7XmXP3XxcshrovC1a+vOJKdRQd4Cr2Sh/qzbcH
9rnZ75Ar565CJKIBgYaIq6tGLIozMimdgvPlilERLmmcaqSrWjZrmJVbi1mM1SAu
Lb3NLJlDCES78ML2RNLwoylQc5mE/cpO+9C8gnNzlSpBBEWAIgEAedIaQx8CAX9R
m8JLK1x/2RZjLx1RV9eK4pJo6fKAM998DEcgCCFkPJUqqecSAJdsQ7rOJlYg4Xhy
TMjfgQuqrTdfycZ9Uqop85qjNlvM5Whd+osbtYlX+ndYgRI235bj/xglDqzXc/g1
gG3MC5V75CmExtOPkOSyQBmwNyn4C/XeSl6Y8K3+JL1MugcVUZYHpmod12ASuvNp
pwFhNQfR3/VvEIAePKUSVc+78nwQB9Uei9sLaTc5hxcVISUtTi3Kj25lnyPI+10d
/oeit53zc5I0ubB5+4YsfWQzOiMplcr/sKm2C2/WzZAo2rMZPog6tOtM72KVrBRf
lGCiuo5Bv13W0daB3X4vG7S786dyFck0YE0ybW18knjadhOKzMmYGH97rSz3EdgW
3e1Qmk5f1RzyXJdDsXQvfXbUPeBlJ1VDJHoW7IiFfQ+oMMphPraYlqTYAb4QGara
+QDap0hKaLuUH/dQzL3MtZUxvikCT5QBR4DtRqNbd18AhdEgHYvnNVg79Yae8R4X
0MVDH3cWbkCuR9PGJPk5+4mgQaAzgPXwJ+bUmLfoM4ADkh40u7y/GNWsi4OhJshT
hv4HqHfyWQjXzj79ifMe7vlsao2x+oFEOnqRvfUaKJ5bSQ1e5bUqO/kkoVqJJEtr
XoIVrsOgXm4mmpc6vi1pOwwfwmMXHBaJ4reHWhs+MyKsSwPRs8vsrTNcZIttYL9w
OPFTZD5NDz5wywD5JfG0sgN0n/Ihaet/6JPmeMgPVtbTqoZNTk4O4b2Wmvs8QO5Z
j4cxlpx1obW3XJVy7eXbydMwlSSgFWabQ1iJW3eyPXe7JxjLkuYj1fEjPQg72IoP
FE6wrjpfF/QE6a2xWkJtcsP+MkePJYorx9HvU+M7s1rW+BX+WXyDs/ZjzjE1QKHu
e/l2SnRe0yKS52mqdT+swKhv8BEd7LiTJgbeIqg6ZWaWvIynFpNExuI1Dj+UV43O
PftyY+9CLpLTp9S4qQS51PYmROKAGotPg9YR96iUxiQ6ep8yi7aGKv9Ia8GK8v3k
+t+dw019/Rd11gbH8C4h+vRxHyqiBs1alMJ1Nqkw2t0pBxJx4LzuW2Aog9lv4Wa3
/hmWkuy5bmv93YNe7dLX/ObsqzZDu9inMlUsQn5qjhBANUytJ9GiSX3LuI3bvNmM
yWzxZb35sFxLcOIP/1ayc/758PNZ2NBago3xzeJWQaN4SHvr7erK465M+lAC/nYS
LMCNSsjECTu/BJjDBEHFVCwvpTfENcMnlKTrILafPy82ohbn1n4O4hpScDBcvji4
uiw4AHVsTWrEgKJSdZ/+MqtSBx5GZuH0ucJmW+VhSuMZlvlO+ZtPhhJuYCS/9twS
IqDVt3bPdG/WAb1hhtQl+wdUyI2aFiCQNzNC1F+AxGGRQ+4QwLbEWHDxWz0azPpc
qmm4OG6ip0CFI4QxGvAOr08HOPYuOnVkJM5A8nftMoPFzZECRSIGjgkHE6C2oX39
I0mf4rgn4ErjBzdi6aMlRyCnXWdjIjN7Fzye90jyDLVscywoGnXhkmoXcYb0T8/y
oAfoaJTz6lM5UEjRRZIQ52zlknqZmOb2swOk0ci7uHla8eHuP5zWXzZ3FmMUsz9x
QQC+KSUGADRbvT13Yp3PlVnaUxix6/qDIAc89UssDORyEkfDV86ZB3HAx82VvT3E
pbNaXt8ZnG4z7YIhzE05l30VQ6OnN10OFm+n+H1r7Ya7FuEFogMp9Lc5ixGYu+6T
qP6NGinPAvqH5umfDj1k8IVfSMhmxRg6dOCrBGTuYabV7BIi8DaD8NRN66erPvHw
7auM3GwNMDz7Sh8CjNYpyfgw3Ul/waPcXIw3Yx/CQx5Zntjrghbmi3JZK4IIN7oM
ANqVMYlv4q/jPtJs/Pg27YObPuhHxctjQV84HsRZF5TKX6ie7LcLsV9cR88ZF4qD
z/H6O6xkKomseYyt/dmRSP8M9gEQLYHe0XzO43f0ugwDaRbobedNYG6X1OieT2EU
WsxOHWO14JOiox8gkkxbPPQ3z9FkdeL4PmRcgnHDHJW+WMGev9LEWm8J1p6GjLN7
siphEeJ8sV+z47R/ZVzltp4dk0vUjPirqSf3IjLZnvkjG163KGM43LzO2qAKG7Fs
0yPRqFWn6wTRC3XeYSl/Wmu8+50yaZqbnZwoD/RG3GJmT6T9gQjvqwTPwpsAm3aB
IZmxUkSFZIj6D5+g/GXoWO4XrLmTjj4Ke+2+2ImiqNhYk/zssTLRVXQePolr12kj
wGYMYmz5aXMKWdwy6ZHilxFDI4T++uBstCw95tTfp/hjQOlzznQoMRyf4jpyFpAY
XwzvOrpR7IdNJ+iXLkMfc6hoW4E3H+10oP2DW/z9mXdrJxww+Ol0AFbpWaCtGPxW
dwJgBVCnOhT9uXvx1feP3a67rTx/J9/yJwV78ZV4qG8PmXRFEf99n8AyI/V2Urbn
YH3FtTw5z1IrUI4yQfbaI2YQf84PwiY1Zf+pwr8GeEAJh+7GAdGqYtKgsjwDc4SB
cyBKh72DEkPr1rUNY9rswVShNsFq6dUL6z0pzEhAiwKMOAA2sDNxUAAhoPY5GB0P
NKW4rH12iz0fkpLsHBIo4fmrjxOg8qBvWJTYoIyvQB8WbZ4Ti/N6KJtxkIkSs/zD
JkLefd+EMSwDbSNA2XsQqOVJcQFDIoLFtkpJXNbJjtWaxrSmX3SHzoAF0TtFNIDj
93P4C7CCG8rXi5NNiUohZghg6U6KfoJj9Fl+ElsQRdjMmOjAUaCwgFTh472ia0WZ
kkI6bsRsRuYUpoCe/XCaLbYM42C13YfMvPIr1YePWc2R27lOUxnIjeA2AhRI150O
W4PM+thr69JjgZRrN3d3Pra9CFD7UKqUXISnfCYMPfBGAWCabF/dOrcA1Y3pvkB2
g54QGMSdvWaK9xTAaY/0kcw3sN5F34JEuJKTPvQKwjY4tfM0ybRie+rXMgQhAebA
7PfOq4ipDJa/FbuEei5IxJtg0wZcc5igOujMoGqYfOeUQcHBOU+zzDEIW1eK6F/x
ozHeD9lSF6dIrzfaUskKjR0Wg5TOEJjgM/KgVnIfMbj4m+pKxYMIqNWGw1uWcLbX
KzXsMD1pkBOcjMyOfe8n2CbNnH7UE91+m+HFHIkxrd6og5U0ftnmsKHBjgHIyPqT
1qBkpv76hEVqDzX7WN39Pp7RnleQy199uG9McA795D1KHFhRzWRmlI6loWSQji6y
2+k8eXLbXpriUoI/6rAZ6KXwjsrqSFoGG3Jgi+r3Bq3Sfs1iIuAfGodzm07/co2S
CRw37ahgv6VO4TK/7wZpgIkXIJ8Tij/K+ru+qh3bw4iNlj7MpNUTFwDVdbAJ31vG
EcP+Y7JzQ/HmS6DVKG8tBX1opu92cRIVKnsu+FSyY7Ujv98H0NhjZTv+S2AQDe9y
7DeAa+QBAFlHCs0V1ntOQOsstoikAdyaKbuyqt7k4A4ZHy3hqs2K7TC8i2Kwlc4s
YegTOAjRRLs8IImSyy7WWvpriD4zOoBlXtSX057esILPKK5ZVjXyf5NOQuVeleQC
bYQI2nJrHutKpbRfT28Gxcb4j1ndFC64QKF+lZY9hH5UDIE6zD6Rs04GNp5k1syr
Cpl4EFmayC4ecu1fiolLZSzGKrRRLfnwipAP1+ZaAZDG1ocxznVAbYCjLoiiuCfv
zIqlRRgXAurxzzjhTpRUpOahNDUZMS5Gu4/vpg41W/sH8TU/8E/FYlTShk9NZECi
EbtmjSow/WaXjZsvGUW+zC1EBaaH/9CPb51mwiJNno+Fch8iUWPP6+1QpTQK0qA/
Xfcw7EVvxibCt1H7h9jg69c7+DY9PYfBRaeLswQ1ueAlRE+EvNydtD4FfHpya7U/
xmEMFQtLrMl902yV4+u/AYLRJdoDfCH/xgX3K7fLryFu2DgDoW9d97QHHVRe6NSF
2QAh+xaoxN6sE3dxrLuecrqUoFu2DydCDMazrVHmIMtGST2Ac3C/fFcvt9qDOAeZ
AgwUChMRFIzDFqTDGr0YpqfYeW7VVAexY0bz1vyF/jAlyf80Ay+HZ4E2HDk9ewyI
f9gL7U+YK3m5BmTvJTrmNvMMDGmLJNdgzC3Vkp8HrejSvuNRutrPwDIlfGOi3wKV
rokbiBAdsihKjpYiuEBmIreX6G/IghmWGOrFt93NI+NnkBFwWD1b/h3SIi1ii9kB
bIzeeYaXIGHuXQTN7sRAMOYLUplbe8FqR9NIQ/MRi6TzbfNeJ1j+I6x3H+hliv5t
3xNvYwNhDZ1X4Xl0MI53VQY/v9vIdBnb61Z6vjgJ3VEKaNnwwSVaOWu6PK9vwYnr
P5XFtNyRr8x6upR40lwvxTuqnzyo/T8qkeOtO5sRQdIlYFYOju9BW6e4IQ1CxwpV
ECLEz+rSd4E4YEqjSj1bcdRLc0JdBmEcjWxG668M6UNJiFiqrcJgfl5GEo1gUrdG
zgkNkxYVrEMKtJUcZbq2jda206DD+womcMDMPKM4DYH5gbvt+JfYB1NS4A055aVH
ajpIUkJ0XjC8b9DiKNvXzue2pfDYEI74evpM8myT6VrF+z7RtVECzERKXWgALlFi
MNV92YpsodQ9pQqO0i7yR3qE/1AgOV6lqqWsU9ksbLE/5qQZfBEwj1L/Io0K8l/J
H4Sl08mtx4QYoI1CincID85I7Q7pCQG4wLXJ2GlNel5ohXtfsezaxoaPJ6upfTa0
Xs9mqSf0j5tr7KgvdGAd/Jgd08SMflbFNbh8snJXw21qoZXf4HzSzd5Cb9HagIL4
COS7/pInkHNp7T13aKTW7o93vb8xpVgZgR8/HkcEcYpQLnrx75r74lXH+yVNZ04R
dQtMAYJmpS/qDHhVY0JDVphxEDgQ0XgWGNzQB9yqdQsXI77jRxpCz5CyGJPjzHbe
EtQXvAsHrHnsRxNdk1X50gyejOfMpb5kEXRWhQkD/MbhzexCE29zg0L4UNd+6B1s
W1lkw1LBSHIPmg81n8KZZT89rsI/zCO5p9IBxviNdxHdiY3Ojyn7rdGJFrx1i427
atWeK4X5+hvcufOIYNsib8zBAf8QGMK1Cgtd2MVVip3aIT3xkkAddFwhZrTAB8vb
zE2LCPzgdhDW0f2OhI5ny8ul6iriWRh/SGLYoQo1lS1pnIkkMVYaRmikoRvZpk9c
m9tOaPxtSuTcpH3W7zdLGgFje/UbItQ8dtvriP89zJxHZln308FSUjzFcVSuWcD6
lNh0cEsni4Ur6/hKu4JgQNK9aSkjd+195Xn5VTOb6A89M/n60okiWNiRDWel7K8Z
oq16sA6RHvG+O0ZXY18lwAmGPkhANIny1FHw7Z6fHm4Jb2Y9KuWarXbvF55zHeSO
HnNMAoE1FHoaWfkt09ajyGPy051/+bkagxD6XOXqX341cBOLImfc3ZC3mmXa+e4y
j06h2AXPHCxJ/v5ONd4LUb5cKbsMHiJkJHQyJFE0DutF/f6YniIWG5GGD+n20YaQ
3EN0wuvM4FVusHXzVXGyraT3PPjQq2bOrT7oLCzcWgrwsFHb9EmZr9XNL82txVh+
TJRWdEbYaD0KJIJ7e3v3mNpiHGvYKPLKTxlCYxli4buuHha/HFzvSWZ6d2PZl0rR
PQ2HbmLK4OcxrMgBSGv1LSuiRQNDH2jKXb/ieongccC8yHdajvFUPMUSjVvqc5tG
iOAOkQDfLV06QqZAEwSrQjLaV9q+A3sRqYeP2k2dZcLkTdDCbtiA9mqQV9fRrejl
6eVp+zsxQTYqlw0CgW9oRMFNdGQJ8QFwASzB3RpuxLUKh2qWI5cMF+wg50gHECSe
iK4RiH10LX0jClXHdQRZZahaNtMEx8VfkIq8ZxYBQZqcwEWOM5B90tRXTW68LkVd
XvB4aeIzl5kizw2PVEcQw0IWLzI5C01G3NfF0pmjQo0QBi6WNn7MgTFkcalQg6Rb
dcrKaQxK/kGi/Ra/pBWZf8vxNUaHAjmNgxkgsjo0p5YWS70dSe+EAfgEPMy4JOxj
++lbnYZB1ypOvJaFgI3ti/SQcgrUVw2w3QWHn1xBV9OtjOUlX13hSRbVzDltu8AM
xOViiMWDj8DMPy8KMYJc8dJpu34GcsX4sf66sec+fAk9HN1B9aaWN/3qP7Oz+5Y6
EnIeMAGWtO0O5kemZXdXUi+F+DOrDiqJCcIeUAuMVj1I7SgIPOKhU1nauV6QI43C
XK8A/ibsrVBdjYHsfBigTlzp1sd9qLpBZOIOcbCbFPV+IZrvso9PqIPQDJyT+i4U
Cc4QWGxzkxpSf0KxNt3ENM71bw1uSlqd5Y6c3jvQZWbvTOwUmCFgi5d1u95NCcOt
IzfjsksKhgtCltVU9kSddR/zWGv5yX4WE9fhEAulvPM6vlfI77O+mk9qJYxg9ZoP
cR1gX+3g9SUSldHDVAskrF4bfN4LhCkwYU0irGtT5ngJP4RmiEoWSQ1aE+PDUTbT
hEHu3LWg51oPHXfvIIUincru1aToLgY8VzN/Il2icma9CXAYeCfpy3vO0BcnvzRO
oQM8gDtFLgDTbRDguE/84nNmMneswYOnu58SzDyJVlfTOuiRgXqVTTlay3J2R60a
0/CJb7zGCnckiRG2eXm4xR/lwdGOqn8BISA6FKEVrNm05uOGkHPX+hFf0ev4cQRJ
EMkZOtGpsDCUqE5lDDQdpJc11/ID9HhiEsKCjoIAUa1WRkyoirg1qiUXGQmNRaPF
4UvKiU5TKWl1PQlWneS5hAgFYzmJOjP+xzNyDLRUsDcZMtRgEhUpmsxMSEYZ1Zw2
nc3AixC6rVb9XJ21ADOXiDBeHNGQ2KFfdaVaLWhosSBSjI3ia764e/K7VHZIZI1/
DbQY9DN4FBoRht2hw5jlmmgYS9CBtNVTPBogzjo7SYfaqwF3URMEywUxqj7hOOkC
7A0FUTPBN16FpUUcSCT+99S5cYSGN1L2+QRLaZxuCXyPeOykJS2Aaz1qnavQNc+P
fKKsL44TDFZEc9L1yLu1knInmHsM2DA6gv0ZEBrIyoT37lIxgtC8NPOO2t1sahZT
STkdOvoPTRdDSdO4RCMuMW566ATotfv/9rlRHiT6XXwVbVgV19OTBnkvfPQELfcZ
qZqH+Hd1388Pp7R2oFEpofQGuoKYYwwoPOx70Z66RTqsoLhoJ7S01J0oTTeQ5rXx
8+P8BKMKcNjtGeiXBDDeKgJ9IsQs8maeDnIuNJNeQiGI3J/LMztkRrj0FizTjlrJ
0HkwykEDtuAusmoRpCr8DPrJvg7CiGPN5NmryC1UEoMszGft2uvZeGaX5n4tLSGp
M8dlDCg7d+hrrLr9n/DHa10wOU/nSMqxlnMn+WPBjqnqoJXmdiI+V4dCAOAdQxDZ
bi9P9QqAYcc/kB6Wbk2rDM5DawBXrH8ams/ryM/fnKhpKshdl922lLU/2EXrb+p5
/NJEWr8gbiFmTZvoj4+Xd6SJCH9rbVRFe8QOvqthq4P2uz2hWVKuvl8qBwabYrD4
ABdHm/Zjw2yZxIPJ6VypCiExNZlx6+ogx/35bnBq4LxdmFCM9S3mFUKreLShhisx
KifRT4+7fc7ppCw1kX4hW4BjrqvNmFOyaVkNsbMVqQC/rdPcFIOGAyqTpfRKA0z6
Nn7iJYo55VnSELHC3BIBb3+VvfICWCPB1vkQ3SfbF/1wEFaU8ZHgj9gDR6DN8Gec
jUbJctPdZjwKSlpoFSJW9DPi3xr7Eg2ohgfU5X6GppBA1BLJaJqY+VwP2lJKkTQx
7AtAw1sdGj/Ywtl1RHErN+FQh9e2MH2Tyla+OD0WAwTdXnHPoJrbEuNyDm3u1M9b
WVVC1zrnGRfjiLI4+sXINMHlMS0k9V/tb+p6V0GQy+T+Xyzn/o5aSwa0YwmzE+LZ
1qJ9a1qkEGbbw8ISvTN76maRqCHIkmRIWeBLsDoVRB+PhJVa9BhdNYGM0VZKoyDl
I8u6QIbpH8BOhz+r/8H5v+79EDWD59WLREbr7JEl9st8xoRmSKA/b77wWr2kZdh2
jaV9nicAHXkC+ouOjafW32D65i4cTX5redEeGmZOEruLANw9Vnq+G9q1Bt3CRJMo
M+eP8Id3LYACMxtSJa8xDWDWcaK2nfWwKUFHUXe9JKShMslFRcExD7Cfb5KGsD8O
vPfe8JAk1QXC8VThQwGaPPJgbEybPEgv5JTOT4lnxA1l6cu8vFwU48Z9nw6VqHs8
fMSX6yL3H7mhoNLMpQWWKfRE+Za3zi7LEfyb1pR3uP90+6QOnDgBRokQHLaV0BvG
VwdbHtt0HHTyObeQp1ltoT8G0TyoOaJRZOnTPRUwRaIlOv0Sx/xDqO8GO+C+FPbj
UTR+ao7mL5oSW/bMx24+GiQDpueBc0oBM3P8AsDRetU3qcvxBKZ/lJiSPYfmhEAy
JLjRhvSz9aVY4JC0I1nyiDx/goS7qH5lLUXcpPDiCUwRDLB7GfwFmnxBQkkaV0ft
TJ0dyMuZV+tmrdHMuoj1a0a6Edi3YOM61B6T3vxWgqGNcXKVYwh3/D4WFBFrLVI/
Ij2q1cnPWLBrJZaGX/v1BKnxfxgvcs5RhqLomP1ZxaekOuuKDmruFUHdGvtDcHzC
iwAl7dIHK0oAhVDi7MGW7oJP26ohNCkdWBdtAqzNB1C8fhQAhPeOkN0Nnc3Yrg4i
VjcxY++S0OJfsYUmTXmQVBB+L7wg5u6RdwCFWOiodJJHLXdCzRzDYTyKBLgvTlSA
E2kx53c1gN/e0dainbyiSBVRQ3UyN1dvaG3mOjgXIRCDHX3UpoczOaOoFWwUAoie
Yfa8HI6itqtzQAN0HoU5tE03ICTQkywiPsPO/lkCqOHu8Y2EERruj30XfiWEUHEP
sHf7uupAfBc6P8b+PyxVtWl4XkxK4bxNnKNo1JT8D0Mlaw4/VA4I3bZ/BniGefpP
NIysn80UPkKcSCmhVW3Mf43z8AvDlXuVjwqTHI5P814MwB8tjA966nv3pV9gniZc
XOZKyZQHEKkNRwR565EBXh1i6usS6U9oEPJVkRLIrrMeYDdhqZjlZnF0Wy6vhb6i
NJA9rVUH26rkXGp3AaiKMDSYT10hkr0nlfvygHJaOI6/NDuY54b+IN6pd3Ue427n
gcbjyd3yTry8ECA95xG3rVxRxynQuiUKkgrrmwV+VltZ0WlqKO5yCFbPEQLBqMGw
KlutZ7Gmx/IAuM81Ql085a8XgT+VX7/CrLfzdIl9ep0smAwYagSHOzzQuqat/nr0
peIpa7e0FAndW9uQMQSXVGUv/uID68phwEh8t25pr1HrscxyvNB5Vexf6BA645zY
R09OtTc0C7D13n18rUF7WLicJ1vY+WtgCVBcLlYgMAXfDfaXJD6yPJ/4UjW8efOR
9eLf5q9Bqe/a0uN4FnQuBzgo0zDts2u9Uzu6DwJeRaoUwezQeoyqBjYIclx0Bvoo
zFfYG37AfZEwxWtf34w4IbthhCo2MtFVQ8Uqo91haYAXnkvxnk9txDAYLmtGY/T4
ZEdibKjrgH7DcZFqO3Rui1zIKwFMfMHi53V9R/iX+mQoRmImqpTu+isjXHBIAZ1p
UJdaCRsVhzBCr/oI/hxbi/g1oKxtDCx+avfX9yHdQvPJDFbc7wPTd2+zfp0nKQFp
8W0KTmgjYPfBt8fZAFnaO7IyNEcKnx+/LH/4/ibPgWn47m7FsynYqVDdhJw6Thk5
v03uXni1bMix4dDHcecoPjk0wlLv93/iwNgnQ8RjLPODS0wrvENMtxyUqekhYCut
cB3tLmIZz5we+2GoLfmQ12yAwCyjdD0l/SuKmQ2DsTKIPeyvKr1Qcafy4kaErqxb
vFXbf8ie8bjMfB15kwty5H002bpU7sUUed2QLuZyJ531MrZlKw4xIgGsgeJCqoQ4
hSUjB1vgxQ6JUJjuTwzR93A5EQW09bNWuw6l8qtZOyRTG2IoUljParKRAY0/95Zf
tVR3CF/qYpYFTxXeQxFGbfLZQMD3jDhlUoTVq8jduS2+qS8MrqOX8hraCpy8p044
qXn8x8mjUexJrgAWygCoA/4VPtb2YLkDKHJ4LRZGwqehD2Y2CG1WivPiwGIY4neC
TBJZtCemFuE/U4we6tSjhBP5MmD9HL0bJ5OHDtd7pYF9M57KoD9xko/l+xKMIY4b
wW/e286FEZKuABvt9KwGw3v6PTWsGWaxCBvAT6q++aPxaJVKjiZQTzLmcsV9IkEt
nFYlzG0cmwWe/7ZGUV+Y075/ZegYnkYD9YBQaw8MMiCEqRBRFG2ejxgwY2gXsNYI
YDj68IRvA/ZjXrlkqZE3ZoVd0AFazAjKfIVCSB3hWuwJanAhbDS3i+v5YkCZb9Cq
Jr7T8mAGJ21BSQueSSJmik2i1osGfcuNOB8rpbzxGU1bOuZ+9qcZEjVV84ZCSXPZ
vWANPPAuK7n4PL2VuyuIbkV4qJAY2IhaUZYlaoiFkLUzp6RIiMk6mzX7obzjl0BP
PjtKMq49yby3s7jvSCg/YUqUE8WSnZRwyLOJz+sKk/Zotyr96TB9dyAJ4Wq7w9hk
99AhHQ8WEAvncD+OIZnbDcjXYInW67MiAPQNyULs2SJ7+28nU+CMHqDs17wc3Wbj
GUsM8W21Bkoz1ozFKqowmOjBQEEchAYw9RHJKDPSC7mo+P3/gUBN5l+oEqCeqI4+
7HrLRJnPRHplb1G8xwnT6FM5FMPlJJ3ztzgKMIsl1YXYuJIGia3FRma39RklOJzd
xbjsQCSd8FA2nSjyUp8BKxl6dp0E4TLtOrP4b5iUnmI8tqLmgiHYRootTz9mnrPT
+iRqrGTLXIHbHWroVIDSP+YHA97le1GGfBBOlY1SyE6ms7ZshXPGzU4A/1jaT2qQ
6/so88QVQ+2ahoygtuUqigV6tA4Jsd1O0BDOWQBjd8L0lp0Z+dJlrzINofYbOgsx
26oe3F9jh0luYjjksvnDmXutR0qwkD4rUWnq4SkbqekNB8xdAGaiHF61wAdhgUI+
VXgRWZ7COEC0Ymd0zEC4on6cVnfKEi0G/qBskF0TNpIXMWQSVjv7kOuuR5SyU4Wx
E04e527xQgiVamFLaNRZbNUnKeSFrg4GrfB4jdgBu/QmWrfINmSvDoSMKiQ/tJgz
v98LO7FZixn/fJMMYCMQ+fJ3ynQG8m58W9N1M5DND3YnxUw6TZNjcNz4N0SK1jF0
Em7mDtE4vKemwj52eUO0irQXmDN+bzo3yr5NzPZ3hJ6wA6yfoSJhuFRYwcCtwxrY
aCS7scHH9P16fewCMI9SCXtRcIHF4LaMoKO3xhpO4ORxxaH6kVaj23H/i+6AAjcC
01hVKflV3i5gHV+31Xo2Ihucn79ncZ+hHcUYkE4Om/ls+heS7umoBwKWMNdCcETU
TCfMJdCWdZV7yyCTrPL61zTLDE3HmGXEqbEsouzzT8eKDp5f8N8jiPu151UnOiM0
5cIKMLP4zCPxLSDfBgIKmTKHyEX0AfUbmbgfUZuBuRsfz2PkNGdwGqu7B9J2In4n
NimALXqUjsK2pHaanopZgdL7uxOJVYNxnrYLZQ0Yy9fIwmeG4ms2beDI9Eo9P5Fs
AlNfoAZB3fODxyRiTVfbaZmPCQ8XgDsERQ90VPG37/G85ThHeKngo0nagj2xQVhX
eDnvY5rcORxivdpBUi7qsm7mkMUVD9179ivATiSIKmLuN0PfQZxDx6ctG4rquFTj
1ouQdBlA5WY+Sj8pO3+KyjdXrirmGc58LXKHlJ+V4VaxqgklxdUJQPFUPG5GY3DK
Q7PmFGTeuBL3s/EJYh7OXJXfWgAH9ejQ1WSmVLBlr25DJuSkArlJ7CPuLqdjRRZk
1uNXAf6eer7jnGcKVmTGWrqzvb1i3upMkrlk4dAwmxeO44HBcysTVhTIChRcutus
nr98tpjy7NVxt9+fQJas7r5JCLjZA9LovfGtcE92n3yJp74lDz8WTgJlQ/y7er4F
BEZp3yOX2j3yi74kzHRJZiU5wFNyTb3lGo0e/U6HBzK0B1Va8qrT3Ef4FVI3vxrT
2oUdfxDVYbL4UxO1e4uyLccxSYjWJVeKaViHLZnErOuSr8PSGQqZT8ADhnyzmIr1
KszS4N2lYvBSxhF3ajm7Cy5l6X7sQ/kk/bNp9sUAYn/7vUcS1pRVbVniA7tMS7vf
BZ2L7XITtXlYgMrHQip1PQ0ZeSvO6cXGDoBMJw6ztbA+v90C2zMi2z7OMxcGP0q4
ZsmeY9kdmmSBv/cjA9a2mYIN5Q2cXcUyS/CtUe8I65EVmfx0mC76Tr1iabZFhV6P
Q31gwyQNdvh1wgPMFwWw70KDScPwVUtmzT0p6Qdkvormyqm2xuk0fXEULHGIOTa0
ZJkf8S2oVqqgQcEY/xLCRMA1/xJ4Iu3UHAp87BZ1IJav+ne+A4zEaGbXAUs+Qjs/
7T4oqoxN0l+hif/GlRAtERTIjCSRe0JQZ1AOhDeRW4EQjNqor/XbhR7DX90o2pD4
ydEI+NUpGJ0kC7PKmPfxJrWIYumA0rTQfeF0Q9OyTKTL7uUZnMLSQ9B+tUuKB9Gw
jmosnn94eMiuSDUbmbRJ8GpMs8wIr3p58oPcBK395Am3FimRO/znvWFmEvaYK1p8
DBsXkkXf6a33KM+7l6ei+HiuClkmN8XIrJsLpeWAIrolcu3rBNQRebOZhvjNhobA
MxXFSulP1709obf1c7DaRXFjelGAGFW4q78CnVn81vNdpd6K+IBsWXBWricKkebe
cEcCZOSfPOR2u8RxBubk9Fxt8qGEAv+9GPoXr6KyRhnZDq+5kdQv9m6c4Np2yULI
VeVlBY+dx7jNd6QkoCtYcm2JF4Y2NQAOze+dRPQNxte+Nije9H0JgLBGr91bRISo
CsvGljmJadLr892Crkr8bdMeNigL9xdtuDvCqS4ROqDacVGzQxnMKowJU5I8H/v2
DUt1CFJWVVjrRG18Ai5Fcelwr3DqWZJUmDPSqglS9oeU28+9h2hMkKNlLGL/m/w9
61QumE+8sKw8OhWBE+RAIeass6Lx1bxpTI6m7eVSaJ2YW/CBUQM6+BxTPv7wuozv
PSDlYi0ugNpXkOAAIuPbo1nOL1X+OSwvybtFU1jE7GrnxLqE0MoCCGxS7osE3RVF
KtvaHUBt5Vay1QrcGGIHw4EFagaRlZ2qpn0RyMPkSvK9MqhJyfuPUK39MYz4EGeC
dE/AGJbsO3GrPzntFpSXIFsF7T5nvSfMGiziG/dWAEu7GDNDy4OeHSELxdr/88la
qygNKQ+m/AX/xlLEFAqjmlnOuFEyO7SyX2sgRM1v0unt0xqRIZLHARy2pooLArHE
7OmcXx7MfHVGo19fCeT4Ukxoza0f5CIGQkOU64vmGehdJ3kkrbYuZ3jNLHB/7QuD
iOUF96W+ykx8MKEjKa1rdLQsGi8kIEuEob1+RKSRbMYizM86jSIgVGaC4Xl+ObMD
VT3eiULlXdGCPMAlTwzn7PCM7amFeIdgy4cCQssGuuvxxUt3KmJw5dfMJPQTr9Pe
sX5mJ3BWKa0FtJ/OtRIg5MBR190EeXhwlZfYK5qS9a9kNJkrmURknGHkAuY+8cSc
AR4yrykTyNorgGn3klrnnxU60BGM/0z8RrlYQ1rkOzxCIOmX8N10OSpOkc2D5NIW
4EB2JsF06hObuMuhRN3SvAfASq7pVDpfG+vDVn9LZORybYz2dr55+OH7YjMnx0rh
MReITvWmvaa6R9Z00IHqjFMq2bCq8zYFy6x3AXh0tc8kOGyjigvDK5RXPEp+rrVy
iT4cxigt/a1svJk4ULe7BOftu4XJ/W4edtHDLfw6DM1QTxUXZ0GwLYytQNgmzuHI
mSfIu+3YH3OfOI8tGV45nPSHHEkHUXRahzYzOTsA0TvA0wifVAxpm3qGJ1FJT6sr
panCO/GxkQsJDYEVt7EU0P+XCYqp7IAOIbCM8FpL4HK/SL6gp+/+klTLL7vi6BQa
+etvfMZLzeCjjAnIZjPMGjA2xzjo/Wwt6Lc6y2tU4EzC6KI5ZNOcP3OYEbeJunGi
oqBlQO/795okgjlUcYftW232OXdVEsxNbazEnoY93FcpLjqmcuzfrOa1H7hbCniQ
fXxs6X4ZJTVo+fkEvUTopWyoTpxcUx1LwAcDt5PPR/Qy8t/rDnYphqiUL/cdEJBM
7HzRx6+WQxi62eOm34+UPQcxJG/nLW3sA3QvA1lWMgsAIrfN4RNzYD2tqxPOnBjn
mdUlFrAoWrxzfM+P9ymYzuex7WWzmdiGYLB+6LbINeQeTNPkhtJvoKzsk4m4zs8f
XaTnhXwEqLhhM4fx9QrTkuEEKnZwnvvzT9XlqiYFyG5OSHViyfu92mKAeMsiVzdX
LyuFyh07QN4BYiRC/zs/Pi86IRpt6eg4TTctX1KC25dHlCY2XU/dQeP1e7k202JP
Ei+W10jSXsv6JMyesczimmMkANhrh+LpXU7aTLDW3Y92y3/z/2cXY609z5//d/pS
CugD++gRnBa4HH1huKUAfW4TIhNJQZKXBIUP3nO2mtHxBlaPAfS6j36m2/wqCEIm
A6iX/5XkgUjL3MdjVE5HZhIkvZrk/J5+/h9MPkKZ9RNNTViltU08mi+ARon8FIRf
TrF2O1MqLdzH5DhRYTI6bmXnvk00kiSSa7u2TMW7nsPRH9Sa9K9e1WezitAfji8T
WPGgxI0DTY+mAUmdyhvNHVpQmLdGhXfkHAj14T1C10ndEfQIFlrlesGAAlJ2go8+
bNt7P3mpUi6xrRXPFLaHBPmYDJnP7KxB6QCnOvvq+gEwyBohz/m86D62cvLRp6FO
SQYeXmgBBGvAYMvMy3nltgWHnmprn2YZW2DnrIcJGNXk0Wj+UB3Lz96FvR2MvBC7
zhhc+UZyJ8ddvLEwOauBDSlBPZCFL9LvwF/hdE2iVHs+PPl8vBkj7PSMnAqIitPJ
ND2QyK/OaeSQeIO8t7BIp55a/tIIMl7n+UegCtSdjEXluZGLGe1+2XyyTVlh3GAB
0CDI+anfglRZY4hsnkeppq6ukReHHhifjmMfEpxvE8UEtVqsrf5pQB7gp5LoTb6n
PWHT95zPCR2S3IQ65UHEx0ok0T7nvenPtcyvr/cE7lNkIovspnNhA0h8HnfSFxl2
xkntWI6/qQWKGRnlXfq3dKwyR6y+3aEev28hi2sYkLLlGJh2pDHtEbrTeLZe0we7
oXUVUB2Bly6+becf6Nd4rCMt2YWAcSeUNdaolR1FYqSGZOftgLNCpEUbVtjYuFIr
XzyrqnSicSSWvkYOldnj+g7GaOAGp7ONdx/QcTsCClTAlQ6AVa34p7vC5gTQUtpl
Qu4fnmrK0QsHrH6slZBEnKnVIEoXqQ+OH7MsgY5oV3vUehXASigXXaDQXqJIKriZ
SNAxubmXgUE5oLSrBDwGnydIz481SmHjjJHw7DVQdNa1yYbUPkfU1A7qQ7laKgmu
9swpL2B1jiATz83dJXE+YynK+ZOLfl+MoytwEw6nLwKnrKqHqpmAIBjNLPxzM1Xf
aQjS8OJR4WlPJJIk3zjJOHgCpm6pmkBvlDJsxJvoznMpGnVhRfX+a9lTkKHQ+GVX
egI1PXkUh87Ji/oZEd6TL5Vt2hr+jJ0Y96J66F+9i6n398mRWYKyIz1IZUqVWQ5Z
xy5BI8vSc1hgTZ0LisGpDAJshWxJT+5XR9om1QFBlpGqMBNqe+tOgk1j9qrmJ/fd
qXWVHH8c2wvGg9zvZQr98wHcHSVV2gp2etdsuUzNp+UacyzNH2WWmUxnCK0zs7xZ
d8owvDipkkchurvSiVDPsEqwxE1p8/PJ3WDDDouTHfcEV/purv17Ql8pG5P9kpw+
sCjDYQ1nMW3doOgKfiB881M8+dStE1ldoG2Dl5idwH7vaLmjpmc5/MSzHXlp1f43
x1tvZX+H8STtSoe+yzvvaQb7HbVVYNGSAqjKdn7iHFT1lINLwuE96CFj0uTqvHjv
dXVEQqvNUt5HfOAmSewNSEXDZmVR/uZV5UPWt6I6dJj6bEHQ/BdB3E4Rk0iuTX26
aXP3kQP+Oh4jwXB/Spvvwsw9mXV8nVeU+BPYxYHtVGShb8nCEtClH+1nhDL3akfm
eJROBChnY3gRLw6Zo6jRxdEoo139MOMkvUWSLfDDAenLi+mkq0ZVSdRJZF+q7GkE
T7nAtvJv0xxCxnP8hv6nSVEHbmcrbdXWjppwTtZUYtmbey/ijKrWgGKKsTxEfpe/
vZAZm/3mdvp40Cudw3zbYk8cYcPRSx/s5UlNeXmL4dl1tkyZJFO5PY0mB0w3CR6L
551xf3Q6piZVFxiPUf9fAxvK8G9HPBDKzRZwgPeFy5nXLMboa14KhdpfHAdHcyHY
QSx1G11GGrTRHoo6Ovaug7J0UwOIJsDVwzyUqFyfFM7r4HgxGaMfVJkyy8dOh/D3
VKKPZhNdWcSsYNgezfs5zDaOQW3jTP7x62vGHUpdmxAtTK6OES6S2rmsnnNchnuE
LqsrxIkB/aYhbuZGaLwW8agsX50shmfzjzs8qDE8F5c5SVP5Lf3FLL8m3bLABdj5
MMK1L5ex185dxQh9C8m41MGqtyAVpRDlzDJiFF5WIY4KecL2vJP03txMxnD+Px35
F2LcsRUCJyYx9UcrY1byCzNryElS694I2fEMSnKuJ0Whg7Y/pihJHvQ+mj9w3qA7
mbDP2ZxMfstj8nob09SwhPRdFeGHB7Mi3IuamePiX77GOe/tQdql5OZIinURp9pL
mBCgcOasj9tfrk6TyQxKt97c7KenXwU8hFzCSue0zJDbsnOjGQ6tvqSwta84Vt51
EsFYMaiifWdun6tSt+IGOZnegu6sn/iE/vrXBoc+1maOwzmo6ZsR5dSXXQ6Xu760
LluAyX6KIBBruW0e3ZG7QZYj2APqoyEEVT/eREeQB5i2ZXPPqJjuv7FzsQ+o1y7a
6bln6c/nPiuWPVXo7NAtE1eIGmyICkVFsUFQpov0nekSaaGecsK9HOqngI3zLyi4
MCtssxkAN9sW6qmIGIVRvd4LZOrFPS3feKtcv5OsMpZu0qyPm3IhtuXx/1a267DA
0rbbASEFusobfs+95/k74NmBHzw8f4y7SucLHYxmCRn4g/yR6mXloN+F5aYy9xJw
w5BVSOurZV3RDAQl1ubaDIN29o3mBY+df7gpE5K+OgCnADz46jGhr3WrB9rgx2tK
o5wBY8VcLMpuJiayj1cv7LeilEgXWozGZy265YeSUm+OiJQ97ADRLZSqhDALPVr3
sMN/v5F/vxeQrxwlGpeCveGYFUcqXxc41NnHthG+E/T2ZI0L5AIsWTzGL8ffvmWX
KwE0GwARFdiMG+Jv1+mZlhRbsK+X4Wl6Ab5Rmm1i20Tp2SFpkiaKL1ARo1si67Oj
VYZ4AUChC0vkBzgXtGLCy/59zUdFwZVxq7VuqPpLujs4DMtdSZClRoCv5/Km21Cm
jpIUBNbprXlwWncRebZzp6g3VvVOiiB7mGeN5SX+yQlXyADDOFlTl3ObhyBh1cZE
sMWkH7YW3pISCdP95wN2msG50jhjqt47RE5wRWRZ+SNzA3rFwjMB5xWsESThZg0N
X2W2JAwEKrNkA7DcUOyFpuxxfzxuAodggi1+u9aOB7akSEIHP/9osqbuMYLAejAp
LZ42xDiqN1L5Lap0aD0RqpwT0UIbuVMfEJ3LnombkFjvjuxQgT353jTq+kDoL0hi
wQbqQlbtSzjJ+dcF2pwSSaiuQocysBWw9HOMsArfgNMNtfi72nNSfX7UUW+dIkL0
x3G/vyAZxZTWt0tF7NdoFVXbhAWDZwTo8SZXOe0M3v6Y0oP2+7oJpST3f840VG7G
3Oan/noo+Pf2gbQ23D8N0Sayanx3ZovTiE8fMP91zXT3FU2DXy5+4grxEvvJ262+
URI6BW3ypTj+m0El8e9YQbQWddcYZOn/tyRWoMXyL84XGdQTNIzGGXx1JvrQm5Da
fBOT6KwOSEtpqF8i/Gn105fRDZ+M2gEWhgLgufDaMcirSJA8yupL4imZi9JN/R2D
aX9XOsBPhk/uGokmBbxXIjfsHw1WGv2IodgLKqi5QpGWwiS5nPibnPPR11UdnLPm
EGtihbZj6VJ5kWOXC4neb8GV3BCEIVPJ9UVBF08yJ9N34PoxiiEqd3abYCCU1L9F
vWBroZdnkj1b2CHdKWgAil86mwkN5ZLjrLxh/97er6hhWfERMmiRtt+i830vhU2x
ZgTWeGwLOvs8+cwu6oA1vwFPCh6whEFwGHUfwAL9XtclnZygMlpN0i9v4g3uhCq7
iSpE5hCyZQNR5AanU0B2/C2/+GYUnG9U0mDViRmJGWCqQWX0bS3fBHPtUocDd28o
1RbY8ALUWN7KXSpL4j+XmrOKXxCJE3E1ly6+Hq1heGF35z/8yzauM1mgqIfktdQf
pMrtb1n5uLBYaHenbHiaVjqVBZfORkgtcdCC3FCcEMuM3oSBvsG7IFvUCrlsD7BT
RdZn7V4JIEVA0HbuhQaY3McluqK82qf0F1T5S2KweDv8sSY3QDBQwQfIlHU2/XWA
quDlRjTFiP1Qo7ozVPGsscGO3Sw8HAMb+wWEV+cDlbNr6o9kv7mFS+P5fZcgqjzC
eY1YdjgdSTYZlODrUfBpO92yJvLua2E4K6Mm65o6OnhvsvepUqag0rQk/ODgiy5I
HnnRn/Y3Cuz9TwCAFgXh6kA0HIvmY1+rVv+iaHpuO9zTfzpDu9cK+IWt5QeGx9cD
GTm+UBQcBrPuJXNyFLGI5Jh0PUa1N99LDIACNilJywtxukgm3Qj5+L2a0+HRz+wj
QSG2EBkTXwKi/2B5mmn7EOIcz5N3SCZ1HpklUdf8kaWuQ01XeRQxuKl+WNLHxzsu
CLriujyS7fH3LyvyxK6wqrg+0BiuReqCOn3JzzgXT/T+BNr6kQcO+mw9TQc1V63X
FLDR9HuF0uKZfVqABWjJFFJFwbdSm2+W9H6qY2HH5Uv9FG72Z63VdAemyGzSmsXN
bfWtf6ghRQv/8oKx9bL4NOSQ2UNlHUOXmSojhEMtsvMeNjpH0wqAHbKIRlUkHm83
5MVsiWLOgbZcpJU++q2jHbFdDRmuE1MEOruouDpCHs0sM4siGR87LEUAMTe+8D6y
MPSqL+3m+ur27IMpygrSV/3/tb+emB2v+cRQ2yu0dghQZVuYZCQW8kN7Ly8FYKH9
ptOs+4EJncxzEgiCKr7dBEintK6+0Ixv7Fwp3TaUQOX6XeoM204U65x5lhsljJYo
6+hYvfFlJQ3jWnl5SYi14jrR0TlYlKgxnZvqXlikuhUhW9OHrwZ2nu1IOkj4UZ43
epI6Ts81W+hMb2cIKIr2v0mT6LKBxu7RJDX5Olw2IEgMDK2x/AdNl5+LVpq5X9hS
UbzOF5CrtDR2GYLrgXV+aoEzYyZfvHbYu2Si0xZg96Cn/PVxvtsA1AUuv3j3F+h/
cSxcXFLaLn25dLibuaG9HFRNHlyJme0Am5kfajHYmO3m65Nng9Y/ZHUzzXbA/XgY
lcjDPj2rB91geC0Z3ZNY853UJvpPNvLovnkEHfaatbpXj5Yg5BTWRL+X0cowwlia
DcpBsxdIbO6mN4Vletr0EooFanF4ZWsJdsVs0XpzHpkkmlH5F4AEAZDIa1rSoJ6X
wU8SakHc6ASgl1+Uuej4xfhs1lMPWNlJ3TEZ5DhcZpwL0R3WFF3bEHP0MsOnp8EA
S8DsHEqpWYRGGx53MTpq/Cm4pi9Sje+FNlpni5/WrFLi/+NjSv7QUlDvzvuTOfOB
r4lHkStY3PDiUyzc95g6UgAQefbFHQyxwfj9mnwyGVI/T3z7PeJo+MtKqL12L0CF
aVc0ZwHH8FI9mTaD1WhHvbrcoutXxgsglwkF0iwnkX1o+PmhG0gtX+lr/3N82EWH
Si7y8F38n+EsTK/NW6cJCEHg3hYEQjU1YgxW0SsVJtSukj6tWWmfI13hsin/LZ5A
N2r/nfe9xIh3YEMKOd4oNJVXQnReTZJjLYs6iD2X2gR0n94i1K4WOXEDjmnwmsHH
r7Lop48/6sSbRG1mojaMshWGcfAZTAOD7HRP3Dg8HBqAD8pzG2axAC0y1ajsuRy4
W3l9S87vfA4Bh6zelninWsgjwWdOY5/nIHLfQzlNjLqxV4NLUPQRDta3T+Or35jR
HcE154xdegZXSTdsJkOsrr7kegR6Zq8Wml9vnl4YqhXRzzrRtxw7b4/XVDHa2eYm
PFrDc0jqiHhTzNHcgr7vk0DUujRKBr5RGuSMaHLNYlvDUM93abdWGVTPgbL17s+9
P92MbWYTaSUkOjs3BPjptjRHLQvmOGacc7FA/Yw06kqlBIKarYtSTeZbA/ilvPUl
llM12zDtmCFQ/WFU4hT3XTPjdxBv18OI2qy+BKDFzQhCSHWgd/Yyp5fi94O3MYxZ
jkTS5WeWWc0KUtyh5NWO1fRHWKoPl25YKJf/jHxloPPjRbU0JS/hCogIaCwEHqs1
BDMn7FMHsM/laqr8nM6LhMYMORce+Y4hJygnyHtL4JCSY3rUJhab4l+mewcpd8yu
ixX35u3Gyh5IMSlh+MNH4XHJHgmDpERjIeIOd+Wq7v7knG8yJnVLOHi3vsvqoypo
sPoNioQddOubxlcLagNPeLA3aGfd0+R7WDTCLr037UyF6vs3Vf7ulUAmcXM+Q58l
/mp+KkO/MKmcIavTmq6lUE+M97NwJRien1vUN4GI9JcXcfjbSuaWNE26Xm/yA8dZ
C7dsUSLE58Yd90yWb3Ff1o8eUtqeV6N0UHm6WJlyh9Q/Bw+vNe2DVo8f4dYumBik
uOraMTEkCZxBYbcLvIxm8XpFUwkosBSWes+/tDVa9rGsVS/wY56Kx7UDniZemvNS
EKgpjt4NATeN0IPW8xU46IjtI+epXtLxAEQcFb105HGvWUjgFuaMWaxoMkX9pCVl
VCmAu3RdZmclmyCKspqTASJ/Q/T8vUG7gWDdy2iJmFLzSZlEuH2mslyg5IhmF+0J
8DDd50S6QXmrHhkRO8yJU2UQJ0hIpAKmH3W56dcTedMZBo+JRCDIzKaRMq5oQTCI
yKbxik57gUusiYLdivpmntoYno8RuLdJftSGFeF+CqWMZ5TBo3T5rDlUm0fpGUCD
gFUddHfsWl0Io7rYnTul0XCtTKifAFLRAdMn4bGe3JOWpV67lIkjupSUFogxGR/U
gG6TicW9gesbJgqL+KXiXznA7CPF095z3EE12F6HLlsPTdq5MhIIhaRd4sO+Z3Xa
FlgTxs5KvdV7vCAfQW5+2LL+1Hbj6qsMuHbCXkWs2bmNpBKpN7GKSDZLiolYQX0Y
Rss9S/3wmOz7fzB1RaCIEK2fMgcST56jS+cYVa4dZSnWZSCpGLk7QYVa74I3IlXe
Q7a3/72OaNikwqTOBuiteTHZoRXIDqsPcl+gleatzbdWoLscmnV/DYx77JnCMlmp
YL1X5ru9jcf5BemGMtbMev9d10FbLuoLWONF2hFAGLyvbGEELGWoWrag+6BwLqkI
gqLwdIKQnIwAuOksyUmTrlNGPMzN8bqdZAqpOLfuSQa2XawkCDGXpX6g2PocT/oQ
YS9O2EcEuAYOZHoqBDUPJC0byW8i7RopSdXXdBx1MSHdIisnroC4uQkT2j92nSG2
v8Em15fNlo3SJ8SgT06C67Nea9dfCiUy/ildQSd5eHQ4btLFOGsqvSUJdronVsWh
xCPNi9pDP2SUlQ6tsS54pl7V/XH7E2WT83BHw2HguWmPQ8MQLNbJh1vJuFyJYYHW
ExA4ele38U1yub0lKankyPMx0xm7lukRrg3h+uTBX9IB+PHKD+nyewOtHCpMXASQ
sn4ULzA5kZwbsI356k2fLR9TKkNayqgO2WC9LcKpJ/nCBeMIOrpq5aMosPc5Tscx
1+oLokXV9bpVq9u5E6ieCec9WWintQGIxPQrkcxCglcP663QaWIAxiUuoPQr27eH
F2rGWbOlvCMObpvUwM6R+JmPe70biMoniwHMeRs6lVOO/kcfzpU8TCiP5uoCGn27
PNBRc9xHTi7BagwycBQrJSwkJ4us8xpNPN9Ifoi90Q1dnnM48lyfFhbngR3lCOGy
iHctXYR0MBP/tGAs5Ka9qXq98zcXhVCz9dFCPhkUqZnQOKICt0Uc1CsWmGy0pI8y
LncwSfJPTJSNxSt5WiwEOgJB8Kfo2Hr9/xIGYY9rAr8CTGG77azkBhVaGOSVB9FN
Ljf9Vo/HWEy9LZ357GOQ3PrZnErGgDPWa+n941/f/zfB8X26c/ebjUge+yvuE5kH
fxLjppmNKI4b9ywVAATddqGRCSByM7h4rjt/jckl8GJ2DnMRH71U/CYJfw0OEBVF
ask1HPrfjzknj5lj5m3BDXOjr8qkdxEPkkcGT/yL1Prg9CNky/ovjEhgak+j3Fzl
TfhajDTm+zJ+8/WrilzZdoovndSmLbxrAc2rM4cmLbEYnnNll3VV3bFlcMaJs8p5
P91E3OXjszksnGCLLtOZaDrVQ62iRSwf4j6NGOsT+iagaD0RKQL3gCqavX4OHEDp
kcSgAtyGbWpZfAORKlKr4QF+FmlJb0ZuycUj6bDRpDhRlmJjEncqCzqyxS4AOOxQ
QlFyTq7S1PktAatTKiXt/uDRkGrsOSR1TKBUbk1X7YIEEQhIcc3YQZzX3eKK+ip5
jq908Ca2yZAGfBpDvCTnr5P1LhQMRdeBo/vxc0uznRqueoOCQSwjCCNL4UcRtbz2
y+JYzKritURi/B+rYuWNeNh5l5Y77svsyypDDUVgEXzC9bG76XHS4DIXhkOJp86S
bXyPtlgUtPN/V+ZhvxpW+dV7FHrblGXyqD8qt3xxGr3b9netKi/ePyvHxXiE4Jvi
Dyk8mu39ZCxDFNmwY/qqd0Vrivh9HR5icoGTH+fKDl5oDCfJfxfl1IbrBXBMG21B
uuWLip34l8gw1y15k2YsGEwpkJTI3QP26j8asfkPa/vjboCujMFkBfrV3qlkv33a
lfcjoGBMRDlgeuYNdD0xG+ReO2iy+abQ5g+IuYedS2OwclbR/RsV2108+Kkt4Z1n
1DUiZlcIADK/RKpPUHzvf/50syKT6bh3oSbqlInOa+x56nJ0YCR3xlcf0NPr6VZg
rpqao3lUSZ/G6DEhhmViZPQI9LOeaANbeT9ONVmdS47W9VcZzzaEl8MmPk4Ueng8
9LZT4hUAwXMw2gndSJq0NxLyqrleXOoO9gR1lM8kSQDpD1IZSWWtn32Kh4f8ZgqY
mBdmfiQbcvr2nWBimblLv17pdlnTlXPIAT8ycZf69nqONbujanICTyWRR4lZLoeU
RjaQsgsrA1yp3titphCo7QuINAEinaLvphYcJTs6IH8eD4IaTJ2yW3dd93UbyK3S
cEO2EyA5tCVeAWPyKRO0syLvUd1gRs/tyXejf8U6VlBB5jmTrZRDecWMnylZU8Ad
xpkuypTkAW9DEKYZD1ExeWZRY87U63gvbGDFMogg2xhMJLI4Y9oFtRM6mJekoNUE
+3SfhQ2M50JpPkoQYyYyfCwrPVjjDN2rITDvlLR9p2zA4W8CfovUuP+h8/w0i5kR
vkLErUTYLbthKC/WwvDDGfqVF0nsaBIxTZQzaLug5n/xh6FZkN9QI6e+2MhRgbcV
M3taPrWXr8Zhot8z7embefY9c/NE/THjI7CHpBKCJM+K7aUqCc/FXm9+86sPKm89
vPX/KJwIiWmLIakCJmyjRTjU/aQDAcsu5zZurfbr/K/pzh3RpOw9Akm3tRHjtQK+
LMwsfe4nwB82tCh3l5qU3LYWFsQR3z8LSZeltRAyHDKf25qiDXCHK79lvL5hS4O8
zFg2/UpqMN1B3h46UVnx/u/bhr95BhwffFh+aZJCBJVnivpKlBZY6D1VDfi/+rWN
XNwMzLkYHOsDITQ3C/Mp3GLPBydqU0sACjF/UsN9FYBC4uA9v+2kuAKkFwqvq/6G
H/2jg59UDl9C6lAsyGZl2IZnnmQrmz7wQ2/UZFxO/71rZwZsK9Pr/CSijzEjHFVj
K4mZYBo9C65Dc26llT0vWgU1R+5zf90BJ2qITbnLF6b/CZzIP+eH+er9h/EeIIxL
9tgrjo2Y1NLHi5fbcb0moldFFNRT+jpzmHnrnqOboTeiryzw6xaJD/fJnUYbtfId
DxuZaL5D+UOjEeWUURz5Uuxa0G0cJ6m9JbqN1ttV26u8W5Wk1cq6F0m+BVWFUFdx
eGSxag/nS26wdkc/lhIgxRrWtf2QlUFDkZR7MIWmMb0g4R3kL9B3jM1tglrv9V+p
igGz5odUxi6z7fu96RaRQh6HyZecWaVJv8nykeARlps53UFSm8i9VMvxTOF+m7Q7
YOHuw08Mz97RU+SsefCcV/q4gW5FIm0BCtaki4W/GjidQMXROyGO+YAj+iLyP/c9
14ZVn+NUDT6Z+9MTLBQZOt7szrytYu3mGnd92uA+CrXeegmfjmVrJ2OOXuN92CXM
CpjMJzSwVKQR3UIphr9JcNhu14+Lj6rfoq24bHNJCIGE9dcXVfC4mlySiNJZCuS5
ysp14CraQOdVyqtn2jNPv41q8y7tDrdJQgiEvFvTCB57sVbRcD3GmiplWWtsfw5Z
mHCBmqQ27EZTyilNF/NlmUEK9OCTEPST7cghuUjHcbSExUe70TPOmUMOrkgN/m9i
gx24OE/xoCySxCbLB3nghut0PlZ+B3LbKS8sZCJ9EV1smEDTKicVxTO3ApIabbkF
dB3dNjtvV9hpKK/nvq5ZAmybFyfdUwVfdCsYSnbIR7Uv6A18arrgWL5wBq6LuOKS
1riYX2sL8Nr9yyB9BOVIg6/2RguZZ+MB2xZXEevuKgGkqlzKbYQ0iB8HDCBmtqBb
Tjd7rq1etWjhKLCHGYaJxIHbCuTlFkmzpmviL2KOS6kOM6bSH2f4Joml6jiGxT4s
CDGp29XXGNwsBE4oJOc3knqz7OBiZDvr6FKQy3/L2KgLUd6zzhGAqZWCle3xh1e8
7kZvwXmw3icbrlGxycUwVtiAPCsPiflV7yW4rImyYH/nAYC+twijFATVSaImJv4z
d5EVs5FDwfYxBVwsurnoSi0rB9FH9P9qHpwxdjD6ZTWtL1OhDXwd0uI8TgbvnAE0
0oLsn9jXqt8JWiBGzLkt5//YS1sQ9AX898BYSmLZMdEtRosZ1ZC+RR0hfEY0N+Zt
Qc/0BoY7Qp04IZlEfTqmo8D/tSy0uZc7y9Gw94R8LwkS0PkDIgtXYBtjSDp9gZld
agZOBy8FRexOgSc34al+cwmbMjnhz91633jyRmjX7a/y6NXDEjqamskxmw2uXsTq
2PCJF1u6PWbj3lBpQj+npjPT76p7Gccl6UD8P4NH8Lqpzfg4KE/vVjEHROOrjD9v
Gj8/vVRU7HQm3JNWldKQPIHrmh0ElSNhmIdiXZ4To6nN6t7r4K4pr4k5l1hsRic+
1SVV6PWgw422gGV4VOsslm07kmt3X6gjCmaBeCWXVTygi2pi0CD8Eyc2Ld7wSEJG
gaKipDxED4GFXydZHf1+saZ8cT1O4jXHzm8TVs0E1Vv6el6pQgYl2k0HkOIbSFRi
sz79FrMbVyW2y9Qrb7eJXdQJEDAHb+fYOsuiawfnAewYjVVmvty//AaJwRej1ZNL
2sUXonlvr5RUfAUa9DBvifIcRJLRK236xSumttWxuE8h45T7FPaxyCHNkxBoClJX
vqSjzpPMAuKyb1fLudWYFhEbkCyXdI1L97vcjHmleY50oyjWGLNjuuL9H7cP+5Pg
REMztfdlbRz5arkEkdzUzSY+UosSdKE6z1h5s6c04DNqWIX1n5hFVoPB92a5wVAo
7QiHe97+rFkVhC0qwk0OWAgeEvxN94U1EaFVYhIpq9WsZvhvdRIiDQQuSugrkl+M
JXNhlfagEflvzi3S5Fli6jgDdjiR3rS7Rzgsp57OHJNtEGD3fKRVOafE+v8kHrwN
zZ5bk/YnWWqTgJUfS6WMcovjvyvAd67XETplwAksFtvqtv7jjYc5qTrPnysABhwj
I3b9NuZvNfJgSWFMDOvXj85F6vQTacioe1+DBntZjY1UAhxwsO/b+5T3OCCz1UCA
H+j/AHjsZzSRS0bq/HMlvneaUGdU2UcrOWI4LR9B0VPzJvYTHoPyqk5HnVgszNvs
Mimzt9Dn64vKMVfJ0GPTtJIAAZrHfVL+2Bh0eeEm3BtFOaj6hWA2D3MdWGXWiqKi
y0m4CKiDQI50XeqXJ3rJ6s/U0My39+W76vHdwlyIztxBj9lrUludQUAtYVs4cGra
uPP7T++pBxLxXQjL1iPAPs2eameZJZ3bZjhvt1he6t4wrQfrj+yWLkhtKunqhunZ
prSneXKIffTw40gE8e2K2Fbm1wMkk56wyP1c/YixyDTWNhSHaCV76VslsqLgkDzp
audvsYIjGgYxlSC1qLAqbHV0Zz6eHFuG5g0HIqVGjT4G6z7WrXVThn1AtTmDJ0P5
a8bP9rwIT6K2Awavbug11mW6+ZsVRQ2umiK2pq74BQPBAuOmEQzwnyDm7Tz61lXt
1//N8JFxkdL3Hfe/LQmC6XPX27fygjgF7QTjlVzrsy6mSQu1SvXA46hWx9vKOGxG
wk9YrB92X7YJyBD24yfuxEwkDtW/4i7tyxJj+2H89g8uMFFzQvuN9wik3NHMFze0
VE2pj97Z4H4SEtrt/DJiRnWaFKnxgEsq+zz9kByyFiZRTSdGs4MOPEQYjharTLHe
CU5RfjANdOjTVr8j10j9ChVWIBkMZss4Lwlokd5cKg2kQTAe9CUctf4srrRbx4HZ
zYGqLPTQh2zdZU1pns4KvF6PnD14q8nPgAQwaX2Y2RvRU35sRxd15Na+F5PvEux7
ROfdyBc5w0gfoOCpCMKjNBFfUlI1/q6fjWp4DR9FvLFHKW/f5I86iz9l1WgIxRd+
/ng+cEIpXyXVMd1qRNLab0KFDLc94XXNXtBFaNnhgLkUcgTbbOWj6stYATSs44//
FzbhQmWYlvHuOg1YGoxk6HT/nrg4etyYGLOk0WNZEvkYMPdMerr3e6Z2K51F4y/H
JqlDZsX5Fw/y4U5vyeXuPk6TIu6NRlq1BpegEenLHrVCtPh5VQ4jAnUNXwZ1s19V
JH4JqsA8El7F3ls7C2aFgtGmSeHfmJeadpy0H2qRWVdatP3TGgbHKkx/8ok7/6l5
LlvI7IMs0rlSiETIDMnFvjwWPJFUckV3g51ORBkpQLrvukP90BJHuEDN7MolQVJn
ZNm8wK5jGVCXuQpdmSHgR/C+pD6rqFXwoq6aSGQeZxMv4UOLc0P/0CpreqCtnCLH
rXH8XoxfDJbWMj7IcMcm15Emv+PKWO7ri1N7EQ29rbeA6GRNh3fqGw37fOS70o9m
vujhwVI3sZqpbXQ3H9vQLstBcSMm6OOgdo2VlSAEFrqqv2DRyrb+eEpHPYUvTM54
mcV1ZkL4a50hkMNqM7/wAwEyusEDjLsM5gOz/DW7o/9TY8YDU5gJrcr4eEOd27Jc
Oyy6scZVytnXwiDrBZ5l7emsyvHo2UV94Tgp4DuDaQt+Ws150eVWeo7gKEtN/nks
kXhTRlAc8o/t1doM4lmfKemUqJZCh3OGyWguRtNwsM3DEMKzHBfZErreK1Hy4AYV
KhAK14MjiBJkHTdO1ZJsyivVrVqyJj+V017LM33Bf+QirsUlipgl682/iIAFlDz5
4Hf8gaPBtI9OkoCHlqnWMRW4xhGH6TxNWRyVdsef4AFvDEIFgw9c1dn3LHIzPsY9
bLDgNT4jmR7N82XIqelLclz6uPphPlssUHA65ObOnXZG/chPhFgg0ptV5QlbWrBL
T83VQ4cE8WO8NT9LaczK+Bfy+IXEnjsNj18xQYixaiNFL9H5JY2upe18WJpWPKhH
7R7emDHiogzQySbOtpqC7E7tgZFvMH+VVGO3u/bHF6d+YnM4Bcz8Q+vroHuuQ8UD
ElxjnNAu0MQEcAmhnDudfJD5cn6E6n+WCWDVMDtpW1GUuEKxXA3VVZ89dEON2rzj
r26GiS0mLGzcZlZEL/XWO9PCKBbikrv8o2gmmP1nTZxCbbFn5LU7rtUBBcXmMMF5
czwHLctI3zYBqPkD7uo6E87pQ8aByEnFQYqXFaK6cnDL8Fd/niVl8Q+5PWJsniZ1
rcmU3861ptv5GYS4MNotWoCjg9g51twb8UpvX+KlTlhQyWUuJXBsoJrqg5EYm2L+
YGtjpn2eVSHKD/BEEGCi+Q0ERss4I07EWNC8ylEVfxgoDkjRv1sTeYWcfz9f3N+q
UU5vYt3sIkT810hq1nZQ1hV/SHX+RH5WXJ7YRfgpf3N/UsXUuL0avcUvkvU00qId
smYHlTtY0m8E2l0EZ+sL+3MuWzsb7j1IzUuMJGPVvpmJXFHDX99PSVLo7KgU0eYr
4VXMVc4Bc6Al797LIXz45Vomg1Qc3W5llIocv/y6de7fuVQK4Vv3SCHbzyqkpLJ/
gbZ/uMhCfQe14GxfadhBxI9Zbr76xWWYpbjuvqtuK9h1uMEwSPvjSw7nJVB1SI+l
+g8GH9HwCcTMhWubAVS8CFBkVttXimXmkqG0HfYcwqGlZi6ED9P/RlWTrCaFUyA+
e5494LuvbKi2ht7YOOUl2dXsr+xbmKLSA/aX8coZRNkBtZ6SawaGWvKl/2GA4K+P
Ovz2JwRXRUmHZwLHzATGKd5Hj2xWX8Qnc6WSC9uwipBc4WQpshSpuo+f0axNunra
nn3N58hSGonuSAa+SfzGlXk9/9wFQ7/CcmShHLg6XebKNGkOocG4DG94kE3buTpR
TRecZYevOVu6/xAUi+eAFYnWMyfqI2AmBvJT66wnwSV4QSazEXyyNXWMp/XAMKyv
G9fDQ+VJP+CGXUfwpzpmnkgpH1Wo9SexrMdyy9cAlyetlR5L7cBxo+kD2cz+25rL
u7o7l0h3cNlR+K0oTQYBMoAR8xgNOQHQftGa7pgXnPl8rgR+hjGG51kJofIoPi5n
+F18NpsrfEwwI5c8ELbRKiDPoG3loHMhIMo+XEATYIVWFlW5TNyh0KhngZ7dUil3
SFe40snBHx3NH5Uk2h2yqAICn3FFf5eruJVC/c0zdEj7zFae8Sv/ECTJwCs7W332
mOGweVpxCqCYn0z1S6xkb9Mmj4Cm6Im55KwENwH963mxa5lI8fP60vE4N8XKXYNN
S6zK2IEZjGOEws6wleLoFC2RnXSFXCbitQ8pgStnARXoJsWy7gAo8Fv7lP7+baTh
yzUH4ueyYbe75CELabEtxam920pCL6fMsnGkTLJaJgMgpXyNY1G5PkIcxvsqP8Im
IlviMnDfTHROnJctgvhBMSSeXzwCylwYRkPatSl7O1+KkSnpSvdsdzLefzI7EwUc
4OHm1Ye6xHXfJLaWhXSIPoVstIPwjqf+wCCNttn8FRbOA4uoXORq3fGoy3KKkiwu
UC7O91yIc/aLEjM0lidVkhKbCzlRGd/a7mB8lEAGzCJN5v59Mp4iJmKZYPR7tqu4
FrpIvIDQEREb4LAkdPdXKlLRDdlm1IMh1NRIreSKPgqV5Vh/9EbaTyXo2k1e6WO4
X8nOCfF94uEElWUbJnWsXQqLsLXWN8BlBBDZWf5xbXj/1M/HBiia64JrFsYzKsaR
SkLsSXsoYNCzeu0KXOYfXtiIHVRqHxS9CwKatpmGa+Uk9XK5be3ci44xQK8lslf5
MlPgT8N+0jGNdIFgp/dsgKNZJbxkk5CdScBgZwPz5CIG0KvOkV2aUUfbrfX6s8ah
j8LZMFbapCSmpD4YLprjMWCb/HJh6/WhcMVIBeBJ7gsmAyc4Ub8m6g8GH3C/yVb6
ipjx+o5HfN/ITTwvMtd0LmjewQh5ChRg2gH+ndnIXpWA6uTT9XNEaEiLPFh4VK4r
ORD7fNeU2xURUtUbujvxbmcq5MViSuxcOr28iKOhCnOAmCPBoWzvToI4HNW8+x6o
JDb1PtA/nRH8HaSS4JE70t1DK6XC827uUQKcdtsSkg03AbpGs04BXTOF1Uj6/9gI
BF2jBaGNndnT7eDRWPg3jM5Omvu2UV/6VkbdFZwX6T8mD+4YvAYP7u0zoq3zWNku
nhJky75nLxKFiwmrsUS5IndOmiW1LxGlf0CXUkwEqKu5wY2V70xtodXtPBqcXFSU
86+6VcUOCNvBcE6oz0QxGcyu3LULCmWXtiHwrzZXitzdlEF+Fwh2cFLUQP9R+mJo
mdAE/r8N1d5hi/cP02j70YkgmqcH0s/GBF5ik9UjnCTdu8hWt/hnXUHGb9EI2h9X
hyvsa5mRMnOMi5voaKqr23lHm9osBxe8PbJyLFltgJpbuEgOkuyENGSY39TR2xmP
ru/qSboeuhDVwcjGL6DeHdrm+w6O/G6VFj2qMzrGzzi+KubIefSfQPtbGdENtUYW
PllzeHkSGWj/d4YLvUH2SAeHYmXm2nLocFBdNt/xYoEfXJk4DFsZD6JNBbVUOHvH
oWsUu3NSNlKusF1mg3XqVLQJLnjq8di1wBNcEZCdOE52dr+PfPAPFdHyx8LKtQjF
rzDExaVPiyG53+6LE+EhzT+vjY3PfInrUzsJSQlaRCFCB5u0tUzQgpQXluiWlQEJ
5KUWn+7cvQO/YSTaa3Gm293olCIi1ZIlmiT1BmntzaVm2wzbMIbywcWFrGO2RmJ0
qijtfD0wweMyGaL0O4kNg3lRpjm1pBC2VqA1hyyPjgkNWxwrpodK5GApt8Fb9P2X
vu5BDiucnJCGH2O28WK2RueHht0OP8GJVTWFvYjRFIe6iPfXASVJ91akfqAmsFyR
Ch5NctqEWpS4d05MgeFkFdEolSlXtFvpc/gD7OdnXybRM9Q2HURh+MiqDEtKVgb5
MOoj09ecaZZx+L95byV6Ml6V/1ppSJFxM633s4VljD0hh1FnE443GdTxO8i9q5A5
rSXr6Zb6zxDixPt7DZs+91Tpg3ABi6g5MuojYQaI0AhZSpHzDr9dwhLu2zX0ObLf
TwtFod+O1lTl1BeriAZFTAOwRt7ehPA3Y1MvuwUWT1EJ3cdTS3Ombqz1oAX1JRGl
WnOHuaJSCrhfNtoeDCsOizHnrO0irOWBUmNKvYiw64u9PJ95RiDFXBrvbVuzcHjw
ty/I+TjBRCcJ7wB9xLtM0LyywouMxzs58D2yfCQHMHJpe/tt4QMiNxYSvLHwPiTN
QRoEQfTvkOAzD5iUKDnB0T9RDh2Gn+Qiqej29DqUFHjg7xBughS8ehc+Zfjle9P3
srgpzFfuDXNZgtZpSUf8YK001z3dZkdI5s581buMFHIbwnsPftKKynDDcVDqXnho
XpIxmGeJToZNd3nQEqMQrnBFv8zJ8vDxvHZM5JqK9z/GZ8ktk14Utektq3hQQXf6
SZSgRkw8W17nbPi6rdL0h342VJqHw9PJrdlFPE/P5JT9SRLwxbFj4WbeT7C2ygOW
YuURnQcjDfiXsUVA6pbilg8hCaWcqgeZYsCIM+kulrvDP4tS1ERBl3EEBxl75hru
vGOfcmkbHE4/BkiRYVykqh4zV/lnAL/FRsnDPnBaxQsToifXzB4IvnLz4uLQMaWU
rUZ4nlnKTGPQ5oRe2tsjBaSRAiReWCz1WSZGT7pVmBi0I8k9xnxWXIZPE/oWxlO/
9Y4u3qCrGqhiVPT8yQknOuMz3DLoucJkoZ6rSa70vvCWo0FN5cpSBR4BnmbVmFPH
8fm4sEop6494nO4gaOY0XbYot6AjDMTZRgzxX/Y+sdtdo/HkPBIJ4oaUAIyhA51x
9nOhM+ENDQwwHnBQcRi4+76eWz3GYNzzBlPByBjLRyIY0Z7zzMi8CoUPH6aNWVLA
fgmyHEoUeB1Tvyj4b9q6uu9JFzQ+6y9srTEzBRYurAT25j4bcYfrIs2l7c4tLahF
PjyDh649VnkFITXbLsS7l9EmudXFrWF8lxhfQKQhiYU2oVDxFezLK27f9vmvxpJL
MNzrV/8q/Y4z9FhLpBgYaR3s9x+SBIIvQa5riq2iLYgm/K9Sj5EPAMS8gugRvYCs
N5BVQ4qCwAUDng2dlgbwq0MdSTTtlMxsSsB8p0yy9PHUF80n3PRuYPxoTHnEZ3GR
buLfXiQDTzmjF9UJHft1iZ9oF60ICb3CicOuO63J22oZYBfBZPERO1D6cEMfoPgR
B/ZyUl+53dk2cPLfx3G+uEVKG/9mnheJpbGUcnB88/5six3K8xw8lYiycJSRwWCg
eq1ZjXjWNu0iuDMLU1pX779eGPMnMQk/syrYGMXYJURsRsHNuaaWPE8PtHUiZC88
eKS3XVu+ZE+Le9g8K2IkOhTI/8Fdd0lE5skCCo5+BqtaXTDAecoF+nGmqJcJjjrR
HElltGlpzpbARDTVJY7OhhrmVEf9SiSvYHpWulYxcIaTd0f0GmOln9wfmFQg1LeQ
OnYfIIxRK/eIlIXFiLR+5K9a6IcWDo3z/i2331hN5sv4C/yyzhPk6qhZtuQxZooX
SEk7VpPneuu2WhSfvt/gT60tYg7I2k5mpfWAYLYtRBDJ4gCIGfUvKN3zQqlcHseG
znaB6cEXZuI0Vz9CtwcZkutZxXKqZISF8VWLAaLltWesS5S4Ru+mpaJBWO4m0FYJ
6QpGAjprL1JXDleKdUDNBJ3hzyiMRgwjk37Kp9j/QJ7Bylfwjk9ZInIF/nN6MYsm
1RyDMu4yyQkDMRaVwFWnCXVVqYzItvzgyyTdcyjkQWbs28NQmVU19wcfNHHVH4IO
rJx5mW4nOt8OT8QCiYzPERYaK5fEU/STd7itag6cbLpQUkcq6MdvMRCisNJp8a6u
8QtaD/52ko2TRGgXSsB6VZAxdnUV//MAxhNhVVUvjR23VBOkXb45yTpeM9VYoEbQ
UQrPv/QEGFs/2xb/zB79Y1PyGpr+ogTCqJuJD6qD8C+wF9XLr/wcL9Jpgo4Xj6DT
UdvRCedNt8MDJZK3oLHEJ80KgHKZenUNANGCG0EQmd2DRT2VFYtA6SBh8NQYRrpA
yMUsELLIO1WbN779vTP0jeQmXkrHZE9baEsbPV9AoIq8k+9R4t98VOyX3+/5Ql6a
xlSgvDmI60RpURJBt3uJMLKGRWm6oT/huapyXNZNqGvxPaS24VIsLoY9cpUPAD4O
b3qvIvnW9Eoc58hwN+8K6th/8soCvXO2tDFpIWuYKat63IWO8H0kFginbnQ/FxcU
GdMkTV/WqF8VAUqU9+19p2CXgHj0tQGRN3/9Cuf+48iQj+FrGoQkzYWhj5w/xaoh
WUs71lZu+bdA5K2mmKki915Vzfq9UDpajYeOivRByQjviKSqaLIgBOMxe3BynkXV
UpmBy/LPWRAy/Oq7eS56+/g/m+c4HYNtBhyAzcQnbg4BtWj94+FDTGeOX11hfPOu
BA2VJTeBkJpMF14nqSGQ9CJdhGqA0iD+ypMX6EQnWSoDIAipVwj6ptHStQ4wla4e
aCmnAWCV+vkS59wvCoFoyi1wSvYE4RZE/KlQNozzSqNcCeqcMzQThDvbLUv/rMfI
q4ooYJ7eEUW4UrxU/klhSoY41+zP1fD3sjnRQqUqbSpsNO+0BHtoY5MVxKJxOCnr
hF9Plm7ELIUKMPcuT1fsgD6jzfJoxLZAbDoSiN/UVshh56HFWWBQQzy00Vz2KL+f
8BgV+M+KZSTsJ/yu+cobqhxrEgdktUjCQgSYi5SvoOI8Wf51EpBJyE8gz7NOnz5r
f3UrIEMoX/PgsXHoxRbipF7Mza0VDFUPQWfZi+XAuodvRt5s+ddyc8l/yS1goISZ
5h4n32emt6B4Nu/N0nt6bcaQ8hlapanuFcGS3cgeO/uEiYcw54EQyh06daFRBmpC
XonEK9UERca0h8Y2QsQ26GKx+7gNDuYi0nfXVKD+Z78PSM0BSxCuxyJCZiitilJO
U5I58C77fpvFk+ENiP3SUog/Pp98517iiVcSuoVPOt/RFxPXWKDRGaeOWa7vDe2f
zXoQQwdB7ryu9F3pOIu1LNv6ahMCn8ahWZXr3ojK+SQlQfwyyHqCAGO3yp07frVs
shw1KBMZ4kFLrjFPdv+CPxiwNtfxdvj2e6XD0CsgsvAx7yaAao77JNidb9Qhphbt
QB6jwDEs+G+9luXRFe2oThPTJvBFLJwCejMgR01Pl9Ho0JoGfP3+HuV/lVRyO0J8
fyc7iK4URmyeoSo6hsGBSAOECdbvoO4SRFb1gLJz6Ge8G75kJMEoQjhhUsF+PaGr
YmfmgcB0Mi7SBGyrq9C/4YaFCZqCY1xP3bmc3QVinUW6qAiT7ROmmbn3r54twLyE
eT6hPwc0riN+4/ley1uRKLYbD90wjdQ8Lo6bQgcvbnjq7dyRrD3eEm8VySfBytL/
66i0Os01FS8PmoXK4XbNQYAPTEo73zB2/YVNpupWi7yYJsn4tcJfj3F3cHLk7EYj
yQ4gNyt/XlLtIv46GV+wBty57ner/lZvFgYtMjEgbBcsQr82yc3kSMfgZJs9GwOn
7gYb72RuZ5Z+RAR1nzZpDMe8hqtl1bmSrfOFhWoOk9rLbsUEe6y3BCClvBFtRN6K
PbgB/GnhrvPBduU8MjV7rjqI5lmwa8x1bIScmHECVOpDHuuob9Gs0mFvbO1XcZR4
/tKMioFklqtw3KXswrmuQttYQghdsmSAJK5LjjzB8TvW1lFLB5+H3dW13gZcneBU
gbF8IuvcNyAJOKUHQXAW3vGfG7vXNzvYJ5cvmORyTSvJUNj35zZf6/9uf73POZX7
P3XogJ66So98FTO7NI+0RO9y5TFO8cxszQyUnQkN1+EElKOkOD7IYTMY529fk7i4
OBAcbTMeospqEAGs5O/E+l70QPlRniSvcLMAUy7wzXk6Cj8paYkLNnSXOB+TOwFU
ayL7Pvzn4LxZWus+qKS9ba8/mZBM7JzSqSFsXx/4m9Z9YTQtoGAjwUx9eV09ONS6
6ZZ3bInqiUm86EZaTz4Ofj49myUZMo2LguVN8OzCS30TkvOQWE4JHaixPeOL9MWC
7kwjeybPgPNk6f6eTUQfc/o/qS0SbNT80kzxku2pTe8EMLpssCzxR9+WHnAnHBWW
/AylPs1AozUbY0Z3V7IKhsir+6PSwiUxr8GIEDi0p+NDonf5AAMvcMSdSKYXFMh+
ZDyKP5+YevQrzsmrTqx4oD2oDCWx73UQobUQEI18yV01J3R8tH5Y3GGMMK41l5p+
CrjEaN3FE61Cxs8II0s5/e+2M3kkyASMuGb38oz+FjctlRYISamIiIAMlCrIQkdk
TtuseNcup2QJl5PKZbaFJ/qxHqPDlYow+d8hRvwm7II85SOAC4PhIFQiCzwctcmt
Yn96cXoKhtSQhdYugdfGn4U2ZwBqRGHTuJFlkHEIj8JRok81JZbabynLDvOcdY4R
ZYsNHcC/I5CrJjG1sp7F+vwhZWxYT6xHT3dX7wNBq+jLX5OFZqOfkv0+ssuVmwwg
QCdZTCcgA5obQj9NR8TuqpCgyXM0pSjp6ek+Vie6L7U1ISvPSr3TE/x/lSSV8MTM
mhG2iShuQ1mh3hu3+J1f4wZhStuXLcyfiImSyGAMyZ+Iiqw/24YT2om0N0mT89Fn
Zue1SrwUATM8tU/5HX71u7RP/t44Kzc7YX3tXo2GrBTHx70qxaJ41xG7oygk+Spp
NbMe70XgF5wtDg7kRS9B3HPudY2WN8Xj1FQTf2JOdEnVwCpxyS2CSwhmB2OlYyO+
lBgIV/8hzx7dLpdEutJwTqVuzD0B1aoxMgFg/QP30vkL13EWnOYeHEjpOv+i5vAa
lXc/eS4OLPY9yEqGDQvutSxfuvi3TgGJbWA+TFGlmR22FITc4rQ3OtZdxz58XOxd
BCbGs1uuQHovI07xWP+gvIpv9OQ5Ob10AK4FLuPO2aW0iHWlDEy65PQDOTX4RWKE
ZvLh9R7Z1mv9YbXR2ZNwuOxjWa+vNh90UvdtKnyBm+2AbYr0DmHVhLsjnUp+RM3p
Q0F4SaQuYqVBD8EieOEZz/+M5jLsevxqXuMxKySXLWtpGyuLhMHMagvJTkB6IMn7
kPEZlm3Hi0qVxawQPJC+KlUVpFRlUVZpDbT1Q97uGhpmUyecslSuk7fQDH+GSwjI
TeKqgYxisYKhzNC6mvp6B/P6lRcliVl44AeumRU8TY3a0mQv3WnFyd/3HIUk6KoH
K7lAE8KvGmCeLgbYnLvmKEtAHHnQf0CqHCfnDWSUmo9p/crwolQ13dzPFJVrvolJ
bFVKLN+gUikwEmZ42suzyw4ypmMJk8V3q6qAV1X0Ww11woH2YVdbC3lxigsIdA+E
GbP+FMxSFqZPNgSQxdJXi0mqFEnQ8o3ToYhw4ovsANfIxMu/P8GcOAJv/kwS9D+w
DQ/FTp3WXGcz5gzp2jNoWATvWiqh8z8JR5UInYl6scGxVpmCkdUrfuV+2e7E6mDp
PCwfqu4hS6YiVQnT4PMn7XFyigH8Yf3TBqRIguuW7bNZUTate+ubVul7TMTfBL3t
wFLWgDQiqMvkZ9qq7XDTjkWyazQOnurNPumfVgQR/9xyfMh1mCUv4wFUiY/rq8Qc
A8oD3Y1efGDo/b1Ky+IBykmcth/JNqGd2jCMK9hVlHiW1bpO7XQiPHM9joVq4u0r
0cLA1PvZdIeY7TZTWn5HfTZ0sbZc1XsogsqiPz7t/mg8PQvZY9VopOs13WNKpD9A
WM/1+osD4PKrc/Vi+YQ+VX2yEO14ljZiJsMeXn4//1puhASsE18eazXrgSeb5lqL
8GQi/oOR4ZT0U3wlgY/qOJG3CaK6kyGgZa/rOrLftU9V5NFfUh9o2QKBM9som9hz
cdVtWqghy/Cjk2Kr14Liv6cj9Dkd3i7q/gm8aaMBSYVbmgL93SDpTHB1INAKkK4t
LXLVPc8oQZqYYY5jeStNDoq/3MQohoSupxSPMB5X3/CTx6IvEj2llgeJw07mdrTn
hznHCs3M9pUsRDiwrr7FjhBADiXYwCXR8stENyKqQubOSkyumfN/uh6GBRQE1c7J
ARkf35+L29fuOYQzAUi/lPuMLL0Z15/qC+kiuJvIU5dnn88knKB7M6S3/NEfAj6G
E5dBqv4nqlRGRmwc9bGCD4mUnzAXhKJUEKE65iE1LGG9jt1vHOMFXY71BroHMby1
KEBrTH7g0Vof53ueHx5+w1/T7qxk8TUYqdZyhkpdPdduaLJrGGK4Hx28ZP69gi6q
tzMp1fWptSsp+teNdsg2Nwz3IGZiq6brpY6ijbnnLUXaKRmpH4uJGjbqkplR15Pf
g/UeY+c6e79nuYKrnJoJHySuIlKR4TWjFloHlSutS2qnYQCr3CU00Qet1vPtiMPq
o2Fxtze14Oe3Aa/uh6yXMVuFwpIYDhs7OawLxTL20rkO23BX9eD2DmBSXf4rcrTD
qRzidTORIr/uq+ssz8o4i2wE2S3PAaVlDTFt8S1SmfAArraijly8DTSIeGgn3EBK
IreGdnHzu5zHCPY8noIe2GI8S4gxRKn1pFBqDEVlEmMO2x1Spdf99GSa/V2PqEIh
Zogf2tzkj4BVdONo2tSduUUnZI88EVT6W6seUmJM3pj0C89d1gHHkQh7iiXU6GsX
Hhij+LUyuvYDVRMOL8pQy57o/NeX5qu15RcX7asiWhOuEMtOv9et84mDZT1FALSi
STlFzkYmRSCXZ0ZoZTjdd2SUmpa878dc4lZ5RhIAcqeo0jfIH+u+wEYNtbliVkxh
k4zcievEgbgJ0jH4EWezKf9WC9Rf3/uuAx4My8NIv90Itv9EVm94AbX1Fowyw9sd
dlBIxMnbqYWEHJIo/kGevXJuAzS2icmkRuV82WpvBVnYAd3zU/iOKzXXyOOv+FvF
KEm9Wp13SleYqkSWFktB9K+9HxbbvUE7C0bSvPVSmGewiU7lxEyqFwk6w3T53773
HCQa0wGi6u2NpzCdcF3rrVpdAVZWAlQC3tYbll6ujOLRav301ZG9MgpZQ/EjX9Yb
BVwVNEUpIZ1BT2j6BkCleQ6SaEc6si+Yk7BCPScRP79l/3TAjPfkgkjIF5XzKAL2
2C8UfWSbALQoFwSh2bDhnYdzww+X+KwdoB+Y/k61BWXlbzWbM+EF3zjPDbqxQxxa
3txVNNPFt6msxywHNrN1Jqx+lA44gI+nEwjlx9OU9/2arq/kDqBOm2OpA+ggzOp4
qfT5r8+k0hJHhqCL+nGVNaElgThrEkLyWb6aNvxTZY57/92tI1hplCCtjpf3zLOu
DrwkBDahlIFtXjYY/qVUh3KimFikQNtWwNyiQxFeMiEHn/MXdb/9BP9Jt7lZhZy7
/IViaPfyUaXSSFMLL1pwI21ZXuJGFy1dbND8c5b2ha8Ynm6aXrLMkFn5i81tNMoM
fUuLEWDz0SZGeD/xMhDpcPNI5aE1deHq7AJ6zRnbor6UgVN7ovMR3AUAvKuOIvCv
QFOFnssaFdHEWw69WyUp6huicYlmY3fn+qXrJmhveIuigcoZj0PHAdNwlPXmG6gb
vlyTKVStMtQH//Vb0FenVjQsryMV9hH00fNkIPg8M8u1yy645S6TYiFni8gkE8k1
kW+1v8j9DfEzU5FIGYp596LFcmiDlmIJlQ/JQ0qy05geBgtqxpojJd6EOK8goQ3/
MnZzsnzsHGTU6HdXWoeDkYZvdUx1vAOCALH14Pl2dR5AhZUT3S5Lre2kJifwUyk9
ugMCyeqw077i9qL2XxM1ejqKj8WxOSMMEtxybe3VYKhEtbmY9BYbBI3w7mhwDaz/
8XGaS0JCwO96K2dum70gRfQzlmxCTBDPoStE1uYuhxepmGmleegmBdGs5DHXFLg5
E7bQJt4Pgu+kkdPXTqOqrlOj6XiGdXpehtJsARX1slx5RuVjtwZITEvgcmeMkl9j
WI8Uskn3BJVCRs0b/fCoYp7YGBOK26JUL02C0sH8GOqQaxZO2CfOn3P6yR6h8VGx
Kjt26n5h4R26hxzkeLkPUt4DpFEurKfdaGhxX/n0ID/5rLaTU0O73jLv18v2pMDZ
Jomk79fAJrGnUEjm1HfnvGp9gnNUTsocQT7w2vIl89w2OCgdql6RLD/1fB3F+03j
F4OV6bSLjdjxfbOkDl1U5bv2N2E8MOsA3keKc8bKeol4kegmkMxlFwc2kCCpRvNd
UkhGFp0WbT9qlm4tT9xffFnpA/KXL23bHx7Jz98KOj4wTtcdOnPxBkWcrRaCNQG8
FwHZvdiblXTY3IsO34S31jY4ty4JAi1PPXFLNEZV9xQCJkNL03LdTubICj0x239i
XeBqQMYEkY3Ac1s5tGwFCCaxEGCN+mrrrsF/yFsJkdzkObrgFHF2GWMf38vVDcx2
okwvtH097Rqs8Rm8RySQlYT/OxQAdZFLKv4vig7uaItbubXUurjn9bz5jIM4br/R
u/b46pyjnVIIndvJ2FIqY/8+SKDnoo41OXwGP25vQ/bbFnWRgUrbP1KRthQedqIw
tqSymZ19IKBWq7GRjb8Dxp91JeK6H753JF/d0gH38qRUYGJFC4GslLx9QHw0nY2r
/0CzaCqzinCvTPE/aocZeJYs3z2D+Kc8vKh9Dyqe8UjBWm/j2uerejFMAMLgvk9P
EsdkwbMfWnMayj8FXVqlZAJOdUc4c27ruGvHgY4O2yQ/sjsFY9sKQ52n0KEiXs69
qPy0plk/nNaS2Gjgc2GsuXIVTFLxiIsccykPmGBYoFMDbs7/0yf9/R/LP8ZGx75N
yfMek4dVANkJXajv6d7jy8+WkoDCaZDDLcGPTA/ceEMjx8GMWoB2Y15r3k8eJSb5
xF7/oYLER1YX+4U5tuorY1/dpGD7ANtOucA2Kb1pyOA3SQjzXS5s3O6tL9Vlgt21
LRqkDUmN+SmyOHmE5LpVeYazPRTmH62WCASRmqzp3PswdEvTsKcijuVJ0PM5YjiW
4Mf5Vu6MePvHg7vDNYUasaP2DuEbXhyTeTeIriXpOEc6CTd9mu0OXJburXszXhTA
zGe/IqU5CWPKE7Bt3rpvNQ3GnxhV0KKVj5qG0Wbkzbbi/VgDzW7ziXjdeb6vsZbw
PdZ5kbCeqxrrLB3X9cApoPGIr0tCME7TvCBYITX6Tn7WkSq1fSeBWIpVwTOqw4jJ
+vU0StSv2uHkoDqlJETid6g6YFGsoCJUW+LEwEkCKJrU5OxfFICzqiR5O6yGE0bI
+KRGau//M+Elnx8goKjABcuHfvXHIO3itoscGGNx8NoEXPvoMyTDF1Ak8aQtE3hu
hMimTOxn3nfpMmvMvvDqWmxQPl5tkDFA2QpRwHt+ZZdkb1BCpOeh5fNM59fQZQHj
Ege+finqc/Adaa/3N8556NmqWuAZ5hbpuCtXbFkY3Jko2TQXhlYaW6pKpqYAbK8+
tDcmEq9Vw64kGTnNAYNgTeU/2w8OSnw+NS5pQtLA2yLh7oddRsq3dmgwxy7Bdtrj
kEP0vKlZmsLfbxjAKzk+40ddbEW1m5Rl3SqGX8qMPwHu+6pGjKt4M+q/XP4hsZ36
T2eJ22yHo4GL1x+1GaQPG9mKfPVtEaU6X6LoQaa7BFXB4KuBuDwLp3D5CYwkprIS
oL19bqssq65O0Y2nZ2+SnhEoMnvwFpsVMN3JwUJ6D1wW9gayatcFANKIA0+rtTO2
i1uFDdW1rpN1vb9CSA8DLsiP8pSUZ7QgG0PehQRXi/015bRG6E8x33zwTd+14SLs
7BwHo2XurN7ZmH4ongiDr4IE72ZZt1nzAg9bgx/hkGsxp3U2CiHwpe+Tv8vqeRUI
cPUb5uQK5vjwlULIE7XMEZeDmr/jT2VP3FiViJfo7TFChvasbrdUggMjl7UILOl6
FdAV2bSDZRVMjjwXyfcMp40jkGCmHIAVIhn0n47muEQR/DsBe1jl9ceQ21LLudC+
4nw/5WhWrprvpyFEVf68M64li5iF2BXfdVfh1X6sPtIPVCOkxYnU4vMmQP0lpQDl
H+fEp4L8VBWCaimuqjMsa1RshF+VH5l7BYrdCnZWkpSGNZYAidEVnaFpVz4YLJew
JyBXCDlgGrdJC7bBUXdpcw2okwanW7QRU81u4SC3d2O8Q3RKrjeBGNo9RlENt9FT
mKQFLRD9MuIAI81y8CkE+mAlrCotYKnbA/W9xm3r7z+PWJFB5nInE+ij0cqD5UIU
ktx/Ad0R3Zq9KW3Y+b8zxJvHdSJHv0+CYoD/l47LnVG4by6OaS9gBiOpx9/M0FUI
BhDzAdrxRIqSQ6QrIV+84dv0vPkFrlembRw8LaAcfTmHWdqua1O5NIEQCRQQeLpF
s34KNaNjknedaxYB7F3QNlOldmB/d/qklZpPLyizKHk4yi7kkIFO9MLqDAMvwI8N
bdi9GsFNYGO0biFjQj9Jz9OcCcEwCvNKbs373X6xB7V73Chu3ur90C5K3Ql9bzwH
YiKVWocvswl18peHRIN1dOdiALQAnc3P6QdkIoIuhQiFcUlqZqijezqEvxsjX9mH
4B0eLTYYPAuCakI4dceNfeqiTR8GT23SWy747icvVeQpxyciEENpt6r+C/z5K8Si
i2DFNGGeG6eg2zzK5sj10QGWUALvePL3zjWBUNZmU+62v+Piy8oCrrgdTii17uEx
hxX/4PDCo3Zu2Tz1kRhdd/iCroe6nVIDZZHULm73rer+r8u9WYpDI0FGC3+2oUO3
stnFrqR7f7suHaJXZ688pJRr+86xsAEUVzcLlrfrB65wvePpDMIs5QTh1SUycFjo
YShCI1zoNp/US4KJzS/SqI3ljQ+CDV6Rjql9aYEAVEh/cHdzfeqqxDeD9lmrb1xR
cYcJBez5A7Z2o5g0XfaIBY1znKAFFx0CV66jpuz1CC3/f9o1mZT5J0GiEdCi/qn8
VjUMRA85za4EByk1KKG6msz+K99cjYlOk8prLNzJXd4wI4h9OGz8dcTyNg7nhw1K
LBY8zaC+4LVOg6+pZr5N7DJ0/8GZtunUBAyHi05xEInmyzjrD/5sH7vwWcfjtLfZ
5NQB93ePMjsDcHXdBOQ98JaeZG3sTfX1jNApgPvZW6xPWdPzuDileQHqeGd8aQkn
DJmJrgLToHg3LtRaHtzs5UZHdMShOUZEu3DzbiIQkE8d8rIQtRgN23UQGRbV/oTL
QPhCXXyjwW+qLTA2o0Y+dv8+GgZtcJ9fRyos4sFgIucYCJ0QWasRDEdRQHOPUZnT
u819x37CnDZ4YnYAghn4ba6xZqj7I1Fp6l/2wHsJHiUT+DPEW/0nQHkSQI9FYwrM
ghTY11OvRxKXAe5U7uMyiNfJFTANnkxMGse2GCLxez6B8/wyXm+m+90BC9cGnBDg
g4tuui8bFLpcXP/fOphYpGUbLzriKqaNwUctx6cBi/qPnnccd3hsvCsOdCDiNBfI
Qfrn5YZzfsUI+nW8zOzpJQgG953cv/edB79JzYgESoH9luiLvP/XFjkn95t6fTmZ
SXrklE0CvQk1ljuHdTUfIfhF5j9ncs77uUAcApEvvtoU7hLf4X36MQOn7EirwcTo
+7J2X6myFJOHfRHxnVR4YZeqbz5zY3HKX2oSSz8Osgf+IwyrwtTWWLq8DpUIii9Z
hCxIUlt2gW2L9vVjm4mcq3IhChAxfALLOuet+pviA188cweypVCuOq19s1sR4Hgj
hXz1C8NBjof/1rOMjydLaLbCqMl1tZ7qBy+TtsHdNz63Gv+9uEG53hTE3xgNE/zK
GDcFwa2v93O1tJ2yiDCvJq2cM13rqtXZibcbq/1VHuyn9tI9zX81/oigCQECpay+
9aFBi5w00t7jLytXjZ9VlihCsuRwJ6wuYjRr7Ega6MjFeAhNbg+sJpotAH1e2FDE
Ar34VfzLMbnS64jk6NVhnu8IFX3TGT1Hiq16s8T8HhEHshS0E61knwmOiOyS9h3b
9hjJ9TXCIBicMAuCdut7wkA0AMDC2IdaX/OaGw/niS/N6GVPhEsN7D4h41c5iOpp
enkFkd44LPxKspwv5wru5iXoWR9baBTZXHlHBh2jHm7ftgKnB/AOCcXqlcEKkb8b
7MWCZddqlC62sfuMTBVeUsHdIQSGzirkEGWODUUiTyAq4cEWQZw0i6cG+6dv4Qjg
AkLkkFfEFPIZra9knqvynh7lET7qHslkQ/uhuXtp6RmOA5EDRtBr6Ip28NfBphjB
D6xP7gvbLxl28cZ9DQO0ymltE0HG6VafG7kXiNB4f8AJ2tMcU7iqlx8qQL8K/vNn
Lf3y38t9vjGeOOpgL+/RXaYACnvld4FacnPlPaFgk59EpM4kBp3YmOj9gv32klFB
dsJ/g+m9sQg0VUDqqPOXrz6PuQ4UoyBq3xeJbDcvvvqSIk6mv1EmTf0NqhtIXK+A
nPPdA3jBbcaO19AssnvKJCcXtVaHMeRC80SkqiZbu3ndk+EP90EzNEmHI6lT2u7W
x8FxF+0pjTebACsAesIsd9tj68H4d5+N/aEI1j4Idlns7QKPMJiJcLznp5WnuBbb
9LucBkAnu/niIHKNPYRQ1h3kcMupQkD0CLODnnQUaRy73gA0s35a6wPIjVnBqLoL
D6ChoJ8hu4QmERckWPqfsI2oTLmV/1l8KRIPqjXL1a4+u5Wzxf256drmNX+06v+F
ZFpO/xiWpSC3l3wiZ1iG1DqhjSuulXnc4L0ivCPC8mpKNQMP/cM+a3ChzrWfjvVc
85B/+wEiJbqJ6CfFqdISMQXZxMR/EFxwF7GggQ5H30ipP9dhOZe3OBKC+GNQ0IMW
o8nRVkKJdBigXytuIPwpNeMMy50KvZNFq3UCmvl8XyE7kbMpbLKPBoqKohlVMNV2
A2DStTR4/i0YnCt0q6xlrGGKuudx+AZGRQa64tY4hsMXcME81T7oLHtqT1xcuqjb
jMKyErebU9j4V5JPWR9mcLQ3nOTD2nECuXk1Vw5FZ1BWho+kgsndTUDeFxzg8ylQ
K817fCirli/r62tOsl0T7PTuvOtuuJkzn+cke+4/8TCFOpGgddb92lv6mEhr/jZ+
NkQ0fcij5bOir4h+eqqK4bFS94yNgOfhEV3LLGV9LYQajoFFwtcO5EwhRmjjNn13
wYPaCQvhEJTK2zR8TCrQ4yz9hNjVuDKIhrJI1+cg+NRQ74tlfldZczqAnTQQgP5S
6zn4uJ/qsTiEeTHjT7GRTPZC6uXOGOhNcqjcKxcQNWP6av3mof0T6WuIu/7Jpv8b
bY9fQWa3gzlMS9INVl4Tkmx6zC63qoMRTYIEWi94DRLSDp8ubttxv3SEh4b3BnEH
eS2TPcJi14HsqArnjACwqvHrgAPEUGtTfTRTNqiLYZmvRl7YkS1V0Yc204jkYJKL
x3dY/cCwhNNoGRNGa8tmSC/a8PrZi5hxKP+Ulfic+Zxwkp7uVPu/7ekWYPP0Skyj
Wz63cACG93znjR9RNaNTm/M0HYszdnA8Ifvl4BKppMxydXeDCDIQiQOLPdrA1gqx
wdIHIEQZfgLg629c1Q2i7V7X9RysLusVmET2AaEJY5KHFbcFft1ks8j9urFUGsa8
fvxs0VjvBxKjhmxAfb//fLDNmlhtR8+jOydEKAbcaUvnhiBxw2Y5Evp5Kl5UJdzv
cIL40i8P/0hOSoBVeXPTNUflueTuziRTAJNFIFw1MsmTc8lzE/nHV8/qkaE4Ztuj
asrHdBuZrGAZ21M+GYbiYSVu0SvwyJuBQgo+TB+Shl2S+219iB+SKbrgNyFOmEgm
hJZ/5IdM5zHp4UUdsNiI1Tr7qk1GtOUBv4f+yABXLn9VK7gsBFulIKBt7nXyYQCB
hOf4v+cOFOkvVN6SSATIZj6GUUx4QtFaNzD6siFPj/x6TIk2BoUNlhVZq8pQ6UgF
K8yinzyDTej83EPgJV/vVapPMqR/BnIRxNeIStT9SOSly7SmcoHA+N5Xs2g/hzDj
vonK12hox8NhBgz6jN3gt+ffWQQAhJ0Y6MeROxJOI8lbbjxsVyddqG4D1VGwkwDW
L1YZ+LdsAUvXySSAEm7UzPS1FtM4wvmdtfQf9NSLVAkg5pggYBQTNfcqg3pd1E5+
nTh0dvBU9sXdTI+4Q0z23UY1rwFUwIbNBOXQNiwYJ1eADFfb5XBA+o228C1pTroS
wKfVUH4EscdTQUbFjDUmwk1LUJzvRm6IJ3GQ1fqrjtEYo5CDPX3TC3AQPpEQM3IW
TDUY/18k3QWfhuwqht8paMaMiUlaWNtjjf5dq9TTcH0+BEdf0BrjO1/8Vfh5uOh0
7Tv/qYcQNKjMifKl5IwinNJXHPhUwl8Qzh81nOo3bheGag7kXjsDekNU7I/GuWE3
I9EhQgmZzS8BPg+BXz962rkX3V6xxOgaszuQnjcmryMOm8OREazWaAf4UZlkKOL+
z3PpYo8aR0r1slBiHL9duxw9d7WSipkcdeXnFdtkk/vSW8KF4xCKQ+AVkogDYDgO
vsuPtQyUgXJN7/Ig3S62TNFcfpL+wnB5wQmyBZkvs+abHNb/HZUQQX8xNhVpiig5
m6lN7ri1KAeRSOqiaRoYwPiw4tEIdnlYqmDs5HPUUnbLn/deYcI4YXFrvWyhLjkY
PCD9BcpjE4qlTMaSTYtT8AV4Zdxopyo5DqNscIcpI3WSL5CEixfYqK0W6r+Acd23
7j2OzfoMSWmjMWEjTAHOufMF8W5kuLhUVgQXq36FALNvDoyvBLMe7tiknfJQ5gOW
ZVz82QY39y5WgYrUyehpNyX2AfhtTPHChtWlIsq+A3oEC8Uv/Ve+oNwitJtdXW8z
lKnTowFvEzhsQ7mf5bJrZgNvbX0LK1Xgqq8IMxEK30veFZbxTa3saxt3aGufXCMO
S5h3bvyDkpmsu7mPIm0hySTmnFyLR2dQVmGFhwSwhCNdE2zLDjXo6hpcJR7FTpTV
k0nLDwKnwQqS7zn/ZW5D6i9iUOM5uRkQftH984EaBSbMzfpXVzRGKYOXwZt/p2MT
ZcIOG50sL7FRFvfT6N36ScCS0l+Hb6HC9JpA/elLHfOgUUEG3V9lYWuUktqM1ahu
iRKfB/P1OQosZ9FVQs8VtMqDqOjEECXdujRWjLEIdzQvL3GqiIoaYzAEOGbqNYbs
hzn5uutWZxt3Io2OzdUD5u9u830S6Sx7KNP95PsZczSGhv8vL0aax31Mv2kQ44iV
G86bU67qr6sHDHBXHxhmPkQ8KQGrR1hz0FyGa4lFAk8bdzKXJCVOJWResfK/FKDO
yRiw/PvUyGaNjdqOBtkSfDCMQjSEfq11ww1xDNBiz+5ww46H7xKBZlc97Rqf0Bda
Badiua+IT+1tTDuS1tfRJ+aTnED64sjQG/BjlF5GW/JmFAJsFQPBnVDPUFO7/k9i
sWCsj4KeLD03kOtlVMdfQtq724piNAApL1N1IWPYBQuEJb1K2V1WrUk39Mz5IP4x
eKwCtpUIw9HQKGDMFLDoNLjOH82NwdXr0cKNH5u5SzR9iVtA15RysCpx2T3kQGV0
GgkI0XS1SGTcfkWm4sBQAManoOaBgttooS0nffTeZ0jgDWhI0she6ednj3VSicer
0ETP5XsbyqqxkIH3gkEZCVg77XqI+AAilwOwN5WCNgT2qfPRZsQXvSwZ0w0Yubia
E96yfKWSvAKI9yKTQ1vXpAxLynRk4F9/MatCWNOAqyS3HieKB3hyjhS35ReZfLqP
PrADVf9jUaCSOStvXGuDDON2UhB70bmAQPVno3vkErzdFZXQ9JTLtDt6840j/CBQ
ginhwP7giA/1hTjT9JNsBcd83Qo+aQA3Ok7Drv4e7cSXIBN/W8pASkd7kyeiQcCc
iQNLaqoJQA/bpdD9xiNEkWOKI/DlQjiLSxmiR0lBrxEpdUZ+i8OAUkiadxhuTwlc
KyObYz0VrmMg7vAWqaw6WDT9ATB20/pnS2Za7TkMz709weeFBGMZsLayQkl9swE1
H90RYU5AZTM8W0+9eC0bMl4Tqa6kKlg+gDuguF/qWWX1bJ/+AiHjc1fKjLGYpTqk
8kvgfAsxV3+EGcX5kxRkB66PFpmfPkhWcoWxvRXu6ZYBHwe1mZoJkO0ftxXQlI5h
eE4glnPNYXjdlTSRpgZFQXWDpOL3Jf1Jpw3OGmhMfWuw6svne68AtuVCqJG4xCsM
QOeoSbLWkxe0WuQonG2F3Z+bMQcdvxzE/rqV/W0KDNtBzpx6INN3xJHtMUMJxNeH
Uu8vVHoreK6WiatJLgiik3JkWbQlf6/wYF0O6u3+faeODNnp/4JqIzY9s1gXow+R
rXgdzgRRkvGtY6SCC4wThfQvVEUgtWWOaASySrO+rgy81JXvVZipHWMGu4XG3i9X
8CTSIvCK0XgGjAU5cWUutigkxFRJ2BbqRxxP7/JayduWM2JXHsTNXnhIqypWgP4v
hDMSc+LRtmi+Y/KTKMOQff5QB0nqX5QShm606qZvfjp5/eYuJzMbYw+dqjRxKdnJ
K/GgP4MQXWm8UJNnLsYZmpAqACBsJiBoQUp5micHMzfupJyf8CLDfMer07rn276/
/3DJbb9U5BINp/02/mlhe05MN0Iv3oGjupCTr5Hy/9ByU6HIK1cPt9CooqePlowL
oNoYNzpHa/ri06InxOmjxgx2PX0x9iWBUPJ8FnNw6LnMlek4QvrAnJQOmnieAb6N
vy6r0R6hhBiAKN8b9XFtgL64C9q5lEavIQMaaHqG86ZCvX1YKe4i3676vjBgTKXp
wPmxg4moPYVXX9nIQXx8jjM/EOaW4l5iRPzhe4kUpv2G3IvMlYDmlkHft5NOLJBd
l5JyPSBTlySdQFEuzsCqW8N6gBiACSSDs/2sjCS8MYpdTuejuUJvhAe4g8PS/6Fg
+AAr8/qNbDh06N/YbqCPw2DGeCZFrGnwR02TwvBFqoy/HnPrieT0QqGgIxSUYsB/
Mqp1VY4ic7pV9XHhE+NQaccJTgoe3+u1FZhFA6RsseryIGQdQQudhMUZ2lVK9bE5
B0ptee8ozdguXIE3CTIMKK8sjBxYnNcvZZ7tlbI0n7kC0FCjaHuelWRTgGEd3fEo
mKgoQ2K6LKJfAaw+QAZmPUiUR+s8GyUIZGHSlqLyqGc/i8O3wsN7Um8FGTLNAjjm
RW+2yC+/kC11m9AgDnRquADqeeeYz+uWloiAht74x+fa6P+id4DwU/T8e01ypKk8
hg4xCVVOtYTsVLpeA/qQbTqmrjfv0Z3rNQo/UgmODzY2Nqvesec24GDyQ3e2x8r1
RQLzUNkDJDIyT1QU51DeXMOv9Q3RBDn8O1wtkYKHEInw4XrHdUdBLTXxWVmwBnF7
acJPm/Q/wkbOUq7Gnqq43b8ASepKa/iBPNAK9WokZeQY4/tdKDynZqVbiKmKh/2n
diAb3Xp3LIWUNTnkysr1o/WMgfza9pMVR5E9X3VYNhOpNp2+HBaeZW0h4LsFcmVz
W9WbChLKbBMfIEhdcBPGYzXuWunIkDsBz+VLNWWVIpsqzvknTZ0+F5TrTcTL4fA2
dzmT+XnLhWj0xoCyo6/hNaRPtkc5dyYEvlw9XO6qjRLBvqTP+P3DF+rHm418RHxb
OvShGJXT7+jPHP7kmu9aE9+T3xD6MbUtOU5hjVfxbWHkD+c9t/GL4QoUsHA8FjIM
5c+8rxqoUpQGDHuLn2RNHRplWgfyvFCu3OWGh682F8uEhentKX0/QFKdfLLnhkrE
HEV4pKTzxcZj5K7U9NjoRy6SQ1VHBkFCJR0xfP8UAcv5Z7r4a7V6zcmM77b2lvgC
US7x0buCBzUs6MfgdR54h7JvrdbokWBYJYjeqF3hZKdCsjNx/2PraeUSpKHcGFaG
4Ybq+0MuyJf0AvyVBVsc51a0euwK9CCm3Bdn9SLdSVmG6P1NGcYwdW0fgIoi4wYs
mo/XF6KamkIbDp1t2IAbPed4URde2Fw96OJ1M+9m1/WXLIwiyhJHXF1bjpBANJ9B
pLDhcyE8yjtm437nwYoynJ9KU06gQuwO17+NOPDr6wcJDYxYYBgH8SDOPdIlsoxm
8NRilRsMs+Uk/c/LMzHTfoCGjUjSchOOmKpL5SB/0l1Ksi/4yziNLpPwfcx4yBJY
uc/oo43Xky5zf2o1uW3GeArWfYs5huKvfNzjlXeWyA06WKQgHWtZQRD6pDvZP5Dd
5i2AabCJbR/uhZWljLy9/BHDYmEezdoJpqHYCtq+p71316Ndvzd1CgVkeWqHhriB
Mk9CSz3j7ig1j9mk01q+xkmIRJFeqjwaYHPEZjXTfMpdhGZS1H9m1cA4mn4usrpQ
SAZbaKTV799J5ExnvmeNIF5PUJL5SnJYDqbPO2zS4BXl480wsWp6UX9kODNiWx6W
IQJp/h66Rd1o+xAxZYWCEYCUqSyfTuDjUUdxLuisEpPsTKIYeVn7prlsNgNCNfKv
4naqc6yySyaYKj0rgE+jwIKu83DuZpPSQy5403Or0M6r/0DBiEMgxVJcl/iEkun1
lNsKLpAHsniu2mVbItCVx6KFuEsMdFbL6owXCOdP86C2GR4CA+9BApBASbKWTQFz
M3Wdpwfea58/PFad9nG9FOSwNs2jArjXapL+cHQNZfqjkkhDozUYNPezCC+wj34b
pDBLCsbijJxn4NThm6msE8q2CaE7GyhZyA0K1sx6CJXlJwVdTzqL9VrgSJGs7Uzu
HJGbgU4ibX7fMOCov8HrnpXLlP6EHQGfmxwwu3ccsSGYyHrz9+6dEvQIPNNRhDdW
/9EENMv11IqEn+XFyWW5Ewh9geBQ3g9lSTlN7JYKD8WSI+6jIA3RUBWZ7t/r4k0l
Dmv4VoU7SVdmkxgS6kDd5/iFgy3P5JTUQAWKv1iZNuJpgGVOIxcIMyRXzdU71JaA
x8pYAONSbmf81gRzvPf872oQGpZ60KD5Puitj9u5Uhe6rEXgu6UNbjtGLm3v+9g2
2SgNTEzm3jsKTIZOe6lBpY9fiNqVVFbc6pmWsXcfU3lhlZZYk6Q/+W6YfmzocFUl
BxlFODn0hJiNzd/6hwNdJX4980TmPOQObbWo2iZlg/Tn+fKvDolA1vdwR9jN4rMp
j+gRtbU07J/6rEITbfUYJrHwFd5yDwj+M1aKGLgyZPO2eU2Q7yFP6kc1yiDx6Xat
1cKkWAzaNZtKK1kN81tS9M2saT4lR++vo2PSJHrwaTSQxBYUSMFZuI0uCfGaZd3v
edCASVFwA3Ox8BVhL2KZgcy87HV05Kd/hn1UKX8DyB2/F/AfE5dCzjUS/aPo3wPz
svQhH5+zuzUaktJhTjKoOJj9sdKZ/2IkIv4+bqzvZ9SpKNRtoVjTvE2DW/nwLjPv
rbQdgnDvGegFB3wJ+pYCbiOtBeLMmK6TyNnjSQSecn75eKDmmYJcqczy/F01Zl9N
qn2djWhKxkeRuJjU7BnwuZXcR3CNH87/P5+rsfMCHqF9hXDnwlQr6hpGjqb+opRN
RtwSidPTPJHVbiXtjIpCbwwOHkK6A8/w5NbN/wdChihVJML5BBFcewR/8WpoAy3k
ShVE3QNc6iNfvVBJItcpx/bhsS3iBFmpApuVv7X6WeOVEnmwHt3dodfeFmv92auW
TtJ6WwZBw1OGRtjlgnGWkmirlxlc3RZVHtO2UEwk05QImFsr9j8O9Qm0eMxYzVGi
eHTVQwMqx27QWPlq4SSdfjSBEB4vv4ouep3FpjMD0gjP289gB8gBrvNSRlzScoTA
25wnREAp5lH7BgUN15X5T8KPbFgG+OwXhKPD/0JerGu+0aiNIKuCqDckwPSX4TYs
S2p60zqA8Gzj8FQiC3jFBEdgWFP8aX232wrbaTWUOd4L1wKGDU5wUXUT9e7r6PHu
7ptnrj6tkFBDHPjirtXvL/3onon0igHQmhnnTvml+kLdMIXbzs1ZG/cFnWYVMMRd
CT/6R/gkaaUed3DbvU/tXWPH61A5dUOG7PC3pNlnr+Fhi+mcACFdw5s86Pq2JwYE
t36png9KSqPHh1riB0DB58fDy1q7UD2dvVxN4ZQCW6frYOwxAVJTXNC31vhqcMBE
gQLLSoFjjvpCQp7ZizjyKyvq7ALkaWbEgQ7OCMrVk6TRz5hW2NcaBXSJID9wYP8v
muAgww9EiE4a2cif8nMuCm6KW6McsFAMFyUwjOpWJC7MO9OCqYjZSEtKV/u3aP9D
8A7FBYsGGJLBZcK37txNWpLYF+1mMVhhUiBcQlIQyjVhRv5ROSZjw+aUelHEpGQE
LMVWzTsGeOqRbRNpdnspaFObOxVJXNYvf8xZ6Zb4ZPcxEhrcrGJ5W78BOLS3NHxQ
E0u0sPUe2GvZFBM/Ap4tw+ZZnfO0QzmFMHDPJXi2O3KT3eZSKOukcR+AzYw5QybP
tKWN3r36rgsHgayrwdut36rIHFZ7bTu7odZgFjuvT6rmGuAdmDCV4hRV3XrdEq6I
Lqto4gkXLNKHxb1NnnUd5VCZPjG6V2bDAz1r4pCg2BfaASOaPhINZZ0WxjlOdMOe
1NfZ1pJ+xR/2msrUnlLJo3WJG3XZxDXwKZhYLdf58guD1BHOFXpGHgef5kmBOYHX
bBAu5aeZArh43+Xn+AMTbeg5B0oCC0n9UXuKFMfgx0ff+F4W46hW9HO7RF52sjjd
WvumMWhgwpeLF/5R+nfG4XGhFZ58Wsi5grwHgXK5ojRRMUfp1R3XkOOWvI8yCdzd
7KE742dgXrQh70O7dlJqNZZpSrp0k2mXEDEbLFMTDo6l7SpdR8jS+fj5lVa3mIvD
9wBVGZ2bi2vXWyPy7bI+0TE4ucu9XfkdmNuGIpVinEAck8+8lPHomvCh9A50Ykms
JYxKVT5EgxeKDFih0gBbpmPaBzf+aO13nfLWDOplTCz0sg7hcv1r4zITSyoab3js
O9yh2pEu+7NLO5fpMCNB7JjFJpHjsDStHDJG41DZ69ScuLG7lwuDh0cXdWRjjhxT
FnaYYE8irXp1itEbZdEUdIN189qklMKszZk89HCYYiwzjUV76aMLKKaVb07tOC9M
5ZwSd4dGWHCf5/N2o8hmaj4qmhTjNYHOdIevc6PsfVlLjauMA+aLsW8okRH+2IWW
33mRXbakw/P2EU/3yA37yfgPDPmPi8abwm72kJrQlazCBopq8XGlvrBGOY9nq7mq
EavCxUTkSDqt9TT4LnKPHa8RF8AeKZ7mXT8R65/hnz+dAXax2DSQ//oQtAO5wdsb
cf31OPnQzuaU3CnGl9b4BGJ2yw3lTTe4CTTsfzUXczRkS71dolMrM/x48qWVzOr7
hZ33eepxoy7rQVJuTPqbw/50T43R532b4G8yAIqXrFFUfNLwrABCcFIPy8zrfy6g
81glhCVFnvQMtSSOnwb3VDaCM4MmhF5LX2JCTKZeCeMJOKOfw6QcE7m7K2gepnCb
hxs8LWuUvX4I3Jinihc6rSIXu/ldO0rt1R2DVxTb57frX022ehOjaFmudtYOVl9J
YajeLikDl/tI6zRSbl31XJ2/WeISSmUaIeX3m6qZ/Mpi4eVPc3MoavAlugj8Z07E
iHWh72ioivletXmRIqX5UrRjasy1uQbJdcnBS2R6LjB/2HoUnppMvcFxH9fhALC4
gQxzxmMMWzKVKMzP+f0axddPBulACz94pZnlU3Y/3nIGZnoFUKFg+VDQsHGfXkRz
41yUdhcv2hhCyYAU9IzTbUvkZ1PNwtnt6e/kLheD27W8ZaBcNaIT4W5fAbh75Rok
5Tkk87ER8O0kmx5EOCuHyVZso+Wn37eQpk4Tsxs+XuWUGOdlqKU3YU1zvaQUoU51
xYwLLzF50TfC1sV/rfr8qY0OBWqY9m2EvPLc9SzLcU0S9DPqPw4y0QCXVdFbVLoc
hW6lHHTfn/orjfXDIQhQNvxWMy1G/gYcfi7BoswaOVvMATNtR1n8bxrAbxdaH7t9
HvSL/6Flon8KT3a4ebEa6zjO8mBdC4pECbgqhHAzIyg/eTsDL86jc0gPewSymMI3
Z8mldzcVjuPS6zCDl/qT19bTS2Jbpjo9Qep1BDgV+13LjiGPggCoCgCODiR/o8u+
5y4BiaMNYvdsbkswR8GZdg9n6HPwRdvcwuoamRiLi6cAXrr139h0TMy8CTtcCX4f
Gg4uDMqnZ8RkKpb8P5m1vW84aXf99jRJKoqlZNv9HOC6JkuQTqEBKC7R6htUp/0x
WFaqSdeWmVc80mmjsRiaoRjnrA47kj7L4kbbG8S6GkDTdwBBxkjJWaN7gYb2NM4I
EfkKRDaCs2xxU/UcjppFkUsRZoqnR5OjTozK4920ehqA57Jp8n1jZpn9broPFfwT
eBOUpytpgPXyqO65GMexv0frFq6+4Vc5vKMpJcZsFLsWUjqi1rkwM71UmogEG6cu
vSzpPsZsWBBf2HpUltrMfJwDb1QQkzYwjWYjTWQSr6qBtgZLeZPuHgSlnRnhQ5er
JAv8rbeyRrUbWrH0GfJ/Dysi24A9CBZNWPlzrgSKgZXE9DvbwDRbcgkyTQrr/+6r
B+GWH2SdeejZDbRi0y5LZvbMZs8WYlBMm04YvQVI2aiVzlw6mdWN3nOHOMUgAb8W
f1d8bS9I9kCwA1K41IJijWgU85NqeQh0pADHvMuQ7lWR2LRg8AQlCZBJR/2cTkkh
xopnCrI+VuFsdLfjstTQBF59lDXzZ6lUYqKW0B7LetKd5w12HTyG4XNZvJWf/hq9
Ls40P4LmYLaHNlXKDvkVW4O7vdIhQUaaZ4o6XSKKMDwduq1CE6WBOczYKm5p/BQh
cj5lr3UHU17kLNMv482ZdpkyRfeNs8+gdYmXNa9H+YB/r25yHSTi1OJY7yo7geXT
SBrifNf0wExMjeO9wVGLDAkzucWnkN43TCk86iTrhIACYE+11ctlrcGvDWKGdLT/
ooP+STNRHYTfhwBhPBQu3/aiEQHtYWOOFApB7Kjj123mcy87VAvryNHyhJuqoluu
gv0gnEHeTO0w8kKStugNFg3e7B+x8bXP5jR9X64HkPc9nYseEd/n5GW+adcRqNtw
Z1g/uTOzO2e/tE+GVUDKoVtPIXho5F6Rje/BxvlnKzPEJTBKWUUdiEtNjcTxLi2q
bPP6d5RbiEPdLGFfOAjxnsnjqE7zAQt4vi70+gxFHbiWD/G86/WoW1pZbyWth5b4
Ltm6XZnkfGdC7LsOoAp9a1F1Q5JmEempVjx96mhmT0DngEwCucJCKVSBVEeQcjGd
aonUx747+ll96X2v6D2fIWsV9eH/H4G/1ZV3whd2vA2lEn8I7uxU4Wn9jYEykreU
zSWwW83Acxr0YljDYMuvJ+VDfZhC7UEWk7NHRQJ0ua+4BNVZL6D3nABCh5pdRPV7
VoamyzgDlAjrwJJFuTK/SqfHdGgjbzATpq8q0WpYdKtud9CZhKFH8ZVNNZTFWlcx
XK3i7ucprr/fRdePV4RLvjxj5UiTMcu1E+UzN1wiDkBBaqqSW8LWv4ek1xPz8f4O
lSF65DsvgLR30k+9sE1xGPfSDGYMzrG9VthH0KA0cmlcdW7ttQOF3gruiAXDUdIZ
0dgKX2cB4iuc+HgzKoITMYYGDFTwfN9h5A/IB2NP9rC/rJ4AlyhvsZnOgs7OczeH
gteIbo7eRbQe3gcK1z5m/Y69B4S0vmUCS1Vz/zEg40yIDrDGWppa6xh2bjEUYV6Q
6gBDPbZQsWXrKMkK1YtpvGLIcZPAOQWAMM10K5F7n9yE8ZTeTLGOs6v1rZSSZj8n
VbZ+azDr5e/dAkL+T+ckVea/SEopmCifb6wOcV9mIP302wemYrcNjVQ7Npd/L5Xw
/ieOpvA4oNpL6ULo7/dpcLdHSb2r9HqoriqIsR7LunJErrRGuKtCHZWx8Keb4QAL
K4YN9dEB3NVfrjB84ybbF9jMZcC+CbgTg6HwBlTasJgNwSjC5MNrpxiQuEVu0I8x
nBB9X78jUco1pcClqXe61S1gawMeRX63YYdz2TSgwM/Ya6Rgwh7o+NEyQUQ+f8hl
l9r+dsEFTqk3pz3jTqR4N3FR1j/j9kQuntXkNQjM7E7lCuL7lDobE1dK/U0aKtnt
ePt5OykdMxJ9Exvq7yMWTK/1X0FEUfC0n7VUBOm3krwDhFmI15u5YCD6fwzVdTyC
ahl5YQT/m12mQW+xfCz5VGPqy8uoua+bC5iob55O3P62s2l2Vo94so2inNtXNfEv
mag2fOMSf7cO2/hbfY6OvlbNMX1utmlUQ+3tWS9s71ucl2V2twqkchm7CCBJraEP
0pVbmBv2SVAyl0axVl19s0VAFT9eEMXk6KpGvP/829tj4CNIq12rzlTz/72ZqOfD
Xbna4l7tiHq+IksnnGWruefPauMijTPPt4T9fz0/3qRkoWb2Xq7nZYavZcC2AkUM
ZcF16tB5vJSitEjD0fiTVazmdn8JQe+IuLJ0w1woxfJWr54fwcN0PxwFOfkodQnq
5WoGUaKrH3UPaNe8/bFbPxyC+dmA1NCWvu+g8rJRAc0rXwlFoWnpH3aIcH+aBfpN
I3Z4eKZfEclkE+xIO4s59EJ1hNRRRNBQ5ItCPmSe2mT1+OC7CSGLOTFkoc7uSgy9
S1tIqHhEY2EISCCPkdTw0FczylgP977Zf5b+sem0H6rDNcCoygC7Z/cJeM+4KTZP
EaPaoAqnUq+LE+6dI/LLYF1zGy2s6S9fZgreWLc6TKOpnFGQXbu87R/kejlYI3vj
veNZVUYGTQ5wVQdNTz7s85vW6b2vSJEao9tuApVvxhJAy4xgmCqXmUtqumfbog9m
L1DQigXj3C6Z/xuLrBpYXrMPTWNMPLUtoAwsxsmQu4dUpIK+1Tm1LuN81X8icRDh
0jj95jfjpfamJp83VwHAlwkbcDa+XMKi2ZBLIO/0aY57020FEm/G5Sf7bjc/8txd
gPoQl36+ULaFYvbOWT4hh1Mw3ymZaAvK0WuaEGylkHyFlHWwpq/bHZ3i8E7jRGMT
pHCQFbhsMicAsQbx8B+ek92fASwidBVpfQqg/ES1wfZO0KHahleA3MvsEJK/m0OX
MeOp146uLqqLkHDThk8NedhOR+BUtkMILnGZKVyTmql7l+smRlLjAeiVM9igSkwR
lcyNnDZ00q6+7GLr93we+WMzufWgrTTDmROGg+cIqin7aV3t51dkLIr+qJWaga20
MlCPGfSQUHGR5DZzMKdvibfSXZjNLTIuWsrygX5lamhhVB4lhITv4Tr/1N193ZB2
bD7B+lFEJk+tM8Q4g5QjgnUMLU1MBNL1VZvwS3qzbWdIFjSIkAbxikfbXtegc976
dlSbiyVEY1k7Nwkl7usxbdwyv5yW88BWxXMYif/7vv6VqrjzFaiftf/fmlpCwxzi
ezDYl4UFmJc6xovA2qQ+Pi1hGDQeVLO4LWj9+UXkA+Oxbfv8Ki1PLu9pUsnDsaTO
9gQL4N+1irYCDy+3lDWVgwesEDhXOP3rXqjQQjt10Dp6YGNQiEHpKMYhtcXgq+aO
xcARwNmopZJMUL2l9vYhKu2Hq22PetWFdYadnZGyivAy9W8uRGsgwaHGwxm1t0XT
fYghJV1/YxgypouK86NLwJmBDfVqZIYSH5eW1f2VDVsPWjn9l5I4UvmH4F5pzU5Q
v2Pw+p2yHNCikb6ufec+888agp+6HkZTMvfFnfVxq1t/vPxL1ie/KrLWqDCthNR3
yat0sYaah9des1gTeqWn0ssi9noHFgZPBdSuysZ8pyexBORfiS0PbQCTmy3fXFTT
blwWNaUA/E3UXST4EOSyzvj87Tmy9VseQDKedziqu9L5wfz6YRuE/Q/oEe2Oa0Vd
VYmOIMzWOzJv2QJJ8sWov/rNlah2FXTbiC+FxHlVwnJOjQtGZp/XBp9+ykXyLgAC
iTtNXf1mSFy1+wQ1JOVon+aX5AWk9TRD0GMBuA11p0lzNrYv4gFVswjwz3fEfHYj
i5wbti9ppVlI0AvJiqlQmDpiAs7fL+NaNekmm6MvzaHAH/iAysohIsTuq8FMOnYL
vf3EasSQWTun+oYqmD/LO7S7ILzwmwMcXYA4a0NSkHuQy64Ed83Nuipu9aHZaCTv
dTaQ30aL+r6z0xVJTM/ueoQB3uP+jX4fR0AE78sLys28v34xunAB38ALfCil3heV
CHX0i2bOdmkq9bnxIlJa6jH4c5W88HBAzwIC4Au5Uhb7OELt3D9oagv3hBFyMGRA
rj5kZv/Va5J360aWGlsogP8gJAFdSmv7F4TgGaQldLmIICsafbsDU2wAUoDmv8lF
VFQv2ERlLxzyk8dE58+h4RL9mWMHZR6pYaIhlelSObh0Ii8yFvPRf0qw5gvaQW33
d98owIi1+m+iXvx+v8SxKlcjhlieZHx8cGHtmJ/HU36qBvvu0stjhR4YBouo7myf
J1HLNuHSAMFzWc9uKKMECUkjy707zTuba1a9NQWVevcWenjDbHKoZbceScQbK9Re
WIC7p6UjG2nvLScZyM2YWBj5QdvwHcqO3bTE4RyGgAL04oFfeMvmVtMzDJVzdub1
am9SE3UASUacxeMpymlM482DWwB4mlY9rkjINn360RXV00qLjqZFkKM70DHdiCya
oThVFGEBqYJ5JwtOcv6OzYlm4g5uFqCM4bboXtwKhg7TA+L1VX+XiGhekRFzN/1Y
t5VHWsr1sd0QS7pppti7JwmlwybnoA3q0aa/5vJTY+tCOvb//5XuPHnvsEz7XE0u
lUwx8O/zCNEGohuSU3q/FPC5WjVmsI8Jp6+YuWGHR8b9XAXCAQKiSemDryrVXH7M
OOoDOqrfj9c2q++Jjf/9Ls4ecaa5/ZCBsdqKPjEmXM4lLYxKnjz+8VVyJFH/mOfj
D5h9odmTkzpE+BN298VbTm/SP8HR6I98cIJnFy1JBwVcUtpos0QWelpGQ3aQV0tG
AhARgivP6jAw6I21adrp66kMUGOuDqgkGP3CnctyfbWcQR1lbPXlDoi6DV7zYhBX
svBkj9Myq2VDlciaqU9x8IZMd6zhQoYl1ifKg2a+dGr7pj5zEandT07bd4pkPpOu
MuQAo7eV9muSGM9t5YPMud8JOuefi9dew/AAD82NVBibXtJSINNfTY2BkhSM84Z3
AN6ko9on8y5D1a/YwdaWEsKDqy4/hpnJBA/zhbDK/kBB+4xSJeHdAibrUC8XR+o+
TUXmojkMe8g2pKLGMfZPQDIdiHIyRUYRita262+yFEiOoBuaGoK1htbik94/BXyV
4UBD/baajA4otD++XuQqbs1f0YWlgav4A+C82WMpSHAi77F5CEVMA9nkysGlHPR2
qpunDj2uteB/jYNln0h9e45wUADf0DsGpACyF+w5s5xt1pdKpI0wMw1h9I1/nubT
2Cw3X0jGGdSoJ6DJuCbWiXP71YZIFnrXQvKyd8Zk9Z1dIA7spLLB1p4SUpD8i2YD
Yi4MGj0bp/CMOKEFbz30TqQMuaKkcU/8lg1GBZV596i9TzFD01quJc7VveCOP/iE
fC+hNMd7ulAq2wttySuIfIA+5jWP8tCRo83KHSpHAcNKLIIV6aew0fuxq1VHo0gN
qV2QIMEgLjiBkTCZmYfAQLxo5MmsbjrUGlnKf6K1gNC8D7GRNEDvpduksHh+RtFX
IATLNYgseWyIu3ldn+kwHN6h9S83HtYq71vaS80Jzo7lJrMvHO/j6HImNEgr5DOX
MWIOIQjCx7ybvp53Gfh5ZmRePNp+XXFoXeXnd5hzdCpyw6dfj9QMFX7RGEbSRYkD
RPyNR90XFPEUO+wgdayl9x0MMeLgn3bngMuuyUPLTLJyEt4A81ZNj42IqnYxhPcf
tpfVaaqjTUbEE2z83KxxOORh8cZnkTCfNQVQ8Nx+H+Kf13D+3ny5vWHH2qrrw0Oe
mzp97GiYCgZbR/orEzGHtYu7yH+/qQ5HnqvJxSKtR8ohDAUxpLtJG5tIDJcK7zKD
7eUJ0cR4uJuomp3ZO1XTEI8+R/eQkU7GEHwjtmKpdvO1l16FkNX4rxh0LLzwCdFR
iYKppStv/tVKErenbdYN45awJBgIP+iAyJowEruSuHSqUPjX/SGVaqGVsnCxWy8z
rjcFmaR0vPavrQKEPYWegrdpq2jZLg4CB1IiGM/qoe5HExGYFog01Hh62cR+wBU0
jAo5KGpoL+U30eSVX0jcFFeI0q9EE744wpZVBxFYGH3MPhVOXUm6xLbpM2Pn1pFR
+TfNvENSHcLwWRozBbVhk2C34ojLlbKov+bcCRh9CFH8HI1hGiD37tFYWLIOSyXB
ws5w0qxYHIm6BnSFU0AlTJGFV3KK8D1DF/sbLUe7nbQsetn2e55hNETOKZMBQBQW
pn0klOcHmoby+vz2WuPXz4Z/xv+mwlxIsnPZNEPJEz7c+sHA/xhzoS6JDhhg/tIS
vX8ob0frvTliELBaEwamt+1NajE2twPdXsL4G6ExW1csGdbiEYURKIb925A4QPCY
WpxgHSKy/xTKmBCPtatJt+leSuGvY5PiYGNKYop4nyXKSzvX7iBJiqqLTKX4PpPw
RiCoSMJWBzpLY4a2ng11S3Tw5f1Wr5hSRWTcEwn60KrSaau6xqj18TovOa0s0Hon
rBaSntSPfS2dYDyglbJWRfDsp38k7D9aPooJRDr/MV1TK7oQzJlqPnTGqe+RStS4
uN3cwAEE6lTFkIaRBTyBVul27cTcc+LNvhoEtPmudGwILuJyDBA6STrpvxAFrH9K
8OAma5ol8enqveC77uVCgZDulaDGwK7nwfD7CQTUNQs1iItTmaUHPslUgn/WgDzg
++/D/t1zLEaq3cpl/S+QeUJrV/rqmt3wNlomID/jMoJcApYotaslKYXkqdCM+alO
fAYEhNVtv3UPa/aBtB8tHdwC8ccAyYfaGFx/13aQm7AGTfhwTit8xoL8fSiuRG5Z
rn4Vt5y6+5wBc8gj1ZfHJzUNo4du73dTpZ8SJBU10LzGnSvTsgdd5/xyOMu1+zlB
hi7sggl/mjFXlESrVIBnmAP7n5Cyu8KulO6b7pmegbgzGliEWfCKFQdp8HOXp553
QQMGul/bRQPOH52koNcyzsJV0JRLD25VNpkv5dMO1WDtCUWidcaGYuCwthXw8Lgi
a+TPPGBGYhFsbkqVtiI1zqMRYU/8T78NmkIPGF/66G/P3nN+zayo76CKp1d8Y3AY
96juziIi//ghr88RxLWPGtBXUBzG4HJ/W79PQn9+WwXX9fTJRSmwn2hsdTiT/CIT
ufIgO2I30e9dwuH522YcycYb0VTxmcH2fxuItkfeWBuHR5Ft37os1oOnpALLf4ob
EUKJKzztoIQah0XqY6mSmRPLItnguUsVfnsvHx989SJIq20iqTyOSCyg0fbpNuB/
uWknNcTF+MyBhorNWQgnEJWQl1veMgPQZatbkPgGRqqXGN8jXEhq30MPZT8/jV9+
+9+HMU4+vHI2UKbcjL8TkMcZ3rWh9m1xPhdXzHDpTO/6Y2ajs/Odv/kEJ139RAom
+3N1SI6XPZVNPV9Pk4n8D8G/nTEjS8ntbOBJpNtB2FXbWf5qvswgyl/VowbQyhYq
dVuDIyKOFkUF+B6lTsLx4huFfQpxLOMg1YEgHwfQHdq1Xd7cO7m/RN1y3IbUiRGv
2nMUOK6jD/dPgOq2DmHV89usxbyXtzdVMGrc1j6iAeHR/oYU/jWKnIj0GKMYpxdC
HByp6p8dbpILhD12avyCyf+Jo4r+Jb1ufzXVB828jH79FoHiujJlKXq7kshDrmOC
1KJ8yOyNbABMBpV/vpvBG96YnOpOaQOe0McAEQa8lTbSeHtS0Af+b3Tuf9qdq2wX
qKqw/+kHlB8l7HWlQQkNRneGC7i8XoRELZZXG3xiJL9kxUJeku/Zxh6OXQPxoMSu
bpUdpOjLguxiizNuhI0AtFBCQT0o9x/sgLoH7QKyxwfmyUZooYCwMNhT+XcRg4BQ
XU+uUtvbX3sGBbk9TW9LyxiZZK0qXFCcKv2bOM2cytE6Y69R20wstau6LByYixJH
lZDf2+MdTU1Vg8Mosxt6gM4TpPvKHGMHFSZFbgZ2ulZq1felZ+OyHw6v6A36k6zp
FcVFMYEUOSGX3pcwdgNZCAQaVE7yk7CJXMiMM87fryOvVvDfjc1/bIo7Z3uOp0wW
l7o8NKE3mP/2JmIHOD8nI4BCCda1x/5/K2msmr7qKDAVilZ7R5ZjDfoPiaT1dGsP
jb4pnRfzIIGO+oTfD2GHCE5Rpzn5dL8dgUn5qpdRzZK1ebfJAfBP14OzmPPMKYvT
TmNAREY6utGgcJ8cSJxgnVxqcuDib+sZDnC5aSRjMIEjQDpdz55cHbMA4D/sHRnV
+opcxOdoaCy3ixJJWton7EeQBFIsPob0TsbOxOeweQMcGZsATzWwn+1phCVFqcw9
uTq2g0kGJNuMJNLjE4aORtRsiYysCXWXYoE9KNfunrB2tTXLK2pCPCaHvXC/m0q4
Q/Yx1Iqls+cfAxj4u8okKcaN4Km4PocuyLVlef6ReNRIJbosWhvpqmyGV5lgwxGa
AlSULCRWuzw5ZtNDblkMW+CvlI+UyMsKdYLoWltG2pz0R+rAiZHRn5RncY5OHJvv
AgZymi+QM2QpHHH8EkQRV1snqNtoObdH1JQVwhV5MD1c5GAm0GLm672YlqKziqQq
90OhNIzc7jxgOoDF1UEP+gt/cIPzQo3hrfM9UgNyhoJ8/NzFuSCBZjPV7SthyP2x
qoNbumY//OnR2EWH3T/qMl+aLIRtjcOn6d413CIaBthceiIGDNQ//NbH0QHb/uje
Nh468PjNu3hfOYOxlDd9O5GJObDOk6MhK3LHy1EWLfW95di5pXKArHzLKukAJudX
MjyvI6MdI9B466g4evkP/ffoQxfXw/g8NvyRhoOX65p4WLiyUvQyc/vz9fF6Dr/j
HR5kPxwdpdIYlj92Z/SW2C0lW0SYm1yd+zmx3QvhOA+cZCcToDvi38xsrXDhjhX2
utbmH/bbwqKY323c4ohrDlUbQBkvt6M+wLy8b8Ztu2eBblGXLK2SG9EyatMIYjl/
xSIBmiu0zyadjpVECPG1mDbQFlha1yJlVqW3vUbe5CB9xlV7081UjIqM0eZ5QByr
UujBA8yzjeKnKzTkRcO55pqLz4m8Q3iJapjh/LHSK8wYUcC3VX1E2xGOA9YNZv/W
p1HBgdHvjwhzuxYALDZHZ5Rd2CSlkRktO5NTRc3aSI4Qz447uL3D11/jkZUeT64B
rQ2Rqeb1WfdPMSERe6u5AfsA6PWvts/CaSmdZ7mf5OeAH8uUJ2NzBTz8QirWuyaT
IwIR9eQA3GCEWx9sd6I1/g1fqg1XvBZsTgtVIvEkWUmVODjRYN9Y/AeuJrEsMism
TsvzhD/KkiQbBmkkm4QmXvSRkGv+yIK9563wBTZcunE/mBFYhk5o0UQz/9KgWv6U
gDtD40CrE4xpynTBOue3AQtz6iq/4bC2424XfGhRa8ojV5KsAPdJScgm01MdItSl
fqbmhD26D9YDGKglKow7ICqkTw41hsgzsHDMh/7ZWm3C/KWrW2v/R3Jm+f4NFuvN
dpGsjS+0o0VO1xazQ0+T6tXZpBBYXF+ZOcJJNhnug/Q45SJ9W+lBdgQI2fPEErwD
yE5ZZSWYuQ7BB76IpEg5BPDPeTK/ni/iT5hmsQrk3uTwAS/ViI78EW2+YoKn+ejD
6zcBSW88zAoCFYPRWJzB1R+IROe9BLJcTxpWUJ/PKL2aU9RNINKaQzeu1MCZ9bkF
r2etsceeqGwY524Ezf3EQyWHcIJiGE9+NbYk9AlJrTXaa39ROWtzaGZX7WrLe+nG
x02uzdFK7S6LlTtUvSjvx3xbufOod9mrVAW3/yZKJHs26qjmPHBc1dnMWr7EA/BJ
VmHcB3x76VAFjWgWPHzZ6Yu787DxO9tqPa6OSt3BahhtsTvwIcMIvgzUVA30jJqy
EBtRqcc7ZqvrPN59ME06MTPsms9kl9sHEGiXeMxBIyFCCoEYsKmNCIkV4RCAyaGr
9DavdQ4Fe6VJTZubNJaHTWA5ukJETPvn1BkOrqvASdFVBoBXnIM5L9gxQ2dm3Igk
K5Nwu4kgsNRTDqnLXwmcq8QZvsXicM1xwq+ZzS1ukJ8h9LHpeqWOPHXQTGPBt4It
S1NMsAUrnOPYg1YmAb5jj4XceJNS49xJgdIcMO+J3LqU05DXCSMsFxUmvvFwzFjR
jRCI5pH6EtBHjZqInP7SEvZTKNFX/TOW47vrVEia+o1nUur5YKWEbgbS7wE5yIim
fh06RzCRzfzq6pCoP7ZljcqDhyYZTi/ni1VoPUGi2V2V1IN/JT6GLw7DOSp08rlu
M7XGZTxRerrE4alXQmSRD7nkhcWKS+z/wGj62E9/2RHMu4MeL5BdJygLkoKgQIY0
sJ1S2D0kqBuVbVk0yEn42Hxk2nmyMB/7IofQY9J8DDvxdskUcYABXMy+vQ+HI8di
XiJWc3YMR/3cdzytmdJxTpjzd5SL78duYBZpX4tAb4VLgg/UpgpsRAC6ZOgRIYin
P43xELEkSWUz7eb5q4vtGNjFHzP29yVhJ1ZnCTVNQdtC3XXA0++pSxX1J4A3imLS
hKdOwhjWFfdPEVY7CQy2/IdYv2JO77Gyx4G9JZL8XjMWlHit6LdoL72KgV9kQxQz
KlI5ZtxiYSsiCvZQNR60rrErSEbGgzls5Cc5gatl76tsAP/+6SzaQ/GCTzAwohGb
886yukiSLS21gs2IRInxt1YHtTDTPKA4RQAfsxnl//+MUwgqMBxQiR6yB46+I0vK
DGSCq4jY5tNhCYoQUjUesjxAPLQdZ9j5EFQHOlWRVgsXIr/Mlfrx7LwJJO3X3WAh
tH4xdIzJ9LN3NTEl6odFiOuFxkX1UmhDloZPfJpAWtn805Zq4dzx/DNhlf3PDGwP
PxQEi+ikralzx+QF+sNlrfywgc6HsyRWBmFUrdl11TCceuZUvYk1ihmI6DsTKejO
Rl4gd2r6UosYqw2gs/6UpJlTLaoZBugsbnYGrLhxGUw0fX1LeejmQX9CjM9ZvpKm
2TUzstgpz6r/SviM5oFIv5+uniUOwSQhmHCfp23iEZmTj4SR/YmDusLtEK16ENav
kBEI9HTPk9Gw5jRovAGiKQHV60Ee3DB5+fkJKj0x2xtgi69kBB0HvQw3Z6QkD7Th
wIn5xuZY6Xo4m5FTELWAUX4+2b+/Smzr9Ln7YYKs02AnUeQ1M6Tqm6fq5xJugf16
vtqAN6kuufclH2Y49ZVKXDOUIAVdNvBpjjiAACrLoDXWn53HekvvzBFwNhwO2eOF
r8n2LIMLn8kBfvZ+EGWmmbGJ6nXXNObb1DuwTri9vcpX3UfdAwX07GshrnGVuRPm
Y9xthc6bwREEf8Y2gPoGBo9CmtSdzQ3o2bzFhiGzv2A86r/2bIYekvXYjE47WX8o
XtjY38FXuCGKIfmrdsAirmy7Gm5ERXTCr7JH72UxtcorPyzfaHHX6SfE4AZNpGiO
9WGbTtVGB4Cf8i1DgxSX3+AI2+G4C9dva6E6fctqO1GLWfIEwXWvzTEmm5l5E9A1
9irRV4fCJr6EiP6dxSCAkDR7EPs4rKgWns1bwY1+/uixPNeVJl+rhRasjpg2ZG2f
ZQA9vEiG2GknP8/iks/undMCrxBVjjP36L+FCwdonOhb6NlmIpkAZgofcUsrfqAT
f0V70O5r1Pc7qIzrsKk1gZ42d2dDTOyZhI+R5ZElWX+yUWJGGoSl04IQl/hBkXCr
IzYLyPqD6jZkPQdjZqShbNUzPTMUPUCSbrdULdZjvAaAMPJfOioZ9G9MY3lLA10T
UVVcFlV6WgbMsj/mpaIV3Vy5poi2XlkrJQjwxNSfUHpyTMFWtdfD3CclBgFu67jJ
n+Gg4z59ItCP2SYIR1YNH/L3TrMcxd0XeVJIhbgUzDr4SlfvKm1sMhHdVPURj/Qb
0GC7py6H0gKxJcC+Y6YfWriqfiGgVuRaf+62ruxgm7npvWTBffE2Gjw0KM+dOm8f
EZ9lnzI4JVOpzDIqimVaOl5fp4p67VwXCANxjB31/GO4yjh8PsdjBNzw/55DotZh
cKDm5u/bCx+DlYNbGuEZQvFwmG6e9XRb/CJ6OaveuNZsdgu5qOFVy7dK3GtzDzub
fbIyVPQ/rPmnW67F0DlYSFN7+xEr+58BUcWZdo4nu9y9T+UVwmk4sR44YnS/qGyU
XQKSI6HKjhhIg7X6GavSjUEtT0mHJ8xvsMx5qw0Pnnmv0eBHPD3nvbVAenSNN54y
D4tTFjEO6ZyzZVBGapSQupSgrWJc2A8l3R5sQeWuGcAEmbWfJ0yvTv+5v4Isyjto
2goahchJblloVAOiVdW0uhc/GcOhaeMAl7cPL4omSyZu0ma+MibQgMdYUkXrejz/
O26LXPNHTNxBL2KlzebvPYHYyHVjw97CiEnHIJ9zLBS9SU7M1bWOI4irCK2D9+Cj
6UEa9UTGxZ+sdCKOpaseQ/gZURK2AfYm8myo1g4FagyDM5BUgL2ZX8fnul91m58X
fBbYsglmh/478M/s4z+fxUuCJhan/YD79yeeYmI3cKmDeLVeA8B1iQ18BKeaEmqt
pE4d21vq/lOJnaCNX4oMC7nDLztwKNLiquUcLbD3elYxMoiStW+KIO4cHasA5FKw
ru7zCXrVfXTIVaCv1HvGN3ojWti1f1y8s8/dvXDV+0O2fvkeKs0IejdcS7ajprVe
NyiuaTwxqMLJC0q6lnla6HMujxF1wQ296EHm3GAq3/Y4jYmOfePr1r1ma/VAEMVZ
+m+mKwWoGmbQ1btQoBoa9p6nWuapcII2ri0ILaI2cVsXiXTn9DrofR3VTYP/8dnL
69LU419qXHxqSy0nITP2YRSCSdhF+pirwCjqmkATnXUEMeAociI8HPlEdOdTgTkk
XfZYj1TThvzB9yxwyHNo+TwC8c61MKddNpn1btrYsXw8OGRb7KRMS7pY4gGg1MCZ
FH9by9Igd0nOikUlUshIHHVLVz/IegRQgMgMdeVaaDdQ2oMkqovbRJS2P9N8djI+
vK3MpqcRcAGhcISCSxYZKKEYQ+nmNMwrrbVERtduU41iTWZPFGrb2FhEvat2ghkM
ekYvr2FJh+EW+FD4WND1H1OqgyV/ETgfUpkIU/ho6OxtGQHflQNo3pUEkM8VXkRh
gFub8Pby63qITTSRVtntIhxkXlhiGEA4KZHJqMLjt4FQIgtQYe10lLGUPZjZ78SR
Yd57MIa8OHf21r4oqrKzBYXqXwS9tpjwFTmmjepiYzCl3lNv0j8yjmiG/lPqZlYz
RQIPg8R0zRRJwAjlJTJjLmsO8LqRf/jcM1ZQPwc5rfL2aMASUfyDSBIZBk6MEzOS
FWoAtdByvyCoOzrK2G27tyDs2Lh7q7DhZv+uDYeTKi7PjMaeFnTozWzLmL0JqwbD
kMI2YD2oO7lC9HSc0ejdXM9FdnXUzF6nMEzTYN90PDUvWlqpv4XMl97caXrcCPXW
S0VUr4nrmZ4CUxKyYWslBOvPDp84D7avpRrdsR6YPdO33O90Cuj/oYfj8eyoIp+z
6JHPzAB9ICfbg5y9Dii4+gUSYxB/TBKGq/tNWwgdJB6BAvg19sV/4JZk7jHlheRe
DcyXSVM9yqXZ03z/vX2UNsk7uibfjsi45CMGcMqi/kCuLNAglPEFoGyETPdfyews
13ltLeQFP94mXyIGj3ZqOGu3A3lodJi0LuWCMAYZSPfM+4FppzL/O0NBrdTmX4Qw
+oJe9hpG5gFBzQK/ykAfXgIADgv7IHzT/b+oHZ4D1Jv7G017R8yZ3gNvFxOH4pra
GJTP6GyyvtMeeVyUGQN9EZ881Y689a7OfwwhsdF4XBKKfijILsonyP/b0S1Dr98s
2Uk9qJ2HQoBi46kFKtvEvf8To8kbSavMxNzOXjdYT/fOiZ1uZplusbXxfW7222Eg
GVfovTaVzi4p1wSuv0A8i7UnKbZzAy+zjLcZcCME952fX6d1j30ZQPjeDVS2knAQ
ketIawDu+aKOLo3rW4GfQwh8DDpklNwNrWBbh/ZsqG7uhk9pMI/WJo+GutSA5eQR
NOc/tY5Gr0Iyz7S1W84jeW37RJFv/Hxfys/sLYh+wKrUAwv4VI3Bd1SQg2PA5QQM
pzgBtGywXgNA6oxZsJytMAz9cnP7sNmMvDb3WW/5X1gCeBrKkqdWsQqUTVZC+fGh
PSpiuZw4LkYxty/C2f12LFeoMWKzRs8mkbvuC6Xvm9545LMSyfAHAJpf9EvFrSEt
Ovsnuni9crt4/jvA2cGTvGXFWP/0FW3u7WYiKpifAx3AX600MVCFCtpJw/MnNkvK
w0B3bYphSna84hH/0C+zXulkMyqF6WVSoT8SF/p84kjBepCjfCmDi5lEDQRTGeEX
VQAa2fWR5sB9wb6aYzCX3zQQM6ed1D11CRv4jlL57adUMtsx25ga2tJ3ygCDmhAp
FNWlnTFC1GgX6m/tv0WVg20Dba2I8Qae7DFBS/Oq0MxadrZ2WXAScMaee+BkVB5D
eIUM0dOIdIHnB/pocUur4eu/wZ+hcsFTkGAjqJHa/e77n+UokkPIjQydANmDKpes
xdcrOfA4ThiKxa+DQ8gaZ+kmImx812rwvcfsda7NEWusCx9jc+poShs2uv53QP3U
Zod6H3YAna+mj1n3Br0h/DF7aE3QNGAN8E3oszcWV1qCaQ3tR+6yWwuMLOOJ9Let
hw9pX2uHvNRwmvJZQ2hgrsJNl1waHNdqf+K9ENzuhu2BD5b5wsKRXc1L8e8ybpMA
72po7SY5X6civMFQ2999tW/5VD93hT+br/YUdkUNuyPKa0YOTMzrAJ++uuYf3GON
JVySnQVqzeYNkWDd0Pu3x61fTrzI8ndHqhomW0wYCvj1xU1+90CWAAAx7tQRsz+J
T6+8FGW0CCL0I7uxAmCXtUfmelHIrGuGSRWjYB/QjNEf3H70xsn4blNXhXrOiV7H
H9REbrTM7uUa1WDbExXoEiA54GNeU9b8nHNWXVeJ7uHVlMkKA60QVczhI+BawAdl
dGho9q8xJp2WHq3SiEGHN62caZOkYGUDEtDUvK9u+oM6H7y7S4H3gKut2LsnXBYp
hNAz/XXPivOdsCcB/SuqAKNqIbsBHSRBhbgLE8RKDCyNeqRoTGZCKsdLJqg1nW65
C2Y345zJlgKVX3Fyv0AkA38y9CsYq1FQcISivfWsi5r45id3UkoogtEas7CrA5A3
hxM8c/ZqdT0Qfn8+rwcrQjD9NAkKB0V9M8wt8fJMoIQK5Ewrhkkxc9ENjUKhxPde
OmHTB9OvKsaZe2YJ3MsHUvSNC7HvhBNj+Maw8xCcBnCA+EHApTFgMEGrinG6Euea
sfrftj7wHLB7ZeIZEOvHxsqZU2pGtu9eACJ0lXPwG9ICr78Q7SXlvdY/6582n24D
UkMOHXzcZ3z9L9XbcEBeeG6ZW63aX0ZjyHBopsoTh60fbeSskFPgNoiYx6jHQInx
KI+TGAEbeLM9w4v7TBf45+n7zCpbOZnSUColgHCsW9SBF9eR6aX2ApkBRNOwYAb4
Keuhv+hbaVZkjqzaeXjzrvXAHtV2mUrJt6Q2P2pmULYjww8B4YeiJdtzL+ETxsMZ
3uKUhB5Ki/46cJYndZZJ0QRNyMB3VpRIzekiZ4DmbOs+8C80pZX2P2Y/SM0ggN6F
6NS657mt8vSbQ3eH2ts1zakG73jfzVsfpbW8EVSkPfMbY73gxsVVkZ3x/0cFNSTY
bWWro+hFExFF17HV+ULjytDIQGtrPBOuYlhKuwiDRbe7+L/Ydla0hPZD3tqgVRev
9ycEetwYdogjsr3KEkX4GwlZuUlD12IXVAMq2q055+T1kfSscyb2Ch9BFLJcsWKg
CrZrfnq+dLdaT9BlTSmHl8q32yJkExyw3+40e4MYRSy3j+ahBb8SP1z7iSBXc3JJ
avVQRdS629XZUffb0f6QAnDTXX6NysG9nF/GL/OXbEl02lw3Zuz4TyTg7Drpi1ua
IV7zGrF3jN/QrO8B+1cCEPcsRb3CESKwMCxHfpkO8fzzLPMWZXHzj+OTfokvd1tn
03mwA+f2jCbjZNGx6RTDGnjHHX35g6O8+ZyhLWnLg/YQGW25FICkYVefTt3ZKUrz
7PEYWXLAryJ+w8GqwY0TqUNOrnnb0nQmiG7g7+n1Kdxoa9StC5L1Wap+KvmjnvNF
LyeeEOyo8xYVWfMtHIYqPGL3O4gUAfITvJPxbN24CbGSqwcprCA6re+cbCS3wG9w
38QBNjWd+a7yMTJR0JgUVjfieERBzkNhmSBYZ3I3kYwfIkELQu7L5Er7imOyDwXv
S46/AvAK3r4QYhR/FRzyNSFv4p00doakzWEJEmLLoJdF4n11msEgVSZov/eWUbAs
91rVqjumrDcU0BA1U3YTdtQv69/uUuKZPxcEFOJJqx23AJR2ugAqv9ChgHkjLvvw
3m5NDDj0NiYYY3DzXmzFhLf0kpoIwe7UW9l7cTG190U62AAjZCeePKWul8q5HN9L
WST8Nm9ixE7vC+0t1TTP1QhqvNOmv5gf7sKMygYuFfKDyaaBAsS/yN6PbmQbevg0
yOy1rQBHGWsy47vWPLRc9+E/JExrrtKrcQGdFmceKmtuMm5HRwxefM4RyCUd3A1Y
fgiMnMWesnKa77vizap5MoniZQ/fnrFwaSQ7l2snGyvrakr9kt1K6ot5EMqSulLG
9E4ULsbZ5FEvpxXV6PB0tVwbi1SI6rJG3G/fz1l9iCkreNiplCo8iY/2/h3wc1ks
UdX4xHLhD1WxBxkTmV+sB5pNsjsTLm4Z1HJLwttl9P7RF0pdOQi4Eyffymcws5UZ
wG8p85dZbONxhfJeIcqtDEY4EgIlMKMvEDLFiXtCD+g8X9ywbCeVGUYLSJaYss/6
lIkLTiwg7d0xGnvQXOnowXC+EnPWREQynTGHQ+79EFKM4sRd16EbMna+65ZdY7Y1
yR5oDV9NP6TA65j+cXLpnIaMgUyMUxro6cBeocExtUIdq7bQNIHZgkFHsjxTsCy9
K5SX8jiX40+A8ZX2SyyE/igYoDmn8Kj7YUCYpiUtuq0oFURTD8+XPYqunmx0Xxki
rDT/CM9SaXknGGD6G/6kLupNjlC+QP82PF3VlV8bar47/Po1PbcXDo6FpjzQw2L5
sLIVPY0opaTkPF243JG4/TKxdxq+sraWflmGP6uUZEVmSuoDfNIjSlTxmdbjVE+s
ABy11OFbo7UNtKDtZjutFmO1Qnu8iOMAzdbluypQbjfDdSxMtvKyp2KkeNT+sEWl
ypdArnz1/UejoUPowLHBrZtLCV0kuIFdKgyuZLbNUnHnfLrgQGCh1wXP83ua2rEi
MIAiCHbyrPCc19FEHMx37mfH8nIOle6oE3nAM2j7bH9Zpnxpl7gQ/0TgVsP2Xi1d
vZR7/G7z4UlY6pakDAlfCLjGNQXllCit+oASkGT4+jPkymar7TfnUvSz8Hb1uMOp
09XhhSF4nwyWvs02m864WO2hxgspglLDKMTJWFQEenH+oPpWpJAd9TDwDcRUChde
p4YrVlB9FtQx0fDWZo7nV4RAyPKHpeUxZ+wO/3O8xlSPtoNekp4lax86c/Z2W61Y
wTUs9hK+s+PaNHIGqfL63XT4lboyDV7G5kqOtRhEkbEXGLUp+iIh2eWRyaJRw4Fo
wMvpFXxAqVOn5GiOkFbFJUNpM57MzLN05RHkIsWuxSNUztGwjvkiclIqDwpidHQj
G/0SRtspBeCi0Dw6BGDK+8Nhqo5JeJFQ/UouhB5Pw95U/crArj4tIeO5fMwVrwj9
icmoWvPHwioRamJh9k1k+iyp5ulEMj6SWvwe3D0EWqHQGmvxS76D0vTeZHn3tqpU
6U/rkKoOWIrym2HL1IZrviElKJvspmt2tHLczyeq9oxI6ONTMShiz4RCLPtErHyE
AQvuLXm44HNaYyi1PkZ5J/WVlghzgrDzkGKAubhQeHO7ylFnjCplGZJqix6goAqP
Q6EA27eJtbGZkqHPPb/9o2gSzdDCE4QLLtn87D1udzOJvDglar4OrJWNg1yek24+
bRWVitQHDN1u2LXihZLSrEKMUJAtEv4bmqstvWxVSso/ZuwIThKGymu/gQAlw3gr
KAFf0IynmUuTiVSBV71Kr6iZwXerTCRl5ZlZyOYLrZuDbAu6osASbwoVpt1g5nlm
ji2889AYRkE7lcDmGoA4UkLsOarQiXUFu4R12gbZWXseXm0BhGqXbPOgaei5DpWS
KP2l/4EsY/lMivzNU3lhZtcEf5EYwh8ch1l7PT4aqTSmU6O6axPkMHx47s3KUuV3
5B4LrMJxxsOKHVzrsrNR99DQzwtrmhCAw9xIiIlCkuJsLWV7bnPTf/b+M0gfkoPe
tmmV5aVdijGcRzRx0IyF5spsyVzHcxkERvAo+Cgl+mmo4Vl45ky1uTSxfRIclG1r
vdQ6F8xWZYnbRryhRLc6v82An2wiFrLUvuKqC5rcHAzSX2ZeXR7knDoiYAQAtuCT
EDS9RsCV0mMh8HQ4ONcdWt6NN8/OejoWSYimOAwEB14f0QHwxguHAhWil4jjdJJx
NXuxGAfBLtduB7VHZ7rQ8uaBdHFdpuRXHcmSHRv/1uBUQOwHWWYG71UqymdHwlnv
R8/pj5KwbPZIQEHptbTyUWe+zPCcS4aMLaDm9T/Xecd/tSL26cU8L4GLaH69JoHM
pvLFuYK9iO7jd0OT/mCyCtvMraOhf0GwHOZCQekFtON2Zy57ZVTTIIqUK7OSVIve
oswrW4uSxG7njSHGeHljyMwvmPGt5LY5bEijjHAGFNR3ZZbhtrQ41ahg03fsGtwY
8ygrjOPZlXNrMJ/9J6qFyvmBrnps23Y30eeeh6yUQ7avJLQDi1WkKru8/ilIairY
8EvJpC66CBElaxB/TuZ8DsSXYQKJhzG9lhPpzL+G8sEEQAvBFU1WsWpWZkPXXEZP
cwTOxJ55jpVNuBHxXXSDBpeD6OgjgdC9ygaFnXrMEpnZTyVsK/LRpOBWkBK2QbOp
LuSZuxXxRAoC8lcpkCmd5vOty/eW2VnHZwbZf+ORbjs8MmMR/U3siTl6wSLpBNuA
3vgQykYlO24W6I6hVPAi6RcFW2vMut5Ug64h4H2ncXHIBLQer3PSAKgxBxnJn0p8
53Jt/4YeyLE31TDFS7pZoYDiHzb8bziC+xQeuqfaIywHDLdI8ryMxNgFhzWhvFSc
Nlagoeo2P2Gd432tRFNPVpStsXxvlL3PjIGsPiLbWz6UkUtsIQoxXw75MBl5jVC3
ks1NWRV0t6NfKbvv4ZEpLhHioWDV4TqdK1Urw+DnDCW5KYmFdsxxfep9cbAxVorf
C06SNOnbEsFcj77qJJunFVHRIx6DcVvDV6/1onTvN9rYP/YT1K2yrzg3QE2xP8uX
Oz1ElqqFwE37z4uyQ5JORc1itigTC7KP3dU3y+jltOkE5c9O8kRbUT2foLKxG4zC
d24f0STev1oMKfzY6crVBYFur7DI2nqas+dMOrxrwCS9zJp4hLSZEj0iykXC4a8c
xF/QWs3rgqE+r+YGYAXlxjCGQOTx2TtKIQxxvShOVSBnzsl0LUVif3HBgbT/JMcT
H6VeXXtzAE8r89an0SnV9EQKabEimBOlLBnKEFb5N2v3ZjyQOa5eSNWTJ6PKhEaw
0WjQEve+eSavKpKfWQ2odMwioBle7k2Pbcz5SZXemk64otOQX+sRiMYkKreZ4VRl
CfJRU/Tu6dK3cRklfRL7f+ZBrp/SOzm+M6W4GZU+C1+RscGswrKN3BRkmU7EV6UL
cwST/IQcfPMJeX5fe5+YMa1QwERaSDL09dmUuz/OoXxx2WjB6HdTBA0A4JoaLgJI
vwd/G8B7OBnSm2wJMAgLvI5cnF+IrLW3Kc//lJYiVMkmOhF2vimKftx/fumo578F
+PGEwEOVgoFl+kJUJM2wbd5+JhAVEXMaxnlQXzTlPloyW85YuuQzhwNjDOkJau3F
Y+0TxxBAwuHaf1fgU+jGkxqW5EsWaoyoe+9htRTqrZ//jmiiJo/zb1qrY/DXH0fK
5UbpgnSyY7Dxs0x3Gn3AhdEqUADHSpv9REoyhE6ybjGhip7919ANdahuDSNXP8y6
DmSHOn8eaSzUsz97s0LxoqUS9i9mVag6wSCeNu7JO6/4qgTrgvZxObowRDJb767j
SFlch8zpPrR3eXTaG7+vveAGGGNlcxiAB1X+2vg7wzdA/DPKqLHAzGbaVNISh6PZ
CH8Ln2Gp80jJh6oXV+SMzzLs98YsXVpZhmfjRVBsQCA2+W37ZDQ5gPxt5cyKIsXj
juxWNlts3qETSZgGY8b1Xicwpal2TyFVpIH9jBLn7UxCFXwi57gF8Z9S4Ad2spGd
lYQtGnfrV3nhahbFDPNXnyLge/yW2eiw2jtAfgD47hI6JrXnOeWe3TX/9mZRsEuT
UjUzZ6/MHuLhDPgvLgDNrnjND72/4lq+CT26ly85y0mhXw//4MhVDjK8Et6b4npZ
7UFda8J+msKTq1H8E/bu5+TYd2+3ueIH6QpYuee3WrVVkFZ3EUjdr6U0Xt+0s+jk
9akDniVSZJoEd6vOXh5Xyo4QtMrZNbCmsYHuhN/h4+UzMhl5WhwSZG0vFUQpDbst
xoPmf+3tnRy3BgvKOWmIuu6FyqqCY/WEN+nA01OOALfqIUpnP3UYwu9naFLeCaQ2
oKvNMBOaOuZzPOQZhYHzp1nal8fXZlB2RtAXvQT4OxEVzEEwRPIy+SsFI7cUUhBC
jmDiPDod75pEc1ko3lOWcQB8C36dLOZ1wIg45zuqgRJRIWTaSoNpcEYW0VelDoBs
X0RydUCV9IoHEwNFo/Vjcvj4s7d3i82ymIsdl05LXT/6dpdvFNWcSFyP8tpJJSCy
BK1S5H1IvCKBUJShB2epzxkx0jFmxcEjst5B2v9CGVkRu7gt9QtXWsERfzQOSfsX
4tDQAdGyswklpscxLgVBxTx5Jwjx5Z4BRxuqWVsqLlu8o9RiuJ4KaT044qAC/9lb
f0bjUg9t6cYTbdzWPxAM6JIfbWLk4GI1f3MDT1gkEnyoaDBitwBWRGpv38eM5Wyj
GAf01uePBpiDQPu9OdLavxx98Fwfu0Hl+G7HfdkDQEAl2cMC+4Z4v671lwEhnr4s
V5U+aedzhfuFk1LJFSeRtxbmocOjn1UzNShNFk5lubCWkYxFGnoEDJUTAF2zuaLw
bntxAn6dJTN/Y/N5myl2aNar1BmP4eigZjy5btJXE3dOQkk8AvOpr36mQaavrRcz
vXUKAnr3L8I0CET121r20s9N8//natEfcPSIZXCkf+B5c+cUTiyuNTMfj8Zh/09U
MqI2TiIeO1c9kIXLpMjnc3RPA98FDL94Pk9NEmc56XWRUTgvBgKJ6mTAOVbzCk6W
QHIx3oJPMDZjdXU2qXCbtbBPGq2pZ8HbtOVqRorxW5DIVKm1oSaPNv01nodgFVho
6MM0Bdnq7I7yJgj3b4tYQ+CleZHMqS0jX5+dY6KoTaOys6odEa5zqRjCJkCNoIeS
+zVmhAFmNtv0kLKUrKCCIJbD24Lbyd1FvV6QEfJinBldHFq8RfCflBT06XReLUAj
Vl+xIToi5zGL/AF34/aLdl54WmTm9H5hm3rQsviSLtBlp4eSMzeEac7uf1CR4MaJ
cRj/kL28rbRW+Sf08t3xf0Moqd8DKIeLwd5jovk4PCPLIomq3KejqzsTQdqdctrg
nm8ihJd2Bfg3o4vInS6KkWvJFIJpGCSbKmLNm0FyQZXX6myDiKTyFCqZMI5pj9WN
gq2xIhn6Nsnp3RfiAbLeESbNBRNnI4W4jxrBOEnRt3OpASCpry9RzkM6CPXdt0O6
h+RNydmIj+uAH0a8VLgTNaME/xWpuoUrtPh4Ff4ZCbMorMSt764xYge8VqcD6mgX
CVc6rgj0rueR74J7N3fiFPi+fVHxomPSMZ/JegcPqc89peuZe4pf2avXWLcpCxEG
7C/zKAVfBP+DoG89gEgpsS5402iDQey8T9S9zLJSVSdiwaPpEa8KZzCYjmWOhZJl
IH2BzDi45jEnO5pY22w5f22SXZ1KZjHfcSVIlTQ0aaYs5WywOz8L/SKSVqeDuSeY
RJ1ReDMW0ke/Gb87ONLR+wj/4bdUZzXIzEQ3PpCvIIx5SzGfpU+AbfhI1TkdqoFP
HKYQqBRGyHkmtjWgE03yTBk7hjDUn703Qm4jJisBC3hEBYuJvuRZWos0dhBZMMmH
+CtopuFq7PHpY7+CFbSGjwxhGMrTakBTb6iubrfCstk9ko76mKTS5Y0CVbjtDe+d
3gPgv0nq7QOQtIMrhOVP60A3L1oe71JJefK3H1kxli3enFYputTeOgQNS59dkiyW
7imJ/XxvsMmgLEoa5RH97hjux9FFXP1kwadxZOO5G7fvDsbljXnCyKK6K8EUwbZZ
rkFnlicoabBWdcSKjfPV+QNQ3HBAXoavhsn0xRXPg9XHAmgM39PryocmqSYFnENj
2QsWdmvg0aCDUVVX6j48dOajRyHlZcT9RsEKQUyvEMG0ygTIbf9o8fe0S48JfZWm
V41fvg59ySbnzPKHB9hdfVnCLhFUilA0CME8Z2o3NJS9d74GCTR4GjtYnMbfY18r
e4vZGvqwExV1cC7GlYGpf/+AdL1GFJvABApUQ7i5E2GkWdBdpY5KCr+w95KVxo17
WjwKrTgIhE785z1/XwqR/h+kD7galTsNRx2IgaHMu1t/u0wzHtT9qpugW/SwuN4X
wrLCENHSb9eyqs63l2gykkrSJ/+k1r0PM1mCoX0XV+Sq8mkD9cdK+UWfAmJUv2XK
vtUoeoWMaUYCZRkJBWuNRM+vevl1/2LkVPw4aUQLDht9gFmP1W7tCZSkQ6SJlVPe
6l0b8FPpMUGdM3s1rS7P7SBqOImWWgCpXNXpsWNwwi5wAuvGJgqWKySdpsJHZxNz
wRWVYXocN9ZInoaH4sP7OrIg4ipzUoeq0h0FitfaFILrsJc0tnqc5eaj0Rc3F+Gi
WOnXu3rDGwZzZVZyTpvH+/HdP5+cBmNSh1sGgeIlLc1nWdosN6Kf9gNQB52dYo8y
oBHaFWBJdBa92ZlOy8qjhl9ukVv/UBvpGYty9lbhbZ1GoGiIooVurF45dC3A5Mcf
pqFIUEe5w7w+GFvQpEWrRGWmCJpjFFmgL1P7Xi9L/79NjDdl/Oxh8+wfJFOHLVdL
LLizhP9d+NQ+pWU+X7s7AYqgYOq0euoX5mk1xtT6yvqg2RN/yzAAXYbQKWkvlr3x
YKq9IdJiAUVGn0QknpVVP1sfrnXPck7dyeKR/CrvuGxzA7RPkMkn/XwHf3OIn8Bb
fAU7vmtLDojCk/95otypkpbZOCbhKmw36rg+MjS6Pi+WYaNm9ycRzsxziITpb9zp
byeP6QRqN0NJSH1uqj59PCLijuRQ6UQmHdp3fOA0ZqnmJi4hghDnufOBSLpZmoLM
pdBdSr9f/U8uvWCSfvlSDLA0FvcMaoMEBgWENpCAf8CsaHtvGkmuTewjR7b5snM2
fWRjO/EJklj6ytTE6g0qQ6H0N5GSMW9nt6ndtbTqaBhkW3Zx44e/ms/vgiibb8z1
chxZW/1UdcPe6Kh8qrKOSb5WH/CZWJMPF8q/VClg5zuA7ozBX4rudA71gphkrH+1
nce+ATt/5QdKRy3hdKTxzISH992VWzjPCzdXJ8dM4GDVx9fcnxti27x1KqvrpIgG
OuDi+nzngPS+bnxNkW+jqMdx1KXKhuDoRgkXSvQOR5sfa3nm1EVp1uz2Bq/gnEA1
PvseKBmHLaNEs5alyJrpyWxzjuSM3quoLYr6ipDgEGuLwzhWaNQcuJspON6PtRDZ
TNumzXgPZcjQC2FK0HONO5qqx4M7UoDcGzWSpVA83d/VGyh2q/ZE/HZb63IG5Ax1
y3XCoNyYdgIOl1cJoKr3piH31GnrgLYtvkg35sv/nmiMOjx08OcM8JZRRXeegEu5
34rYfy3APVImSED0xVoNOCwwrqYkX9dur3sjPXBqg3AjYXQYvEq/FRaDpcaFtb2l
zt2Ght+OMYgKlsfc9KEMtZxuoCqY51bFHIxqDNxErqOrUNzr3plQKMuzMLN7qvnU
tk7ny9CIOGiHESdtAiLcvbV0hqYlIfAmCVFvX0tgl+iZbN0MX9YYfeiiuClhXZzH
nmS2F3ccsVENhaYDcrwEE5b1UhoXZzfSQBZ5JmtVVncF1yxnO/RtrAN4tJnpByr5
RG9jzJaVZM3oqqVCPYYmtBDKCXyPqM1K2ztuMVHNueXh1e6kaE5hXR+Icu5/uOdc
ao4NK6eTQ1OG6QMIJnNA8iAKGh+l5XznmiqwASYb1zD6byY8nluJH/pOzlgt83yt
UaS2Ly7sAPxmpcAk/hkxDeypMfxGViTog3AwOpH/4XjGZHmTZhfqyfl+k15ZA7as
35EAnKKajXSsCqIuT6nq16V4W3kzqJwu18JIz5frZZbSx49qBWE+hFJKKpyWQd4u
XudWCGagsz3CwDUxVpVnfEqZxooDNmzgqeCTtBRi3rCyZyLWrCvAEPaCtbqTYZLU
3Af1FgAJcwR2gDC6QvUFGb21CbEVm4G6sNO1u47seAyiW13QXnz4+mPxiM/cR/Q5
bhCD4ynNBjdXIN2xZKQmUu74iVI/ZSamh97BkDo5LcLd6wizGqFIkVy9g5j1yyAQ
JJnI5bDTa357K7zgFIp4WO00H/+Y3AgjNqTKwU5r4NaUiT8M/CZKLpe9dtMo39wr
jQoSIFAbsW8BCWhi2MN5G0p5h+DnUu6Wua8jvSqXcwgaS8gsQei8hohsAlftguLK
uIv1OoPnWEA4b/4cOZtTDdH2JcO8A2TTiAbbQ672kUe/Ai3Nw50MmBWQbm91aSvg
SRjfildhALG9utMaKU5/iZgRMQcI4gRZlSlgZ/+BAzqLLpPMK6SA6pNbN1Cby5Ah
bsLWJ8NFZdxcF7ZVxd0oddX16OBK4HlmeSaNKvt9abU8tpviyQn43eaLAf+BN9B3
oj+vxK964k+gZJJmAfSRmce/oocoHaILpnUtd4BgwhaFbpVDoDCC5acx4JvHTVIN
LKBKOxlkb4PsIeA/1gmURb3bb3uuffeNYCgMa5Ip+1YB/s0vAVhT3rReo+5GHTpM
8vJPgphBSBdGKf9ByPPQayrjBj9qbTfkCxyJN5YcPI+h69qkHTPI+bsiCB+J2SED
VfZ9YL7PeJha2c7evG7JMmqI5AT8Zpt38UxAjy8JoAQC8ev+T5DKdaVfv/i0r9Rw
EYKvQw2vwzd0i8ku20uZ5k+Da4LrfegDwlbyAFjm+gcE3xCKqgMDqaTVpmBHL/rj
ckmmTCZFDTsGX/x+yOAIYBITwO/OGlsV4RwaLBxWKcQPq4D2iFqwNh7KiUXNMY8a
6XCxX66aW+33dm3Bj/GeIiAs068dOgqR1PZJ5NA72iys5FhXXOwzvRce0zaPPnPT
k9RRj/O6fCpF8AFa9hyvXnYb1BRF5eL/YcMoMj2s+E4GAqF2tDxvghdulL4zWi0Y
U7Ag7C/+e+piG/Smn2yTYbgjZ4NsMxGkA/8xf3+KOTn3TDUPQ0UdD4hbbBAzPupo
2YpzhK3f6izbkb/l0AybZSEdnOm0wOZEnIhFRwDLdGqkHf/qP5lRgiUPGYSucW7E
xrdrHhxE/uA6dSjpAXFrEwv4lQtjVXQqvlkwb3WiIDHNkSsKIqr2eXK7m4t6V+J9
zjZJQdfDewaz+FQD2/K/0eTiehgDFYPpnftx44GtOtE/k/ck1zb0Jq+P66truTE7
voYRoDE2wvqym0VluvJ2ohraKjatG0UfYVoPvjgQbaWOLOzQm7lZAh3kZZfITuvb
BTx0aYefHbmDk1LEI+92BpLA/LLS4PqVGMwQIJjmzm2g8ET4PtjwiQhaBFfVnV5N
v4tejbPkIQKZ2zY/Rbg5P+29jQoLy64YNUcy3yrqW0ZBF3ydMXeZ62gkRfl47nFS
m/OKVXg6iQE7RWgOEe4yOnLbKpC4BYuzVMKOGBz4xmN9CLwI04Wx9BxQW0YDJqso
9n/YHhEoe7IV9GrHhZN6Xe+g2ng0xMLJaUoT/be98biHBh90jTpQu2ux6zbEStvY
7kWcfJeXCLO/2kw/fP46ip9jAt9le0T2DpeGlLvJD6xGrEx4IPMgiQCYs1ecDkwk
0mOxrKxFw3ocqTrRMKaoUTw/2GQR2fFFT9TkoIToYYi7AYObXdLwF52jVZ7oN3xa
v7nymsRsEjgnDSKDpoYqZSDdWzZZId15n8QW6dBJSxxCdrvfe4MMjFMoj/KXnm4M
yn3UEeCb8F59y9wDlWtwOIY7k/XgkBzHjvNQZkh5JOe+OR5cELTpg/z5i18aIFa9
xK3LNVFYKWmv4eAeCuX84B452SoXtcYmATkIF2z3TyRW5hfNGayeUponmZQjWy+U
lIZLS/Ewkj8yzlSB2nNh8XdkKpGAfb4hJNZkoMaDlfarOoPrsEh7MOWR/ZvdjqGp
Z0Jf3kcLfOwMYfCHTqpurcMnSEbGB9iMQ3FMfJxOY4gnlLMq85VL37o76wB0vmAz
CEoRYdAWY4oMwHBwmibtpEcT0ydnzzIqei5gb8DQBJgzl3gMzeS8fs25sDy9NcXe
GZU+w1GTrmREkdnRsfQD6DBoXxMUV2NoBjbRrp8yYcXLtVIoZY3WEEsLIQ75R+fK
FC0mJ039PE/49Y1ulE/wW0UgkcFj4cQa0w/N2nRKsXQGeqrhDJjk9zgM1C1jWou3
JWSSpgb1TmjrzXoO/l3Iop6e1Q69B+qwywJ4SyrMJExHZwLhHf9ICC52Kouo3Ndu
SD2EryTNvfp/YKyXfZ+yvv5wg8TVsu82BzhUDDqgkGdDuR7GQGYMFrSWfJS7Rz7G
C5gQ1s/eUbGDW5XzdKQ3tbA4xA48oJm83E+adAe+DTp/7lXWz+wRkQUC4qclkMUV
6PTHiBOtaH1g/SnEiuWbEO0UrpspyivnXQSLRR7ABDaAUEy4S+yc1FsL3+f7wA4y
C1fROIDVdjcTporb7e4RNO65rt3LMv6ARcsh27tuEXv5yPtYLDdEZXETnQvOfAkV
68u82twhi18YvNjSn0d28fhGP0GGAjQsLBm1A/sBVjFgJQgDWV64I/JM6MRzkMUJ
veRILcH8z8NDAYF3EdXzVPExA714obdZkFUxvnMe7Ff21IkjWonzlH7W7h1b7YNZ
lp/SROVYkBFuAQBRsHu7oEp8diKyYfsN0ZW6usPW7Jx37Qc9pLayUzBZkwYn7Hua
Akyv3DbwUigARTaxtyZ4IJGpyip0j60BnqjCxQ3lO6WZ1CJkKHR/95gaQxr/v95r
HFNuXzgduU7z8N8/q3oWsOenyPR9Aj05auqS7+whmR3HdIA9AGWjO693ISApPl+M
ZIrJsp5uJJvzfEjAUbeWylNuVHITO0+6R8PZc1aWo2ogP64fP8YRe4qkb+fASGiy
L8u7atgI5SOIdCgC6ZsZLl8po9Y8ohtyEtFOiJtzaPs6ADSU7DNeXbhqnVoyo7jX
o2gbe3/+pWbV7PdKXmsqKL6tlCa1F6lbzuH0NW+QpU0mHd/3F1U1wzMwfFtuoLU+
ujF92PSS3vapuK1sZPCAU40riFhpQ7Zw2HCzLwQid5zAxARKenY7Gjw3U4wN/Dhe
DmSs/MBrT2CWEGG7VOtSu7LsZIqi57SpFUgRlLdTms7OdLOriJO6eDrXkfHBpNSf
5V+N7d48U7sPqWtMyQmn4c0Zu83oQ5n1zSBHoksW3j9hlFNqaY7sdUk0V9lUx5q/
o5j17guPMToTmrc0ltpBccfrmrLH7j5MBHW37gPQYBZ5bTkkYhYG+eCF5Z7VUZoi
o5yWTwWEN5ozgnVZrNAr8Bup6ZwGMcWLXehUo6k2pEpHOjP6+HHic9e034k2BLll
uSklJBdHTd+23R5/cOvVafm7cELqI1KwMfu7iHpbdQE4P2ZkoaVK/+qLJODSOSEs
SXLx6lBNdr8bOBUiMUB8jL+sCEB3RQTpGg9NPeBVE4Af7P2w+Dxz+QQAEYPGA5iK
lHEJlf1bjwPgrdPJEvH3eVaUKWFeda5KEmdUbUgfm7KRFe+iK4UXa9DAtVFtlwZc
CfD5tNlaanlfcTa/LBaAlk6Voo2ZdVi1r9msK0ZC0WY5deBsGC8aUDwe+3qLUaRa
Z5vjjjFz6FCFv2xANrhpGXChc4JSxgLSxPri+ciob4a0NNblM843j5OgDC4jwVpv
IZW4Fd/lDHy+j/+HkQNS2jNx05gC/i/Lggf2dco3Eqv3/XQ/5MXZh+AtMx0g12sY
hj4GPoIApmcnSGwZ+YcjP+e/GBKKmXBy8/Femr6hMg3rphH45y1FSDhCFJLGINdu
BexeU/gjSCWbKh4kHwaco3EorsoBbqDz+QPnHhAh9F/cPXidH3cyLOmF0ML3n9Aj
JV52C3f6E4A/kSr926GXwaATEiDkinGCvHwKfAOU0Mjr+ZEZW+LSZPBJRivpbkf+
c5qFBI9Kwwa8NNyN30dbLjO7xz78DAD+azL4lcdEejbxzaEpnI81Xqnxo96mk+6a
AY0ZUUdPp4ES2YvIuIJ/0tf5hF58b0DeAUot8RWSDlF04eDIzap+ebrU3A47DVkv
aTXNwfIfFE0rFat7rhLbv/oYdhNaeBWb/NNc+Oljj77jhG1z+VtkZgo7R2zcfHi5
jltHVARRVY8k1U+AUu5XTdpuZwSpapkHdSYZor3SSAhojlb2c6UKYW20Olw9Tp4V
bstiiOQ1RFEN+NeYtlaQdWsqzpsO3IEkUKrCgZihaObIy6XIDLQ7tx9ChI9h5XQS
HaLp4fsFrhB38LZL2U5isQcedRrCTxhVvd8Kmpv0q+o5jRbexeHSgJeeDjMPUqaC
4ST11bHJqhaAgt5KzPxJT2hyaCz68shPeJfjX2FUr0pJXbxnS8MVsiW+3ueUEumk
FMq+6OD3Wh8EWtZ4H2txWK1UGB9OR2b4P498KtVkgVeldLIH4vBv+TWyK45I264G
Wzte2hy0w/mvy8x5RbPjlQlrR5wCSvcM6F+8L4L44o1RR8HOjMyuxJFh0QCf9Uvq
CaSB6TeMVfU2nElK2Q6jaaNmESgoJwexURBehDylFJy5A2VHBCwAdkyNd2uV3jzw
j1glaINRcMqiXWUA4RKKFlem15u3rZur1rcoCzA1g8vXCsLXZkYSPWgdY0MMhieu
lFNLfMnVO4hTK8g8p7Njb4U8rPBE3sKbepYcJuYnY0kgRigPVZvIztYDKhOHmySx
4l5Gv+mcEGVLKUSlw84gNR008WUdkzOa+QEvy8wase9r08EHWKJ1JlV59OPqOk1A
asHWm3Fr5vs5w+qOGVuFVLtztpui9h0tjIoA6lNYAgC0diFw56cJyK8x/mEJ3oje
l/PVQa5GTQ1teGte/t2r3Ft1Zo+as3lBQ47yyt8eJnbccUQI4UEOjaiFeaAHIr66
4zxgpqDpkncJfPYOoAxeokHX5wkhXlLTzNDQN0hJhv4scE2CvgXMrIKsOmTedCd/
eJhmtYgBKeoV5ZMTWnujo33xzSjs/Dlnmy087L4qpe42ydYUmjdBEKA5IA1Jkg7S
3v/Iqrpx7UhQLp1rKDZfuhbNymkvVuK6blavXEbL9zbsiqokbmfHvyOpLv5TlGbV
F3+6mW3LS0HR5x71ZX/jqOczQXY3jMW/vfzvuCjEybqSatqQev4TeLv3JXEJvp1u
v8DFlRHsAkTbv5GE3o1W/23zSTEylzGMzYpfgAu5A9U23YHEs+n9w1d39daqVB/p
VpzB4TkxDBg4No8LckG5Nqup9Bgguizd8AwJP38Ounx57+11NXvmanpUVBUoLWIt
Ok7Qqq1ZCxMg916EVEFI/lQynZBCpg6LLj9ttxqbwxiW3J8H/1lP54BX33I37p7C
DbXXElDS9Ao+rUikjg+ULSWyLGbuqw1L77Y3ldmkydVRGr0nNUs11LcfSHLI83CY
IpYPhk1H2QX4WR5h+IuGf4j8AFIP3riaDXN/AWx7KXtaCHIAHt8B/+Ytza3PcQdS
t3Ds9KJW5jxWOzjbcnG04Z/h1yjILzLpuHvbzF2ioUfIs49W9dW+Ofi7s9X/7AWO
ielGZZIqJb4q8b++eHfWYD9AxY782zx089e3l80Bguzn+OAAQaQ1k+1m0zA5qEkN
Kaoc2aBLca45ocJdeuErN3IhtsJUnWrDYlizAbU7CJdt3iSNzXIGqxWO+ZGpSv/q
bElpa408r9FjCNvUsxr5ulS7ucFHLPm8g6AbwHWAsfTPpYKCefULHvYW58l5+Q8F
LjcklrL1xaSxMFAbUvKGqyl3UywtEW5eEg0mzRo0gpvk6McTFYO3jM4cDmZJD3k4
gZKNdwPjvao8HNJWfIuP7oRVHPYYfi+1dU0NGJO1iYy9db2pW2wqGFSPYYATN2C7
8yr6fuq0seCVUpoKp8LK+2yKMRIcw5RROyu5Pj0ZbJvYgFR4+6ev0yX9XZOOK0fy
DAv4fSnyHzHtS7HdYu6QTp/PgpiWuYJSk0olrR4Xoav204lbS6jw+Yv9sFjZErui
kRfk90JngDV85fqvUsxEnJywTmbWZa5J+pe7crUbPhg9fHXrFYEmmkD6i7/H4xkO
p0f0zJWBcknNMEDvdqT2GJ8PEKTcNHhFlQpXlDKFOftdzfmfhkXdd7pQA5BBn/fA
TkTjOzM4wC8oixxR+Bq4tbKEwu2mfkX+89YVmF9UTq+39MgkVU30yRTT95Q+txZb
+gt2COCgWIdEhCd2UyjSxD2QR6NwRD3KXzea05b6lY2qTefzVwmO0SEBVJpTEbyM
sqCGGr75eue8wHOr3dggS4X3dHi89mma4awE3JgwYYf13NY7BoLQfWJu3yoNuLHy
8VW9/jp4AN3jGYf8wPKAz0PJNY+rlvVV3epl92JqesaCpCQgGhrk3aL9YOOae5T0
K8YsMsZNB1n7qvREFtIwKaOQqcIvPEeQsWT348nuVKRh2235zdLv8iZ4BY7rVMSc
YElJo0XJN28cPBedFpYkDsvp+SzgjRpnhM3DdpyhdzPKSlKVI92vHUxcP8zQYS2m
jNhCWqEtBN9vvD5/44Hd5CQCtG1AXXlgfM6yzOhU6C7n7PpX2KhkqpDUgpBrOFMx
SGS2bi2zZ+t5Qx+AqdZe9jSQUKtv/WpqHS1rE3TnVjimGGTdiALKhCHh3YXRVWbP
EDubAAWwYIuHOjfWw03XuPH2wDLp74yuoEB7CyGqUwDZe23YRIZkrC3093KxZ5Ka
3+YPakOGJtE0DNN/cz6H+G5TyC/mxaC0E4lZer3yN74n84PazKXs9DabwFxa699R
k1gfMhsP9s/Beq+jf2UcZNot8JUMHY283Ob1tr092Sm8Q9jci2S0gCdvLKU37ivn
ZWUkzC6lgBCDfo366twNMltuhfP/w2+jZMEF2YDT6RVkfvvLJuaLQW207ijLeVC6
UZA8rcQ4E7YtrP1QS7jsERIJsCcFKf5vbBf76CoaMy7W0y0N1RAeXiupHh8ULbWg
W0lFKOP3rzi7bkZSy/rFeaAyTb3yu1hELf+Zm+R87HyEh7jc78Fiw0IjmjBjh11d
JiPbKYMChbI6Xq8uXcbUUfA2rj3jUkbXx4hiBd7za/U7Lgcj4Q/oej1FJ3cizMSv
sCrlF3btQzt5Xoy5a9c6wk6sOslaqRTCAL63NCncsyPbaJG21QPddGbHJyHpbG8B
YGoj9AtChH/ZtpdfvRKNZwtTXb4o29qbX4SidyK+KR4F8/jOow97oJuE+LoznRSx
WtmolprobV04IXYLVagjYsXANE2lDwFRtmInN0RbiaO+d9ucAZ1kSA+8wUzjSn5x
JhoAEo76ZZfj6UVAPpUb8jt5SEk1CDWGe2RTmT1rKI3ME1h9kgeCL7eKyNJR98/M
fke/Ybo14MhdQJ10gegiM5dd/+Ef88S13NhTxKLvjo5uN140AYfGdo/MprTXoAZu
4trqan94ZUM+F5StroppQTxBr9DDAzJvCXK4zmLOHioHKvydXG44dRWyMKW/+ZdF
CVVcd+684mcYiQqPYuCXqGm40xAh4oIxdkygtI2W6e1SfdWuapGhZ6e2q4ZkPBQN
47Iea2FO8MX82K5y4drXNq3Cy3eXIvKzWzFKIfo8gUq074Y/wQdeTD79aZaoV0Zp
QU8z+F/ky5+0zoAArtqIr0ZG1Suq0X+fNoYFl6LHGRPZBnyaCzqe5BScU+6Calor
DVltJ9ZXXH1ae69P4+FGT0Ygf7tnMbpbbc/EDQK/VVS6vgVXHXe8xFHVwXhGIECU
3GZyViLXFKfRjimSY7ln4hqu9/j3TEJmE1WE8lNq4af3/J/dfHYcQs467PqZRys1
YQL9lUx1Hmdh+XfLkFr9Ma/BSxfiO+QohR9Z8OFppETKfIuDGzDT9Y2m4ECDmLkC
gh6Y2ybBS811ZATDgBBCdkIcWFVhaC7eWTVu5so1Bgdu5ONA6yaHHVrsBEoyADTs
E2gN83aTqoUFu2ZEO4Q/H5pFe/EwhFGOITlR4oba9Nh0bTUmJB0PS+gPJ636m5RJ
nc6/2+EalFztJ4LAYKsxVTB1CjRwPmM8A9Ua5mo+ZzCujGsKKmfZef9ImpZDFE3d
I0F/RaF5lBrxcj97J1QKkArxR5JTSdxbt9UiO1t9YnCKGvgmSyF8qIelH1AHVg5M
BIQ8rxH9Fi9LjT3J8ske7gR1syLaBVbyR+MpM/mGThJEn6xxb4oS8/sFbK47b2c7
hdZBJA5sj+QNzCYZFjV7uFVoy3HtUb+NCHEeYZ1QDVX7I9O+/sX51xZLpDnz1wwv
EQvMBWiB3J3dNBVecUsL4qUlEsWeGxV2SRzpwtCDEI0zRSvKAZj0FI8qonkitnBP
eXR5uXbJMJtnLqLgPVM5xZ5j+tG8tolppaj4UZHpojvmBe7kEBjbGZ6hjEHacZse
XigJm6YDxrQlHYxGiv5FgMnyHwessPNPmPYhb4R7HmwQT9HHFSwg75iZMxI8OLNr
fjmSBseIjP1Apco+7EeyI+5N6BsEdVDe2Wqc5I00yWi+yDmyKRvBajceDAkQ3jGM
LwGxniSX5K8xCTtxK5jVZ4ABY01fuWBvxb2j+trWyyUMgC0lDxzY1SxVuQgSKRDa
UbAxfqG/WVnNBUkRQaTflUGNTIDyf5PY02tsn3Q+cmWdbIV8yPxiZkgxUygQUnc1
sM7PsArZYY6xP2awXlhRPCBy97/+3Dt1i9TS6+SZqRRNKzRPsx6W5WD5gpErI7Ap
KSdflqYmWT3nWcH4JL3atGdrHRBSrZqtT7gCqQ21lHWQF2d/kQAl4Uv7RngFEhU9
H9pd4rmxgPRbHjOSksNdkYfK+H14Aaev97AjDIPgBRdd79bmuk1tigay++r5UKaP
/hcx/OzRFC9+dYJtd8z2t56/N72D/bTMEjPXptGV/LpbLpGZYfna3/w41ZmNrhe6
San9p5g6lvqC4+DC74GxUcjiHAYVlfmrroPxOctvJ/Et9gCpRfWQA9kVj0vqd6E+
5qG4fz/lcPFQp4YuLEvpx811ZJdnIhlZqBtWEEpfm1hGIbEy5mS0YnljgwTe5dOr
nCzUhoUA7mYW4MhpsHry0pOCI4RB+rqBZde7kYqgpZIc1gsAi2YXh8wEi/nzcq5r
4NhJ8Cu1dKf1FPGRnrHkl5BMCMmSQYcWDlr3hwuj6Mu9OIN6fjepBR3O+HmfrT0G
xYM10mkRTYjSgCGUzNdrJnhQALNkcZE9KB2juJNt6T+X2SfeHcUblgwnEwBUK7Oo
nWroHqOY85aMhnWGlbaWqbxURmX4AOOmOjPWon84nkD9gBde5wsTIAOeYU+hPSnB
hJ21veGVlMX0pLttGb65kJIHDI15UHipFPP4ALmGa0D4NFHxWTaILhrLkgoDa65s
RedrzszN8IvchCftXIkbp41rKFiKXae1BS+werzT9j/yYpEAJdJr9Zve0nfj5muI
0fW/GaixOliG1f+qGAdJJPWR95QqZWNtVdstGZsIIJPGaW1mBUN4nluR7YNVqIw/
hq1wB3Pbt9LVucXz8wF26p+67KZvalCfWNxpD600SNlCZj3zYXS0qipMuU/oV67y
szhQ7WFHNFuOiEFgDK6FbCBms13hldIg9f3jTRWbm5aj20alUhZ3R/aaeRqauOoR
Nrj3xTwHRFSghCO20kPAKiWkGE5OiNyTjtz+lvHzVysjXj4ytXfPBcxALRzFWsUM
XhEbfzmtIUgb1/QVHiMThrttMnTL03fIMFA685HE+Pqw5YlQmaGvQTz5gzmUMW0c
oaHThQ5v9uGXT/nh48gUzkQxoQqbxDHmhAZ7sFoUbJKoIIUWEHGIG3nUhAVApflf
7JQGgRS2+8HA/DYvroJHPHqRUlQnE3XVmawEi8OsIeLjxlY9bkdO5h4BRYe+xCok
CW5KknONpyglieXrvuUzcaIVJe9cu5VeISobYrX26CeX7xlaytrHWSMadzsuwpdz
TJJdgV3N+54m4SGaGHv0JMEuaAhEgI3KzVCs9AQAggIm5NbXY9k1v+ayRFxLUioF
c+NfLSY5A90XNhf3wFwWD2z+TR/xiD7l2kLAPobjGn5RVv4FvuPy1H4bJWdEbyQC
E6sKyaWs7r2LsKvTROGgHcTtvY4Jjt1OEF2zGQzzYIBRYvWbNFsPmIL8YWpBT62c
5sBr6iKsEhQ01OeckCluRRrqxIkpzpazyDRGMN2QtBUuo33jKCIi+30NCULFQP2e
pZex2seiA/AdG43gnGBrfx+LzRdf3t7WvmTTFaIRTuGpHGdtWcNCVKVTmlXsO/qA
obdmMBt+Sv3B7qmCR8mbkX1UveETgJNQPyEdVqitYAY1JmFou0QT2KgpbsrF3F1b
Z7zrwdlRIiJCNvEXwbSoFcJW9996E1BuSJ5b6rftH+l1nsLiJYke/3fkqyd0woLs
yDMGuPqWubbWIAyH/GkiR7l8OUV3MC45ArNOGg2FeJbs5q0lEEcDZWSXE3gGhd6g
Wgga+jepN/tz3RHXogSM/xz27R3yALvVrNjb2B0WT35k/T87tBd12LBnrVDiwCCM
/5wqQi2wedcJ44oEOYINwpStvj/g9m1JDkLQEb5KMIXVVn2AzSNBX3B3CaIkkZgu
Bc+xdj3dLk80ZRu2e08qYRrOVBxPsWjmDXpgjRslYFxKC0TzjhGQU49E3RquOn9j
t22B73s/oIuzMkR7VzQ9y/kcKZl5BrwW194bLbz4/U1AVVwFQX42euG3irvpLIXb
NtUPlwDIMwbHsedDDd/u/Camu566Ich0zIucnXI25SSXlus/QXFAx4w3lOI48g2I
mb42GXkz9XShfO8m3FUfHrOiQvgrEyFQvH0DY4z4EbOJWbxfeINYLFaQQ1IXafAw
8yoW4WnoBadex0oFfFdNvVjdNsjdRTH8yhtQY9+1/MsRL+gEbDLHTLL9XpFaSWBK
id3cIYpYcotWIH6nKVeJ9CMeixRcyk5hvl4xE97dZd7IIi94wuBZQAhgfzQVrHqy
K4MZnN3Bya+DLGGYTllppO7b2cI5l+5fIcCmYSbyPPM2I4LygB6UD/ZtEvCC2dZJ
E8oolP2Jy2e27SYQ0hKNRCjGIEb3f+0rjiHlMUBPBqcwcqbOX28HAOSaAypvWM4r
lD7MwVCVOXx+G2ucsqKWtKtTZ8kpvGV0UBmq70990qScPi8+CxYm0byqqIPMlerZ
hfk5d253wdI1kDdpQ6eERUj/XBoLAokwxtZl3caRVQ0ToXjSZv/bSMhRRaHbk8Hh
DKtvYF7jlKTHQYuMizkBamZ4fAgU7rSl+5QDMQMAefT+0nsTLqlRSstpwbcNs9MX
DKNx7ybDkG28iit9OabbCU+40vw6182+zP3UO9lHvKcovTwhl2H78bDL6hwjtMRT
wSbYIiZC2q9Efm1TD2z6JU10POuPqgOKw7+7QlAKU+r7JrakGi1wt11aNiocXSBA
+JkGiEoEpyuKDhQY31JtG7fOvmB1FJbpdK11r62vGmeif0Z6pY4M7hOIbffmF7Y3
lgEjanXdStQp2xzwMEgBHLjmT9VO5SN1bANSHBwh4b5Yx0X2bcYCN0kFa8c3XG8M
2qLw0k4MMelb/QSgCbR+ACYlSfDmqZloGQofGhDJQMhgPsUa8+iuKGq71ZoU6QLi
lwFGOsZ7Oa+C9uSv2BBnfB9MOBb2NdGjxg0UhWpSFDtBo5xUipY3l3NLI9OZoLXP
dGCQwxChYlIiFwhnM0p5CwILu6Xrm4cA6jU4vaKdfF4E5jUD4xke8AwT5TJxMOVt
IqmgHLZmEbd4fiCSy86TOeRzCmJIwqcwtnTm1ZFCHQ4NPVGnmXY+LC1VF1xaq8Kj
92XoEciiR3D4f3m2DcIKU8R1uLTJo6Y9mmYAOjck+M/W/fg2ZuNP94CWHxNzXimd
d/Rw6Z3R/Zk859NIeWGCFfGTahFND01zjPN4CEpg+mKWsyPmaTIm4rMyuURRJTIL
ZjrwjD9pC9FLDXpdVi0ZMnLgmZBMGNCRNS7XDL0q5IvmmTSdDOwz6qSLun3EysjN
iInOr4aHLzt34635Ic8lJOxeXpiFi7KyxAXFEIyeWIEP+47rkSwSAO/hdtiCQdmh
ro3Z0EzUpZtoK7Y/8z5cK/at1rLpp+wAjs+eWMVz3goL0Eah81adKlog6vSFJlxp
iILn36XNVvU7IOjA424Qha5GeYx2tfyAyMgaumP1yiuOyaVKgoVf8sYDFpylzK3L
NcE39guEpY2ygkUs8e+8GsQbc92mJ9JA6KbsTgV17WR0EHJo0Iaci0aQkCwmxSYB
q6croxSwUmLI+hhdcFeLbCT+5yJ3rl47vx/su3t2sDnxYjdTwzog9Nne65EHB9al
VSU8birq4VOiuOyhxLr7EFOO0QJzAfPc+4S8tPkHACc+DEH+cJkpKBM4ANKXQaQp
zOrLcWbteJ0txrQvQzou0vRxpKF/OHwtYkXWpdygpM1PvasKrr1+eke5UTprv9KN
mPzB9EXPx5nnr0q2ayuwl5XBXIabLIc6vVnvcdkwns7mccTdy3fkpJ60kAHhM1+6
PnJuxohAtsyAedbUJ0LuFRMlbt8TSxU06QTzwvuP5X0IOexHPlZpLPbCZmCD2z0t
+OcdxIXVFvV1jT42qyk2b0vsmZoc32Jtd/rawsrtgplHqatulytMLrfcDuOuF2Ex
69wS0qJOzUVxLmJsDTBOZam+Kacyc+/5vhclsi0QDKxqRuR1Zrs8IqxdsS6Xi5UP
x+LZvTcNTdqPc8IL12JXTfG2HXZW1ul4HCYeBUw79gGk+/kWL/ri4TMLDKoNPZnw
TUpx78EYQbf2IaieKqHANIF5hKotED99ps3mbI2orpM6uh3y1l6BjoEfBOY5y0Q/
aUQKydG9UBS10CWU+QPKJ8EsQ8WwTOT4Yu16dscuO8GTCbGCJDypJXdKi0r9Eodg
FchS3l6KkaEDrU49W/Jl7wsxIyzjXdLCcfwPewBw9lfH/GCCfFj23RsEc5DHIhSu
XWjB9klrQhUCX4eMMlXsKrbxTcohLaBAQfGpL4q0WDh115hjnEjrBfJBS8C+gCtx
Gz/LCjbJeuoZ67o/ZjnU5BoYoeyuGUKI3zAIrsEvYEjlGW7oFMlyPwDSoS945JeZ
8N/VhvbxBiwobGD1WZLASQIlBXh0wI20a1ezkhg+zrBitJNpXlydmwSD3mjiTKFY
cc37j43hd8WYrNMmcuTh0ZwwFEjKXS8RGvX4iTRXwtwu93KgbhThk+xhNH+OUofo
FVSQIbHzuPnc0M9UAt62ulNNjUI3iZcW4sM/uKwxNYmIBPoZinvg6oLPpjCFBYGP
Z0DhWIctzImshTQaPs2Eqe443y5yUKCEnhPezIjNAPA2QfHGzti9CvjVUCyPCuhU
sKRcYh09so85/lIQ8hsqcvwS3OFdZd3e/1RHFjRfaoMjIcYn5NuUtMNjs1p+0IGo
bIoqZUEEiXKIGE7wGQxxYifvb5lU/8SzoEFeBfnk6krWzxsq+3Bq0/NXJGE/Jjc0
01hJxMwUrXUsEbCmadrtAlCBKvap4Sfs61rM/V5xoGdYplOAg8F4ROY2Rk14KzIx
SfXpn8nPzRgIsjNDAXn9mXAehssLj20V95/snEKJ7M4bhZuFYiv9ldLrrVhWdrAN
QP7q1ug/hMmXtjFhoPGxBJyTvzuGxfyp2slPr/QeGKWqRWJyvybJ0yHSShfPkiFV
rNxKQXMz1AZ6bdQbWPyzBbY1NnFAwgCf+EZK6HW9hK1spwoROeZwqPqH+1pQ2aP1
9XE+G9b2Xt7FdEDyOWm5Ws1nIKoGrUtBGQDLF75gsoPz5IrRDyPVbKhaZLXGIlp5
ueR5Oupumf7kRIvaQdOjneZoj5aeEvgxDnuXFXfTPr5tGReeYCur7Wm2a030rz5i
Oawi+qWjbfFV34xjbQEHf0Pjkr9u3wBaJMDcSra3z5cPxtui4q52pmRbluhO+8HH
HNT0CvsUv2FLbGB7Md1/rSMPEXU0y2yUpguaTLXWsNJmxx6sr6debMJjL7cO6LnP
xAi8c6ySo9WH+e6hTT1ieRRbz5CtA7zas+JGsf61swMvBQWzj9qzNeF3dBbcCWZ7
hA57yaw891tR3XM4A/OVXS+hq3l+jrEXQxbYpWikgXpvPpyLza9h+86ud89N96Jn
iCg8Pgb2rkFHuU3Sy+R9XS3Glbiie7j84MQDwoUqIfvPyQTw4SpVTJlMehKc8wkw
VYQ5IGK5wakmNLJMFrpJq/5G5jQMmrh/P9TrzKj06HL9t0M+mVef/KUjwiNcSHGU
mdkQk9A8a2AvXJHH0nRR/tTEq6XV91oRGOSYyxNulYEZrc4MUPGqlr43nlrRGag9
EEV12VQdDWAuKIFE/cFAwNNh6P0qmyxjA/sG8E5iiQWIz9qOi1C9DNf+/oGLKUjf
2Ir7kT6OkogfXcFWmEFd0Y14YqPykKXD1GXkLA4MBwsP+ZutwDIgwIV8PPPsqhYB
K5LCHUxZwfoFsn9l2i8IsXZdG3/pzlPHnrCILZ/lZWzoGGNTvOg0vKsU+kIT5v9r
RsmrxdQVKwNqHWsDif7Y0ZME11f3ZZvun2AkkXChuNDghtVNWIHORQHvN5mfdQXi
GSbHtvigF+UKzqRxrLtybR2WLKrBZtHQDSUR1Z+Lo5JOuEvTjxDmOB0mO9b9f9im
uRiDmFIm9Xu1BS4x9P4vSx5QBnldumx9lf3w+Ya4tCBRkpNjIEflDaqePUfuYJnR
DzA2vzGPPkgk5v+mS2UU4HcbE4UCej74hhzGGQO/hD/uaHd64NCe8h9O2mGC7xpS
EMlGNy/naElbc67ufIcGiApmxdOeSivNjwdb7mOrg0DZoApvtK4b0lSy9YTZqdWc
Owb/juIq8KdooUJW69WM6qcl3tGgb7lf9extYVT6nCVrwWLXv7VZJxxDV6Deg9aL
6QLEO1+byTp6/CkZW1gDwI8adbOV4j94tumc/vESNZ9d92CIJOFCWpRT44js105Y
Jkd2MazmILV99ajfiOkxs4zXYLbHSknlS+32zJvp0VMkxPYvvveZNDF8KYQ3Amlk
YnYgMCYfalKNfqFN4C17TOlRyGpmpj+TADG75eoCWzJ+zljuK9oquwfcUlU3Xa8C
5RfYsH8UY3JgI/8GKqDOYOPJdDhSkJgUofJTvzWVlN8eP3QaYVTB395eN3P+QlKv
HJBAed4zJQRiXhFr4aZrCeDHFZbKW3FbcH66icMCTwrGVdfIAwjFeSQunR4nKLsI
OI57yLJlOf+ECg+sLF4r4NBCHoDKzOU+vF9+jDdGzRngfz3WZgGH4ZcxAvomTjvq
J2vUd++7DjA09GaHf9NshvUcj9qfkwXLHb4stXKIxASBDcCom8DErBY9t59hkCFh
i7v+zhPiOEAMs3JZt8WO952oxLuhehhc2RDMUPSuqTOGA+YRveX8Z5+b4LFMjBmW
LVKgBp/Z0aX8yAiw7olClQokjxWbET4NuJImx1Pvop9FfgiAFUlxGdGJEDqIyrHZ
/1yo5iK+dMssg0vA0IO5GrVdhORVsgAcFZ5f4P2jLF5Jpl/MPLE9sOfe2bd7hIuI
1zwPLeHuJQG8Qu9TEb1UCizP/nrt4EkI/RpCrkxmxHJSL7OJ7T59bBbYkFm9fpIS
wmNY0Ga7kVcFjYjHdOtwkdfUtCowjgGc3x84Ciig5YNmRx25PQzDGB+14oyz5A2O
smk1s2EX5FWua771Zvtx6m+tbVy6b3jnHgGSn1IcML6qK9VJ4jxq0t2euezNK+ge
Z3d60djtnRdQ31FxTpaXwtjhbv7uUxyuc0ACrbdBg2jCEXzxBODxnABRaJy6hzFW
eDpW3bTKghWzMnC4Tfld5qvB1zG0A1YKlpCy2pZU9A66OCx2T6b9SR2Wlzz+DO8F
2f2VxhP8yGTq1sK5taGroydfIX6YLpmhjtKZEM/mH9EgjVHRSDYeiHLbm0burikj
v+IBiBWVaxVRQyctTKHYbKiH2zBcJ6d0tt7+S+JDj7ghcfo0NXw2KKcJB9J1Z8vw
UyV15C22y1uoOzdgXrSkteUEGF9hup+0YejH3gaCOPAHWHhYVjjjkW4zuvBRdg+k
FZ9sbCSNMrkbvrAClgRz3omyteNM9lR5s8Sc1kpbBsNl0wdOJHhE8oYxcSVkdsDY
N0lFPhySErtXaqVGpYQwYtLRLNrPyzE6luyeTnryqaoGc4fx0Z0FEYmHFJxSuYly
A0qXGQvUuc74iuED5JYPQDsoQDRxEBBm11Pwa/oXmxPxmBNVlNFmzuQbpXvHv1uZ
cM29qGRQj9Mf2BlfwaPg+y45Az5GpXRVn0CF0g4MEeFHyw7RR0D+m4hZt9kE1+5n
iWhGZCRTz39oIDh8GtGZxveHjTn553ejxebwNi51c9azm5U4CDKiOV/O7tQGYOPE
UGu23pPF4wH4nIHj7CoKjujfEBK3TvbhiFMT075DpZHYRA+g9eaIjJMKkuj2qAkH
VZvktaWBjbayT7s26iFqKOzMMTzLWeDPNuYK0ZLDMNDw4r3Ks+FSDwB1wcSxHzUU
vQLS2HwbC5N45N2E39JzO29NdiAuVqA95Wym+WNgdukZ8NpY7ZB7xpihanbqSOAs
VGigibCfKj9SythxmxtNXHf3J7Gq+1xKyu7qiBVlPNntF2uqD21JeSCHeaq7QaTX
jJjdn3pJy/0ePKJN5sp8jS3f2Q0eJvmGLWaNRf0ZXGOZRdzp4bFwHirG2LgnuJNy
GeBXUjz9muOm7mAZCBvcCADQKLHjNzqDx7PhX77kdxfmKisNizAcWb25NtiHdo2T
Ii4GE3psWA8rTFrcjhA9lhXbEIJujkFruRPA+liGmWQUKc60fHNAGm/luTdv2vSl
9tfP/g3794GGc329IdD67c68c4aR6jPxhlgt271GR2iYRVzMaWy+b0/sGyfSUvVn
T5/4dr9/mnJEQvMmebc2QfQPDZU+AnypPFnzBCRWRMyK1QpXRcHumKWuC3AuUtWu
13weaZybt5CvfoPIS5y9ut/bLrke4c7MWGzbGIdxB/VlFyQvDDfiq2sxcSBGJrne
KEpBRTeAzhNHcfcE7w72ESzJSBpse4B902yWWIv9A81+YHmcUhnV3H7ypI3X/Uqn
PfS5V957gbbjVd7GIaFNBYm3MjOCbSX9TEkC3x8PQtLTlaKJb6D40MAcwRU8IyFd
Lj1DtnF80spx0cta5y6TiW1cBLKzIHl6l3I9tPw5E8roGCoBHm68alCUO6ORVntl
L4wgTtULXsjEjv/PrrDzz1R871ywfg5FQtVscLpAvGDy6mD8ac1+uE8dYQu/aVmk
3EOUiVGoYwGrqBaDj1+s/khAW16yFrt5kShafwdS45oVHl0pMW3sG4nLdUbj6MR7
ph/pabnVJOKGZIObPR5SR3X8AsL+fMhP2EA9dV6cgLynH7P3qhQNPOdNnRrTgr/N
9zg87EKmPwqpbIz7LeQYpkAS0ky3bVYiS0C6Lp3vAoOjXR6siJgjx+OP+b3bA2K6
t2SDWRbio7Qi9a6DJ9xaxCyFqr5vaVDgFV/Sgyuc3MVgCZVnar4V3iifpxZnyeGV
8ARyCfFgkLu+Ukt31I1CqfneMeddFPMPF6IOdTXTouRFBvNDybYZplE2duAJV1J2
wp8i2X65KkkEzlX+u6GRga9Ywx4RWZYUIC88VVe5lL9tBzx8uhidbh+e9Okg5lQB
Elu/q3lgpT1HGJOgoqwUu+Natf9N66ESfG4+r2doMr0oFKBJYBizV0H7Gh+WQ3g2
dCGNIDxpFkpRXrM5arOU9UMElFar/a1Y3mz1l9hRWQ/XkwW8c/zHMwu9jMXL86Ao
46zgNuCpG8TUyg6Ac6NptTPBMfdyqF8M8VKHcK6tFI8hAlh/vCE3P2DBMte7KGra
/xBeNtvMwoPzvzYGg240TEIVWIxIoEviVPO2siRT6GAQsge21ie8Ucw+0PESMUyF
t5pck/cvlUjtWeG0uw/0M9u+c1f6w7m5L7ByKgD0XOj3tyH9cAQsjQPXwm68tN3E
oLGeRiBGlMH0X3/YTBPqdBkEOBVQ2JS2x7IswDN5Uv478/MM2yUgqN99a5vaCgyK
wC7lKT4hSDf1NBKhsQtMDvT84ny02ftExNfllv1G52IgFaXa+XFxgSuzlQDA+FBQ
Y1W47yszOTjxLmaqMFKOqg6zHdHGiENLPVPGu5oIAitLvFLlw2Nxsis+Zbr8tIle
qeMsloODHtCNP3D9YpQv98Ey6GdDGCdkTylzKIRrbpmXET5jiYB/WTQl9FqA1fCV
m5AJ+K6avEZ68FatIK9rg7IQ21bcDtDzDDL+trlKd61RTfZsPGc1DXKo5bmdOq48
rsE9WgcWE0oJ5HTPu3FjRqDWTJPgWU7VuIoz8nQtOEOtND5of29+ZigliOmvLpdt
KgeTVQkFFflXzsMlZP/MgGuZ9fvoGMxOjgHWamiIkFvhZu62F9w0tk82p8qsEgUk
QtCsv/2Cms86DxjMKm3itCf7NqcXE4vN0gD40wNPcFXFp4Ei0LbAMZHxCc9Nk0eE
xKEOuXW8wGfFkJs23ceBaTGN5ZQh6mNouFUAf4T69Ey757OdAKx45qy7DU5zuaHh
y1btTHYl1JP2lxGdqLDFgE3+Ymo1chdPFmFDLYqAcsW/NohnMKtwst7rGUSQI1fF
uIJblsFrxz/B21FxJ+pXGqPiqde64uhKgnTJP8S/XZgwo3MQyq2P47PhkLdY8Obn
Pu1OpUpoX1Jyq+StXifArL1DMB9ldgtc5KftFxPo8JJOZsG5SrzgMzkALc9CMtpw
jk+XjSvIqxoOOwxaPXgo9aG14f/lP/eMCO+5y3ie4K0k3IgohtmiZGGKtJXT9QBF
ee07XcQTP2/n42ybqtfeKupZrhA3mnpxAAqCB/MNZeJ0kt7CkKsx+V9Pt5q+MdQK
i7DLMN3XwWM1Nn+tJlGna8K+/TqLzwciaNdBmnsXjAiMSVuMqto43BknzEAN5dWi
8Tuh7tsLxE1ynxvaudwM6ATK4I+3EoRnvem8Da60JniZt+aVRsb2faSK3SxROUtF
Va4AGsYblzlyBnVgo5R6Qm685BqhXrqBuD+t8Y3W73nttIzj4ekNXGNNmy06ejrQ
AC+9j9gmKLfAvZcuc1VtvRMLYF2XQ6YK5RFSl14sfU99L3AI9/aAU/1ShJrJvfK+
0GTNy/FGbyalKKiCGA7EATHFJ5on7RltGDDl9E1pUAmJXC14NYRzpumaLDxoAeUC
Qmdtdq0+b/5+4FeUhSlu8JFih3J6V78OBw/dgASKXe1v4jbHOLolovjVcUuQJ1Ko
DnLnqdp9lW3+iDVkDtwS26qfJWOj5z+6K5X9wVaqrYw3gIvL2yzQR5vUzGM3e8f/
hxrVfHEHvF2ytX2CULE0BygrSOUWb+W5p/ISAKUgnqUXqDCviI5eJCwzGvhhtUh4
8wTbdxFt6GqkOMyVp8kXKLpWZrbNiH0zKswHy4Nhynf5zrsUiodyUGgoJ9M2vMK9
L3Qt2S6hmKVTOAYTpKmX97ovlOPiNiU201p4pWV+5l3EaTAr6gCuP7m0/E0zd4wK
5/5hJEzxeRVF8nyR7G+lHdUOC2vfj73XVF22+HygqNuly19QkcOUMHGJigJQcHgY
K8tplnOsTFTrBEKUb56EVxT6Zvy49BZthmAFapv45BAMhP7d/7I/v88uUYjuPuDl
n4URFxqis9stpl4JR7z7rAMWc1+nKnuzyHIF4Y5+onGfpzAnoqJbYD69bGJ+brqq
vmciwM5VyPzfWHjXxHINNoZHk/37rNlhjzW8lh2nN/jH+3vV9FxQwj3NyPN4xAaE
Rw4eaxFQ+IleAwA3icBfp/baXj6Vnl4dh7WggFx/qYMbSUTsnRcCbb9QH79YNBrF
FrR2dVohHAZ0JU9qD8vh575xmebM2d+WFMMNnEyPCxpurWZRkNXRXOyOatEQn3YN
kQH6rfzJejjhRYFEViLl08QC6SLyKlBA3e5kn58yvrXeY44POkN5g9KGS4vXX495
Pd37myTC9+lac4rnsOhPy3P2lWdXrPHsA1HIBkS1CRANz/OXtt3kFKxOh6fl1Aly
yC3GzIf/TO0fuLU2q+FvIQ17AtPzWhs9Dhx3ZWh3Hg8UIyUDGRMuM8tx18friKsW
j0j/p6I/qGdeGf83iCNmw8NQLI80UWlbGprENFLh1mJmpmduRgUZ1YjoYlkqQOwE
VUs8+GoWrvrCOQlJsXswhozAdhpDI/EcWma1sg3kglOuOo00Z0Dn46UmyY9QNwUE
uzAf+vn1pXIBYiY2VSBMOjFNACrHsznSP6Ppb9EGJmqoyb31QW8GhtqLA5sFJm7P
+Lieb7ObsoWMcCCqSR8whgyCCNsJ/jPGwTv/0f9zJPKc0wKWuWEhyIw2VYqHAZUl
4kuXbCFWtjoxRYWZ2RoKY5iyOO/oZUF7tgK5msJSnzFFIxiyIAfTsNjkthWt/M5U
+5oJaubdAJHrtpy7yYcJT1L+Aa/ymfF80xbd2vkjUnvV4J6je93loiSZHfSPmsSM
LB87u+EEnFHGazusJyzCgtbNuM/F+imcALMWeypzBhQFJuqwvxDNUzB3aSoDIY0J
HMrel/p6bFf05RsNhntOX6m1KtXYK+8MwiN5OwdQATYhoimczk2w9PUYBHw2HAuB
SYGDY0Yf9D0oPMKz2QNkE5Tc4CH+kTjBxGX2sHBOlYHZPadFlHuJ+XTvTfSJc3+E
3BbDHagkhh2cMBGB6I10VNMV3sHh6kM6Vg5ibwY+tVwVXUZs6c5uVgXiu0cKQudr
1t3rxPc1yXx2KRFHxPE234fr9OMJxrPfOHhJyjQSvCQma4Em7n0ic1c+XzgCSNAI
wMpAKMevqL55bLeNYqWMMKj9SWU9PTM9r184CFXXoXhpj0R8md5Y0b+ssjl9GsD3
ZxlAHNuKptx4LiVSggShDc6edm5Plm2zt32sZ901eiwG2tw3kroKiAVqMl8UFLgD
sSzTmc8+RoNjXAuAK5KeicJVLQdIwNcQl/fj3RH890MslOKZOgODgtNVR+mr19Hx
2h5DoKs5chKRiOWkXE/hoKrGE8Xjg0onSXgLzEojSwNE50XRhk4uyqtf5nEx0fSp
z8VLbBY914C3HkFIELr6IvdsvJRK/q2QaUleBIuysWZeaTBbsbqzZnXE3bfElfhj
lT1Eum6mJ5cWJss3S27nDmkTns3UMhQR6IbN1J7FsfamWhbGA0qqJeb2doFwXIRT
M6zbzCxfdeDvHQgZhJwU4g6CJ0nW1+sGIeVRsPQqRnsuIU129tP1AtCbV90mmoEY
q+1lX0UI/O7lKBdxenn4zQfUldK4wDYCw4In6t/VTK8wHOu0YhkQVjzZUlxaVpDE
aGSfXUrCG9a3MxqcR9/tK5fgARY1g+iTJKyShEqRpVxFVw/J+haGtNeUl6ozG/hM
fCy5EhkmbJYb4M8wOFoEaMS+JOVTpczKZGfqIs5NE2oWnugW2ZDQoTan9+FktRfP
+zvXBaGqszN/X0vWGqc0iMw3suvA9PzTMHO+bBh1RCWGQ60bHYCHGBGqRJ3ClKb8
jIGqzF6fKdJdIXxfMDiZ1dmtj0fuDs0y0JFsnwmUj4avPaTPI4i/9VWDRqmNKGCb
tSezIbmgDLZGpPADbDaUShCIk2et65PseIp/SMswze+RvxWTlBhOwjezyZIzYZpG
ctbIkIjBRypegnTQYEuROhKTDgO8JzH7JPe65c3Yk9oqLjnmxeHBsAf5m70OMRE9
RKO2GnbgE1euwWZmVwgrdFuP63unVuLGvDydLdfrwWDvvR6hnVU5Vk3u6L/U4icU
pqN/w8IK20RVbU63cfqL6E6qtcj68a0+IAW/izRySpneV31P0rd1qkhNiEKgF5Hs
YTZhOE+/AH2elsMaJdP93NIGIKgxEOmGyDGTf1g7O/r4JmETRyKHlr6lckMIkVFL
utXPiNdEXRJqCtWOCXXYgqkWdvVfhfyCCNthmvBXE9kD3YEN2mS7e7ai3UscSIf3
ncRNqFMBUXgVHh7o1TuJirgaA/cLHkbmz2FS/METXrpO59ib2rKR3XPjLLWAWXdo
GIUU8k94aioFjRmdVhwe5wPDwPB1T7hMZPZQYy4xwqypT1yoMNxi6mye7ur+Jdzu
jg7AwUXxEX4GZmzb+mR/n0AWiwG6cfUDdS2IF9BHDG4J6B2I/bZ8V0D83367dS9a
uXTIAD+7+txsYelpcWFZzvGryZSaQb4l6iMEjk0xR2Qnbu/SXNYgsIfVVOPaZyot
sKYuKo7Ddz5J5/er7+JvMwXdSwTIqSbgcNmGo79JOhQwEFFQnXghEbAa5IkVUxjO
sJJex5fmFKTJW0cHa83LVciZDBm6rEZXa/G/tlUWi41mUXzY9mQ4YpSs/ha/cALM
8mNOk5+ILmXFhy4wRPY8CuvHrsWH46RlsErANj19ubIEXLJW+N1V/gh7vdkdcF5d
Ky+kGeAImaQhwptNwL5ielJRCebaY8r5poxas0LDryzC1iCf+JWc7fiVFOWwnFIM
pQNz5tIpaSCyYikJPRYlv8sBoFaA4n2M3TJsOdPduiiyp7jP5so91kgnB1l4R1Xe
KzQRAMg1Mj7GUxbX3H9Fbm/UPPK3PiAVKAUaCT/7qjogboCTBDyN+d/JbEnwToYs
hbEaVWKoEIiM5S5y1G/apKeZMUgSjBUxg1d4ysK7FZj8NrYoc4JMhZGe9e6bJsZM
SBO4c9dXBl9wE7/+++z9z1nM/14ZIYzP41P0ZzjYC5KUldhJqhpX/0tO8bsRjR3z
L3ZIrhDoXZ1WNQyloIvH1D5EBkIMdK/bsro4v2dbAbLiRDupfvxX7NOwf0Hy6vs1
b0R2SU5Lfo8qWA4mKy9X3bxRRrm5Yz5qDAlkfZs1xFrzCVN58M6HQojyKK2mKJ/R
z3UySgRSYw6Kd3yPxInq9hzwXkrsHEPUJUuwgF/SNhMIwUL44bKa8nQ6m2JcmvtG
RPqTLztM5ses/JkObJI55tXQhJ2DU+VuQWowuv5wP4Ha4vjLs5sXVfRAxU3mrWKF
gLGv3HKfjeul1/hHwdGLui9cFCjpSsJSygZ2iNdvs0aPPzyslHmXjkzIWqWellek
G2YszATvHxDknpMyBRlf/T32dAFTujmSLxKzVMcDu81mtLHryz1DlEFaF43VGIMn
564wXY6kGRRLR8mMX2rOJbmUwu3vB3UGvVvRpWgsmx2dgvixQh7ePkOd6dIRxhyv
b3/CAnuyJl/6gl0vlEFFC+zP4REdEENFIGrnjbDgc50uFXK/A1ErErdttkQZai/M
YS9GG9UpBe6+KbVxEFY2/L9LikxHGBs1ivngz9A4dGXOS1hZoXNC9DJrg1kJGzkJ
rs8KKY4p7jBc8IN5P7hwariJyw2BCE43IPkMSMbCDEGEZ9CeiyREg1Ch2+nAJS1v
l/yvFzq7ZO7sOjzWgXl8L6s8UjgpvftWOfeRCdexZ+g5T719HBFt/eCi/1L6wxt7
d6dkO/YZuLDW90iyNeiit4cBCwMFvc0xgUCMB0G8n1vUxpdlZXzfUf5pzVmUchlq
9OenQPm7jYuNMSo4liiAynmWZq59q2kYyxcE77tczAx5k/inIgQ40zB0NqlRz9c+
p5TnPW8YgpJfVhkkALTS9h2lYUhIFniTxwAmflKvVs8bWCqBT1Oe4/CoR4+bVbX7
ERJ68r2c1+UkAt1FT/Ooeen0Q6zhhlUAmowANmW4UYeAQB/+SHN1q/eANL+9n1z5
XXtDDr9qFR6/mekGbMIROMykLZ1XGVu9cD3J36ujqoEKCS8O7mcxLq5lY7hCYMy9
cfKr4zHk+b385/mZ2VIUB1VQPxQTx9AXh6fFukC453VheVqZPkgva1p9O7rdaXKW
LIOhf6oEEcxDToRDzfIrJSqE5ybRJH9btLf4pFA4jdBc9jwna2NDnxiRetwkGpW5
x3PU+pGMHXN6vsJ0bYJaXlns11+UnUu/ZhFFjGTCaeF5KSW82Shi+h8ZJMvIZ9uc
afhvvOtkdAVcS8CLsFylsdZQknP1jTss4TMo465ggVxK7wv7wxwjfXakWgpIRpVj
S6MStadxFD7QUSJRWkefmCES0havtW2q0Q9D7/YOI/j22voiH0Jin3gExTE7bTCl
+EfEPiYizYUlB10H7ChYTTLNvvrTEN2NMYVJyM5zkSKq2xkrgIeVpXelm8i3/6cV
8T5G0CXzQ/QzSzwGWI5rPwZN08R89RDRMFHZ/fa0Ie0BADqQRXTBFO3c4dyQm3Ie
WinoZKmHmLCF31sANKHDkdY2p0/irGtevkRoTllKSsmd6rrJ2WEpPXu2g771GuGY
jsLU3V/svgzJV3NQbx/aqDfXLwwmk28A7/USRIWWfV7/JgkRxpOqbXIeAlKw4Ym8
K+6aYhjNF2AFXSlu2AF6rnk/D6TDzkkNWkpbo3L8ecMWmOYpwfL2a2ennVqIysO3
mD/mNl0lO6FSkfj/K4uyyY9WGlAvA+ZNPiWrbBWrpTVDackVKVy8LL9oEB6wE4D+
7b5U2IndqP/FcQpKBL4SCbUeuBtrz/QaACkTi3zRQ5fBG1w6/oNIC+DQ4ORc0m0I
GDT7Evi3ij301SXohH6AxkkqOrICN0Z5G7RkfFm4eYtbsMoTRHL0r9hHCxuSSNM/
sji6lNyCmpZK34akfQoQeClxsjvorkE9tsmaOgR2DUuEH0KNUI4NDPS42sBGCWjI
oA/GBkEUahBOC+2TCZ3hneoNJgQryeMHt/GvuDUnyeSqPxvuAWJuI8qy5aACPMgA
kEidkpIAcZe8ZG72+p9C+kwkavDRBYLz8winpawQreLF5lzskt6k1SYI6YbuGP+O
VLS+U8Twlfe+puH3CCN1Svg+meQ5PkziLnCyYzWLrDKi9B9wXttffsXm+Fs7HSu7
PdZJvVNPZp7kx2wktvWtiT0bxoFKqyar+EobHkHAKdkHtRffmFDRaecx0oLIfCwa
/WEeUTfjT3bRld62ZXqWEyyhSVID+O3ldWwccy15+OpvsdS2WqgA2e1seMVJ/qVY
ZVTTwz3ef14rTNrJxOEU9RZBWtdCBf9dT5v2NknWo8WlLg4tJoH/3wkSx3EftbP/
eiPrCqrnqw8CDNBll7wiOidDdn7GvuQ7oSqToO/lLqPaIhyDAZbQScv7hOkYAeE0
UYwUsSZ2A3CRxzSh+lBbLnqh0wjmhWhPwu1tBTlWtqeTX25CkW2+5t4cTnC099xC
Ae1AZuLfsnbDSVtq2RKUp//OC86X+XEuVdWqqKxtBYurw9aWOzGYaH6QPZ3swe1M
XOFNUJIXDTz6KUwmM1Wq4+aI8QYwzpGaiCbOJ+tH4UXfJ+Z7ay2Sq2KmJeVEUBuO
PSVTyRvj33o9RONuqMpFc+D/75tEWdff4+zpeEgSXYpY/8ZJwWLM0FI0c6cBX046
kl/adzr+mjU1h+sxmk04mjy46gwkQ1NHkob4+9oxijn+3fH07ZPbvUxUxvwtIOes
tNULM2+8eByvToy4XKmAWgTw0CQvhzc3KIa+R8TtiBsAe+DW13ltYthYCOhFZLxQ
hpAOwvTn7Yh/b0ArQyzHxnRFZCaA1pco6RSX9KiKUquLwt3r6yC8DF2gY/U7z9SN
P8LX8SgR/m0+UrF1qdS717N2X8XYXlyvHy4/VOgVEz9oHylm1bDJ25Gb/2DMCTDh
29aO8igA9tmM7dFsBpTcWV481P1cA61zWbSX8vDR4ezs32U9pxThDZ0DjFm/rQlg
uwwK5a8hQ1YD1lBkHFn+msra+ZuZhBgZVqA5uw0VZtEjszOf9cg8GmkjCdLU4yha
u9n11NSGJ2UJ9aX5J38+XI2yA78iEPZIkgmhDZ8jMtQsR+4Pf91JeqzKN+NYSoHE
a2uvXk1DN1MllQ0NNpSTcJxmBeW70RghzgOfP8ewceWVQGHD+acHL15wssbwxkm1
mG0QyV3AE6uzC2fnl06HjRJzOvUrJ1WI4+djaT1zDof3BTf8xjWHTCdVOhFjU0it
jfWCNEfZ4D5D025paI50qkKrSPs2rr9xZBhQaB8nhu/uPBjgM2RvUw5shBob+Ug2
RQKvMn1HDjYJKny6y3+P+fowvSpWiTg1szwg4wezJCp0wYIVWVZTIkBhYK4klmRg
Z5fbftwx5NZo1GxJ5vpSSMIO5kQQM0s2JkA+0pKEeCathhYRGNKEhZb1URL/lKb/
wQ8S5Hu0nE2vcuOsDm2G6UIUPuvrnJnzYt8sPMFPDQv3bMoPiAAK7O+o+6FffLIP
vjtM0B71TQNIR53+3oCxvzHN6JooUZKsCI03Aci0y7mduPNgR6xodrDlKa3MsiBh
9stHEbW7J1c4QeVUj5gjnnilRzV4L8pIQOAsR8Sf4x6FfS94ifYwEKAjXGZjRqSa
iu1Qa+DP9VAm60f1OXntgVRHDMPSODo7Jl8fHihSTRaLJz7LlMdsFFVj/w2L/KT8
hr3m2ovV6WR8mhgkmuuD3W12zF86t+WxmLZQ5UD+oDHrf++W7o8tpglVGNQMDPMp
o0kXwPOzu6BYlk9dNxlJaQrmQ/E+ZULxNAT866uH1V9gAJEheNp22tH2/1QHPFkr
vuzQfUt42d6fCLU0VtRERLY0JruqAREbLFE2LLwzBD3WO3WZfqZh5VelXUThrCyn
dMM/qPHXmJImqY8K2EtoFkjPqICXhxcrU6uj3lu2/RXJfRElkTm1+qh9XI1mZQbS
vD7uE4/A8DRAJcSpu5ChH9QG1b5rpv/Y6XgDNwKBu0EOjn/yJwn3Rdxx5cRLazhN
h4jD6ztPtGhArvjuxWnJon/VJn9T+1xLeOLI2doQaNLmrMWao8WMjFGFO2Dufa3J
kPbL6L6iMlcGunA3bDbuRcZ6jlHFp5RnL03oTHsShugiTkAk5N1H9PsJrLQr9EU0
+BC9hVORGFZX3+sD4oHDLo/RxojxQ15rOBY10ZkIoVwEnvbXvMtnvzxQqVV9u7iU
msZcN8kwVs/9CDSTm01fdR/Oh0TNxTT1p4QvZEAziwZsKpbOqB4zpSdOjss9ezFi
lKwKah7OjVOUf3I1xejsrcJFx7sebFP+NcWroZvQqvbz7AaMHPb8MSRhrRGRuU4W
TfzYlsZxKkV4JSJtwz10BxNLET6bIaq8azRFCRvKymsfkcULle1JBKUV9lwdeZU9
RVI2bkEQvoKpqTYHytFGwr1tG+sDftnahW3w9VO1b/nxWXrgLE0Bf2E43wKpOMm7
FCh6BBGzrRv3hbKL9HgscQOna87WbKUxGOL0VJxhbXKt1Wbuj5m54qFUtJPhQ/pK
OPIPL7w76oh232sz9Bypul16gK64UvwClFJdSYH+RBOVf+rjGj3jR37rvObHusAY
O3CRn8vWVTHG+SLmuugPnV71EC2epKdH2qbu8M+UQ7IKDdoId+q7iapq8GsLoH+G
gEP/Db0SbbEwJJb2zZX3dC+H9BteFtUpT51PYb19sz4hlL5gFTkn+zY/aQokU5g5
Q41289nPGIhd2V3s/afW/5BkUQlZib7fl8PfUpUp52OEFXAMRhIXi8uuY3ANK56J
Kh3D/K0zig2s5+0YEGJNGsVwb+xkCZ1+MrdCT7S0EZUPxQVG67XHcaPvcaAm7JA2
w4NyiYO3xh3AE2hPM1DJrQHEJ17BMcY7Q4CFQHJCSkOLic7+PItyRTBw2C/3AX5a
uZeWzwfaFsTaY6ISYM7pYxd15gwbsk+07UV2oHbQipwry5rfI1U/PP5NktayVV/T
cSVyZ4640BCAvKmXeS9bFEIEL+lb864cPJu1zmsJlIMIXSXKoi8sutz9euOHzt7l
IWIxFasoGMgSIq02rC+C0NDG9UB4fzssO1/Yg1qOCfgLrXeKloJDAKVcBZB3px+Y
8H5jWN6Da6BIAu15Jg+reZrdgae4tl9UK3qs5F7Ljqa4GBhbAgNLdA700Fu47C3y
tvRb11ci8ob8hK/VF3DQZLuwyQzhLoyem4VXBV/bPBERB7Hi6u9ZtQubUjYrdQSv
t4PDTlu3UnRLkoZKRyCScA+kp9wqFdaWAS7ugxN7I78hFlHKIUuxfrURCVnXxcbL
ZIh1wATUo9Ahq2A0+a149s53HUqIRYdLiLSL9AJ/hvHYx7GJ/kbjJL2cCyrcR8M9
LJEv7o5zxA5VM2nfK/5qxE25eIFiqevjKTnwNSVnn9cbBUuZLJIRb+YqU1yJYNDh
4xKvIZPshK3gdflyGhDH3a8JL1QR/2t7E8DgBuUNgdl8N2aOSK+sFA9RsvAkueZJ
lMvM1JQcmkVBQCEbjnC6HqUBSaL+Dlf53sOEnAaMrO9wR5lcA0OW8oXpxmMhLtiS
nWpef3TUwN92eAwBOQBFnbDXz9WaMhMKAY/65/5oAlZ1+xkD4gocX62lxmqoGcPu
8ltE/vT5JBKBeclKbnCtXZDcy8mbmZiT3C+uOpGvEuDfChF7yB/h6cOD4Tq+IZMX
rcM2141XXyJg6N0+Y/9l4s6VDkrDQ+n3ZGm1LTBTQyioEe8qrhVwL8AdXiUXj+Ar
lz4Zjuy4uzmeEDdefFTpv+7xZOSK/kWPrlIY0D3Au+OC/9JJJB0TN3nA/q7UWwxq
5bJxJG2hgF0BsdS27XgJo6KsqiXJYJL3BEC9r64nEs6+LY/v4GtNCyXRNoq8HkY2
MDFE9ogqx9HBb6t3Ft0ym3W2KDUueh84wCp8CR++9Agv9Jo0BFhEpEXQYckw2jqt
LqessmvriwXj+urIbhgrYhsA6Ku6MPv3jcZAjmu7GaRF0zYmYHjTe4ohNrEo3A3z
SF+wlNd44ZrvTWjjl3YLuopuWKOonGpRCBI9MocMiNyo/4STDvuoRhfWO0YR43Wj
qXKLAEzydpTuVKmumN+dVGaCBwix74/apCxsJoP/MCl76s01qfWeyjEDkRpzLAjo
Q/OovTGUqvjBAip5XNtoWX3MXR2VXjYpF4VssI/Z6j3cmwFuAkaZ2HZQDL/MGwKk
g7vGCVXPuyp1QfOBcJ+roIiYmmNon12eI8paCHqXtWg6hX6d+JdXgQ5j8t8poPgI
/bBaSxGwbIFo4LN7j7YTRjeTEEUFLRqNMq63qBMfKuewTuGw49IRq4iGw6Is2ytf
PEERLuHSwZjJQmL2VI/l9602xhyE6Fd0W5zLbT1igx/RPdtg9XzQgHTxaGghU+lU
3VKzd8HqcCRa+sy250Su0zoaeSsVA/Qni8TgFE5kWA3+a3MoR6Heb+fjbfV18TUx
000j/oKxSKcfXcRi4SxmxZKYCHIiMiazgXybWLbclfjWurMkItLqpGp6rH8HF6jZ
/qqdaDlBaPqdvF5zZzWAXyFEBuK355NY4dHY6xTdMcS4Rvizl874yx1BaaOH0/xd
cj0JMpkIG/oLkeeMAfaCMUdnS4bWUoNVCGv8Y1Li0VP0/t5V74N/lRquhuLQXCiU
KqBCHknH+stIMxs2uEtFGs1eWoC3EvT1Wq1vn0uQM9zAlKc60N4WPQJFV6q7zdUs
r97HWT1fd9TI4A6VIK5YlAWv9k/xCZcVkjy8Sonv2gpHgRFw3bezSNU1CPtzg+b8
RqpIjfsNtPqF+Nb3NxQzAhfZ2mTAJCkT98F3aLPazfWP2RtjqBbyTdGZignokMbD
/9aQwll06OtskYKyZLm45bTPhkrZGcbtljQWiiuRtUk993jJr69w2VmBe9SbgdwX
EHoIvHCR7OZ8t0ONW+faBMur/ipkKFguUM+Ho7hzb6ZhkWVMKih7x7EVJ9L7pZKD
yvl3FHJ4oIRgovgi1LDBd23jduCYCSJX9cx20Y+meDBs4NPKfjxn2vQXI6WFgRFo
ST6tCWLlMb9aKsVkQZyFs4t0JXQWFPJx6hboHoEQS1NcY75L0aNamAW7yaMR1Jh6
dBGb2bW/mPoJ1GfLOld7qEnI8k1c/V8RT2L2v4mYCsOL2tsUsXqZGTVGuxtbBVaA
hyjASXv9ceqUV7MzsZTStAUf6Jgf5OUNSU0JgwJhvcNWXLxUm0YDSUco5TJ+TKWo
6sd8ICN1UdlN2p6g+ajQCZRcLmMde2sR8wk5JUF2XwORxw9hlvXPEWJtrgluoTKt
IA8YhL0UvbiccLPCfvElGSBtL+rAqK5+31o4Za0VMIgf27Djn1rCCg3X07IszFa7
fLN/ky5GofHlRLZR5eY/kuub1dsFGfNh8njkDMMCYQTugFpRfwGRtt86DpczJhCA
C5QW5ZD5V0L4wOH4y49gXdX/oUk/V50znNMN/bHX1NWnunmjWKkniN5Zo+He+/Gc
notQ12S+Sxi0JJapu0xzlSuwK/SlPc0zNYLrVUl951Xi07UADrsFjFcEIZG1w7gd
8Eb4cOSQ0qXgpq3nt66/7b5TQz5ZsatGyCiBauYTx7b7q8XkQSWpvocSpsQrBauf
wylzTAMQ3ccmrl1dS/BWidzsKN2Cj5N6byknY9wF8a0EE49JOUjBl/YVTOTCNTVm
oNXyg+dmQrGLmjb/qbKyzewRQPEfoZR0O5cMI4W6MnBNlpRvEIjU3Ug7ng8hpu4R
X/iEipGB4JHZzEAWOHc6pOULWTh+/ujZ8vOukKcKgyb7UOE1End4qkxtTcphVxXm
TpDULxCayDLOhaZ5qu5dMMrbiSBogGJ0aTZGqBl8D88UNnGHfMU/SpV0ACTWxIif
/xvCvEa2k2kpeTp5HcJFABGL76Z+q0ezvSx27hMsiANxeV2DtpgenGPVaVvo6Gml
KWE1ckrOk11UZRMfGfA5LqxtN0AYMKgcQfw+EgpTVpp3iIUftouXkcGYXNv088NT
w6ULiC4tCbq2QNLyAGyztxPkjmfhg3D5UF017rZtDycm6ndULdJxC/sx6csnzFtQ
6TpUSDHK8Xei7H5uSOouqLFA7ueo9UHfIADzNuBWbwh5LNwBzWVdav27aOu90EYr
5Eqh0GWcLsqWwbtVebCCQIV1vG359cxj2uhHXTWOSP6y8eFD9QTuHgD3CGuHtqGg
VP2bbxZGgvcCfAc7VN3Rp7jIw7Otdb4tF0LMQ5++OdxxQh1EE6SCLsvH+7F6l1gC
Atd0AZqFaI6Ee1PyGySZ8WQ4Kr3aC/rB2SYusGKTdbTlU/g/O5Y8MKcDhDajpIfO
p2NnKezRyicKob7lJUhBZ5zLIAXQZrjNFmAd9YU8GWVP8U+1lgYz4kYZbEAZ1/7H
AubdSrUxPuwdsIh7aN4M6pOy7WHbzExBBypUQWACQ2Q7DOu621WCN3SovSKHM3qB
kD+EBInKhVVgAYtw9bWZU6eCPajpqypmey+VURwgab407lZeLwlssHgTr26/Wvvd
coz4ShnuevVhliaWLKwzDswEGXT7IP6Ga3E/Q4LeVvDXl/Z1+BwHq/jNOmWXYd9a
Wiv6ACDtA6QlKfGBQhjXJ+9h1JP6dpEM6C9uShjnMqgNde9tb20mqZdFGrlMk7cM
eSNhVsTNOAD1m9mVhPh33fp4srtFzTaXbuyimv+juHljYQSeszKOyW4B1+imCmYD
OtPhxC5QEVnRcGwJS0uOfCW21BTiZUxmCBUTuO2CxkiOSxTtqEmwI2qjFfEGK3ae
F1b7sWHlkYOwiceY+CGkH9FLzgcV1biDFznRXuVcHyRabbuAaP5MkcO/VTjBgKGz
wCztT59JoLb8VEVCmJ4gaGNzVbW1hAA6eP9t3e5kqw7Ceicqu2vseU5nnRudxPyc
iXMAfJLRveXYk13zoYP3h7YNtO7E9V+mo1XUOMIWqh9JQnsQGbxNJHcFmEkLzl+l
7KlGQbUTtW3xEY795KuH/glccOENbjmFUnrxOBxc6JlEuUzCQVDozAP4BnznaTnV
E62TsQOYE+6mfUC7hLV+X6NeGUrEg7K/HFtyN+cTWoOTaPdNe297qSR8jkhVk01m
xhwS9fijLvyTuXbKtY4NTcc4Qd8IwP8vSUKZ6MnCeFljCZN46xsSJZPJQJhCvXMt
fVueHLutaiJYhBFPW+s4pYAF591TpLGMV5LHttdHC2+zv0sLRbRhqvXx2NW/o0Kf
9uO/Pr58TjLlKzdDrSFkdgvS0V7gwy+lM3AHTZZOt+XtIUrgYpEaUO4rA6bTyUX6
YKmE+OComZ9JN9eKhfFNdVi7rviuNMlgUACYPAOIg7K68/EKX4WRbmVu2FoG5N3I
QlbcwwKVsitEUm4x9sW6oPPeLCTDJEvmfWFdXJyH9/en2vYOKiqOYGMbWmyawZs6
4h5yHRU9dY5HT0IwEikbcZRoxQMi97cq9kHpGiBBXzShWUW2USmlqfN94yHTSG0K
nZ3DjRYZj8z/4tSzyl4wUyo3tszc0DRigtSDjqpFFiHO7oFN1dhrXQwND5sOr3FC
VLpl6C2FTkTC8XY2vI06rAElW/quZG4OJ/v68A11gpKAl38E9IhqB9UwFdlXzXpP
2A6mvNQJ6wkBoaHnaThJsz5VrD6nVNmGp1LXzbdwI7cUssCFFM+nDk40AkUZWy3u
14j/OWwFEsmrAB5rGCtsUb6dyMxnlZfDnEQrhIp9QYhQid6y5+PHiG4oV1mPo8UH
hWMzW0wPxoM7xNiTMAdRPVx1cA5EWx5cGWW3eVZLn2tE4IaoBJJEGkh6ZLZUiXC6
87Gk3/ZVKiXbzkMThqgyK1xKu+rU4/KK8zCXZiqUeH8LUDyMK1KqYJc9R0qxIlHi
oYgH3lvls1j4+2HXLA5T7TPkShOcYmw55gnQvCxnm1UwM/tfX4Mn198kcq7h6PGZ
gF3DTJ3tmQBNSv9iBeiRRZCCzJ1bUOlIelZk8bY8mlU0XzmFtztU3sxPkIHoVZod
+D1tIcLJzzFZKlzeCSSe2g6mybYCrRkQbdFLxv12AjorEIGLWVbrleoYs38fvYi0
YTQ6jCPHTcrumiVUxzmBWiPgP1M8zpPoT8WhdAiWEGP506crsWkx7D+F5xUqyIbl
rhOeyvj/A4bRxjEC0PazqPEsBxcvsxd2mHcMWtWQ1e2QZI1FIM66VuAYTyFNIyET
WX2sa3BaQ7QATOUGk1ptAKKSArNEC9GjUiKkJ/0fzfBTAX6UzVnoTA/UUYuY3fBd
XXTCxGr4RakxKeI/v39CvdGHP3xl/OCknEF39T1ZLEUA7DbQ09dA84Rymk53D51i
/CJ+88k3ORBk4krPfM+VbngTHyk1glI1ICa0peOS0zx/iuxKG7b09jVQADTq/z15
CuPH3hpw6H3cKiraQgJ0f2a4Nk6We3XAMuezA7X5zdurwaDQ1w9uQtBPgZUugGgB
hknZ/qojoXvkGcG8GAWugfhGm/n2I0XktBbAOjyi7iYrErvnEhnJu+/SXn1H40XF
rwwRsjneIx2RNsaL3ayFN6Etiun0Yg7sKaXyO4UsSHlG1HmE6892FkBepZnteiBC
lB6+/4XZuKjsUYJlW+/tqBV8gK9DqmDK0lS608vWP+enxoYz94CMltVBKPe1YHkU
tjtDdoON+oZoYz6vZdbg+tw66dDbNkZXMzUOrYEnLOwMRDn/PfSXmtj2pVCH6JlV
CW1zt2QE4KSi7YGRiYGdKZhKK7+FVTqNWMsR8Hsw5ZWGknmtpkzDw4Fpn1lTxzLD
HjmwKttgSwkW8A1UgQAbsY1KquRmTsBhvswOL2SG8/ndBPmOpe/e7ZWirk+31hG+
vNW0oDkMMCtaqe3MvcTy+Zd1PQD1FW6L26up8DIKAjT9Del6Ac+XzDJUd+sXO+5I
YzQiKUnbmn2lDQiQAaUzPkHgNPRT7QkUgBIwYugjLbcWFL9GL44pF1slIhsBf7WF
YJke0/VMPWju+qMv+ewUqJ8ZKG4xsrnQ2f2LzUdgc12cWfxWyU0Iq12tSwJJoYlZ
PdFxmPOrq0YXJ79ubJ7C807qaRw4SNmMIWtLmfirheFm0Buv2s4F3ICt+HPOWRvk
TmdaQSVJTu1DrBrpS5YhPrvCbEZ7tmx07+Oukyr3jZergkFPV6thTrHGs25E59D1
wdWVLS+aP11wInR7mqGZVR6o/TgFyCWFNRDHw0Y+f7n0xYH5uiZ8axQspV+PWH6U
vrOnAGx0V06vqaLDGYVbXRuOM6ZeO01es78DqhiQmq/VWQPOwrueiGQdykiJ96hf
LwUHbVD7mO8q87fO2q36aLo3Kh2UKqwfKgTy4QEAsTsfutEegh2EkVZWDw63orJw
gUU7AZr1DOjjgP/i1/wfNf3+/kpHWP6ZKdNcC/4LBtJj3vLkT9rmpdziCgsnvntU
DBMqga0VYM1YyNI17q3P7JYDOTchNF/OnbMoitGimRwMy3pAheLizPTuU/vxD8VO
QYlp1mB9HMtK+Az9lSUqqlqt0N5t77HvuP+ZyaEcUCdtVw/le9lO9Lv3GhVRbrA9
p2pwIfDBdgO9uEoD0P12zy1RdmHRgP6jnTqrka5OVSI4jZUx4AiDPdPAsyqUvjFY
1Bxg1KC6g/+N26RuZpBOfwCtqDonCjYcYgdkaVCDTR9JVsM4THondffBH/Z5kWzS
LK0q334eL+X5pAs7MMAZ7JUSAoRQTkQpHVgng4RmgjY4kO0x6R0uh/bSv8drXOY6
DoeIywDSPIQq9Kd+cQlk7r3lzNetIPxSeE9MSQE0juQcbZtEPaATJztkkrzBCnFM
B48OmYQNSn72q2bv21OAAanYE40f7jyw6PGwhSZoADM6olXNWvHneb6gvipTdV9+
Oy38eRI7lWASU0nID549DUTWox9WwxkJxwizK7K81S5nRyCb7KdsHgQ4sKVJDNfY
i2eQYNcMuNiylpYBmwaylBIothStu2KEaX+HRW4BJQNvpqeIAbwu4Gp+rZUtvITD
n0o99UYsPFZNLiWdH5dUQaE9Xvot3FP17RxDI1KvpW8FvF6e1xySlchEXZUk+CaL
4ZZQlyDCCYUapfOA5vWhbCaM/6/+3LCZJpXYLCor4EidP+913P+sc/+9kvfdtqEg
PrTLWfJxac+6HHDNPvJbCY+ZcWa1u/8zqUMvPc00HfT/EI91iAoHWyfQwTsqVzsr
Aurnisvd/burL0d8qmoHQsslgdxIMYEXNLSeiBX94asJJwnebMppnYD0ETDRsy80
I+Bqb6XfALJyuhvlRr5ESyOrCpzAos5PXdPFw+MTbc1BYebf82OgUs/lDLBksU1y
qNp/82aCdr6pRnhtCSJxTqKgk4D+Q+DNOvxv78wXolqez9XALExkdwzJPw1KrV5t
TDD2ReB3t60+qHa6uMQnvPSWmhZxT65cQVoUFhGIrvPB1twiVfLYfNhqiCzgAAgA
gYpwWRMexrOIE0Uj9JtmphfTxtVYrARmntIVT4y0h+gt7ozGr3nxPmWvJhWaIiwv
z/96+3GzJmHUkmJG3bF3qvhQ6a9IIkN71g1m3Oe6kuGn01P1/jkrXs1ToNQvs1U6
w9SyiF9lYAUZILuXGLCy+5+hdr3qG/YwQ5CmVoV48A0GQQLtBJOzS18mE4zjVi//
wg/IvBhrrx5xscskjXvPecyC1v6+c4RDKcCKF5LfJYz6CZRaJ/VPTOsHS8AENdJ0
busa1yF+U0wYEAlTzcCs13CUOU3x0Ry59EVVWJPwh8MIpZZMf/TxE2HWJ6OkWrpi
qocGF6gBKA99+SEMLUxu7oWUXymI6iNIJhXeyjx4FykLwwZJ8mvUazxRjz4aTqjz
0QO6fglC+NIluC8G/VKcAXAuRDQtxrK/JWDnp2GKA23RQobTAzaaTztxlOweqgGb
6jPIw7gR3yjAGdOpxinxdkxiME0aBo1aOCj8xjCbvgR1kAj3pHdUcbywgtaiLx+j
BmBjQHSsULPwnCGPb3pQbtROs6svNXgnmG/cdxx7HsqfHC431yuYaQyIbS/KNXnT
zYGlKA6K8Ezm+fsMAw6tE0oSw0OfyRv3LAIUNDJiFwfVb2RyzB7WpJiX+Jde5HFi
4pDtbGWaij+5hCwHGIjOb3et3Eyi989hXfODADWQ34drkvFTJSrluph6Lj3HRoqq
9fatLZ/hvu1imt+kvnmx67OQJL6RL0xFRbN5zKKWC5ZEmEKzS9SmJQi+FCglPOA2
VNUa2CaaRsA/kzEU/HcMQnZSG3yhLCryNwu1iNaWxV/e5hEqhrYvSapZNHTZkZ0N
KDynu2EV/obr9FehbAgdmanLA1qKBJAAFV+nNXRb3dMH/41Mcn/U7IG44rOLvdFy
xw/ld0owUlR0ugyPJaiLzb2+hn90KgCTiow3jjhD19eDCWp+1CBBsTYO62qmiDbq
Luge3P4JU5/sIeRHddsNjT8OM/40x+8dIDM8eI3TWxXH5PDLWLMOq1xxJh8B7JfL
Z9x511Ehr0aprMvYtYB1zDwIVnH/GH4hi1x3qrd8EueJyOrhTVuBTiOrpPCur+Pf
YYLdLl1/MvGpy8OHC/war9rIyiTFfXZzHodicRefOpDF+XYVOUOK2x2iyKF1ciEl
ml6X/8z9k6PrxRHFMNPzmPIFwv0+ys89nsx/MGUhZu98W633sQ8lL6m49PuV28yU
W+7sfldVdHhv+0XBtc0pggqONCr1QDxLfs16ffrGayprod5Qo0iE7zdg259UN3P6
UejfH4CxyIRJiS1TX6sGP/7chC2IbzcjE3LD+/28lNPStXRGVQKA7Ue47xJ0Bszu
zTOdZ5p90MJKTi1cdy2BlYQu/8XyJqGLfr/tZtxiv3fzx+4PHy3RXS/aOqm71DZL
r2J0ZOOIb4Z9nFBCwAdBDzCPg/tiLxDtkjxYZ/eH7Cw+YnGiLTE48Xi7Fxkjx4oS
IcjHjg31t9+KE9ijcSbt/V4vt5urHaaOjvFbBcJEn0gdGvQrRVGPPrPFlhusAyKw
ecB4rnzB3V6oXjJXX7MmhH3j6EO1i2i40HonkPaLLorR3EkCGuSlF2WXArU0YcVB
uW64BylpfWZwe6qsIXwS138Zf0WyVPd7jGknwOtY+y7RG7ftKALxuzC5mGONwOfl
b182RUm7AJcCW+IqYSNNNVOwEIEF3m2sCv8N3Hr9eGIQ7cTUz/KwjTBihlLAoXXH
bc+iJUSlQQDdSOmiCOltaV5XeNDMD0I/h/wO4r2FJVMH+PHbiXdyEPnn24g360C3
MaFFySLlcXG2z9ZSgDQl1zTgXcKcmG4ywbClyxbShep3KaI8xKKeezRpVyrL6SBS
lUgsWiGucP4q4fjmLaQH2qViEmd14rGz6paU4PTuJi57NDp7PeKka/MXm6/fLirh
UTzPhwY4p/8pZ9fSJKJBQKltemWfvVeiyI/hN9Dzl7gg70YsVxAO0HsYUrtwm6xg
DHwBcdK/jORNqx8tNS0H8vkOWy5GeU2lBx0K7AFZwDX30SR/us6Hrm9i0FqA7Mhk
FbOEge25HInsNTbDc8dip5XtQH5xStlQRaI5GkuWEMuQ2bYuuYFUmX2hQbvLKWmD
JXITID2OinzcsxsqxfumkQQhEb2vxs6Ymr6vlRsBViF/cXV2oUI8ALm5c9pzTULx
fS5Nwj0xTbSeGZFQsRV02oww11aBnemsePu/ZHNjlJ8ansl71T5WvDpSZLo5xAKt
knHw/GaeuHZe40UI1136/3mvw3beSFmY2jJIS+L2qax9RIbqULRZecfM26q+C7QC
e4LyRo1bYKMDQC6roW45kOWI+120fFAOOgBX1bs00vuzkgOoS9bN2jgvjV+DL8Qk
Q2pADBae1V8HdzLWrcHZMYIqvdSopQpoxR5KnIN9iARdu6l3YCLfsDSmz5213Bp9
BwrqofcWvTYEHPCIC92r4nDIZVCfqsgOEmQe9aGH2afl9WAJy6Q9u7wsMneuGo8z
deUSkP6AVNPYq31kJQKmWhB8mHdgzw+5jLDs/QgyJQdWjAZMtqqD/ebSfHrenJvS
/RvFqOzD1XUxSOdaU85ehELKRTsy1IV/99J4JO2Z2m62dgWPO21hascINIyXxmXf
SDCf//xKRRSmuHT7vTAdi6GAUZCSLsGXS3av4UZBnajMSEQJNACjkGCUQ7+rMenw
sSOF0ZJ4dSjZNH4n0jVShbBSBBeMMJ/ZX5H8qYZI2fdliGlKYjwQ05bM4hyiP8ZZ
Wb3XlUZDBHGe/sLHyl/RtkbbwSWGjVk6OGCg1kxnXQwNB/i3vX5HR/Nsy2PMBPxz
Enuyfm6ovFE8lb3mL8yyZyihHTZXyfoWxIKwTz9zwbgXSIur4zM2jPzo2R/e4hEI
osoV/stQ32aXn0EEaVw42Qy3Eroq8C93SHkw/PhI07ehP7biSTJF5ncnRuHWVGfu
knq4bJFKxO9S6/uDGEsULjg2MSmD76YYMX3DnoLufPO/J5NYZgcjDmP5cobFWxeI
KVheei8QhzWc9I10BoAuKXHgUqvnhDLNMU4rI1vsqpQDisI0OqJXr3+GNokA6uq5
vK4sAnRyvr0hJf43hf8060V6sK7iEHIil/zf714+PqBygKUWIYzPtG9cUIRT9T3Y
FxFGSIgCzGE73VQjSd03jpAd/ytzvknKRy3yg0/LNw1HEu0X9Ypo5IoJtJhnPdOg
PTuR0SVxviyrxLXKmPj3Lqf2lFq70sbcNqfU8AQD2/D905ZkcMRzn17U6+hEWsfx
1tx0OE1RIC0PZ407XUzv8k4wzJUst7T2fGc7dpPWJu3GalLwNG0uvgb0N5n5hpy2
q7ON7J/eba3fKPaJ+N9+ruFfEmF2/VvXlU9pc6ylZUfatQzrnvcaQRNBAWkVosz0
GOZnzmrIyOssN7TtNoKNa5L+zl05vpPOs7PD1odRAqFSbDYaocJ8BMtcFP8qM0Sy
uXNsI/ITkEcntKzzOJ8UBPwuOV4SLMuusNVum5k7TIkdHMb42BYKCYjoTOh4czFe
c2CLaw7LqdhM052rlaevNO5kkCB74oy895RPH7WFjzNoX/rwLEAnqufzJok0+3/p
sOZ1LCZu9syC3EP36zFDJR2W9rM4r537H9SfHpDFFuvEpdoxwp7gCrO0xVcsfKlL
b/fSmDFAROjniq6mKSOmrpx7jIf5Hl3HKlKAdHCfnjvEprk/O6qNemSgHWzflmiq
cvOxi/miksMrmfcHJp/4oOWXzMYoktK346+28feP97fqLkgYamUR/lprEkKjNNE0
bsf9NyA7NMoyGOGXAEWLelgWbRqT01JS1MIt+OzSRHqoopmniaBlL7VnK/XP4AhQ
VMii0Y5hIVYkb+xNJbufK1kV9Oj+eZ6aNClgcnajz+wP6rp1sh37Pi1UXNf16Oap
YWptNTFCTYsU3vd47X/jnu/vewRr6Pmi7QDF+8kntoOVH9Fcpv+12WKbbRXV4sSW
HdfZvYVMq5JoFTftMy3UvP1bX6LQd3yWiPX6kgsGq/2/LlqyC+c+olo5WXMiao/y
f5PHIWwgThTMujr/7pcJjTh3gQ1IktTALj5a4ivIysSTKv3beWRnBS0sHHe5LNjy
ax4V2Cu32l4Xdx/C6+0OAhMoXBxwAqNjKay0Q9lwf8kYhBbwUoRN/xc1eXOW6CNh
LNQcpjI6WwoNZsBahPg2rU8pPzd12P7vNbPpFt7Vse651cINntBCotsWN4u9Ul9L
z+qVA6VmhpEyhkz7zph7d6+Zcl6N7AUtRgbdYbf/IgzQSIi45Wk0WVOnDZlOfDJd
uKlvjW45+CLQnJg+/mTqyyU166WTcV3Nvhn3t/+RNueRZGjahN8fxzuddrT62pKG
B1MDNRsoIPUI4K1kic1Sgmk+hKXCrpP4pz5tleO4JpI3nivnfRO8c5O9NpPcjjeX
IVyGa32FAueI5cbfksmrubLNKdtmwj/1CjX4yHuRkArGoTYrAIKbuEGDqO+SAPjZ
QUfprlkQfKp59smdNcftdGrnQd3TQEB1CQurGOthC5/ZY5xivRaffoubyS7parVK
6T9TDqCclFrNvZdK/sEFN+Fdr7dOObaG48S6qGbJlavfBHPavu3PycxUbUaXOy6J
NKX9oIyqjhfqObUs4KDj9ac5xmaRS/yxfwT/ISLSGwoYdiocvuqh1XSZnObW1jaB
0kNUrB5wY0k9hJ94zvfNy5EKBJt+OzRBcEQWGBojYdH3+7lsyLDaZ6LnRnxDQlew
5wmpHyvgjqUhg4R1PdZ4ZAonJb249GKCExA2+2zCVqhG8VHaXJElgo4wYscxIfun
fyindq7MRQN7BwDVnzy+I8nnkMX42TgC4UNQpo48WFft8Nrp+c0kbPWKI8n+C3st
3n9cvHgQNMLt7vd+PHUy9dBJpHUXBVm4MiR0ltTB4hCSThBgCIGQce9bYYMrhzyZ
bwWL/ZXX96XHMNA7OsRsFXU6mI1nd3B30gWuYoRuqkzRykKL0/bnVly5kj8m8WKj
7QYxM8hxEZ6cwzDn/sCQbv209b6uIrOuqEX5WemadFVNtxCWn2z5lSVWuY0Sv1YH
RhdvZqJvqCzCAmB4UAJj+CHoQizpdhL9lzTKtlOJf5tT5SiFAeDN+YjVvs4ygFMF
6klqj3cL/BryqXTjTA3Ks1Z/bDvyA6ziT/Fo18WdqDQgQiJVdZa2czRhkuArovAq
AUi+b/jFDVSb3TqS7EZ1cjXlJMglWt1VFkDBmar/8x/QFRWc9LHcHJ+D6IDjskmo
ApOVUGJzjubIdBgO4cZiPZwVsN4PdFln1l6bcYL3xNBfRY1kJtyD1FNh0y/HIvxb
q4CdgQ4GStG8mfDPTKYIYKsmi/HCWVg81mW1uPsJzcAEQdY4bdYwvN+Nfjr+40pS
MWLSuKOAq+UufLJQ0YXAjdURQcms5IMsSRFJU5q7+ijZzA7k4mQORGes7yftFtb1
i9H9ykn8x7QznFaGKJX+iPC1RCl8CgpAyU7uJh4VsSrdLkVMzI7pgsYQWjpjubjb
f7Nx1+79JrVMnySwpaTGknT0VTh1Y0BzHfmskffWgONAYa8cy4HAFEobS1WPG0Yp
pNx6o/uEMu0hnFzn1rQnQy7mzGodZDDiQ5hZI8q6MbLCaQ+39Za3sJr4f5tbhWvd
rq9ui5WDQ/mBUbwKTY39NBLRTs1DCJyXLaqW5ALa8zPGNrIvbWlF2braJ3kL4fBW
QXQRpjep6Z/X/La7SrTxIUyDmHoU70JE0iiDH+hsB8bU86DMWjIo2SLnYQKw4jQU
8aEdIpfyiBqgMliWKdlcxKh+Mt0G82kOwLTuMqvMCdf/gFQzGDYvqw945/rjskmQ
MM92/+SD4EoOApExdMmATza4osuzSoZ32bOb0vasIdx89isbavyAAWgsYJx3kMDL
aexvRTA/Xj7RNzbCuHjEPcrBg7s+RykWM8EhKyq0HkSwvI5vBLLTRiN8aZBMQHMs
bFZWywPOA5wnAOgsvKykwzq57k7+Ci2+ZNC5krQafEhZQYNUj35yGgZrOFyz56Wx
qkd9ftgZnZBIoZ69Zb4W+75YQAeh//SndRS8Wj44DYZ8ThBDDzLzr0gja+sMEBWX
ZWkXl3oj5BzPNMgv3RYn63jFhO0hyh1XOJAVqRKbrULfRCO9aUCw/jVKptxht3iH
9yPbjvsvDk59grPOA6ftDTXecUzGCOA9tBsff9U8RD7dVgZP4tgy7QBfssatzPiv
wGBrKVxR/Xctxra/sEf01d+T3HbNy9wIgqOcHJRZGfBCWZu+02pSZ2i53kEjakmX
g92BK17b0jj7HALhs4VHm3fXeenhK4C3zEWCQTgj+tA3RhI1EDFuX5edqkJgwduq
nF+XqNwQ5UcPe4UAQJ/42FPLxamU/Y9KoYsFl6AwiZiSb2Q4hIOzshT6EHGvGHsn
FbFMZumLifhQjtuJZst5MWNvqnXkaq9olrym3G6T+Dp3fc+KSwDqDmg/jQFyI6Yf
fcYY8+rSOCQvUPyOERQhIJOAy3NJ9H/9ZWNARk54X+d3u1V4gQ1FDoM/zh+F/rA9
KwQRB11dXDXAzIUXk+ic/CW6oyBmApT+8iEcpFbKgEo64G+53D6hAwyF2ujK1gRL
s4tioZoEUTesBctuyXdv7UHjmI7rAP2E7xNtWzRshGSIZrS1PMsoKnjfYkxgbP2e
VMWFGYb75duEqnDmfHQecUPy8mtAz6u6l9ux2QCibBC/KvLpb/k5X0OqrAyEUriG
kdiwgsvctS8oal5RgoS4PfCcQlW0fwtz/rufcSLktlkqOUkL9xadPWxNp00JK+Gf
zESZd2y55louNSYpzE0kBU+Uu07bwO+ptk+ZT6FdBNLU4mgT3tv0nJWeyVd9yWGu
cDxCXLzQ8gpNDFkbTUHwNigHRoHZJlHr/5tIfUB9L4oRRrllu7USPmckOVoli3Da
i5YJkCHxQ2rH61zwQ21F9/SAUufshRYsvl8y7CU0hIQko68jDKRu8VpFVpHovgVS
CKqIy1xXSBWcUGuv+FpAUwuZaXE61V4AaObDDaqaMP2c0EQZrdfHd2bEL+H2YhN+
kwo0pGKvlbUlYVY37So6H4JVAP1+bmAoTSKPwKIjc5TP7g3NhItQc493VQWgVCwW
BK+/OJ26QDKrtAu1emxaHSYs0IRAbTpsZwrRSZUAKFbhJDtPH1uuimFSNtKMwr9s
CjRW9rwejAXF1WL8SQ0Dom28/MW3qCO5CmEdjSagdrSJKqFZMnDbf9aP7hXWy2OZ
ziYzPnLL2khADUC+pwLm9JB/MF6CoQo7iCH0d22NXgjFAVL1oqBwvfoDkDt/vWmW
peKRd7SdOjq1aWdfz2cAaGMVMtuDNtUr51wNRWTh7iowW0dXyPsL8m23N7Z03kU8
4K4SBlofCWU17fAco3B+53I7knv3wQ37Zqpccl8ICXrymR0hef9JuIkplL/YEh/w
dkVKHy0xu0iG0U2WHOZpBjU5SgkkFwKOYWa1o5b27AutqFnqv8OMTnoGgDxvJ9gV
rTMcF8vQlAVehT2lR3T/Jrr7VgAYSvetv661xByYj4Q9VzfhLIzWxtLTcHUCdW/b
S1KSgLuP2MXGigYrZ9W+A1edNvMeldcXnBNdwimDPUbeyXnvVJR9nhM1ameCB/t1
lNl7UeiG+PhQpmdSdtyIZf82Z6cDSuBZ9C/Ep/FT/urPfVGoiFUQqmqgEeoCsHJI
htFT/UR+lIY4lu7LdMNeF6TsWHzksAWbh/XAiG/G1Stco0MaE4zy3NcjeiYCV6Dr
rxMgA4yHT5B3uw9LEzwb3Htg8gOSea1IVi1iIgS+JpKf0l7tUY+kAQys+FI0Am2D
qINDW/wGoVhp4yrz10wXMsKRHGRckoSsKwMjzXOJ9KmGlGoNmjL049szpljrWec8
3PQDXzZr8v3kYHziB6rLwjXx+xttvN/YuckR1SiHtx/ZopSsVRNusIcwlrzRM6xJ
wTZQm7Y3SpqaWytOQA0GeOgo4JDPFDmFFkJSUA/phcuOIjkYXOJ5SmxSjLhSFAzL
quxnbAZIC8WROpWBfE+05SjumFcTZ2rZfvFuU0ia2gPMnyU+Kolb83xUWbr1V6zC
9/WdQ/uYdeYUzBShMn3nA7Q9MHDZv71R2mKjhX6MPDfJPJZPKUuo8Q27WYSPqRKm
57phv4q+mV/wzDjZNvw4Bm4EzP2rPZBGYrnjI3vcuzUWzXMw1wZwV9y1NXMLmhbE
F4ciZSaeWw6HvetwTG+l2gBIwjcfYWOHHvp6znTIEkBtZv9JgYCVgkPnOgsZdvEb
knoQULo2GCM/7Ffm6tbJ6Wq2oOvPODkvSKfmVBpIQKSZ8m026it3V2dp8bgvkpCT
Ln35wRjEz1kaSn/dyQwh4UCtkattQgfFlH9a9i9pXGROSkopBbP3JqEvtEVJ/iJx
LpXN5HXiVk8KoqocHqMo4lG+p08MfUZnnkSuGH0LxkJ+5uI8N8NVicq+gNG5Fh5l
+rLI7EKsiRRnt3GB90Qp5EUFXBNGpN7TKb++7vMzlqlu1NpZMyzlSZJZ0D2KNpG5
gREiBGpZhU58A6EKlriMV38u/4BZ2mOHps3O+Kvy9RPsiQN8IlksQcCL0qiSmiyT
z06bSg029xSSp4KtQgHXlGc9W15JZ7K5PakHDktfDaj/h7OUET1/2zoQfW0VSSBt
eQQOjSNDpygK0uDBUJ0XuXq8opy9c0T+IxyuTtXnThjXjCrGc1XYXdjregGTjhdO
R6Mp8kaZQu/qGJGqXdpZ/QYOGKZYd1O+JztNCpi33PyutpaDturI40jFKXDIUxl5
vrv8ozjag7/KAXmCAsU7wGXc90oR3dtSk5oGHzyOkQXNqnMdqoN/054ZVUfJgbF/
RGgvokLBL/epN7o9GoAL0mwHgeQU11AhjvXErk5+Zlt65ZdHLvJE6Wf0UHfGyjzf
maNTECvAOK8GNZT/SIzGQVPVKpenkwzdUKM0G1fh3lAncz6WS1evSGbvYv0LOoMc
GLB0gSFnr7fxPLZsowSb96iLAo0lUU+E2x4mdnNyjACb+tKzNt/vdLShoPp1Qqew
jEEiLD3qXE6B9An2+uYZwEACEvhPIqO62aTJoivojur0UDCjmZzmFSfkk0kjGiQu
m5PuJPjLDDBZ84DBla7Im7UcxspXjXUCL87N74wlHwNsNDxvjyt4jQbotHBJwnMo
JA+Kau19XkBkYA5rtWiMczOMuIapMtE8vsbkizqyjindAyJtZkcN7IEpW0BsR4nX
jshvu0Kj2psmNN2KCo4hUOUbooI/f61LgH9XFZqxN1vUpXuEPQXelC/JOUSeteAG
mxyH/pM1qjdjP6GKtznFvIRxk3Qj7CANpVjcffF9VkMrKLYC0+XmXl2dg7OGUipa
QIOOYFeouX7U3gwZHqMNb2gPM2xgmWx5/j6C8+iTiGV8+vV82FJwWvNSLGlSOUSv
hcw1HfCDAS5KzyIhGVkSqmsffYhSG/J3XyqMu9iKqHJPnuXl5K6Soc+8JJ9eAhSw
JOB99IIB8SYOZav0uMxrjqFQBCaZAiNbrAGfj2h0DB8omONsUX5gl1X2LYtglSVq
HMnkibdhwcZ6OBcpeDd7kIqxaS4Sz0vr+ubRE2Y/WvhyyGUgVjpf+dsK2fY5Yyov
W2hSnyIDsC/55R0pQAoxu7ggF2gXIhFRwR4ZuvPcitGm4+zYxgYC1b/Pg/NFjTnx
dY7ZngcX6cKvkCIippJbd/3AaUV6CeG/wTZVVHds8THlF4gAH6ri3j4XYw7A2uGy
ZGEiIBP4YoXG/Hf80cZr3w8S4X5PM5HgR7aUtayr+8ZxMIo3x+ElijWSL3fOamIB
eK23njMd/UMuRj9RMbwrMRYlqNUYqsHSVkK9IOs6oa3lGHu4NIjDERAVxcppYMM9
mTqGCMnxcSp2zpy7QgzibryUySjaF3N3RKRdGXjqCL5+BJJRGsNUTX9aRpg+ocVV
WvyETOtUN7qKlwsJleQTLnJRKRNRQG3dBkIfbqudWQGG2pjfTYqTE1x4/FK/Nh+X
/+EkEfX2XSqV7uveHKyiiSls8o3S9sXlq+1LQ3cKpEEpB/k9OQscCoKYmmau9qxl
Cm/wwIpPhZF/TCWlC7+giQtH0Ix/hK1lRdLQWJvOJiadzFWBYySyJh6BDqN2FBZv
n9ov4ExNGDS9MNHGg1pFeEsJfzWPKS+KTIPlcyDTwBYHH2MOOY2Xxn7EOV+S+Mq5
0/4GkZK4tQuHjd5WG0er8XlUgcOiJMxZLNcZd9VJZnLHwqREnW/v93BUvuNM/Mm5
B8WqZNddB4ksaHdvjKcvTU2RpVPgknpAgMbsYxzQcnji4dTtkJXXtAOpe29ACo98
rfz/GTc8pw7fkWXiPai0cncoUnKAW1SWEQG5jUDEt+tebNeGAj48mRg229drFzwG
URVRrtYhGHSTVY8WDtFI1kEkI+qf3AzO+/iNOatzduLJSCdbL8uFn0uEHrZBUXB1
uFeTzw3tKX09QYf+wsMiw2OeBB3v90f0MYzquhZDXZTcjGa4gfzpfQsgwWo0DrHW
Hvj62v0dSKDotH6kTafUArhs2cozbqiXtxra0V3oczvVADdFH10Yh7xuSZoSEODg
XotUtmlbw2aGpF5LniCIHGOQM3cb7o+hLqUGyG0ZgQBwRw02aN9imDgn+SImPeGm
TF1B1l5l3p2uK9DeN6e/J5Hb2+oLR5hbgkm5sf6wcV+9TytVHR2k8MHXsb8uyx9n
tqgqqfeXJCvjZXe20ztEaAEKalivDgdkW91HrdFESDQN8fq6p5LS+5XpRqlGV3xY
ym4ZaNESM1F6IjJSjL8KifdrlTSltLOwyGZQdpz+rGXqexmAUOHFgmrdTUOP6J3w
J8FQ/fmcC79mc4iszyegeHDWLYbunMMfnf61VGLOfbQmkv0dMLBicMQCF0QcyH6W
Z/s58qdFKepKgm21N5vJz3H4yHQHwtws5CYCSHRBlAYWgMOTfQHi4zZjm6/+EHMi
MWs9ZM4l4a1muvZCRxp9CgqItWJjaYfEZBdCXBoCcR9ypa5uFZheD42J8IxOwfW3
BGHmCI9l8f+RwFJdG5VkL6EO2RAVVwm99HgW/PebPxyEg+77X8UiN2iPJ9YMBba9
tQUjvJafBfG9VoZkjVIN5Vtze1gsXX6+4dmV0zjkRl/YFpdunPV6uR8U0k0FyJkr
tIyfJGzqDLJJ1XPoRlAQ0EUMlIF+FKbNq0Y9Y1rRw2D1EWhUrd6gbTySwkuHYtGD
cP3V0HOrp/qL9pdTb1fC9X4iliKEAB/7X56yrjHuQsKEjyspqtE6FMW0y3lwgFbU
PhAaxtKx3NMXfL2lbF/bmgiXAX1F6V2ujEPZBIQVFAEgYTYLUBsScd28VJjqcucO
GcZ+EwVzDmHkIxw9oOFA9uyaCnIG6mpMhu92Ka08f6ZmGNLv5laXvsCAQPd0ELU8
WSdKBxkJAWcC91B94ht2ssES2ovHGW8bck43roRqOE6lqJw8L5DsMRzbJcS1+9Z3
dAALLtdPNSlxCElqChV40pIo+Fp4CPDIJjjcaYKjS54B0yI78Qyjd0FukF8iyEBr
p3upoVH0hOO4qPMoE6tbSSRuSjsxu4QiunU3z7GKAyUnW4+rR4Tkpt/ezycMNmbM
/grIqrU/xjJ9fPZHhpjg74+3n2AAZyFBamXO5l1Off6nfkYAiU+vNNG4VmFY3DnL
fD4yk/KZhzC4TxzVEOeXFHk4t4sXKaIx02KpLnJcqaCts+a4XX114fqp9cB8seQQ
m+c7GGs0zuOpMw1fiS1G+JXHx/mgpIwI97jLUJN+ExTT1l4i9DJtsndr03kDO6hq
qeBGm30RMpJdlHRcVlQ3bi38h05IaKwclYlmESko2aOSjIXL6V+RRCfj2Ojymxep
x8DRVqWChl5sHSOv8y5lBrlObjYdELbQIdZqAZrMhUWPYGlqgaefbdedbfxEgNkc
dvTYBmuBCTxYfcQ3n3jq43CeuEwdoFYKuKVO3mt8hIMx0j6LpHcR36Yv1PxKg6BV
Ss3OC1PR5lVfliyPnUp9XzcTMYatpEvmpRxoOuQa5c7DVoZO4rWFdyKs5UksgIxa
jSAznK8xSNS02qSz3tv3E9LqJcmU8a69PIMoxwcA6WngAMv9cGlY7/N3Rx61NfDE
S57w81x4y34AviMscgQj13kmmQV8E353pIrhOd/eOWCIpXAi7o1X4SiUF6sQJXX1
ChUem3uroUQsB0rkYtzrgYBsVS+WiqYUx1vMGGeJABuwszkPikKSwu1HC718Luhp
JH8r7byGZ/1C3vLfwMosAwvEpa2xXQTKxcS8nQkwHX4HMx7zbIj2s1pjo51KNp9L
PfuokutaGslagGAA8LfsTdCD2aWUOrVhn5JwzRHiBQgl+ZBOgmlFaQpfS8wnmdJK
yiPaPUxDD4jlAHYYB5pJNbAetAhmOZgZGKIwyXpg6BV3hCLPTxoNuYTdByeRGo9v
FjpdeI3i52Kgx+PGy70lCIOtbbH8N2UCCP1khtoJxRYVGodWyhKHoKZ/BdVY8HyU
CGfKt4/wq28DAN/2cK38XWNZ2gFp4DU5S/MewjFxPY7xIlyeGzxrZ2vIQi3mKLoP
tZMT2QEfKLE/66H/QL/VxzlZzTRxMI4ev2y2s835GXe9cAQxQ+MgHDFB/st1gajv
aNBzDcuQ6I5Mi63b64u1uRj1YbXHtG0v0bVJAhKWiyXN8W3xtUlcGdyZXNF0Okm0
lTgNd5YZCXbIApMParaLrNIxkvdSixFXLLNiM/oyLoE54KOdzNux61N1q9E6P57e
wRUyLBEaqdQN1g7Q/xoVSPFS0Iqm6ZPJTv483V/mJbMP21OoPj+3KvyAKz4NfgVa
wj46nuuppUKcgMkigC7fCLY5aVuPAKf1lY7hUcBADWkXxtrG2glEZphydBAdtX/p
svmQlvxGzkw4//e+x3DxFkHF06X67wPv8+nDSJV9eCrK9bHIPt50/JMGLKCpSsgn
i6ahUDTXYL/XH9XSaB95Aocorad6VUt+XOpB0gjVvCPlCqM5+KPkYq4lTQVn+brt
ettjJ7t+0FuCPLCU38VUXH3gGRhl++LTNddNmsqKNVFOiU3F309SWrZ4X6PKmMEB
SPgyF4tAegAgBI1/FvhdS4E71kXeIhhX97MTS88H3JRlrsatPPXVGkQXdC8RPS9G
+5FmZCrzm2YOcupmECRbmmluAZPaQkVGM3Pw5QqyO5AFVMNqtgUYtCTU/+rR3U1U
7phA4hTDmMwwhElx+nKn9EZrW4t41LJY5mYQ7svdSoNxWgt/uSD0VQ18OIyuxe85
BanvwQNUySCMhe9BpzlBY+vQ3vGshcUA+9gz3it+W6mnmA8ZVdSLouKdFyQ6qIU6
A8Xe5G2tv9WuqDpP70cG9fhgELUPtPCClzyO8kztw/LhstntzdJ6M/kATO4PFRbF
8m8PDL4isvq4VK2z8fXcIFzfQ2jtgYXM3FO3H41XzomkOb7/BtgewE3cQqaNa5Ow
b/ZfZ6FSEBjUHJQeGYp51KDYr9WYZ0TySIdi7cQLdIYHZEWZvsoSerZAV1as5823
l79psDne1qY/R517N+rjJcsg6sl3AFVYwBwbe+D7thiaHQLpn8EVuyy6r1HkwBrV
FtjNKx6Jx7vlx+kQoOGD1OUmHm/syls7yoxVK6cpgBzc7TkQgMvpM+SV9/sccZCN
IyJy2/N3plBOafAsv6rD0nlDOzk8n8VckkWa4o5eMizEsq6gRiaxlLfTt7EChERh
6smdRR+M3H8KrLyk4xkIW4xbZTyth9e/xzmI0iWVoP7xJ8fRK6xxbunjtvNbj1gT
f3LTEJfrxI6B96S6l1ODBF4dCYRPL9ww5noKLgXFUqnEvhXX1DZF1ppvtJJSM/OF
f14lak/pd2qZNOgdvrkwi1P7vj6g6Ilz4R59/MlteaYPRQjM9FXnDEdwLF0HOxJF
DmsaCiDSOh4De4giUY2u+bDe95fS5+Bv5QzIXZtYHJVJMPT57z1DMKakLWOWWIBV
tKr9i5J4hUClNaXXY80i5WHPyj/zSLVYd3qDnYHf/MV84u6IistJImb4qW4G7xNj
+L3vrTXlEthbaSFLYN0prbh/GZVeRhi7IdJhragEx7ZBsqRU245hljIGmr8LJ5Ih
ROKbRb2dGoA+Y3ZC6mdyyUIoRk+xZivCut5AgT14yBOz0BDc0bdctD39UdmSkKh+
oIRuMy6RGsYqUwkshBz+jPR5BkpvUfDPyUGbmqaCSgjd+/0l/uAbTHqOvmbj1sht
hIFa1Zytom8l1jMXSuy2yGWfDRuQFP3XIWvTSNl+fzVpWFCNTUCNksUcf+o1yDrl
RYSbt5HFm2+zw5ClNPqOT//X+mdkxOBRwjMoTvJBGfbdF3Lm39WDZPJVl/65aS66
kUv7+P7jD047l25iDJku7mZ1ZNhu+w2/IPnpoKNVy4z54Aw63BN5XLWUkzgngUOv
tRUE3HtL+d0+57MlA/cDb8L7axlcnOghJT42HRBDU6NucEBWlogRhuYlll1NIEUU
CyYdURE9kEfkBt2JKNY7fh6wqT7/WcPihCaHRArpaeIAxSZYsH9GKTSrTt5v/NGs
uZ3mDu3j0GIHyoja+ebaM2MZEhPoForseAcsD2GqJGeB57pQH0XeB8C0ekmPCqvA
HCzl4Z1aYM0TiyBzTE4FFOA/YPJBbfdJypbp+97yjEu4vJGTDBI8FAwhrhobVyal
s5Qje5q1BPhRs60Cm5TJLQiBw22pyaBhs3En+Cc94tBTj/RgIl9LrraqN1UYGptP
+TYTrEp2aj4ju5GjPU24oPcUuS7SIT0Q2616a6FSoAS0eSZgLu3bZVskklgHRhNp
8wPkqHrBD/CMZ7TgSuRRILYEORcyyB04qKiRSOsevwo/JKYgNkm/Xj4wHe8eaOfV
2iQMeW/ltzzoYj3M9JJdnVNTNwBmUk337HarJmVtVM+tB3gw2biKGH8QR5mZQV1M
BlSjPrSWSb4b2ng2vYZKHqEAescWhqXem5tMLI4hziooLt6H+8IdY/CvXxtoL/18
gHw6KyHWHcXpJ4pqoHcDWkFryru3jagL8XhFJcfTVWRNJzgoyGAaA4DX1Vb0H5q9
CYpKnzUhCmT56QuavFg+u8KLT5K+V2HmtJssoys62nZrdT2/hISG3Nsr5fLZi9d6
eVC1djoHF810nszZjvaiNRjPq7C2gYui+Smxzhpuwvz6WvOTOG1saSg/qSBMd1SI
4GdIajyJVVBQq4osrT/192MNbkVLD3xMiu1GQ91pHfNY30H4rALgKUeb4ZOrpgoR
UHbbgaCoSJHMcKHR96Se0Arg9DBbzu6gWduiAnuemjE1v94HrXFU8qQ8QMy5w1uL
x8KTcEHyOL54qXRYWopqrb0NfHGYTTYLu+wgKoOSAy4gwDmGyAtxsU+KLOCLhLBx
JQshe0Mjddinzd0tcJVi/vvBt2X3o0zjWKjw1rKzEa5WPRPvx/1szGQziN5UKT4E
rdx7cVjpJojQiB3ZKyvcO4SSU4GYSie02imKHyMDZhSqI0L2jubSzUqU5a6OVCjk
pXY9IahJQHVQ/lM8e6x++lswPM0wozagsmehLMyGjU0c/sAsdHfYhIkK84ggfN3c
kbpxX1z9O8A1i078g1PPXUff+cnV7x0ccv0pSRaSBftLryrx2C8ZNfo1KTb34sUw
Q4kqwfhI5hubEHdFF0LOP+4NN7rWalDK7W+jxAR1FMB6NAPHVsxiuRGAq2RDzEFc
A175SfbbIWlXUzKS2pqf3rSYQAnNEb6N24F2nXOzA0sq9YZPMOjhKvdkyk/UCgV+
NdTSWHvuuqja71/akteAK4XtE2DLFapJ/8fDYcSkH3MlMctP3PgsWmR/I3Wi8oDo
DrmXFs3gRUbWTM1832gNUX2urptbPfMYmqEiC2iulxM4/hnd5B+du2PPG5OppiUz
dDZvORxW7IQKnKQHkeOTTyOIGvU54F+c0w+KYJSblaBrN1E7dENfl8T+BDkTvne6
Hd/oGSPv4u+4rMXYVig//cc2J+Dyr7GkDZwn9z9T3o6fctmX4GLvccfHPOt/y5gO
zatB2ISH/GoLuJUHAt5LAKNZ5dt+q8wM0iHoEtE1X79FYravyW66w5ZMLWujeC3f
P1wGuMfDpuTjI5TJi33KqrmfSLqhNe48BsqOBCMltpC6sPgN4c/Dg8ia2q6t7f7N
oUU4FwSiLavuFK2l8bcpBBJr1EEGcrV6QAOf2FlimefUqg5AAI43HWH+kG5Gx7M3
wiZVP3XYnETeL0L2oiu3/l1SJ2Zjrkdge6NSLa/9wEPUx+X2Qxi9s9J0B+sZhpCa
thmnc1fF+4rCjOFafBrXOO3pOc51e6CAHeJtixmT0gt8rpR1kHoBj04ZZP/xy3oT
f93EIoVAp/1PTtwBwsnIxuEFnhWYt0ADr8AGEGRdFAnjfwnGlPcZSdeE+YpCC0Qj
OBSmOPzS7FrO7RUuUb3pZzu0WV5kIIjRtJS8AVRHP2hb624jafgdxmj4NBhKEttB
J9Fl06WCHoG7LmyJzrPPB2F40Hkdz0g6fCa/oYPcKpC7GG3ZgX42wVsGHiPZLAFg
2OsuRGq80iSbqSMpqIPQPnN5xAwSlAzRzTkbbI25/5Y9jgKskvrAPQuA2MeIkmnl
0QCvYi27u7DMYpWYVmsQ0cUH1kJiF4jaYE/eHxM36DJ43yV1INsbyCQ7kGM+BBY7
o2qIocuJJqPdssemgR7ctuD/csIUI9xNHiMN+4PQOqrRrYuJ99yVTLpV2TiSw5vB
pOMKxi9DUL8suEr0knKtq25D10oMAsFyEQJOZc3mFA0QcUFWSfGKGdBl5SlZwrtv
ogyC2NEkKAZPnwWaNvqQNcUsF+Eebc2Gkprd8sAeGta4gQEvhCXdVCgGOtq+T60g
MI1YKpb9QOrkEAo/H1+x1BMlWvqeWP6V9WT3w9lAI3ePCT5lFnxAk45sY7Yjc3eY
4MECjIquOGQFdR8UoJQAMzeh1CEi/cCkS1w6RRewS+TfkqyPGJHAEuix4sjYx1BV
poNhQq0VJYu4MGkWH8z/dT+KU2Gri/jb0YBnip82WK2Ce0BvqJxNyXNZy2BvWsVx
uUfrHnDGgnBSeq8Am2w7ekojnwjzqoFeZX0s9Gv4w1EG5Pqnyem2eHmlPPDQ9GCL
aG72LvvN8DMjqHnzTFxMuuMPekQDzQeMcl8QfK6urvNcIKcNe40w5XtWA1UwqBIq
ZlBE89rCpzM7g3ycclTM6tQFqVgpZzk3GKEST1fKfwzPmfrpjYY8OStL2xI+3/0o
gMH33splIo9/GtRenBorFqqIhub1UUSLcl4+MHlv4q01RBNitR03+lsaVzGikWX6
A0UA6aFbeqQWLrf07qS0DfCZgaMFvbjLAItgqJWzNV+MZFcJilslxnBDuaFPxyN0
NtKeyzymbFHu6vJ8ZuhDruwnuPpQ+Y9pgpCczx+0ZGjy1VWWn24QNdaJ9sS7syfi
RPazJ9e7sSPRZHKfdZ3iDJJUeTVnVTRwQP1vXBBZm4PqbYPyejgrC510pnbT1wsY
5gMU8jHDVxQM/3LlDjJkp9KTsdMaj0v2mjExxCZj8ApLyMxjlj6dFcf1t4KYm8hQ
piyIf8kLKkdeOVR7OYbNCRr2/aYEUMsbZBnLp4cwhOPH/HNNNvToZDi2DBIGxFAp
4mn/LxtQZvnEvklTYFXCMOsW5f4C8iFyLlaK7v/D0B8h5i5Gnnx5k6aJlLxLgNEM
L4+t+FJeYwGNl1p/ENCcBCjmTDMdhL5UzeoTXSgQlQ+OOX7C/oknu6E+uqIXAoOe
/0HoRYpMBFidK8j4s2HuOsmkhiZP6VbQumIWIQhd0btPbRv/HMB/Lo+7A5DZ61eM
AHOfXkcLtbVL/LMb2dUIY/UOIMmgdewfujNVbDCjajir8hcVQfjucl8vqBZsp5nO
cWhpPH0sJ9LRVSJJbPiW7VEskN07H32G97h9go5gxU4cevqoq0/toFqeNcRnbZzC
9HUdwZ++eGwNIajsyCGfau0UD8aaR+cwTa4tcaKnMo5u3TwdbhxkuqavcoNlGgNu
TbV8482YKu0hHNtN/EIZ2as+OBNfROXRPbJ8fMkzhNmHzVt3J+bDMf9lVcQbhfZp
tSAFwgUY0Xlm7Za/JwIev3GBnvmyq8N7RM5BSfCWjs/P/nOXxbMVHB48QxVa1MUZ
mBBpP22zXFhfH1VH9xhIvHLa2xsZD10B9ZXOFSvOGueXn2Q5Fej92mrc+enl8Ink
hW7/y+lWsXr23IWPwFYKDYgNKIPfYzRr7XSGxJQo5qe6TJwSXb3IYhSi12LZOeAi
Loq56WwXBibKvxdcms56e9OWzt/fOAz12jsOY0N5FiUsGf2iyL5NLSWTsJyoJagJ
LeCWHVXRFgsqzOIIaAFU6bPDvOQu+32bXZAJoTBZSfoOnrEcB9/nouSE/RWqqdSn
lRcU9Zq+HHWembenf+SD41pegEQxJpUOYk01z2HS2wb2qXQCYzPEnpcEYBA0kiSb
jcrOLp6f2diAJeXDunRxDHgLPiiqwqzuMDb6F5C8ST7uymqURT3T2vijqWdznw7U
zTHyXGqxcJuVv8XySIDxTt521dfVDdKZOI+yXDWkUjhCXGPH/xByuReb9OEkQbtP
ol62syvPSStf+CgwCeNpBDJ6kKZwEzBoOkeO9J4LrtJcwWy0xLiZlzhEdHPL61aE
yAo7CRs1/2HTJmYW7o65hO21e2BJISoZN3NZuQTMhqwJq8Lur14o3e0Qo7HcJTTc
LDGZUmPX+9NzRfIJShIvabr14XC/Z1WZrJd1c2oCW8iaJ8yAcI/j9XWHJZYlv6gQ
XqE55uPoSwNDcK4/LXkxukLXwTGb+glDaxhs4jFM90fsvIrH3GCmxK6TTOLuP+xP
pB50h0ip+1bhx4nxlmDYv1sBF2wIaI4qtVkHBr1Df+UOokwePs11GZ6JEqSwNYO8
xdjaEy8lGOZ0rLKauhY5wjvhLuiDe9GWRQOpzjWo9LWH8fWO79RKPYHFd2cPKGEE
4uSXvfbUGwAHm5oorw80ZPzyulFfldT25S+4GjLD6OW1zmueALCm1EmGWOjK+RKt
0rcTUT0J3Oi/76KTfZLH03qcAZNevJOEp3aDkGN6gVfm2xBXgXJ8C1O3/nhiDkW5
A19axeh3zkVqwW6TUtkHihh71GJmQ/HJST5J/fMovDPLz3BP5mQlkYMaFK5lYI2A
yMs+hM2w9S3JpvloliVJWZ1wF2vjljCb8w8+oy49zR9PbiPGkn7fBkSjOrqGpmE3
ej5EZ+tJPDVVtz0zTvh3W2M1TJ/pYb0EbcMECl3hLTxXg9NkEJ/VLRVWYZMOcMFl
XYoXjwpOSjLdB9nIPNyro9Hgn5RL/81PRP9j0hv7oBnK2Gd75VSKDMa4+lCkXZwj
hhsOpWxaXHwbI9NJgkJ//EmI6SOOfcA+TcHkvEeKz95T9XT5/EORVGl5DLNbzbZ2
LXD8XFKYzqbufmDXCohHewhaa78pj2SW+mI0AaPR1VJ3h6EULU3oojb9iA5Fqymy
t/CBKHp1h8FKYo1/BHh7YrU4Ug1rrsAtp9WuOzwMUFr36fWcFYoZpmN/2m61I9IE
SVYvi+ze6U9vesGgWekjXLxzUHQyT5cwZeeigyDFZaxJqM+oeUkJ0AZBIjeQ6ha7
1Xwr77YxxM6KrfxYq7ACZ5VZdMLBPAvISteSGfYpW2MO4hdJD+tPYcBIzexEKkQ6
cbZ3wWBBILM4y42zwNiw3NuZuuy3iZFAKf+iykzHJMki5qyIB9FodIiOx708Rnx8
lRbAL7Itg7fhsqbqiQEZ09SgEEjdx6bhnw9hxc3L0wi+SG0SzwnB3tDoyJEgjU30
P2gMZIaOeJS0AnomQZrwYlLu0MCzr+SSk6eB5bgOSgkxAw/W8zFpKjTNshsIgThX
8d4dkyYdldLshG/tB8SCqaMzR+fj30TGa7c6a3EJeySIOcK/dxHGyzf6jS2oh20H
uMqCo7VvKyzipYQGa49EEVeu0srT9B8sFkgrgfgSFOH4EpMlJp5TVXj5Eexf96LW
13gqtlqA+M9Pc42BT0nmEGNgm1TprL2UMCe+34DCc/wz5YBfwHLWVdcdgrnv+qOX
54yCg92vhLSzq8F6iKmAWw24+tLOh1ncT+5RyXcxkosk32RKF+s1Hk5epxllmkef
rxttgdcHs5YDj3iAr+9AnCizn6ANp3vfgKS5/11js+D03EPT5y2vR8uZ9prNTTlm
Lp6rxo7wyOZTJpV7/3Zsxs0M4xoToBvVuvKQavDl82MGY0RZPUCmnu+Aq1RFnu+F
YXCUr7WvfDt4F3GjzMijJ0JFYOsIWh1Lk7c6v5QC9hPSkr8O3Q6H/rkvIR54GTUU
QvPvQw/s25I1iqN/BYIaz//nNz5yyyvxivM9vRjmrZjuI4VsLMZLGC0CvWOVm4GS
IcCoIC3JmqZgirs9Bp2qLai+hBUT5KEEF00FLw02wzbZN2NatbzUNRYnwe/NGXD8
NDXp+FVaTrCancCwVnhq3OO23bf8jpAVXt/knMWK94zg0N3+8ieueocF1l8vmPSz
+OzOzESyK7Xdje2di+ohLUz0vYJABAjQ4ftopoMXTRbqGQ9f0TN5SfnhXeYKzevO
WgTKGpLS8vDLgTVNQEdHBJrzWDY6gN+kQLowJdy56wzwBB1/Kcmq7cvarOEJSsEl
9hBdQr9IqYtWfPkI0U0dWzrH00eCFXkpjmBWnSJrjBwZ8LakPl4SNkFUB54jCJmv
czMAwRUyNuoHbJsIihzJ7Iz1AjygE5Xbe53gtHCbsTiwqNpcn1jKCISVG7shJSzq
elDwhMO8H2IG+P1KyqW2FTloQGW03fRlHvmlXfkX8sqI8ALG3SxMyigvCZHiiXNu
NN/z8XHFN4fF+X4Ot4/Dw6hB7CIyjacvFgJCSo68j3JeDlEwjEzIB0xD+yEDF1L6
uZjUQtPCyrEVx3CyWBNLF8p6EuMQ8+bZ1cwBNIgJ3e1LRBDXuk16AdUU0mzIYp79
WEWlEf133XsuZ6jSRnDhbfeM+2pKHg8BsM9PGDMZI6elhyo+99s4kJvISebxA1VQ
DdG3y9TjmB6tFq7p+INvK+FHcxzbneDNmLUoqnro10ibsQqVISkVXBrNggqs5RHh
jteTUAoNYcjRNmtacRXQelBQUvDZMedJ2TpOwC6oEVkH+6GAS/z8iTJtmDUyDR8H
qgHzSmGCNITeqO7cp4r2SVQXf4akMVdBFYeyZ2rkNaIjKOT25A3z200zYPan73W2
Azlehi8eXFKwkkreTSYKzTFZeJ+iV4oY8HCJQaMSPLtG1+q3bYeMnPFhu1tHFBlO
9CUSjwCvagNMlFwnC5PtdsJUmC8W9awlP7UNCt75luZfaqwvqGqviwt5dIPP575l
NyUEPwwi0DuECgqgUOQbU6W7Rtzt6eyrLw4+yMyYKdcB4seBNyetDVX39t0VrOdC
zs0Dh400WcQcbiTNWLgOn/kAhTYE48+gCRP6EGuRXbcCtNBV4Y2Nyc/FSzpPraHq
5qqdHY7diKQqZmCpzB9bWVQ8f8AaIqlTzF2A2xlGShRNQkZvhiF3Kq9VcVdv6Dw4
RQ1m+BgpQ53J2j/EuiENWBfFWtBzh8HkdeSeGOTUOLWuEIxnHC8WTiE59hE2RqwO
wAXyM30iK3zDa41RPlr5Gp44IWRtIZtriVkAs/pmG/SCVACwjt8lKTSx72RhCWUC
Odv+SgVrnyo4E1mnHa99UsfRMJiwThThbbnZ84NI0XO11r46Jsci8KKwEnJMq859
rp+CpbyawQhuXPN62Y53Nj19PXdwh3uFnv4CAbnk4ldB9bJjFn+Z8o9rUyyj0h1c
IRvMaQRPS47vAXU29EXcJtagfA5D3pHmaJnfBjDC2i4BDn3Z5bwRBlYCtkjbLvSm
G6hhohm3fdGrCn0iUtMSeruMKyYLqTNB/KHP/V5HhicOoKuJdPrjox0yR81HQO1W
U+jv0zLegkv/yYsJqrk4FrwWZDThRBDoeqvklRkY0NZbPpxi5Y/N6CdS7xuMWspt
D02mYfK9tcua95hryzhywQD2NEyIIg5xWloLousVZISrh+XtNTBH/f8I3ylMGnNr
Zxw0IRfOPn8suRO8+gyTm6MpOpWLRUrcGP+7swzNJMJBJK0UNuBmvtbaY5sAr4AM
jWQxu2Fvna/VwAN8ss70ly3o1vpnnhIejGVaZ8p6B1Q9Hp1TiSze8b5QOlXE904X
36l7WopApJRbMaA3Zy+eaENeWiT2IejuFzVP9htUsJVSdzur2cSK8FVu2dv5R59+
Z3obqbUTvLBzHC1C6biztQtcqePdi3daGRuGvrDTa4eSD+tjWy/OpSgIj2U59xVw
jLirFF0FmyMuk2FTQzlk2YjQmj8uS/XiJyNX6ClzNvIjpOVhl/FvK1Pu5hsGPCJY
7AZKBCma6gXuoAUCRl+zDJN4w4355WJK/k6MEoVOHEYI1diCck+gnAoEkJCx9kFA
QNi56mmgUDLbZtnAGi38Aqxmf8nOGIYytJnHWEb3wDrzHPQTAkxbM+O0QjH1pvKq
koyUVziKK5qc3miwwLtx3Eaqpdm2KFxau84AdJy5gwllW09hucg91AndNbWyp+St
P3C5RKo/KvXemQfcH/qPsuZ7m+4oU9bgR7zjuohtCl/9QdnABZCFHqgShZUlualy
EPVBp0FCndVj10JIYZzr6SJQ6rgGC732qmEoggPaSTmwr76BerIL3Nz8vmbd7vrz
TnNRPNDMre/971oh28Rw3r9XxONC35wYUKf8Q1/k2ACJZOnaK/HJPZjQtFlhVp/x
mugbeQJ8DN78WC++NsaFqdfqctN/xvAHmXIYFMOWe7pD5DlTKrXAw87Um6XKKi51
Fbo/PO8qlAcQA8rqPRvdynk2qjzmzL+0DpJY0BllUdZZzB7YiZCZTzzga/vgvZH0
Xe0UT4bUeQminE69y5BTWlkmxzOy/n1CFJAQwwgYhKQGIwKPvxEe47/IhbddQwyf
5EiFytFvpcAYz85Rryl8Xcu74clbAAeXuOXGdphc8top3KZgKFlSOcAISXUgidiN
Xc5uu1nf4snLDzgf0+qAasO95JmKzMsqsHiLwjiMI/c6XfUa89bYn9wZFjPgOcWY
8weqH80eoh1FVuAW+KB2USeYMJieQvJgzZbxnxf1XUpD1vfwCWOg/cTqVLKHBjHN
igONBcolZHU6vwDQI7WMKT3seig0EbfTlvGcJ72NK4IjSAvFZo3/AT//fRDb0mMW
yN2I5f4XrsCK3nk9xLsQB4sw54zbH35lSbfdS7PnnojyQhnEl3Yyx6qkeK8ChFfg
8D+gMWf/+5WwpOiOrWS+IwnvE0t59Zyzaf5CRrG5zFiIqeJXvPXHlG0XcEec6W+o
HPpxP/1ss3z/tvHhPPjKRCW/e3d3iAOYYmBgdZ186fd8qAFc2MDe4LFkHsbneDK1
hSSOFYBERtmnojrZSAr9C7CkdIO9KKOK8nhox1QD9yva6oL/uBQ+c0CLkoR844iE
xYoXR6hB5SSU25MM9AhN3L2kchnC9lt1H9rgyyOvH6kiByDwDKxOGNclgYRBfemy
QTxEAN2PK1N5dznLaOfLN6rXQdqtWX0b9xCIpFwaldxrTJiV4hsY5hwW+UT2yvZt
esnnhqzmBLAlGZ4xsFJ7EUp9x0JVSud89xowYnwq/OZsrDPCTNrM8mCi0ZB7OCnE
Xd4RSZf8OkGf7WQcZLtBODjWrGGrltQKmr85bnF0aAbTPCCmnftBjO4avwGMvnH3
WrFCrsxq+Ss4/yxDSSDGKLea3YyX7PHR0nrslWJYAWBsxYVE9fLC9e2LjRtHomSZ
twYjwX1sQ04K+djlzgoT8wIqm0aeCsa9BM6JzrjEeYjAhNFb5hE4fmAft3+ZCfpy
4e3l/uNaj07k8fHiM5M7lN+rKxDMBnIWZ+NtyUquG4eGjRaWpqhBHZkmsNFMsnye
fGjuknie+KuYJOI7bfoJl3QOFniMK08SljLyJIyOQ3of30h3k9aFL19oSksdfhSB
eBGkAj4MPKZ1qG/JmuOvTnqPFFZrGUU9O0NwXW1xdk+nbRnNiSxjwFx1ksZPoqvG
Hrjrz0jSHoFkE5CGYyM6qUmluNCp1rbgkH9uWlGa/VUSai0d/HyfQ4ZcwDz4dAhN
ePyoT0AK8kqZtRhyilYzl5hn9Jwqx713ZQnZ2CB5Bp+wI4QfU6/D92Ohy3+lEGHq
Z3c0uc8RyzkBS7QlDZLr/r3rF/2E6qKUwjN5sepMEQIYNyEc7Ea11ES/VrKajMoB
BZJY7Ho/rZQ22kGipekX9XWy2d7T+6/KVOxMURvyuaaAwTW/awSuLc63xjInLrS9
gBU+22p7Cfg1kQWRsQhiyAZ5Fwt1u7nWIOsic1CmU5OWJq42fj8nhT22RoE0BPcC
3wVlUvoDP5vCMrloeeY7v1L7ljY9dPIuHZFynhaP5s4EwEbI1gS/OE26DSOMKbk7
yxR4c0Kn1sunLHLvQDFSynl0FPFiogwrT6N32uhhj3R+Ls0WcD6fw2CB607Wtk1o
3tWyayB24yLXrcT1o2dukFZy/Z96kCI5Su/OhnOn8qBA8Hci3gebXrm86XHlh9j6
4pfzPMXu9Dmb5A+1wXHOPqnPUF/gK9NIRAzih+ZcUZuJU6isWWUpFocoCXH7J9Lu
ZJkaZ6T84rzwhijW6FTdBJydQiFKDL8AQYfjNn2e6AywligduzqfPa9ro3PvrryQ
B1uAE1yV+k8+F3RInuXPSQ64pCDycYaLqh51Eq1bXSZsI6wjaI3SHaFnASIFb46k
W3dYmimldib/xmAr5htMqeKdV4SD3NyBHenW6UNzzLTnfI68zOZZEoPixHDXYWGO
WZs6c/wsQO06Hfxn95h7/Ek1uWSrjRhGNk6paY3awLWK7mterRQI8O5MDeeL+vIf
Yo5VSC3/Mcy3MVfUwT1h6TVUMxtBf5Ht9nIbI1uy1bA15etYT/4MqTZGlAc5hKpN
llAhhMVhiWNkB4xrO+CAUTeWtdPifIoJ6ZxEXCbKuBT/wKQiybGkRaTxmiP40qls
I/zKPUmwSlgF1CtFe9I7BcjpDGeDA5U0NSCybAvqG1SoHhhR5tCbBRVsF+CS1l1u
rQXJtalZgmO/L7JlDW2CKFuefcvOLqUFVriL24QQv0C2j5OBLVngINdbp8oN7Qa2
pP8BFFK+qa89T77TKOOL29SNWzL118vNuReOIsemQUCH6mvq06b2s6Hm4TWA/pBQ
7qrnysP2KI293NOFGPXtj52uqvRS+Itr/FTPjfcWeDcRBIbVbzIKqgUm9fzRk4s3
xBpMMPqTzwwte2RXUei4WAynAffkeOVYo/SNPr9CGWSLnbnznGsTHhuOkmbAFJbJ
bmjKqAzH8H2859dyXW3cynbIZlCB4kVsOfNBmpP8VQxejRt98vc2IvR0PTAWPkkc
eDdcBy69t01h26KjQDYrBzsy9KH2EnlmqZr2DFepnrX5x8MzTGzFCJkM59hq2tHI
2R5ro50oRmZwtD8CMdEsh++PeMp/hxybvwyucSf1Unm8f0qy/OO7TIqhm17wMSn+
22sRtRHyoqpEmpzOPBRS3OFduI0aZypQGYfMvMp1MkS0tjukHVif1k2meS4eSSZR
u7RC83isLslD99F6niWzZWTWlnbtZf6Do2aWRsE3tIUvqReIYIqEwQSVzNJVd/Ek
NJQ4WO6oYVIuHIdoP1ofSLiMLmJbWzqVPdP4SYjlFXRs5uVbz01A7KGPx1yGCHp3
2yMd4D1XgIBfRL8xyBIYd7C4jnnGDHRwTsTY4XS10MaZF0oUoqA8JqYr3dOz0fZ0
t81/Aw9BLWZ8ut44IRigUuqLsHrdqOGaWPr3Azt7ccgBU87Ar7Bs2rUoKeFssw60
JucH7OnnT0TGMTkHwBfgwTcJNLsHkaarNha3eojC7El3o23BwNFrq5qYnNciXnli
Ivg7Zo/Aw9/pEAl9P+HwoCBQDvJV73yKP5dQGa33zXX35/qicfEQ3oC9vX/m3TPo
trioMLbiItDz+sqSwtfIHetEHVOf2A+VBdrpv+8pfiF/i+9Zz+Jrs5O/knxY2w1W
oEXAUyK9vrUNf/5kIVijkj92QZacgswXFt2TbIctVR3ZzrfGtyBHrDv9QekzcL+T
nB1Z6wD+p7GPjNrmEJ6DSB8OPgaw5zNWuwDZCeO2tX9uWceHfPXfwmL/sMdPbDpL
8iv+pCzYJDp1T6qO7iIszrJDR71dghPLEMXegGckMn4kzIBntc9G9/WTxn95uY/T
GVxUHPFC3y7GrwDb57yOVDuCgxU671iFI0oa3ioImfOXz5y52Mlxf743/UuqCkyX
wXYXXjNbP7RiGlqNzpBw8jlVYs3WdtIaSEqxO0i2aPAGKfTKt/PxiKlKaDncwaGJ
GWc73F65aJuKFc4UVCoQo1r58Gh6HH36ldj6/gH8HySaQEQwlh5x2+J9x0vH5R0n
FrUMs/cD43MmuCmP4q6doMwUkEua34nmRt3akpAzYlsPeWXm12QOhNbtcr8e6MEG
XHPZKK3RwSVRtGPzRHj606sLH/lM5AIuCagUDm9iJ5+ClKcE334LF4KcLFbr+ch5
ZiK0j4EawaBF8SH5X4C9DSGjxUVrtn80W2zap+XY8hbvtYx36R/spIvfYxrUf19s
S0uZyc/svNnxGlMNBsPO10+DcD7QkUKTrlzS4WW4TJJGU/Tm7OPbA8HdxfWQaDgS
Igyx+vImDI27BR0rTIyYfIXiNc/BVUnigGHJouRZ3QBR6/if53gZIIlAdrm5/QYj
MHybXlKFvd417iXk9U8KXYyqCujSmiFYbeDtPK8JL/THM0K7lPWHjyMUC8UMbccA
yfSK9aca/m3wN1Qls+lmM21sAC7cd83YKca9cYbgUsjg+89S61aw4dmEry7jI031
ZRc5igoA+hjam9aW58QBfmDudgL+GZyXGyTzoxpR3Q9IZ36Ytv3EJtTXm6iGDueQ
aEoq8ymkXg1JJ43ZLcozJquqVddSSDlzTrGMeEvB70RRXlKD9hypq9dUvlpasUbZ
lc7MItONgtSZU+yo1ZlHMx1ipD5fNa3XxMWPYgWOrLBjjRnQGZ/ShowxFUxJSNpK
cjIIjM8m1eCQ0c8Ha/lEmWUB4epvNySjdJAr/EVFCw2pQsEU4YdnhG4oggcjeRxg
Sl2dZ+qqSVNNrKQSxuWpwhepkZHgFIEXvueeLLQLdPcrhbUwatYwHaqTNEc4VgH/
6B0qqW3Oe32Z7Kv72KozbtIqvq3xATT0NagcFBo3eZDCqgrF4+FKMAsadmPkSzfQ
/BUlz+t1YodyDUHdrdrspuF2YJnQHKXR/PKiH+wW+6fXncwL9SsEGP4USia89tAf
Y7zQv28vG8I8mmA59SQUaMIFjTAZU4aL26S2ljO4lcCVZWp1nwhLGVaJ1BKSl97r
00aITu46ITqtAgp/ugsHcEOsR6VRZ9ru7BWEUU34vjFzOENo8BhIJmXLcUckYbz2
O5h8XdjaxSZ7r/Rm5FgRIUN18GHfcnZWHbHDvh8svlLh6/QU0KfBMmc2fLyDRYAC
9SyoTbNOvMNWQdiv76LOhi6q+NZ0Ph4julTdgl9jo29sAL/L6gifptQdtCizWPlx
+bR7rdPl8zwHxIxT1JVDnF7NUElASUHMKilcYooBRdKUP/bqlmlLBXU5C8cqCH26
+DFVSoDMmwNHCjPhTDBmgPjTXat0FSEp9ukRzxONOFzemGXdj3MWtvJvBkF88XM+
RF0zFmwzWbzpbn5FrT/+RLTyXggaFZ+ZY+Fifpyaoc+SxpGIofDlkRfrxEzDVCGY
KUZ+Z7ulVkNCjEpdwnA4A746t6V1u4GjE5kUQNBVldG+9BG7gy4+q/RC3JS9jR/I
fRWW6TrqucuAAZXoRn1M9djfI+aba5tsCDvmenvJsIH20MXA1iI3oaoGAbwEEScc
rpcQ+NdyPOauY4Jjwnm1FuvdmR7lKBdfEa7j4RWL9pNWgbf/1JXYhLasxRF9u+Rd
Q5I7ZANR4/OonuvkDhrIWznlgCI4Doug+GmDpECb//eLD9goxPijP7TIIO/oIkv9
v4pn/5iC9nbsDESWXgcmqrX1FwMpbAUbJD+NoxRfyWzh9ZytvnKGGvNOOdrNNziO
7Hossmg0cvf1vlqhaZYJ5taPIrNSCzbYas3XUSmoRPvDs+dK4euvF0T4YzLz9yCQ
uncDctpsLcBcvPu2F0SiVKTWuJbIsglocfclTEH4j0vbnQKb5c/fgsNybxCYVpb2
gwl45VM7S2RY5Yf7mzbxsuy0oiQWyy1lrnHUtUwyqMxJVKw6oJOjkVD8YbF/WZWC
tQbjmN5G8dGy1SdAu3gcXHt7iqBACrN1fc2SjfQ+NTi0DXO1a2MDH8c6L6M0tRNe
Mz2mIN+R1RyTfF+IKwWy2eyBPb6EPnQs4AQrURwHm0jx587pWNByQYCdwSKRs1rc
2scN2LwQVJVCnfbkH70Cfdn+fB35wW5xqDArB5ifN1WNQU5C0nYoodhsSGlPp7X5
Y/t48YYdqpdxQ+3HvhE7tJnmDelPGV32j67pyqgd+PiWW6o0cssyZPUaNTj8lZHO
m50JdKWWjmGfPQjFlG0f9q2ilXF3oDXqYU2hA8qQ33t8YiEvwewkxp+jHI6DXwlZ
eBX9z17DeZJYrE+q9aMHCYmo9dHH6IXRo+Z3WCLB5miH0UAl0YApyWRure8YbMdN
/LMasx2uMEBJo3Ado+gAuloLJZmS0JcEGFBT47Pr/xmnOPdzexYH3hIaklMFGxCT
JjzN3/O7hFsdWaQDQAXyoguDSkRo7RQXM+SX2MKIs3tMxyxvVc2W0mrMBwqppkvB
qDaW7nETA79QVUm257heetSHP48JvHpV+BuYdPM76ZpntmUQ39qlR9sde6zNTc+N
Qwt8RZhPw5f+VvR4JFyJC3Q4A4CCW89bnH6szKY6+hDTUgef2ZKaCgI4/McP7NaX
AW3mNsIWLo4QwtENzaimczyFL8K0+1Gmkj9ExzV41RkynmsGowVak0fyO5NIoZQC
+y5Ik2KWWX+cHC7KTejpfeEZ+jWsvWgM83bp89vKIyc3dHKL+hiDeq5tKeGu1Dim
N4YEEcufnYPGgQxYqVqZ0ALuxFig27hqXG017M01P0BV9U/p9GbXID3GdRw1fnf9
3FRaS8tVu5f4z/n8O3cuWXuQA3MtLHVk02lSBvScVBJ0Vj9sAxygyVGJ3yPVLL99
AEt7ZJdHj1HKVA0DOVL6R1jXoZBRmlHrzVdnqI0a/MiPT05+wQHDFbuLn0Qf77tj
zP0o50of2V51oBwjfgYzTIWkt4vjBJGe1S+b2oZJ+Tec1Jj7dqil8nIC8SRl7E/p
/KIidCp8T8t92zWxMd2+xZrwdg/iSWF30FMB/DGJ/UuqSw1Iy1iKcYDtnnZP7sRy
M3Pf3j7pcvuSvQX/toguAoVDtUhweIgBML7/lI8qauuH2Q7MTi8M7QnYhTFsX6RN
ymF+ORRUdTfIJe/gPt+U4xWhR74c83HXO6uW5eqDwarUGblmSBdRkmL5RaDMtTIp
+KbkgXAUXyXjFhRRg144csdWOLBExzD5d9l0c7Z6J8mk9cZQN3Z5FUUEmvTEgoGh
wrNgr3I6Aiz8Ce7lcj8ifULxO15L7sXxdnyCOuyQp4AEVszcEPweTgfaNVFXaGOS
XuzsS1eMaRB2jC0Egmc4kPadPR+6WvcGv/rz1ZAG5eL3ITJ0v9qUXGOKsh3sd1ZM
JyEhTaHGndVuxGwWWePf/pmMFtzV/XUOn9KVTDDjwgQrcdFV9CZG7YeIddPenJNo
e654XCQcrytsVRm3xJK2VnSKE5S6d3fmr+cl0Q74rI+JCBdgxo3wIk+fdZVdQckE
2EFCPe3s4WWQ6gFgQ2dHB8z1SoIOh4ojdjr5HeEXPa6wtb90bkIoysP4YLHu9neW
y0fcJQtA02wKwgxPfVLBx0gb8Y1E/MFYY+H5OCF/m2zq9nPxi6bWmA0HfF3/Ib5q
pBe/47y6gCqJUjJ6ggUK8bzvQRNy/ZOAezW3TMhqHdj75Sov+n5FA6RyebNOpEBp
ws7Ao5IGKfo3/GjNC8HJKMDlUqqHV9EBrULQ7EtazEeweoi71CsNtrB9+nwf0FRE
YHXVFVGTv2rZ+7WCA04kGx51p97YPF4B1WZ+3EViHSaehtA/1WsdHbEiERd3uoOJ
hnhk2z9YfO+6VeI7BAD/+Qe9nNcPylyxnMLr8b354xKjRut/RDGn2O6/L6WOJ7N5
G9X3Tnnj2+MNkn1yUERC9tFm8pJenDiHhr1eRcCwUfAdExMhC4IbBDSUpvSQxzva
mAs8KkGfXEwSDR6gw4u1TrzdRj1iIvFH/4I+Rd57D69zjDFQbAloMGhn8wrrcJ3d
cHe6TidOpqCpzfQfxLK/LAYVR35xK9GcvvoSd1PuGYz6/L8czt2HmP4HQPbnOsHy
F+v0pZp8aSJTEX47zr7BRo79xAIg1/Oukulzzpn7K2fAIwXLKSDbom9rdCV+5stK
kHl66tplUfDQUoJrCfsjx0ns+HPQW0y7JeGcQJr43wwdcgJCw5XOPAd0EjTfwmRk
87R3ZHmIAG67o2nCmUrxm8v+pxDZNuKl0g7NdLeZ2btwIA/fxunN8WftG44tl4zj
vz71pGRpA91boqKrIFX5hs46lZAjsTnBXMldxHoOosbM9PnJpKAqL/xrZ0JW/V84
Y1XdPwpdV/jJslQdcaKdS8gzx8hzGdbxNv677hqNeQb2phw9MyQO90cDTpWhBoyn
CJCge3LJTSt6+naYtXinmahrL7UEHwRheyW10BDXVvTHsJj6ZPRkbsZvmav2s+6P
NcbtXboK3jQqja8TMkzQPR8InEmPkGyg//ncOa3zihRT6BNgt1A8YN8qdHl28CuW
rEqebDM042xTpdnypYa6YWxHwFsDnu2nnlKHunRVRcVSf+Xb161bI6nBA1lrpwGv
jL86hZ4mHQvVlVPX+oTCbXT95189bhtIf8qsd3kpX0KtkFK7rEZzozPbNzYvYBCl
u61tWG1QoSvCNRgD6tlpl6zdyIAnmfGalaSwlD0c1D/ROs9o32DqriTmFW8UJj7P
ng5KJM/VY5meIVYPHEnBI+531dRTCmMPsyLkQnzAUjvHbH8JowtlMd+PK6vAii3h
BgWCKuSMU2jI/CbW95Nxh/iLABT1HGV1qY/HdnBsydYFp6Ms0poKKWU2XNiUmWYa
epqRtrnmtJqO6fAOX1SUP+gw/EAoMBdS5Z1N6oBjNKYLbU3tmpIAT7MOa/Q3FVxx
0spZiFNXyoDC4qfc+At5drJ5wuOpMJqneZ3QRnLBcHcTgYa6sI6Qo9ga1z2M3Iow
kTix6lmqMXnIqofsaUFyWXuYFiptFRrJ7piVd0jVc/dW9+HMPbPSsPzSMY9+DtQo
KqVY8Cwyh83V4SAMCu3GSqxoJ9GeqHyiAnO9cgQjcsZzozKRYNq0YE5X6d4FNEzv
MazvsHK3/wjLY4z5YT0oGrUtiJZjTb1LLVTg/ZebyJtIiFH0eM97pHxN7ldccnxd
k+OFTxsf+hK8Nzk/iMPelYY0gQGQ2Z5DeXx5i/cwCRLU6Ao7AyZlBd1h/kza9zj1
KK4sWydgaw0BCu9QDGdCy9F253AC8e8MZcxcwOBQyiQljTN+Nsw0eDxg50SITWhN
d/CIuFPYgsHNFL2WoxdgMzkc5UrPw0ZH7p08FZKMi89K0CU9p+VjQv5coha0/C71
0ccFJ20Fqa5NV+DvYgv/oGPJzqo+BDCznd2NlWIR2MI4CxmUznwKKNTc7A3Hj/Jf
JWyBInrv7aqFu8Y7E3a5bK7vOPJjY5uLg9P9Pm0CBkfs9YCVp1Da6KANMb7T5jt2
6jzyLKZjHfhmIiLT6LeCgJvEaKxjXe/K056DOv5ZHzHtGx/poxydvZkF4C6FTkpB
DHNDTUd7fleiUUKF3NeMDlZKY/hyFt7D/t139NjFX66BrofzlQPHXjBTim/Za4/m
rSnlNsU+RugmmiSC6xgzS/WA7N8Ox9eS8OdeFg/YisTMAFniPz0iXGt/u09iDutH
WBctk5wb0R0OjFbxrm/gT1u9An1/WcomZBwH1zKqaet3ME45REDFtb1o7+URa04t
vv1ioBjOyeyUV9yX01kjig5EUWQzzGhesxx4zswCC7DzvHwVUsG+++pQBtcNl798
cje8QQmeTJdiHbh6rUwPu5+WFK1Sdx69t7CUQEulyaUw6495T3pdQuz8nqgvj7g/
IihXQPv2nHWo1gggEMHK1jIxo+sED26kebx0wJFGq4EIuf+6qHEJ1JOj5t5EYg+y
CsaelMayJ8lwWl/UE3nihPpk7mSLQQVZLs0trO2UjhX9nGunOKBlvNuuwOBnBGZX
zfEWQ9WZoIiq2x+aHZ4SjkfRCgH2Ld8heTq5C5D3ULN4zcH5AdAAnFo+qanWcrcQ
lKBGbVQspex5rBAMprgmmQTihIBzHYzi0oRw5Ob/wG6pfiV3wKto0pk1DAwT9djA
PUkHqFyGBCwsGRkfLhlbOy1w/HDMHXDdBXhvUdtRTvPbTziYR0HvPEmzUWXnLy0e
/UexUk3PVi5jue2muCyu4zoeRBeZz2TrRYt4K40KTSfLvx+GgbV4H+u+66UdNk/+
G0tTO5f2CktY+BbYmS6sugU4kABvdmfvU8qVTSDJSB4ypgjJsch8v0N3UPd3uAvm
H2DYF6Egm0GA8zLnHiznH5hxZq8oPI//2LR+pQ1hhFbQJrv/1MJA205ZRWdBNdMe
0gYSM7+vGFghsUAuKqJpFZMgN9UrfWQdyaY7ShS59vibNbWWAJI5CmjV3ZBnwhxK
HWNuJq+qWHvlXfqLPJfZpmGAVohmJejvh6NZaJI7vlD4IzOBv61UmSDTf8fYY33c
p3paWkxQx4v/cCWwg2vOcuMp2Vrl1z8iYz+eouYV0brQGYZ3r2R7pXnu0HZjW4vR
PWOmkKtmhC1nl5d0QkKtTYOhzt6zd4n5BMxp2Gm1AVJFZQVgnd6F3TE6MrJs3plr
CAca5HoDthKjpzP6rjcw167xzZjdlb7pdL+7bcASYQF85maxxmZ8A8uCLXCNrgnG
QPHH9jVEG8dW+zRHLR4hvEVua0vLpUmHimctRc9fQvTquc4c3hpF5bs/JGYmHSQk
2BrE/1pel2IVAlGq/3/qYuvEoJDSdkVtauYeJmGF57KvXfcdBRolwEc6G4XPAfGx
Z3D7Z/vyQIDdtFNN0Uf5axB24CoPrfqfWDwy9lDyiZpXNZejyeuM2K4mOB+KkHfV
V0JlQBNJtpfwRfR0r+vu7swKjzGhlRf95GXfMQ3u3DBjfSkbm0FvUvowFZWtJNSJ
ll0UTKOQr+V53qSpQ4oKW0IyDRLLRX44NtkDUxhFFVHKFd6Bgp3BC6F3/2u7o8iT
wUvrj+sR0ichgrJZ9qzvBj28c+efBtnRnM3YSddMhGBMmxK3aKZvQ0ubyJMSsPIZ
q4iIHpgvOYfIi2NBHFU9GuTwHPnY0QC+fDGXcbRKVSj4UwsFoaXY/shH9646Qyxp
nUSSazdF2al6tWYJu1znpswk4kiBT2t3wNatTzyvlPTzgmtNgiVAiM1B0kgRK+dS
Trl3342b2WguXnilHs/8HdBwRDElw0EyXa3UcfyWjfmI70eToXcOpl15M81WtVUl
BC6O5sYUlc0m8xTaLEy3wDFn4DV9RFgalcq/S9Rz7gcStMKoW/cSBePAeWHTNp9b
tsdTQwq56Iu4ewXaz1WHtOH3OdKCLlop+amkdL/6oR+NSUQvaV+NYMmMcHKt0jJl
+FrATfAVVyIb2NSMvkZzV9xMIyhiE7Xv9sztKdtw0JY/5obGYkR+JWdrxBJhYKd7
viKLEk7XLRfG0RuyvLDHhHgxae2gTBUYcbQ6BHCjmDatuJcrrhtscJ35LApgjft7
7uTuawyyniECKlB2W4gQ858/R4RdVkdc9aC0/X8e7Uw6TQx/4swlszxLzD57u7Or
IESIGxx5MlOniXyV/tFw2UFPRyMuEKfjIJqjHYJsltb/PDu4oaDrHxhQTBEcOfAw
2ShG6g5n2PYxOtPAFreoMZRqh8Q5Fixn5CsLIXxIEMhkvAPS0DrwVxrFofR6dLRH
Ya3Y8kPtLVZ7amqhfzkerTPtLBOrf/3XovkccYdiOQHkF3DbXAE5AeGZJTQb1lFE
SRTlxrRS+4IMz4KYxBG31Lp0spoP+apDmsEclTDmfWl1c4pIDP4fLVCWazur2Mbi
p56H2pKEIkzVchBoCysTORpDcQh3dYj5TgyIjsaYKcEl3P7Bc8cqgdqswjEDM9Pq
d+X9nEEF7mdIYdGpsWjuVFcsj9Zco+DLodvdCs/GusW+vLCYQmWBUmxqLY0ruvnR
Sjike8fRxMtq/7lReMrbtoAOzB9Z5hieLXcplIfGkUmi5CVydIt0MP4hUW9d5+Gp
DSaLWHD5REy8xmMO/8DmyhBuTvez//GBG2iA7VRNEtS63NROu0l1IMnNc2ooL9Nb
HQfuFyS2x6zKNAZ/+96HrM34zWEQWUu12lAAn2sWNdjW6ErVkrMufqDS86NCy+0C
ekAkvqVDZNZTEL4sSegbVXYRt9SMUgHGWByRsM00WXzA09cMqJ4INMhM26g48dBY
ebqe5/pbbU+4yPEeloT6vXOTZAANseoXYuly41H3IgLG5UVpQhBUzJFK99DpKc7j
trciJ/sDLk24aH62GUONcCE6Ko9GuYIN2R+kekeBbiEUWnC/7PeGI+cnuwkOamMk
Gm9ul6Xqce7KNSWU0ypTP1AStU+Zv6IzaZBbhEh3ul+uMyl6Kc4z0mKpi31jx6qo
+9anlFwOuQRqX0ETTGo8XwqPo5YsAjW4enbBAIwGTmLiL87utT1Jm2UmVSu05vf7
p6npgC1IcajPOwuZIf9DuhQLw9+SrZBedGaSAfrkpdole6jZNQdFsiLXs1Xj0St/
NNFEM3fYwu6uRo4HHsWQdCLV0zCF8jyD8c4yX4bjCMlCv9QGTHlDQZUuQrOd4RHC
Sp/93qPVca93Xdh+EATJdVoyHyJAEtOr6Kh07jaaA3ev9lwbV6lr64nsD/hefE9l
emsia528U4tY2+itWu6SYsNIEXvHFj+wSpmWj4K2KRS6wEDbLFSdV56pZsKUbxmr
eLz++Pg7JwMI/4hCbR2wLgPLYUtRSFvNUerAEeXijp2epZpi8QnXEVo3BKsdKbqr
PpHk3IIcJMjpLTtSKM/m0xr4KTOLZ53G3kd5FoOO4AXyHRre8Lb/GZ6aQ0W2J0HH
9FnpAPICv9ibgG3NdM40c4X3mE6fIAq1slDiq3zF4AXgBJMTOnliC+Lm6+46vjkN
OwRoQI5dyflm+4WS6kcSVkyjT55hr6frRpssSDuDz/mi04gIav0ZtTarcQ6DwTUX
O2Nbll15j9AuaaA/BAh8xpoMF40zZAo5L9nXAP1Go/Vu2BrH6l6rYaewh456iv9t
AHkdQ7VPKzE5CedlcN+AO+zHDU+cMCURqGofFmxHMRskpAFCoXKQ5wmIuzW7r1Q4
pd2AuWHFNrfHxJ8cryYukKHSzfpPMsT7qnrkKgfWdoqY+ur4bll431EAuhjhfyDx
qCFjJ7hVowIl2yxv6vL9S7X6G1xiZVolQzhjI1c0/zjFa3ikJJNd+gFvOtwRZJqv
X0fmY67h5/PQ9c5JvOKjYWHnEYHQS8NtcElZ8+czh4gNEf8Vf+8eHiMe8ISzOtgt
Ef/MAuM8a1ArEorfoGOgqbsnEKf417EQWPfdzPw/oIkouQK9dINGcWLh4swDMp/D
cJ8YuTeVt7k5AuFvSR1T6kzgkfhamUY9zKlt8QRacnqe0sgzDwlm31POD1klRp5M
M2IDE9ZED78sHd4gecl8YETvdt4VkQ53vlNKe7at7LWdU6YDfu2TSVMFztuzHXfr
RcQEoDDHVpxUXjPtloQSn6fsAOR06M/jTAXSOth8HRPdNs94pfNrO9M33NT7U2mc
6OU/OiGysr8Y4QWBjxiF0OWr8ZXRJ7KuiW9uboEUFViD1lUg8PzyX86scpeO39jU
SXrFKKvHcabH3afIFhlPaDZTbSWbsmOJeYAoPkc98y1MXaG8fTWrVEV4fbNiQGlB
zClbGWOG5Kp9FzO0ZR5lp/zpMw8w34JnfIhnbjKT5qGLqRednVy3zvTIK9sD6FOI
96Un0U8277vYmBW2r19EYdMszLAc+fAiJjowWteAKSnpcJWv96knNXkfUOFBGYAA
rXA9w8HImk5OEJw5akBtzoaLUxK9OH9P2w+6IHeAIF4rzGQhSuBZJ/DFidko4sGa
zXFncV/M6g0VaxipyUuQ7QcFNHScuc/9ame3f0NFDEFdQy6bnmIIKG2ZO+gLh+37
CjWU5jbh34wPny3ogyBXyGh2PpquEOJJ8ArE9nDDdJ6hmNre0SJ7YndXFLYjPgB7
via7ZkIxBLPIiMjKFXAPxeLeff7z9ayqCzGi9FEhRQpiK1/FIBFpc975Wsojcr2e
2a63FvvuZ7ZebCkdM6JiNn8C8YcylkxtcXzNBrJnBS+TiWjr4SdauAr9lBhf8ebQ
+FBFlJ0FM3C3lYHMNToMiDhQupV61xHjlVIbxyCdTBYH7g4FBY19G2uO8fiL/Z2Z
/R04rl6oRX9IxbfnZvwSlImiEr2kekBbDhuQxL6d/JbYHH4MwVmlrPF/7CFdVUxv
W1GKGeXW4h4XQoGE10WWNajLDMfk313EBMBwBWWjb2ZF6AsEsuvcXB7lEnVVcXuB
vyHM/Aq2RTdhHyJl9ir2LWryYkTEogLzBetJPp72WxbIughG37SI8XyANYaY9rnD
BgdGOnDNM28ciXVfWV0R9oL69TWgtYD0Y2eY02cfJ1ozbtaS6kikF6yFil+fWinZ
u1PxDUS5OKsWS2eODz9qHFDIwIHJl5r8u7Bnn34fvT0jvgBC08mEYg6eZIbQY3LM
GGLdGnLKyipxaO7vPamsXAs+qCgC9ClQAAR5ZBoVZKO5W//erkb2Fqust0Ng1hL5
+bbiju/eHR1L4xR9AUZt2hsa04RJypHJNieUNkoSfmLBvzQ/pDHgC0wE4HLBQ8Vl
frHOZWqgmNfhFd7l7ttODYgHPnQdzP1Wj3nVaoqIu841Bd58xSBpb/X2+rXbfUAv
S1T68S+RiEzH41htdBtYvxVSoWAK0fVgDD436sqxu4cEkWn3gEhfWvrwWNPIf/eG
ylC+6zDeJSyjfQbpdIygxiVncya5jhjPUugpWKg8tUEeoxAb8QF95J4BvkDj7he0
nQ1YITTf7+UcT9q5HTigJoXdBBd07ZU5b/ae4C29iS1E6yWhhn7ezDpWULS+0t+L
ry2EuJMp7rA+iFDQUjHSyyktkdcIWLWlezd8FZHeVGZCwN95yFHJRzJ9oKBvaWH7
DEO/Gb1x4q0Qg4mKfm3qd7XWjWGA0ahO8+YfW17RHVaotxVP58xp6oeyf5KxVh0x
0pSJqCRXo9UGMVdN7MBkhcw3TQmuE8hF2q7Zml1sImVm/+YvrfOtOlpNNr0j6Sb3
eQK4tAmB/J/6iNEQnStywVjLcr9smHNUUGI/nU3fQ2k+7iVS5UBYXOhLarndARlQ
71Zi244SO5F4Q7k30FCswsrrIMnrZZL7FmCbEl6LkVA5rjohPE8bp0OoZb5H9Vw7
Gbixciz+/0W+HrjprP83yRRmg7WUgZv34NONrHX4E8Wjpg5y3ve0AfIs6zjagdwW
RVBb0cjtHE8EQrlyeAg2/3r1VbKmHG2zXrFEAOpgTi2cxREDSKbEceYEgZ2vX6Ts
5J1hSPmOXpOguB5/tOPRquv3KPePjjRVEyHT64f9NVZ+Bfi9o//wPLV7VSzmqh1v
21wr14jYEtbWd1ewHjcP3AdulAhwrM2qkCy8TsTeNQjmZ40ScsPa3Vj15FU6f9+V
LfqJijsHCeFdXVQW8vXHiq1thK0JXOWg4MxLIHzKjkxtBKXstHPmLMQtSKcP56aP
kDIV0RLBcou3KmsSekS0Ni2MuJwKc6LR0BQjsZqG2HpT+YBgz7cD92k/mT+yjqkO
xWVU/dfhiYb3AV4C+RaF14xc3pHPqj/YgNoTryDvKPeCUpbD+PJnABSExoNwSa+z
j8OaxvHp4JLc1oX/+o/Q5+FrY8XUYTnaZMeHsS2ABtSb5C73C+JtCgtpAfsbJ3GM
lzDQCwNo3GWT/IcFbQI0QZ9SpG/9SbIyyZsHw/gBzYPwzZnvs6EADmgl8VnwBtBe
TwjMLZUNNrbhszhFKwudVOJottXCboOPj2pOBruw083dnUo0jo3CGI9qWmlllSlt
/6wGnYaDKlkS3obRtW5yH1cIv9t/Pk/nPAUe7n54tATBUdxMb0W1bfmc3iJoAE64
3CZe1KAHO/dOnCsOPxk29A6XYcuyMYhxrgUIugX3sIOzwI5PIpdysC75Va4l2T1Z
Kui8nRPxGPHrRmyaQSqjCsT05h85iS7EY9DYAsCM6o4uLWe4hhQ2xo3vEcbbDXkT
HaiPkRCShKx/gjZ+vElZN16BBiEK+SX47eCiiNhojnXirBuhIw3dtez600brna1d
nX4vuyRXYVYQbBfgjc75CcGxH+wXBkYXnbUy1n99JKkS4sKQ46NezK12dPSNcD7j
DGnbdWqfFwdJ39fJoqczyqIpji9xTfxYRGLefo6hfBgSny7jYvnMwYcRawnh/a76
2kKMyN42uV0kQP4+GkYU7li+iM70tu4h1I/kO/jACoA4iZMq2Au98+BXtGUR9HAs
iGvW2FwOq/46KKzzvIGWTwrOsTU1sSmsQJ2E+r/u5v5o+jaLuqpZX6GglE+8RlLs
ApBhjIKcYgjWmcjRh4+7P62LFnQcjMF7JPPYiIrWZ3EwZAGqs0rCzStLgb64YCsM
f+8xrahfc2QtN8iTsRcB9hC5vDVfR68S9Ma1nIAB2dnGa2XeSu+/D2d9OLxLsIoo
OxujtgVAjmscD4wdHmKidw4hxq70T2jju+c6Zh/GL6OULbccZYmshKKzTVpi2Aap
NFm6g5bHXuLdubMp2kzmPgZRzMWJgZXc7qMDWigbLr9vHl0n5+0i1GIWaJZTG3uj
ARHIS08oXUy/Wse1OR9r34uMNSnQZSs2htXCZATgtYPVvayHDKX5+1SB1PrZZPhE
WYMr1PmSwaqL4H8a/3fpjH0g0w+VkB1/nk4Gl22XkjsJ7dUJz6J5gu2Bzt/eiRyd
PZ9rC4C6PNmPOj7bs7dxtaSz1ydEOeCEHHagT0Myda3/jb7KfDKJz8AvwhGh/CT+
lLgJDUeUZBzq8xSKgQkFxQ6kw6Ga4i4uU+fYxDjEgycN2bZAUqTepYuKeQwaMsWp
lYfnljTUmiFgo6w3MEOlMuOPi4om7FkvogVVWd4zOZmpFazW8pJCjEG2J9EMQSK4
GEbXM6gXkiTTW3GQzCQOGeFdRlcrE3qgQNgFql/h+qwg+d2Tt3OrK0jr9SbI1KTh
ei0EK1EFfZmwCP6FPhcdS2HINAwuV40HxNSrIuX8ywGfXdZm6EOetWAcfLZL3vrX
MtOx4O99HVe4m07iwb+wKrCEFZefMdBU8eOSTQEKszNX/LqS0PMXaZO0A1NyfVcV
ez+E9J3s/Z9ut/tsFTXu4Xk+B2Vf1GumVSeU96BQLPQ+d+zFNCvmUum/H0Z156mV
u9vmRY0RolfuEW2+b8dYb0k2BzQ//2a1J/3n2+ncQkPKL1fnSs18qQfgFH+QMM/n
91OFqq9BwpUfSwlWCUdsNyD3Nwq6Ajo6hUu/8Y9dNOC5/FivPvV7S7of1hrArFnm
FtkVfbKZuzflPKQYB6v2RyB2zW1oDPxYpuiqifvaVF1CmOzeaZkQnZzqxEDa3amx
/zkAGm58Tq6z4YsiytRnDbB/Ofb1QtP2hVwGDGv/2ZHZGIG5bkrbV2ZBc6UzSQ/y
ZYqQcOBnGZUkPT9bMbjLdOzvkz1Tx0HKfGJQYO2bxlV8BzZRk79C6ropXxqoMr6R
WraU7piVoyC9cuGdhq5gYXXXWoJ8AVEmfdAEdtalx071hrX7PFEX1UqVu3bXHgtE
0LFSuj2K+CjFaHyuBMpitVpkd9nkzjyx+h6gV407yHuUOlUgrOVaJh/siv4Bl+Si
U1NzajXlUT5UbgOsfTiXpMZk4FbjlylBIYrvWSMyVjkAvyvedtWsI3gsFyQkJ2sO
PZkNFHQ8d7DD9x3EFXrbmEoeGQv+EtdUvvx6aGcO1nqoNrnlOPtghQzevRUxwXOw
WYDIz6V6vr3mZYNHyie8RjRfrdIEzUe86AfCaB8/mrDe0jFIitMNkfctPYZ2Hqpy
YPgHGKpk5QpJ5Ac2a8bb+Z0J9d1U/bmeHZryDzq+ZB+8KZJT2mB+XYLkHBYXFkef
eBNQMz3BEwUuHRIh/9DwWKbZMcpodAPxHND7T4LKnJ28p2GUtee0XnGsdcnFhG1z
UrsILIbi9oMPxXsEgurgeXcWSguKm7x2T5PWCJAtE6eYP7kSF9Xk//+wm5FGjuJM
wM+NLXDJ7f3/uOJsvEyTp7DZSCDL3jzRMCrG+HZKnYkBGoQvbWpkARKkDNxpQfbJ
kRF8CfRplW2qWVYf55xBDmgVq1GNMLN1DFKFl8fALJrNibfFOBWmShb4m796HdwH
i6tJMQCWsb90vhEhjawZwsVMBzjhOULkeLiIIVf/tHr35x/kw2TDBL4UUWI7hU8+
SQotyK8m9UZW5Jpjv+rzv3s8uCafweCz4UNFNmWPPmDmCUvJjH/f/FHkrj8RY8Q9
Pn0NykxYqH1Ok9QPNiDvcmQJOrh4Y0Pj7xlw14brLphrFg+vxCX5T1JDx41cqSCE
/en6ivuu8uNXcs/WBo+fU5IQSxLu6StsKB1jYvqhPfVerl+fu+PpWe2yEWkJf0q7
BVXhfcvQP2RNp+C6L3ZUfJlGY5hiHAKLvDk/1m0/QN26un64nVjgtrVowaD1MBcg
VTtEuqpZ0bbQwVf6dmgES6iDUK6HWqbL/adE8VyXbdmBkFO8XkHSWow6mYIlTsnP
qbjoFhJN1L+d2Ttxpr784h6WZJG00S9t1dInNXEoLH2nF5mzYn3HWHp5mceFHVZn
ccYT9tWTg2d5cD/a9o6tISWd7uI0pEeDou5CXWNqUWCzf2rEfjHszMUpjEA+KhrZ
sXW8gYZbo84u5Y12p9fhdL37bl5jL5rrEqX4/fgoI62lpu6jiWCv5AoMEtXtj0TV
4yF6qy4XplVXbX2Tb9OQIE/nt0FQDD++PgM7xWTCBpSQ980m+bd4Qm8u2vj+XMWP
z+be+yh/0U2AlbJe5t6KLAFg8Yf51Wp/zq6esfDN9ZUdLgkMUuC6xF1/6qw3dSc/
JnovnnSB2rF++F9AXpUlBH4CymzuOZFvw7qbqmwKqNG8dQ/vTTG8xX4r2bwH5c0e
Jdiu+zNHhKQ+WWyeZuKmmV5S73W/rr2AToVsrtpWtt+EDV+1DkaUSWnWDfBkMr2h
bHDt+w2WrIRHenPS4lqQNUhgJ6Oxuyt4R9IiU7wBApiRhvNNpOb9jJiUR8zANaKE
VYoPpDlaPSIQB8R53NWIaSRzwFK+a079BCvlmPcw4BedzhFcDg4fLx+Qily9RNm8
RLSeLTRFTt8VhvplKeVMcWYRLy4sFDtCpk8i3dtUykToLn4qEXb/gv/R5ljXS1xJ
ZtfqUC/TnAeNNArfxEw2IalEDpb+pnUGscjdHjrHl0lNCXRb29E7rRPmaXvqnTNI
ZSyfzqml5VAmAcPYi27ZuhfWhTRmuaXq5G0orDicvVX7RjN+SJp1XO8vB47n4o9i
QIHiaRWPS0E4/Wl6p7J61ya1W82Jgibni0z38K8uPgiECLJg3LLGb/hO71AVihoX
Q/OLqFJBoDUeyBpL5Kjri1NGaPqYzV8qmuMy+s3yVelryTWO3shlIv4Y14tWEdb9
OemVo2UpHkNcij9rKuTI3ZnQb8y7UPE8rFDwtfgktBQKiVukD4jIIcdzsiPSqXdb
Z8c3EzMqQkKrSHjFesVESm1HGXOvyTL59y1+DQCAxM8Knw2lgquzJ/iqNExaLczC
xsoLKSB5VEG62dCahWdyEGU9hxe4Z9R89op06vGbak4QKRfhItWDj5GGYW3AznP8
mBNpZcq8ZwtVoF3Snf043M6dCP6sy28yDx+eyF8BBlmqHQ5RGA4Po9cD4ZKMy6bq
utSA4kfOpg/0X1SAvl2eq8DRn+XyzbFyKwy60QrI+e7b0sxIFLms4S6IGachAj8x
9gsN+CHIiE7MPVlXlO6rfUiZACRRBKZdUBwKkYWIR7xNS7zB1sw2ywljWGh+0uZL
RQl2dzYam1KR+vGiCACW8a7hWyacg1UGLGs9Bo3W7tZ6DTStciEDIIERgW0EGtVj
6BPwbWiz8zwK46p0fsxhKdtfb6vLAXSgemWTc2EUtljvDEi6eXm38hqCQ9mepbak
mC5oQ+KkIXBRXffhId9PuzuEN04sABW8jKnxNqfB3kxRccNMqZYx1VDQV1T8W518
4X5KEAXKwhJmZjz05nAsNEJIpb8WrZlz/Jg35BUzpQVNp9nt5meNUyah2CqSV6JF
kk6Ul4K6+aHp3YQrodga3pKr4XGSNjVi9skdmsESn+EO6SRI+R9M1QQKQyj7mEUv
cI9R2eXruxkHjmbXGafl+P3vyBIkCaO87hadQ6nkFZmRyxT1k0Aj0vdYMoYI6YIC
uxztS4+z3d1w38Oe/NOUboL4FEyhYUHED77cEAQ60AqBEao2D6tkow8u1rqHJXKS
sDzQeDQYySwCMN6skftV6i7/oTsC0h3gS3jeHzNoh6tcPQCRhQttNljnFMGqdyPw
OZ1pxXebIRUT8RgJIWOFiR9tcNUo6ccGZR3RM19ou5Z87de2YfcPFaIjSbKLV3GV
18/tbIOYsKwtIWPUfKhaZUFCnSTDebyGH8gbBlOXlNqcqs4b7mwEFarpoSziUS0C
d4bn7ZHxA9sru1iBWLrx5+fSDZxdX6GRZ/KM+AKw+46tnHqvbw+xQBJ25em9yr29
kU28XGHPkqwTmu6jXPaOLSBaOtoVMrK8nNdl4R0rh0EAM3IASxItUAJ4hBnKVTGt
7EEs7kMmbdh2Dn+qifDwHOcS3lVvOHxKeXcqi60OcyhO71cMFNpXZWkUAiJH+81K
Qr/p4m/Qrg4eUtM5uSTzE/kVofzXmrmk10mmCBllCEklWqAqvrVlj1O4Ss2GgW9Y
yFRiCgnxEantZDTz+/NXjFzxOWoccTyR/uqcMq46rkoONoX4mL3BgAgD3292SdQ9
WVeKGhdNjudKeldkbuuVnbuaMFlYDbpg8I4pnbzIyF4rwXI8sUY2lQrVAsp0Pdl4
ajLiGX1kP/FrN5BztXM79BY75pxlDqL10hgoJ7p+EVLp9d28fIWaUPpyM6wzT9Pl
swqev6b4QQ/q0IWHahQoUnjXH3pobdoSCqdGuHsCPBvd4s8PzEw9qc7V/NUqcAiA
mMf6Fk7lXHydRO6U3gmnf4WRJS0i6NFZv0XC6viOd9wt+6Gq3bMkxFqv3soIQRu9
t8w4eDErMvGf2jIBo4i27nnye63sQyE2j//MmxzH5pjxUKoNjYO6V3AiZC98cOg/
PzZY5uA2C9XYl+ALbfmWXLtpdWIWGoaIFf8bFZ6RqGpsQBhG4To2wJQPnbkSjFfx
CFxIJjx7wXwaxHNlpMa05L6ERk765jtTqqSpUCUkHqLXai+vo/Bfzlo6/+fN62Ws
8liP5HNH7DWiSx2xbPaPzoCwSts2ko403LJRFHR4N5CLJmTswSgg4LHatFh87nhz
CxganLqV5DKtsfjKq5XhP6tmoQJEub+4YTDjUFcIbPL1DmKX+GdDBMr8NVaP1I4i
jgdtEdiwNwwiDJGBmES/GyBiGefFmU5YWo9U1aR31Ub6CngUBbHqpNspcAZq8W6+
3h4vpUHBjPxCpTyAaNC7+eFF1vtbBrk/Q6uXEsC63akUDNMduuH1x2AYS/Jvy7JP
1sbVbCyUiunSRQ6ZhkOXl1jxtVdhNZKSbPMcHPas8o4XlE9ZIza9/BEfsrLBvoAl
oCvuI54/lDkROhCk8w7l963FLMiOciRK4gi1NuykanqkeuktZMJ4KPIW3M19pgUV
yfzogY9ECedcjA1kdalAiGtEhesHIWwgaXfWw8tjSg3fqC0UhNWntdth/PndAD7X
WOTZlQ3YSfSbi5/pUggK7PpzmOpjMV1PhNwYYv6AeH/YM8Ou8/v3vMla3mnKTMSt
spJuOCwXEHklvxmqJJ+nW+DfDtLctyzsiNU39OP9IyMl22It6oAGU3FfMWJRtn4P
OsV2CiyXTxLKpe4YQGckhKB9uvvTOUcdM3rFfapdYyhY95SvdcjF3ZJJpz54/fJ6
2cbS9qc+6etshIlgxgsBHKMBCirZGGVl9kK4BWRKb3X6oHQQIYQ2JaTqsfeU2IqW
LFrut1D85vhCICmijL1FiqFzTvkZSXK5W+ys+2WXpwKokAGFw/xIsvX8jUsyznHV
PYibggc/LU3vpGiv+OV+uCU/x55fBZ2IVY6ODZiA2lN9ssvh2HKUVc5lNWGBxWEz
wjWtWDTJtvdCpvXF0iu/I7jHRxd4nSkjt76rS30SFuTaBN60p9xDe3wWLu6rmGxL
zNLdKBh2YEBLDBQVKJKJeDA+46RC17TuaMKuqwnAQ9lS25C4wjJiIN3z+kBdkruS
PbxZbG2fpeCEvWr1s/cMuvLIiVsJ8/XZWNa9QO/kyeHc85oapfNyRKuz+erApvoH
77dLxg3/E36qCxd48qsatodTEfIMCDCfcf3JPwUN8ZZVZTYc4P4+Gen8kfRYLBwl
q5fecd+/M4YbPs8T2vB5akhM8m56S++xcmEDY7WXxSNs8dV8NqcJ8/HbmKbbQFz+
FscSkWKQoIPX6vNEAUuO61cl9XQenGZg1rz0NBiIpb45KCNLu5GgFHH+16nbzuyA
tspSASr//kjcU2Y3YX/3SaQnE+nAp7EjmcmZoVv+s3rMRnLvaQBerFLnlxb/4yx2
4/NbjC+Vd8blgbwpB5wBWISYImHfji5xCOgkuBYw8svz+Ao4j5OvaKXM90OXU5wf
LYEQOIEqGH+mC3Xg++HUDhXS8/z4vyhAmKZosRNIQHf0wqsL8eUg43aE1TxXFN30
yBKTevPw7WwcUnUUUSLdTMWUC+fdROHzMpKd7kVuo9U5Pb6/KCkJWoXNBCY5DqV4
aREfZ99nS4D8bE5B5WWVQOYmc7HLGIBEhJCu0xV5xKRcBP7eYVe3s1L2cWcJJ3o5
/1PXvJmnZ7vMXfiVbvHiM+DhCro+aEs8mqanf4dTbwV8Ct+Cn8rkMg7/XXm6hen3
5WcRKOM3tfwIDg+k/m2q94Fys3ZpwTUHQIBXGtmG69da4u2c0YZpbcX+sLRM6w2r
lAmWC9UuO2l9sajxcmsTwtRBwALUqWFt5N0Y7Z72Tj0XAPMsrWdrDsfLxefMjS9/
hVG2jJIqGQdOv3HtlVSerN5xA5BZX3sX9ZiDssKq8mS32TcIDusSrA6Bqlks3LY9
ldkKXAwgxgTZxz5Fl3hWrwY+yY6fu1RkDKYhoLGdPSn8LKm+YQ8Wv1fEBmip3h3S
S7ZKBYmLV8jk8yxHdv0NUYwT3wAf79TYPhzolAh2I5pXPWlCaPbA09kKlqt3ONIY
SYwM+a5RR6aVVvgFqGP7Qeosg6bzlfFsOlbVqyVD6zaqQC5vUYQl0s4ryf/VVMM2
3D0jhu8FRkmewePsey7Q+DJns4p8Eb9cqhxRbmllVUjuQj43l5Wc8EGInctfaWhn
YWglb4JDZSL5ph/holrmLbJc8EgaeMFJm2kjni8EEamzdpSWBHdFe2iasGfOuXyx
f+cc4+Jc524BR/GLSR07d2m9KNL4ebg9qJaqIekMuSVtuMGLRDUirOC9Sa1efBsJ
ptD63LdbQ/O/bGy9GCSB2uojlA2sOinf7nQtbwW45K1JLsWWc3X84ZBAGp4CWgyg
n3eW7S47ALcE4bAn89aqBVZxX64gd+9C5e1IFshsianpBU3kjlEMOOfjk/eRZx9k
WjfJxvBFALTyAGQnRtycGqzvXez0N1X50UBbuWC9on9L9btfdY6R33YTqEc4gXLs
vSjawHRbTigAg46QUUciW1WrdfUPpROBAp6UWYo/nk1RNAfdQuZ6w7v8jVCEBc9i
CteNV5mxa6Lq0BFsBh5UHxRHDqmMWPmlgVHuGEQ+YHLoJPVy5yCpSbgtt+bRsAem
WeumDEzeatco54yCXFpz8zHrBtcWEea8M03cdZOBLgEoXZ1Tc3Pgc4+UNVkYz7Un
065K3lipMurVt7B3rVMSo14Ti0ZD5VY5/x9TWELHl0EJRwpxS/oRdFnOa/vS5/iq
yiZixnTSRKfokywpY1MxWsY5/lmW4lQt/S8JajqN87GhEUC3lUS2zhZW8JqI5Ubb
+80p9BPXTG13B7dkCaCLYeP2S3aKPCwJQcinHsVNyEc23IX1LXfo1hUEIkD/Xtt0
eOja19OzkbgRtmlBrG3Xx/npMGJDMbt2+yAsBGTKUUkOB3cWcEASqu+L3TMEjHy+
Dotb1Fk7qjeOibrf0qOx8BrJ6Q4Pgw+17Keu9D9sDrFtiKLdiI73rWRFPWug4vPX
6BWKzPanRIDupjhV5Qj6q7hQV8XERE0sg+bZQvVZjzLrS1LgLSA24nfJNhEj/UuS
lwW1nald+vNA/lm+1UccRhzd9L7BqyRsQCGL86xhG9fnz7HTUuBQYHQMLcsAVIAv
8Y6DAA+I7vZXTepjPXH4c9WfxkVpxue5hMOt1YxM1wfzY9H7uEx2lDcdV9hQwcmL
TmN8NbgW2HPgC0vFaSVsEUsH4Veuxn74nRyleibdaOBpcmT6cAqanIbTtImmKVD1
SZdd7y6IPyaLre6A851eJgOIHiPXHRq9qL99FAIZuP2d3hoFdcVvX3J92HvXbpLH
veLnNVl9+QABDvlV61u2irV69f9josqz2rMAbKuCxKhWgVUaU6rgcEqSBTF4vxJ3
ST8mC9He9+A0sUAwx8ZDoADnkahcp1Qw3We4CEAr+OjyQIQ+jNz5zcjV3DyXZH6d
oCGoTquZtrRg0wgBOVIhOI4BL1WkcKOYgXCmmOyIHogj48Zl+KSpgWRfeqlLsabb
uKscJtMWS6n+iEUoN90S4ANy81qYSrqaKWqOMdvuTZUMc9ChG3wIBpBmEgRtxTqM
msmDzdx2ZcXvLs1kNS5rVZt7szDnsPeGPznmRKlgfkELDhSQl2ZcL8DMGChvGII+
f30knuHxzKk1l4DDwxqzFKa4fcTIB0wnc8FUka7L7j5xlXIbhBJKWmSKsTm4J/6e
bee3DpzGqloRjNu2Y08+8uOEDcj2ZBxRo2Fw8NRx2zx9UQg4cxncCoU3wXl9yW9l
idZdCene7tHLEOtC+VKADxfw/jv3hWxbP0D+8CYC5Mu98v9Gg186t0omWmMqsPf4
yN6YY0dCxvEJR7jkjN04K5qePgViRWpQT/Kpe05Y1eoCwq1uC3B26g4gtct3R4VO
XkqoF7auLup/Qh2jmEYPBMZi1P+REsHu786qKgq4kyxj8uIcosjmqIJ9I03HQGeV
8Q2vj57YjZwYd7ZUe090UFH5ufGSaM35GfgSt9ikoalp4GlHkZlOj9ESzOZ/WsM2
M4A38fEad8U2J/hoIHOS1Dzk2v5AlAEJ2PqX/PjHy2J8Nx7ZYOv0AL7jl3+rI4/M
ufdd9KU8Y0B5PycUlt4x6kXSpp/3Mu1t5YYZw4iMmPYPbMjVfaEVVptg+1BKpsO0
+KmhE4t0vf6U2Ci87yuOsTL+CGqnccfFBCaQupEfiHii6sU7wS4a3r6cVbaVXBit
ZaP/LzP5rqy8bI6B8RMBVxh6M914b3t7xw2/8A9R+2+70nj9kVqu6XZNnZruaDYE
n4DOdEqUOrH/ZRuXIx8l9bANjPJGFUbmUk9DX04t7rxusWEtA5cAWjpNB2jkBd+5
3mOp4o6G7TJahbQEeQp1sP0fgL9/eZvHnLJ7cbdUECoUqlQCXMuomqLL4qEQw6U5
adK6E9l82H3DrOJGbc3YcjbJCKAbPvUoKOIj3I3940dTTilbfHf8u9vd/RP8xQtf
GV3OnBbEi+yg6pQ/9Jsbdgfaid567K+rHI0lCC4psfiEDElMy4NLgmfrzIgdQ/ur
WzfVUTisokOf9l5H/AJPk40PkYplbbQOCLtmkGG+uEYy7r2pUBnCdDimbEOLPpX4
DBi80Av6wx5pSz4EUrrmzZqOfS7eTZ8/wmiO8bKsEJwyFYqeeoufhOji8wvfFYmB
rBUN2G9+na/vvIZhqLJ0uySCJ1LUJHG2chEtl+EEZSQi4lLTSU/OKQAjDDTv6JG0
RjIMFVVX5cDRTxEd9EL1Y/44tdbi5JB3SP3UfTV3lITgWbUpTAc7sDKLLT91iE4b
kmIYeLKY16UE9UdzVJqeBSKYjp92BitdCb264BQ2T9MHSrxGd3FBG/Pz5n8nd5nw
7cCbSLeQln5QF1LqriuqO0gW+ut+OOVbZXzW/QuCN4Ug0bm95Kzt1EaGlxkdEn0g
fdoAoMdYvzT9thkpDRyK3KbbtMGxIRcdtYHjGPQhDyVQuajGlk76qIylG+xOpmg0
OAGBF9T05pkvHI2gfDNv8A8x+QzCEyyFcxVmVlbeDK/YWnTzNGLyXCRrKoQysFj6
mR6Ysi0nbbeK/xAOygQYnJsl7Fw5DnYdF07KeK8fuEEndDO4Y8AI5FdQ1lF8ul6/
CsfSDvDDzac2e+v4yJ7zjpYfH3MSG3hwg9A8MrYrt5uyW7QLtTfv82RZ+1j/j7Vt
BPxv7dNcZSRUiTew8QjmaVa87J9rNnG7Xfs5vlxGKKtvzBS+DnCQU529O9asn3/R
Wr+WqWF/DMmjxEjOZliTgA5FXjS6EAChg+FZnKT7lu/q4WdlvQ0Ll2TJmxMGED32
RWk4iTagou0ev/966cWNIkVWHWM/PkDxfLt2tnw3RnrpqoQyiNR/OH6vTffGvmls
XQ75CqNzccvlSoUta4G4FnEM6IOY11Wd3/6Zpo+jjkPZ81dagGMGcCcQcsTYdALN
tmJq+xG53aDQFJ/k0tx/JVOkgFYOp0ypqWU9ZNtXK2eOIsdQ+4D6ICZr7Pun5JdF
XZCteS4kZPKqNP17+tKR8XCa8mrg6Y/sp5YZ7Zpm8pWZ4PZi2olzLYwEp2MnhJit
U3XagXI+4TM8hA0y9HfB2PTiOrepsR4Ezfon/l2okgSFXlHQD7ALirs3tplb+D4w
KtcZ6KkPazkOluwV5wKO+zltrOyqTLM1jrkIHJXm72IEaRamX3I02AjxesTmseO/
ZSD0fdNnmVS14i32puh8WovVtcN7wouAB8WNlQbvuh1RO/PwABV8xi+qPVPGBTQr
nMUjaiouSv77mVr/vh5NQx25L+maM5q1m98K9sC2IdtJTIsGGbJmArpLBCVDWkJm
IvXxEiI89f7+ssp+NV6xPslEbv1DhNDS9d4sxwnCQAQ6vZ1ZjCTXsYwx8YUJgqNg
ThEpTRX9vv3H4nDJhxkj/fPf6jJVbG0JV54iq5o/80HFuwxDxmKQL5wT58hAhoHk
0d0xTrft1B7yeC+pUa+whUz1v0NV/2uRVE0AaMK2IUHWshoELQrfQoXpUBdycwVP
xyZ8kBsL42wwcMDesxHhc82HCj/0el7RUB2E1fs8b22H9H0eTYmuO2kyeCdgGT3+
pAUWkSlchOVjuM0s3KhAVbtzEUw0A40uiXJCVak0+dW/kKTs5ntmIZWvW4Oulhhy
2nf6CTnroCVinmq6uNBMIca5EUI88ZKvet3iZaJQzlUjFrrCJNwsMDkYpOoJR8Br
AfmlR0QNSF/Hu2dU9+IxUJujUUClYw8JwZo15oixtYps5wEvIAp+zQVdNYawUEhM
TGb+httXu4UNRHeF73u5se+BYr/AWXJQqV9ZGzaC7zeCtFWdorGss9tLOYBTH/WB
1u0H+Sb0qfeMVxy9gABOoh5DmtQiIkK8QwWvLCy9r8YRx2T/vOynJ5LxKYhEghyf
nr7Dbt2y3/fnGwhq4ejedOTz8GktEInjDfuq9BX8SV+iZ01APr64lTOxluBlRwXY
rlqOOX/AkFK5DoQyr4QTO8pJ3kZdrI6t+hhO2QF61vDY6h4tcskwxED0sCSQ55rp
PYv202aVGCKLABR31jRcY2GA1jc4B7dxzAKdH9yxkmaBLEnv7kWuvhDneY5b4MHo
tlCXjH90VawUOmpDLEtbsY1whyMiJMoz195pgGGHkyXIN7cmk7JUji5J5fIy4t80
V5wQP5d8/eAT4uCvYpYh7kXxWHVx52C0XX2v1IALZTS/BCV7dtikOOjvhq7c2pXC
VerQpVeatvK5w+MEbg0nfBzT2doH+S9g7K29lEDEucmQlpSKd5YVan49/DtCEC8W
yrJ74H/rX7vnngWQqkmDvFPc+J1/WlEii40fncw2aM8Ea62WTdcZICCCBd4rwip7
Ts7CVtZdpOlWufCfTHp6SqkuoZoSHcycOHqA67hlXLpZisu2pOVt0k6XtJ9eU2w8
jg3z5BF+LBB7TVdCEj0kNt5AX05tdElKLFknf84P7Q4GPqs+iFvPbwdBBBSBK5GF
ZzK8aATPqWoCN0MvFUJKWX9vZrV6iN+jlMmwhz2BW54azi56f4jiE/p7akVm+1rY
1Z1tc2SrQct9/wXbyyve3okQKB8d0vwdt4BvMwHfEwiYVHoYJJUzG1cvo8lJW3Pj
7CzOMXc+AZnmiqVaJElGAD+HCBLounYBdeaNC1BLCjHAE90nwoFxT6Fv4MhiGoZ7
xdrODiHWcOfWd7TGp37mtIWXHjMsUULPNe6QTC4xmanJCL8DczUih4V5jQY325++
G7vc43Kvujepy33dQtQIld+02DTwOZaEErDo/QT995QeAWVhxJPbNK8DTlx6pTrd
+6qRYFN2JziQIqI5yUWuTU1YP+CEaxRi9OnivfQXvZ5m0S7YY/LRNxXXyudXCn4j
9TK9z+2BF6EQZ4U4TTmhhFquMDG8lzx+lWB++5u3Y7QPEsUQeSLYMmnA1zSyXEGl
rrz0nYDmRW7XAcW9thQPCHnJJGldB1xl4MiKbmVUnPEJQQPU4/uJoMtvgWRN9Ssg
PQvG5QlnjQ44CdyUo2CMrM61Df5WVnJsejsfvVE8ofK4OcNFEl8QZX8XJLN/nTAY
rMNNBrasAnmbwmqWrPZ+NhCdULQSa2QaiGV9lyE68ZWO2BuvbUJhbbjCdHry8xay
xpfj/V6EG8YSfFKLVpJNKhPvSo4JEhybmAlnp87cFIZT470KDUFyFH52PP7RswBV
oqgFbfTKIQIdEy8B5Dg6eoEkCCthxCM5uZ7VM1RPjVueCWlzOUVf3WeDq4OuNzGv
4fJx9XqIpQcr5fl0EBEzlhwhlN4LvVhY0gHaprT/ErdZbN/wSXfKGA+YfADXBit5
bo5myZAkUrspt7FTQZ+hJd8PN8XBxC2Lje2MxUq0osKuieFdCZVSIK5/dQu8Hv2e
OrDuVUgmFzY4IbPpfeOqnObp4Czx8FLjBClaxK7Qn4PsL0i8XB8uHZlg1YTqQJS1
8Ei3Eo3hQYbNG2luCrpTbX6ihNvbc1ETb89fKwocIBJojBlF0xfdWgNprTGRXpBY
TZUUHdbplIC8/jE2d71jUlg2m+4+wLJmhFpLhXNFRlzHNORGVv59SBlNldodGRSx
BL+qODeD6Av0401EooncWhaZjUZ/dzDDuNCvTBeXa6IiHoTRdIvan/zzAyqkU3qh
HDYSQtq5meRIlx/jIJ61SLZcweA69oxsK7OVFiiMT9jlooWfRWKxW8+3etTYK8Ox
p8/rq12GwBCiariNUtEa3iOdHdjz5SzDtwxcyPB94D4V4lLZSA8ln6uHMu2xx5CL
9hgF1xDQwxwVYzQ03P5t3Hf1GcuJjvjTklK/VPfVNg1gjKPA849uMPCpgCBzINxJ
XNc45N1IXlhEsC976sLxdoXTbnej0ZPnaGqBInOcLJLsIXf1hcqHNF8jH7AzSj6R
R9IdCJpE7ZdJ5EoTqMygah1EqeqMgmJdfh+R6vD8gsd0skkFXELWhdL9RzmAREf5
4ZDwsWtXKvSCnNHwIr6KCDeUgJa7TDsY9X4sXTQQTZBEbU73H2dI5x0V/bJdF6gi
72SGZToLPgjzHXejKuBjfjvX1WCHIj4YHfBxXVIn8X7GOvJENi2tiGh1M/gkSgMa
QT/yzG9lv+14nWYwnPIUhs755M+Gzk0GHojeDMvnF+Qfxjdq/WVtypo0WwdjGyX9
Ca2ZZxrxps9sYIZ1Yb9+ViZK9yca2J93cvutBZfkIygUssNTEFkJjV70xL9OPxFs
sB0N4tT06YK/+phQMCZnf/k9D84L9jBtdqxY8fF8rxgge/RhDme9BIdwTuKt5kwP
FjWjVRySmHGSHtccgD+FUtzQjx7UBCCTm75kpFsFMsvjw/lKOZQx3EesPgQmikr1
AVtuY7n+KMKGrWeHOTXct70Fhgiq0eh3cyZ3Sbi7GgGv3qQQeIhVVq3qjyFp4Atg
c/VRbNQnRAohAEHYe1hOohtFj5cGzg4CPUjb549fABZwl/poztZXSjzHoh6ecfT2
wbrZwvEHWqdEnQFKcTfVgW9X5yR/1Ol0rWdyK09xYmu3cDMFsezX0lMGFDTHBFGT
UoUXvo1JzRuvaAmVWzGLTyVHyNZgU6K/f/mq5ioqT4qsrHM3UMjBnWG2tILLbWsG
8j+ZeixonzL3gPutZHHWlkjBNErgX4nm1H9r7BZtasf9kAsrvesKAJwk6xxUODHd
aKfcCL+TQpXHcCRCKp4fK9FO3M5/fD4b3VLBskhdP0miVYMWMNW65HtLZelNe9Jt
sblNKI00Xn4k0y4cpNwh4a2b/JLg8lsxhkqnw76ZZaeiMvoXXfBKkQgeQ2OlROvB
JzhrBm5FsseChYvSIdWcIqGn+7jSFdn3cC2+ISxb+uFUpuPZMYUcCYc4o/RoHkq/
m086BrgZXmY/HgoRcqtNrMuEXWCLcRvQx5tqW2SOWhJ/539B4sO6mw/RLzaEyMpE
9O72todmObJwd8nIgKKCRODCOcZ8AWLGCd6XcleYK8ghHL9Xegmgvov/3zSQlyNh
cQTtXV4s+wZM18lt3C+ObZveUgDjTQCiFCgnmB4Zi+JlwMa6fwH0EjdSAuV3cq98
T5SDTf4iiIKeAnRDe8Jodj+KKD0Y1SGpej7WZ5vDtqfmcefFpzqqJ/sW8yopp8e8
InT8PAOnjpCH1moEufAtWdSduSnfiq1+0gApPauXPEz6n0LBnX5Qwhho2TNSe1Lm
ErU+uyWSSWlXL2D8gxHcXuf9SRv4JbWSjCEHFzX8TMUg/ovfPKYKu7mVGUy7a6gN
dyEhkOhA4rXnV7bCizytmdqfIuBQAYt+FT4Ds+IoQgKuZN/LDXfhVOqnH8f4Q0M2
KFQjM7RT8JSv9BKO02ulATA5m+WJKpDPyDGx2oqjt3fKrlXBzOPLLQxUcV1luGC+
rHymetT387qoS01GgAHAVvhn3myWUU24uA4+T//QsFefwG1O4JSj18+L4icK5wR4
NCWe3pi9b60wpsBXnDAtGQj5mbUcFYG3WRjDUcHMoF8d++kokBCLZ1a0MA69iYmZ
6toV7w1yWOezdAabSGzDlfA/ipgAqBWjmw/yu3MmB1xvjMA8lLInDCJSLOBB4zW0
IcdpFWO5wHrbLu3+RggEwQrYxwucbAzPneSZjFHVVuraPZiYYRoIq6TpuYyahD+1
PMefodNn7eAKWsA/uS14W07hyJn4qdguuWifjsQAl3do/rHMiCTbBvCmxU78UT34
Bf2MFYeX1vDhNQvebgT4qq+S7tyrdM/IvffWMQOsMaS08oh5S4KVelNShmsxFjFR
2UjCzjcT/EPs03y0CauWksaWlmCKOm8JYy5riIhZEcsOgz2P1VD4OrsTv9ms65Ja
AT63zm6fRRXsRCV8jFelZi9VBLoGb35Pddnskk80N+iupDwVlai6bD2Jh0a5FVSC
jcnWOcBKz5JpXeMYLC5ck6DJ6da1Q53SfasMwNu5UG+ZSMiM2eBve19J5WNArBXH
jk4ChepPF5+r3RbByRZxUMqokbXTOMXPRlMDykzn0An8he9JvR1shJZ0d5h2ULI4
foDtKt3BIALhPFxA3uBd1eZoyRCoPqJ7oHf7Djr5n2VKgcVMQlbzK6VwOu6Z7NPb
qUsQxX8cdsacZt5Cj6NaIJpdTonZ4A6GCF9E82yQb+2N0j6sE0bzw0Em+j50Ik7y
O14JLnTEf8w1MxKB/15tPTr1Fer+ocTw7M9piOEuqzwP8Ml3cn5+V9n3gLs+Eyej
8+jGZkv4FVK/WWS1ya+z12dSAAlgjl+frN22RjAy5d3LaKcqO2V7EEAjb3mriSbv
mKLim+eX66fw+yAsWOLBkKQLaTZc6hkpzdm9g5x+/e9e+xy2XTpgjEHXHDKNqbCS
Bjn1iTr/iLwoMbE6WeoxGUSdd6wWHOnCogSWoYDtNukwPQt1t0tDWvErUVcl3m3h
XpiCNL1OItr+JRhMWQ8BqYcHkcd+tHR7q0od0dbQKrFYwFQQiNZPACBbNY7JEFjq
55bQlEHCGZaf/468jJ5m7tLWashoAIWEW1wAX8dYwTdgFSJjDDN6v/Yhir8gf2gn
fEVlh0vLMJnXiIStKXitxAvXu1b6446HKof4KHLyz11cskQmXRhX9KYWB3iQEQyF
zVqn/QkANBQhF8/2J/LJ/0VUIMcezz+6vq0XZRXUD4AjmbObSqko4Ydze15qh1Qo
rZlNVy21TeunIKJWRos0/5tb3OhUESXFzJBKOjyUL12yZl3f79/QaEw7HBNl7P/Q
sUkNUcn7MCz2QBH8gubU+yZNG/FvDMgA5vfDBHYy5vjdRj+mzsW310fDSuhZlIpB
XDKFPoqRK+ux5tMTJ/lgqpfVNvLmS2Zc/5B9HFe4ES+8QtJ+tHa65MmKQLdVB8l8
J7z3QJGPlScul1rXO5jvgDrGfNAgs05RWB6nwv/jt6bSiIEQFY2vmL3dsvMVTlIn
2CxHcTRazg8QRl12eNgj0dEqaM0QzSiBazxjmh1TTo76XOhPwEvqq9LZ+ev5Jn/a
j7jai3yFDUemX/OvexFC5WYkRXdEJsmODbEXDH8CaCXWi+5lcGap8xXZNd4OVjSg
GRhkZn0KXZ2txB1Pks1XTXW5ghwVfLYdm5UtbWd/7JBMOzHquBR8GwB3mRSRdOQ2
l4skluOE8ACDBzQz9XIHysaBXX6hkRBN9P2sFb76u277+oFwEXBg31qkRc4lcI8N
vdhFNuqQe87TGRMeAvz/kXDSnVNyqiLSZXH7dUf4S5HI8llBLAyS51VirlBkCWpH
tmknpCci/ZUr93Ozh6xP9wAAPHGVuA8xlzOTTVpVcfvi8OAsDlqwF8WmGKA81N9s
ho+n2xgWwvuA0sL8kNXJnaN7ZfBuxhf2bdAIvmqnNawAO/YczRzW9evIlaBY8Td2
TgiKW66wtPQ8/KDCXp+6ba7aD+ubPD9hxyhbAwohO6c+C5anr0FDwqNhYu8gYZFg
AyLYli748wzAAuYh1MRUM5syKCjzx2Ucvv9GJnRWI4/ZGbEUjGLmsyX0MJBJRRHG
h4N8Ji8uG8ncJr3DWo7Hxtq02w5o3drR0QD7Rvp62jYSVaIMxh8ncRo/JCDLZwlj
5vH4+rDwU6LPehGaZI6H7XPxFhmAjCSIU6C93RBd6JICNk21eqRQjGpfzWxXcY/5
RKbgL7unT7TZL3MrcNrCOeCnKyRgKdZ1z08QPoB2A1VZRvppf2/3HCWaB3+LEr4z
IwBhuKXrQMfjeepvVHdhx0kZJz2WbURygpTSLD3FJObsBu8NRAqmWhZEfVZQRifn
1XiteHZGhGW9fGm/RyJCemph9oaKUvOsl4l0KWUkefG7iyWu/A0whFOpHRGpVjX1
xg2B7GeaqW+dL6myOsDYNMz0p0M45BMH00HvQVSocvYaddl3UxG9B9+VyZ7iYWXr
RQo120oc3010c/3Ah+OXlXrV2cFSMykp9EgNx7wmLD4RsN/2k077f1Q5DwOqv8WR
/LH5t2dbBO6jx1i6gtZeRh7LsVegqNN0orDIXYK21oAisxqr0IJXwfh1b/0goiba
+A+THJs4rwSBedMOTidtteaLc/faZLHPuTpqkTe5xaUbFsUkJziFA98MlBiS6m8D
ZjnOE+ZLYxTWJmpDRMw65efzxfc2Lx8d4PGd1dkGOX5KfUpIofnBpzpn3ivt71ia
z3hKq0+gJtM0AfP0RoLxs3RQxKy+QICs9nO0BzDuKg5tf+eGoXzGdAfOhvXJn1in
b8x7PK/v9/3uGJ8YEo4kVKxEyTr2rwRd2SmPo5qsMQqZUk1jPA74HpEtDbIxIsh2
pMpsSaKfB9xo4LMfCcD7Nzi+o7plfNMLDbZ5cW7+5dNH3Ch0FbpNODlDoa86mkWK
g6lnt4spD0vSjVdo1A5zYF+eVX2hUnzRlTx6cKBYZMhmlRsfQBOybK8ifikOBIzU
/zEvSVyKg/fr9S/DWwz0IDBZBmn3/Ya4jtZweg7yAQ4FAGZdDZeKYKwwpYs/EJ0Z
3uaEOKLcTtbkhcj+/IjLVz/AqcAYvWIJd4o7sbx7kO9WFvpeJUsx1vu/Zi2/GF1A
HVfUEHlas1DBhwfi4P9vIdeZ9EPDdZy6Fw2CeTcAPcb7k6t3QXpJV6PEG1mSQcYf
eEpU9dBvv4Or8AGmxvH2YJhExzbff1bN8vVY66NuFSVmHjoT1/1l8hyA0xzNQMDR
vDR2q7uoB9jMLTykyqzVIgdpraBStuyXYu6yp96eqAThsqK9ptOfeaTPqNpo/1w/
dFAB43mTVnXeqCG8dCkV9dRAMnWFxVOleSDJN803+y5U0jpJC1RZaEwKVVPjvDBp
6KNkySWOl3OsPhe7iA38ExsLeaQ5p0lG2e30nqfRuEvu+k7dArkLJQyZUQ9KVuSF
SXBQNkIYJHiMwTETu2QwvI7Y+yIiihtK3Achu9HsjjTF0mywPIPgmrbSZmmHTboH
Y6lbWCS1t4tc3xTsFfHeGrHw5FdThgwst+CFwtQZG7KxwVCeyavXUr7F/Km6Ksqy
jI6IBAkY38ojZEIHKuuIPJV1mjkbtI7bBAiAneeRLmvb5cWKPQ/+sSLCL5Os5bgj
AgiCbj9dfXjk0I05K3iWdjEAYPUWYLsylOqSBO80F7FFkwoT5Ngr6H5AFWqyMegG
DHr7nsJctozMD+FPHYg6Ri+LcIfHpqIXGWP/B2aOf2IUoTYRQzmTUrS43ZB5HRkx
5OGWI+YDdpHXOhoNHgvc+gQTNFMeVVXgb84na45BxusRQReF85xmczhLeaNDbpLG
cd9aul8oTBuqhYE0vG0olxpeir52bwfSIgqetmjPAuyeRsOnQZ1iZ3/rc5RtOG8g
V2eu+G7lzfvuylqFkAp8YUdWxXzQeAqGTpsIYWQBwHa1+585dVt3FGnqoIDgZ6RE
CceHo5BJ357Yr65S/Qn/qztVTW4NOOTbcvT8vE9a00zSPycsH1hP6YicNBG7WsOO
Zgc2mQQF7TGCr88s0XJTk8zR1ZQ83jVyocZMohKAveYQ5hFJB+DCYJCunWpLBRBS
2PNYJc2LrXFEaf1WL8GCuwTnGm8vVZ1TKmiGN5MqTUhnWoka9rWBLVzIYEhMfXgc
5oNBX/s1UwAsh1jA84gRI64kB5kL8Byi1edMizivFqYcfR57dZbM1alsQGlUaKwn
uJqAChAyfC1rzoVlzXuKD77o9Q1VJRGc+ghb5NvZKB0rx6VA0C4wLLcLkBDLhhAa
k9lyUgD49ENwknNz4HPM7TMRvaPwHC3D7XObevc6a7m4/PPIoTn4oPbgengEBB+M
OCp+4QZRKa8V1AB2l3x1zBZPJL0KlxfSTZaPZh9B+9054KMa7tPZTW5uW/ozQ/w7
K29+iEjlib3k3YqrDCgG6ITrE7AiB6fAem4ZMqEz1HEjn77YsgfXUVXai3LvVLOh
sSNdcTK5PQQSR4+cKjbczei9AKp7qC2dOVGLYGF51plzH/CtHiWCVGD5ghppo8BB
DZpPYxnU+7ZSyn85gF2HK/qNJJo/FqIcCpXZ090xdIpTu2eOL1AGRAwuBfEgHc43
ZruIyZoOaTL0ShtueR5NSlkhXfKo8ZUQaZ2BU3o174ftjR4tslBB843SMpe9DNH3
izkVF15MHj4jP/ojrrOgn0pkqtIQnG9pmq6m8IgFxR8Mnp2HuEkXzCfsM75Zj+/R
GBKBeztZcnuyLOS8cSWPoOjgCFH7Kq5AR3xe/HwsDaDwjufawFmRi3vU8tlT0uTm
T5C+9bTHCrbY20xJLS9LTCm6X2mLECe+ToLI7c1B57Kp4FQ8737+Xq0hQUnT+ZFJ
O73LoD4/JXeaE9QPyTdv8djHTlRAiIwZq6DTNDP7nQEp6ixsnzvhcESi+wwDmpOj
dNTYh5hVFrgEjf4/bHD/5d/c0IA3Q4YdzOyJhhYeePM17Q8oS4oPGtAagRrWi1ax
FQJ3L5xDE0hXIb8/B3WJBEfDZ2b19slrMM992ZwxyehV3EmmgF7FQ9PxUUO0ctKw
zuIlPGV/4UEr7eh7xv2vc2eQEN/J1YFoo3CGkwCLL0/6VFbn55DHFnf0JQgDnrqz
XpMlLxohq9yv2BvI2BFk7DPZiXZJWfd8VJTARIbjvZWtGlGBSybr+hDzF/0EBtB1
kg8hzl84eMqrKflxx8+jHuqemOU7NlarHiXiXOJX6zYnvUMX5bGrkUh0FImmZSrS
Ars2e6xBzxVxI80jXikqi7B0o4POA96aQIPguObVqRSoeDkrsH9Q0WqASTvubOq9
sX3GS4QfSnsRQpVS6f5CIP2Gra2AjPkAre4ZNelAkJpjaMMotW/D6LlJQK+VwHMw
s6BG5xtCyMtSYSoBfFncOukNjV5l0RDUScsvzJ45gsv1WKLL7MdssiSF76EyXh8y
xVJtsNQHMMpusgh5UeoxQoeN3uXDkMfJwuAIx5HppPzlZJaHrD57ahry/wfPuQjP
5+ssxvriUnStc0pipvUtxsutc3Jbs+/6HUGZLUEc+mvLhkS94joORsmPhyb6OtPz
XXTwa0mkQgLNXsFe2SuAdXlA3jXJxlV2+zbCTHhXFVDeBvpf1e5fCJORWis8E8cX
Dl0xz6cs9kOP761z5z+ePxQL/dFQNDtkalSbHY2MmrbmukTa4zlP3SHAbYAqO1un
t7LTt1gzZVkunG0DOj7+XAcyZt+k6Ia6P+yF1q9DzBlMSzlr9SPy5zq7MmSoemwY
7PasJJ89FDGSfA0uFBnan+uUfZZkwAtgAEWLZdS8kn6yEILTqcvA5I3jhjMSs+NK
V5+iMUA34YNe7LxhSikadxClyR+GOwMFAI38RycTKeS00TdvQN4KU2AZcA0ffsem
4/X3KpitmKGhkKSWyza13L4qeFYkzFMCoga5ezxSAgRGwd3NCDiEW/qHhvTYTd5f
Ct+kx+KMRKXv6nbzOBWXSsN8k3IOR3Z95u/feFIdgVmfepTCwNQsZDkVUKCuBFB6
BDYLEdIEj0ASf3cO8fvQ5MXwtIK0G5L6ttpRqF4P53bIdSssvzXsJ8hWLiYtGXPW
5GzZE4sW69yXLu2/Nz+QbSHGipeyB/eveCyQG8iFfGfc6JixKrh/S3lLZv/3eiiU
PmmYpymjPxe8H4yHVgTQQE8C96jO2wiseMr3GVlACLQZEc+REYIVtxAWZ+5Lok/T
GHO6k3Ut0z6nnvA0u7iElSlBkfOYzF4AzMCGW3DBNdG6kkY5FDRJ0o7QxeNWvtz9
xUwTC+DckuVMgoDbFXg0WhPGxcMBFvVfo4to1WuquBWUs2aJO4UdAEZcZf5N+utd
xLoTPKZUziKXqWfe9Xa+Y8/BvUIx7VMPRW6skYS/RpJdLQCjQz3anxLZvO2CBjr6
Oc5fgzGqqeqAaYPn5j4oY5RTYGpc90G9mUvnGmte5EuivRMrnxxnGVVllXq0ZUQ1
oV7cZHd33i4lOY02x4cq47voBmzlFDnix5rkN3Ql0p4CfG01spmLYlUVozpuDDKA
I9Y+igJdotxRneUmVn6VgspnP9Hzyvl89rvT8otyfSIkQe5nRIK7/A168Pbs2gs2
reCuG9Lkx3Q4pqgEXZksqNbdatFWfQVIOdcNrEAZQ5zVsotUTvjQpzN6RGJX/LNx
MoiRNVNpklHwgsm5cQiKNXvNHDMxd8iIEeP6OWJ7SitYnwS94GTqGoQkiRIJ3lWi
Zz/9lfPsRNqEk3ZDBdaX1MyTEJxqZkF3lk9mj6NxeXG+DUiO8Su/VryZrFpdZE6Z
3I8YwHF2M97r/lOsa3pr5ZyvA+YtSJaBpUtSkJ0rKy7jLgj5jJI3Rj8dBZhwh4Uh
UAbOfnZosa+rGXQwo+2s9hq1YBmD6JmPz8D44UBqIDSAZw8jNFGAXXB1S39Wgtn/
221isIajgunV411q6NKIgmQ/2wnOgSjo/h+ysVmd1SYeEeNDlEQZ196SIEBVnIHD
vYqbbRTRLuiW5a5ORL8ZXcvsup8vrCImkz2Bp8K13XoN6QvH5+Jg/a9DPYc5TetL
bH9TAwBGjlyiwJulVy5Bklu2oWEEGujGcjGLbdB7bSfy2YapBqheXk3RAYB1cadI
uAGQKmkl9oFupRj4MOURgV1khNoVDVT6XzF7BzIg/z+slXrhAyxnC1sFes+xVyps
ZAngUUM603B2VcOf3idTapIHp9NPc225vHRsb/WXSjg1QPJb+tgI6jGivsrfMA36
Ui/PO74nQwzgvoAW9+y8SOn1KrBwrCV4IJZc9BWGjiz02HLFjA95n250Xdi8vkyy
myOppy8CvTayQt6Yo7fEfKRpsGsD5e+d0DvEZDT4JfgBW1WnivNAAgiPum9c5FzU
513Bus0gLmy5BUgvZDYdJbdh1BIIP/yzEzgCbsvkOJc4kiXTdBecK6BJsPNcBcdl
lci8E/NtrgcZC0g39E1bVdnJL5p5uPlULYa39fMOFScvm2GB5OzyvM/QLvpHQU7X
QhFI2IHPUu+O7IlUD622eT5YvwIDCR8Va2TwUrWVA5tadUMUMjfG7Sarz8QMMPrS
8A68y8MhM0jIwc2T6WXFOPn+vnmEokL4IH2Ry/9KhwjVzNk/bnX7/Ou0AiPDAiGc
uJ8Ww9CPsnuAI4xYD7rDHwqbTPcUEaEWuOfvHX60EhCLThH88wfXI9gy52GZ9mIL
39MbLbLYVFuwpXuntc5GNv87Qafud7kRkhYYEXAQcfNe8TiyL7e0r8hzJFlOoqbw
v3BLSTWpAiS7QdHDV42Wznbyb0PbO1ZKVlwkvXHeyRfTlEtTgluSIwADMNVVv4C4
H2lrBgPDXAqJksfUebFcGUfSFDOs/Ego5f20EJwTxikU0YyAkpGYDfHrG2Nfwyr1
t8DXdRAof5LLFUC8ei4yH7VnLwajqSycU9YY3bNDlh9B1IsVNj+Vhu1D+YLMMiME
LRVKU22V9qz2H9MPR6PQ1tDmjiA91yQubRe/wfNbXL2tdWIZwFGfAONiWmVBZfVK
xfgUnzTNDVD8shunE7FDN+Bo4kDk/LCwEZIw4JVSwLUWJh49MY/HNqAIfjDtAPGv
N2D2nnO2TnbiOZhL5jnhdd5AfpCj++Oh7595NrocnZwQMxTrb7RGxkwjTLOYsQqu
vChUpw8QReJoSKyK/Kc5YaODzRIDMKWNP+nJqDjYRRKbZO6clFCW6HywSoWY0Vww
/MxQt1TEb7t3wxsLoodjhokHsKAzuddsFbxCX8/4X6G4qQ296uAPeI53ey+188WO
IoUZF9E5VVqGEPzPI9g6AYqynJ6to1D2EDaRV3dkaevVgiPWCNTVbXJMkEBJCsdi
srGec1axfOvYCXDCU1UoMW5yfeRiUG0035AfLMAC1UuGmFI0++jovPIrUTxDZx09
gLY7njCRK3zuEM4Cg1Q/k1qgzqHa6u4CqB44kHYaS4B+QjmD+39dN6lAIlqK/0uc
V8O7ttwhEwJjisKBYDiIm7Xhgzf6rfiZCwk60374RRH7d1Qh+/tFFFulBl6cWQY5
rlFERuitpM6lbS4Y41XBDbCqqgLYlPxe0JlXAstvZdOYHsuY5ilgnUbW4FLQzfH8
2/aNMi2uqtF3oLVMYLC0ii8vIVbT3IdfoHTjmHBSGPrbYmg0GCEwhlR0AVUZMyMe
x8eDrM9/ziqCyciU1uZWTy2GaK86WdItI7XNnapHyq8tVJ42OTPYhhQ7sgRBDVax
3PWMEdk2oKYAKypnDLvOano8+go9W40j9VSyyLIVITL5dyHO2nFyCWzK3GSVP87R
PxKLT920drBA5rulKQEGGNwPQhCFMEjbmDDZ+VLFL/Ora6ghQ8ZPXQmNtON7cXyO
svbUwspsS3MstM6aW95MwEFWJadVUy6I6aIjIj5cKAnNzE0Y1ZP1sDtkY/hq9GWA
CnrbZy2OYG9aLOMSkdDCdTJ//UtDkQSDdFrZNIHiDJ/dfti8u92D8KzxyUnE/j1p
u7WG55H1vMd9e5+QxqNcw4tFn/yb0EVfy6cxARJqsuJU/PEueq59bkAhJvrBJwnt
0Ozzqy1yIvbu+ruPgXLVszWpI9CQaE87vYvry+eAMqhUBJ+EpctUtj9Ii4K1OqBO
FH5Kbo1XyCAkOWeMF/OGWwyQHDDw2tnrsK41i98GbXO51lg2OmfWTExwGSqZEAGh
UFBKElRAkSCyqdLHJtptp5+Y/T3+CrMoggbqwX0gBOO9Cd9Goijp6PNbmJFseEsW
vnBYv+Ap1HSo9hLDXmTcfOTHdAVtm7mb4OLo2K8OMyOoasl/ETyfhMj2ufQGj8HJ
07z81ylr3rdWaM7+jUZ9NgU6hIqNFT35BAM5cBC6hw8GPHbj1FSjrY5M4hjPbp6w
3I3EU3ra5zJ1IWU5J0N31NGJlkSsX1RR1IsuzjKx9tS/PU3KEMDp0Xh4+AzJ8Ju2
RTwjBANLDvmZwJA3F4ThluCszMp7SWHDVcQwZyK9uU0vCQaovIl6F16GExZhmff+
v6gqhA07DX7WO/La2mK12CRgw4DvW6XQZenuB9Fhkf0qHa3lAc1T8rWutpV0dB3I
q2CVdhWwTcv5ddPfDEF7nkSLA/jZg7tc/PzE7KFKdyVKLPe1uTphDG098omHbI8h
lXjtM1NX9378SGNeeUeWxLHxRwyA12UmA7EPIDy2Nd6sW6XOJMQstVynEo2YWrrf
0ztZl5vzFjN6xZ+AicL2b/G1jeEM2Y6fFGMBil3YRklowgzBaojBkqfjANCDahd7
tIrSeztU5KM7hxiqXrkFeiWCgI+l1AexkLgeX0MzAGEC01Hlr0UqTu+O+YZLBTEw
Vq/yqEHnCV28TRybpgrTRIJV8FiRCtUI3ts019df3WW2qmPqswMOrHMhndLSupGF
3fNp6iawT0sxNyNqmR6pSmGf2v201kj46axk8D0pMT5soQn24g0aUdR9pFmjrH1F
kA4D71EoKq+Vod3owJSslz/A2tSYobCniFjq7Wp9Qruccw8T31O2x9Q3+KPNfmgW
xsX4ti6+bDKKjZrvZjnC4r6IzFaOlwnoqIFhn34gj8K7+/Vm+hb4PrQpBJHzLOuJ
txqq090fElepskNCk7mG2iKaPTRhHGvAqB0zJZBmvVKkFIxuzo9xBLZIpMEIEo4O
mP0ggrWNNVv1UcD462zYqxx0DI8Y6gruOTFfsEUhxJLQ9Tt9S2nVzHYk8Vk6m37T
bdR/sBUBZ+6WG34+hIymZnTYD4oeWwthcsKz8sL07YbyZVixpZREmtcfJA4WRpC8
w4HgB+PHlM+X5sGJSZN/YK+jjGDA3RjTtzt+MZ5V8gvgcqAp4PljFE9iXsG2OPjz
UQ355bCOcWWMmYkko5ftF5lEDIcDotx1xfu9fGZ+gUMxvn77QKpMhuAlrQW8Oal2
3Sj8gP/v5RXk0I8+EDV+lXY4P0AM3aMLh4Dy3jco5cyH9p38R0sjNJpPL8K7J1wN
xur4coPRY7/DVcfdcA44xTNfRObB7KTY8wEOn/wATP/nPFYb1vh+yjZpCm4HlBg+
mhdZ/Jun7hn/3wTKYXr5qbSc6uw5jat9Q6XxgpFY9uhX4Ofsu6LxnJZFCmfP/B/B
H8cBXIRliFxLl9F7u7F6O+OT7dmppa6sWmVTvgFT71BdtPdVc4KV15ZnSRlnMDbx
izJtdbAUP751EswlFr9AJqP/XyNAcPlMatFp9VSRsGR6H+OYn1b2qpwKSeR3dx0t
ipiguXl/T3OWSL6opO/qm18wBps6jBMR9PeONZksvOSNiurCWUz1OHREf4bDEoXL
jl0HBgSU/1rndFIwddmUx3VZcntCoaMZA+8lz5sciwcyma/gWWRdsS/iXeRH+L1Z
pSHhrek/9STlFOPUD75MwebTjvsw/2fLmH/Rz1CWTl2jN3wELAcVqf+jTtT8ny5e
HV7xdwGs47F8HXNoooRsOPPucG8iPMtjlM5b0cjylzpkIxvfTgiUzoFRBatDl+vx
+QWwAYdRBpiRB5xJNgwv/jAqiS8OGcfnj9tbJYk3I2IBH9Wzq6Oe7qslQjNfXy9I
03UBsoocjajrV6Bmpj1FfURCK2uNvseLGGrFDYUPqHs+9ASPS1dcgv3zydUjENx5
lpK4SfE+xCJ+EYfjXtWRbUBPO84VRFDoluhsPSixSosITb1f5ETHns+d8NDcmoIv
co6HYbMndj7QS7Ks1O0NgFpAa+XweV9C4UkeonMUJuIASHn/U1cI1fKSQJb0+qNP
85sLfnB55P5oVSMwjjwQIrfAJxUn8Q2qu7MxQ3o7qsr3SNjjMhDWh6NNW1WNazzZ
wbCXGtGsKtOBpCz6PS5A3+wEyustudIVRKFPVO6TddEWk/z0LuHFZO8epix/3tdT
9BQc7Ox3K82XtAiHkdN3BbKW3j+/2Cyoz6tyrayFWFXlp8EkMq191y0WxjFFAcRh
dPYT+rMztI2Idg90i6Ojn4zb1xJa8YbCGmhEzqf8ujsg2ZPwnFO8PCPucoYk39mk
Ljx8hJjFVLFk9AZF8z/zwA9kAFKWRfNY2u1Mr7kK7ZjwP5450Qpglq4Xnc5GYW02
NvR1QYtkh7HrW48vkitn6I9mU1vsGmCw6wa+JazuzvL4scpUIeaLGaTxSgsZnt3h
l65aD4rN1wh1T82PRg3Zg4KEpHDXqALJ81ajlarf6LRgcvgaMUNdyNdfX8HXTsP8
nE6g6bhR+CaHKvtMcf8PW6fgREJmAnhsLDnw0oWachsAOQmEC19ecdi5yQODg2Dk
Io7IseCwf8vNvztGAyvwKoyOuzoqqeqlPyBIVpxojmm70/dnnzI6RPWie5rVYPGU
OqXoQ6UgN3GXwMUIPGgIL8RjB0dvhLa6lRftSywjafcLQIGIK4/mCX+Ge+6mndY9
06SHxVK94BO7YwN9Msx7+ItTRoZ06qU9weiZLe3T8t/NTE5wghSes5qgLe5CE6LG
1QJQo3FqwdbwQAM0S9wI77p8GbLdA8wG5HogKz875nzth85+buJlXHT0dD7ecLKQ
Hb6N3fziTN5OkWIdJwEw7BOWKRzqeSpc0CsJlbgpSZ0fS+dnZivEh4YPjWbbVsEP
UO3itAGDRWKGLjZbXRlRsdZT1g6qiBShfGQ6J7oQgA7hvU624PXP3iwVYOncjw8v
k17+j1oolnJq34Hx8/ojnsUFvMkWc9AFw4//9+7bEszTmaMyclUZGMn6LSf7dUuh
y/cmU41ezo3plXizAfQVTsnnYvo9gUAQkXqCgZiaCAtQ81A6QBmZmIpnA4vexwmX
DlkVb82bg5G7D0hBdgRuXfkK2F813CL1KsMzoqeX1HC/Z2MPKQfj0i05hnGh52W7
s7Vt5kv5ZHml6NoU4GYGi+jFpl2K52Rd/kLLh/1Or8d68P7RyhY2T0s2NQf0F8v6
JUCn7Cr/zOH3Zbg2f9u/WmQgsl2cRnWSnsB33TX2Qi8hPNiqByb0LWuenPj3a7SW
W7HEkmPrebwBul5idFe1Pd4DF3PKMrWwGAxNp5vuueJPOTf2UjGs+CrgJbtUXI6+
+g2XJgnkDjyDcUM4mutWfqzcB+rQYjyRacXAB/8Fx4sDR+DubpVS9nnU92KuPrH4
RfnEtIWpFkFw07Or5uFWPobG8gvqZQeqNrzOvlwzr2yVryw9JTevaJWNbklO/HyH
8ok4p8/vZYmQ7MDd+URTECs47NrXrLGXSGjiOTvosYQ6MOtcTO8GcWzYpTAo3D+W
kdXc2N0VvjGGscbOtF/nsJ+1hNB2smakYYSTygjd/KUrgRYYw9FoW5K5d+TcCPo8
c6AeQHt1nHv1lCUgtYuLG98H2aDzGcW75JVf/wPWiKxhE/fC85gxx03krLCs+kLV
llPFmXcop3eSEYqS3/Xnc5LKl+hIreUWiBjBNMrnKjMtUkMLc/yS0U8xzmdxv3Sh
63xZrdQdH68NBWovyHl2yh+71um8jxp7kwaEb7zdj0Is0am19sJEXxwPK5oMim7D
piz5W4YvjNv5IGfG1PLX8MhKnPniQFFWNHEyK4YyZtr3LYPFu0ghAPL4TkNTQFJH
/M+Hc9Jlk7b6FFAvxqAledKMuHNHwM8AqXkM1llgsF7Vv8oJZIOurPQhrwzz8zYm
ZFmQI/zvGFVgltoxULhstoy6JW3cnwYLHkm2yrrzsMwFqLe2bwJpVlXY10Z5mBZf
4ntTDoI6SXOkXMGUpn8dSe0PjT7IQ0Lz9SDh9/KxBQ0ZNxfe7lcsMxNu7Fbun9ce
4U9OMdkg5noYQyNACl/HqpMZz7RaPFscXDCjoy0ajDkIzoZAIkvtoqX8UklpCp13
XNUAv228VXBX81RDkIA7HO8wgqFyxaeRJ9+Ke4dNHqkyCIJ7dXi5MT9n/0KRfwfw
wYMgpgwmZ4/9cleF8+VnmGE6l4jAr+aPsxsQNRTqAgRI11IU7Cvfv/a5rqqYzBwN
vwTlTO1vM6aRBsF57faPJAdjUj20ElEg5jy6DPCbzDcSF4VUgMUDe3NAngtrc+JD
4BshSFwB2w3mXUtbtCQ0uRmngyQkQ+TO8F2W1fbPBfe/x50mHTVkKUWB8+d635+S
27b3pqmcpBdw6D6HwJ4knYKugAQUmy1pLpigYqJo3RIWEYQfhmqMQgdoJXOhWb7z
Insk7ONYe4GFLCks7O67/bBRGUrNRueUmS0T9YM5i96EVBq+nYhAr51pweEGjIDc
Lbgyt+F4hHHxxwGzep55mrDp7l1I7E/f42hZkkGJuzHl7ddPcrmuabSRmWouZzk2
S9Gzl24DUwICpoXugmMrjAzgAJWto0ZxmFji0UPaOW0o/a/Y0p4gzVeJ855sbIKW
2+zFQRC/CFjwiyy0kwG7Sz3EdVWaGp+C4D6/V73XPPjmi6TlQfIjQ6P/ER1OqhQ5
H/CgnKRTj+CXz32GXrPo5eOpdPVRL1wbRh9QuEWIIWt6ty6VXJw2Tur7r8BWQ8gk
K9PtI9wZfPoZFGfNBOcPjplREmx5JSRAi0vIWcyXmCLr3ke5hzHSaCcWmyH3Oq5n
uBhmJxrKcxwHxerYEr4etvKjCUm2ngoO+h89T0klx/m4L8BhlCwGnDR5gYaT3zSQ
pfy626l79OPdG4t6sMjITlTXAQYSYK8jiXfC7HBT9h7toJOMDQlr3xrDT9x/bOHC
idAjn+D/1m4tSvD6DADzd1Khh38jJ87M5GWCFcJIzNCem1DMFoGcUdxxzfH70jVb
PZ5P83hTzzervx7X43LFXtf7L6No3Msoh3d7TXTukezP2e73DA03sV5YmaozaYvr
8QU482umWHvPxDOziuuKQ5QnCjy7H6DWae9hI+L/IxwYxchS2/oWbYwwJGWE8B97
RXAqEQPuVh4ErRWpzqowOuDuWekY2RljEx3KTzo9OO7w8rFRevUaygCdJaEcynGX
lvCFBZrZUlXhBY7pgQUfrjVVYgVVhoYC16H5ScNC9e3VD9D0NYX8lfzgtlUBCrXz
rdQgflTeGx671p6nCtRWIpzO4UU5xgjS8X6OgK56NxYWYGf3y1RbH5Mf4eZwM7kg
Cj5TO2/4ZbRWDC46+glmA9A9kdag0Ggw3Aw17H5Tt6yb7iDaHNoiqugxcyE005wE
9kOMn3od79wDQ1tb26L4t6u2b2gDjwMCXtCINRux3omJc2HXaX9GapeVTn/eAG4q
fcz1nKSB3w1IcJvrsHsJpqOcKtvZFWAN5q/H5qBjpU3wO3fNG6DneaN07TiNgWuU
3IDnRDeMOkGeQ6tIKI+z6G10KDHxIIg7qUmOqzlq2SCckEuzlFV2ALPTMSe+HKvf
weLH9JQUudqgjZ7R22oAdPy8JdXfhAfAfdq4Vnf7squTKLbQyoPqnJL5NOtqDnJw
nhJ5+DpJ8pZ0c1EisvdnE+/mXSGUDqxTK1IBOvlJaEmCcmyEZPp1HakFziPS3WKJ
SJJXU66JjUK6PdFcADXv+OASshXQpFfQHzfjrKeJhw+rgvfldlmwSKyU6r930Npz
cPnLc+oOvRY8yxGt1kfOKRHmwGpeGyZ9p+sveUYuRZy8kOx8PuSKFtUiFWK6wjv7
wl1CgWJmBw3FbINQBcV7hATewzsv82iVWRVEsVBL/qTRUEDDZ8pRPsNyzxG59YQP
wr/FHs643eX/QO1reRnOCMjdQR2cnNYOJP8O0oWOhuah+6GJ3i/WFvIHwIETTSbA
y+CAj5WixQX+zSZSJtHkwoF9g/sN3zb6Een23ihpxtMjDJXa5dtGukQ5Zv77v/qv
1iDUEV6UjdQaEOdsUEiC9GqeNVq/4LuR3vOhnYv1zmN3Pora+jab0zei8Wysziet
RvFj9D/clNvE+egxQ83LBkZxtP71jYWrKBbI3lGtw7xZpxI2wMfhCxI6bsbFB5RQ
e5E7gj6Bcto+OBXuqYXh8Xhcm1c6M1UXmzPV6JChNFPIWSbclJUZhbDCGUrNbuJ1
DjctUGEdEcUfdZ88Efpqmb+uDoi7Xpee3K4dtNR+LqZZDq8+0xelJgBRSPenaVLs
czm8npeeZZ5BzYqYVoJ487R8wuTF3x0gvImXUtRfxJqSGRYoOaS0trjHNc92x+gl
UK2zuoBIRSEztsKHKR59LsHxCF9308NDEZ5RYVuozmcss4GB2QdsafB/WYc+1gxP
RvaKLmlY8HSb/xod9pKb9Ezhq+gzhBA3hp6dVbok45U1dqVblHWoyJm+0InPvcj8
4OVjsaxw+Qt5rDnS50dut9p+rIlwjzqkCElcGa+RXxiPuHt0/iFXwJYKLo/75AwP
7KxvZmTZUKknOk8JBhpNwxvcUvxTDwt+0QgDOOHqkqiucGXFKcepU+bt6gxEOCtl
qh27ktg2hVmVacWGbgkicqVCcwN7l3OWBeZTZbheK3kbNFb6kkEqK+8k0v2H8f/t
DoXRRA4ycHmWUKlLZGcMM5TuLmNFmORg0iANQhmjFZIklMIl08ZQwqFjygSTWe52
s/sE5q7pUPXsuzLeQkdi5YhFiXt/WOst44wTGVNYLCtt9T5Gtk/iWl5M4x4BvYSj
MZRRcKwZMu+o2wT6vd6+G/4UkxgJBn31bqovUyLOWu+mqtIBUef1UTXaIJrCYF6y
YUJzOVTUrPZmx/2sXkz1gVSA/sA3h2CNiC68BZ6XZgvLqsdCki731sOyqt9H1VJB
h+lU8eWWdt8rERHYfDznTSwChVcyG6PFYy5wdArJ9E80X5Eb9WenttQceHCPvpsb
C46JlsURdN+8EqSglq2QGXSyfd8vsuqpfPvSPhmHJN0PIDnqH0vCeNNom1nt+jT1
Z26ufW18KRCUv2loWzl5dwBm+z0/9ThAOvATBzBVRresqBdjr3VB2UuMpbhk1/W6
kJOrSWunAdlFZ96Iv2SKS6uCjW/ZnXg30yREYE/LIvoePabGGLhqNnS6tWEi2+AU
I3zZNuOdph1oUeAQwgZu/Ro67/bAHWzbARnSJ4WdO/faWogI/rtm1bIkDYghYf9g
GYbXyroQeWAkB3Px58Hm/hSbPtAevzwLJWXV3DQzDcBXygoXDOKTJ/hVh4EtmLRD
aGDj8BoxXWvrBo+HZzCh4OVC3iqWK9ULCeTaADNDK0kfN7AUMn+oEM8qRDEslW9D
XBVpbaRPUb/PNKirPaJlEOKQ+82RV+dr3XKH1vgilg7CJOWrKCEd4hWs1AgnTrbr
bdkScBSljB8axNjKRVP8oasR864LDpW+NYBW8DZjJoxg6b9RGqld4Vf//nD+0rNw
pL8KOI5x49kP5PhUsZ72tUATsAvwdoCQk5qonHEuVp3S8H8/+mfvPylhOHSX+wHk
Jt/D3u/NAAxKJge/+yNKb+NLrACBt0N25rRiYr/NXxkmE3Jaz4xPLvAKypsxsgUI
J+rZ54Try0gYKlD1I6dpXpf3PJ5daovYLsboJXjize2PaIUqZAAS9jRScEnzZMRw
N8azaOmdwgxylm3BIYs+C/xIz5bG0xLukLFBubq5WKD64Y+mpWrBauRjRcTbIcYE
fm1BzMZvDdukWI12mvXVfbT3xcV8OsoIeqqtpzKNifvSuGXTdzoKz5fZWaEqKIQL
mwZbQJNHAUz2wELd3Eq6a+MR2yrieRasq2QyiMNn2r2js9XHR+VbJtuvcxdFVC8R
KVykHupjnim6jVHXDY0Yitvcnh4vo779DfAS9AzaAwFJKJiRT9VUr9mxWkqyCkXL
tHtJPgFXi1iLwDghcXj8sKMhttip/RwMI328WqLtaFEUrJT7SfJFlVJBQGizp8/b
NgYlKKKkUwWFsRQBRPXtOGnXm4I7W1b8pOkJnkwYZf2YApSChaY+EXibCGMxQhgb
2FXrd/QIelFh8EsRCLJ0bepNPE+PTptDIx8L4BotPB3w7MKzrvX7ZOhATNW3KVIn
wRbvnOKmc/f/5Gz/tISDiJEpGyCp0W6WPajtW/hkI+26/aB76/00wZVCtg1vsbgU
C/RuvVAmKbwnkKKY0cNWJPVyIzaI9RQjFG8WbW3iNaXzujL8zHRkBRCqF7G06c+0
t0ipBPuWZuTnG0pN2iEfpqTWtn6TEED2tkh0VTvm6BV9KXwh1Zmck9VftezEqr7/
n5uVSJjedGBHnoFSwaXWrDCPTWfA3+5r+N9Kgq1aB2JUnwOyNoOMQm4K0qsSHt3d
I1rp+BRMX0DnE6zD0aOhiy1Wa8WD65v5UW8xj8INGXiLFgiQYgLcnkqCnM4yk37a
dJAX0l7o2ph+arDeOyVqbC1IdB16DOtghPVd6pSzgeoWbI9I7eDpj4K4rgh1wzA/
b9jv3lbPbvd2pO7N1GK0Q1BjfAhljhPknKmayufzym0k0elwo+kyJ2x1moS7fxr6
yW2canCscdZaJjGPVVqK/HcAA405MyARShp6T7qrn9FNiLVV8lOW49ngDkTFVGa7
O/ApSH4mpse8pkC2p/9P5z4vY+Kzp5VdoB5C+YOvzGEpB8ZwUXHqRWHqi8VPSxfc
ZzzNJYOv9UBIhaSakml3c7CRmEvrzjtaKrrDJ3fvvYoWy20xetuCNSie+/NHKY7j
pUqo5J/AVX9u8tBpcoql4+V3VUIF1Z0vl/k42GV54SONS3dhkXE6QrY7+BZRLkmZ
+O3cH0TTMkYXUiIMC3X752/mRG8YR4uhRbNZ/ELlfsDYicYtIMh1zCrFqAfkG0VF
liHbSk9Ehl9+Q6vGVx/4FIsKM7KH2WYVBI+Y4UgZ/+gLkRxf0moUDezjRianpP59
3jI97cQQCsWl+Tuze3Xqjjw9ANnsKAtIWJZa46rFa6ZDzIGrIEvSpBSL6G6kAXge
DD6ivy/tGy9Osv4dslSysrCfcAKvb0+ZPMZHkDTRrbcU61pF8pAZu37xY1fJCASn
WoLzXM+lbM0If1KMfz/xoy1ToH5lF8EflphyVcvPbZlEveRHxAozVhutDk5yPQR9
/df/0GuC6ezhmCX44morCgqsX/8vnqiUXHJGGazga7tXxdL30gqxGhsdYCXURm68
/9h7Ffj082H2kO15EcDWt/WZwGIuNhDEu+FoIOAP5rVyWMgAS/Pi3B8cKqJTX0qW
g3GYzRz4FzYXBKUYyhQZqe3hcwzMctDrpNK700KMNAkfDvR46xPOpi6qMshoMC2+
pgLPjoFUcGEpbr4S5YPIloPGukMvbKwZoQg4dn6FQBl8K1iUj1NtTbB9pF6Dyhow
HJ8raGo0oUEDT9EenIT3ZwYKVwE03rLTlwB84Ny0yTeq8NMBjxxU4mhxIP9UzUp9
eYvYPqaYDP7KPbqMUlR41gAY0dEXuVMcdlZFXbm60M4PNVxQAsCKv8+J7/vdAYLW
U3CIlr4iNM/gtII5fFlx2tsct1fZgULFUhOnMjjXcIEX/ZMMp3ybg24uAuGe6E3h
k5mZ+yEB9qAhvHwNPqDVWeQL6jrR4ix8lJzLM5wTQnX5L4X6oqsCaIs9tL7e2oO3
AwaCZO+3L2mPDopTnfzLx5RhUnEh0d9LunSqnve/+Q1mm2p0uP4MqqBfh2PXwBQD
G+ZQeAW84ePYJfg6k3i5+uQBso9WEZWYfETd4++w0SHeusrHFPadxrp9byLv4hyx
Zs7SOLKxXc73Q+wPu+uQCyFkRIaW7pBmapFf6iVQcgWHw+9nP658boxZudrrI0nm
63ox6MkBTRbmBG/4WCkcT6k6EtUqU1SQqyv9tEhYZHjR3PQAxBgLbIVO9Pq2lwXs
/0w0lhHsXbhycapi5FaeqrtX/qWhxMHy3+vt7YumIZXz1NDTTkpKUlAn6lT1/20Z
kqDfDHMTu/uF+7BR2DTmRgrrUGQ8SKDHhg8FHNRdVAXyMz2LzTofkelnMqZcQdcj
uVlpCOfrWPEzs6bge7qM8Ly5j3vktIJlmJizv7HMDz7JuULyrAtV2YKj3eCI1Dne
tP2Ef5sw/5Iix3VJ1An/LJeZtbXoXmtnaBQj3QZlzGy2t+4KqOh0sTT5FAYnBONP
axYIYtPmsx9OLWGIK+urGQ3X0EvfASQQGr1ANXWaCgWzVOe/WXyqGiaQ8/YwRN4X
rK6ATCKFmyoq4NcQ//zvPqPSyno55GptY4I5b6aGE5CYGYQO7/8PGBZPzN+Xnzzf
i3Tw/t9Q/uFEirR8DYWH8HNrDx4FhvuwV1/Fcdx706zHJcPmsphhj3LA9oRQrHqx
YnQE60sb8Fn0ivtKDlZcVoATqP65Y1BHmDNTrVlES6OGw+KIoENP0qMuYWh6tQdK
8np1U3+/yIic5WdQnvJxh88cCdpPmQBZfAA+TSeyY/3wF2ljuyi+EYhV9//sYMLH
yqPWpS586tbAP31D8lxqjEU/xHUCJLRXv32MdI6MceMtT9Lyc3TNrSgyuMyUZiNp
Z+N6Kfc8NqginfL+wNnUEYJBpPU/L14ynEaMAnJLfirR/Wm57OP9oTOMn83yZktK
GXkC/HfweYPJrHKaNbsbU/CLZuNsZ7BTmOkIoy3ovs/ZrG2djJYkwk1iADQYJbJ6
2vUMG0NAH/9ge0NBYfWzI6HH2P9NkHdkjkQxMqY1MGaye/KF7aeqiEKe1Zg5GX/k
VhVITZmIbnYVqBWVn/NlauFnTi/f9KlCmyqiV1k1a7x9bBKqjSWgYnjJkvnFba1U
zIwUfDiVxGFy4Df9cBhcJxryKcbCL6gf4A+raZw6F1cpWkGRFEQsGwuF0LLXDtN5
oFStVUZWJdyghOr7SlaGOD1kQQMink5lxXWqSE4LtPfPeyamg6S4Q7tkgUpFWqF6
NtaGpZf4EUiTagDI+D5sSuy0bSlKU38e1OZtfnJ+IKVvQUCjIC23lUDoaZPOEY9z
0KT/DbQZO0gpTqNbbfbpTsH6E+jMtgYrm5RdZggYV5qdp340OwTak6R3mIlg03IJ
J6Vr1JcGVOFGtLjkUU7dsT2RbNGOD/jptm72odkEPHdpnzOJNwgbL0Z711rhlspd
FooDOZszmj160GkvdxoXv/gRrcDPaMzooH3lXfZboMRVyzT796ICeHfElg9otIQ2
1pRV2dLUmDo1w+hWLXjqlXYluhtHiSYYavINT8bQKkQSY7kyH/Jp3eVvUgvcF6R2
X+6bVOkuZvt/6yBWsGukrfSysU7OI56AwwlAhMirrn426UVu/ySI0oHv9ry5D/YF
/Pbu600SPqvONzTVlha3xNKKyEZqUnAnQXYyDIqRiFvYAsKQqnVXk8yCC1lS8lT+
e314zNyfIVw48pbrml99yJIcTWVyTmpEsjF1LgUT5AD7ICBe3E5zc7nxGVmqvVAc
nSITNXGTwrUbEn0tYRxKJ7BjdXXPz86ZOPuyXl0UQ8Egtr15zkUuj56denUb7h7I
Nn8GHxAmElVE6YsUWEtCxdu4i6zSrLqaxV9+5kADzDxdPQK+sDIpVZ2DeO6b5CuB
8P8L5PBwWcDhvAucBoffEX3Lq2yypr7OiVEjnkd7lIm6kT4B0uqOEp/05Mxxe0QP
lvuBl81biJpNxXxBuTAuqCCtN81OkaKWaACX2uhz3v0zV0WFAnMdtgeTjuwbT+23
pwX3DZpWwbMEkH0llLThT/2kDnW9M8LMlhr2JjIFG4is1+Fo34Qmxdx2gkgXStLB
6EQxtTxh3AmLlKh4LIKOwGGnHijpNjxIP7rTeAhV2CZ6je5qj+RrBRs9lvsUtPby
nQtq8Edj2jlS0jidT6C/0NwvxoxU8+nBvpWyEaKbG1le470tnWeOX5BiVWVtRaPp
tG1P9Q7kZpKIFDMdg4EUP12VLNKLkMoPiGJANS1PrOh+JoHhwhcSSJpAq5WHGam7
8xjKvZifreC0QauB8jPlOwDDq+oB44IxCAgFDD25K2Qqo2YddDz8Vjftj05JonKT
Y4rn+OYNIKlvsjbhqRAZSmqPOsjGpFM+q5VL4EZVhKUSVNr6f4CEWZcCJivBhynH
gm3Kol0B2YgigU1MjJEIVXh5DoDqPmEg1yD5suuDjNy4zurv02V7TyIQZg9TOpWd
FeO4GgfeJAUZ4reO6Rr8Be5hYhsU+csPekVkxlFyHEncuBWIeXquQDTv4NdYmdwK
vvUw+rRDXlyCL5aKEgfVbTtM/rPSpjRDrewfy8h4NnmMbinjKMW0U9Bqnw1f0aBf
vwK3iU2FmB0Bd9xhW7mdcN5NLnaFAcaV3p3Z5DX0gZm/DGnmpWG1Ab5Q2Kpypkj8
7TakFj0zURMqgcRJN1fzIDWFrrLYhmEqUqt37s7NJd0uxGY1rsd+A8GIjy3h8ewN
afGjg0HfMyrusHzSNdMypkdZJiSomqmQyU+1XJiWHC87BT9rvN3eigmGGq9XtHwT
K2W13ITjJzvV8KnEGci+52K+LyXtd5aGZfalLQWgMIfOdI8ZFqhL19W6m4b92rem
rTWl+JaGW8cpRbDbhusvw70RwvbLqNVVkfhFmAx5fxSBL7RiET1Kdy6mpQO1Ks5z
vjURBWnGKQ8bcDOykEKaCGtlUtOdQI/CfGVkkFWb8cDIxXcg81K7S/z0FcdHZ+S8
l8KNubyDpNw5hG8rnfPxS65BuUDdU+hHEP8d0+NHbEmnF5dfchFv+dmK+p0XQI4S
fzIr9UKVraGzq+9WwUQGEQyUmxzm7PncPgskPnpduOG0QwnP1rGaaX3HRl2X5OZl
6HOHS626AtmBiWFpHOg7S5VPZtD7z/mf9N5U1rI83+mPr2/geuU2e+pqa+n38ta7
L9EeXLryXKfVHGq//oFlb0w5C2MFTbmCUqlAx/EDdRkUIDixno9aAH08XdrKV/ug
zCzSR6PzjCaL/BUp3OIwPBRbAo5gkasN6IwQI/xcB61+dgBXsB3ZLYQpgt6FceBj
2WLLFwKdZqeQeosgw6hg+2SW/IRGfC/on/C6SnIqMgbuHWt1J/Hu5CoCljhixkur
FrZoceKLucf65/OI1EFeVkuSb/vLtv0yvY+ThmJE8RzxXGemJqQiZo4swaabusQ2
X0feROXThX2gq+VGApNtJQ7ba5EFSTXt+0cIDb5TYVQs2WlU6clYcrmrztWEciZD
ISh1xpWavugptq47zDCd1SWfDKcL/7o629dFnLF1WXRir+PzIW70uqnT+VrSVtkA
/r/nO74rZRJI9tzy/po5azdjI0mFBSs5F6l1FhlY4ExUb2baR+6m+tqEWy+4sQu4
ZUMXk0OAmsZF9mXtR9gAF/KvnyGr0RiwYb4DapGD6/PoQK7do6PNutjDT0Xd8Skg
HOfDHsgMJ+yxgxMBeP44WTxDQVTu/6SqnAG1bS8lwku9mzmAxIr5x+D1lfZMnz8D
P8Br0uVEIpUkH3QQqo7ZypcXj3fcLVoPuCvyrQuHI/ppzSNRTG6PgUBAmpLUvtLv
JxyGHNgdiUsNCjU7bWtZRv03ukG39Vh1UwYAJkNyBlkWcEKNMg36zmgqYEX6eCbj
UBVyl047foIpDH0pXhbz6q97yPvZOHxhvky6sIOonBjuLEEmBljT/RKiyXxkwyGu
PXD64UrkhrTWt1CENB9Zpg+96dtQ3CZCxx4ZbvjueRMNrN+JzqbbZgaGhmWwbmCz
JIKIsef2/3FfL9i+Ax3eI9t0I99XRcxcVJxf0Pbpp3xpkqWdqyHqAte79yDIW6FO
GiaD6af4hBNb4/jZMjD+eqa8AAZ+mGdZvaNKzCtl0c9YxWDVuhQmPscQSQ51w0Ro
H2mUtpPxIYVJy7mHUDsfpLgMwIM6EOh3oojx2723E9l9kTvLx1W60XE32I+FlMLl
zgGhCO7qP4Q7ERlJzmcLPGGoqrHMnWJUCn0Kt4otw1S3hVYu6x7ABt7Gz93JwEg8
Qf9Yhb3Eej6SiDVbPJMj0N2GZOdjot9Wl4lDR3hrIpUeuszYethDY3xW1fiZKrHr
78Nk8LJIAXE/Agmh6cXjhDTCS5EKqxJ+JaRtI1lQyywHPMvO4gmRNLDhCRlxyN0H
L6QnGzbseVFupZDmGOtJ5D/oJJVvErR9LR0y/YcalI7oL1zlCQHYZa84MVTm6LAv
NqUchDV6Dpxm5xNO2a+DHoCAXrYxdIEIw63EodxlZCi/JSEzP4C/q2DoetJzuspP
arEbkTc4DXfTyD4eBv9DZqthIOsr3TzUI6guCLQe7bAXHwhOmLbl4hm7w3QLUR0d
+DbJEJZ0xLSFeEhnTApF6C6dLAuzFqyHqD5zWIu6/pevFc0vR/i/kniMxFaYqpRu
V1dP9PSZCLArKIb9BH37RZ46zDtIpfrash6rmMJcGoy2jhzKrQh2uj5MTJuMcriJ
R13YB+eIgdGackdi+hu799q1Ak3eqZTbzbfm07GyxbDk6yWGxRTakm4fUEY6SW+S
QGmhI5UGbhwoh02a04EHLfs67BIqlpN1wchkKtZyrd4DnYUb6Z5ENtNv/zhfwdFz
+Cuw10g54T3rf5TjbdfsCkXkMmNIhe0Qys5bQ/T40r5zR0IrRfSOMjQtE6NseOgN
aILfi9/pT7ZSl66r+ACXhhug1Zb710z0OoRAT7957bicHMWfYt5DDwRS5MnDRiRX
yf0hu3PXWIq3erhyn4D/FjFRPXtlThSrkJTqiT9OMx+Y5yPyf2XKdGs7ohie0OHz
30kR+WxUnhXVeDBy9nLilzRaXBVtA9AGJE+KlyKyvqxNJODhZG8qsWM77rhXxGdj
iSyEDB+w+qeLYvQ4Q4w//0GErFvRBHoCd9wUmSsjXvl1bMb3vjujpT5tJeTFrXga
mHxsUe/cQkg1wEPcXIamX4DWoU2JgB55Kg+VUF9pCtxim1/yaRF/QbSO/eKM7uIs
C+MHwxV+ShNX4ivFHcHE24N6inN/YYE9IdDFdL3UJF1jmMl3Wyofi0rGzEs5Vezj
2pcZjv+i0Wd7B4UcKs80Zk1olwz2dFXxRZMgVPtY5VaxKBLQnnxgJcDBJw+ayHp6
5XVqghMPEehubVSOJH3hdNNE64MhqfTQ8h1XT4WI8+5U5XSrqiZ6alwpzLQKZ6Zo
/H/uF4zySqw+9a8ExOlEmlip/nUEkoojPdm0V4TRwh3R2RiH2Ex1kM8d9Mk+aFbX
XMB5gsDO/QpN4/Q5UnKr4EkV4HL03w7N/9ckMfZMn3a3BfViotxLtSUujNaItGe9
ZJnBXgdH5gR6SfbAMuem2Xr5pf79+1eee3y4fxEKBZ2nHCTjCJgG+Lqi6MdfMeXv
0o7fytEJeZsHv34JVATI0o2I45TyIHuvLJUtXuPNOeiXrI6chaMMyRwLNY/yD2uh
eb5tT9KCWwoeJHkeLpZKnd9PZbYP4idda++YvwJ2IZRYwHDmvhkEbgR2mjHhD+SN
/zkgywQhr8ibR+kcpjV6IzyBrl5B3wkpNRnmf234SKZRIo8DW34HqUuYeQzrTsNP
7tJumJb7nZz1+3wAMLpwLA3oZ+tpGC7Fu+Azq5c9KhmJQQesedVLeUzGaAET1xKH
K0gxLZwXeQ2YwfeCPCj9zuDyIgwlOYlpwFjey0J9c7cihYnzqVE9mfSetXimbcZE
o0dWqu6+vfjx8y5ahFOzjHzg71ZROLcKPsoZXrvDUj3a+D0fGfPyynaizr4WIYC6
F5KANVLxdbwZmqg99xj2eqwr4Rbj8tovZYSnHVIVQWmAaQt2q72Ml6P1J/pOlvoR
d2/psc0OQuQpqIiGuDAboVK82QhLlSOXo7pWgnJH3ZJi7YRb7YmJlLZMflyHmfwu
U9I2gljzWYd03dHzf1ljZ3Bx9VhVe45BVN0/fG3EOnhmFX2E+ZLbcRe9ADTuehGL
8GihgcUAO7LJnf0jqHQSsaiB/30eeoSLCkY8FAx1TtgndLTv470sqKNEfp/BBYXF
BqNsc0a3rMugOfq1pkZOPmPCri8TGNhhJMGyBgPLli+OWN7tNVRTMsTAJEGUHV/x
DaZRpZylgvSFoaqKTWbBJRlDrMHJfIFEJyWcO+0R9mb+HPhagZrgwHTKzpACsvuW
AJfuRVT01XN+/vHC/sUUypZkpe+4FFCrB0tlVIekn3+cyQk37+ihGE6Ew19l8DoC
ouSSG5vW22VDB4iFlTBWirm/L7PMOfpiuwFwBBePRR21rHZ9hgy7zEp3jOpdkXnZ
GNCQZ7d361S3Vx2jGgmWrmFAg6X3gTT5R5gz00rHoNXm/iMWz/bEnk5tNuM/mnqt
Y0f4O/3DG2klH/1EfrpyYUzFuG6RrKGB+TD8tBrSNpA95dkv3fACEck07y7mjqN4
E/tqWShRJE+E9q7tK6dabN//sNdzaTtYXBddSxkFTmqh8yeVnkRfuwv1SGrsQER3
2i6rKOQ0jbNVb3/jIKWvTmgPws4jqTGGSr/vTx6ufpGxemK3YPtj3T6Sutg9FBSu
Ke5k9i50njwsKqMyonaXDtKDVsShNq96FBa4DNnll9O7Bj19NATx8ks5mxV89Roc
cUxeOu3/z6FlAJwqEqvKD0Tvhc3ldqzCt+7N3UcOF9rvTkZ4I5zJpUby0xgpe6/j
Uo/OXeKIBxe1iXnWedOcQrf/O+b0ruxAKgvFZTbUKXP1wOTdS9DtUUxL1dwu/4Hf
lH4ZY4DmWhDN78d6St9KGlY5qjczoRrlDnQTELYco32JqGxn2IPfzQ3XxEMLItMV
9aov/jJ8KnjUWTIw9O2Pplvd+OMpKZgvnJ7nSrkOR+rqbRF+Km2Pmcn5v2QrlqmF
qzX2Z5nPHJt4a8RW+QyrbYR7+SVObLOOx3NYL7EWLWVVwAZwnYfAm2eRHHlo8sMg
7EAluZBuCFiFy5S2o0zATkqCXce3DBsBu4WfqK+bh7DZPo8Z7clsIyXm48mCY51e
XhVdFFs/D31uhKx106Umdnc4EKCQtdMSwKMaldn/Ym9RmK2l0Yc3AtiCuCRFfSzT
hp19/ypM3bl6HMQRHNQ5yl8/nC+3epTRKYcJv7z5Q9lEZMOBZ54sYdPDQ54OdG/F
QWjg+bY/O1v7fqzCT7cMRtqiYRsHyBHdOC7BoDv0/q0cienaSJRy4DK0yL9G08Co
6bL46g+U4QP4n9TIMve32fY5KReI2UkKXusxagfHqyGOeeN+XzDeigszK70mAWhU
qpgK8e2/b/uiikbzQtc6jfakC9pReeqPZGFTq6FZaJzUM9d9hOFGXhJp7m/bKDMD
7H6AtUpXxyvfMmToqnX6rZwwVPPh1HKcy7qjBMSlV0fbYwhn44im0Euk+aAN+Bzw
ythLap+wYwAU5Tzh3p2BLuSTZbgtlLK05cCpzwN30XEqx/mhFoAB+qTeVvzjNYHD
iy5Hbk8o3Jw5HHhqNIZwevcYmfXDEeGCwUoTIGV4BVA0eZ8ryNM8QO7uPv9A0Dj7
kjrDzS255/h2Xz0bW5ecKgsxCBfLAI1lZ3qwWXw8A+VBGxj0jYc2eLpvdQMgr+M2
AsnpnzQWIKyQzhKEXbstcHivXI6O0nUO1CoIuwHKVxhxV8x3iFOQBSvET2hWhG6l
1UM6p+xXThqxgBLX7lUj/NZmwmLoTn6B5ifO0RNxL2unwa5U8fgGWQq8gym+6f5C
nYJ8tp6c6CTTsZWYLwQ/Q3Z8jt+DI0tc1W+GwbBAVZDnd310JeIHqIqj08xKuejo
9BCAZx7ObHvXLNsPCMN/Rjncs2ysPV1RHaBaS0ek6NgzMquwTlDxz4P+4kjJGYQh
xcjfGytdE1cQLAH4yAGkMimKxBR5lg2O0xlWp98QGhvQb0gVTOJ1QQ51FrdqDg4S
Mq9v14JlXWEjj2sST4mG3aLkSQT8gQdaEQSL8m48eqh8apjE2PMDBfS9AvJ3tGQn
rDYVhv8Et7jElyxqFjBcbj17UwFWUzz3U/hQI+CSh/iBHmOEkbcJIInEG4XYu0MZ
sOUdLDL3vpdTfGwdgBqJruTuGVgVCxGkMCnA+4idSlfnFcNus8FD1N0Dop5ndqYp
YKS2QvmF35+0vS1IYX/oYEUhlR5xWNCUrknBNSP5MD4Tb5i9P6aWUkZqO7jkSIbV
lTe4xURj+3XKSrqhsGGrO4cuiNiJ2CPqVat65/hXn9jNdQHu7tNDlk6igfjSTAFz
oitJQ+Qkz20wD2ASqXCP/eRJZzQfN0LuiXGQROp2AdDl0FZqbZtIg3rtjBQo2vkW
yqi6JMZa2Fm9yXtxreFeknWxbFpt+UXZ4hKc4gAXNzn2zs12ezu3A6gntbkxuhrg
1l0qmUZWau2qOMvCozuy+8FWWb8gVjgnKqo2CPIQW9L0iAnt2yMPgXXR0/kV/jIU
thxLWeO3VTJjuOzV35gIAOp5ciYyTXritz/ET5m9OfBbl+cRepXrnOKSyrB3KR0W
lYhnfIKr8uWTmWayXGyWOEUge79Dl2OPqg9wQ2EDOGW/oARPubbe+2yUL6AJBa/B
Er9NdC8+45vfDdC/HYAhx7liwqWPHHlVkQFEyv7bDUOlJo/IjqaDJj/K4OCN9sF7
flh013zSq0pZkukiHGnOyq8PAGMhh5vAIJY8bfZhGSXlRjqAAIgso/+wwUY+Xy8Y
KxeR5y3rLLzg5ss3bvCYLB47igAEPkGWe238BlECOIb5vH6N8vXYvYO8uMrXLIyh
vOuXpIVmuPQSvWZmBR7GFNu8L8pkp0npYl/bkUNZKqLeQpkR0j9Q4vOqqgHY0HlM
wc9Ip2ouLRUUMSYyUdCa/H6zbuJT/zqM8LJ0Ms4WUvHgzYwppLf6RIAOFK2Bi2+h
2oQwul9VDlzCG29+n90UAnQUwUdqnBEbUu/B+I8VgwUHBYaCK4onVPJ7wPwbCHUp
6xto/7rqEKaGG4GpUxqe5ow0FN1pp8y+QRLTlECFhNG+meifx9b2BgBpM/ghyAEj
xLOBUBJmhhMT8vN1Aa4qajW32EqMEqCPxfPwIQ6KAzvA5UIY4X2ILwV1S4Yt0ev6
9iWif5Tk6GTJQLOVyt58qLmRPNt0Xni67SIe3CMSYCAJEH0niOHcQafD2HzB3dK5
tEnxn3tkjGK/WfwPhpnb0EuNiYxdQjOp+rhEG0kCMgKPQSTejV6553XpOvqxSxZZ
pY98T1xc6CnlLvXqYs2GKgGbqYENaek/70FOJIX8Zec8sIhb0wrBOIPrlTjUMbyh
rnc68RmynPkOYtXYXOwyaB1T/MjNlvUoppuXOCcHny1Iizk2WEMXm6A7Gbgx71WP
JmJVD4igwwz5UnasFJ/8WZa3XUuCvu/2V+wo89BeilJr9x27DRf8YizJil6vqDbp
YAG58SYDlF4AGe9ATdcFwDJwQ3Yh4mxFfBiByFvqs4sJKJw2Qtqka9/VQ5MPqLv1
r3S3fnVMiDxHaZrnp9oC4O5rY8araTau/JsKj/Tf0Q1Npq0UmxbJn28hU4QVpMjD
LnrCiDSvaPouHO3XvqPOb82dfzbQzcGDrtlsYH9AABsn8IgOMbW4JMXqCyZhrVwZ
Cvum5CPkm4Rn7sTo6ceUg14C6jhngyBaZPcRaaRkuprRgGGP7wBXqzEa+avfqN0p
1m1Ad4y5QxePvpHbt95pLKzKgQbuvaTUkX7lqh5Tf0t9vVgEs2qY9iwKs+hd19MO
fFDrNqc5gdv6liJd3jMeGBzzrB32hMoDSNRTWIwTlZyicrsPI3H50pZioWrKUbb/
S+IVib23/62heJL83nFE1W3zTTN9hFOb2oQ8wrbQj9izCWERTgyohFGPeklSdQIa
GsCd8Q9lA+A+iKEC77EYgv0Adu7WQ8rHnzc6DXFwkZhxK3MwWlYd/3K7Un45pR2f
UVot8QxExhkJwSd4o5RpEsjtLtxC5cZCTTnpiE/+RGl+2PrUO+e+ULeDwAAR1RoI
V1gkUkiVx9EVP+Y5gYz3jFpeGKghmQ64HQdFbBeSP4e06QdpSifakGasv7UIWezF
zhzvH2CAl5oI2DbifBFNY3KtHVCoBNxW+aQCsQw6wunZni+T2gnzmYZCiZdwEOJN
ytUzXkXjEiUF3B3hwnDtbBCzPcO2LN3V2PiOcn5BOpGmTnAhIQBf/NO/nrE8wd5f
uYnLyRSLFaePF7auUAKwPZRSzY5QUWbuXkdgNKfS5Z08fXOF8CVpUjCM/IUXQ6Jn
OITlVxTk0FvDT8FKpsQdBgjHMJrYjTR+3AX1UJDsBJNZgixIimnkMAWBkeB8wfFa
UDIVjZXgklkLo6VOqg70nCZJEM8vNUBdr93dnBbT0rYbR0+2sUhUO63de8bgM/Dy
L26UKjdOjpTNKRmbUICeAKj978Tqmg9PcP1SSYw6l0LCxSpT/FWZQZgT5w1hB4Yk
cPOic3pZHfOfeAAJVQAGL3R96AlxAq+Hu1MDcFze2P0wSdysHveO8MoFlmVgT3sK
uUiIyyNXV7PEdhWjVg+mvOIHLpS+QuQeVy1bwl0Sby9McaIqtH6jiz/vm8rCHOcJ
4FRHD+Fyb9KtQ4lDMQcdPLNauqFzwk0AgxH93+eyEvEjUOw7y3UEwasLN9NRm3iQ
obEvP5v5cHA0Gn+WdmtBuDKz3Gij7RwCTVxHvrsjRjSU3ExiLpAgzoMpJGQlUNQY
/VQ2fNoxo2qZ0oexa4pHGgao82E0lJi9Koc/Oywvc6atRbxG1UWBYwRTBuZSVgd7
n8eCW+CqMeKqPgMKyhBysL+2SSJWNVr/VQ2Do325oageXfgHS3/6JzHqgRO71CPK
EWjrBvHloSyDdFySoWjzvnCPNTSA8vfQVgrjxxk9X+xxzo+ZA2n4csXSx0yVqhbh
7RKoYaOqyX+ZrGzXCodAOiD5kUP5Ob60QqvoE+b1HD+y5ralK77T8/syO8P8abqg
nniNw1xrQeZH4LItltYQgJzp07tB9OWeBiAQ5TFD78TTh6vKVpg5CkePX7yl0F0E
T1qVsXi+WuelSHCTYQp4wl3WEtY44QUUx5UHtHpBSa7Xq/4wajP7A2UviniAMx/0
QwiYDjv+VZTdT2nhxD4lwzSJ7b6kqfOevBqXGN9GUOhVjNLYAw1dFLjWuft0N/Xa
WrXlGcE0vYdN+u4fA6ZB+LBVmIPPM5eOMuF8QJNsQyiVgI4sAR4CM25p846NCHzD
BFjs9oSFOMzcOMMopYWAcGSLtIEuONgNcAVNUWr2wLlVr7IL77MVCpPpaWC2gV+V
cIa5P2ILayrdmlBEYi7RrBhlTEh5lkR2piWsvSwDAHJ/sC7S87PJN1K+jmzIDvHu
v9sLCrBQK7xZeHRgdLco6DsPqpBNc1teFLLfTnlXct3YFUu69NXzlbYzUZTMiLek
qwqKG/2vesz21TyaDQKbEZxtns4UPHc9lnnCVLsKARHV8VdnAGW2gC7s7gQCEWPR
HyspX9kKobz3ENeAcZJC2VeD32OX+Du+qSb6hh9y+3x9xxx4NWvYYSL8O5+bCum1
E5xVGOm+p7IJ5Oi5v3bvaZO4O0x0Y7WojUJ53J8d6v6pn+xBSIdfkkQ/hY4qF9NG
jhpIIXjDM07wBMrofbg2pw0eC6lVhYcm1IERzXGu/LXTqSckiEsFtFTM6iJqGpva
w2xdEvz1iTT20CEw5F/Xx1oeH9MHrCizodsz88oGHChcxiSEzwPdZa3zZfauaJ/V
KdJ6GciJ5nQYai6zgMicotrieHqlVSVyC+JgVm/MJ1ScSy3LlsKvxGQerNP95oWn
qKKZDfvxOd1PVSakBwtnnXwHAiPHF7lS0EqTS3yZx7Oh7Nr46hLmTvdVdTHxApZr
+J7gD2N7BmWX2wiLZJBJCw87tVc8PSTW/mUBf6LdrMuH1t9+AdLZ+nyfwXJGMqVC
5mNU3iWF5LFEw4aJGv5kGfjwIMcJSXYTPLlaAGnN6G7o2sj0MWWnUEW4eMQIi5Eu
Ev2ItGVwm+5SJxYmpVpMiekPQJPJA7+98NbozwOPLBWfuMLJ7Buwv5y1bNGRhqdw
5DDqUCd1mpwh5qgs/PNclUlfVWz1DAonGOWsVNK6g13g0miVLoQK5njMmbUbOU2S
MmVeftoQsrPhurILuLZr76jw/XJTXhqH1XnilcDx7C1OPyrD1KYl+39MsydNEs/i
BtahMSlxxGQ+O2b+EXSK5FeV/pnkp++DZ9vT8WcLFNUd4beLkvWZFDj8AxjRbB8Y
OAivA/9grW55U3/Z6ixaFPEMEdRgUtTYYDxjMqRKkpyj28CkAqcDa+X2tXqnDmfQ
f4xPBNcfxLBQ+C+dX80p2xlDdF9SvDGdqt6Zrpd5kclrBwSrWb5TMR6PPNCbtYHQ
OFkk+pXpVQTZPMbeD8/pWCqXsitGYhkXz6TfU1ojykFPvfbsj30NNRYkYOkIqok1
Yy0IkaJKv/sMihAbkv5XV6AY7SstQ2iWKqWOP9EADNIFM6CiZ/X4Vj/7ZrfoFaaO
2x9VzaOm85W5a8TqEW94yYrCHfsu9KjzJ14t+00AaY4JOahlUL3mQmv6LH9GyEJH
UalcXFtmp9GucKRMC04TR5iOQKayuFxlcNqDeLwT3VrfVYQA3kHFcOR2yZ4l9K+p
Qc3Awz1rTCGes5V2QBRgLTMJzd6LtPVuCCu/LKZ3vVMoyUgQByJCRbluIq0p6jmt
SP/lBCvummFhBsxWv0S3NFmopVX8uJyMnj+UEXDPswg0rdk1Am/sOKIfx7yeTj97
59+dYquSo9ALkgnLuomVm3vqbQw5PDeLkhXCnw3oghckQaG21acREYXzOE9Uy3US
PnPvX0Y7eqwe+MPyiTif1yEA8rg8+WCdRHAOWtiAb1hXBSAEhtAo3napz+RPAga3
fk9hLRim2aV2w5ECMOzIiqSYihw+on1oT8oBiCCL5jWdAqIV+hh9zVCfz7kGXJpX
xn13BJuUsGYJhHK1VS9NTVyBeTcNJxs+emtt+4ujT54AJaOYTZA3ckJq0ObRkL6x
1UnTW++jZV52+xStX4Nyo97Im7h4rbfR68PrQZC7kmifsZV8uhUleQ8/6Y5Q95tU
PbT1gePF6JGHLs2+k4edEu9wO7xIv08unfFysVah2OphkiPTbTwIU8+cpL2Jl6fG
vG1q0gCiaJbB9gTKk4mrDkhV9jE09iF5TvurIDHT8+OvM3Hn6tRVX2bXucXnXhaL
XY8xKim8rKV2FC4yBTN0N3ekALQkmf+Wu7d+KfmLoLtSa5gctoS3uSdtt4G4SSr6
LpS4CAudJRvF0EwuSpTNVEoE/rTAMvSSTepIhLHrCZFFSYEJomJbqVaPA5/sby6T
QHgdsNsaTxYaHdoH7q5Fl69vdnQkytcW+AW/En2lF0zdeSEndLho5rrYtNCUYsQ1
tGwBQYn4TNslQq/iO1C7Nxnz5mbJwOJvvoAl4ldf25pB0NjkQt2dvrOPFr833K8Z
+Df93pac5w4i/nFwAk9WN9l7I2KwP7k4sapeFEfPRjya7ol0dXMYWeHsmJ2OW1DH
OgfCh4UbFPy36LCOCpNCzTdFxyqUNGB20b00a0EMHXQEEBjiK69fqnk9Cn4Pfp1z
slGkG68tViVqsS5ljPIh3xNGfNthvj9Dz4yytrTHTzEvQxE8F/HlNZYupSj+6ZRt
89CgAC+PUhAxnaDFpj7ugo8dwX9NGWXxCDYm0z1gcB/v2EdyzL477fx7A3iK8UrP
X41zszU0puZSMIKQeAqXBxL2/RPP8BnlXL7oBFdgVI6fnTw/JosE7cbXNjOh8xXm
bN4Yc3l91gQr2SmQBbQZUY4/YBcfrv3/pqUiH9mLhRS2pseHpXUS82MNexKjfwCE
J54f9avLR7G4TXfgTx2mAB54i9VMGSs//cxYVCm3w/Bmyhr0ve5R39yBzGW6KmuR
ql1GduYs089xIuFBDzdVXh0l4vEWVHT0vjwa0lzEe55fGV3LY714XGn0dQxBSd56
fXWbP5/mAVY7k30ybaVNmI4rk6cWB20HyMMgbHBFW7QJTWOnO0szwJsdswxMse3K
ebW8DB8jkPmrtQ/oWlpOUFtnuSqctkAdUyxUysHm8zrt7EDbo4hTb/6O9cby7ibE
m7OZICBCMMLhkHrVk8AoGKIn71IdaVbsVDqmZyhwAGyoTOgrM+ussSxyrN4opgvX
kHAiGNUN8iX0isXNJRwlV0prmn9Rv4gCVopKpQ1RHReuThx0sAh6/KmCRimkcvwL
3R1ohMZYTJQVa8k62u5M0JeVoPBfuHuqAQQUPRrMXlzZsw8aAqfk/dwcjjfvwYiG
agGDCbeRb9MwOQ0qcv6vD9MaxGqUUdmqIWpmR2QmyHvKhnThWCwib3nfrpGR4b6M
yXoO88NIll3c0eLIRoZoSWQ69BA4jAqPVsqQpjV/tktCL+BkjxU5hYTuSvXWhHtQ
/ZN3ZePcUlr9UFBO2fBkIuj8DttW5yV3ej00SnlPZY82gaB3X6Wye1EMyatxyxcl
WIWWuRUZZsw9+yM1mIkPNYf7hk+uihbb2Y4UK8wfob6Wd0KLP0IpypzLeW58dIdA
jnA0KFuX0rmAxU16iVhLTlle/66IOQexmZBNBxRCVgp+edahw8yt9kvmMM7GT47F
nxbw01EEXnDxnqrcrfxmUnU71y8ilpCEpFxDmbsfwTgAiJBUdepcZooLcokkZXtb
iQooYuEVVsmvTjCeLqjzI6CIdioiVx455NtZJafNlttml2RTeRESPKS5cOmnZ2vd
KrtZWoN43K/iKluehD6+1CrtdKKTxbsoGU6ytlKwN6WuJHQitl0zHS9kZkJ83U9N
1f8uT66I5vvu4mex2+B3bvjveaF+0Rw4qxHtrLJA1WOb/V+u4piD+x6rw7PaJ69j
HLWyHaEPuJ5T+5AOsSBJHc1MCB8Es+VCO5222DyaJ4Xvw/RvZPYlXn/AE/ExvUvb
VS8i8yNG4tHR0QntaAAXxl+jvJEerBY6OhQQaormsspAwHt0UoDvVtatLWfEoCaN
7BDki78a9usTsQHtLXeplojbxcdsvD0dQ8IqzirbJB0OmG4wRolBQW0cD/RR6hsw
bbwA1sYvutomxoPuK482aQNirX18gxGCqCt1HLtBK8WoTulWOqhNgyDdmT+HqKCj
mB/csTfBk5TZxqyBGgirIHNSp95R99D4rmARaP+m8R9EtgZotj551GNSavTYjw4R
WMB3QVVVtXAAO52LGlRCpVXzywWxDIt8HnE2oYnkUwpdaUImzKXvtk8a5l779vMV
XXCHo0ZZjfnGoPQh4gtfZGuKZN8ILKCeBJb3ZTQY4TI6IKDws6YiM3b+0TiIjssQ
YuQlGNAhWjQjEoWItEb7nshHtXWkQbvh/ONQUYGV2RzWEvxU9PinI0hRm0FRf8R9
z62ZivKJe2ri9psBg4RH7qksulotRxuvknPs1KrnACPrPi4MmZZlB+qj0E+e1A3e
w4Tm9hZ9CSesJgEskz+F7AACX8c+oy3o/V/VjyQeqkbVwP3IybuD1Q99q5II12Nt
0cLDKeSmry7kpdy2OlMwxgrak2oXLHXzVuNNANL9diqqOfKZaUM37Ccz+mIae1vU
mZKvjzBrcOg8SNhWNhrrnJlB+eHhI1Yfrq2oyptOsIHmHb/jcy3jXhb3oIl6ICSz
K5pkuyoIVc9s2kw/+fN2+/hxKWBGFDs6ChGAU3TNeH+qJNFqfl211z+Uae1W4O9N
7UbjM+QMQgxY1Hsj9zdlRfbetYXhMsXOYtVjHXJAMBnj0XhFxjm4G4NZqrhiKDoC
bW29DKorh7Ze3+PpM8c32ey9tsYUmUe+Ys5snmNvZEf1oXXAS4waAwyt0+YBxDLh
TYgj2ZpcKW/wc75L1jfEGv0zdDpcJw6YgA+Jrp5IkWlXuoudMkhwsQk3d0WF4VLr
1sWcsD3LJVuVxO8g6oPbORQEA46Gc7AR5W+TRbxzqOKWb6oZLWoXSrhm4ovbUgTB
JPeyzCpxb4XdIbnZ8dtXTDboKcrcBWfqM0ubmu36rTM3/Ko9J8gy8ULbymX3/NpY
2q+s+lKtUSWRorI/PdKBrfUeO9rUPeDeHAWlee4EvTLtyf0Ld1393VWNsrIblsyn
si2Pvgp5kWcKUiBvCyPDMENwSTA9+xMzeGsJuzBwM8IB5DvFNcLutkH0RwuCJDZw
ulk04/IyvIUVbSXK9AS3ZZE2bufTMN2ZfEMsjmvKpAQrEp4ktG0Zs29B56Pu94zK
pYAnumgs7rE0hTV6y4ocZsa70Vz1BTmpRCPH/xHtMK80aM07D9BX+bPVa9/YIC6B
sWVnzezFGBGB0dvnej+LiEpHpzNM9X699CnDlQ0MZ1PNHGtGsPSpgucltSVwY7R7
ygtNr4JJRxXx9kJHSlT+KvnuxHGQE428Lc6a2uKJId9sRnqxYW4l4jmfWYSvWnIw
1vDuLF5Y6uzUhiFai8WPbavxMdezAm5Op0zcljkGkT49HmK5RBe9YyQVWbQ6stp+
y23KkTrL3zqm7/oKjZlodhR2Ss8/EptgsB/Rik58BmlMjKU41Mypic6Pn+lcplqL
xQ9/Q00vd1FFWCc8Ecs6zwqWcEVFDB9BcaycpdJA+RWbUBlyebp7tL3tTdjj6A6d
KBIzPCmRlM4r1ITUM3RKtjhGRjUpacFtpaRzsu8dwxJ+g/l1jjJ1RfhvgaIfM0lU
UakAtVVK8dZQ4OmgWL7hHKN3xHF7+tr3MpebX9fdGTOs0ELzjy/t0fy6iie78J39
8c6vxEW/c6t+SYkYVhJ+rCOQIEyndKYzYMdYsPCmzLYS7Ursl4j9s+qUZURpTV1k
Vc/pyi6rhGOguSb4xEfKOAU8Fnmha5mKC1aC2AY3GllNZbpAALDEJGQGVrsoHREP
kaflEFKlPwXwV+dDb4ZS8Ln2Ur+kUWbt55L6Flu9JZATC+g1c+M6WRYun20+Knba
eT8K4aSvwLaQMBIFCKuoUGeuesZkEuDn1NFbeIdMST1IrHoR2fWyCpMztqBjYraB
j2TeYEtpYhfDGyLfwU3HkccEfhDzhXEAeLojjL23MG5b9VFAJ0HxJkD97cY/C3sB
ffeYKLleiuffTSOMY2yb+GQZ989wy+CI+cucQJa2/BMHXErkDaolyEq4G7cikA84
cQkp8f+0fD8abmIhTfKYMx2mJtHr4AoPZM666Z7GfDSNVZ0azcIrRwn9Y+tGv1XI
dA73dw2wxg7TwPk8cPpiFooGkPRCIg7Iduu9JV8rx3dG3AqZFnCkCYGAcloQc5M3
IvKAXprYIklqe1TDUkRwLT0XQjrIJP+e1ZmsWMAtm2glmEDlnYoTm14kj8Ykr7B+
taB+Cfdie/Jm00Y86+DNUAYeicajPc8xou2wVe5MPgk4wSS37DfmSYHG5aG/1NLw
xqu/5BcLqaGbuBWRNPDn4XPk9LW16rmTj0jHj2fZT4W5MPNLnotpH8xdX/oIivYf
Nm2yLh5JWHRRExcY1LL7gtVQfVAIBfXZoHkczAWAzpj5zQMjrfxTf/bv2Ck72QLv
+t5Ht4hae+C/iZx6aKUH380USEqT25vqOKxpZ+7ZsYzfiskUpcjTvCA2blLmQMjc
/O0gLS5PPV+CJuWThXzJfnQqLKfbIEr9jB+DRBCvJl5NXpz7mLzESbyl/zHiR8Nv
Y5JpAsvuYVZfz5H/+ziclVJ5DI13V3aCEaNKK4z0bD96rihQ7CY+p8SFhQHMeA7d
dvfboI5EWwrAVfj6snFAUA+Say1ywrGqAx3Vw6ltl0inpzI7ZD8Z4iPiRFIfGzXo
U0PPpNEwgMJUkDQ2EdA3wB6ACn5HlCXIgxVsbUDQNQLgfHjHJ/kA/Hz+m1ztzxyY
GZ/buF0VFJX71TB0MKJheTYyVTOPF9KEuToxovM4VLVlroWDXoU1wSwp69tbIVEe
amTSU9+zypJ5t2dhAL8DdhCND1Ws5UUEmI7t3j+0onlqLyAnAfrUuQEDbl33Je5I
6oYfLKxH9omaC+QIb0+E+VC4w6AqtnUDxh4IsA00fIj6HNyDFU5neU76CsyAhGDk
JFyJJd14p7sDohDPTRdg5pTZa3uEsdhNEHroc2h6N2ZJr3ZPPy/XvD0xAiNEtjpg
CQ/pIdNDs2QkSJY4VMRK+3t1gidPrgcFOIRzsCFoa+VHZS988q/5XDOYCzEvh1c3
oV2fp9osfi2ruIJ/Wnu5d3J9EG7Z97jBfsA4piEHaFq8srGNMmcUyoJlR2XyKz9Q
NfUzWAVMifUfw352Eorxy3iqjZ5Pj+o6mnwByoAmwygdzesqoT9BAn+TUKeCLz0s
fsZza0GYWbPICMWn1iEr703km/7eQq71K+2l1gKH46qUfh98+5iaHtxcF239d1VR
cmdGipSlXcGTMpKcUeQR71a7e0NB6CLj//6eXNSrK/0Ba6ZyrFaoaaU9NsPsSlnw
u8Cq+LElK9Xt2JAjIppOWX85iTlD8Hq+EW1Gq4dZHghI1BwDEdUSeUM/3bbWVvJo
3S3QRpMWWj1WHHve99Fd2m13zXc9FBaIMrj/JTR6wnXFyZ+XljFJHf/w0+EtJ11X
1FQMSDakIOcSp0SS177atVwArPo13ydPDL6H+SqqocPAPkOIy5mTEOJk5bqmk0HL
pjm2+oHtjswQlvinrf7u0bTpGejwHgT5qyCWlzRvFTx4ax4N2BS5DQg2WgXhV0XL
wJJlVdQRTOfA/9cDKbpCfDS117k74HhH+rGjWn3yoS3bx5ZjyaAhhzFfbzaOg1bu
Gjp+AOeWdx1fw7hbwgzWUe3spSvaV1ZbVuKScZ7lGR1EtnDFMxJlUEPgCXAzyAnU
b1cO6w5rMjN0AogVVTZpKefcdn4yPyiY6JfH3kLEEKP7uzEBuXypOuZvwWPntrfk
iVnDKlVFwncPQ369T882+GlneWPscwDmTAucag3AcTJVuPDxydQTljB5nvhpqrz1
tTVTBPiFOvQGX1y0Ayfod7eLxNAOYMEF94JwyPpjpenbzFPFIJ67L0XmBmNvRz/l
iYcovfPnhWyFln5vUftvquZVzBJct6EH5ML4i64CsTt2rTZYL8q2oozdi4YeA3nz
a0nAqzpr6HOtLJHK5QA8XgXPRnHU3y9vg3Tmcjd/x1HVWwYFTx/1RmKNOBOv71JA
oHb0tQmlEl6JyfkVm2EfPyp75nq9Bk6qg26p9nSPGMuHYg0Ib7xcNSkFimzE4rD6
szaT7F7LKqefI6BuSWbOYe66WMXM8GyXHgDP9B1xqlpcQcKbO3REg6fSxHNcyBm9
7NKCht4r/sI+1iYyUdbHzQKFUvg/Kxb8PrxaE3zuGnwYY/BAGXy8xpAq0o0h3Vij
4szDXRCTrpCV5rtkji8qs92dBhKxiqyBGY7gRNYjnIbk5h0xBDbUzszWv9l/CrWZ
81wrXu9OxIGymA7q6YYBO5Zq1SaWYCmkDMPY8BFEW2+2ipr9IQz2jpTmOq33tSqx
mvO+ms4vO/oNU/YFTF396iOpfuXNF64OLY2kuU/t4WyLwkFKFZOdd4fsWhoGfUv7
YgsRRGanu0hwX5g1hbqTm9RhSNs0AduAz7RQowtQcY292CKC+ahrpkyPYtYKiPpL
20moClcMLCfBuuevEoA+AWGM4LFOqH2AAhtb74ijjyBPCq27vRlvnslSOi50jQC8
ApfcUr+CzvOiNkySIvKxjHcS6XSJJn/B1Gf1bDwDy4C19Gem0dMiAunVAB7jDLYA
mRD+3MyiFmvBbcZ71wQ/cNqLZfLCils7MKDzWu7YipeWEXFlkBHsiJJz4rlvma1u
UF66OqH4/vEok6oeTAEa8DTL4OxJmRAj954TeJl2a3m6nzhBuLq/50mtmTBpA3Ih
iTqRf++08sXkTmViq3ha7aX5LNxGcupIW0e+6u9D9qMXH9ZjW+cwhb/CoRDOquAv
N2UdImFc6NT4eiAuDFknZOnEYkgjRoMee5xRZD8d0dJuZB1saGQbmwomgQI17qqC
w+kb21x2lfm4CJMngEWHZ1zlFoqvlPf8EXN+1KObatN38tKk57RlFdmFEVag6WFD
ASjvGAtaUnw1H7ZZHEeemJ8S5QkTEcKEELpaVK4PZ/wdf4GSu9CFe8aIO8ECXcJr
nrteDi+XegITJuRNkn9wqADj8GECrePSXS+F137ZZKkAuWFtVtR2zD+jQndHgPrS
1vlX8YQI1DLbal9CrQEtoGMa1EHGme2ntfpQ5CHiQfJ2BF87T+zaIupXk/Ho385N
tgyjwhao7qROAqKPU8OIMfcbBfcH4cazcPKYyhtaXhDXuPghIGmH1dQ6PY2wUluI
/WH3954KlBgNzxgbCBgO6NJW2w/R9s2UvncGS78+lyiXz1Z9uYeOGb0Cdqn2broj
DTzLNxmYRmF5uUYULv7C9iB5Pw7jt6BrvZU9VEHDMcEGS2he7fVJXos3FJnaFsNW
9xda5u2reEk4Bk0toXX9jrI0UvRusOwY7Ou1Hqjr96sjQFWKO2y4zi4sJRVTjQi5
MJleBBpTORLAy3vGQQFpzmYJmZ6GioHX1wjdPOlMVzenKibjlS3cRnGuJ/VjG4lw
O6SbG+EbqwRKUMgA6fOAKY+dU374fwdkZEIsu19KunzvcZ6m+8s6jkLesHcPYJ8S
StHstMdTfrFDq1iAPe3IpwqpNc2rLdpnSXLci8+KaoijsbptysYRo0IwnMY/XSh5
m94KagrmfK5/aTvWIyaGoGt6krAY7gz9ZENqBKYVtRVrJsLLeZOlTlmFbrfNDFAC
7ECBNapyOjHV2HmgtLt/z49qu2x+uic9XYfa9W4gOb3EKOpUaY0/aDwmKvWc3QQ3
7WNPbl/3K83KD6CvBSh0LHHmtC4JQG6KcYhzWrrBTZ7Aw3yh+YOjCYksjFE/k8fb
NtsOHqIl/gJb9n2fn/TPqk7tKHnSnTDvY3B9B0JSGbLXAS7wYCn2/++ZhBZYrGBE
6WgXpOEakRsm34FHlHh1hTFEAp58MRu9+y7U62BItnaDXi8IRTwSNKcY27kUVyag
Z+89nfWePDFaibZnklct0IT0GLlYT2tpcIVRiFroqbFmptb2Ue4YsnS2tXn48XSC
4q9qPBiUbPmN4bSJY+7IGfcBSRT20Uu8oeKAl5wFRX9mjzuOhRcDi5xIzYt88uyn
BxjYfdKv7keC1mDMGOTx1CavozpmmmAkivptOvvMEftvR9aqKkFJ9nJpkljXNIpd
Nu7ymcyBRGRe4SEq3UZmqCD1z8CnaqpfSGvi7I2PikqKz6k6bNTGUC0hWiHT11MR
Lrxk5EziOHpLWP5BvRTgGefGGRvQo+Y2AbDyu1OVY8F2o4XIlhLUC+vYavUJ064c
cx0S2hGn9WRxMtR7UTYZRS1b7NcmGR2AQew+NRPlzwlEcWSi1QK3rdoRVHFAcxir
ZqN7CAm01w8vSsx9YSrH+CpLEA6RyqmS7SV4FmZ5TBcenfkyrkIJoa6Ro8aRUtpc
ZSfTnyqrTnfO2JRDIEsjpHlkt5krlYUcLaCXLSxCdnK0+13PJcCEddvfGgPunrRX
kvJBR5oGCHG7vNrXrHPhQD8fW/c5rnx0COEvm/wd+xoGFwcxcip1iQFaAG9uL/JR
UTLv1uUao+W0xe+H9lgLOI6tfI7e8x/bCPHvsMLIBBKOz+ges8RRj6oVCnUu2FG0
F/EFzGuOvLLKg+lF2Wmym2bItQCEFJs03fjP1nJHynt9bC+LoWsbC1uMivcA84hb
RSBKq7b38AWjru6ghQZwM94IaZO5T1bH3ahXciUNHkKSH1AEZ1N1A+c8MhV5LG+N
XR0QF7TzX4EQt1AKIafhlz3gA+vaCoKV9GyzxNi5kEzz0Egm2UWYF67tRleNAGQQ
Vh2+zo9nf1gr4dWyuPgJhlS8a4DldQoVsgtbgeQIYNaMXapVur6FnWivOPrK53Jc
nBytFkiqfZdh40kz01NzJxWvFjAEQfQ2LCwe0xw8070JMybYDUt+AR3JaUP8EAME
TJL23W/ZvQyChRGtx+1bZH6kjlaT/3EF9iOlNKUsQMpf5Nu3ktWSJBUw3BIpDvNz
MlJTHi5H8+GkyJr2jsGQ6R72leV3vT43+os2cmlKABM23QlhvMMJeIFYFBy0bBgA
fPCEEkqw1VnOH+Lqe2ey49NMTpCI2CpGcSOEkpdfQvVw0cPi9d+t9kTJ+kQ6RJWK
pkIXACcJq00gUhciBEXQJN6ESOZc5xnnop3o3KiUavprG7NhhQbCS0SptKPuLOnL
cyXVmpgQwyj2OJ1zpargU3ld9zmSIAoHOaGiOPb1cuo+v7HBP/02jlxzNITBlK15
2jrKoTAN48glZXg8psqtwBdnfcJ2H5WLOaIOojlzclO2OLmRds/zkMd4WlY9necs
bY8n+yGS2ZumjepACemkgrfl19ZOdj6LT0Gy7kbYwE3mtD0UHGaWh2RbsdLCukZB
8AvlozUQadwtAREanidl2Ig743XdVx3qWuorf+u6ovWk7BJ/r0yRP23Lm+tFhz54
5vd4aP8zQxxpsWrngV9DBZmKRGOhlPcni2AMjE3ZgDRli0oWJFnjOaCfoEFZ+xeu
Zav8mnR61loctcDJK7D7+fLxX0hMS/3Y/+2X3lRKI1GL+yjypFXftEGhvmn/K4rR
A2W8jYhFcoXcdcqc/sv8pagFh6Nnzt6yQqNKgApRX+Qg7SNubB2BWuLxv9qUDItB
pCZKAf7/AXB/q2Aj4SAOMnfN/38x71TZjV6H98rdZwDvOuCI4LUnvM+i5WiC1Tk4
E9lhpHvqZHhXc4VcmpCal/sK3MKzazbubmCybcMaa5lw5rCCQ1GOLxAKVdQ3p2m8
mX3THZwsgnZ2jofEm5KmjX5gqv6ZF5sX/5t8GMPfdIzCbi2IEkfqY17JIe0NrvGc
do2vUcJzSmt/33AMotxf5NxmJoWkrJieDSFBlBnOCa/IiSftQjMOXUMeeP1twncn
DTVRGISZHAxDMMTY6N3GogWG9AsKKE8pTpS9gJYnc5ze4qBS8WAWbOS7dn0I5C7W
13K9bg4ISpMWA3uCYqaBzkeS68Yn3jmpACN3yGmTXjXOTdqvbWWgYNEl4C8cb5r3
/B2o/KAULUNUt9s133zfAT7Wn9cCrFDr6b0k7OJdZQicEd93YwCJSe8w5d4sAGYJ
xDGgztTfwoF8/wjSuJgcwLzqY51mQl2FQLcHZTDmL9nSX694U+gEJstQkRrNHLUm
z94ymykUTk9LPJVld7htrcvO6QmOVLbTwedMw2j8rLnTpiMrMgsEvQELiSf96zPw
zHD8nHvbHKf9ZwyO8z8nJgtSqkIF67xZdom23FY2IgqlJxMc42UH0ogFpO/GWeSn
rK7RmwIuUchr/t29ILzkJJI38WAVorY3GV/dV/gndaYvZybqYbiulHl1Zwyx5j2n
wGTtOmVOqlInm135qRfcMVCaorUQd2ZadNoGcC7ShqwbS15Zo1RS1GnSm8wV2uCO
QI0UkEXh3yFV3KqjM/OifTvDCjnkSMh14Yyh4RZNV8z+GzLdQzrZow5nlTgytYqu
uE1wuKhDAzUIn9336ubeF/0fIf/D87bYhcXDgCP0voaMe852j6N9Y0hgShJmPjLy
4JPOz3wERnPl4RRt4tLWSEhgan8IYfECuEstjWuYKKwVar+e1/OQyEUKO4/XytFn
L4RytvFTn21AhroKZHqEzCHj72ovUxCddlsZqpgpHVOOrWYBNUjOr1sxQAAZaQC3
laeX/BPpqavv8snS8qo051JFA9DUGQ3TX6Kt8yHn7TnGbGMuPWYONpeT13gfYUH0
UNMFL9p4proXf18Npkm9fDbLhSCxnLr+vr0VH8wchisJzLvp8FF7u0rMgNjaA9kK
B1RRzK9FC14GkfNO7HKdqRSqk/FNko892QEWtxgDbU1rItgqzo2XrhT235Wt7tEk
RpRbT94/2Vb0nByRVA0ZSXcLBT80LQXZbDvT3wTBduVS+SeUFx1IOhRGCCKmkktC
gMo71oh7pueS+aP45cmdBBQ0DpFR+h9Z8hrtUHaUROVN432wPZTk/Au/Cshf6Ps4
IdD0K9mUZizeXqIdu/bFKffRVkY0nw5JoO7vukQj4/+Gpt0jzeUnYTOWfFWQBruO
et6FLgyE1f1JdPXfFsLnClzB503AQfvgcb2C7hOUHEFmzO7KvxSXtEbXe8ggBikQ
z5/o9hLUjpbhKHFsTRDT/h1lDASw9JW2Sm6XF90NX9spWrOU/rfTN7ae/kcW+Xxy
mwd16aLLABqZtZLDEmSmNOB7EOolQO1eUwRgN3OaYdBx9n0CpTpJMg28gf7xzdLl
d7jU3jhhq0Q+na9+Jybhs7eWNdeB9qXhG63YnS4f8iZWdLPEEUGBhzQCIZjtOzWa
lenFKEEXFZyubTwGtuwJeHhtgm0PTHLvDy5U+puyp3fhqOH/mn8gPysfgUhIs+x8
tjLD2sWjYkpBixSOWOSff1mOtLzzGOPsjhAHolx4rz9AlKO42j5v4cr5EzAHYARw
0UQjHGhCfOYY2NMDJy7iOdmrp2gktnNbQVHheZA6rj+9h+SIT0vdi3A2q1ooYZXL
HULNYgtAM/6fqYBM52MoysQbdfmRz4OhYx/9y/1d2J0+wq+R2WKUz8q+h/ecvl52
QeM10nRFEbWwBF/nAF0BPEgcl5jwM8Yb2YEdnNVbg6RI1VrxadJA3AqLJxWtWnQS
fQamurk2V4hw9ooD8uT6+RCEZ7V56/MN/SbpRZEkwf+879CriybXGvIf1XTnbezF
DpqXHZOwlM6OzWXd9K6JJoX3Gp+PiEKX59FLZ6emT2Y6hRqBPWHpRpu4xthkEKdI
GzXZqySLmULtfNh7xDDg15LoTXctaUerRyV3z87fNdgSN5muhon4f0Ar+WRb08HZ
7fKhupFK6JLHho3NVKimW1juUcdNs0xy9kslpvh5AEo8IT3Hdox0gJjDUaWKsvlI
HM97T5IVnmdiQ6sNskNmaIBwOgzQ3v4EaVcWGWE3inyCRlFBFL9rAYzO+LVVbmqI
C7c+OvPHLi6zcrwtX+16K3233Dz8Rs5xkFHZ2GLheN6R0xacfEyO4oo/C3xyS/uy
BOlEMYd9Vn4IlY9KCH8QFblMo9hwNf37ry2NxYkKoCROXkioAxkUgL3bcYASvLpl
HRvw2cvfC7vtDGNDhOiVaPSWaeT3lKcPHB2F9qqFPgots36iJVOiUOqA/1baOeEk
HJr46IWRaB4Ld8ma5RiXMM6GuMWUOe04f88fDu/XNSjAKw06mIM5TE41ifntUwnp
HQnP1jxPRLV/VsBcikwYb+QcJxqJ5LFHPL7eDk6h+5m6hLVWo7H3tPuFetOZ+zs6
WlG1MJyJfGQpDixyZPUgwusZfSU2Q0kEoKtQV5JzKIvUIC0m6bLW2bvw9gff1WoR
fr2TPitkVgLdTRRT9p6e4yfRLmGKxGvJjfQIdKbGrauY73vARhQhUCrGvWAXUm+X
/iR3MAWHoB5+ijJk7XG6u2yFDh/OvM0oHyG5Mls26WwZC5c307wEzApBfHeA9fi6
9Asedt6nOG2tn32ks1g+NegQ/bG32W8LWxzubJyZe8tJAX5sOKotMnYIAvDfMAQN
LWmAmRngacEyF2bmKK3HiEGa8WzMHhS4rEX80MHY99zVcaguJttZR1QYtlzD/jZL
dxKvd0U2B5DdzA/F1KhYq9VN24tee5Db014mt9aq1qLFegzNt/lrtT21q7svy1Ml
Co1Ky/TEjVLYAO8OOYU3yAb3orovS924GCw1iAWNrW6LpyDkQS3nxXyJMfAur8Vg
yoE7IVbuQpXgTheZ3hCLX7yVtw+gqhrnq5f7c2nBimciQglKqPsRA/964CeZ1hju
udsiWZ4XY+phH0e9ANAJNhaE9oapCpM5zG+VGxXHCFp/GWhN2j4IgHRJB3X1LqJ5
Et6LbNSplXWqUuoeKixQsOlDQYyj/MqjLnGQ6VwEA8NZ9qHrlkJCKWXUbG1SPvZg
REBEdveCiWS43W5oHNLtm0/Oeq9gXLBWZAei7LX/FPZqcTFBi9HXduY4yiVRx3zz
L8gzLnqWAdQeYDtLZ2aqVFMUDE0grHgjqIFSLqGck096G28pjh8LeW1K+2QieMx/
g8zaczKpuDoW0h44morf98BInSXN1bkbozWOfEq3xD/+WJo4U5skuxWmFf3M+mrN
iAheijeiv82ePPHQBV5Dl73diNrqdhC07LwhlbOW9IzwtkZf8QBqjxBuM6xCCezk
glJY+VkTok6nb+A/wJ0iG7fpc9wvcKSnR9DAxH1lHMeF3rie75Kg0ZXQQKHZ+cCO
DGYc44ZD1RRDwjGVYLJLNswhfPOerElngl2j7mZzNt2G8/g/clTjTbyy5GwY/LdB
4xxK7AjQ9XhZLDQpyqlIMQAxagq8/IniULaPPmkcDn77vRKtF2NPdh/TqqeSqNn0
jvWnn12auj8RD5XSwChfojAR86pLHVx9yerQRAdlcdGrflgd8Jyhz997n30TNLTJ
wm6skqgKYoFo29xqeHiJl9Mte1KppcamVppuGPd/PjVzS+G/m47w/tfmVAhDA7Sk
ViiCsXE17hFWnVrm3GacpSEkUYzh+40QN1W9OuN1A78EAONSMQv8stl/3G1XAdOT
KY+Dl+cztGLWwhgeAWF/Rd7cSXQpIbzhzyJsM2SFD1hTamtsTUgt8mtkuiDtle2H
MKi5/WVFYJzzdw4fBdFiG5pYMjj6VsprYrKolZZ/4Z/urSd6Q+Y+/OHdsUkEnGnA
c8v/ps6gAnSTNULpDYAqEgPTgS9l94f6sLq8SGC/pt8ed1yTDU4Ggrw7T13486zu
tEHvnaSwPYvt3lQE3aKlDHtc1LWThfXuztUk6t04SfYs/8LpGWTqSGtDkhFy63x3
8sPD0COlR8MtIp1K1SZky/tmPc0jzGBWt6zDkfWF0TKf9p3+gR8Pym4KjF3ErGNg
cHDAuq+K8GBJxlXNmHSWojx6UolEssWoNE0G+mqNopNonvZ0UkaPMsMfFJQsH99l
KtP31sGBuKxjsLezvVbaumIRCjaB5DRQUG3WnL+YNLa2hDUJc8Gy7q7HJ0DekD84
/aI3e+BqePPZepDdcPLPNGEH5yX55Tr5KH17Q2HTelSP6F2opkHG/LcJ5iOYFF8z
IlEB6xaeIO7/GymMRr1VRqwVtnPz5EkY9zVSMhl5tCpMyLJjcawY8d5j+xcS56Vt
QuM3pF0lxzkGC6b71M2c7p7QHXdTuaDf4dGh4FyoFWLhVQ2KQVCppoivIwdE+Pr6
WogJQ/wq9KPFwK7acEY+FRwm4vvhH5wUL44AqDSUa7SDFsrNg8p7wwefuX9cuVFn
sgfEhsaGbxrkpGDJlkC+io5On2pu+k6wjCWDs3Qxz+AS0W7ZYRGMKxssNM1vWY4w
QrZZ3/DYWus0vY/xMuJoIRZM5KD9dfb6Wf4N03dOF2QV5pNJKJnbvJJPQk+ETcIO
beri6gUS+Mi+DnT7asHhKUOEW9EYfKt+ve2V1ySKuL3V2MmQl0khQmR+Gj7F1x2g
TCH0mExhEr/ONCee+w/vNMuJqUvFPxkfiZjCAGhHKG245CgYUL8cPAXvNBqCZyjd
9CBbZS4ofmiyVOIOVVrZrocGVALK9rho9X3Cng7bOLLhheI8FufYhyCRmoJKmtdl
KDY8kQrak4OyOX9M1wmu/YFhba5RuFhg5ZtUdNA7AAU6VKRtJg7gFkTwMxPh2cSM
lIBIiU8YFIfA1VAjFbV2fwJrKW7Djqx/1Hq+pqOz7kD2Qd6YyN/zAGIM0qdL/MhZ
MBkAmxlWhlgV52tDJQkK/m9hHVA6c50GdC9wKuz1bnaLF4UfPYXDpHZYJHT0dBfQ
f6Q3W3OXK0oApi6DCwq8zMRguRNLzl+o0/9qvQsCfBv9J5RLIVgIo6X4/llYdXOY
l8VevFz8OOuA5s7rCEeqiIkPq0liyYhy0SE1e1XAvfOg5ds2OHqTFMvnNyeo0Am0
OmmPkCa3O3m38BfuB2HXRR1g5pYkoSzEPA9MsQbxOky+Kffu/0LsLr/qjvNgd3vp
9lfTq4F6IGevAONRBaWpP9EF05wlEweSbohQ+boopEEOTX6YKtcLXVoJRsRTbiLq
onwONlBFF7LvvZx/I/3Y/D6aj4Jn20o/p6oqcss0Wc/TKAIRAYx6mTKnkq8OspLd
dPiulZqaE7z7mbvi2OVTqoUyyFZSgV7J2Uw8f2CfEXLDKPqHtrGz1KAXGzhF9HIf
lXYTjwS1jzjHuRy7Oi4pELeae1LLjlg/LwRBhUDVh0p5vfaKnF2Q3Oh+Pf4s4GpF
AG4R2+OESnBrNBw8dch9Z3q1WTjMbh5ISxp7rRtpCnlm7XtB+mQA9U9nDFjrGr9j
svEHqk3E1M2WM1CxsA7o+SFEdWW3vodVfGX3OHyrKUb/KKLZp7GeBEUcitSV74Sc
RPmlX8F0iNqu8QMHFLOEBQ3KazMn839N9o5XXljrGjPgpAnl4kr9sdAtQFx+QkCR
VJafE3nJVoPCMEZ+n66P6NSIRpbWrydiWCAdiMlFg89YWpV0O6+bn12ppwoBXQKr
8OGWlBEuCNDXmmZht+KrMYluDB8sE6Dv2YG9XD6qEMsR4PH9vCBLrLvCA7mIgZNF
BVQwLb/kxtvGCP+7Be2beJiSz/wFC4uosp8a++DjKXdc34Daa7hwP1Tz8VgynCh5
mybGyxhoxXljA2RymTrEJ7taPfIg3LBfIqgf7wlbBkXom3sjX7ibIcjUsibdgPfw
FbdaxfscScBiH8kuwjvjT3HIu61uklk+3aZcH4d6/3xQKtOzMW3EgfzxhONwmWOR
iLgTr/gFwQg3WGZ3KlZv9nI5AbxJWXgxLekAfQq8DRZIKPT6kEcI4SeVrPKsEK42
5oQqRddKzM8X1FpLYtP6CsXUZIJ8EGBxRm4TmI4O7PtwG4E1IJKGfZeWzKQanqQh
xe1CtKG968Vg5zW+/hdkunGuQzzwhPiLyj9mVOyVe3RWoPid4fxYRLK32pG49yhp
T/wj5CzmaqP3VzV/D5RxxnriFTgvGbTAsUUxBbevWPf0+YF1yhgrUhflsfHXPl8L
jUS+41zkoqs2uDiF2rPRc4OMDKBymnXZ1ZKGpfvGAWwkyKb4//X0JU5VHBTrll7B
UtC4NBT2NucYAAp0yHfxCRpeTNdwuounU92l3WpWUC2Z4F5oZzWwj05azFFyHttJ
87EUjWTOmo/U2rfsRljvDYs/lyg4f41cn2EkPef6X1JnKRIqe8lrF3STFESQuxmH
XUcheFMgnVoMUA71zSSCkLDW6ob2RktfpGC05E7Cg1tfZdP/I3TQpLKce8X10hYu
XO+d7h8tfkNPsgwPwbNJ13qsFfnd3mVnQuNJ4y3GV+njwHU62sXXBpVTMP9XLNbd
+UahMoFiavjjEtciBGYHwnHQ6pVCTIklXYSsuyPAxvq1mt4vkPMZq8uk7/eHJnVf
qO004I6pKyC2khLlfRls7UHmolNxRzzYG/fKs1wAEBlXDX7aGzWucnpVpbU6bZnJ
ygoX+VOYmClI7mrrmPq7oz40Q/+2hRAYJJoZZsv64FGVS1lE68IaBKoTAOPntLtv
p6O+/7JHp50IvLy0M7D1ehnqvk1d7+H4m9JOBxLT61k1Q1swSEOWukocAUu9UNJj
BIqlpcaP/+HjZ2fcz5zg+KdRGTdAIpPOjy/PJCi8v6NliZzaGMAikRzB8/2QjoSc
p8+wC1uZNnss6ihk4wDkvcsaz06H3mt73Ve0n81Fe/vy4mmI42q4lfWCzEDjn5AE
RFfrg2qITopq/QErlyWxuC3PG0ImOYDCQlbQCZ7z+zMabPDwBfljQbbSko1vfwaS
m0yQKzc3y6XVStSkgpVzd+nejbfzSiHbBY2bNz0H3YmTxWban3qTVaQRyyybXeDy
ZLrvhj8VUl9Oti/k6BjOCmA5uCiQ0Pneqo/USSUpEud86eo8Dl8L1Bg12O4FZ6NN
7Wg9NAEa5TJZnyH7XuIvmT52s2mowB8kK+DqS6AFBpMFFjs+RBWYUN++yYVLxtcf
YpUiroVI5fwhk13Lo8bXUQV6V417V2SHm+JKbAwTPsyUzuzwVofHbdsVwpENRGAZ
TnwdE6s4GRm5Ikp0kzsretC3KMjHww484sf7ZkAhY9whrSlrxA2d6Y6u410htI4c
hFLdXXlM3qWEhoVDpyhBxPGDJfDvj/Z0z7dj6YcU53g8Q6U6iY07QCAPbPwVNizD
l86rUmBjbYekJ7jM5UbGuJoz3aeEZn7/f7A0gWOmBHkPnYRLRhX55jggzbENaCen
JVP+FpkcJ2Ki0QS6qcko3W6hQ1Bm1aTyMJe9LmJC//tJxKs8pAAyw7ezxH/nq10u
2f+pLkYudIKBhrOBEUJfBXPfsrMIY4boQzvUOs7i2AgWv2l5KvXbsRY0nfcp2Jqi
+1lowtBwK7FmRpN1VlBs+E0eiMMVNTzhodxiyVAAU5a9FaCX2lQTq6xbD7QAgXf+
itMX/ZJP0ZLCCLJc2T6Icri9cJvU7nCgtoH2oHXCZcNsuYq3ME1zSntp/vKlme3Y
mc23B/0ds3o0E0O++u0qrsqUmU7Mei0bmsBy6CUHwRpFyaEYP8SWbwgZ4bdS6vKu
dyOyWt24oCmfQWfs71jv94Oaxdz4IzKOldiRVXpqzf629mlv102MAkToq/IMRWU1
HiDvelEc9epFEIFw6K7sFHnF2MF4h+gkXvwN3QsljduaunXCpbSj7r6U7atRUGqU
V6H1ydH0PLaOOWHgHHu/KXB7jEpFj7vyPS7KCoK6QSlQZRDWFiUNHQ3BhYvHwTS/
53ABF6AlBJqvBbqRe97aecwr3C3dhRElpn2SyW1CQrTIO6BPU/I5qXSyQYLyxA1X
VIx0cGrw1MeI5HlXisMTWXKaI3n1AW+PMFG/Wn5y8yH4MzVbxbETs3NIS8NKJtyu
SQmlOsq5IfE9CxduQ/IYHa8E2hRrxGEH5tfaJ0vDYLvfGAAn4sQQRE+mdokn8WXX
mRE3K0xr5SONkjwLC1MdoysgoTJDtCURXtm8uJAdGtgqZDW/21LrPnvnHJ7/rKnz
OW/L9+k2ph9OZIEQ4I89bjaC3ng22XCDop63GrS1/1RpdBM1nrdvcIjgqnmYZ4++
syhvCXsE/u3lAcvSZNIC4mB+QD6W+DcZrqfgGtyJxGN+NaQBP9qzZ7CO2MlG70ko
5o0eWd5o4fqq4hj1wxyKnb2PrlX5kCU1rGpza9XlidDNWc2phbJ8PA0CWGxqR6Hv
JKBFhWobzpfZsKdMYShTHtosjJM1qs96xXR5FH6MsaZp3Be47cCz1OKrz4pYQzwL
vCGW/Hbmo1BiJa5nyQIHQ02Jmz83h7b4fDx5r5185gExXMzWbKZiw6iRHSQFHj3m
uVZGF+OxynyBDzeMkfWXD2+Xh5mXFI0V4076xuSmwCUYh0p3UWaJAI/vyFF2F1Je
gWQopgqHKqY1py9LrOD6tztbAs4Lk5VHJIUqX1QYuRPthuETmreqSWk1TO/DBXoN
rS1a/tSLnZNgFdXrtAjmrOtdrIUE6RCI3vMMtugJL5PVWBlNoReBKj72xORQQ6zS
A1yX7T/xx/z9TigdR6XgK7jdtBWxSqcKvuPGqYivpfdFEaa+g0J1FlFvCPLSQIey
3VJxhG/pEOXGAGL9WHiZ8T1XRjohjYcMdRzmimXv9lcuFW7/fBOm1pAUIqbWXncZ
vVgav1LpuqC/PC1NXoWI0I2ThG5xn2yZ5INR77oxTmuHjC5dL//jA5fbCDiMm0NY
jPTWlot3Ib/vUjAmXune0jXlMbADWgYaEEWUXwr57nBRCC4RHqFTV3A/uMlMsQXQ
9W1LQd9UgYfu+uCNRr444vCZ0auW6ESBvEu8UelYZ/kOGmSDfWjYd9bIx0/mBfJY
37GUC1/mw/tov4mO/KVX33XSa1OH5PyoovNofPRsDVtp7gMQRbCKmAth8hGuO4rY
AccX0//U+o48lpf/m8BsLhSzvnGAUYFpguEll5uCgN5OH+z3Z7+uYPh5jXcpUujj
k4VDhdw56iRpaLUVGSFpZPNtFzlk+EpR4NXYoaQqUUD01WT+1RJgJwsYGbdM4czF
8qPv2+fHw8Z4G+z0H2eq44sy7i6jGMFkgRCBM1j9ElwUBv5dWlvldH4V2mKuIAtD
aVI67ZmuG1FKgYDc5JpQL9oAoMIQ8DlV7mhcMc2aLqFs0VnqeSlbsPysQo/hrJmK
MH/W5Q3z0hqmNmpkOp9qyZ72K76xowPVPS+x24yvn/hABZmPCDPcTMbIBSVNimnp
xTvD7CCfZhCgtGxHYAQE25jVhgE7dLgVDz4U7A0LebBFCmHXHA3lPePUgSVP4jaw
TKO9rCw5t3wG3CN+ENN5TJdFYXnaEIQxU9aDbl7XQqJpZWe/jxGYzVwkPj1HhENk
87SVm0JlOAdLStqBZxfFDK0u3HHJTvrpLtxG8WVRmJB7eXydi/L+ESd6d5rRKEN8
Suv5vlY/uF3LZC28mapni+itLFsASIL5BXim6x+uOQsoa7QsN6NqHUP0QBGqW0qS
SFxbi6SnQA1OHqa4R86S6A3XS0C2jJLYkNjh0Ld7VJXMgdSABhdJUUnQY9xukgU4
0tNYl+wiUphugYubxBvZHhsfVsovcZyfm/LyMHkr9SlSj8wf/g4GPDn/SrPWOElg
d8SS+apIeEP00KQE8UBbs5ZH2QEoI5sGblL3/27AHfumsuCJJAmW/XqMHcQOL66m
mvVGWvCmXa9nJNBfF89Rtv/WxkU7dvg8NNOQoX35fVBjPXcFDh1Tq4BspCE3BG3E
q5sCg8JJ56ctX70TeZgIp/ZDqp+jImyigdffh253vMZbTiSqjOHBQjleR5jL672L
DYP5U41QI05hl0O+tGmxYdnbEZRkY27lscKyni1XGxDQsb1v+CoM6X2b/DmfuNfo
ZGMi0sQ0JSaiXWR1m57IPGq9mkxZsWSADmQZhggh8oH6RGj3vjHuTtCZbF3i7XTw
6a+XU0ggXuqNQDFUiGyXhF9HuGL0gh5pfs57WI8zZQANlgceu99mqtT71YEtgQAc
ckXHjvuP0T/NH3wROws0sQ4o/BN2OWd59pepN5Cj2/0uGsVBak3vlZ9X6zKRyZza
Oor+Y5nYijyujrC35JSGGcWpyw6+lTX1rREnNXQhgOFSmB/WLxTtpctTTiUmLGN6
lTCfOQLupSuKL6LQfaxEmjOMVe8w1L6KLWLBPM+LD9rmjqiV1tJAN5KLluW548Ki
f8NPXJ7eXqyd74XYxS2yLWTEv/csHehWmnTBXmrgGy19nzQXKImb4NDGOxdNd2rp
uZr0xQz9EBJgBpIqw1iERRwBDjYuYOA3Zxaj/W0hui64XyLJzIF+gQO7ENPPXzHt
5L0fOadxupNGyUcANE1uy2JLRHwv0fD8Osx5q2aC4gCeyvxmu69ZcYFjPMI6bbyQ
fske93TYnW+fAJobAlmwSOvPPQjpjEnMCMgcztOVOdwMvbpv0vL9eCIrKfJV0LUT
b9BA6jdLsProubaYbGxtAdZbCVEuPVuPUAUXi/QfDKrs+fExG/t5LNUG9qzOK8NK
rzMVsoHXuM4sfhbk1/h+dDxFHskHnS0QESZulLIuvhTj5cJW7ZBi253lx1x4quV+
K5NQauIcZcZcyxWxq3UqC1jJtgQcN15MnCET0xpbE23XhFK4CpCeM5dB2Od/Uiyc
OpdNcSSxkLyBbDcIJKysrYPLLrKsLjx/BzNzQQ2sezQigjt0+KEXtD/QmNQGnqnM
+j1aSVQAcMfxEgY2hWQWQNjA4ZyVFofG89eLYGzouorg/tINROj1Cb00hp40tf0A
RKKTTdUfKdovd/ojn9ebdwWn6lKuSHZRZf93iaA59sL+JDJXK9JVSPrij2GR0NYH
MhrAVOWVqenfB1PJkyI4svGAYia38b1lqKkPB1KKNmbC0L6FHdgKDOT5RQ8npgg1
tP32X/dm2ha7urMmegfAFTUPLB7EYuAUcxRi8EBBJW0xjSsl2+P7H+bhphwgeTD/
Hife4nOLvYahNOZEhmJiUgNJywYgVb2HSqbTQE9I80J5GjbcaSV8KwrNVrhWqKXK
QINUiQT/iWabfcBWh6zW3IQ5QTvnh+2RI19H9ErcxIYGlH6UhnHWq7vwXm1YrN1y
jbbIUxZQYEY7y0XoTzD/dxWm1pnssnzLa1a/RpolGUn112awSbkJMpXR6dd6KcUW
R6VizYc9Z75fthdi4oUbsD60ZseSIVrThbhCTfsBnkF5OjgT3fbo7aLST4p73sGR
fDKFhFK6atsFUjq4hW13hRvJKs3gNjAkQI940f3TVTuxl90vg7boMmHsb9/NkSYD
meo3XRrn5I5t84y4HeZbenPp7gB9DF9+qitewBwWM1g0M2xR4kjRy4bSzMuHRy7k
SkOPO6gYPQo4IgzEjSsysdfwsfvj6IVrzv7z8ESaRWFt+jNZgz/+NQ7JCFVQHADK
z450c7EHlccn+rpHE7gnqcikBz9uRgZVMVKj2Kryhn+UsFUnLm8YtZOe8I5kDh1V
qb2H/Zh8tuyW8UNd294nKbDZibTQV67DaCoaLBSFCqxomh6hIPb8R53kp4UZalyl
7G86QT6gSZIqpNjv+ElCR/7brcq8DOz7cLHCFP+glmMy4BP8q7D4ho99keIgLu/+
yPT2hQFqA006bHinYqPSkKrpRXrPbg18SW1igPZljK9BilcIOsUbQHK2hvFHvK3y
k/f0jaP1Rba3/tb8G30OIefD2Znil95IGToy+K8W6kd3YZ6dlk7R6PGPwDv6TGHB
iJ+6i1Hphpx0C/R9fbjOoNPk5T599/PaPAV6JdBpJ7aTSP0ExNmtCkksr7Lfz7Fc
NpnFPQZjBIfcwZSC60AG8m0W1GScZcyKqXfFbrBmYW6EEPiZdc2eD1s3XlDWfs4A
zw5ixv2I+xYIIuY1nPjChCHM35w14eq5b0uv0AFQ1AgnRy/92uC+A1C+CS04TGbn
3Sg/Noqwmi8JpNx2lvQJEAVpj4/F2zJQAK/BbBb5cc1JtgLxMJZxl7/j1/fydtTU
x2fUsRmeNDlm52jG7xJAaXC1e3avxzQKvnejT1RuKry07qCkhh4Bvm+KgglMLiSy
Ua9Z63uGrwYCRwJipRYIEluRTuVABYbXhpZEyzCHllYmRiJx/HwHvflkKF2vkmRS
fa+EmqLreoMq1bZ+2PQCFEnJfJ1joN2E3lR/nW4d/75cyJdr8vxQ5+D3DVyJtH1d
JTVgJY31gmOgkbF+mUB1nP5/6Wvp/KpBWj/1OUI5mAZYDrl3ajTNDUCWmoYDE0Fe
sPyyqwIZeqqUWTu729WkI+vyJt4Jn+HVvmq0OrOgaCvVA0HZ8R8lRACuAxL6rJfy
NV4t96hASiZbIfe7/2zSLT4V7MxBeAHR0+5/eM7sJU8uf8+MyX3Hl/sZ85yCtNwh
lzq0Lw/atYsvFaVWMobo6XCTvYRiawl1XjYBQunayF6xykWdKeMifTEU1q5vLlQw
+P8Q0ZzYKN9oVvAWVGsOaNj+ECj/I/5RjhNIr5cpRZqRrTTDMMIUx8IcOKc09r2s
qaUDO6XF8KuqMs5WeTYEaiGSVGKXeqru11ENdDzBvqAl3Awq5QS0Ec8GNY4ZD54T
ArtomOYUR+MbgLnZzYuQ0you958KP2gOQcMg7ORy5oHnRCE8HktSVXWzNJlCnh59
Kh2129wRPFO9D5yJjBhalP/4LmyEHcNl3sAndRS/LsJgXvMNzTSEtQqiMk5EW85E
tNZPOl7Wgl6csSZkfgQTjVmtKtT5Yep07vte37siaXC4Zjhc9tF87pEQBp0jFnqV
m9AOddIx/v2fjQi+5pTts4FuH76DMwwHJjd4wSIIjWUXcx8GY1Upj7/lFOhqjpgH
6JP2KbJl87WBoVPXSSLPGMfxrFM1EFhWw6LSw+FwN05GLzinIHrlaqq/7Obi5dpC
7JpyID6AZtTjEm1lBYCpLA7U2OC+gllJPzLs3ygiB0PIMc1mzn4/qH3On1tuYQRX
widMFHiXtjQ0b6d+cGbzSfPzxznREb1Sr5ggzYOPe7Q6pcquQwJ3W0h0hQAnyZpS
USIHVjPcx/53XXgW/N0n1sD8XGKEKqXcSVp+V5lhXmjZPJzXhBFIkz1TEhvBzbDM
GZ0vJkfmNCBo/EcRZGeYyLOY+YqMKNERjrgzqP0Q3TQ/xpU6q/Pl6wRbvMPfOyOK
Sss8LgAwyrieM88ZtsfcehpRuJ6rU37b05iSrFHY/T6/jmQqJIpXawPMA+9m4/rv
XkDsSNpYDjcSSJiGuxjBhuQyGl+Wbiwz+hFAAJX+2+ajEQHkoy2z5HudiFNox4Ck
7O65IxNlXsVU1anKzlliV5nXOlJcnB/9ARWj9bn1PPeWO/IOD0N5AakSTuoKakPf
KHxGsK7R4jmhdo0hM9ng9Hleria+oUAm6kNwXMhLjkBtU1KYuFNCMuGphTSSUkzv
leidHQb0dhWvUWlm30+Yq9NyMP6es9SPWqyxxxcswk+/tJT11FFt7Y98Mqgne5J4
sytwcvbJkfPbGXF/aGdb17es74HqVtSURyzSTJvxihMqz3s+SnQIDmIwnoc6z6c1
P0T+YW9r59pJqj1H4/q945rJt04K7zuZVsTxNURQwEkNnQEcJg61QtkDTUfsfLtF
TPxYO8lBLtnQKEY64oe5vD/NKv97DROP7yN48C2vciXPUvLU3gb8GpZaMAuaogRa
yU3SGiYEWWHDxtvVwQARwnXMvhLvwFZSnyeZDFiz5CuzpichHrqb5MWW4E3CgPhi
zA7NOzFASgOOmDlGOpQXqWvQJ+tKiz0SyFu+1Ie7x0q7o/TWo7K1FVYpKq1dxmbj
JK8S8fvig//Ce0sugvuFHpu7mAZVPyvrV8nXnBRg2IYptRkDy5ooWQGUj/inTg5G
txD/IwZdPtXk1kdGP2s6IcwrnRhLWp5r5kwcetAmSYPOCUiTKw5w3bZr61Ij0Eqg
/mkLy0CUCXEhwZ6d7/z4XusILbEaxkU26OXbMrMW936fvU6vC3GpU/bwgqotSN11
I3QwMlSVAnKFBQdBcC4KyFmaOQffGplmyRO0gizj3FQFJMUJeA3AIHOIJlcjxPCf
1T4GCfffJ67s2G2E8AZ3RBN18LEV3XGavlHbUe1OYUXxvdX7YlNrv0okZU2ivPsp
KJVRhbzhynaoAenJ5b7a4sz17rydQapg7djvZmPDYpep8hM/cOhufs3LIY6ziuyj
Lj/HlHfR/BEGpB50DKHotDF1Eul0yyjAdgvml1qBi5nBmHoGrq7ft6VtdqvxlpAJ
i8M83Lb10fzIBbyA9LQUSYAPSObyCtnJwhx9puq/RKfQyNefsSQJp1DQN50RoZUN
w2mKkqiywNKTvJce0uMkbNW0ZJTfEgwtujdQYBWX+zCWN9rUp35mpneZ40h/ZWuW
UCOSRR944koVqcVt1z9Fu0Ej17TxdkwYjJKylYlLiZTZGKs5g18Ykz2QtmqybKNE
UVJZ9y8BAtVV8aLxvyu/nK2B9koXpsmM6BkRUpaRE9R/PnG5s2oLTrR3ImtNpZoW
XHzK2r2RmFMk7kt1UM3OoEaXosXynSPfRqfokMBcNEUqZ9OTvCLP16s9LDvNqqZK
QmHzd1lEROtunDTm9gCC0wKKNX5xKqC7XBuzV0+Vtru6+58f4JME9N+cZolb0Wgj
LBH3+PzBF6wqxPppZqz+tFiIYKAaCFw+lHF0xpM6OB1EF9BnvamGrlykvWv3oSA5
wPXquJIF9B7BSqtMQ4wNLaHDMRNo+ehVgjUHXZMnOE5mO5cskFSaNE5V1BfGrYfR
n5qjtddZ7+Ok9yHyYzodRBg4YTusoVTNk2r4UmMOUQkaeVzSuQTxtH29FXJP/MBm
1bzuEfeDkSf5khFVGYogntSTduo4vIwJ5wsTmY02NlHJXMivZ3NvO5u6Y8YQ179l
0NIcTovK7ZonP+8Is20q+WjNDrZ3QQHLt7Cgcjc7+U2FQAI2asNgjv9YcRGRsPmZ
p5ZIzGtjcioBWW0AKMQDEJFRbrD4o6yDuoxIzBgxWBMHPl1o3IssSw+uLsVC/Gfg
cL8FypcX3Dgus6bEt2l9tVKNJdxnABUdAY10MR1JOkOkqegYVIT7wP+XD7pDkYkG
N+VCAfaHneuX7JzOQ4yOqrrZkwgG9pbj4z8HS8bR0BHeTb6H/wJXgpCxIq4rzpy3
mmwA7tmKJ8l4kqnEtHPdSbiO4IcvYXrW1B09h17x5sY0h8jiBwGOLphUXTSUwFDR
yO9yiPpeNqg4zjxnJCQAvZu+SXjtcLf9tFYBQPHCg483EF/55Kjc9BMeSEaqA/wF
cVMW6Y3To4PotfgAbakLlmwo6YT11ZKQIJkWIAuRygDGpMjQxnDb7/VWLhDcNDEo
Nx7rseCPzLncpiw71w7wLg3Pm5VlvuXTzwBfvD7x6lDoXJx63ClJtfpdhtfpA6Zs
oSSt3e+6WMAbUk9PRi6t3JgsyBwXNLhud9cGGLxu6gp1z2Xt51wINsCOyaww26j0
TsNBcrEfVKvUaT6BZvQxVFefQ8rZu0EATCF7lTrQGq11W0B0QIMMKhCQQXKrIPCg
5DjT4Dq8gQqQtePudROiATLYpwW7UKIJqnzEHF8PBq0g8vXnmXsoZhrg2i+yqPRm
ausDolZOD7RvdrvdGPMf/sTfuYvgf3f6I+UjQ/D8ZLvTydyHy3/7Ht2tBqOz34Pb
gbCWiWdfIJHNPydsBWksuCwjbdTfNAj5xjdFUNZhJNBTk/bBsd2QJ0tG+/1qSyI0
nGw/z27Lnsi1UIwQe933BqYC5DJA9fA4DxY5TwMWtkJNZSrR9LlIkCaHkeNzR1Bw
6XFsd+Aut9CmKeDt7lkPCtMZR8XfVg51piOJq11OR9wTPP5azM7FizkZqikwCFnb
8RcclVG7RlDciJ0sY9KLXRu2wOftTHzbSpQogKIhyBFLd+x6JYmXHG3LVswmufMB
IZEw9tGYgOFcznvOeXrOyCQvVlODQVYUWq3DlMp5mnmrOrXKd8W6gFbR5v0LOygG
LQA0FeM5jjHn9wlukOrAc8XR3eKchmJO2WePzwyHsUkYHqOzAYeHjr8DuwOqmvXY
702qpAUJ4Z4saEcqGHZ8LuLjageGiFawKl4VyQu8SBuTkgbTdsL0IMoHalOlvUlZ
m59ipLatlfketrbVtvHFDIrbdJGmss0XJZX6N3vwUZnc1xZec6F6WxO7+EuS8MT3
UucNSKkdiXPwS8mz4JV0OxCRQ/+pvHckYqcHSYS7t23j89YOk+I6vjzfBDqGGMaX
OQcoqjLqNkWp/tfSR9WETKJpkU+3D6KHRy2WIC3e+9dJ2cjxBBnSQMKeIgUCqCsw
dU9YXCoorBSgSEk8VtCGMBrL58UqZOYxNabhr+bnCAk/87frAJTmqH9K75F+yLLC
oXJkIwrh9dXY8yiFYwwZhrXlVkZk1cME2AdEDo2aEBXtNMiW9WAdlJpwenQ0WG5l
MHSzOkGyBjKFZLLn3HeFrgZkUA+KV/S5J4iSzKkc+uHEWK8Q3SB/nbnJGGO4ioCQ
Mqwp4y5/p3EXE6eQJlH2odfJU87z+3S6sECAFx1/jmlEgxyTa2XJibNg9fxTHuEC
jgtZWihL0oN1zxGxamVKnHLoOXwm2or/zpjISuY1Jd6mBOsPPfZ7DACKgskdWXKv
daqdrxygBIFzazD8H5A5PDvojOaOJtwhizjQ9adW1w2YIkEfdGuMRID8u6pAgVx2
1zNC2sYcO3XV75QK0q4bURs9I9DGQuP9FjnunEF7niTWfT+ZnhJX5PXNq0e4Wbq0
oB7xi2Hc1OmZKw5WsqU5KYNpsmXuWxZb4e4CyI88cTiSN/uqwjrNybADUqlKAG7t
vqFkJLpXpxn9JlMtTYQuuVHsws/kkZx1VIqm0ePiKwfwiyxdlaSKAtCxBo+lreSy
utGjVnjFBwjKxSUOB1ALU2F5VGvenH/yikBGUh24OlK8ZI4DyCMA6/afxrJ6SA5s
PtBcJgpC6c/unE23R1xARV8yBCiLHeau5fNVVbIcpcKT+z1LOLkxYKwZ6ZZ3oJcO
dYjIFflcHsFrFSRF8qDYsLj1E+L9R0X/lHwMaha8Q7UrBch3rXKIX4WLeMoniIxP
AKlug7heaZKwrNqu0WH9nK3bdlEa7JKDxBn7aoucxT6uxJN1qMLiaZnG0a0MX8o5
f4cgamJfd0PGir3cu8HviVnsZ5gRAiY3DcEX9roG3jwrqAxLhrdHUsjC+WOxkoIw
OOjIB9IXNHKYeFt1hJDJNZ9OsPm4AO+TtjIbmNej3VbdO5s7NUAC+YbuRmHOF86k
7L0shugXfYae/qZ/aEFeNJycRLWufyAfUgVroIiDh+piEYPNEpR3U4AwN303Ns8+
nhnFrQiMZ1ml2Z+m+J+j1ihPJOkgCG5thj6zAproZ4kFAQx0+yuqwdPGUHB2uDcY
SKrNZC/Bdpu4jmLxQaA1D6yHSWWmDY5OB9e7cQSm8Lek30UDznPPFk6eFbWahCTi
QBqs9gy1yQZMiX4s+P/CdbluCxfs/TiG2TNrGn/n/wtKXTIThwFC8bhOqu+BBiAg
yzFiFx4Jijzt6z71xnJCVEVFqjMgb99WlHrQPFG2DaRndmJAHSfpxWiPk1Z95Oi2
YLN9SRKSaSSnPMvUWJgD/bh2RjTW3aZwMI2KXakYFwl+ZwsvYmfG6NziBjsxuJyp
swQu4Znx4YKpF9sYsZhAFBd8FUZoWU2Ot666ZBQ5CJl+MuIFXhbpcmYj8+zUTcl9
8ZPEu3qhs75s92o4tY2ANkyLbXWC7jM0xM1YRHZqhx5r2G8DEFDQl1R8BDCVP9l8
EMTTfK6VVi8QYaOXB+QbqYm/rZBqNgZbxU/Yj/1yZVRT1RMSdPtP2eh6F2NuS1Np
rI4CHJXnzKwhjCeeM312TzZSPkBOj9kIATzzmJ7Oj0SoBbH04yC13hXaWKjhwXGE
L86jQqH+oPsffi3x+iXPb5ohnQXm5Udv4kDeks87iZkhod4alXs1OtThwhq8Jj2a
rbwcqU6A4wqyv+6POrOvbp7ym71jh6lKDqeGpTUWv5DaAOZv7Hq69NORPJ3/gyUF
l+TEAx4NIg33FhJL98Wlp5mXa9x9DKdqMNW8qYYVD1pNPmkK4zucGOzOrjjibkBy
acBAqYAlougCVVwFm+d2Wmf4pWU9RtLXRhPVSoRmgAUvgMIYwwFr/9/li/gDTs3h
0Gsrqh6fECTg96bKH8gcBj4+5um4eSqhjdWUVgbyUDQGt/R40D70n1T9Rln/rUKs
lh5/kaYYHWzaTTorxCuWSrWzvLJB/NqaXT4kIVPfrWXJHOaqdfMyadEN/As/viAv
I2BLLMG6sEliQc0hRSHBnCQGn9yK7gm4ONo7ABGOX4Jm4sSzbBZte5ytJH4irDV0
yU0OekOmsM7sGC2iQlTtdsi8CxMtN/oRcFMHG4SEwR0hWfGBq+XLcZ39gJvFui5y
zuMuKF3gGONI7thkywwn64abhZP+sy/coxOBUuGDuPTEXjwy43ZM05Lv4zGatIC5
ZXlsUHQOGJ4mJZgVzGg+N88jPWjRa26KfUmTLgLvT0n2yu+CtCSKKJeeVpMtV0uV
Rx5Lm6OHIDUZl+H9pWvuLOsM6obSbPO2QCa2dj6j4XT68GmCXWHxkM7yOS06z+ig
TpOAUMKIZm4YgBs585iiohPbjGGf8v6g2wZ6wDDMZXwxSRlowgvrApK+DyiRo64r
Ls2Yap2aOTh9yBLnRUs7O6vlDWrc6X+S86UueEy2YPG6Qm0iqDS8x9AWqOGaBsvc
VNJIjd/71Gy9HncGs62SCCn0368qG4DDLrMST5nKRQdRhnW9bKn6uG7Ij/ek0nRl
7D+SZzV2JGoVqSzXMV7aGuzlAK/uYYlqUk9tNwfeqz5SqxhIA0tmo6OI2WHymWWj
CfbMBkU8pi+ny6S+g4kw2D6bYs4LnUfDteB/s1N9ANpt9kiEiv2ndwusyMRLSYDd
fzZm8aLSZU83pfhSxhBF7rrrQqLoGU2Aybei8tTokZt+qS0RW1rIJBvWN/I9fSCg
/rYDY+SyiLFr4qC8GIY6sPESEHmMnbd8qGw4tNfaRL4uDDxpLDsLBlV7K7KqQbw1
mNWKZ2nHDMmK6khaiA1j687X7FfyE+BJsMIgD95wFwnnObgmD6UKMy34v3T5G6k3
x/le5af7720oUhIvt7Hqk8cbZVT6jISCcCRWbneB2+HhL9mhrGiempxEvkvl7ALi
cWvsXlaq1dApZ+gJNgH8e2str5LUrlWqsBicZUWNmSpB6qFwxCyXbNTUEIxpFmDT
12NLqh7qjLtYFxWlmdUgblzIP7oziTA/lwnJyDUx6uqIzozg0bz+BmU0ZKLrDVTV
Ql/piT1JgRQmEhSyvMOJBruN9onoRRL4vk9j7g9nP/GJUx/Unofevq28f27O8kvl
wC2dfeooPHvZxGiJq01hJVnv/nteQUJQ+wJa6whEWFb0x4XsdMLsABc8UqkC3F+s
a7hKUXj9w7qZPEgfcdSQUWVAlQT/XMZ178APvzQMRIK/SHVzWoV93vmP6e4N7xgy
I2V44Veh4sPWSX+OcL8/l5j/XL59AYN/JZ2Yc+l3QWr2/qYLcczCFhqciHhNuspi
G7Ii75F1PVG4zuJH6ne9d4QOraw0Qpm7oiLPckg+filttMXwWektQij4IOabzkwC
gHw+IeGazVsWgegeHJNz6qr9n/rQoGZyt4j5ndSErQiAB816UPxgcgpV3j5h6Rf7
D3DgvDUok+O38TEtw8YSZ+qvCQBwV93TWMFbD7j2tCx/zpsOzztWK0yXVKri7qUP
cxUOgmPgZFvhbb154xkkWb3iv4Bi3KkNwg20q4C0XPY0noU2dn0be52HY7kTPWdq
SQ4BtC/o13yrSmfDWwE1HKoOQVR9fVNj2/1EapYXQQbbdLhgU+/RSiDNpgdIWO81
VZ2ww+U2XCFyY8I5+8WWB/RPQSfVbR3zO3KnCduhdMdUf0sr6Zf2e8LHPd4iYhKH
ALzEjkPPPKS5Yg6AJfRVuPpTa46isqNoL6ZypSqayMjxaY8+5YfuvLQDNvUSLSJX
csfVPBE2A32WFUg8G3jh68slqV6biBzmm8gKZaFujXT1UYZRRg5oGEHjBAUfhOQX
1aPohFbREG6YaQLh2xyTKCA+hvaBCtC6uhuztJexnMkYm5ihP3WqK+o3oafHRgJO
+FgG8Elq+N6v0p5eaEaUF2tw4736dG7deQpwYCGEdXShRiBR3kobYBKbNINnuMEo
/P5pmPpkhI62YjnUV19j+89tdNL3LWfAIB9Y3wstiQb43ceOl+FwFLcc8PnF31Vh
DhVD7CBgsaRs2y/37B4AV+rutAybkNegGfzQro/3RJvQwSimR0Lw46WbPVjOtekp
uMqom0w58MpeU8RbH+abd75lEHZqU/ZzB0vgFdupMeyIu32QlJABkNW/aVeOj4Mv
EYHBrveZtwNhS7DFZ9toqpxrrA87AOZN3Xq3HjovPVtpR7rjlZ03e6QH9xp1TKH0
wDrgBTMjXBrROenC46eCKelQNVkQS5XzcoEWQcoWumYmjrhBZANv3rrmo4o3FJQI
gcb0bZe0aUryajY/xoIBxOoLN9MPnP/QyuudqUqeATBUHLFjFaraQvSWyhajEQ6a
qq7jJBwotbm1t7/eLXEbmy31tYpg7XjA0/GrYi2YgpFz0lvqsDr9L4PDzfeJqLZm
+ExKQMv6T7wmUo3DDttnpwAb/1p1fWczuzzSdbMqhLvirP2ppRu+t4RyECquuIq/
gU3UV2LRftjmHhghzIgEXzsm3KUuLQLViYjcDYTcvXbgsTR3+uOLqVB5ppnjvJOz
ZJGFZjiE0TsqVQFcxiDKnMaX8hjoi71VByFk8/T+R5kz/HICJWYIz9qhZRFx4lpG
6FM+u9TXJqdHRYnBcF6+p48v6OjsoMuyPSCO8OFzWmvtfROaAeJzkk5IbXEeLsSp
2nKQfvAoBOg27o1dsVuzMV7jbaD1qKugPOhZCo+DaoJ0Dd2995+BRueHZzFaHvG6
Bb9u6z6a8903QUqNLKKWBCWnRW8sBTMQLEyojgUgU/DoFJcQaTlxux0W84BtdiZw
4lSpuFAoyMkvyYg/Wk9VhnDPxABldfgbof4irtKrCznYi9hRVLguZvKJ71X0C2RB
MMIZP0+zIWrY+IEipprUdO+dYEHxztUUqWhJfuIKdtqPcCjzLzoCsmPOZw7ttrxG
xDB4ptbfQND6Z/25xb0/LGz2isEPtdfPsablsfly3wyt2/VKAG1GM1Es8G74Kig9
A+ED1MHfE0Qij1Bv+VtoZXkntRkmMOG3FUxfNJRNc+CpuagfjrY3gfX3Gyw8sZae
Hv/LCAEgef1rPxBkLjP2e/veGZBi3U90Dv7HnIdTuVRUtBjS5EzQjtWYFkcuX3DN
1SwI3M5jK2R6VPQyqEUgaD2Ehs1ONO89tycf6YjKR7t9HY7i2D4O+BScKLbQpBMp
1RaN0KK8sUopesrbeN6vnJ6hUSZ1LICftSJVg5K1KRCVcEtawwhFaT81PdMidDfA
iOLhIBaFsDa5wFWjn5y7DnsrCfmWzFGBgCXZy33qAFW4S5vnMgG0lfLQc7eim3fo
RR7b/DoGKGej0uaX2b1n2S3AWwkmatnR2xeo31AcDE8R18Fggc7o2YvVBi5KFRwN
mQXKKTd1UbH3S4m2AqDA0xyTLMUucbd9O39v254oNA7leF8TcwIUGoZ7wt473Ffd
nbVZ1px1/3o22GJ60XJjRdm5ddnB44IBeZAbPAIxC9CzbyFv+KyPeeGvUtMM/jaB
9bXm7sLHDvTWBGIQvSdBbx7Qk48prti5uZ0tDKpIAFWjLF9zjz7hY5L3E34yNE+I
T2VfoXUfvIE2Y+9VM6LYkLclVj5cnlR7D1CwxRfZG8/QgW2hjdyVeREIBhkurltl
eF4YMMOBtD1mhAJUYxo9isSDMgpiGjr6nikG6/EWS8nq7rVbPM0+mtUq6+u+kWBI
Ugus6Xt1+oKcFNuUJCC8c98HKfPBLm01k/kLR5KTzJw5+/b4lY6JjPKqbk5ons4L
1H7stI5f4wPQA24djNVNiUbXfV3z661bLs0vPWQjHlrW2CQLRO8GHQdcalZaFtXL
vwHtptRk6hXiKS79Ttw2Bif8t8AmyfgkIcc9BAZj9HC6BL9R37NnFiND4qNpaJWt
w3QQTTOtXDADRyD0KdJ9f/LAN4xc60CToVNsptF7idEllgHTBNztl/pfFNxUo+fa
vq5HDJwI/tLi2XyVJ1lipldeKOx/utPLCVqTGX25lZIGUX3BNs0U53B53F1HdvFQ
x5JX8RezgZRwMEkHCY81eY6bPAqwGJu98LmrJxVPDYM7aXniXdB+c889mXyq/AYh
FVwdZZtxcQ57ZKMSUr7XFzjTLMw9MB0wY3+eqAgXlxUKEpPfKZ7+8q5errOtFzwP
7MPgvLEnUpXmYZSC2VOHwmody5GPlBr8hMNWbcthdVNbrcmoYC9gopcq+l0C6mQN
ObsAvf6PWvmWQKTXU7S8EEyS6y3Lfhre0DjOiC53IPcf6zY//oljjMb53MSAiVCO
47LTvim9NFBNGyicZ4ySjsoz7iCYjVmlYIMK2Tocqd7vXZk0PuqbmmxDhCUfjP6Y
r34VS/mjhBnZcd0QimC51eFwDG5F4yfJRo4H28epuTITomvb8WZAVYxMBmyTjCwk
51u4j0JkLDwl8ptQF7I7e1n5aZP+k/J4FdPwFGb89ASWw0Yjh9DfbkTyjSc95Ffo
KfdjZPI1USJs8CKMZGwqMVpH44/XMJ/Q+nE3HPvlzYyd4Tymep3gpcE1SCefTFjT
7Hs4LAV4KR9TTk0Hwt8yQ/OAuCq5k3LK1hjVa93MQjokzwN/LDcbIbo938wbMjlx
bUVtWnLICap6OK6oHZkkPVKHA67mqUJTDVLXeB/avYAWs+IqtkVhf7wMpv9GMu6P
sj3JIyA9Fu5sKQX+9bZMzJVpRUXbwhwP6hnhuJ9fn5Jka1Jrftf1jDAvYx5Qi6FQ
WXqXA/b7RzcJLBLXKcSRfG/aNuNBqFIwklgMeBc2ilAYaCoiJr+9t9Sn3RImIzBz
e3pSKwV1h4RywyuzBd3KOQ5C6+cq9kUi2q+++sgZlD93KbPRSIidI4NDJ3iHF4Pd
bXHdGT0L6TtmzZxwhOjCdpMtc612uvHTY+RFMJrj1/zgbZMJcI8zucMawTTV04xg
l8+Eqrldfs2iXvvUdHWT/Z3OR1pIU2SdPC97YElpNBOQ7Z6lxJqjilMoVJ4hbW02
crpD1ywhVYXc31XIYy6KrNCsG9asp7yiGM7JJCgnzhztdzNZRi3MjmmM7WnJ6M7X
BmqkJ6wHHVVi3ATgoF67pnn4XVBcINs57nFQtWF8BVgVN4AujodZoV6u05xrMxgk
paasmMxGrR8gDTL78poSIUPYNpOO4pB6dN5eWxnt1nwvbxAYwEo/NQvJ7IXDANn9
CqcMZTeGqpc+JnOez2pqRAWtt9AKgoNqxIDCSbT2nt7Y07OWygBFoMIWBe4BBB+1
uGBw4EDPUAd0H63vlW5JoHpvqg29KjkKIuLnBSllNc8hYzO4a9ozHPxh29ln3Qks
dyV/NBXDVfCrdZ1QQRd8Mq3T2tZTBH9pSeA/yGIEwC2xBXqqnUbTUxSNiv3eybV6
KI7w0HodwtJ14lASnwZZob1uAzaFsBStJ33fgdYs+1MjeZ1n/1w+aeG12aEbf17q
2wAWuoK2NF2YQi8YCpafsIMXSG34LTflRjnB1hJ5lmGPyU1+JnKINw8sNnXRzA8g
g48vfnzrinT2JU803Q2qemyBpI7WNBpEjU6zT6RmmwQnpdU5a/+A78zoqrxv3/lO
CDJEyCmC+OK66H1DeVUUUsBUG5/Kl42aaCKv7EmJA+C5JxIOmcFnEUazzNlrmb8p
NeaV/ZBxNVBVKSOWDbkW2mMdPG4dOlQgPtnkCW2Bi3KKRywEh7KvU0XzkIZ72Ve1
ZVSpVwnv2Mdq+8HRrO/VEnTArbKOmLcatoShdYLzWQkZo/XPDqonU1itG72mQrAF
VcjOOcOgZRLj3vJbrduZPiwPlIay3ZvUqROmu6PDytspnaju6zpCiku0pprYZkzN
xzFwC1XBxxMC3GpVHCpXsoupkG48fN9pdWGQzsPkZxhGkzTK/Qh7zpycunMOEPKE
WCGJ1ShlRTQT734Ad6X44ADcuh1Uk88iUN702uw+Z/ln0T0TtK9kB3qamqwa7oaf
nOTJK8nKz+4RRhpEyIMwrEB0ykCja8GND3S/U4kfXvfNvHeWxERoWgCyruBYQ0V4
Yk/RU6XxTOlYQdJd8PN2BZ7uh/BADNsX2kSzOVwMOmQdqH8O0LdozSnYL5fIbWQ4
EYyat58+yavowxwwqIMWrjduBmr5NOhjQkfBgD3GfUXKFHVreNVgupCEab+BqLVB
4ic2ugMEurGDVHutfUasLhUPs57tlQp/CpYgu8CSZGS71rKPxwHxyVDPVvIoWIJI
87Fndu1wRklO1WuYphqgNMVYaKyXR/IZS0iLbukkG6wgXrjcUp2vQIllXQ88xPnM
6vVIYfGWcfGfwqCgbGbONmkHZuB26h9+GBgIp0b2DNfDm4H1o63fmu4UfaZOsMl+
rHp8HJdAcMcCQCd5nr0gAudcXCp8nqxJKMB/gDIgCqVj1cXz3igy0XwYZTsJZ733
cVVfcTSV1/clwST84OK/w4LoOq94veg9+74ry3DpyelYgzPZsrX8DYpsSPdoUP7I
3klz9NrrQba24H8U3duz2K2l32yJ/54iEwU3oOXOUIbJ27uLbJsIbsNfNTB8s5nT
9pu0d12EOwck3/+foV03sAIJQvdeZofjg5EujKq9LciP4DIrextF2rn5cNEjvszd
OCfVSV+0HkxKi9hGcJ/1OtFNPbK1PpqAFa3OQNIsW8VL1nvYjxAxWp3dXU1Kej45
Zu0lFkNOeZNTstHTyHgDdE2CN8Pft/cbHA9pFxkLDAwB2PkkK/NJS3dTTPBpPHDs
fEfOpPHiMRB0Dq1Anm/LImJ6K+C+H6k2kKIMl0J/wx7UYgAqAB08RjC1Sdq23qF/
aoflE1NyD204rh7oKDpPEgpb0dDvHeDo65zF29dFJpmiyOuJ31l3qQ1ZNL2et0kl
1r84Me9Ca7AqC986ysGQayRdnM/lPZ1qmxRGTd5mvsH3PcYvGLT0cfEfBCe2gAq8
IURo2a3QTM0mug4HjNEthIe9xXhoAlv64m9piC/yUoENYeIkq94emdposCnlk/jc
uyORT4LsOV82hHEGgbKB808D5r8y8BWyImgGvbqs2UIxDUiLyz/S3yQX8C3EHkgZ
QfaNL/vc08OVbrMz73ytxFJko06eOcmxdO1J9GbnNCj2hKNv4TWHY8491MWcChnM
td6J38LdAdGXneWxloxx+Mlq6gTVxlGdWLQCXJ70gmxEytC5AhwOriheiz/5JmKx
avsZrMH6l3dKMFqUKuEwisyOCPsmAKlnOgxI/xM35faPqEd3+zX7JBjNuNtvUbG+
k9s+eE64YhXkC1qpsNEknOIv0KGeilJDvHhKaGoaCiEfLiOzh+zTJQqjzFseHUok
IQdna6adLKtB4XGXX/ub7WFYcENDAYri1uGRqSSBXeKZcaebIPOBVs0f9jYsM3XG
wCCrsTj6FoOmy9CzEmoL+2xs86W9Pxo8gROJEv684+9aQIwByTtkV9TpNJ/8Q0GL
Cg5HPnoj3JJxavycHLctECemI0QvKyFyUxodDOjwQ7RG2uRx76e/w6oMX3K7/pCY
KiTZIZH/+fvfBW650m6mF7DhT/4H0s9RCyFAFN2BK9uOYD9S5Vy1rEwRzWOyI/p0
VJaRqLI0IhWlmTFKacWwdE77axIJpwYJGEnsGtkwUA+MlZTlpjCOjWrzY7qE3pGP
/RyBbtCQ1GpJTbZZg/7Z/d8z/2ZDBzEjJ6/5hevdTrJa1xE8x1RXILPPSTYhsH4D
5cTssPv+O3GFV5pzxYvCQCc8qgusS3GUmsEdFOtUWD/3+kQKzOqaby2ncr7+Qtom
M2owH4O1pTBhDPlBGYxKLtNEAzlr468NJQq4o59yiW82RMZyxnNa5aCJP0aeW2VJ
YyNytvCpqgilJRPdRniFKNzNcav+Kr3XrynsZvTyxD48O24H1tUFul/mE+LT9sLj
4PUMZtYOe3Ycxv2mzwL67T61kq8uHoFxFMTRH/j1YPNTFF4ttYei/Obku169orM2
YX783pniSR8XP9H8KL5utHd4JlPpY0aOvSQfI/tFRj7TGtmELYbXoum3mVxQizNC
YmdkFDjVXDl5UCmr1C0SrELLEVLrhDsoyzPeUH3Xb3B5vnYq9s+bbWClh6nas4Dg
eahWkrqsd8FNVIsTJyQWJ+zPYG7XJ/g5HvjEScihM5x/TYpT6xqTDtG8JxeLtnhB
kKsQX1q8Kb3l0BZPHcvQ5EXUoEpG/Z44dffVTXW6pBxgZjlKyT3M7yij+HQ42c8l
x1eJOGqJaUbQjnxIiIlaVqqMFOrHx3vBF2i/SYMhe4CscOy6xA7gOwQnVWaOgBYd
qUK4u2qRkc9TvnnqGeqJ7UGTQrPOVAxWaZIItBX04pVQQxhjpTMjfU7G7/JwjV7A
Jxgsx2RuVBdsekGx8l7L/Pw4hCdOoaCTXwrBHjHVXf+OVQBEViiF5/f440V1HBgc
bAe9CTYeEWeWQN/yO+hyoJAw2psx9ZpfAXz7gsC3uOOviARBHr4MCu6+jLDoU1BS
jF9VflrEbqqXhzs+PdpgAptD5Fwybi6A3yA9ZJ/fMoPDnhp7a2DdV3OFtZVSkJE+
fZ3I34pNeJOLCe0GiGawSAtpDWjrMGDYoHyhXHauj5sfWixzXgjtloFDSFTN4bV+
RU0ePnf1ig3Z0T7CVIlm8mu35T7nxpHb+lGsEiSD2BpIGS9UhugktgAGf2dhFZdZ
/fEsxeRUyncugNw+WOt8wsrpy4X8eD26nbX1zMwOq6Oii0C2AN5XpB+5RnCvjsi0
xy1z5htBWBngQUSq7Zcs4CVIRWkc0LvynDfxmEEq3XFK4Is3ef6vPUKE+JOfYWr+
7nAhNRKfXf7dlvRtaFRs+pEhYVkxcSNktNTcb93tRoJazJmScqbqu2baK1d5PQxs
6DdB6P5EfCBtkJNi3rf7u4JMAgTnh4KFNHAEvj9vULov/b6ny3SPKqVCWyiaZhJS
44/pz8hzHdvUO/DF9XmOaXVfMlz5gmFTmu812t++v+PHsY+Eo2Pxey6HNwsLjL+P
1vVyf/gOWWjd5vGIpSxSVMm4NrWLKvvi5lp0iXuEbvfGzLGI92mkVnzXnf4xzAk2
0CqHzPi2TOmm9eOujU8G4kvad2YgkfbmylHNa+/uRLiOptTwwbNLoZH3Kc7eZcwX
hxnhHHif3SDLbfPfuCJSTkFd1Ry+JpSOCqYCJInJSkR/oZM/7WirgS2g3RNsUQF/
e7r6IRWSDJi2oQOD9MOXopKeXMamnPCuFSaTCBELdmF93FuvyeU9qeG1VFO/77so
4TsTcwxzDx8yN6YK+iV1SetQGMquh5jqbaWXLVEXXt/RApPd63oFW/vkt1osFpco
xSX0CcHMAzCJsxmb/6kPI9TMZkelvawMdu6+ftAfYb+TDsntdRAuoxGcTE73I0Wt
rQoEO6qSHkCeNMMPfjNQ5rnxWYBIrLvArlpzqTM9OWZWUgKflJcGZj2+FC53a66r
KHDoast7QoE3xwRTGeFRC2vIgfx4svCll1P5Auc6MtotsWtyM9XsXyY061L0zhHj
S/jHqBGCFXelxzWEic/UOL4XXLx30hls58t/WM3dbZ8F2w2lwxriGgQYUGoPAed/
DoJbVIgn+UYeVPTJMo2Dd0OFJs8v2ziGOMr34L25RuTSVQBiYJcAL96N7tbzyE8r
nN/qqR9kcW25/Ok6JXixjhHCZ/WQxRAoeu01hLwy8GrQ4YqXNEa+5EPg/aHaqiqD
h4Zc5l+zI+PHS+/HVdteS44+XYLgJ2LdVW9HW28ovslQwpdGLyr+btcaH6vpSIA6
rVVsTz1/4Ahw4LLTtRTA2E2BIRZRKkcHNDM1UF8SgaVGunfMnPlkFvG+oOE9y+a7
B37cRmzqKDftypZZSlWEpH+XGYh8g6u4AQxgLM2UBMxw6jfbpNmXbJO8gPoZqO2F
IJYh59/dT48JJEKPTPbXw3jCKfl2Mq2jt6sIIIzMRpmjRgbkpMm45SmzVzUs0bW8
SeEl8Ja6rYiTmt78H15eZH7u95rkwnofloa1RYpw08nM5iv+bMGz/VJOHIOkHZTZ
ninVYkeVyTNKWays5ik+KHVckk4Uwv0H8t3t4noB45UTkxv+Qjh8b0hutdzZFQQl
RB4BJONCh4xmic06ViLv29eUdG0WYDa3mEKaYuc391Hxr1RteZnihPk8MRFqD3l1
XFlJDhUwPynmS8YxS09QkA0hXjU5FWC6OeFq9M68m8lc9fkg2g5Os4SVbgRtH01d
ATMfY5ESOTJJVy6q9z+FxzIfiRWokqNPlIfI3P3da2jRmuj//xbpkk6zsgxfJe/E
hprN/KUkKc6UwV/lVNtQm2slV/JH9ayYDFa5z/i+wPGF5vsnP3ubbQxegDQkwFcu
gCDN0qUwhgB7UPCyUNvh+q5Og69RCJsN5tLSc/CWkWuhhDNWNZaejQdj7Yuhu26J
rHfEMJZh9vSStx3Q0ETLNg8E+Rm88kwNfWf6K9qP+Gt7eflT5LZGW38aQXTzASM6
hwU0DLE4ED7EZhL6pazHWI0rZU/CdhWApnNtrIUY92oXj9cBNi+p6at41lTAD2G9
MzyK9b6gTjI5NFj9kr7M2g/6AAo1Fa6iWUo5pP06r7CKCAi9ikUzFxx8Xc1Smv1g
Nz2eHPLdunib76QjcL6ZiEmCxetPqhqrXSgjmdbxr6qoQ865dpYGJqm/26/YF2GE
qJle88f4o0XbbcdfUQEHY9e7hrHkyDL2JLrDvz4GDYPI4z7DFzfXt6tfW2mPlVwB
J40a4C5h7rlAivSdu5ow6zLUvDEvMtSE8pA1w+bIG7AjTRFCkXD5lun139JuUijX
1mlXpHn5os8s6kOJQeFx6RCm9rvjxdtNzVK5nFyUNs9uJKR7/4Cf27SXnUr3KQxE
6MB1pDm9Finl5hdtWxHushXC9jTYn2SfqhGLy7dT2zAt3wVoLGNty4aZRbmDRbF7
OhS2oLRvjlljVuCwRhEB5+xnOmwmOpHGfXhCKledcsfK0cgE+bjVicvKlIdB11Lh
mOnw5c++4Yx8FKxgJVp+ol9SjoAt9XH6bYl2GIvHsm1LTn7BL4VP6hwGHOVo0YEk
XkHpRyxkpNKEdC0fGRGTZEc0eCT5qK3bicGDU+RRKheDrBn0yPCNpva9CqslHi1l
b2BkZepBn/WUbq4L17JXPTewAGFYoBTzqMHXKmKSXZJOvU7Lo6QQ7d3BRh+hOtAF
ga4A32YOtA2BaEG20mxnTF8FZvY89RUlRfjipczpg5ke/Q5m11xN8ScwmJFjmV19
ZMKzoeptx2cNCVVaQ4sR9SvQVCxGciLp4UxWK2TmqcOMTqcOOJjislxgnLPY+SUN
kXPl23aQ8Sp0qrRu1Ab53VMzwy8jSnRLfW8MwDmbJwr/aNpPrdXVRvhbuCVb9bHp
inCNgIps7i5LgyZJkH6bllnFpqMmSZdYo/Zdrn9yE8QNRg1bmE2mg//ZDW/mp5Ug
uP7czLixsVfUkfpFfaPWP2BiDnZ9ALHoAVSGWA1yGCkmnnjL+Mt+OafJSfH64pMY
zD5P6mbmMYtEivLGkYhK8KTxHvyGNR/XiZSrPPPsIVMeVWU1YmWC+Ukjc1ue+6NN
5GAusc6IuEroSclAXH/HwOUwKxXhXn3t+zMpoWOReqxtMTxrYZh3jum2phCLa/nG
U75dTydcOhWLbHbsPrEaLQhBd8lAqKjseuVPMc4B+/Ksq6ChvCGGE8G5+PveFksn
pMa1GKwRF6vBnfH9jboKCVP9xIwSXu/wTfvk/EAnq16dJd0t76JVe+kruhx1fcAw
a0CQG9Cd2vGoo3RSarkFm6yzThnUV3rn7Fqo8zbl8Q/QYRMRjK1YaxmvIHDxutP2
+9G39vEfQBQMx0nIBGtTW0WdGx1a1SPneC5gjhdF1i6jAzL4t1zQwJXXLnkT9zIa
Pjt2CgcJpNSYcB56YbtcBsnk6fnaTkuwQsp0gMc2nl5BbJYlTmA9UyXcpPgxZaeY
vy2DQ1+jsU5oE9gTUZ79UA7GZlm9oFKTo64FuwpbDw5SCiabVQLMEDMfXpW+kKrD
Hvcy9kZes+YrEZbXr4v084y5wF6/5LMpJRyy3AZOJr7g5NpT90wybE8WdB/4Z/S5
2LfbjBPqVZPJc8vTxcFbLhZkTdB7Wba00oLTyIxZvlS8KgzJZezWgwWqzF93A+vJ
7jtT71swiG5+UDciT2MGLbynU4wYPfWMx67cEr4Sx3z0rQgVVAzS1X/CMIC0v/es
me/GLei8Pjj8L+CJUPdE177lEGAfnb9oSAg/bt7YrThmvvKRGlCJcKroJ+flpaHH
sWAq/qT2ay0LtadG5i2d07FvsmeS3hVModI+Rag4BsdCnqYA1s+TSnT/4k7T1Wt1
dpyiRkUjOvUCcvK3hBDmB5M8IR7bdTRVmXAtiDWdj3sghqFeI2MokvDBtiaY9RmB
FmdWCxYUiBOYa7qkXdZziOqTM7UZSDSOVFIfjraV21MSFKKKCR3Lg3hCizuOiR31
QCbzETV25Z10IUX5qNpPYI5LgQUfvipkOnxgUXyhsGrxjSsI5EA3sHnUwzLIlSe4
YhUTmfFV7qmMl4WxYqj3A3+7jbVJUOUuv7UpsslFBosjtUgTOF4OSHIxRjnbc1HA
QHP3IYW3uMR3EKb2DFfpka6Zl/8IVeJU/zsE8IG7tc7LTKYJHm6P7KcPIpXoxFQ2
b4KqMkQBWm0Sf8xiW1DoyUJvlA9YV/k0pTE8mgUL7tBawWwsIheOzNfw7rdYhHuY
cG5UONolv/K/CrycoYnTVWwNIJi5fAh1GHvrgsJ4LlvbdINdc2+hyMG9TM4qnGJ9
dUh/7EFxw4BUQefo43RjlnAjJWApDH89hkWVZ6zNSGE6QTHk8iIq5LjwuIeVyww/
tGi+TVMHW0lhxjf2mRcWep/7ZXtaqQp6c3G7Zq+Aa/Yr4nPBeQLA0c4n/hLv0rSk
7U4ItTOwkY5U/KfRDO+LDo/cdODVLJm88bFZQN+cE8kS7r6vwT89Ws2OAdrCNm+g
nXOtp3H66o9rcWLTxg2yfYfY4fkWk9t8lMLSw5awV+f1EwplDfOFvd8/lcE/W33x
TD1AUuCgLCi9xqpjBb3YxUgKHCW67UzQ0HO6XRprSV7r60vMPvptpox5FXYMocVj
B9LYxDjNREtwe6gA266zuryGItGt8DBLjjENqSJFWrNYGraVIJ1K9dQ+qIaLbMk1
2m2L8+gGkZ5RUc8YACX25jFU3nsoa8rbAScwNowOd79/AqaFmWg50bR+PmThiVsi
IF9VzwIzehUVmxD/RrgDETsFaTdoLVeKv888g/Zd0fknImJClu4tkTGiexiz6U6M
nIOSjH+1SVkx6esdQsM2rkhQ3sBX9JrgwbPrmbFjiO78XnmE8L9bPQhL0dzHwN8W
4WQWW1uRUyzT9U3QyR2pEQupBqK+82jxhlOQ5Apew7m/f3GNSO/g8GFpVziwlBW9
3farStozBzJRFueEEbygqo5huT3Bn6oGiKwDUP9DvJ8I+BYLE8rwlMxZJzsj2f/O
+0ipaTjInNZ1GVSVEfzkkvqUOXHyKJGhb4YkQjw+JfgugNB10CXQg/K4fP0NSnWc
JHd7doxPIuXpGb+a41SEgrs0uzEgaTsqo2GwdtQH/RRP2HoTyp8JoqJBmyEZ6XS/
uYhbT/FibWt89iRCIEi9fkN9iNV6owPnvl8jf44HSzxEmgcage1x3lZ5ERsJoxe8
3qyORDLAlP091KrZPa5ctNm8e5hi2eQ7Gkt91f+xk/XnykEhqiDGGPdA8j+oUqOI
jmfb5bwG8TUETGKJsFKnGOyr3VhP3b3aHEOKYiz583UDYC7hrpUC7+EDcUiLZDso
uOcv0V5a3EJj+M5WgDRW9MnAOFNxhlkBLz3ge6YHRfEBVqCJWO03ZDkDqOleQH+C
cR7E0E7L90yNZ8h/MNDZWpAMngGInYpxJNlIUiHnB92mIGfE592jBJ5mgrpJGjb/
Qn7du30Lk1azzYyIxVT9/HsjnU13yCiIaPgluquKZ4K26yEoD2PQATGAObn13CLC
zWQjrB92jZF2AYBmP41rMFXgrbcBzO51u3EOjwAXAhzxxM75b/1+IJDdO4FI5X5C
LI28ut1+k9Hz9XMglu7f1Atvk3LFFjBaKcjmQuBn/NTAnhnDbtxa3KI+UGr8byLY
hGXlPkt7Y438TJCYW6r0/ezrV29K6xyv+IiKZEV/s75n+0pz0Sjwc+ntYWAWjdgu
RvEF/g8dqRVnfwzvpsvq1lV74G04U/4YkYmUxNiXBSF6w4PLVVO515kcnbESBFDO
gLb4zNzak5r9xiAMgVvWUbezvu9vyaVdez4+JXeWge7eDAyyVg16JshPgQhTe4Ws
Wza3UlGRcLDmzgvJG7UUTyATEDtaUaU9gi8x6H7ACwwIrD9y8rq0hlklcvXW/NH1
jp3h4XMsN8lBuMVHRcOVUrxyLCEg7C4drllgq8GyhJY1OQx1D/imGQ/xDNEsw6xS
6sLOyROKObsQ+Fw96TjSCl2OI1gAx2KYodUHFACNfXGuIw7S4KJ3rsoFH0LbU5AW
yASIQinJqmDF5MpSHOECErUIG1KAsCaIX+71gOxytfk6bFBpyHKUqZoQHaYaEqmY
I6Y0BYSMO4b/lDUJVRYGclet/L9vI9xvFgCOG9AfqBGaeqds96htRGkcn62C7x8v
U7BdxJStAYSZJyeExSt43ge6HOPgABp77xUj61sWuI446F/OPPog8LhOZ0zG1y2U
R9NmAUsJlkEZPYLUr8+Y65dq4XGTkAT1xPvnMtF2mwSMfxFiGvGiCAsCiLZIvAWA
bwd06MWoR47LSBf97hgtor5PkC5nhkDGvWG1H7Jk+0tdqme7UtQ1HOL0J+eYiovW
bxwLdzclVuvL0i/r/cXKenN7o39l2VYkMCbxjPrYXCBUxsErkpEaAyQyWDbjeNht
iBamQQ2vUek2AsVdGHBXSUN5C0Rfa8LT4ez7SkIlPJNOgNwfFs13iHH5TaF63sfE
3qzd2rUe5+xI4LUYoAKx7w70PHcywnz2CqFUfZoLqMJQYIACsgGJ9cZ0+yP1CZRl
ezQDPSDDlpxpS1nOh8HdAhLfBr46+t2Ja/yHUETIPJcHwQRY31cUkjvmWs1sGPOW
eV8Cm8ePxHXcftbU3bUC051vInyVmM9AmBGTKLPlu0q99wFoZwohpA+Sjb+JjFfq
dfYgVyin6RNaMghAP4u/a2FkPE5AQY1SWL5K2QsBxQp3jWMv/fsLOns3SsTMmT8n
/1yYKCFCNP3IqoxRJ+y/RLr2HiXAb5icZWz3lHwwl9j1M3ykire3Nin5MfA1Pa7h
77tAnbmiGE6VpV6j2T9ZDpa2Y/+DdMVH3rS498jfZjs/QL5PRyPJoXGK1GLSdtLW
cGa1NoRXrp2OF+haqPaFC/MSaGJRkL5p0NL/q1zZHvgxltboNA0JbGxS/UCbLYVv
th09QH1WT+LGCfmwnxmnxRxGrGHw19vDnWindJteYdzxK5ZuHW4RfRnXXJ0+XPph
E+iMuAYHaVw0OaIRjmDy9mJ1TJIkriFEk+z2qCU2vKUIwxkH92mIlnQC6WmrKQif
C7xx6FOT25K6/rXnzspLwofihE0O4S9FxubcZcb1uwcgi7dIY+XI0i1grUeytxAv
Bm3Ow51wR+FAM5rc8ffosyhdchTwDZNQsuBNFnzh0Ue0FPPIJLzlrC+9QoaUP6x+
sfjkLgNtXfckMQpbPXQdNYiTmu9VGfYhHfCQNeTrlsmSWxUiKXrcVTtiDnL4ZtQm
Ec06P77pWRwEb/lAsUTZzHCNq3cf9EbWeseJ5jNld0rcmyz8RkW2SqATfK23u+BW
SWtsFTfttXhzwCbWP1QSGSBPShhqBempuCI5Rrnx4OKh9vqWhf0uFPDuPbIUr9ow
XnFUMTQsJXVNI6j/zmk9HyNUGVx3GcNSM45a8pZTuRfwNp1Adw6TyqHqMj5VkeiN
+Wo5AVh8XS0aQLlF7FE6N7fzfLsC6/tdFfUCgKea84e1m6a7yyIqKKpTR9pVT6FB
UTUEFyzn3CyWdjeckct/QS8Of/BWj5RwgN70n21ksfzhUW5szZqW1tBVhGvjyPea
/M4LxGWFNWdhSRA0PUgAPbGbx2JbH+jinvL42vBJBr9ugjby+jsOO7JdWKSblmZr
09H7g1/roWO8+UuKXzCvh873KgnxMSCoMK1ZMKBa/Imiep0LQD+z6NqqyvTCw9jd
D3AFJuG51aNrz+5O8DYK4AxjVk1ww2KYIngtT7ujXpdNtPDUU2wSC/sDKIrhBjsl
G6bSCU+ZnXmXh5VPKrg+7vss3ApRCJHy1kOPovBJxgufMY9CxquIpQHtxx3FMsmE
IFRXOWiro9dQVHCsxhYE8Bc0Bpclp2hUIoqEASphUF7MvY0zyAdae2+1OuTxcoZZ
6RuJXSKLpzv6V6IvB1qaLppzrbdy7DAAh7zhzunpVjFPbYty7MKScq+NAbHHgCs1
QEFua03rblZRdqRrIeOL089Wr5GQeBKmLAWwCPVwZ1MaYB/5Mn8BGNtSE2IblJcl
PvVD16ZSn4Q6S8lyJkx9kFdpel204aAjXPeRY3h0MkjvcwtGKmrOi22Ehz94DGzs
tV5cXyZkkreFd1euiEDUPA2ip7e8S+JDiqNGUXcDvc1hr40zViFSYzEU3YiPKxsh
QjobpfymYr0eu1HV/CntxneKwEm0HjlLME2MCGRd0MllIlprWrzgNfii+Hk3s8DZ
rE5/YnagsiNIw37d8qorRvZiAXIQ1pu2H1WVIvgsqG8Pl6Z3ZHaRyb55hY79HTOr
7EdHHmbUuY+1NYpWemvJuDdgSBmzSwP50MOpM7QsUW/RxlHbotcU+KJrF+BPxnxT
86hBm41e4UQk6wJjuQDE5QGClfLaWiLpvmYxaD5uvMnqPUrsbbIAnA/bpw1W3C4W
egKDNiACMzDZQIgmXk9c+Vulbnlj4/8zFEuYMHpnXMnVVn2ZGmXYXioMz2Whj5d1
sq40Bh8icwiHVySprMwfrlqGDHh3qJ7iIJENY+kYhCpu6weei4rjkdmpI36/HFqR
q7ZlROoaQRWAXbgRr8/VDWVqeYCuyAqpS/TRIlaLSDHzJmSSyfaVquB3ad2p9iZ5
HN6q35DkAXEeRjIJdP8X9c3EZygR7hjWS2NNhg+6hI+5IrsdLyYtgPQZSSVC2wo1
87xaCHrx5qXype2bdGgnuj4QzUufPMTIMQvshZbL51shoHoPtHXp5KZJ5ruUXELz
SyCBzyAjiVH5M5vnCqCzLTNK0BYe5cVAEMl0Hc5qs8PzAWMRSAOQywGofuC/zFqV
1e6lTdCj/eTaE5+kTdZpevrI/Tjm4mylNJWnl+ikkcm039xLiDk8t6hbGndizH9X
gXFQFpRFA3uTVeRixuygYKOsDQM6bn4s8XosB9a5YfDtUgZUSvc+4lHdxOgYoQrB
TS/K1DMokeTZQDpOZ3K7cc3su8Ryli4D0wE3mvJyObhPZdihUY6+8+IJpitKeY44
kx0P7Zgavn3VVugoitacAWvOVds7a8cRB7YXMtdC7tzhrAs5ofkSWui5H01IsKTb
nnB42bzurKklfvCpL869Rt0S+8Itn6cELgPglDgSn6PSsSSLesk6XZaD6Lo4Wg1i
sUKaCX6+RNkEGEcgmeXszfl2utu/V11ypE+GwwKBGXjTH7H81HyOvYkkIz552wl6
HWKFJn1QsdMY16282IGkr4g7KoRZnxRfisN6NHAUsBqsTWZtzV544cJPMyaUBVt+
DvnGYWeZQYBrgWDjHAAr1e/KDzqWKIaLR+o3i/Umz6Vg92mCd2KT6ANOMFBvOsol
abxWls7D/1pqlzIS7N2Qs9uu40DrG2cw/UMGRfCZ7+fr+MBRl8ElTdeRWdWxTppW
hshc0Mjv0FAlI70HW0Rr3qUokMLkxcXpVtSMaWUF8PTicDYpiCV9E9w6byRHO1IN
gi1CR0texsUGmp8bvQc9mZzTN4WtQ5Tik9nMz1eZHu53emvSNrtJRs6PLNR1Wb4T
gLWU6AwcJUK19ni4IhT8p0TFe99TH9sVcv088T5m9Tx5IgUdSSIJRcS80Z+vMiMe
blJZASRk8RQSxz6nZY2AIh7KMsYCLKFyjlOEAdkWTRmp5C+Ob3C89xyu7vUsyI8j
OvG6DSN+hQNg6MVbFHUGO4+HL4pldzj/DhfJ9jgxznzrLIMb15iA+9p9WkRJBJcu
dj8rrhOfrn7spgWgE9ZmCQgH/URP0VOX6aToc/NWtHE5pL4uXGx7M04o2Xzn94rD
FP7TvyehcgWJORNUgDfHagPtawwH828Vvx/6WNSub7XdNMVfwz2Osy3Z0RFLbR3I
ihHdGtJW5ilQX5m3NFCRQxj8QEgwh6Ak9Ruy5JN0o60fHa0L/FLcE8rRTHcZaSRm
/G6lwXiPcpDe8MJ752Avj6HztGyjgLM1saQolLyFciSCoq1pD45z+pC8bPQWSOe9
miw8CyS3YvlFwwyaAdQkEB659eM8AYFCWJnB4SwmTr8F09XfmMOqlkLDmMSUgRIf
jfnzHz8azyUey9C1OeIij/ybry4ptpC25s8NqtfFdccNoYKSXmC85ncAiMduPpMC
qRs8u2DXv56PVktSceybeE2QwIF4rr87rzGrYvHKcaN54Rr/6I+mHLpHtOxjC7QV
rle58XEYWwsLQ97FSdcfgFgtLntQL0fqKoqLC9XZHpS6i3dzI6Y+V4X62I51uKrI
Tzgq+EOZnzVKy2DgDjMENIWNz+NRpBlxuN0LmpY61QJp1/5sXamQAaPZxZaSK5vX
J7yN7ZemUxLymzMROudQ7wa/ZAPTNazIM9TyW3ErDA2Xodzzn1LEf0IO2xQ4DQ4F
vNSu3wip7gtoP4rszYoBqiEQ2GQFyaveeW/IADPje6Vf52GmxpneKHQhx5AyTIC6
IrJcbEvBl7K+/b9EvJN5d3zPiPRFKjLVAMjP+Pzk499hp43UhkgjAuwTedOCY7nu
dW4bjtlrB0EG3yAfzkKdQ5vv7dRfi6YyXb7f/Rg8BDKstTH2dUq/4Z/YzMP64ASs
OXcmzAq8Tau688IXZyIQ3ldJwzn27v5/skQFmKz59kEJhlmyBCgwMmk9CnkUY1HO
J5VeTkKtQI5WJCX6WELMIfFY/xHHOF94+IaB9xT+ylc8kOSFnmnXgNHQ2+0KLtmw
sbbZSx/mSqkFklorM+hVZlXKQt5uq2B46gX15IIR1bRaShmXsj0ZoWWrUF3oFqAB
9W+qQZpXVEcOPfnPFp29ALByPA9mMxh+3NJrws6wG7eTu1KelFG7UX0mcOXdg0fk
9lO5NH6mxS0l31/6jOhCTLT6qAwgB1j1i2EvMuzGx6YueaLbsJbh5QpJ2xXGhQ9w
qu+FNFeC5ndDW2NktvCQepV4nTxVhaOfleXSuhUp3rSzqS+FAoByqT/VWDewUwnt
+Kj3woEu3JTwX83cQwvUdP5WxuKed6XoE72mXXpeZUK/JFZ5eE3WV7Vm4b6FD6t5
qD2t4CKLtlUqqQ4cR0DUgHQpzmpRUINkgx5zcQAAqDKjuDbvcOLpAbWoCC7x48+J
JgIR4gFzD3Id294EPVfqITNNiSKWWXDU9S4WWbmtaMQjHPOGLEpBS0qIvWZb7HGS
Ti6Jnmhh+ZVDTItztVmpQR98HKPRASuzRT5gofaNX1hEMgPdiQvAFV3QCffCBtpD
OWkJcg1vgc02CLLPm9e5oihEDtvLrezoFxyqlNtTMwsvRk/m+ajIojRUvfb/J4wy
BGEEAurFcpvspTCYZWtMY4tcrQHOZ5j/ESj+Ey7WctBgWGTEM+t97hvncSzpByfx
bBhueAeeDNpeVMY6hak4P0cOuNBfC7m0UKXSNau746xkMDbr1Yq2mfmQk/bcs3Fk
F+q1xoezRQbcXCd5dxPTQJyL/w0bzjK8jDqXgz4luw6NzHVFHPaESO00F9A204bZ
VdwsOTVUdkwmtW0ofN10pR7MZUPb9vj8FKJRqcz0ChGqPFTvt7RX030N6BsjaWnC
sdqTXog7qYvXrSwBTtXEqTMgq8Ey2pIHTwGlv1G0dGsSuZGPTRqMCkr+ecPbUb6K
wUomZste0Zw/kF7vHqYXwL+yt6FRAxkusXPwkU1rl67tsaiSU66wTav2ZGrEl6Kr
7gfUZsfyhfI22Yq1dmChiFftpkZshUoQtnPNd/VQlnLTohZNZbZGbShB12ck2uwH
D5KUKWN2zeiZ4rBbQk98CItiwMVajR9JuE7cKsPsIOfa7tpCfpkEQtXeNcjklh+Y
xw5mYnBh6jqze1b/emI+el8jXnJ6oAR/Y+4WvzufO+mKye48J9SSkecDgAnnGJQN
8ZfOT6E/vw/cGTrcvLGUOpk6mgph2OdUKhlEaTYqGOi+1cvqsjdRX4+QxVxLJgZz
GCvrhA8fwgjrLsNX1he/I4G90woT0+loA1CzuG3sOoNN9RG2oCYtXpCB1Mw4JzgA
vaF4i7Whnn56I60gF6M7YLfhTouXiYT39LpEILL8ZW7+JFy4EyoDEOiDwikWVsBF
5Q3baVgIKJc5sMT+izN6dZyxBRtPFV2hTe//1PT/e2FJbBXPFpGq+hbnga+jE1GH
wHNHiDs4dk4RdCFnkP25xAoXEud0bXHmHBv48+1YMhoqjNY5wry3CTgQCzNGjwZU
EKifcxgjkJuczWhbhDP7/zl7jH54kic7y6sahYN6PsN/t8UnmYri80mYBLlTjHjZ
4aO7YQxtW4xttORtZci1lcLzBuQkzev4zVUDYnQEl9ifgolpo2ixM+KVN9ydpYtI
zl6jvVmxV0SPKbVt+NxnJExrM06cuzhA651S5w89P50U4W0HYIofLEycvb4eY/Iu
L0DsRAXPlvNbmxj4wgTTF7+CLjmultvOfxthfAo8yyHJ8JN3WupCVL3VNTwmvRTk
3lIZJHnbWr0B3SEdBvZf7wAvB1NoHuTIwlg0FSEmMvN9Ip4c2t/hoR/8IFLNGO4l
GEH+4VCQULTOqTtLQCwb1XApjai3kjkimnGcPyrd6qGwBGswkG53w0xZSgE2Lyl4
lC8r5QTIH/71o+LZ/b/CMxzwRGRkC1kKdOEX4NN2mrcmk2/QkaCMSzrgHYk0uaEl
v5+kxfQKGyrh51sakqt/nIgEkPhLUqiHYP51PPF1EkGZgeRkp+pw5T9yBvlSuDYz
UFUpQcoQnC0vT4kn6lDAmmpv7HB6ioqjCXMfyxK5hG4CK8vV0CRAY6UXRfKODmJY
GLJmkMXy/v859JiX6148ZPPSayP8mHB1n8ntZOO8yT2tdak7lpMXaM3zs8is/1nn
CsBTUG6AlTmxbMlZcdnzsZp1d/7mqsQIzQsStDLg720fWWWpeAzsMPBfG7NSmO+6
ftbwbfV937W+xLRSVhgqNxAeU/LZe6Tns11W7XNxNvqlqy3ujoVpVb69Xemtr/oG
g6+Bn0QUHCoZjdSHCgoOemz7o6TQogj4WFuTp70vSyMV6KVGfuzjL0xWp1cZKlID
1G/9wBVehW39gP2U60DPoKfFfzEgmeXZW8D2Po2d6+mONYdNZNW9pMFGGzIV4DgE
MAWfreT4qwTTLv4698z8TLnl5VoVpI1tfjU9q3GtYnfNaO1C1z8X8tTo14Qmt+Be
NJCppKYjHXDNKRSVBP1C3+YKNMKvv4uyc3Ppyz/eqdbkz5UsnhwBiZKEiZRn5U9P
XrYCKnnGp9Uj7SE7YFH7VnhiGGvR3UClQtgGgUmdbRP/ds3XgLuxRT3gTZFJXITV
n1ZIp6FAG5B9UhIpHSPinKLmkt8ZPpbAE3Cn/BwvxDX1Rlcnk4uW6i7o1dfbprr5
Uy+oMLmEsGsQy4SOKPulpUujipeIKKE0s7PEO9WOzGh5l9s7qCqdxlO1yVTlAaip
7o5jXFYb0TgFKM+nvu4+R1R8SlYWpRH9CUg8s/f1STDr1ReglP0WEFWSnxSiH0Od
jDtHI3EqmGehg+bZMRf5oxjc5PZL3heK7QGSuYQh0C5gcMq2ihQ9CHCGy8di5Pu2
dHvT7h+ZopdsJpC3JXH8qqGhYLA6aLd60yUHdwqsB5H+VN9GlMfYZo/aL+D1UVqN
kYrLxe1ZOpcp6+/p0i07cz5+g1gx7CaPa1WZ322UZuE11XyJ3VfFvC8liDzBw+wp
wTqkqT62nzdFAlgdtwmIgVQSXSNofWrThAVJxET4SqhFyIvEmjSJgXTXzvJDAsZc
YT/nwqARj3vmCgozwEpMcy49ikXoGJUFi1tl4agt2c9Jc5xYLp5ssn9AB5ngOe2E
qO0+Hn3uRUdkqu9sGd4ZyelWwoEiZ5/KShieGiNuLQxGiYKOESHTe8f+/iMxCTSt
HE/kU6jqxRoBQTwNFU+DsMv8yAOwGRybSy8BzWwXPKIYfHDLpuaOiztEHPjmIeWY
ky52Mx75Nw3uvALKFfj8UfeerO0c40PzoA/44dRa7Q03aDPap7lQKF9q+07i+Fmv
Dy8VInauFekFile8srXFXJ2+T4VjxaMeyhJi68gA13PxBTgVMt7f1ulseOdb0BMc
crDUOyuvwqhHXAVGKisjKF7HMvrSeWXgINMJZf1hG2t08VWSZSCzNNdhgf9c7bmi
mabPdNIj3KCmn22bXpjhbX1Dn1e/hPIsfzbd/v5VrLlo4htHKkv/INwAKSJaCvup
opiL/giSND5Jz99iX+yyxmdH6m+bh6WO+cTCTPevXN3TcLs8nX6XM9vFYVCpq58/
hpQKIF2Z2elGwG4QSvVs0xTtM/tzM/gl9P+0turXw3cqYz53+YASZwsvgUBDAm0S
H8GLavh7r8oPohTQJE7sV7S2FXoWl4lZI5vymIsQNpWObUgwQiVwxXtie1yjfmB1
V03srmYmMxtn0bfT3R04QS15RaMN8WfM2uqGqa+N6QvbFkZs1RC8umL267dwTyf5
iG3SavO2B1dxUh99N8rsK/ZZQd9+k25pg5fXmnS8FX4KtZZnWCnESoW04I4hRnHs
B5cCmMuupANELOgbXzigpWA9y0W3mdn22KKfPvwvqIdVKh3HV/bz6Kh4x7bJfIAY
g29EOsVLYLHdF5T9SmL+Xwa4n+Sq2Yz2OCx1vNZGyX3FNWIb/mQNBXq29MDXYgL+
AWrs/qzKMz9bcT62WzrGBUZ1XLQnnZiGJNfeJogUXIEUX80xt0QEJWTPfDFSZnfn
cJKWsINSakPwHSHWUih0kw3e9VVETXqKAZrW31FqPn06Ft8RdOAjSKM4F7S7bFiC
VzcTCTQM7xOAL4W/4t/LEpWxNKm+zA5REj+yLFh5/Vtpg/6wHeF4r9zquocsqvPZ
6iWBVygQQbFn4Srba4QKxWmTEZn9RuRh1UfF+aISY8kdE8qqHAjSVV5IoGxVHYFm
68bc02h/JqgTiBGCSAUw6R4Khu6B7jQi3wK1JWZmWNqNygaMdp/cuRUCDVMN1tD8
s1XAyoXr5tv7TUwzU87mTZREMqlWeJDIlQEpzxBKSGT/ys3+5pKyq7kFEcCE3+Cf
QYzHi6U1uliuohtjagFFgdzXrOfJTaU6N8DKFjWpW7z+9WEZpyvX0GVpgn9+MTqH
ihPt0FyHNMQAnZh1/dm1o9Z+gqWIyPv3sv1pPiNFSvowtYzFajBA7Oa9apIHg7/Y
kibMNgz52ECRZ+m7h9kC0p+DxfVHDvJWs0ALBvHv+QNCefyLAgVvSXDUNWqrBZLR
mkvtFwlRDkGOfAy/+zmLPfgYDew7Tzl7Dr1acEHb+rFr7mtzJSUEyWVQvJ475JXw
lndV/4INkt5VwcMR0SUsEJraKFSlEjiqHYyc3dbRT3cJ51riC6Xe0U/UjVBgKOZk
QgyXYEx1nTpWuoHo3BTvg4aqUiqf8GRg0d0wkiCapClX7xmnz4Kopv3OP0dqPAKS
JeviTQWtnpIJ1HKyvAaAryQWZiTOGmXdFFrRvbKsSyXqkQZcBgKjfTHS0ulqrrIK
p81+Y2K6LjJWXUmKVDE0Oylj5RhQq0bV5peDnIJAT1VWLkxS+/L6vD1CvMlAbRYb
rmimRU1ohkV4i9yjuZwMLaRiWu7jDOcZ7TO2jOPV3LTzNZKk5AgGeAxO0sGI8dHK
bW/Up7g3elWKVUjD9uDDV8nBr13fkKgMYPJ8HKN/0deUWrPtUHiwRnOhjsLSN3a5
H8DtNoUmzozvK4D6dpMnXEA5gl4NBhk5ssKdxE7S+sk9QzmwB/kmO6EDnDaUWW8P
5ylUHUNJRyThamz6y7r51tBeD/n/1O5OuPHoST3Cgc6oxPAniswVXPvr0BJt2/dG
a4mDptgrZDk9i/NW47eZIVG5HbQW8Sb5fqial/SgcLbrLQTOoZBW/sZxItmWCpyf
yZxW6fDtBJJHmK4mmixSxu+gGo8eaXDnuPkInTR3uJSEvlkdOJTeqVrbV9ytC6Eg
Y6nNAQeB68EZLV9ZRlDkrCzc/ukmsFXRQQknJfeMTzmyrBxt34pMejbfZVcMcZPB
jhtw1O8FKObau7A54IFL1InJzdZbPE4fgmjp3P4zr2auppgYFABZNTe2ZQZpEIxR
FNxsnAe6OxdYZLWUatdl7W5kFjOGT9b8xi84Qd3M6+WayEa5cqFz+lYBJ75+j8j4
qt0kCd7HBwgsfaYsG0bWTDzAPScW2mYT/UlRKtYDkkfS342cw7BdRXHzc6SpSzeg
ny3L1ADfvkqeovVKQPWowKBLLuYY930YZWpM07ZREaCt23QfLc3DUDFeKW5qoLoc
Are4HtjJxIlwbffdGoMGb0iP2/5xmsZjmHpsWPDG05G/w4zI2w4OxKIuVH3YU0Vw
pWGeFxcT9KeQ/IJgpoUMOwoeF6z/hxliiquAAgfd7GlCD0Z52kqgjVeKoVXhs7HF
/L4RarLacXo+7J5X7luvKEZDpYZSff81qa8Xj+iUd9IUpDbi8QGNYDq/9Vx/bnHb
UQLKzKBj+4BXqrZBWQwXJVwTyEuC5jR8e9zbLRAGsgfFX580McHLNVQkyG+vRSj+
otqYfvRK8mTsQrGkM8li2w65h0Ghh5Rd7EjnVGvUX3rRZhbNqcySA8eDZnwVFUYA
GmaElHlMsv+r7fiZpMLJFZJG71wqFieshtih6KA/XGEv79I+L+QbsDdmNg9yc66J
WqmCMfFVABFGI6qURUv/7XwyntmtGsKq4Ch5RmdOaX3zDERHK6F/KZlMu+D7MANR
SNSPhuR8lkAwo4/JNjQI8iWkHhvv+RpkBV6Ux9x/XYsHECSKjoUixiqP1beBm8nZ
XlbDhEHcg9lYemWTlCXIpd0gpBg+1mH5gJ/+UiJWVM3qEXmjAzYlqtzIxaraax1R
UlSG9RJanuOUbVGtCd8lPQFohKdk+4SjOTU5ogah3ZI+hIdLM4hMfvOmCkpPPc5A
EzWjdjvMNUtpgsFWN4gk3ucam2B16hA3U4HyfeEIIIuKLd7vCYRsndYmi+tQlEBa
sIBoAfbksaVe3HIkY8gdHZHI1bb00nRSidqlq7BFgEO0AeKRVrFZKdQhpOWEqLme
H7gSruuENK2YX3P1iut2/IQuaPzFyrDRwm6zLtrwUhhf4LK3a0s8gcHu/R7m2lef
3y1Sr4CGrA0HuRLzaZyfsIhrFgC2choUkWhRWX/4/3oe0n4XLt/2vAnWlYntphuc
RTY2T1KYV2wRGPB0QwYg8gWgEviGwmB5OUfyWlrldDQo3K5t9A/+UCkwG25Ss+H9
MfPfdrqbZg62A+xs8lsiZq09j9FHz/pJUZJBf4CYEPXYLy9lyW3c7VhOreDPP18d
13lL+MjmVfDu/W3BrMwBvaNi3rDL+W3X9XmiR8ATka6kHeDuZcN/Q5s0SrpTMwGY
lIuA9bg6G6BSAe4kdTTyFST2zZPTT2AwNCSksBXt8XiNXtdetv1h8+J/kUZ2CTq1
HggzweE73QbN9dKfKByCd0S+xdZFGuYL54qI0XgZb/LXQlYt/fhL5Pjyhy1MjgrG
uiOdpYdDfhUiBGj7iT3D5KJ7wARUgus99tNXNykaF5VbFzt6FCvfijIVaxKKSpJ6
ec62YqT/3HIqAYmdgQP6QcGNrPgtvYkdF0CEaG3p+z1bpJhbgGRKrqZG6m6+kLk8
bZvOfcvUHt4unQJDdZxmCzgyw0zgjRYLRwvSRMKnfGPwEbMbRdGrWuC7H9cAlV7S
+GKjQ0x8pHcHkVuXjH8dkJWh+WDe1sH97736tPOv00iiIDJkTBTrEOx3l4sN+q12
s2qRLEsAFBJ4TBJyrYyGqZXcH+aCW/BplSoQe94SQ8S2Tra67fJ77ydL7rl0qbsT
+Py5wdn1HhFBGrHrOFQsNjrLk2zzWAu0GaK/RotQdZGkqIXlaadytWAB+HpjcmOv
6j4zlYpcYeCUYqgRQhfefu7r+PFBXzcwAxaH9XR/GjZdMQifwHzDQzFu5fBeauqR
JQMe/xzoLyQrrEi+C7CN7GaOW3/AJR6/krQVsYECbAmWJDI8uoHhU3AKTzN3Z0Z/
rX1YpLMeduuY8s2iaqwvqK1L4eyq8jsMwjHXaC3fFeNJ8Ta8HfselTS1TW2Npfab
Qdw3cc1T24yYbQH+3nnb6R+fChuj95zMJRWSKiS6799QzWHGSu4YfEdQqB6yHAm1
CvOHDHHCkGZuK2XAHo27XymgN6BXBffV8/EF00+Wt+cjFleSA/cLid6eK7vHE84+
QCig3xambBNJvCvHBnQ6+M7zWvAsuTeu0O7QGNWs5sR83MJ5p/qrvqt5hOexfEdL
7OLUivDwvtdgkz+2eKsdSXYqXwGtvDATss4StHJcsdZCgwNvwMqmw4WY4scudsyC
bMAaq1RTkVXBCwVaEr9rKUln0snvaY0rZFqf3611ARJE+KRl/tMuSPqLUPJVIkcp
4RDp9FFx/gFvS3iayssLuO6rQrb53AmIYKszd8lR8hfFVVS6NxLnyhCZfaKwTibj
2ZzIlrEclnBI2DVYbn/NVKhyMnv2sLeAISXEdKQ7oqxuMk/juiujHuMR/cfpz1ag
Y98ouDVCIfgfXFZ5nI2noRjzqMLHbfXqoC4n9ekhcshNKqlXbJtMApGAMqfW+EYG
ZBG5GyZBmIcSLBOnj63LijbaaHw5Q4SQeIGJSrrcvi/3G9PYQWuUS2l4E7UpimR0
uW68LwYkE6jKSgZOHLlqPASenjOLdBaDPlhRkyxGwlLdubUfqTp8VawjNkbiRMRt
31zqNFJ/ZUHBgpWi7I4otXqDs0T/mo/tGJeJjuwROxt9sBwJoQmO5oU+zILteZIs
DJdHDVVAEQALw50t/hnDLagA/4V8Gor6WdRYPfX9f4vrHel+wK+gKP56VqpZNaVS
eaHTpCxKIRKhdMt3Ok2pF6+unSxOfJqBcO4VczcrAr/6J3zuj3f9VfSkjEfb/DEL
KXfLxm2LKE1tK5SVS4Qk/wg7OHc0Ys6uH2qrmU51RHvSIWv0PQ28OgUqJqEykloG
AYaJDySDb2SsvHGDIwRo5Oe96evavgdsGhjAB/MDrELRnc6Qwuyv9g0a8TMWtrap
hH2mZK2yinTpRodfejz22TqggHPljR1FEIvG5pGmSoe6wbZ2KwZE95F9aLfApWil
SLBgKvz6G8Q6Dr0ihdD1rDGkK+fDmiLWg0aOJRsOVHYzooJQpDziLXNku3lYzNY2
LazRbDJBNjGuguhCpSHCPSRH2mF27OuMav+PIFXNi60rtrbSP4e9omHowNuuQe36
7d7kvcBv9CSpQRRKzDa5GiGxkAsfn3vZw8m3z8WoD6klGvAX4/idUpY60GXxIWjY
ZE5vPQtCB9WFX1o61ZyafEGwFOVpC8AeSi9TqOShZNJwZEyWKdyyBnTO1IpkA/6O
zmZlepidVC9HbDcSyFSmjDNTJyf+AdNHxQgKt0RncPe7BLEV6wc1dBg0GsSln0ut
PaExUS2dKDdt6l60mIWWoFP64Pr2TsqRl7BUoWSYSdGGAQXHJu1qcb9AcY63hjfc
3MHCgRLN6voIm8RX3aL7rtXYcUxEbN2pEZgNuoznCgh62PFjKvt714rm6E3bshDg
VvC7HXaH0xAkxcy7bnSu7rWqQnkeieT3lK6brGDujDoo9v/eIoDP7ps2jWOvTw69
SzMhwJSVnKPIP+cSZEjyeVb7zVi4WhNPwyJHR+R7SFYJJBSWPW7FDEEnugxho4r2
cTHpB6RE8Xkj1zX81g3IYMQfr2qcLjFRs/yaeemThWy25j6HLCNvg3pgHRCm9E4+
1D8NIXs62xgOT2NyTLMlbKShW+jiH915JOlLxd6KTo55t3aPlY/XEzuzQDeVr2/+
cz6cZqKnrJG55kHIeiK3wSwanXCi4hHulKo2ermjXfzste1hZtW4HZmHPJ/EmjMe
8+HWGHSBTlnyPjM6ogtHtB6jAsBQCYDW+Myc2d0UPNvS/1r3js708i7/mPwCNexM
s8TqokO8fgd7zEoQPgWi+7zGFwMe4sjUO0gGwiiDeCQ7b0DWhwIGLYJKKAl21rCd
UJPrWOc/fni0OBaUZh+gCSu2629GLNcKR/qNGmNY9zKv04Qy6z0bu6FmZpRa0scN
8w/nENcaJ7DnE+/9wRptgw8RwoWsJ3ODT3FCVYcK2Mdpe2h+VPgBv9PczbUuCj7p
mASoyZHaagHlOHxzaCdchmNj0uD0XZfP46pTRgePjx4XjZ0Zls+sps+zAXO6Ac26
+N9NsHZIPveIlFr/BltraRTQXZzGl7etLzhDMTKDVgPDCNKKzuLr6ynDkRvgXQfa
3B9DvA1HUb1IsPd+xxD0HZF+hi08M5ZFbvzSBGRckUF3A0dU8UQaFZVywonADDFn
/WBb0jemS4sjAjWMy/8/7WpV2NfKwzD22lEPTGyYJYyGVKESN2fHG1RZ/CfoNs6G
go6TD5jypL6HnHTJ/DCpg0MpftgBFSvNYrp/Tceretpl+fGxP0Co46Ip7SlzMfqZ
bQzySDpLVtq4WPalbKQ3S2ACfTV2Cspebx6Sm5aWTF9Ke/cGa+v0MK3Nn9NVpIuN
AH8AklxqwMh2eubrfxtYBly0R4szCdBfW3zsDPyITdiq0069gdC3PCiLgNl2CZQr
EB9g15d7iEGZRxl9gECmPA55UUcJFvZFMSyfWocndKyJm4Y83szko/m0BSRxn2Yy
GpxM7OxhSsP2ngHeiiloL3NXjR3y70Z6jSUANGuJ+OxfDubUrCM2cHY8Xf52CDER
fg6dpxP4tZ80cR5jpSBsTXKhHiuQ264GSVu/1rWtPXrXdiQWbOypf0QmNe4CRZ+3
wIxW/ELDq7faj83zEjzkCvogU2acs18NNqBwnvIyrdMv4TI1Lw7qdrY73zaZZt2n
MwNo45M1ehCJ47lZ19WnMhklgoahOGgp+yi/+Fcb2xegf7m4KfmLvEDu26Igz1nb
MvzWro1dWN/hZ6jxXF18nK1jd3mk41aD+xjWfcX4FHPLghiQXB4Gv1VfmNCdKhxI
3diSwhrH6B4f1DZwrLswHveXewqsepVhzLbMUdtYeAyGYnAntPcSNtFHsa9phdNw
fOg4Wm3raOI+DPCudJbEvrOtT4r0JSXMKYq5ochASZFG3u5P+g/upzql+Ar3M21t
xWwsXuYgmpjK2xi08b5awK2qBLU2539FvORbxrnSnLOh7cggae/i5Tw9NKP1GBnh
Efe7mNt/PLKIo3R+2fCUEHq8moMTegrhVbp21F6dsTV5SmmBaEM13iVTGKb78Soq
Pj1g3G/J15dAF0psU+bb08q7isdsqyJUfjC8b3Vh3CTz/Xe8LrvBTjMvky1ZW0g2
xjJCfKDrl2HhsfNZprwOJOhAqadVzn7w7x5ol/Xc4m8wuq0hecfRt4mqZp92FXQk
YoZTEI4vuh+tSxmu+MtgmC6v2+qEgiFcMwBmUePIDQXeA9NqiQ9P9XQdOHXQbg6g
OknUIqbAZ+hjeYMs1xalaxG3u10Zu/AsE536SCq0m9Uvj4uF9NPNUN8cd3LP6V2P
7sgyK9GGfcvj4SUdoZfUo7aH9rg/R8nRXuslDCzSV5USBGOLmLoE7/EserHE2yCj
Vc7yBmesDyEZLlbNhThWcRYlzjEX7bDcDICo03S592I0DcJTDmW1KwnZvvtKdtB7
Xrz+kfgrJ8oY3I3F0Q7KJx0YnYtKRf3CTy8/Y605V75z+VbVYAR1E6sIDajwQ2/x
fWH+pVzkr2+BT6Ju1sIHkxLUqvYywv1C5ow85QXhpk2F+GzLOZV/vq0Bdr0k9Pdy
92brgEZpF+i0pFR5ZC/zYEfxckZEaeDejhNnPAYajA+F12C6bSwP7kABhoU/0MuG
rvNx36N+erU9vzMKqzIiImSyHFoUmjIFuEhktZ3QGKmd/XRDjhJ3wHJTzEMlBPst
B00h9s4B9mrejEYrwjHqch6bOw+1LGRDHok5Of2KMA7HBIjVsSKKVgYGASSeSHg4
MfH7/IHwT2cX9g+P1UjJ875vcDMFBvygHu9MqqrNOxGaPRL0RN60JZ5ShknmKTNd
0ZU0/6ToBV8J290eV3ri7oQ61roA+giC6jP6aNaVRfOdrbmb6nLAnTdYf9Llnq0p
tTEsHtpDzKhktF2HrGzgnCmjngzYzHddRPzHPUDZI+FsLpkx48p9UgyfIwRoBZHV
CaNm+t+MOtx9RsrO/GwcT5fWYXMMkVqV6FzPRE3yX3nnaPHPiZeZJhqWVwiYenTj
VjUPyDydAcIWF/ZGl1pEA5NT2iJOnO0BmGPyjIujxK79CL6EJ4Gt7KoOCmT4Z+ed
b5S+uv5jdyyn5uBu1creEuOcZ5+NvTRH9aF+Z8wMbPBs0Ine2avwpNub2I+3PPa6
0T7tzfJY0qlkq6Z0WpLRH97/5jXk8sjtNN13WWCd0t2ssv+XmkRFMXLwEicN89rG
slAZ7+SwXINvngk29YybweVCIJkk31g6duWIs17R1e3ssGOfejdQe2Z58ZIWkU35
FvAiS2pH+bdgktG+vCkB0NCN4F3CINs37v+1KybTCqntJua7rO28ZHkZrQ/0yn3y
HU87TQUURSl5PpJVb6iZEfiRPBR1Gwq0oa77MqFPIr26ncuQjq1e9rdabmAO+REx
cUAM9F6XBtwmMgHxQ+UyH0Bpf3ylWMwN/V9tQL0Ov+u3lojWYpjHjbVNs009tjHb
GUayJPIdpe1eLjvIp9ZAsbSAwIKY5IJ0cH4mn4N9IPfOT3ot3cIayaYpl1aC6fuY
j6WbXT0WQrPg7CoNtPqbNx0NwBUwQ/z2etBVlLtAoHA6fidPrtKgPX7hoTNDv0oR
8NQfTcJHV7oCq0E8xHsb80uQOZ19c5dMTX2JEEOzivDkR8AWJVTqHgWgih1D2D2W
1LODJTXgxPdYXZn5BFt0ee1dEzkgc1gn/wdCJTXjbK8Vu6kbrNSXhdAZ1tVYKRac
UlstYVrTvRhMpP9dtA/adD0f/X3oIEmAJsSoXTEzfB9JoNP78QNSF9ig4lq1d78W
utq6mUgZFd3EX9lvt/2wO6NTGMkL0dfkTyqShzhgc7szLA+7N4guG2fMKVlswmMa
ECch0Hm/p2j6VYipd2bKJUKJxQx6kObcSmNO9fcTR4fzvTBsdp5VPpQ+V2W40Xab
isPNy85cWQPY/vNXat9Cobddn8lzPOtXRHoXpo30N8/CsV4IaAmKM0qc86jo2zYF
hsHYIpaNOWOkR77SJnbrzTbmVYTQu2L53hn8igkRUAko0AifXoAP4beEo+0A+UMp
iJIy7ahlu8NM4lHjk7hvK/+cnWVQRgbiTfVHqDxUEkauXtbYwuVjwoyz6lh6mPr4
HEvapRHttcz/xgVr4jXPLuTAraWxAGJSd3PexSsMHl26fEc1b1s59dL4dDkHy8E+
QGpH11Oc6lVaFN8C5oE0S16zEAhPh7P/uiRSbDO1MDkTk9C80OzcnBS/bkXztp0t
gjFbtpA994E5mgGyeBHxAeOrcRpB+qlCRBsJy3lsVbr/8b/S59Sz8/1OBFoYAnMj
XF1f1uQccjKcdlXkxwtsCvRVaC4dB3R8GU/G6POrQQUAI47SuGPWlniKyDNtjjp6
TiFhtOI7Aw40/eA/QUMGVxtt0r3HsRnD01rQAD7FSf5zw+PdQcEFKEcov+ryMWAR
7ta0XQa0FLaKr8GV2rSYneP3TzaO9nhudCf+gQ5bxvEUHgBgPwXEi7/ev59Wpjx/
0Sr9vFH0wFhsHc8dDNJxa46eWwJufWdfsbXaQKJloJMPOPDOHnJ0SWqM52Rpn2bq
Mx1XZYz60D5s73inIGHclz3IEMPMaYGXqZ3G4Sfvhsn+D5yuQ6I0cBpGtM3YlyjG
lmIC8dnG7ylTwgDckEkMQVNkooXQ19E1XOy4WZZlPNmbI3X8Ssdf1lt+7y+K/hOs
C5awB0lU4s400T/Rq7aRa6oD/b00EqO9mn6Gm6Y9ymbq8JYCPnwiONGApG23+SUs
Us7p/rOtoKN7IBQYQNZW/upeaNZLfLJ7D0xra01vATtyKd7BgwDylFpl7dOJ2+QU
EJO64yumb7FfvnFbIYP0DuvxN+yIvxnN0J3fGlhW/CcGY20DU0+8pKPO/BIoHg20
bszZYln278zf0o6DvlmMEX8yg1nfUi28j5feV0cYECrbkC1BQAixzmRN7Og7gfeB
7PYdNata+m83yT9xxPizWGtxuL/eQGV7hCX8oN260NiOHCr61shEqg0MO9aXIS+D
TrAN1BCyG9oTnJAFcOzr6ST/GcMezyCUSdagxFipNGzWUf5WEUI2+vR2xKllfxvc
7hh06F/QSvHZnknWzLhVScN80xYrTHS+CsJesI8+NVfgXtD7bI3yqrFaLQuKv3rA
bI2vu6mSSv8BfNKoCZreM3eo+CYtttnBYaPJ0Y5meA6nzT3P/kVepaBPzwjTLts3
RswlPrGNkSBc0VerLS3+FpeCPk34TYajPAUxJtDzbYq8GMSbun339CPqyyr3IuBV
HjJsja+NSr7XrEPRQ34Aky1Q5qS4xtd1Jcsy6YPzBSd0kldJMJ2PGVtwrNWO4uZe
MqfcHJg1LYntcPBYqqVBJWIh//LM42XrK1SrtKFn8ZXWbPDSh6AEopOayzPEIwSf
32fNED3kCCDYpX938avfLpcZBmR8JINa5/DnWsxXZyQgKMtCcmdziQYi3nJB4aeq
uIDFBhnWgju7hrHFdD840Dxl3p2Mn3ebfkS2h9GYKKAy8YUBK6wGGFx/a63G5yby
rsCDjWsFQiJAjdBiO8hAJR2zmqX9hIuvaxgPqyoa8wZWWfVKh0EppEG5lIvday54
rT11iHKVITylXpf6eSEclZmqM/BVnYM20gcXJlGVMuuzmV/T0FFywKEE3F8t+AJH
4QEST4Ss0oQIzWTCNi0Q62TbFYXxWDxJL3OcW34A9Hwx35pnPe+yeiaaUTrG2t3y
fjPDBjWX/B5QHN78Dn2cDHUdgVLhjji2MMCDt3RREUja+Mx1ve5Ju6J3UdWCdD8m
wCHTHx3tyDMEccLE6UEUH/QPVVAipWQwAlcf5HYSvP6fZKcKUdqDH3pgNHU5mcx9
K74njTjeh7YoZEFtKys2RrhcBuBIhP+YH1ZMjVNEpa61VviDLEtFQiXrevCrBAvI
tWqoTd+XfKkRQaxbP89lQ9BvbY7qPmU0CMYwoX7meWLdAdI5Kqwcbz6t2VxLNbUH
lAOqyaorDFn33zpJJsjVAUl10t2EmRaHqdGxEQWYEdX9P1atlEVL2VpA96USbHGj
tjmUFbwVmiTMD2G5JaRaB5eX05GTVaf8DjKkghSAyvcrzHp22mKS27a3snsTDTth
u77P43L/EjvB+ucc2la6mgjngx0ow28PFcFc5WhZ2EZZFSf8JbHZ1ES4hu3HP/Mq
4FLbpjfGz5I7IsO7nY4g2xsc6dR5g3aDELUaprbdMvXvymnQdReeSdpkLelYQliU
TNuIaleQ/4ZBZePuAt3rMq6fOWpFZgWIYA59fCGZ5naTDdEsU+ZyFh2tI2mgCHDm
AyjACLq+zSEXI6/tKAScDz4lDPHH4dtUeWXy5XP96Ok/DIpHcFg78KMj8x0qZMRa
gBBSAty0MWYDbOIaUc8sBEl3s+DfMJ+iRVsgo+UKlMsXQgWaGlZhO+uj3GZfMMkm
xsfNWrYJ97Q7MK4r1qCRn7Fylx9edC3C7PWLJyTP971EpB9qMzdOdD7V4KVLZA86
5ihOi1+cBf/7Uu8Tg65BrcjTAx9yhYwJtoAe9oXpRe8iUkYmNH8T+rgspfxbYoj0
uZYiS6Ztk/GciK31bBLsXHy0VirlJ9yE0QyoD4Yr0Mkxe7amdZlKTS34CNuyIfR8
h15JYHmgjZSKxHD/yXf0+Y+3Y1x8u5LftV4xNurSj9kucpF7TUZRkgY/c+56tSae
BeLSTmADSiKtIS94MDgx5Rmnn8cFbcWFtfpvSXFHViA7E0rFb/JBI/J5Zi6BbNFF
haYCDS3XEZ+X5Lh97LQoLD6aMMSfo1cY80rlL44d/Az2uYZUuf4dfbuLpAJ2Ep8B
570qF3XxkKdTy9U/HW8JwPibDn5ynKxwxrX96uk2Lz1bX+7r1MWFx9QWw1QVM9l3
pMCqa4aNB3XCkMWZh+bNG1zMBEPY08ng5csv7UU4lrBEqS47TANbNQvlau7zI1zM
tCmdzcK1adGht7FOuOQh+ur+4OCq390km3XIEuCELlK0+KAMvA4GiByhBZucM9C/
zC7K2dMB7cKVCwaGJkiSL4HIpjqjeQNfNgGXvFd4HXrlGSZtaJslvIyAYQNP/y59
UScs5mYmw/kgfuuQGvYe36+PL3/xacmP+qF7AignbO0fud8oJJ1j+t6soCIhSWDM
NNwt4kfTppoaPAQR9LnU8//jUaBFt/jeDOooU3/Cf06/AeplcfEoibofQt3NJvCR
ClgeDhU45YFrVUTUPYJJbYg630YMU5QjmMtzNGsYxBW5Ctu78AOCvE6tp/xPLvEb
G4fYcc0L47PCxhaw3nXY5qPRA0b/I9J7JHdvgwQIivzM6AQkjm6PewkMPyvRJg0s
4i8ZFqHbQjIMlPHiM8AyDGsulOnphFcCIFIewGyhF2X/uAjw2s9kdHjfH0Yfj81R
R+rJhDBuLatrkzMbJT0gDUOcvaRN2K8OhEYflZndk1ekOdilTe6L7JCT7c6exKf8
BMXynyrtKt2qh9cdhrY6Vd7wKoHDjNwE9fo5913XcCGgQDVJCrlNIPX80np0zw8x
EnZ5RF8NezWO400zfZSUpmgSncq/uI4uetDwovZdkRc1S1UqZroeE61bVWYboGfV
+588TWQX/jH0wYzA5MeKjfAg3QnkOBF+r9ICVWyP9sU5N8KeNInng8pIa+fiwOiU
0l9jJ6W5n3+bH8PUPdIhp2+0DWwJHVmgjKQyY3qR8JGilbAJPQFS7W8g1Hb5ef9k
9IMC3Fvbk9AZ2Lvo6j6zbD8bhaJrPb8SUUqtICrgEtw6JqjemYvQ0RQZej2cmZWi
5QkKpNV5xfMAPsFOJiNVWFwDfEYKCzNl3vREfggqRFSoKKq/haQibE30FI/5yEKH
32m+mfIucEzWfqiSWgoM7IDjmKZNNX+xOCk5x6jPtQBFWzppkI94GbzBVKPfEZnS
uW6ja6MUpel+1sw+9gtGCdEAwFPHNYhGbxY4uMuVhOTLWSoWS2nY4UUb+qLG06wD
t7vIC/lnuTezRD0aF1T4YDptKj5nWcgG0evgp3OHl+c2zjUSYM73SMMJOitkvnsZ
4jB/5jndgnNzOpXpVuPPvhlgWmBYoivfHI3T6oTgBD0/fgeolWIM7r8QMTwXBq90
5VzjSnv0eDeOeAqJeUPkXjDlFxJrErJ1qBsqArHJKrMM3KTeyaWCLY7Z5Lu90q45
eDl8FIKBEI4+q+cstVarLx1uv69Y7GZIXbeX14RWKY0/DvV9Jy2y2seK2ut2ITUh
PskeNjshjrad8vUr7NadJLm+7z1a7U6M4/LbagyPEZ3pzeTfW9V1yTyxGEDqBY0F
0eoESrPm7qQLRFxX3XxBFjIgL5KKuKrABRKtWjpUGvTRWbGCaeKI0S7OYFx/1QL9
MqVnquBdP0vNi9zNCmNakFaNq9iiJ1FDFwoEKDKLin6nRk35mj3bXjgCUBckBRUv
F0wLFRz+LBIL+e9pCaFd6DbWCp+V8Mtc1uCwsIwQ2QPGZg/NV+5+qdTkTqbJvuW4
UxlmQJRe50xKAafkWWsKL1XDBcrjmFvZAzAUFBphAR5Y/vvgLV4M3KFXcjhXgh98
+/2qGbJmcPz3KGerG59RFTRu5XeQmKYH3OfYI3V+1va/dmA515AY108yDX8Wrviz
/e9DOL7XmV7B5cR19wg3NQ0PElmo31JRXgkg3is26VMRwr1gcgX7vJKDB+505CCQ
webvcZv6qBJP8KCs/7iLSYybcNVupAsk+ghddOk4IUHXvF0yo9vzwT6WnVF5/Se7
SZpE9dFrj1WER3XxJ1bqxp3BzJIt6l3GyjIRK581Y6AYdNy8esGQhey6blKOgmBL
5qDPmDAFqzcczTqjap1Z6cf83OcHCxUk+J8XpwjKaSgbuCdglfHjdEPpviUCY4iT
XCzxiAQr1YaQv6UMKkucRK+LvAsj/ISdIb7TZYzuYuRU+rntKkUtVqFmzghfgAAN
rjty8ZCmC78V6G6zGK9W+aZN2CcP+afwH46YD/lXcx/8L5bJOVGRIPSNMUFRERKL
c5fOzio/Xi3yNh91t6oFkc0i/uTvOK6xrh76Jym3PDYG2tBYDg0NX04OGZOeJhj3
t0JoEy7UNlyeWhvXM2m9326ZyAaTkexqusdg7KdTLr9AyXyKAL1ySBztR7vIO+Mc
CDLSjPxJBg8iN0vOZp6+eot6XiGPSc+Z9Jn7mDExZ1U9zrozcIOYT5V9/QvOQbr7
FcITKMQpSZYTuAEHSFXuDW345SZY1sg1BW3nVJpsw8zP9S66SmSs4R7hfV6g4hqc
RHek/24ozChjed8oBKdmA1ehM1BV1KYgXwpo0k5iN9c+N/zY1mGFa8pDgwZPpj3R
O8Yh4uBQpa9/9HHT8ZuKHb/GBJ9jM6lU1LvFS6ylyNGtTpvWvzs+bc9UVA/+AUq+
N4tcG4B+gPHaIyYCW8Nzr25o4q0r/bPTW8eEfAaR1x/sUVAGw/0nwS0pPiTH3GxK
D+aoi8MgfKGY5kmn9clOmu3cSrsBDTUGD0oZFlAInG9KPSJeXfdpKpvZPrORVrtH
P11MRSI/i5ZWZyxNELezSz0UljRULsvWO5ijNy4QT22q3g2EXPaJIU0fzas4Y7Hj
dj/hhAQjbHKHhbzHH5ecPohUbMYtAICONE4tyCz9e2VdflcLkzEs5XI7jQuU12a5
Wv67m05g0EZg7X8gHq4Jl7eHRp5F4IQLZQrBTTt4irbeW0J9YAlhRAwxXTdNqcQB
zSBtDZiUkCcyKhpBoiDj8y7mue2V4nxkCW6MeydZ8H8Ey3dI7R/NN+LtJFcUsSrH
deMTY8xt6kgPuKgeBOTai0NBJBJp9NsJ+gLLrD2k/eDMaKLmsGpuyRwN4j5wecUg
JOdjxhJWzc4mYppykvP3HQPWtuMZXQe9kXK6VKFlbQVr+T0+R9Q0FYAzP19lPdQV
fZCoixPqyPTmYysu5JVFMHM+cN9QKpb5kgpf3JWpODc1Wt9zvBZOONmwMtG+x8Fr
GUX+DsvdDuTLxuxmjk40f5cwkOAPJvaxaE83w/f6Ktj1fNjzHXRmYxwOLEGeIjdJ
+PpfLZ6LMFweiFYimMHUMpsJ0zhaioNMm9VJie4LWKt4QepzXib6oyu40qrL2oKR
TTcqRBlkxNN2RPCaA4u+1I8Sg0TR6cNUd4v/y34S0pUboP0EVkhfm98x5cqsZGl4
ZDSQE9wZk+T38gipAU79COVplrjm4xzaf/lspjSJ06QJaBnknUj+tIJLvSlpDb+9
J7vn6nMHRaVn81Em1FGRkF7uYE+zQIRdENqGmPNXEHKtx90VNrHqNK05a8vMvpm7
MhT1dJFdLkw+/1FfpLgochEPCjr0CyYEFukuComG3ItmiPVLmO8srro3O6ahxQ9H
qJpBgexZv58DL2Xk8/lyz3fXImdrlpz29KIAg6JSv7SqV6ertgbdBdt4AI4Cbmy2
qOa/tTLfh+gPXVRYxmDGmMj/ayRipf1CwKPVa52DfWnf4TTk2MUSvzH2UHN0K50B
1WWh1lhyzUzI8TJhQDoUcOdqAtTDWOk3vHiSS3BAndSC+3YKz7AO5sMcXfA5g+/u
y6z1L9izX+uZBpZS964iO0ddJFj+Y1Zl8r3JlQayYdlx8Mzn6RWo5aLS15wlx/L3
rrm6XfUe1AFW0/0xT3eL8pd/AizZ0LquL9xxFelc5Mss8aaOXFggn3IXFd3tlhu9
5aTwAUFhqaAFGSlcOKs0c7nLNNbiINAJ7Qr5RCdUot3orDuSmX97wBA2Dontq1Gx
+eJlsBEINI92DMjPifA1G2UDMVU9sMwcXe8XimlVHsr0VgROzJiPihMHqfGIqE5B
WQZSkbYEnibrFP5ML7LJi6wSspUEDb8CHi8Wv/iJTs4dILzevtZkSGmSPWAzkHq/
BLUdwdDKwyDvAs8VL2t5TOE78y2JOL87G3+Rx2QL1EgQWOuM3/viMuvjwJFDkUzu
8UQb4HO7tGzetOVxp/J2jIQGsmm/XtP7LNW3uazVrI2f+mUsDCV1iR7thzcZFKwv
q3ysDlRU4yD52Claz3d1WZi0hTdqlFQeoDhxEhgNzpVNHOS5+TFIW9tnWnEzTaS+
q2JbOV7N5Ro/ZliHS+WSLLEOSS2RXF9lBALR5gy/2DPHwo7lcwPoZsC+aMk/KprG
/AifSEpyEOpnwQH3A6LlmGuk2eWdOqkcyLaYOeO2b5JSdbyp8eVTtkNwopYEHiXW
eVWpY5hxHaVMQYm4GYFslbltnAim3NmWr811Yz/4rKbZUja5awlYsxNu6ecw3Ky3
4GWU8HtAj/bBN8Fh7Ge8Abq5OQ9Tq+jKnhW/qcLyxdXPSyRMqnRJQpdqjOUQJeRI
ImkyOd8+Og5G/Dv2aOwJ37tk2OrxUPmTAkn4pMvb3w1FAG/R78JOmPimo/N32BG8
49WDyt/Xt00EJ6MHbwfSBE1Jy8gG+Hc3zuz2i8aEpwHzsDwet0e9XUJgLTMFuJSl
f3HthH5b15Dtu1D14rgkd6WYUUHZzBnIAV2sO8a/FUUmMF5gEAfUrt4z1z1G39kB
WTqAfJJDlz3o+BjmoK2yCm2eGtdZ0aTSyU8xGv6CN5s2uwhO8c0uqVlT+riBxviV
flEN0z0E0GPHt0xxrbsU9rb7MouiWlz2hcujZdwkXiE63vEq/CqZnxxU27eqGwdz
EaywGpp0CU/+3b/vwr5jDzLm+OoYTPBviZajHuNEisZ9O+nYFKUqEzt44jbJodch
yBysgrY/hJnGOhBBDRGwNK1DNySXA/hoP03EsIqOGOQMA3syu19e4ylnT4dmL4KE
HT3D5xsqL7nx80F1ZVE5hCHTVM3JbQzDcuWvFQUfmasQKLqZYPXDfBtU5H85zRUi
We9vd3wSUM8qUptBYH6NcSG2NU5+bBXBpWaoTgoEMHTGovt73z19hnN/Ll/8KC57
DsueYh+Jn6Npg2uOmNPJY8I8I67/CvCgd4P5B0KTqzw9pB84iIJxdj8zGRUQCKfs
yTekmAkma6FU+hQbyKjWSLej4Z44BPaOIi/hESySqt7DdfNuvYwCUi4RRNjIMXMi
tyPr9zOxCi9bawVD5nqqebkwf89zR0EOy0IO2hd/GChgN/RfY85ByacyLyNHSFhM
k/Boq6bwYwOg4eqOHCxpLAzJFi4XprB7XQxKLyDLYRpeoxWen+3bZLkQZpwMMu7z
quCtB9x2qpPz/Ww0GG9rwl5T1K41ujG8jTKnjgOLUSEm8JazM25JeeRzeI8W1y+a
R4YyId5dZvxunZ/dG7FfdaRTQ/paQkflii5Ep9qgbmhZ+qdGAEE5Rb5qQ9Gmsnz6
GqXcJbpwPGzkltw0H/pc5vbiERl1uUkA76Fhr3x7yDXox2k6brYjBPW5vFPa/RB6
UVUzjkQbHZXcMJJxa7tC8VBmXclrcGcr3YiS7w2+O5p+xuiD3uyTuxLGkC/L2ly4
x1DeLeMSjyFRiMYhUC78RPWaSpxsHdnicYksjsxMzKWBNDRTOEHIR+ak2hpJYWLV
H+RboS7cLPMtiHziIqXltJ4I876TnPZ+6pPjfUNrMlgGH3NV15mkwyfFTA9amxdP
xxV+dqO28VDLnbacbN6OIbT4v+TeTfsQkvkMmK3YolucfdaBX6zB1I/HCfJd9NuN
lkBVFtL33KKJ7CxrgoeTQoL1PHy1Rc83EN+D/hiCU/iavOlGgGnox3LgXW0tjbIO
vHygCLDUi7Xf3rxPudLRSPS1o0JUclWb8VfH02AnIvSroWMeiHay6M4wEynUFGze
6N8nyvUkVFXVYPMEXO4zQqIL8FiJnykU+cUyS19XlFsliuJT2iNz16B8dPyUZvSt
MnMhNyuptplgzVec0QYcZjzYpmnmPrpIN8PH5sLTDge49HGZ8hlbixkHYTmv38bO
W991maJ33vRubfMQUGFqzQZdpe803rbiOpjQsu8WlgKl3WqLvMtDZFKtOVee/5Py
NGothsAWfWIScKc4aeVXyRl5vX0ZK7/UA+s9y4vdUAxrmQlQyKebl2J2ETUh7kGs
FEs0OFsNBqfMpQ7EFh6M4N0aSAuauf8w49/1HqtyZPMDCfGE4iYnEzrMIx10qZh8
uAswq7NMXzV3Hqu+47wOR2+IWwLGZayoYDrfOul3M+T6P9g93E9ufEeFqg07JGGB
aNJz1A9uiyD8SeJ2MI9VgIy8VOyQkh3nhREhPKzNbAwQ8hDAJdL4QOcWJJ9q+I6a
0ZuO+0fAslHKSmZzI1XYGfJrkH9BosuB3EXHIcm4p3EAao41uiCuiMu5S5k9AJAD
+szvV1483LAuY02kG2aa23iul4DZaDWF3m9eh2+DIlU0PMHs7SdQc0vJq110EwAw
VUtH4lkbSPmWSb3SlB5nK/O0YF0ntbylHsWg2L0bn27n37toraY8G2nUejNfsTEK
USygzLWxQ2uDP8C1A5CDken1MK5Vfj8ZLLAVrf7cHCSP+RrJ/NOgXiR0jC7iEmpf
ebMwmz/OliJY5ebYIfV8Y82/vb80cR50h/mcg3chFeDg2+kqcFev7/5dxZsc/sua
VX2gF0hnWNnNgGgE9VbWVii9l4twB9dI5RYhyjFl5QgUDR4CfvXxSsj1b+MV34Hd
smUWCe3IpVMHtbTVFfkEGGPtsJm8CwwLLLEOZiNjL7r0StvXavWP6t8ovl1chXr9
7Pxdu4LuQZwvnSzTTOV99gd5nkoZLR/BY/eYoild7OgHJYvHzMB+DXBM/DVM2Zf1
gWUDnfGGndT9xxmEqlIkb3HYGuXAOmDyauCs/e8BEIcJKQ4zOWH49f3JfhHyFAsh
fS0DrwSM8f1ITXuHqpKOcpBphmPF0VikoQKD92PFQ3Fi70LkQBc4DkriZhVVpHWi
8rnJUwZlMYlj2DgSY5q6bqhgzrA1g65A6iyFL2B6pO79RsYTchcnEr/LWOIq6kTo
zcYYWj+bBbyOhCs1w51zdIHk8FQAGBK8DaMeu0lTCmPGl6FnusbAY1C5OcWjmMC2
e3Cp5F2Ik8ILk4rGxpAZYGt/Ujd4bY9uilcJq6UVrm2LD3FbNab9YulJFDRjxasT
fFxeipsT0Z7X4sbz7TdVlz67lRvw1uLKWup30L5wNzmgYLqKuxxJtDs7syqLaItq
b0xf6rQycmzxKXnZG+2PqD6fs0qayIkHFnIZZiS7K0RO6H8DkGW5jc2sBFbgGTL5
h54+EQbz8iXw+Ucox2ikKJl/zIj20AnUAEXSRGmpfcbmVTDRyJzMh4hKv8C/C3UE
mOmMZxfAj5Z/kJJMTIRPYYuJRcHNp31IevvOUVNbLMxrWSyYsIXbQzQ5UZ1PlJGE
1Hr0vjyqoviqRxvofUm3EdANip3EuligUBEfvjd2b68AGg9gwmNwajNoBRoi7Ibq
oMQVekTrhZ033psyxnSleF3VzepQpsha14FjMvsDfmMhenqf9NLD2ZRZ/DoVruft
fH6W/nhv7HRCSit5E1QRf+Qyy7x7XuqDV0nBMih495cpW5UQRdiszgSVI+TlH7lD
Yf2OUApcQI79DDOGPeenlU2K/z47qAo2BDNhkWTDn1r/PIJQ/AuVlxm+GZWXPD1w
wiDHlFk743upSVtzOEBUfSqOLGcwXn3UjUSWiEHbr2wRhCE/s9Kf7g4ynSEcYiOW
q5FM2qrol0pss32WeOh2QOePzqRFHmVRGqCf7OpIYXzwJSSoUMrDRQyVpkVJYWkF
Fek9NJu4uWMR6FliFG8r+XJbsRwA2GEBn+8Y98L6YwGOSNQaaUYNeWnRrFBl7wrZ
CVkY9Sx1i+YeSWvMh+tVpbYt88vZ9Z7rwP99oSt15boyAPqW7IRGRoi/Rou7UTtV
U0f4neGtphNPXgX/wGuyPGuXr9HjWJzK9W66QJpOkqhuArRaUdxiHoHmrYJ3KJlG
a5t1lqkf0zU/Cq1WPqYGCxpAySfFpDK6SkIqFDb4WkT9dIXH0NK9cUy2UdK+Kokj
lucvPkAg8rASQctJrj6Fmck7L8VGJuVVpiV7Wnz76/tmIbd7DnrOQ9fMWurTPkgB
EmGrFsjufTNT5p1IEGTih7F7mvgHqTclQCX1wq1ubdkYJCHoAF7HGH9Kq+yDvMAb
er7tlVtScLjXG1WKA496h+Ro0VkF1U+w9VF54JmKQklaiyeEc1lQ7cFkp8nSRaSk
Ougc1GBI5k7Hu0cSdXO6iAUZDekxw5mpbrOBu9PJinlU6zAaMRVfL/p29QWB6v31
SjDAIm79+A+45aZkGr52LoGZiwg5MP5g8X8Pte+iwzVaM1vjW20VTeLYyWxFEMx3
8ec2Y7/7ESNpd/rpgwO9wuOlA0+PdO3AooGxv5+emPg6e0et4QxU8Dnz3hI4XxXp
3fKnfL6hjHVPN3RmS2VAysZfZlUZCU19SjIRaj5k41xSN1xKBnYRjg/a964zIlPd
wWYo/zyq6V2nR8ChpS2/LVr0xmVRemLdQfDhHNhYjAp7v2i+ChtXvQVfsvoJoTOX
BbPpc66NxaahR3IN4Sp5gCFJz4Uopq/nOWR8/2DOi7ePpAI1aZxlQtEEhVHsBqbT
dnMe3Irq7A2/RRFSv9PtRL6ANjzXTs0o/TXgo0QJsmwQbVBug2jMEP2mWUeM+ysP
5XCYGAiUY0LM3Vrg0DAaIPytpx4Iez4hIwkRNYdR49FiY8zMfC+WexPYAiRSXCCP
voBl4OEXj1tSFen3y8w2splitJMfk3R8SeX4v0tU8FqaYHIS+5MmBEsdxdztIyU9
zSqdW4psshMcHGSk/akbtnF8w/181RXA9IS8XMdivU8aa1hnIUW6lLcguUx1nJZw
YbhSjT4VqgklsO0x3F61VfM/vexMRYzfZahbxGCW/vFdhkw9eSaYhSevQoIPlXTo
CcAOBhK2QQNPet31aQIlAXyEbceqELSwlvjee75AjZfJ8D6F1CpgSstW1is/XrV1
uX41YPI6mkQMcXF4+jQDF07JVDy8q9Pd1V5ZkPIvwTKUYbwcAPfg1LUxYkPXdsDh
lUObrUQG7Hr4pJpXSUaMPhqKPl8nSiaAsYKOK1F+6ZTOzZ0+/xWzkKJfYn8nAHtN
VJ88p6pcepL8sIik2DiHzjFywRPXCwd++jHo+wrJaaHgQnmbIJBLiBDUtBssca2E
mdpsCfGgp8AGCEcv1j2Rcj0oUIo4pbyZDRG/wXxBlsAHBg9ol/gbL62jD0n65djo
VAcOSXCIzr99grS+mdaXs1Ii/re2aeiMYWFb4RWxVebdA5o6zWtnyphUbQy1Qe+c
s0cp3DrOVrkxW9W1hQ70andPepz4x3/BqunyZPp8bCibxypl1U94W2byZP7FoeCj
X/a6NwOyTk8/RCrbVfgbv2EYbNZWGeNktXO8R0spr+h/d8bMLRl3pH1f+/bQw6+Y
9oBYSgEQKVHjdq4sd+81S3IgKVB1ckEB2DgDAC+9exQDb63y0Lg7r1wObL8QLjNa
45igyv/1HSDMPQ3aepP3+ve2Q4OepGsPIxtUoi/oBdaoCW0QHM6milNSDnRmJQAj
5bJQnrZSZRheEE3+CW1ep/yomF+sZPaDwMZs+tSR3Ms+4G49LXqHrAO3hhhOr6gM
uVJILZRIwax5ME6TWVIoSaMyCCYVWW/uIHyc1YgMxkQtAQsyI87Z8LobEYcEDx30
Pf0GbJO82f1OWn3mi95SYmc4LZimMO+xrJ/eXn3ioZf6Oi8dy3TY5SGFiZuYrR3B
6FB688IJXw8vOmGKmcaK6ObSJUIw3iULfrJVl70TERT1VzYVwYDCCSc+5zwlYGNw
E6Edof5NGcVeSW6WaMrwpQduv1p4bTizt44Uj2pil3OqzKTHK4xWos2t95lKPhcS
CDSMUH4x9HIZNX9HGzExTKVBZv3LeMyBIim1bW778yelFM9UDw67uy2S6FYUmWnr
IVGiIuvxZSm920WDwD/HQhpOoYQfWjMIiHiozYl4mxhwmPQxUrhGtF1CILfVaarc
8b69AdMIcWdE++5cHlfDyr3AbAaKDE6WJOjY3gkLbIOoPQ73tuk4cO2VY1fRgmwk
uvAqbsz7IlFSDwm4rC0debXJPku+hCWZpiONTuHacKa9bHkcOMJX3mvRn6afVacV
JoUBIWGON/FPKsk+wmcjtuh3aOn59rLo+RvMhAacqgwYLhDgDVFz3ea+PJF+jMkd
DwMMVoFi6rYsy7OzIcPgW6gLYeTsYyH2xbcMptFsWcGZdzj0dkOPud0xMdaWFHS1
H8Xk44hTiNUBCefIYQP/DeO0c+bCKFbTO3F18XeFij7Av03VtHU8QJP8n9KSl4Zv
vCWAwAPY/+fUQXHRMWIc8OrQAn0suSKeXh0xk2oKs7YRrnRV/2uxeY+g/acta+DX
u/n6DuDMsZ5lywGTvW4JW082ukgvDPewfmgvMxCOQSCijdBgpUjnk2J2LTkZdqWF
rnIB6AwCdUzoIekQmfGR9vWjtFFgzKgiAbPx1/0kA0Zg+Y9ivXY+sJ0s9Tow43Uj
+OMX74DCQVpcR+vcA+nki83pro0IpQmKT5NP724qMCh1c9vOSpo2KayghEWKrXzx
jB2qGdN5wpyxgpfz7IS9Ztu3s9rgDW15lQb4vord0eZWIVPMEMs0V37UgVcfhsLg
sTf7ZtMJZkbVM10+3RXSxvbxGbAwZu+XcuvxNXkBI5A2Sjk/pVRdpu3GqEwaQytw
WM9y7I8Urxhgbmtn8Fjg8Bd6x7qiEnYatM8VmVRiqW7+gML0kZYywY/eZ2mw3zVj
k8jH1Ob5SMqno2LONOkFmH+Rfujo7eq5bJk1Do79fwAYHHrxiG7iBdMD9vMbCnCZ
xUpqqToaI/wPIae/kwrt04i+0Ii50oAOYj2uq20LSyNV5G7e8UKMu0TVpTbi3Cls
r4NTelwBeaWvlpL0ckUQy9AwDTYdmYSs+fBknHQoIANT9QV4AD7ArJxYskgtL2vr
QYFJrWjwq0skwrVPdav3c0iiTniNX0UUaFdjh7FQH4m7VhM68iuNOzxEQoXMBkMi
/cs9i7C/wkAeAczthHr/M6D5nxYvvtDmoNIh9DH6BdvgTJ5z7/JeICQt4jZPsEC6
cZg2+6+IjgJ2rFOmmxLRWk6UvZxbiQwu/jQqC+LmaG2XfxNu9BlwJtJSSUr7tU7R
tDXGIAWOaix4SWuW/Z54ZqGu7Uwpvzj05xNEhXuJN9+7hHeLThI8TEbv5V8D/ken
boxBmDkgzWD+xq/6ST1ASiGHBGqH7mdxZIZ1P2TuXTU8KNvZkteAtT7Y+h03DvGu
7Ez+i5gl4TAs/Vu/3tTAIXVS/L9cKiGqkUaDf7g8mZclURS2ZfnHVtxSKiSGjAjJ
phQQLdQ8tHIuRc/hWvV/blG0tQAlXVgRI5I5oxKy0PrdcBHEhTANLp7ad/MztUOR
GS+UvOIHfPmawG+cdaVMSqprBm7ORdVM9xrQhcX/I9nv0Zy/XpWF4a06QZFENaTo
3wEgsy9aF4LGyZJQa6+da3xUJJIH8hqzQ5g4DU+Byc5eI/MBAyH/Pq2ovRxMwzan
k8prBguBclAHLchQC+MKO+lUBgPFMRYhefaZcKxmQTlCDslt12sXHTqsPNbeMDH4
XZEEUyRU1t8pOzd2LHI09Q7GmVwFZDK3UsD1w2rBF/zV2tFsxJ0oGSgTPCw9ZuTe
DJ5I/0cyDjYGveK3fqvmxIX+8Co77dJhlxQL801xhqg+Zm0opVCrqHKymJx3KAQQ
LLQFHNdYFnQk6moVsOuy1sRt2EcjLQYLkmnMZwC441iNFRII2G7xeAC9P7chxwmZ
bOomFNaOsYgmBWpr4KMY8d2JCVT4wr6uVVMyEjYa9nAEHRDbwACmmRRlCFYvyGel
40YFaK96pvcP0YLirSaWtlIXNgg5M7dTm6HmS57HhgBDLtxQyoCgW3Pqu0cJXw+7
2PD22U3G+wLWJO7DfzzhT1JgSVvqqLQFRyWf2v0S1+/pt18pCNqJVgDChSA7BYCP
dHT1EavUVnl4nNIfK4FuTFucoGE98n7+f/Nb0naJGvk5jYVb0R+Rj67R3Oa48A3A
3r031Xea5rOzI9gGYVKRITLClw3twZpDW1UjIbvJNga94PlG4mCmjxcRk+q8HMGL
/4EZqYKJThD9Blh4cngXwmYIwoNP+kprbKZ0twYI+tNTAOWgn7fBTIAVWFC6P2O8
ghBmRwxiNH/KAOzd6V1mBpDKCS+PifFFiWWqEXIsqysEMXzL7ydzItx1QQaE9wyC
NSay3GffvocsJYtaO7hV7OWgYEtk9TUqVCGA9w5FQtzALzNOGfIdE8usCCabPzxd
b6rzJ0i+5Umcvte0ElFRjrTFd6qqO4HJ4+xYaR9BB240bnwX3m7c/PBHz1mgYIZn
yzUNoseGOthM6SqguAihiyZz0hxf26d/BJd5p7GbhU6fOUeMb1Q0Kr2Is1rH/PIl
XGApRPwgfgTyES7P+Yz35Brz+qKa6BPopXmDjcf65ZQr1y/opFlM1tQYYqLx6CtE
QP8gXyxAtxnwTR8JDNdT0LanO6KuUuaLqrM8/01/HMR1E90ZACK8IAXIxAeisLZG
eY8LQITMig5j9PViepRzmhjStCjG3VREKvKqePr9UFhTCro3XJbeGz/ahp7YPuL/
7CTrY0Im/GzeJQUjNQAu+JaTHJRN4sVV0WtaQpj8xNaDFDDsIQte3aOEHn5uU+4M
G8248OE2NRjAtHpl8zUqtVx8LXdcC+YQLrn/Rlq6VjW+INZaf/NmK8CnLgCdjoRh
fMJv4fUQ78GSmZFhEHqF+e/MescvD3LbhZPfLbam7CBXNb/zL5uTXvr/B0zf1iew
xl5RpFwQmdAs7OkymqiAcqJTUnoZ90S6vC99PeGMXUAZ+cVeGSxBFWrpcVxigYP4
OTIiwMN99pIU6JX7C+21kqV+IE03iKfw6EV5OHnlq8U/eA3dhrt7g81ZLtRo9FPB
AfQRuf8bujkZTiHn5Udv83Nt8oY/YsBwnV4Dk31BACIRSAma4+9UW+EmxcUJ711+
wylpOFiDT3X/+euN6dmPG3qtUgqnqQzARgmYK99Hs4lfMK084GLOdpl4wHPE2ZD3
yQF4hfSUrePpB2QcRgbULUeNM1ly3hl3ZW7dN7HzBpf7Zc6HN0/VzYptReLXLod8
Y22QcFOJDV4YzNlhL0L+DCWycLOrrGx+gzavu+zjfEdZWej2ddbre0dEuUSv/Yol
OSzu7bAreHCWF8t4AG4bYSoMDxyRdYm1gicROlYS0vomU/C7t28qTau6X4gfuEJJ
AmME8V+S5ERmP0zLZQDn6wQZLUVx3myuZ5FiDGEoJpZhGJS6SQIPtE66HBiOWYVy
wFDQbOrxx1cVfFmKLBtM46p+nalbTPuO5c/ZtoJqEMafqdumxYMmAXXbHZcf+96Q
JjzItMZ9ibr4mAUfCZiAzfbUOARmldrf+acTfGZeg7UlaahJEHgeEYvEex4YTZtr
xgI2vbpDN8fi8TfiGakqtdEmoF1jho+KyYGEmeinD3xUoWoT2mwWvVQhAo5sDjUm
pbX5oF49/yQZsOEs1IoYeH3kfsVkVwpIbpDeTEx7CLJJYUsN2lJWzXShPKdb2Q7d
kgYikWJtfejHcWXgAJc3izc7GjwF+OJ+jBjAV7T76dgfBzt1oEkCNXlH5h1fPgC2
d3Xmqf2G64J3f3w9Ah30iawGNaFMJhQXxtVGW5r3XnaT+0CwCbF4J/Q3MAAJFru5
sDJVAmFDcEDbZl+yvP8B93ISduc39zGPAJUdrhuiWzd3HszdjuVR+p8X7JVTIQsf
NaPffjaeytzScL8jXoOk/HO3ki7PDe+8kiabzZ6KO0YgcKixhFlDamYX3D6BpKGT
JTgEaA/uJxK/JLYqmMA9eFW65Qkuogm9KxiklQwloMQqCgtVLfEAFbWJK47V7BeE
cwuiBrzBGRMfvTBPAoOVfEcGxidjxlzvwoh9J2uYwyKkBxkssw7LpL9gN777wjZ4
9tog7KQRwXzugTvRUAspBnkSL+lOBTR1+4ZiDprII4ayYwKmxth79/hTRtnwUTPX
kRX/UZL2HRqqjPdauOROFs3LkxIoKruj4AATx3VKdVQOLTdd2nnb6MgTDrBYTOjt
JVUsPJj0D6Q6zkakdRFdNjYjHmbXpGMxIRALQdxstNmP+geXM3BjW0M13mvedVca
D19vHmTM0u5B+72Fh/qdwsX2bIp6/+dHcD/QhG4bSXtKzyzSVwO6uqkti6ZsU4jP
u+qeY8KBLpOwlFSwA0SCyon0TPcmOiayqjscksl5QaEgJ0/FWgekosOroOyT/h2n
iaUXFmeLMq3G8m8t8UWU+l7tWv+eWJPb4OVbHGa/dHHaXIYUF3ZJf+pR2L/Ph5bK
JIyEmwrCdEr8KZPKTWsLun1fK61nUaiKDSZk33RzF6jkydMn00VZa0eH/gylbbYq
nh8v4bmGGbA7DtCak3YcouUkBdw4PSwQJybbrEzuK3cfqRBGo8Ie2c8fmP3Quhwv
AXse/0U/c8fAJWKUVZ3J5dIvVlUMcegep+3aSGMlpSHrwe7DerivH4ba3HaOAzUt
fz1v3MYtOSgWKb2+bKrwq5DY/LAa1zjozJM4pNQhnnOsCmfxj6B2uQnHJWQnUO2J
mYtbZu2bqhLojI7lQrLXOrPFLNohQRN9ync2wYmzk712Ij5/ykYF4YFnH3xkjDVE
R4FPzuiHBeScOjB6XXl4Dcv6oI8oDEvcSkwDey3BtoPx1bjTLwlvdOg7DgO5olOJ
V3xrrFPAGsFmz6N0N2CFv+VuK5Z+CiiM5DquvuNnRQ/Kp4Q6kcTi9elUNk62Ukzf
2kR6ntHk1JAXSA28956ZMhz2MsDfMMtqdzbLR2XF5xs9f23EqAQlyjIlI85/yBAQ
87vcBnYOog2AU+51sjgkQ9opsHG3gLpDzk7syD4bhPW2PzgyGSOmDxO+6ZOCQuYy
Wc/Gk+qW+0e3rVTIoUb1CByrFxTKLwsWZZPn8l0Au/dT4lUZ51KMAygdTKjN77tn
/t8ZqmRMuSnECr32qFBZIIOmx7izgmdTcwQNnIbeWbfw1Te07mpSi74pVHNN7imh
wSjmmCTDFRul6LtSy+7hvfA7/5Y6JR8uOI43BVDXiv71bVvWhjnTcfc0m1tgDEvT
s1MEm7QrRnyHML7UTy2q6lKeIsqIA0QaIHGXKbhIaZcs+buZdBzM8K+06ccYHb0J
bOMzrm857BTnfbJ5vyGJ7iuKjQGTPpLTqlseSmeDOswwyEJXaXYQMt8xV8qhWlDe
YMuulvDH/VNog2dHjot5JezITrcagTr7T64q1k1PdESxftLlpulQOobLwAYE5tW/
8+ubFHtAgvAZHpAPI4SDW5HjlGgyHFROR/x3PMkLHGsMqcA1BsXp5LHurfkLD3AR
NWirkA7jAo6rUqldud+/Jm9OpQpUBrkI3j/AGY7SJ9EEPOKVRd7I/hsexPuj2rSV
CGTeBWOD4V2duYbVSFaReQeb5xcD/EZtaurKxQjB5AlbKMY8KjbGXJKefxjV9T+B
zPS29bWqt+wg8Cno5YVAVvlZQH+jrVhBGIOSksqmEg4sNc0AmoAbnsoMYGJwMfyh
Mf0o2zMUpalNgS4qD/IH/nGqkyciB8M2EBmBQhM9iZpmxxEDzGAHEY6+8WMTJ7Ap
/2gr9NRZ7uuPOTV/iLbDTZ42kpfBCeGXAcufXIbUKcn9udUZHhCSNE8NB0h0Y7og
PgDfyVr/F9LJT22fmIX3OgWZo1boNAfXCrwibLwckTQR/EF1YcV1OgkpZGxxqeGF
JAXitc9mzCZJ/e8O2StL8nWWu0eRNEU6bCaVW4k03zuNVzevYI2Y6rs3w3r2p2Ve
uPSpUKyRVqZyi47KPoB+dIomQMEnNpp5ijROOtemAWPLX49n3H3ipJoisK7ZM0CQ
pV4uzURkFdHYA7MaxUhbmHFF9anDGjW4JKOXu0jMa+kEQv08+6tnA/HhEHAdL4mF
18AeEn5Dx3DMg8eG1qmhYlOtqi747k1CtitjWRn7JE/rslZk3c7THsuOpVA7tRkC
kNK2p6CrhtEXeu7UxH2vQHX9GP6+i3ew9FhOODjLPd+U9BNylbTixJ0ij7TZylFI
2SwgKf/PVQJDlSKmOg9g3IRcCEq4EnDFlRfBN4ufZsWnDTRTCTME+WwLa10bZAt0
UjiQ/W7S1Svi+Ule04nh+FrlRrSXCDsp2QnwYaorw/NNLGk4LccPW+fgfWxAuVaa
cbbJDhhb+eAluvE22hxZw/qinv0mfStNQmx5XFb1oa6FELoiyrZNGtNgrzxe9wNj
YOcT2BRxgyg+MOrySXoHsr7OybPwYVDGyidY/lK5c+uN0PE9HTcJQWLW3gOVKOW/
MHX+d/ZAJFReZ4hMN673BODriyzzcVCINYvJxcQ2lYpbR2hGvxX+BqdTN9bHeyFz
2UNjfxtunMw0/NdSBIwAVadwl+aPhiwVkQSMIW0cpSTRq+vVW3DUh8pcpKaLeEf+
eMgdrYMT9oMROKOR2a61bHoOljnyCYZorvyVvsjH7KL2JoCd0oWviJWlHa0A4x3d
PT5cjR3Bm8xZaUjOX//QG1WGPYnueeo2II7ynbHR2V3AZs1l8emFXI7Acbfwdc9Y
my/73NQ5aNLQ5VA+VAnCUIqEWXfaW6SINynjqgsPVm3Yws6RdWU1CFT4ZfvW8IOy
ik9k6QAfmOW4YZPQJs7DIkkRDcFUUOjP7CzY6jjL/ID/GMTTAhdRTrIjgRLp0+wZ
ibJtg2wmhwl3XAFKLn9jUoHShrDLZO8UAcjs1WFb3lfejW147tu5qedA5Tbu7qH5
dZoiFGxEvsTZJ/iyZ+JNy+f8IQPIsex1BLLi3JgVq36Cgfxv5lojlTTul9062yUo
nnNf8VYOW5aF6RVPA5f2vmr4UQ3Q3e0BZ31BxSGen4cgoMVnc5gN5DHbowXfRGUq
2OiqMuWwRQncQMcFm/SPN8UeQ2h6fDAKMR8wHRYGqz+Fv6GfyHTDyyAVedXB22NZ
wYVp5wlcx9hOaf70mPK7r6wd43urz6N1xs+6yN8QLfSOYCqTW4gFUtuwITRIAE2m
AB4j0QQ95dAu4YvtwG8rInQ5ATYoQsZzHV+bKQvsEBtLNEUM2dAWiKfSib7s4fVW
DJtpCo8bn4Gqbjv3XpjTHeEDxo08BTFNus+nENbQAf6J5t+b3dh/z6tDdZJyjlYP
uNspFolqxpYt0ac1t/EIXa1Bmo2CLd5BO4tUXz7vRZTt5Qa9N58Q68w7IPtlF5md
GZ0kPe4pEAwlwxLk0+h4psLQnaS7YQgVtBNDEN0ShDJZZ7RPVXTm4TeP4XAmR8HC
JiOPrHevl86cmrwFkCMYtLGHf7DSt/W9xvsyWpTEVfctfknZ4GBSyGWhOP3tqFLI
nJ8Us1c9jFoRbUkODKIL/j9YfD4vPCQu+2Xh5qbKjMKXRm2mH2Kkjy4M5Tmc063n
wp9xn26z0DayxejekTfUHJTyedpN8wv4kYVBTFIrPM4RLIh4hL83nM+ZvBDyaFJc
DpFM9R0GJIfLhc5Paq3rvLPmQeP3TCULYbn09pdK19OyieIx1TQYlkqQ7lzJt89F
aQr+v4VdJb767emeEPqfJ97OHaCXEBz0UBL4jRENOZDqekSOkFHUuTYnKpMBUriZ
YNB0alw6YNPHQwu+W+vIkafZG2WxRsy3fA+4QnTJZJXaGQ44bQFD3L+zEHh5+8j9
xyF3nzyBFeYR/AXUk4kWTMEvQngKqXaBD/31fJRCUpcyh0KNdsK7LYtqBef420l7
NPiyd+CiEdd1fBUSHS76AX4aWUqDglQezHnKc8uokmJt/hXBaFfGef9Nlx3S6fTK
soQK6g8QkTy2ncUOiRqBUOF4ZNISpW0xh+88LZ4S6ptPPIwyYnY8madc52ZMDrUJ
YcqLwBII9ZY4j0enqT1Aw3A726DK+8P8hxQI6sfttH9Q1eq5PNjPgqSAtlAM0x2h
BUbeimJXnIgJbqP7QPH9vyl0JwUEY7CcKr2yCLVmGQ1N1TqxW0IfK+ecutAa8fNJ
1Yh0oEjBg+apMg3yltrKM0y8tj+MPyqtL7yudBuqaDF7xCaHWRubVWSlVdHrKYcf
cicBy5Y6G29SUFBd6gncova0xC3YyVdg49EjrAI0OmokCdNk3R4zKrIwFVtayS9A
RbJlDuAFGYOLccLp9H5OOON+QZRrh4KdY4U375pJKr+aJIko/63dCC0g6+wNF0CR
HAo4FEeh5810NfwNxG+vm0ODR62ez/tRU6J/EjI7hcqH3vInLRQ5bVbHkcuqzu4u
DfQWIw9vvbdwWoi+irccx04sKr5j4bT0oo6Dcg4Gmdp/K66DGwYeGvhtfSJnE9pI
VWFjHhOWkebGFKgOXynCiP33nHf4Ya3zzM5TykmmzsSc+m0t349iey1tE8GP+e8b
9qzvIBvtnSRNzF1e83S6ssK3xleXp0Om36fW/6ocda8UVCCI0AELneNv+YUK11SS
SNaLoXU9A8t2Fm6lFfRKG5wO+gDxWfyRezIZXfmoLP/xppf2Jk25qGWtizvSR9Qt
35LI+ejdo2WvD8h7UeCrFe4f2EIb6JGAk/q5q2OeCFsAe0pEGFxWiwi6Ly1+/Nh7
GzFxbJTs1AHowrJ6LisvvfRhQG8S/zQtjdH2EZyE28wWQif0GQbx6nuASINFTLsD
TGVCk8AvfDFUTWWqsu2g0Q8Pbv4o+qr9qkM5gQ+T5yo0I3NFaHdw85V7JJ6HTmzB
CKjv7flcj5isAvaX8kKn8mX04GPDpsrf2S6gkKyFrOISpy8u9SSzvKwSKdw/wv81
5ZxFTx0zbO8hdEXmOZWBOpq/fH8ndcrxYpI2GpqHuVep4sgC1/k2UPB7R4nib6u5
nCHaYpl3/87j2vpiTxBLgtlg0sRYo+ylYGg8LK+f+OYzr8PAbk8lY6oSmha6a+Pa
wp9zHLlln+xHxJ1NwIWGsx+0rOe/l5AgarM/+z+SUrxbMtCIa3PPmeXURKXCQJrF
SHOaeE4rpaBcHAICDvYSGTcD9STX7OcXWvtABSROpZLZmSwXGhvAJ5wz/HXeD+2k
wewx5Ya+1jJdqOx3QNiy8ARmvUajmaxQERr3EpJWjXKvp93KxoHNaAlGyQeIkRsa
KHAoGoMUfwgDftc2hpo0WLQ8Uvd2GBcE9zFgx9pOgSzYGRIa0TqzJAYjFTuIHXmr
HENC3LUpN9a9opi/ZYrh7WbsULxDyaWc9urHQ4HtjpCmEzlPz26pWwYqjJj6dAx4
qm3R8Htpw7hdKt0B4bttQfUp49/vLudqz4jmOqRWCVvsTllPyfHCEMBtDaM2qkS9
1b+c1nvk7fz8jL02ihYgczCoTyt2CHfu0t2XG9B9daQLi4zCOoAhIIJGnAfgbTbs
vizKRYNT6AncFbzMuO3btri13QIIg36m9foSso27TZgtIARmiByyWQUjARRe6MCI
FeEzAF/EnofbAVQtBGZnFqlWerUXrrzNR7R+8FV++lxKv55wSr5DTKcG/J33Kdv2
ie+dGTxZ7m46SdCTfLJrTfx8bLR7PrDKQObs8QOxNY5zF2aWPsCL+96FzgZySdpR
TwznFoWYX+Yy02FChvIp5NmC1TFH+sefVAUC8D9W8RilfcdJl+WFyzXhmbtYfn0v
QyIZT+MNQBmq5I6qYfMg+/scJ1oy9obB18AeSOxixAelxo+3Bqv3VWydAwlr4t50
EgV9u4+VZj40gMAF/kcaUzDUS5Gz7R6gqP48qrONKF0jwSX6oLEE76d7w74Rej9H
6D3zM4VKieHNYMIm5wqe6U2Xaoz1nsiug6SEuWdMt717KCa9u/lcEVZb5DrdGdtS
/nmnMq+bDGnc0znKXIAO+K2CQpaEYJyFitWZIa4KDxOOchmmao7t6DatBZAgZ+J/
D9MLfU/F6FF+rYD6WNhU+DB3o0loocKzuJZX/wrTrsUAWwq8kahPA1uh86FwtmfD
rEByLepV3sIrf55VmUk3nRzHetfgSAUQCUP/SYAPNtQfkit553r4LpGmz2aewJFP
tpQsO395kvXKeCa+eaQ/Hdkp9gzJXx3jZLgN8uLNb799jFXSDix/3oSMppQMvyKh
zoeBUiPTovhs1TSeD2vU/hRNcsnQtXpxi00LtaLxZ97wTDvD5xmknf/wHRRAo+dd
o2vbeSfhdQvPSmNHe0DHjoJEvvTSxCvllbqVNqw/ENcIKmn9vlwzcTnKfQAv9578
6Kg5IbDf0ksbVurE+0c4FOgBj74xuo1wXp7VK9z97F8Xb6Z9zCLNEroxAqj03JTs
p20JqE3xBLoPAs8+oXeMm2gcmW6AX5DG2f+cheC5qO4lPtKd9Jq94NHwBq0rV59z
VtTNH+IihuNYo64hbCkgoG0ubMocslR31Q+H+bKsEPHTBXLMRhDDiZfpMSoVZZdx
2BopOOopkDPN8bAbPFoaS4ck4kG4J6i/3ULLg59gyy0VlwPAXVGaPQm2Eck0sRff
krC3VipfhIDlQnBZaLj5CllgitsCU6infbVG5+h64kZFlGLcbtDZgDnyH28p/WI8
S1ruzT58EZ6D+v81Cjtmv9pYZDiDBnof3n3++LSBXwq8GvkXd6i8bZJHOklEEJ/7
ZBOcEBBgeiT6D1KhyFfWYchD7nxUZWo5Dk3cETcG1ZiK79gqEL0uxEXLG4MUCFWI
1G4FvEnurPf5D3F5/czD+K/fK5vvyHbDryv+iK4C648icD/UY4wbhiylVrVVqCFO
iTc/l9AndQRO391oZfsk4O9D/+G5x6be5spF8SGzfiHpSLjH69FP1DXuQGAKTfku
vzodELNZyOa6LP+2OPrVes8gov0FrJk5RmcUxgQb06+fFhKr0JpKMZO88y60z785
t/0bTJVhxL4u5eFwN33b583uuxmAv4RnOAXGj+5l0BzVwWRLLpB9s/zJymiQ4lhI
t3Kb4zodrXWNR80G29pl4b6pgq482crdDNecvuBB9zePeiQHN8zXtfXs+0cqasFu
L0RVrMWdwfIj4pHAPTMI8evhguDrxO1j5g6suSiqZGZ81pDOjLmY9ZDsFvugM52+
gQMnaaL0QE57oKUAemQD7xsKzKeklHPFTOqwx6Ibt/mjvq96HYoLWzV4UjHfgOQV
aWKUDURVa/cKYfojQ+9nErWjfo2fv1m3EDEtrwjHIvX7hUI1CzbsOqVxjRM+6xUe
gRgABA4Ir4AoF203dG4eWqdG7yNaWuavPKhfDXp+EfSgxKecOl88YC0MZSO2qe0H
HqPq/5Mo6xlWiEMAvTHs596JdgMGAG9NTZugB9eJZUEaY5PhzhgSJP5aTjVE42Xo
BOG8VQrgdivEe3pRLjqHKVRJqxAwudAAS/cI9yIgF0zu86wAmpzbyJNk7TqZk08o
U84epg6jFa5sXO1yhQs7AQusqQQBcv5R6Fc6UqnblSTmtmwrZDsPgBNBcZNpZqbp
3e5kGMyDDlgv8Bm0wzt81fMWRqA/2tFs518QINXmDGFpjGTjVDLe27KWS1mhPmKB
ar+hNOU8zRPH73NVGP9IgWbQOpGY4hiGt878Ur5OiBgqbNTZKfrXlwkAcnLDpsZI
8amkBnou7cDlbITnSv0wpIeC12t4LZ0RafEIz/6mKbyxGUdkxlMWVYLvh8Z58Hx9
wOBuf3AFYjn97r2uGJjOw3tmqgv1KOJrvqC1SzKSQUPV+DjzxQxCiOeZerc+Bh9A
b36dyVPBvW3w0bhlYEF4y3R4LSR88R/xF+Xd8OfNfoiVxOL1Caa2nIdsWxSQEGbM
QR7nKgxmOz1g1sZFTIwftMwGt2qYoA3gwVUEOL5s7W0vfyqN3bLsYG/nA3P4z+Wn
H2fqJ35hcV3GDCm6Vw+tlBqP4D82+tVlTvCxYhgdLSpS2p5Vqwq7vYJR0iboHe0R
Kn0MsmnOAO965WqAiGZNO7N6+Hc+5bhtQwnum/yi1SjD+BfTKI8wqV2WHtpMUJ8c
lylbB8+0TbHzCSlrzMWoEyfUGIHxclzyXWGTbjVku4LIyatavcWKW6bJGlWghzAl
jEoEzhTzT11X7+NxtcGdM91x00M526RtLl/mhviWQLucLaoA+WqqwKc3uZsjpE6C
t0tvcjJExZ1Balto0828D+NqpfnFpeqGMObDFIm95kK34qKuGgQ7ZV0H1Odmp0Ca
MgcK+p3H9Axd1rZU68Lb7MWl8S5jz+RMHnrEMRXJxEawH8RtIqH3X86VbQ4O71Lf
s4AaKjXrCgub4Y6K3/BdJ/9zCbTWoCklivr9aoFMker/L69ifGrTbk66CyQTlzkl
ziMsFs+JZFOfVwCU3Gd7BeOoKA2+aRzpR+4h2yHzVUyYeI1WrWExYImdhqwkD2t7
2JvwBfguQn62Uie0q5xjA4RdDwtiyj5Uq6yp+dslE2CH9PVW+4X69IuJKwDYhz3G
ww/ezzTGfXTYJHr+m68ewA8Qg2MTZd2WX4lsKzcXJeobaUD+pncIMz2ta19f/9R1
RZS8931zxHyGLgv/L0DGrfQrFmgZjMA5alyTSy87anCIqwFufM5lB22zTFYK0lKh
29qiPXHbVndJSEmZS9dh8zERaPzSutpVLw9FbTKZkPheYzx6SN2O6yCxgMmDxukV
v/P4lzx2FEVx6qNHUOBYTeM6+eHWyigl7UEraOMdVlczVtfUBPTruE64+aQEsIaP
KPBObbKPvtbROFXAa7NiOscoz8ewNS+g4dwBZG75kv1agdkmOrL/mJDw+rpi8M46
c5YEHS0MKaOnlzvaeIMFQ6WekmdR6X41gpYbfJFdqevJqQ60Vua2YheeLydi+5El
07/q/j21GkCaBwlhgUD4ixbz2kOJ5Rqe3PIfy2oTkxVpJfE56+sLSieeOT4JXmSK
DwC/NvadZqJsYs7uvW0h9svEdXeThz0paMlo0e7sf+fsjfPBs/6ITeVFMjtDbivk
r+LtBoq42EAWDgw2RIUXeIvBc5Ud+Ay2vmf0Bsum/+8TF24ozhe75grtr4qNbyjL
3+d7pQxnoo6b2KJj2FHPUShEUO+b7uiiVX3oTNX9T01C+t8EjPH0XML/CnLVdVAo
vcXJclKIYvTzoR03A+gqkC4zz0JLH/wRbzNOnCVwNmK1BVz6CY4zWNBy8482k4fP
6skPckpWr4ewE+KBLxWX3s7/ySFbir2b0pPgV/gUwoj+liY4/2zdfVxjdtPNjOK7
YCEtswiiwpfZX+jemmlctaaKipYTDZJ43sUDd7NvZj2d4Q3V5u84scAzbVOiEOaW
iA7EUKjhOqvvDSGH1aqj3QM6QR5MJ+gUUCuqSZsxnENk8V7XgrtN3kfNp7ZWqzdw
Ds56OyK1P7DUUKDEVC+5G4JJdvkLiFqFATpdd5XYOe8MNtmRqEn5RnFF53sZrjS2
hEbZSiAhF19j0Z5DafqmHUdgEpsD/CXUIPKHi4eeJKaYbWbU7VDTd1Mj0bmaLy++
+WQmC/jv7jRiua1TgXSAGJ3IOUxgjnNu1KUlHAa8eTZOw231G1F8taPI8bAjRRir
FMqsXUm58aRm2YmCBhnh7T0GS6a5/VW7R0xHr5tb6OiqrAFKebU8BHsG0U4K3UYC
KGWvQvMcDdRBp/Jy4JmPwQyD7MWpKAuNmBxA2ER2vdyIIa3BqyZMlDLe/sVUeAzd
RqP14TPRuWalbihpPndoXED8xUGwLoVNBXm81FCq4/mC6IwgBqqNekWClw0fPv7n
Tgfcr1OSxUXgm5XULM4teDJ5S9BheFGvozt7k+hJV9+X+Xr9kgtFIwRGfCXP+XFt
4UUKv7m/HNVVf8TYL3V9xSrYqsDB9otzYTBf+DaT7O7SBQc15lt2S0E4TBj5Ghtd
rBDDEGRwvYogZXvnEXh3BMcYLfX0r0LSKWBnR7DK+TNHqMyzUX8hDaKXNDlmZ/Ao
UtKo36NIgx6NBk8Ifftl+FN2SRf3SldgDP57mIFeFT5sF28SSqZxYOFv7zdeIBAa
OcJflgNZzGCkt07xS9f27ylpV1wi9dRf2OADhLuXNQ9CL4ttSYX1b7ORiV77zH6C
WVnGPgq7go1oIsXLxBbbddZYJBXPNc9TQslibnNO4ndJ/S0VPuroVZXCp/xyd1+o
O/GNf0UNlivbKPMoND44iVEqOa6+DCbCFX0yhUvMeTdt4WpOz11Q8cFWnOo31kEA
ad3rlvbn2ePywwiF/fW8zbe6aaPeQdftIz6IybVZNpL6FigJnHIv8NteYiCINGUa
5xVOA7cCDGnarHXZkFZgbSbD5fY3oCLNF6xDsjpdo4ygNho9H4EZl1pWCKv0FPLV
Ml28Fim6c6fSuOpwcDIeUSTu8EzTFHZ67SZ31aDU+QSq0SHgcrbBJRPE8BDdQx84
xhBGBSyyD5HNAK3eJJskC7C8pu7ybxFO5l6o0916ErmtbrH77bvQWgymxANHY6Fb
LLKUvXjdpeQn24RSPDXDdS/qkYZOtFRUtRD47vamgbI9eSYOJD78bUdSSdBXTYx0
5QXhTlfj6IxMSTNJBEsHMXizkz8yaCIw4TqQq4V7nCakPxpOnaK8qScO/rUSRbzu
bM1acq9OtgsK698RDog+AQc6oQtikoAzWjyXBc79bX940XA63/ReGyPBGGYI5rXq
5aTONxuxAxm7NtRMx0x2JQOLp5im0tN5//8uZD52Qw1ewhfoDOi/lrZaGo2Crq6K
AGzRWIlfEVdM5DUBj53KUnblCdxM1K9E3J9fZ3nM29I+krEynY+m1gODMVsEYuuq
W60Qfnb5bDAAxrgAzD3V508VVPsib3ivNC9pN4q6A8BhXYAcAp4BuoJWbgp9ihoc
wuSu+iPIJ8K/h6NcrcvliZFgmQrUo2rmWnfLSkxDM08eZ2GXAajkDBjSxFnFla+l
I5imhFt7LUaRlqTERP20uCSydBXXwc8soVosbATaQd6qCu8SOpFP3snp0uVI/OXd
t8E8m+KVkJxrhypoEAITZWFh7LUUOH5HgOsb8gv09GRFy1tKykmz0lbFRnCcTx3g
T/iHl0G8UPou+TjUOspufXoaE/Td5RtjV5GcWANlWJZs3yotfQEQV1r0QTyPeHmY
Pa15RAqX+DTabAk7dIkKGevKHV9L4TN7axu2SZ/F0MeWIKXjwHvG6ReVJrRZ82u/
6OvQYFXRWqBaNdft3LgOPWZLMNEGJr7QZccPGLvxUoz8wtEKs/OcelsJrM1lxFjk
kL7RBq9B+gX/s0zhLYhNuooW2PE9JAv3WUhB+L5z+aZT5RRBA/9cpIgobtmiqWTh
pJfKVUU/GXzcAwoeEVxynXCsjuYYPxAmqWt/yVMNFIuWL2TR2PLe2xGsaIPIgvhl
lw2/ofadOW5j71yIEJBtmXL00+at9o/Ap7yLiqnKk1jzEgxbOblMo6YpAcOzsUpE
6bRhfoq2VXO2bDGAlnnKipy6JZS8MB506wq5luCt4x5wOrsa1DvyKwRWizbdwpiR
l8DYyNXEy2RYkvqIXLux3VCeHunvDkx+Lk5IbcpgNsDEM0GgLeNsQzYDd0qU8LXd
21x0Qo6gCCDsGR7BcdLMXyRJAobv/CCpDnRlLBjOwv5jwvqM6+1p4qaSXbpKAFSt
Rxd8lL3lncj/LVdg1Q9QZAqyLZkVp1qFYh6muVpgmhHxmRRVBj3oloGHoWoogNS8
DBraw05FeJncNYCjM3tb184vXnD0ex76/VmHvjTp8DhCeyrPbMUt4bp43ohBAS5D
YXAMVimbe56TN0iPwIkRb43KOhEWGiRmqYXxiusUIaYlMpXtvraOzHv4L6o746PW
iHmYWK+5EZDubDvJ0q3WTV5axrlow9mHeMCzMk0MsjUC9zPceeu1um+JZsYh9D2n
5G3p5uzwPGuqwfxn2v7nSQHTuW7/gXSXelNVlIjGH17sFaXoi0iLXKnKNKdGAmrW
Ce3RiQitwz1eSMuj4d0JQmJxhHN+1NKt2yaZ5h6dPijYGhJtnQei2ffHMlFMHaUF
Q2zdB1vG8s8bqjc0j+7eHdIlYOQHIeKdrRpdvzIkCEzyj05/sy4MVZs3PBASvEHd
CzGGR0I1vEpjuYE102xve443bKwZn424rt62po7eB2/XNgDQh6u0fLqAh7Kx90qn
gvRmZRR2bwOhmrx8WeJZ2nsocH8vf/z9tnqFcSBkv5WUvcGBwIdnwKzAi5P5lxDa
wN+HWOOMTPBM6J2RknVKFKUQR4/a5BVIEL0/CYfpNtDo5gkzsY5IvuqqFNyn51bd
5uK3opPRzEMiBQPo1/cB5t9lg7G4mHOelSu1IrMFVQt+nbxlccWP/g6tpdXA102u
6yoTcT99qqfhebDbQwJJF/bTfux11WffE9iY2/ck/qSHQItthBQ0++oifoEfRIlB
xmLL5S4YwIaDHe6me5zJPTghgeLWvg2phuegqxsy4580aKh8Ea5wzQN8yLoWe/9b
1KnHpzgkbHiUX8xraB0hXHPkaQ0Bd+lexD8Oyck4wVV7qeCExgRVJji21p0eril3
G5X4do6txzpddyKtZWjZtQ3W01+NNySo1R7im02FMN4SbRe6cEcae1kcTBfYSNCo
Hj3Ox6f67PwoyIiHjENp88q4x9mkgtr/A8arHP2PT/KpbqVOJoyWVgXMW8unUj2i
cSgAW0f3N6rmwT0vzNiylpdlfRhiB1d69x4npumhnuuvxKPvMj3xssNnYFc/1VN/
8VsFjX6VHV5lSAAfd3Ri7TNXqYThcB7xZOHZu17xo3ZyxBrtqmU2pJ7qczkOeOPw
fIjQh5jJEQ5NJE+N3127bItK+mBQkDHkD02QiGaLsGUFS1/Sr5hph0Rx+nvqS3LU
xKKTrYTFAbSq5re7NARLBBOwvLGyIp5h8kGyPeq5/+q1rH0Gm9IeuPluYtV9Xt+B
SXmhrKTF+ix5EfeQ+Qt17BL4dmzUW0VzM9F5pp52w4DdH8mXJdsc7j3oXmsSPm3i
MmFjtWD8KIvAmhjmxnYUft+ZwtKE33cZL7YLilBuFUOUEg8Zuji/tozeuUMmt8qs
F1XFQQR8KizNZCZ+l2lrmHLBgc+aZb2pmmulm+bxBzl772dPI9S0lcL1lWpHMOd3
oVdYWdiXKPVJxLvgC6mrBKfYGlvL/AjLmYAXx/dTjmVUK2LkWLaPMJPMeTH+fL7u
opDIZoCGJgw/neRFEeg+edg4af6/zZmJ6REFxfDQrraUCmvOxV9KK3EBw3qZS3Ky
7/rlaiJSJl+f8HwHHsNzt6NrV83qAIxxt4UnYmXBYSqtA/ieJV3LtQhbU+o+1d61
UWGxUyPDB7NCUoUQ+1Bp928IFfXw/P8s5eV8RHUGnfBXe/Rf6sZu4cvThAp8pqQG
6g2QM9S4fM3tpazJKlxpDAV1m5fD8tpB0mKBglVoFYNDf3G5kEGC7b9Xx8aefhk3
WS8l8znVI8VmEXFVERQsY8HGiAVUtclTCzRln+dt1kMK/baSZZLPds28fFMMBpVM
Q4Q1/jWakXq7VWbT7P0VuvCkqXlYL6yC3j10FECfJgcuhNEH6c6EQiuFu1z0HqQL
PWkHOMZfyfalE16PrnxAwyMczrWXByg9V1SYI+YAVRZ4OSsBwm9OhTv0vF8+OWZ4
zEqjW9ymig2bxbfeb7WPra5Xy8YzLjcV1UpDy8ftGgWfCiZGQBJh/jRGUhx9Ljwu
vGNCmyPzSKTDKJLeG1JRzpm5yk6BkzGfa2ASfKYM8/ts+ALesi32IikoNROud7Ot
8fUhDOqA36dz8h4/uAVhvkcqdqf1WQaDsjB6yWUNjZ+7R4icVgU43msKnBgGegkK
AWR+1EaCokNtMBCjODwaswdjDEq8WfQaeyv3cvCxsOQ8xbP5doPGz8hBtRVkWCnk
KtGp3vetDmcrVA3KE2Fw41SokixzJsFvbLLv3IDLkmsjbcRi52vnHp3XaUN8OAWl
iksmogThx1Y8cERUvOUFIA/cYvueasdRfHxaYyhF73NvpSCketcAgmyg1+jHZw+I
DQr7hpifox2j1ofX/utNyD7RTD/gLq1W37EdTjngIM1A+BLQewCoGkudP375udyy
ypZIuqhYFxfZK1BIBBrxXYR75M8bveV+N6dp3mbV9obzNEV0QtUdlJmO7u6nuwD+
huDfuhfqY3XxDpDUOqYJne6cCRNKzjzJBULWhHj1Wd3MV2/AqesL+Cy1yooyX7dM
8YNG1gqxubaH8Ndft6U+EqIvrie8vPUzd/OLKiL6ObKlMQc2PfnWYQKisvCM/zvu
GJ13fvtJ5e6QsEP0pVAgHwoDG7jxnD9SQ+JRaPBUIe5plSrh8W+RaK2K3KRuZwNA
PNccagzPBXdshs6yJDk7pOVJNfgpVl1U60EQGfALiY5yYkkB8Xa3yOcNZ1tBixYY
Duk6HDzMdUOAa9J5kAY7KCC3Gwap7c65ORkdH8e+2nk9F2Rsj+GtjzDUnnan1ni/
mGnWf1MF5wC5QdUTdL1YbkVL5q1uCy9YIkDeRWrpRClpSzid0kCVSmdSkrcrIfHu
jLmDCt11xKqUl51wm96mb3xo/Xxw1b8cAlxHfKF1sDamXpPhh9Pvf2dypoiX71Ip
JklUL38vD1NUNo8S7f6YjPMBG73WFyAcoghwL3OYeIMRc1LRbgFmxHILHpEsxa2x
uYXb7Q1TWzPzh5QkFXNRxIud9EC/dFi51vwuVrkyuswYN9iU/gqbhkxwZ7svSUcv
aXfvrM8HdqMjXmKp7HeRfMtn02WvrcftjIVEongc6d60GPNhuwG9UhxJxoEuNPW9
an/Ghw7A9opTwz5PERb4TDIHVGJzdQDOVhmhSpWaeJdf3vvNTiZ0w2sozVTeVmRy
0+JOR0FeB5XTDrxgl6qMhYV4cd0Ba/L6w5aaKj+hdkoI9Qnz7TQ4tICQyv/GttJe
ArI8H4HwFXqF9fS+nPUhd/KanXNX8Q4J/phcIYwyXDpnZ0dE/zCdoaj07JGgvHAe
C/aZX+fcjd3/6WO0LJp80LBaQhbmv0mvqth/2CC/AkW2anoQfq9/xe85xEUC9Rrb
PYIGE45U5OqMpFCNV/fhuPZU+MK20UMA3l+y9pqXllnSBLABkcLBXTA8kpqpatQy
M+dI5wED1soBLRj+2YBG00FNsbK1bC/KSKSxQHyguoD7qiJVfjrt5mmowG1V4IP5
/+PwB3U0Lj19Z4jKo750QNxK5PGJ3K4RqFrIK9r/WpugNpeofphIXIuRY6q0DkbF
Canf2aNfppBad8BVA8Vzf2FVaqZTVTPVOCJ+7M/eNVtqWE20Ch6FE3U7LkKRSvlp
bAEH8l6IMJ6dtaIGW/3zPUbpHw+jeBmjCtr15fP+plnTDnrJPOSGG1QZzqeE3A8v
W9/fLi+utvy/eVfM0cLz2rW6KTWshI/m+XZ7tKT+xFLu8A/tixTfEo4LOkPH0iUo
ivxXPurPCFAQjb0WI0iNetISBuI5k2X2TRjLjsw4F/x8R9tw9SGgUP/sLBXY96Nd
R5ZbIvFPGi7vm1tlUHTWc2jrBwiu39EE9Hfy+LhrHgcpovl4vvcJVxtllmAM6mnP
WnRtpgwyvx7/MwaEY8N5wwQSu2Tu2qjNlF6eYFC1IAt08EnDdPpmZfGIlAs0Fxbg
isnml3bXey6bdkZEjZc4dENhlJn0GsgH8omWNUIuPvoDLVAlC7ct/wwXyTxSddwr
lLnpjsxFehHpexzDFxn+h1+rqvw+epeSFJIku3O47tqU7Lc9sg4GzgxaUzAMQAKy
ReG1cnFAlEOOfoevaEOLLPtQTu1RViXT06uF1/qsSW4BObpZAi3SZU/i9pGzo/IS
MA0ZoAYn50hvaZtWYAf0h7vlT5O6wbsnJyjT82Hh27Ue5VknbUB78BP5vQymGHTa
BqDbfTbIVx/dIIJfNrMPN8gE0L+SWW1W6d7uoXQQ2DFq2skBJmMs08MSPRHlaPiM
v0uikjy66EpxExY27canWeFjPYHWfHyguwPPx6IqicYeF62htvLIxMKnIHuYPZUX
vR6dqaw288yusAdikn+Ub51NfSaDP9uUlLxAyJYlAP69oCffSFqjN8eS9m+k/Ugw
EyC28UNYBe5POU8Uhj8DOQjmhtYPv9kx9qidce77ddNm3iUlLeWZlu4Dc7OE8apd
bOUFL9LNwn4tE4zUWoatIQmySZaEMPhxQWJXKzmSPpVtxWHhRX1e0iE1mvTM1ndL
JGXn+BICrx/cNtx99Qn6KaAPmln/zUTYFPJMVvnUdVTlyM4dib9C2MRInMIuEod0
E6P+oNOZLakuuTH2xDohD8o15wYLOxmxi4OIOc5iyLIC+lAfTc1uxqYL/VZw7Xty
twmS/HYiQr/vSc7XRak57qT7jeTer5fZGFCsnL/7PGGh6OoVrfijJq6n7UnfRipa
iXtiI4lLvKFxEw5f0B/Y2EqCjRIQU+C58ApRAQvCGpowoJmEr5KHx6/RWrXeIvhU
0sScztteVMonqwSB7EPIbarTJ8Aw66ar4Eic6wANM24uypTv9a7h4jjxU2NUQnEZ
jp92OySnSj8OuGHAa7gySlQnVXmpcNohPU03wBf8A7R3ydSnGlf2Xjgzjv9RYLO5
PszipKSkBKf+s8OPxp3VZzaUpdLjbQz5HDj3kr+tnJy3nyK9O6XbRb+OLDE8bhy/
ByGp/+46xaGpGU5WMuDBIAK+lhrkz5Q6GmJZ2p/AvjR3D25k85oapuW4mr6I2JEv
wVzVPlK64fjCrAprCAg6/fZ8N7tntD/F4s/b0dpe91bd4WhZAA4oNpUAntX1SmVe
/IOiAyNFOXb+HvPxf5Oq9sl8NNe001IjNYtI5JNFjY6/o3MfV/mzLLTKkS8cdoP4
N2Gpjhrcfogwom846i3agDeFMNuFbiQSvqduFBLl4ZnC7G149bczeZmVFU0OoDSm
ExYuTO6ceKQDrZtqZhk4jEC2lp7tMVpPMppYxHyHQbF/VxnOhnKYjlVc1orJtcLX
epDm+o7UMqV3VzizOCIn5uzZcsyM1tWCl3KMy6CtzLP5nSaMXceQCnz/4tC729VH
C4EaVmWEHtXaaZqxdXeRrCRLz/OLVS/PuNKKM7JKNopmNweQtb0j2JJL09LYdsq0
u8+YvJcPYdFOt+M8gttHZS3kNB9Csx4PPfvUl/9O3Lfvuy8b/rKsVB4mzEBROKhb
0oSXdL+v4ogdm2fiOwLDhToiLIInXwBOMvNBGWTGcmwPcqfjUDybDBSwBKjHqavr
fxDkyA0kv8IQyglm/4QQxbjSoEvZK1I+0uwSRpe2PCYaWW1OW9FcBqUfcoxBAxf3
SbBb7O8k00t6VrdeFABC+l0O0sqy/JhsSlXQzUbWzP5YEZ+xo6WQs1vatakpXkN/
PkKXnf2cP8C7bFhBQACs7Nwnh0BcDYisy6KAwDBeedYlnACkHiZYB91thVg5QsSR
Qz0Fwrn78iotIeo9flwFnPaYWJ7t3fWvmq88EIp3iDpd0vsEdAeHrIArOQDZdeS0
U/Hctuhhy7XreHgEMpHqZGhuwmZmH1xFfSn3PsOwL2+DjtWE2uCm7kfKli4E6X/R
g27KHVqcC8y/dgAmuoYyUO002L9p98x4/xx7ZnTwto2YuM5Bh0faMFCMZYA0IMhG
VTHJMq+jVyq19+9EzSZWmkSYuKwMLO7P2ipXfIaLSJwtp5p8JjobGdVjzumEiGoQ
fHF75mWUHKE4VhBhcjVueKqGC4c7hidv3LQFAqMQjk5aXpVgspfykz+lxgs9SiEv
bWW01GhMhxPpguULk/438Kq4JUH3d2oQkRPZvQ+BySEzX9Vfxi6nGNRo4YnhGW1O
lv9zC4jideHZ5kRd4yij30pgHwcfORH9rKK7fEFaZx47+gMq9G1JJqBHQuU7itJR
Gl5bQmgHhq4B7arBrqKUNmCOGwyC3pDc+IUuqKfMmjI12XqW/xX+bMgTpM9lNTMa
/lMoNDV3jXKB7ac4eo1XEez7MtqYKXFnwLt7p/i1zt/Yv9tiXXLo96xhXZhi3WeQ
DI4Oz/vCqUgzUx0MptWf+FgU6xOBajcSr5RrMKxlgfvxE+/aTGCLD2LMFNZr/Z3l
VVM8Cs3/lGndyQqgWMv0JHzPijVJoQgJ8qeIRtWzEuMHxdoaolYIAt7kLvaVJKu0
U2GIjAXqC8q4NRPxbaYI3EclwHEe4VL17HSiwVjyY4ndWGr2+HJ1qeQIDXvfSUui
OxV7+38AQOpH/LJNBpiDkY3i/PBnDM3LtaBvPThLWQ95MwF/A9KtPP/5O2pbEB9l
FEh1Fy21a66xKh2/dDJ397uWwmrdbvcBqe6QsvJ/zxUD3DIYTrfdSPfHPOiuIElv
UDZ2E3EbMgC8XiuYnlafxtJ4UKhtmcArs8VZSmWAxo39xBoSKiF2ym3KiQeBCIcH
eP0VEQnVUrTh4Bl6hMcykGYvovUJHufMAQMavTRRN97nxk++9UCTE0EUA5/4FMVc
alRXZOytOFbp9hYHhJxWlYTnDORbpnZZOVohBkfmInYnwwcxUtNtkFvBxcENOjgN
+ttFw4ilR+pBZPS/5rE5nvZluTdQ49xzbQhDyYwUrtXefeFIYmf2rlMYSN5SyQbd
oZmOenxZ7n0At+BBlBu4bbn3FQ6Wl9xMkMXEZrqoxVnj8yDSxc8cEA9s/n2gMhY1
crILkteymA5vpbxQIQ0BctyNmNtG2Bvtp/8HET603x5J98lAmnz9pCEeq3wdkWh7
y2UoFE2h3mlJddwtKj81OxoQ/BqVHI+8p9CNeH3MqxO3rdRIaH9+ynDyrIHemb/1
FiSyRDsuB+/OkiCNgeNRTm7QodZD0+bY7ElIineS6QyoiNx769WRPODZ2qJexM2z
YZ6rq2fMkCM/9KtTOoKhdjhP8JZHT2FPBzgcPAHcEpWuvsFrvL56gnUme124ua++
plRGo1k+EGmx7MhMoiqtsgR7+PayD9zJEMYFLXmNvmAqWetyBepYV8l6RDrS5FtX
hCGIXMPdvpLf0uE0qlWYvJRrxgZbMlohamLSiMUv4pS/m89gUPP/lcP8/vXP2Ddv
ScuUC3M07FG67SAGchZ9yOVH3XVagMBXDJTOLN8dmGyjIV4+U3ll/vGAZAX6dS9i
q10jRrvvRS+WUSqAW0VITE6r9ckdwYnRDQvqWqWFv0arU0TmDaduexPPyEi1dMUP
9sYXTkQmkv00LJnAm77Ecf2aWWROvcde8ZUzt3m0Fkixv7sRARs5Cw3vb4tI7ZdA
uSLKPUHKWYWnluk/4TKiPJLSZ7q0PQ6MtaCwgPfmwaHT6yrAixReiH+iPeZI0/8m
LuCUrdAR4+StkskHIkhK4xeDszDoWT+oab8KFhI7sD49kOdYeDjDFRwT0GtIApVc
CXF/IYHYwwXu4eTqa/P9EMKJ0n7u4dOxO2g5Clpt2EBb3x2Zy9yuspayM8kKF4XJ
tTtV/anvq4XH4uyZNFGsgIDG1tvgr9daC6oik/waJ4z4i/kJE42tS9s8X3FLFczi
iV865f58IpRzWa+UCnDilqXVPw/97ItbU/K5X3UJdNp7IZKqypHUAkvptHMt5lmq
oOKk0VRr5kKzEcbRjdjfQ5pdXBBDW+zyEIDGbCkJkbVAWO4zy6XvgViuFqHXxBSz
SKNRHMzzenLLRPXUZI9QpwaXNt56jetpirk60kPYuDnhvxbqD5ab02lbHCTHrPSH
TFAXS/7aGnp8DZbCxVhAWiZub5FUcK5jNFTnltY76NGoHN/dg9v7S5652A3FT0DM
WEBcDltjWC0L97U1zSCZZmQfDvTFxXon1EMrmiOdgM3t6EyeU/EOi74LC95ejbaX
bziZZDEeQ++NiGOUP4HyyXU+Wr7o52H15mu8XcEIfNoxnXKkIr9dktBaD0HruQvm
8f+v6kQMLQROF8nO2hx5xABLGu4esQI/+R0ecBLU0WqVqG6kQaRNUX3XSdjTf2mm
+5+sBselxq6VJxrt1zts4SDvvZNYsDJtZzozuNa2bqSZRIrIEMxyYB0tsDCYpG+2
by7JpK2R/oCt0omg69TE8wM3TCSgYY3sgw2vzNxZPJzA617sIVxfFeqaWczn/+WW
+XkHLdK0fx5IHPyaBUAvXD9PjQrxcSBd8fjJXtL4MRVTR1Oyec4tq7WvZdVjsncG
4T4cjCI0wC98i4VCG+6KLvFh+HeYHyQ2Aip0UpDPQYv9b/+KUk5U45St3Z1N6Xgm
mXpiU97yoNx36qIRRE0QH2fk2y/NSv0D+SwfVDc9CGhcxr5+P2IZiXujo/fjmkPc
9huvwZ/PCs5ebuXpiRen0qOtRqyamiiiDmExMwky/e+pB1wUg7Rg9ispejEBQtaH
edfjnv8IRE1Y/+0x2Chmydy+GPiQBO1TuHr8htswXdKkhZcRnfe8ZXwP9tZeYqdu
CgRYHwpa3uYGKKsCwiX0IL8wbBIDC/9au8u71gTSmZBVrjHylbhvW0q/UVDPYjFI
pARjDHeVlD8Q0GYqQ12V/aN0LZELGKjYOUpoFB7c5WTNDTQ9RUqBVMo9UE5cmEgE
i3QuuaUN1Oul6WGcPP3IaFeac20pbB7D2jZufBOHh2ojwnCDgcq2K7L48K2+JFrN
rYrd6ZKPfvR0fKWxHu8KLwldUQJ8x9PP9IRo48z9GjUOsv4fH+S33NL36/sHvqDC
H20VFd3C/w5dekvGfsyLsiWOT3br2CCL5LCb3mNBsTZFcagqGCGqLYlcqVkn7c2g
4EM8oOVgFP8vbroBgy8qrWLGcoppCyxa5Y2HawsYtYGlFmc/0p9poN/+JoHtke19
hBMyEhmhFIAF9sZTDFzhrrS0SUYn7RwjLSxs7sZ3UfyCu1Gj0dfrE1knZDnXxVAP
yhiTWtaFJ9BkT9oKic3ZUaAMSaLk0CrebK+7u0wMKoSxCENcL0I1E9j/EjEmtU5t
x3aqfbtkyqhWlumbvk6Q6ctDwKzcSEF4SY9Wh72/r/NKTfAwoSkiWM68t7H0U7r3
So2vCswjBl7pmrpacNvkSs6Z9glFg88oIetSPDOxb4iiWmvD7tUkPubOgNXMQsOM
rs2XTbWcRMPd2/rlNMZqBfjvDanctxr4Df8wKfIbsq+BGuDHh8cvGvZzyU6uUe1l
Z/PCz2YM2jr97jkJrvNaF1hTZa81nUxQlnI2n7QtcPj+WYAESDSwj1jmPKUzEDyH
sLqVzh2iHSu/SWGHV1wEthM2j1A6xiBpu3ED0FVv5KARw4Ercrdwdk84lTLGP9+I
7q7ck3IEJj/XX5dTIp2urLd6zfpHV+42ukcwFVh2unIRZhF6uJnYT+eDOjVPANeL
cpdkdryKgu4Ri5u+QuPUau8xaGZta14pKn+8KAmRrPo9znrhHEuXb/37CisEMyIr
QH7IQwAizeBWr5i/gH/PY9+uDGTBrNgk7b1IU/MjTaM+65CD7i6LJKNEq/sSwllv
LTx3k7LNtbxbrwld7Iv5Dh94yvVCmZkwYaxQumI+bbkXh3q8W8HFI4UswAbLpfGU
egpAxAsrrNupde9KfTFZGc4jJJZc5ophTNX4ZeYuI2DoXytrRSF7kVwmcolOm32y
TfXG0TLIzcW4ypcfJo38WPaNlgIfcLADDwHsB3PcJ8cUuiIHLylA3EVfeEpLYMwM
chaOJdaJ8bXw8JmI9OpF9Yz3LNajzOjbD3/qIHcl5nsTi43u2aCuiq2/kDK9I5Z0
cSiOjyI56qzOByf4ca4HGQUMgnWLVw4HivSb6sf2X+EG3WNw5QLRDAFhJXiLx92D
UvguXWFtZQo6JXeh+UsHHAeH5PNAHHSMnQC98lanRcPppacdzngUGPlAKmqWvpIR
+rRduqsshR6bOEGEYS7FhmZ/UWUiTHBas8JxhmURglQV/N9QUwYfF3Q9YQYHRCfa
zka8T266h5cW3fA1jSBPM/jgFJVhX5SV6lTlCjq7Z/YfWA2sTLQg1smNahK556Pb
YHjrIKNxQAsp3jN0JdHtgMf0VcmMbFojzdpwXdxurMlqnm5uOVxp8TQx1+dr+5GI
0/ujCpUqX48W1zwilNWhbnXKdf9j+nydTdIIssBfhEaLOTJi2nY/M0O3DiM2x1Da
M6WrfNeZUXCKiOx/p0n+YMj8q/AcZoKmmoyETZonTyBaHbdjaHyfBNWlPtcyPkJC
pQkLMetbfPmWqXY6o1uDwhqR5BehuRLy+D/X9neVaEZLpOuEBAPhfqSeZIcxUZQd
FeG03nwYmv39sPOVqKDzQAdLU8cKufob4xx8DNaZRo6PY+GGRuAeuKBR1s+HDAUr
ATZlzqDTOw3xN6892XeCj5VJ7VhUs7pifV4vzkil8b18oJgKDfWouKwlcyxQk1jn
1F5vGZIJIeQ38G/4Ywh23N6w6s3WFdLnS22nGvqHYTeVfxt0daALhLtBm7W2qYND
nKjACQcAug+WcTD/S+W3Dji/xJ2nv8W/ei3a/zp+jzG2T6yORRYLn18LJsIgc0+L
h3w1t57fdizRYfSu6r/DaD07Y0SsALWjg8z/F8DdPiI8U1YQsCn11qPGm4VsFQjk
Yr3nbqKE/UUHHUmKOj34Cr86Ls9fINPr11Iou9rm6YGqNH1p5jp2Ik7V7ft85yrU
Av9Ixacpp6M3L7d2cRvUj986IIf9dmyuusJ2jaKW7x7oGW4dXvvYFk74wB9OxaYn
wC4xyO3eqeUfd9xrHsLCVIWAVgJQIz7eniAoE+4e0B0LKJloRXjX5ypl7iGY/NLf
UnP7HcaJ5wr79w9Zy1FarTEJEdywCfU/e4ZGvKxCyi/3FfFfzkGZNFoanUGVpJk+
bPqgkeJTJyQgLweYKTu9SPO6qvBeg+z3gSjLpVXNZReHbpKO4Kch7SAKJYb7guYx
Rxw2iMU1Iq0BbKjqTNfobAk6XN4WNHyiXGwgfQaI7ofhwDdLo3bNnjaqET9elZ0a
wrlTbB5wSpQcNw9LxK+pAfJQG9U7VQguoLYbc3Hu1WJyutuRyzZzOTqASzJSz1Wq
RBHTAOQxZJC2iExWFhW2zmyp4+FBPJjMnuNBDGX12ihoKiv5UZZW784QRztS+Avh
VbJ8sxEX477HqVqOuJgRExrxrHiPRMBxUgfSjqenBEtr5AovRfIJZl+6e2BvSGdB
XZUQb5MwRzuCbQQ9DOtGyDIiSnZIyNoBDXRTGFL3YPQ0KUXh79qGe9fgsLtUYhFA
DDNyXM2NQTp0k7iJWBuT+ngcefQYApV7iAvMSQHJElQ5v6XXRA6OQBTsVrYncwVK
54dZZT9G3fIVAquOOcz8gLUkZ0jIRS97zGdQVkX39FwGVRyXSgLR42BhuM7gAxR8
Swuff89IcCR6evKnIEkEnYLylrGiyo/C+D+OniStbYpZAxaEoTzx9gYqEHSb5ozQ
nTKcWg1KctMYdi7tWP7WyBvKBG4fG7RzREsXbPwXHJoSXsNg6GgywCgyoklidhbW
Og9Ozaq1+fj6QkFHSju51IZYS/dx6aLpIkpo5Zy0zOyk6WyStrX/NNH9NKgPR3tw
Q8s4wOWtEztlM1OKGq5aiNJlSc+WQlp3htzdwTXN0mfprcR85cU7GmwzoGypX4EN
HZ0+L5XB20eeOysWrDAT0Rb+GVHQ52c0OVc6EaZO1PgLGG8bO5MUII1ZyQTZx4AW
zbcpeQz3ZaQRl/ZmvtgPwMDEcfLT8yY6MDVn/3DLT1XWZI14A4u8p1Wlrxd56c1U
wb3BCJIt/4PW1z4UvSLPYoIy/itiHguxmoL5R5gJe+ABgEva88DT5sY9CeVJfQsQ
qDEpWPdvexgEhJkp55svIuIUmUlFtNKvxZSSHbAfuAiVGapM3fP5shsm5yEHXqG1
5CyXFvZnGROzC63f/WUu6vTxt1X8/ewCoKayaSlLXXN0GcBwa3nkBY9WHROL++zR
X1ihkKQzsoZcwe5X+4pXfrfv34+M6IsmbmQD/FjchzSnB9NBRZ815/e0YwsxjOKA
xAkf663thZol+9dQnxvnniFF00Y/z/JfrYgb9LNHN2Lyv/Hs/PgXakHI5YZujvcA
oDjpzk+4Y7dmH0XEfD6nytpElZsyFzKakhONtWFnIdpuYdjHikndV5Id8Fk+QttC
ReFpyUfORpHDA2Dl7o0FBQGOFe8/30MrznVAn559KxlLuNAi4/0YtB6pnWa7aaxs
gO9QDbMZ0HUZIf9XLwjxAz4cy1gViE32c6n31PxERrgcaT0zZMCOVY9oqAewalQC
jJrTjen2irQRL4B+5wWUIm8A47AyvpGcAKH7YKO0fZJVBLNOc+4VMNhnM4NRI3aL
g8XiuIa+ClhEboaDruTqVjORykydv8hHD4ivIa/OU5d8udenIQ5awkzCOLI2Ruff
n3nHCnoEvIzJQBcfuxjF3PZyFuN+tbJFTw3KZ//I2fEYA17xj02xQi1YJm6oVlri
zQid05CNeFWTdZXoqctQy0tw43rlEUTgAvvolucfDByk2dtuNRU03pRkSUs4tld8
AtHNf4nt8kURlmclH3BE2iSUm2UEZpN6V5k4g3QLdUXjicBkfy48Abw4mbxjdRb7
5oqrKJSFq7MEJGwoIp5G5t72+p1PZdc3L0omUXe5q0RI9FlaBe8oOW7tV2ypS2Yp
5lKH+KSrg5QrebHtqT5gssL7XgKsvCb9LptuINqMh7/heSj+vdMowbQJ3k6l1b5y
eSiUItoh90A/2YNtPlkA+5afcXuaElOdraD44nbsi/xy+JJrCS6cojvkkUEhabQH
HqoQYyTV4tCRgxyY6lRg9kz6Us5JtJx0eEW9Vm1TewmH8GD2aOyHA5smP05dl3Y6
A/arpF9zIqaQK25+CGLBOmf1BtOSpvaEq5L3FbKvc945Zt34i12HrP7PgPUIPHmW
5y8Mdq71HtG9LGlFs8X5b/811ffGR05S/LeIFiObeNMRippXvs9n4Kqn7iUwB7/a
FWgifozoHb6w4kZCeQ6h9PeWaFhGTKbLU+cxDnKP+YFKU+JRo0OzUkOtPjNCWisl
ui2+tDyu/ZjSayFzSdmFstI4JTE5xmtKPVv213Xk24abBCNRnbPU+rYdi96Uekbn
p26PUPTMl2j/4dr0Q4A0k9cgc4YusyZVVC5RiF7IjiNWDpO+lHEeQaboUxr0cRlj
6c3YZ0xo/mCQbTmvHPEq73LeaAhzj2jwemxyuyy8x0nJXbVYJ+CQi9EeN/JEP2fA
M1lcEPo5zHhLqp79FRiF4WQreaPd9tOK/pTL7aRp202a+Y9EoVUhXe8sEceuLhh7
Z6ex/YmNyMkCF003WDMoKEBEWLXzOTSBbdxA2lbCU5mUpeOmAflMTVrIx6czkQym
gbDBUEWTPZ6ntOwBRC970dEjZVAhyAgX3yVuK1ETk2WVU0MXXayBn2L5gw/5o+Hq
H//PhOdVVkjJ30Raz/TVr6T3AkOpC+o4RLe53jWaoUh0V1kqdPVCYh68npQQ2cl3
FT+Uh5ZpeIF+McE+k7gyiv0amH5DaRwWR8aHeaMLFLHjILDPMNMGIZxTdX65BJId
aFyXWHRvipB9brXxzlMPUeE1gNp2hCEoPPv840uyIW53Ilj9WlxKXS4BZEzb4r76
hth0s5wy/2YJDul3EYoYq+ggNhMLfeOmfobksPMZmTV95FgISKqmqFdAjZ3utqO+
hBIoY7FtSKjuyB6L2vWRAcvXSBXKxbQIiXHSSlFdWWJFH/Bqh8bQCHf4PYBpv2Bo
1Er7cuRMMoEfNgXpdR7r2aHrl/Z4WKlVbFOTmUlL+S3rU3ya19V6pjoYe+YIUj97
9DxeVaVCuh/og9Su3REdi+W772Uh3e2hUTUAne4Bjnc9H+i03tOsUn30OpCfHQYU
qHr21sIeYqsuM8cXV5D+pTjvXR/c1g5HsNcRredd+EJg7B01ti6xeHptScxf009t
Jmg240KDfeFXC4WzqV1al7o4K7kcZXL/M5lchoNUF7PxdFoqt6tqUpsc2FpwhM33
81f76PLPQSpY2Xi5O5G2Unl5dWqaeWd8aHY7pdB66dgI8JzPxhQvkYhGm2FPPS+X
MdVtf7pRIy8G+0ORXDW+j0+d10iSwO7dRrPQkVRdFkPTIkEIgmL4amTrZ2nzZlq6
8So3PMR51KKlGWw+ce4Bchharbiwqt59xOGZ2HlcsrhBQjIQYY17eayMd+QAdMum
hm4rM+rXBbiiglOIX44wIqShRXIKlgs0v5nywvHVwn3Ja7eTy0kVBxwBstNpBO6D
yF9aHi/XbkTRRQ0E6bKJsVxY0UcMWnijlwmLkAHa5Iqdxqro+CEuDXxXcS2lDafm
J89P2n1ZcQ9l7olqzbmx5Tim5aRpO1RQVOKbb6eITxMoPso+jYa1XgFOWXMf7O9F
rnD13FnbY0EZuZpwj+VTyEUJ/IooNWrOT4BuysGG4PL59nVqmgYyC9IXS6pkXbrX
om7Yr2Wdn3cxm+hrP+PUfxIH2LhL2EYLllkI3wkGXeUez/r8ZBTruCySsDorJYZS
wBMtt9qby/m7YilK+OI2j3eI1OBK/4qjdFoO6PjsksAuHnSofBSAoRR7Yki0WgqW
tRUx17JAZ6kJ+kZgELkUiIS5hF1DepepNBOZM4flqn2tvwLnSQrItEK8CcOxz2d3
eBaIyjqkyVzlOhZ6Gn5dxJvIW864+VyGfyEBMG6MnU9xsQhr0R8roPeCEgc+COy5
NDr4SbvDnRXY6mTrdRPt4dQbR874stArfIXWQ4EUEkeesBi+nGCWxtZidbGRz5Eg
c1qLu4XQs7pW9f3xT1q1qS7c+nnEXjvnooDNsE0SkPqnpaLVifmngUOfRaA+gwp0
refh1/LgR8XCi9eQxHssfuUdMaBEv820UcesBVzUNCc8n3vwTKo1ejZEqpzRCqbM
QJGObXz/fGEOctrHHN7apwGJ1iGb1NNhvE5Sure3GwXWnL6/Vwk4Dtv+M6QIDW8D
ygtAJ3HsdrTZPRnaj1A7IPCYphwdrWfBb53KAP0sXtz7VThCFPDZmGWc2VUgSAnT
ouVscXoa3P9vlHKRt8bn/40OqKJOR29YnKmHz0Il+okO83Nn7S0WYKc55YmIq2wl
UITGy098M+WJwnMrbKTCGYXee9o/0Xm2mvBC5NzjDi36UYsFuwAKopwInas9Yw3j
mm2H5HCySLDIV23cLF+64mXJPhdsisWa+5EnpZfYGKG+sOUN19Gz3tkO1/uNwHK4
oym8zpa7YVUPWkBD/MH1zFA3iSrFa0S+hnRy4sG+TA/fxg2iyYr3XPHM7XszJRwv
WVJsWM5lHp1NypfYa5Fs1hfvp33UuyVSPAfdMzIhrV9jL1V9Ld/f0c0wKlg8gYMS
9HvsysBxlPcaEk7FGECKA9wA61Et8oCIlf/BBC0VxVopG2+1IsiLX/lYAUdHYzlm
q12Uem8tFqXAjEuqpqTXkOLMD2F+bjhS+dFmL1lbUV2xLaJfdETkKOz8CkozCdNc
ovoSfUCRYK/vHS0Wj0/A/0NofVhazocHPxELhgjdBMeMWSnpm0gxeIZ+Fmwpz9Vp
BtsFZ0kX2uT5/ANkkeLfvuUXoeoQBmckHmyfSoJpHH/5i5E5nwrLQ/eqJn4Q3Chq
X0NOd4vK9HPkupIvAigym+TJ/eZSw09kKgo7y+BQ4xbZgSqJ6uAr8UzRGdZa5BRc
4HYn2rIN91ISmBiEGPfBryrXjPvwvwwbwxJovgUe4nzjY7HtAQhPzLmDWKMYhIvj
f3GyJ7b/Zn9cAXp7m+l3C+30jfPDSbZegKMD19z1tqMRraG1XSXXk14qPs6nW19e
h40L74DX0PsQGOE+THRwFhCOGD5+zk8G9EZuS6Ps4PZKtMxtRDHLExq5ncYPWY+o
a6zW7nqcZO972vREfCyDhVmkF6x8Ob3GqUogKOVwLRFIfqOoxtgEVtzy1ZMZpIbI
evvj32Uk8fboAoGX+rmjDabn9zTrYw01dMsfHkTA++V+2MWlcOMnoTZQ/Ma2rP/m
8Y5fVvnEuTqPxChjbn29ZWdGJGmQsN3d36X/NJvL3hTu4xdoGDufLS+v51Tf9l0N
ceEU8Koc8erv92jRaByH30CgPoGFiu5/PSL7bMQ3g7Dz04RhNE5cPbGExG3Us8Gw
aRUwG0rPRHuJj/jMLw1dacdap1u3W6+iXJZi50cCEqGQYHOj9YVXS8ivZlTcYAN5
o/sgGAfLs42+U5O/nKfADenwkm/mK27mP3ZiQm5EVQwrdvOLKKid594CZ0Cu9PQe
nUXlt3XYM7BgS7XgWnDhyrqlPZdbUg9dQpZIT5ZF5nsr/Z4Q7r0qzkBBUYUiM2hA
eerXkBdX9mhIW8AMk9bS/hOpIsTNB5xVuQVnklQ2HdbgjQJZrNds/xFi4I2p7uQH
jaZv6wzu0454gANAd8DV14Q56fjisYkvHBCf/b0f6ZuMe8J5cYyCErLbwirRqYUH
2KcQaL7g6k0z6GRJLQR4ooiMt6wnip4+8FpxW7o8N9PnJPQ/3rvjdahlq3rLzNlr
QS6bfJVuBrOCddPhsttMI/NzJ0Rb3hBkrLF588PJa0vjGz8R37QIcIOoLA4b8MJL
775mpCFECHoXG8z08XksX3I6AG9zcB84qD/Z7+7a2wnpgEJ27twF2zlX6r7EQN75
ZlUZea/BKmxP0BEsPGzQ/3JBYzIwmuTg3sC1Fh1WK847QBJjGslg3FWKhvvYecGB
yOUO4dRoaEoMnt3/4FxMrm+ESuU+q5pKe34M6w+FJ42cxSMGwOmsA7UnSX4hToix
PyqyvfwIPNXsji/mLUEITzOgyCepk2ZLkAuX7zYjSO4Wu5Tra51ZBkMBE9IDHj+G
mvenkLTAE3mRnPX5rFKftB4FZtqIcF9gW/V7p38zK+bxcf10RiJMu/ufveYRbrRF
Oftv/QKrbOtEkhOX8tCgMsusU6hr7zHGq4DwnACjrJuwRsvzZqP2YNtxvf21rA/6
V8kTKKXctSUMXg2202Bi3XaBeuPDrFMjWzpHUoaSUkOC+jGon1snafYQQz0pPQGk
Zk2dquYkrlHCfJw5HRFYzgdrfpc3M3YKhRKOZ6Jn1kk/ZCvPgNlRzCb9Kd1E8g2R
7AJT7JgUKIKWZjqlibJ1rMQRCwMmQtP7hp3VDYk7ctKHCBuKlAs3LHQg5SCCSssf
+3sRgNDs0P64Jz9D4+7DwRmbYt37v6cXEvoO2iwATgysC9VGwdra0oCDCfOv5eX5
Vn9YQ9zVAFFNvH6LQArwK3XHYq/s31LttOW0p2YDU+rMjwllnJxJgBQJ9U9tZkDI
YvI6bnQ6pnCd78bwVCP48ZImuWq4Q0Bl5QYYdKFqtrRf9xAuzmSRh7dPODxB46fP
oWGi48K9b94dPJIms7cSNJLZBWaN8Th0sKpO4s/R0490UghYr9lPiurAItoQ+p09
ciVGPgLHB5xanPkHqk7npXOU3P3bExgghfGZYsDn1zCFYq+OvZDmCTJmnQGM+kBS
DYgXCfGrGyjVR2yFw0szUJ3tfxX8FAi2VvMSUtFNPVrBQdqdqLBLxr9EVUVspLdI
VG1pURNxXQerPFDvloqHqUu2lmUYdSuNHt1RjQ5hmPLIjP3o8zJFnQraqTpXM2Gy
KRfGEEHQP+PrRgREWjIS2gRbLMk1xh6LIl8ordp64AYcTdaTnHnQGB9jwanwhWKn
TirQrAzIOSVNbqbtL26EuvJYlVl9flVjY8QlH666n52b3JKYTC5nDsvnquhXK3Vc
yy43pGnqnZs8XWEmkZGhaKHggqIdfiF9ar6auqhqCZUehCWSZSkbtyTMOVLaYJIH
wHb2/eimUzaRdfTVrM/TJg1QQ+mRX61ZL4mmxOBzHQ/p1yUrt3uhvdzWt8XBktbH
nnogPTjzgYFjmXsoawahbzjwVBLItxEQsN9llNyLHKqjYyLhM9gsUTaFVYGhaUS0
lIML045Ay7Bam4nUmZ4KHb7AKo3Mca17TZ0mgkjZM5MLB+tJqY+9oya4F9DCMyvI
361mhW27xkG/UvctY9uwwuBZp/U+lGaBMTFemP3enIROPQlfRezprfPEBtxM3oh6
YOy3fdOk/Y6fpDYiJ6HFErcikDbyVIVZwo5mduc1+i/EdOylc/bQt4fq4CU4z5uE
1Z8Ac27cAlAHl0KCPuq0v/+SGd3zL2bp+JcqnOuTjBJ28353jH26HRJKHaZXcacn
q5Y3n3/ifn/zxtfZ7uwsCDbF0ObKw8iZrUTnHoZsnfNsF4ptSOXMXWrg08NlHy17
HfaPx1gsyknPniyIkC1C5cY6561w6+wuCJm0p7ekZwqPkoDOue9BwtN8M+v1Q2db
bJ88QBrWnTuByPfoxjAAhplzhXsH8SX8x0058bihGEve+QOUS02u+rxyLv5L/ZjV
I+vOTIN89K6my228e+5LGv7IN/OmPH2wZPfCuXjbYgDfggJF4T9mTla6hLgg2UcI
ZC3J4mG0rvHetwhUi6set3Nfw8+xGhXRyjELskmmhjkH9G4E8CoHDgsxOco7w7uG
9L/eiLpowMuWulLwbcvxEhbFzrSpe1MRy9p92QOZ8hDr73pjxM9nGmHrPRLXSABS
G2vi8xUNcqG4lzl5j5byGX69HYEwBZpGAudlxAEWBltjYLdvxaSxnmDuMEXJT3Sf
gUvM10L2/lCqthTNARpjeE+Q2iOvOdzZN5A6aXnTdq2PHOvYopUawlMkAwIW+UUH
fL5Ng3NDIEEEDccKh7HrtKIuDD4TlIJsEQDY55xIJsT3FPh5cUU80xsjkkIW5EtB
4BEhqAa2ckiDR79uuvFNtQONO6+aYVt5GWGXzQB43V2o0FcQykZf7O6Z+CPmczhs
aemu7pV5YHqrRtvMR4jNCiFGETzseFo0tB5rPoDl1EWqlMS3fuPzTLXXUKsSd/ql
wKRb56zW0uCFQ9nmmkCurw35VBja4d7RUa8kVrrPKo48CllUANvOXekhduTfVDUo
yJnziFQpi1Xda/gIXgD/VRYOUsxBKt0zmYsIRaw1VCx9JwuiLahHwEm9ZZjYzj54
GKxvyDG2qkWqJJnWopewUIaXk3CaegRpKB1FtQDvd/YhIXYoG3Cmzl7SvfiA6M1L
rD2zkQtOEVXBqQknyoqY5O/6feBUHhU0ECKrrGKt7BRHuUc+Nv1p//bkTc1rpEFU
It7RRPjvE4sPZ15ud3OB4dOVh93yKlcrwd5/v4OKKgaGhRjYUTguEPcKpX+ct/O4
QoR0LzvTJWLVhtSOvHxgu9ok2/uZUatkoOPDAU/B9ymj5daUTMab2Dg6CDAI8mMW
zqkwd0bpR7/0M7REzmAmU+xqOKAfIOTb6kQ3ihotPdfUwy6iq2oZ+Bpcm+6YV7UP
LBiCSKs2cJPCaEwqI7EHRe1zbhoMGBLnegBGoGfYw7/272232Rxf4ybZ0K9O09l7
LzIV3psGSiro92423Ms5j8Y/7qBfyV8bc17B9ddocIviCaOHIaq862MWVB3szUyJ
VrjlGStM2jsMMximzTobQ/+HxY7qtaZAxDCC1ld5g9bsCbCB1WTYohEpSj4onnQ7
U8Aw+PKLw+vvJFFJnhe6KN1v8s2HXRgMZXRaOQKJLiVo6rxjLLfT0PeMCMSuzYdd
F1rV5IyGE8gqiydy3tywDz7Hg4OjbSBnC3gTgn2FKVLTYTX8szCKkli9v1llMnHX
7W4x4Y2/gRLMurave6U2DWx6F6vhUYdTmtyahoAVZVHa3WUvu6oCFA5rKRHi7Cog
OYuHgGutVDAZB5JlMRAkedSFqm0z7EZC6t7H/gsFJsmFdGE9pOcBIB5AMQPaTyD/
HfA353xb5PWqJqbJtAsMyXrQqLp7YeOQZmJoNOwhcT0DKM/VJ/5GJsFpwm+YkaBC
1jwjk3FS2I3yXjvgaTuljRA7mgxOLSuROgDz1H/ovltnPUr9rfdxeLUvACFNKbiu
KsqdewP6g3AKYhRVznAMd3bPx9Tsbl8Kzye7PP5Va0a6m9yx8RoWYLFafz051kaG
hhM5akAxw52BIheNwTAFUPPrvJckYZwdYcAWPWxJECGdQpTwhlocR4oKtW9oJLYo
RhAZBg9t0LjcJt7oV6tz6xaB0qlKnaWK5AeCphtaq3PsgySacN08TOZP2hiOEWxi
xsC2bamDXq30VjRboQ/EXpXoJ4duxo9LpyCdYzqCCwV8D/vvmfez/cKrHWIfdHE3
XLleyH//d1ti1ohe0yaN4gi+Qmc8yurSnAJwp0mjpjeX9DN6d540iuAFbXIMvFFu
xkDY9fQW5p3GLwJsj1G3Wr9yFv39dZbl7w6f3gPgWxmKzea2IDG5dWwXyzbbrNNM
Vhg4iqBRljQOtNCOUQwhhKZ0ArPb60ISKSEQA2yha/BGiRWvZO16XJAhtzo16zSY
gI7xNjHDgxExUFZuNbKzaaotHDG+i2gVmVo117MzLAQtQKs37sxQuN7xjfPrF0pJ
yInnuVsrxDbWSFyrubPB35YKEpX/KaUgLweFG2ePBQwsiQ4lc8GoJ9JKNeRvqYQN
mFdGJACnyv+s/vIgSkweQEL5Ug2aSb4mVE7j7F22iMe5DbRsUqAfFi7bUMz1XKZm
aEJ6qdZYNDqSZUu8B++hESTtn9NKx6OfnCQl+V9pGSYDA9AkNBBk3ul/k4j8k+8L
7o1feQTqT3r7gVD9/2i2vCyFL9NIWd6VM+n1HZtt+OmP+YzFkseSEQLS4by10VgB
Gm/+YT8ixgWuCndv7OmlbcuA5S15m/4eDnb405ksKay9vumF6+Oph+5Omckt8o85
mlvEnXkSTIj3wR56bf2uTxv/VDKRB+1Q0Ac7RHxiPo439krhzk1hE6cCNFFjcmOV
8ZxIedCGuaRQVpLu0CktMfm+qGNcNDUk6h8ovB+I0QltL40iic4JlrFHxm4bM6MT
Quji02g9siPrmnMIAmX7MeSSEbiL6EtTVeMtNkqh9maZBSs9M9foVkA4uGz2jp5l
Di8wn25GV7NBl+BLoUl67nl4ZZKcUyIXj2br3ODSQmwoMEZOGnAwScbu3YZgqP3m
887NVxsp/0ZOdvP1irwl5zNSpSrMD+jyqYevxXdxNPybCcNWQl6pBdVI16mZaR6o
AE85qMYvvFanl5WOTX2c7XjTdvKN/GfFhi2Uf/MDu/zkVYTBTpQJrgM9yr6TMUPX
O7/UMPjZbzdmtRhXDBjrywNZBb5Ozqw5c1/d10eq3NPO8AxzWTGRNcmAxXmkpjdX
aPDxIJYLIcjwvnIoji9YU21xS/7Va1Qwk2HUja3zsMjfz7iEW2jko+9njlOzfVkW
rwRCgSDCuHLWRWN1FqxQCjnuh+b/RTsQXVER58IZ5AsJAcykqRNaKGZFWb8T/Tkh
W1ETsFU/SqmCYFW03Nw7VpJAWD4R1BjSkjDz40osxHfVRIixkWjor89Z5RBv5tS/
q6g0DSJ3/aYUpO6jA9oUaGBdxBsbd15Gx70AkOS9r0+YSrzvAhXHgH544HhfVxuh
PZOyaom6L/9RUN7lXdK4eczOt6Mku1VKQSCV36JS3e9rB9XXs7tMYI7N4B45XQ7X
3TbrX/HQdLfEZWfaTs4WULvctbYKCM5rrlw/AAioFXjTlXCEu6Z3iEu/3vqggKHJ
K1AQ+KLb/6I/7955Rlw0ZzaeQyMEndOhnineQpPknxe5bvz1gyAqJMucE0G/eVaU
PiONV9I2GTO4PrTTJRub1CPFGdxBnrTuKw592XGUaUPon+aXAglMTJMAc3lq3qmG
lfgYRQRWNRsGdomqeN2RCEOuGE/jyY4u0NkCMfW4L+RyWAylxrqbTQgQeN8RIj/y
FJMdC1ljcu6jC+xYOiwuONOSPxdymdl980xW4+yVgcPOOOK/eisQ1WNAfVr50RIN
sW+657Llo5Ft2joUMIsr6KFpVFuXoRfXaEiV5aTaq1h449u5aVuryE1HsidrNU3b
RLS87vVHK5N7HUNohW/g4Aj2BX8c8OUqMYMCYHx8KpMPUJLtAa60DMbDvIfo2m6P
UoaGjgEaOcbJK5z+NRVGc/wT7MyOmV55cIpuW8xnKdjEUoaQ29QYNg6hrIQ0LvmB
opFg6hIB1MQ1IeOu6AMjq29gOqc0os9uDYJFmtouf8IHUETxBhZlttnm6J/y7DBX
qlt3YAxA4SJg5A0EdSKYtkStCpsOuBu9nz1GvbkJKrc0vHlfBPanImouOS7hzpAa
gEnL/m/3pCr61Y1L2CusBn/tnSiVZDy6bomw+tO+68LX1HF1CGMK66RL7ZC7E8++
Fuvh/C/N6HkieG7ws5vJnw1+Ww6DdHaIL8N4D5CNoG6BGu6F6+lQbOjpAE1I2SrU
uCKkACweSUHTFd45dBvntdm7ugjhe4Z6NU0BK5HaCZjQXtv9efdyp9o3haPYrCSJ
b+OBWE4NsAyjDl4xHym7+e20od90vHPA1P1UphCNay6oiV/DKjpyDTekCGu/Q5GH
4/ljJ5kDzMGIpy1gCCOT57Zhe1TF7q41lEj3ot/+iXPGcgSLyA0cQG5Iod7ayj2w
CyNMNc6HOSVBunZBIOPIntwxjz0rxaiiv1gyncg7CV7UcVKDnRWwJvCIC3DW1XOD
yJIOcpw7W5kCinim0MqXeXDF1mEQYczD9oL5THzoMSQLUg1LyyusOn8Miy46Bhdw
2fmF0J8Ijo15ANCzbpltFyaDuucLsr5IK8dlRHhpvPv+NcHa6pcjjnJCNTrUB+vk
Wk6vsAu+fN49nJq8Z5mDtcdclzsbUfsn2TmnF76IWlQngNAFY66RS65OujEPwlDh
KvonAeMNC2f8yTloRTSESm3vC+XR0KlSdJ1cmx3yPVOVY8FLnYiQDyESM249bnqS
Q2pfBTOUDeq5NKdHu4aNrXJVWpylcYbtmKjDR4BoXslwcaum1JuKbSRIXxuGnmqR
7J04dMT66DpcUm6/8AoadN00UqVMv4xHyCXfsbyVMNB8qJXdYZlpMXHxfAgZJ68j
sTDPI2vTxpwNBPu3FyZG7vUf0+ru+xSQ5PxIYjE6xxEYZmLG+bzlnAPN9oUJ4aPb
TJD7ZPEIKa8+uOUTBct7nAovHSc7nDszl+/OuGnfNcybPHBcxCb/FDn7bd6gXjDy
kl/8zyogJ7O1d2cnvyNAPPlxy7qXAvVOZxCxQtKX6GXOnH57CcQgw0PMCMWJdgmy
smZxyerguVSAHI54+ykSFXQG+xm00SXGHvchyA+cr7FyXzdWDEGLpgwc0K8y8yAO
vZBc+WoF/O4BF8UyWmQGDKQlKVwObE41qpHv+N1vEVcp448NdxFmOme2rQBhlZ7n
VXRwsEtV+/90xfML1xE9+bgBpadbKY6EwidUN6Rr4d1T73WonvNFrTV06MewWZxE
EP36lOB2171EhJw5pqPfoXaxtQkyqtS5gm2k/6wbvEnbI6OfNX4q44qCtOmFCQiP
Ga6xJkF0EXIZqYeeRHDdbU1ot8ZNzv2lZZ6fApdnuWpxVskBySlmAQ9lj1d2yjwf
A38e6DXQLCQPAwqn+DwjMTfd8BqD4rPp/YykWrYHihqG+9lCVRIOx/XbdAH+zmqs
MGYywMQYdURGLpKfaHulPxhnaBhxkjGfH7m9GZrtRx2X2QAGeKZHypxzG38jtOPt
Oe7JnAsFnmg+q5td5+wdn5DIrkiWskq8cXKchgBoITz9QnWr55tuMzX0zOjEH035
B7/zHm2SymXuLiHCg3SYUYIN9/u7DxvjnH5/5Zj4c+s/RuRo9Ia7m+y5bwKGMxFr
Jt1z1iGYo+GkcBAwGk8ODAqMsinPkVL4Wj5LBTbtDEqa/wo8NXfCU/Li9JSE8Gm0
F4F14oYCc8NF3SEItgUtN1H/ZjzAB5VTkwuZ/QKvN0uDHnd3tIxar+V77RgrMi6I
mdggvuKjVd1VEjpP4PqBMUiut/6Qaln0Ov6+w7PDI6orics//HZ8A0GSYilcUU8S
KJZkyy3GuzjWsyAmvS1hV6z2BQuhIwXpJgaORpVqX1G5eLeY4JisWDqPzAF/karU
a+qxsKUMU1TO18AQcb7FBpNxvsJaSg9srztjMhMpfuNp7lxGPBjpsm+RdqC/rpBd
7fb1V2jSKFb/mhdQTh5LTkLKN8qK28CAhncGHDvnp0B4uJvU+N/SsLLiPiM1lkNK
l0Epf9ezExYYahzgB/Te5wlyO3WpQHwNUyACy9mtqavWsvlqMuzbPK4RkUrSwrxj
c1+RXgP1/I6uVo2UPgrxIk5k90R9ZoiAEMl1ufrKhZt0hZKuNuwq7PSJqevEFl9F
HU+H5smuhWq+k+wC/otYa20n+An01IuKuHn6zjkZj/Z9FuixA610YJ5r+jdBhA62
+eSVHqWuTZnbZl8iudLVOmj5xHo7TP8gJMnaRIMPEHl+zsUENSTgBRT7jt7Kv4n7
SJFiPZJcU35nrE6YxpL56tfChBVaC5j03vyO/Ut0Bd7Vni5uXaqYhAVrYFp9rGOx
FYhCYgVxizPyL4h5c0gTzHBB912jE3Y9G0bjPy8vOjSl0GV2tDc3Dltcq/q1X9vo
XYBSawuLviKYQFKFn2sNBNJPYK+jixSyp3PdnGRhr35lwWXjDiR8zWVx2OLMT/Tj
VxcqtyykYW+Xhf8V0UhgowCcK3ZWI66CS85WhIi2fz8KRO+ehO7AYAdrU+Zpv5bF
5ddXGgH5vJJoCq6F67ni1j/6Lc3L7DYUedDSueJUDinZZ8Yuy0jQnizBuc8eY3Fk
+Dud8fQebR3n+9EP0HAOSkIDPtXNUhTb93DuoKHjIgTVh0JQ38I21y/QjGv13ZiV
9X9AApkb07q9Scmj2OvWlo8qGeWK99m0XDz9IwgRW5XFLXL3ekqskCvZrLspK7Zu
1yxK4s6xXGOkXwxZ/Y+4KW55A3F1IO28vy0Jd9PGEHO1vRubDj0Hcy4MO4VFALFo
9kk+zKz7iABm1DKvQ7i1aGiR7PSiH8eWMUhKFGoe+3toRr/DlYASqVh2nBDVMgB6
jGac5UvzaxZmFZ09HGmSKfiuxlJhjz/EaI0DvghhZzx58eNhAApS6oUUvUBrY21z
HHVBQ+qqtWt9WYf6Mu4Bg5av1qoRt4ISA+IfQpH57xfc0DgFDjs5/GmguycOcjac
H45axnk9EuU+tiQIGdWbhk/WNJcM1O1mrjlIMscIhJaq+5itvEJCVfmk/i2RLsQv
9Kr1nkEH8oNpUvwYPIRb5fpyfL1KuwObsWpMBFk1cpn9VmWlQTJR5fypPswLXpu3
+tKjYm7MzDH1oBzedZBfcAB46P2Pvg6fJ9nhHJUm/BSAqAfUFMtlUxS/hwPp2Ou7
+eZmIyzzg972dsZJUWkdKHDgC5EGqeN0gRLGnREJWEXV6pgt4HnZP1mkZ3W/roT9
x0HsxPFKIyIBIe7v6+xz0aXE3rBTk+CdJq27jT82R58qTD8Q3CgXRmR4YWge+6wf
/Vjv6iHVn2+C2yPVSM7CQjzpgn9rS10a1RRhyphekR2HpHloGDIEiq3xVT0eR/SG
nJiwN5k5CFXq8Nw11xeabdBSOfjq1AmUsKVckDSb0uBFN7HKM/PRp8QLnIP9L7g/
AtJ0jv0lhPl1lx5Mx++6agEOwxnqqlmzF9moqrDF1eUj3yCP9Vnx8umukLOEU79r
fHLxxE+U5JQK/QXbJ9tBQ7RSEQWC+I9w9TxBWEMJfhog3p3+CxJT8gmke1eh6mCy
anoMYCqjztzePSoXEYGo9eowA/9WIoCin7V5uFM+GhP9ys2uohWLDD0SW7mgA5qT
oUe5WWQ1a1lu/WO3MMrxL/OAJ18d9jI1HoFJ/7KmqG50+qLN0lsJEf/35fimztjt
pCwFBVBWUqXESiSMd7+4bgArHT4srI6rX5yMLy6nde9YIEBZCinla7739aht7WGu
tD8+3B/4UX5DJ+J2xHbhvMrpivSez6O8AatUlW69H8DR5RC6rxszJUt4ij8xIjbP
FdVpe6I6woBfykCR/a4cu8cvQaLLJAuZYi1A9PG8LJgYfu5GvySDooGuT6B0n+Ry
tH7nAq4AlLCNIT0y/LaqhVn6anX10HJ5KXji3Hjv0LfTR/HzyWF1I85LSpdleEF3
kaPy9uHaN4K4t7Gi+w+4vxdYP5n4/MNNrOoef9FbTzo0LttcjW374+4czJCnpU9r
wH4sgSSE+7M2dz6HA91BlUfi1/Sr5KGFu/TDWY64dlt3pcEvnLSaSIi+k5alfCP6
DNS53ecPuZ6nXxs/p3LUDP9wuUEWvudE04uqtIEK+oeKgKVFmJ76JONWJyL9IN6C
ueD+kdTYJzyjr2XCRRcLZexFBsspXibKcCPeQDwRAolCQqyQsEwkGpYv0OtI4F3j
aquXeMl5aPGOFkFxeB+vRSdpCWdCG1NXjcT1rFtRptn0JoJzQVdek2W0C6CkGJq7
BFEBR4ihcbVRqh14liO7UXn5JZUlGHEG7JoPu2ZY0+R4wi8kenTaqAmeo0j7hkzJ
vPQLW5bfQ9PX/s7oe4rGDJbT+64ElCcdgDiXwxX2q1QTcMrBGvvNGpgM/gmyJror
5toDjX/9kWyW8VfwAu7cC1NjtXpQWPvle+lphnqthypYho3+FTczkJfHFMBUT4AE
fb1elpxjgJ9apg0AHNmkgLZr9nvvvog0eA6Z7M7hMDbVCJ07pZWLeDydo1NJj77l
sc9/ZQBWCZ80Tr8DG5JmvN1yoEwq+34FBRzJ1cMX9d6JhXU+kHL9/P8J1V+7jXmy
ao8rXPxbRFTqu0WlcvMA+hCDe7MRgebYv1dVV5/bcVHijYb19sw3BRYijAgK0qZT
0rAHcwSRWMwtQX/HmZWZ+6LO+moQLujc5KIdmX6v1kxp3Y/vehwOs5rObAenTt9H
MACHzcX1ktKJyjt0RJ91d+kmDJM9e69UjSwel3K/HtbK+v4Drk/JtM4wqDg5PH1W
xtdMJwP0gJZ4BgnU4vHH1/o/38RpigGGF9jg1oKGZBTxXmdiFhzggXlaBIRjXQkM
nddDxA+B5CjERkemG9FePnREPeKLgjpxSmJ1xEadnsCdPIE6vCWKqBAUq69gB4U3
SO5oaEK6Vvpr1b0Xx+KQq8ux7ClvRF18WJSuAHMSBfs8FjlR7Uun8lhyLlo0cmIO
NocbGrPWU4QZiY4FYm6xNgxcm8/GStRp05DPEVDBLgIHKoGgLRtUx5tOVTywKS3J
GC8Q9Y1DMbQiNjgt0gCmRZ1C8sHv+bkJGIF6r/YVdYWiuOHw3lzGwilX653049eG
KB6iaKFWmTTA6NkCgwjwU4KOuQWw6CXHu26FkbYtwqiDVRA4oW97YzfC++f1wsr3
h84zY3M07oafAYyvYtUpBtPBXGLpAlueD0742lIfkn/pgrKDh/x1ATdgf/fgaYiN
uwmIMZB7Gr5R97fyq33m9D1ECC0K7rhUkrESUwyWp8Dhsap3I8sutXLYQSGxICtK
qp1jtDt0IKc3ACE2QsZflSRQpeuy5wCHt7Fw9+/gd6UkF5DqCZWsUE6n26iltukl
agHMmlEiMhGd09A2dCk0VOiTiAq9lCt6FbRH/GjP0/onu0cKqV+bKz2Ep8cNA0oF
d/kJYwRzCTX9jYqH+zdNLdD/cEJPuR+klC8oJIodxlQvkAY1sMAoNIjvY7ExgBYC
anzq0X37A4LiznxxCkvOn2MypwSuv5OzOndVPLxGdpuehO4qOTOc0wErvKQO1uhc
ySzHb29zLY22adWRB/pF2/Pfao205M2YHTJ9UnVblKiIG3e1jy9/06CnVGurShtA
esVFvoOAYihvGjSeoG2ES5SVg2gVzlDbFnV/jjPkDFoHYn5comddjtSDo1wbmiD+
3pVNAxJujsSGin+WmwQkTSdkeCty/D5IzsmmuRAtY6jSAdy9do6egohTA2lg3LR+
jeghC5JvAhIlPelko5XicR6HmwhfLeqRvkzs1By7MF31iGaZRHlvCpci8tHWynnZ
lxdov/Irg4cC6oTHtACTC8//otdg+6LPpNMe6Yr4L39B+WiZOLKWtbKDoR99VK6r
nAKXMEVIpB4LBRoPKnRzUciULIpgeHf5PlEk2MM+8dbPIZUn9naXN8si1wHqnjbv
qH5HFdolJe59zH5fHMOTDn9LEzANIMK1RvYhYqvlezRLw5hQ4iQk1i44oknp1SxB
oZTqOSDnaJ4aLmQobSlMUzlkFkfKREYSASvbgn9z8DNb3qVr/OnNIYxz1doSxOAx
8Cdl3pc5xGF/fxeyCqkI7bPxHik88sOWFwWk3oc6aRxNJqtLD5lBmVle3Z6RkWwN
UrKX8yaZH61b6T3fbq2USG9aFIl6tUFzCJJk6AgqaLZjY+ZOq4US5WVatuQc3Xzb
HrJIysxQIeUe6Bg8AMpnNkek7hMUbepOzahWvMSsjcUSYq4w510wcE06l3awjBlB
mp3JVoYs6CDNSKV0EQHk1W3rJ1urxxNeCsHHDWebbehuSx9I1MgOKsceFSkD4dXz
9bHhlQ6dgRTcNzwxu0/NX9vzSxUJjUk6+802bqbzd9iufwGXhvaYyJeila1h2+KL
B3r+PKet9wPIkln71wx+V3rgUqEyZ+HsU/99j+Nch2bwJtJeTtNaN3fknpzSYbvQ
iI/BxSFe01iOGpFMYRG2nOGqyfXLwJxCMQH4MR7Q+x4trZyoRTUq8u7QcGgguWL/
spWQufIneO1dCQlekyQug1F+d4tOA71UoqAoQliP8v7SVBV6BRzPAv3c+JYSWUw/
hy+ENW9NGHl9H1eXA/Pp+L5jrlxPj0OGvPv1g36pNXX/LKLeg2HYxGwDeUSdNHzd
JbZryKy8mgLOafv94TAjxVNND5A846iMRL1IdbUo37ryjUv0FNXDjNxjkao3OTJ1
La+qet+XN6X4utXKH9oHp7uRdYuM3DdK1Pi55OMvFwtTpOHqyeEybw8QYavlJni+
iVCLisYPW7qhsNE1OpacQz1Z6mamXhu7YpW/kxR3J/pD3DjCDCSn3c/Q1WPb/Isa
mf099n/Rij2FOKqLsLmlmfeikP/UwAszmx2aoIlrdq+llh5PpXF095kaYoBFIAdI
DVAhmXh92qeKFz4uXsDnRmF/hYcv3Xjq5h2XBFYuEH3oASNGqDbkLyT7QzN17U1b
H7KQ9Td0c9UTdRDpaT3SzcDOGy90S9C+fJD/d8iMmhMFLhy3i1iUi4wlbhP8/V2t
iTnqy52Yq9HHE07pNVZEziUP9FPrdCMRlzWuVuJaPaWIdtcYjHUeCIoRzWBjC8KA
xyiuI6FHvfO2IEarriFynILP8kKBKUdtUgBg0EnR7Ar+t59QIlwc5jSzWIhQXo+v
FffLFcOzOARsmXymKfUCQi/opZUQopXpn/Ft+3vd80einq4t2Z9qngb5PIGmiS5U
eO3ZiPdGp3VQA9okGcNlehdkmPwYG4mTwpXl0Px4HOkm19saSm/CIJK7+wRUXjEp
ocQs5ghpbLsR5C4YUnj2L6i5pSvb7VDENO5p8Q5cgQU7UJ6yxrpikQdEzpMUgbqb
Fe64CDMLQTxaV6U16wwIlr/mubEIxTN5wJslrRrn6PuIW04qmA6iZ7vJZAdjwvun
LkQfwwlT1lyIDnR5WbGZI2LOyiSvBeLkxhSn4vSwEXyQ7V775HIXo4P4/tux2R6e
6Wqh6Nhd2MGfJDfbYS6xGdKxj3deyiytcU5k/Y5KlwRoICVktE3pxOoxocm9cLlC
dm4c2ExDYrz93qBQ6nuDFWtiAsKmGgcH1euOgb6CtTNcGsosM3aYw1V5SNODFZkw
v+5wS1hlN+WRSdjXgg9NkJoAmAeQKt9etA868Au2yw5sdNvAfkwnWO1wjCkQr/gc
jStlBS/yQPDQh4DeGOmmCiUKHZwRUj6hWXc7vZKpfgmxwwBeClmYy/Ga9pY/TzYh
BYV9ZsyW00C5KDPlsu0Ga8QRZRAvbnwmU2HjxwX36sp9h76gdv2AYnUyO0BEGUft
bkDgEXUmQcH7juzsoM9vnAWapLy/V02vpR5vu4UrSETmdh8gi6hY22axlsOPDArT
bZAzT8oGxn3iB15aJdsNKCI+YJIfFqbo2mnn/QoQOzW98hVMuq9rDSDZ96KAbGIO
9Cy9P6FSx49dDeH5ef0Dnzg0ieh4jXKhrAiOP3QRp6Y8SJMXEeaT2tFE7ceHdr+T
tRRCxjyVZxEhl1oj/MGOqI2MdEAUDv59NJr9H3eFPISP44B2FvgkIt5uRk062amo
vnTr1SH9Yl34XtO9MeoQ3+3knkyuDWg6FkR6cQ5UqRADouDlpP4wC8zqNBQF+BEU
8JBBb+D1TUBZVT7MyV5nMb+BOQvS5FQUGhYtCPTWRo7CasA84MoxTvbvviiV8PEe
yXfBoN9hYC0vzmpkv9EdV6FRZewg4iGvQvhXpN2EGKMgSMNOO0EdK2votO5uLXIg
vXEBzWlIng0GqNSgrfUdX5B+y6AILcXTWiejHBCHO3Av0T3LFGLu7aTgomFEgmVV
cotUNcsqk9JtDJi+LEe+/EnkTyi6CFkLJnnwwPw19q8SpgX3AWvI5LiO7Ky46+oJ
VI3T6q8fvp4CXWX1C27CmhoUCcX3ZRfbS/PurgbfJ+uu2QKOBYEi3AphGVwRD7PV
ueKXsJ7VrYjaWYSyutCc68EiChu+qKW0o0/VUb3u5EFT+inzLHnQdF3Ak1xTmqhe
K4MOavI5wNVfSHJzMkcIsTDgBbxA/LryqkyDOAtjfHxsMJM3b97mTJQ8yDLrYu9f
qZ6XjK1nmdXxCGK607CZy1xZLtO3gaRegSCKXFmoKlMYsUm+/qn+H9IAH4N1VKAI
Z3RazHQIpjj4dulbwgjD2Lydl7NLi/wLgKuPHyv4j6g7KRhV7v09XKdvkoGRje6X
bdCUxmVipM/6l1pFqv6acHV3pbEU45jKDvxDPY5KK8mEDD1o3iMFsthX2VqcVPUZ
XpLyqHsWH0XYyTFE3tXdRvw6SQywDQLWiqjZyg3lsVLH03HQk/6B/nqbZvf45T2F
w8BlW1HgHbpsRqRDddJMEHZzVp/Lp5ewTdwGazNIFlVhpsAFE4YK0VlOZPuWs6aX
1f6+XtfF7kUfYfHm1jHzEuQJWZtyDzVuhy54EwZcrXb/iyWWh7fqCKXgFy0RH2kA
VOKlG72jFx8KyxH8VRRjkaJTPdD2ZIr1FKPBLK1+3dAtiCnE613ZuFaengI5UmCS
+aV6b3TOq5voWVgU2+qMc827Ds5+QJJVf3UquNbQHQAib/EVxrAlX5h4nYY6BNP6
uDtdcBfuu7xYPXl4WbBMvu7VU35YJMGFQcVwqShhzqMJZdwhsJHg108eczkcrwJX
W/ufeK6RLoDJm+X+dmfr2sn3Ty48dV7+7wq90vKUr/LNnVuIxkY5Invtiul2E8Zi
VkHeqPP49UYBUKsJC5Az/FawPNHcA/+ICKNe0r9ET1IegjEZw/2/NVDtNWdFa5Pq
tf5tyOG54EkmtjnFvpnzuMQDeX2SV6cvS4Nw+VucR6blII+Vy/JE3+3+WwT8tQhW
IeX6q3vcthmYfpyYkxIWrXm17mC4Pl4dad3bDety59yAOb2njdiTGFKolToTGdAb
FeR6Zcg80r3x3oquFEU6qNWC3+iQdYtCQY4WBeWnz+yTpyJB61xyKRFVyKZf4R69
yP2laYxUy8cVQZWZAxQKTrR/rVHLnJt5xrLjhAsavrE5pUQBSN4SnbZGUdsUXw2K
1fnW4YqgJ26lyGajSrbk1xm8VuHqDTO1K8aCan4sVY8SakTGsXn8p5AbHKJ1fAD7
ZwxZaL/HvnyUTCOwRSFpKa88VfvBS+FhWLO/oBdBh1CUgTXooDNGYz2NKJz47bgx
oYMo6W6H1g6KPkEY/FXa3qfl4580OTYsgR7XzkyTT93QtSHQBjuAiccviw0h0ln1
oHpO5qA3bsGReECFeZnhgJAuhMIGzyOoe330Wo/Qigjr6MuNRzU0AZXMRfvSzDHV
iakcbVUy8acXVS8B5apid28XQ2rD9tN67I6r2NEe5y01J9GRygAT7kXu5piN4Psu
NvK+xFAZ7A3cC2YGQNzNWObR8k3SQWo9rHj03wGH1cAzA9AOWyRkFH53HGVloda2
s+pPKTLTWgeUifeRnMGIr9FKc4m9DQSNk3Y3+/NoQSIoaiZ8rtRbI1hPbVDxc6lZ
WaxgAgSM7rYovZQBHRObkN/0ara9Cdfs/kGtyhPETUF3C67GAKl9lugQvxyO6kZp
nmksHHv3ypH/M3HfCxzEyEWiNm+PxkyzS0y+48WBU4mZsw4cLWfOw6czEud+/pyM
n9crjQhQsjWOSlpw7GOtdxg7fFtjZ5E8u1FiwkhcrI/v2eM+RYWDHeFsjuImssIA
3Ch9dw28qnnN0GI75tIY1zVjXOHHCstCpHu+SEny1b6B28ejrUMz/rTcKcKT7CdI
i2OWiA46GgcwF46tLGkZWr2HWPL4Grvy8QOuJJSS9dlHXAvYgatloQf4qNkPNffb
vpket/4mF+SWIZRyMylXycRI/geaoGB/8jy/bhOrHGXg6Q3SlhPX4CCH83diGX7f
d7qyLBOwrXfdXTHx00SU/MbMSB5IhW3PPhMqWQAzqYINTVV646zGk9ngKAex6ODb
R5/t0z0hBQ3Z5f2YBQh7rBOBThjDG6S1W0P0JixmCMZsl1TjWfHZnMUziSq4KjsP
xp5Hkk8tlMx6yG4BEKVj05F2ZAA18wKtUSAAtZSxeiHHaFEKIr4ejIlj825Da51I
wTxD8Cp8ryZUkNhtl77KXKoxH26T1J49LNGeZZXeKcc2AJwrn/LJziuaLe45Yv81
UOazSLDCUeAez/4gn9t8aZh2MjM+2nlvITvyWXjSqjZ5NW1gSEhY2Iv/1nge0O9j
+LKJEZWIZi3gf43itzbdNbIo6rIspljYZItp1zIjqZrk7PWbSQqajfFk//ZOd9Jf
rpz/spaSlEWFfDwVFcGq7Fsytf5B927VnZLChcfifft8UshGF5RhqbPLKmHgUzxj
gX2TwGFuk7gcofVPqjn+QY57XurQy0BBjORQr7kgG1qhhRry39nEPPp6fFZ9bnbL
fnCDTQE4ZTlK6lblk/F7QDH01GXX2WIQ45dXPOWJtL2ZQLk+lUIkt5kwrjjhe/eU
Z1syn26p+4zQCDqsg1bZ++kkkCtv8AAQm9iJ9MLK4ird7MyAQQFT44nGjRZ2ttmB
+rkes0YSxZalFGje6JCXhjKrjvHpxAgURkWvmNeXMAAbnXK6O7T5TANV5Eqrh5JT
f7snrWpclp+2u1FSgYOvLxpk32QNk1fVFWn/69N27q/G7hXM4Gok7PEo6lKSzorg
Mxu6J0MEO5LSDrhWjMUfl8bu2OaPbSS26Dp63rhdW8R2T2MpngH3JQRiH/pgo7pm
LBm9wtG3dRoHTPaZLmqnrQI6xj3LqlM5B15ohVJ8+HWFKN5kTleq+UWL2yTX+/ox
UKqR8Bh7AzhAn1RcE4+ktp2b11PG8xiajjd+amwA3mGbPmdepZBmRhsXASLQ3r2K
XAdmmSnkC1/Mlh6rPRssB30fA+lK/sX9zpb/ZPFkMlAIo/sAjLOXPIp4EqXII89K
q3G2S5sqkhrfgBHLW9veGKWcct7y0gxJ/RUJ2+vAEg6M/wEKedaRaeo1OLPjJFaC
/MJWqAimx4NVVLvhyZ0A+XASADi9vvlbf3QTyKAnupNo9glX1VMQbC3KO+ov3gw8
pqsrPVMwHNdn3kLM9bAifbT6nPEbKu4k04AaAETKlimlDDWAa0xjCHz+0KS1YA3x
NCCkxFqdcoSlFC7ANkClIOwn3/z6yGiYVYkxSGePNDboC9westwyzCjM7ZufV2Kc
d6rDv7O3cpJsqXtoqX989KVCG2XmP+ekh2Gx1uF6aKX38PZhbRXZv6MV2oOLzA0W
nDk5XD1wHm3NxQfhuUQ8gYNvF6fEHowa2233E7vRIVfqtglSC4ri/aSL5A61IUCP
hc62Dk+68jB6Uk97hXGrq8A8DN/WcDcASmF+DQfO670ONV1NTLPHsaXAAIiUOrPj
jTF75nuEhIO4OPI2Aht6xOUAWIBbKfySlZlSoOcWRXh/x0d97UymhmXVXOge8NW7
wyFlnY0TMhR5ZtOq5WB14JC97PB9p9++pm3H5KbdyWz35Z48ZJO+cJwsFys2nCgp
jcmMDz/IV0TIbPaOYAqTTyMIk7Mi7/1zl85dRE0WsUlhR59oYZnhg2bEtLMDdeC7
/G1XpamuYPMVlUHcsXZv7BCDnu6Y03kksRmru1R3lvIuzl4wgSDwNRttpO0hwYPo
/YH2TaFbnaEF51V4HeHI3syc4xS3+yftALLJiT0sxjqkYzR0RyuCyP3ckot1Qa1s
hRderL2rVFJLJAToGjNfwYpAnfHDYib6JnxR38WkmNDePOCRH9fmZTQkWFcn46Ui
JUtAbl9FCPEYtse83paCbsExdVcnW1cmcrv3Si5V+heoCIAFOGRtfvLXKQv+7WzK
0KyWPquDLGgZY4sEXEdPQeEsRklLLIayhPXJ6LOYKPgIoDm/CoIKM57JrMy7mbib
zZziXELmvbAE72lTtGgcN/LD0MHI8Olrd/93GGDtYNnHz3JhkLy38OVDVGPWhsJm
qmIE+wS0QhYgDLUTtLAk6lIJmHQFJAFTJ1bS62bmc+K9DuD529KXvUKy5DILK7+5
4nX6l8hSMjLDh5qso8sa3gxJId9BVeM6NzAzpxyyEU9X/Iqzal0ZniqobwnACZX8
aSac3ro7IugaBKgUktim/VM5tYCTaobofSxfqC6ce7fuUyFSExBqnd0W7k9M050G
uBQdr4OHrFxwxPM0Q50OjxN8vmL2a+5bYkAVWnyvsSR0RQAxcB6Gkqt6iHVP4IBT
J7KmUIcDxsf4KYpDgYLlvEx7p5mte6E3S6TjY5gkamedPiU+mZQB3ZEaM+qdya4Q
dBSerUMqDCYJFVkB1aFw7HsS5NxuDvUsmCMiGAjA9rqBc+ttVN5rXh/iQVrku+VS
YRA4+c3sSN3y3F0ESdhGAKGrPYoHpr9bFNkaTJ8imgTFwpyOTonpptC4CHdMLYV7
vWRK3YpjfRgKzdV4IG29qPBTmJFuUi/9XyJsVwxYdnD5Pzb5s5tlO3TEePolle69
L/V87VR3D6r2ydxqGmbTzMaF6N9nN+YFzC2Lc/EPqsSZvFfb1I9zBB8sjFMiVlVU
iDVK+bXIZFqfYETp9uH4YWJwazaSOrq3PNr4vC34K3UJed3vQvll1U+2eUAfUb6p
wdiDNypmWMcvSa8cmJeX2cQwJ1CpBRm/wy4cxF2tg+YgBjbFpX8Rt7lyqo1UIW0R
f1T5LnxnQwdGZTOt/B2t5B4exbdFe4gsJH8QDrkpCXq8dqXuMIduCWGDrnXbJpa6
c+uDsxMlUkJK7utABpL9UQZHCQ87MgZzhmPusgI75MZdY5b4ZrlX1cmOcoxqf6SQ
aUTDJtW1IAgEBDMT6Cwt/iEISDKlFDzI3aWSxdtxxmYTC44tksfsgVQYpRj93WO3
DxtfRCgdEVtGlrZOtbdot+P2GhvXcue0ZU2gI2rZrXcrVA6feP9BamMJ+lhfKl2G
Yt9zElesUVLm85t2BrGYKKTYq+3E3/Ang1buemoziY54O07W8k+rb8ZV8hYdZ3dt
GhNUpfk47FnpZcMirsDPnqsCF3CdEzRJG+zm66ppOhsBbfITH+c41AGN/fu4ICtz
4DJfjr2oV8NsogDrvO/PClUEjv6mlyM4NsGjUQ9t1wJDxzdqflLxQto5y4fL0YEI
zhxgA8ZfUrPPsDOOfMPMy9x7soyEVlhW+lRsM1P+VBCuugYRDJAZqQoseifcobjF
B8t6TgZp2fpYT1DBUEfEkEEl4SZKr/AlXW8j4lCCAreBDxfxDFtXXzkYTY2a8TqP
ipKwQ6Mzxn+VLaOB9lznAPxg9AaNXTkMg9XpIPTZLUPYVD+xwKg7LUSQOe93MdPZ
dYXRmNreRyHa++UxFiL7Esqoog4RTUEmhJM0ODq1vmEM8uDakFweUoiDb19lPXO/
5VbmM3dWIYOvGIltY0W0pLKo6+48BP5fyG+aBOwIXT/FTx2czrfQGqE0ObS8qiXi
bV1Lcvh2pxRgJJIzQNpub/1VhAM9d9Q18n1TfWk3BpufWaPzFlfg7fVUlDOs1jsv
f+vmlGhmNGAuVSXrIUfubmAuuZEvG9Sufr6f6iYtqeUCrF08ZoBbGUak1W7myu9J
XUdpGFJbMDIYzyVazdkPXJq9XThRWND3dQpoHfZnSz5eWodIkYbSFt/fg/qN8mpE
oTnCat4e/FKjskwdiGO8/1M1FpV3M8knX7kYZKiXxH2uqn0XuQKUekyO59f0BD9E
JYgpqexHYEV6kM4v+msFIuxsgg7DxrGOWUjmMwhpMqFYwH9m6QqzMdJm68XKxOD2
YGBzFP7cNkQxxocEvoK9bYhSHUnM/dHpnzFybrqsxEp7j8uYS4w6obTiMQT88/MA
aB2L6teObSQKrktOa1BHrHrk9WeMiI9BIHvC+RUNvYdZ17gysOTJzRKvxAItK+WP
ppZidwbDampk+PC0mhL+WneylE0UApQDIWlNDc206KvjgwOki+gYMlrCqgsV2qng
KbNqj1QzvmAUYD5ZCbwms44xkSjwwFWwpCkkR/RaHD0IG13HHTulMd3CX9jHlO1G
dfjkcmR7vozc34KQ848dgpXxoTZsw/aKef/qOgOdhgKBjYG4MrthzFF8Wuq+hnK6
57FRwXtK4ri2cy+pVM1Z5tbqNIfnPcyupfGRzcEMhQ9UaqQZBpTsGsqjHOiB4H64
iHu1BTncKAYQE9dvoibAJUnQlzJ8fF1+mI+CVeZEPTX8BSzZrBHibK4+GudFj/0i
Dv+o50+LonwzEf/unzMwrOg1re7YRba9Z4RlGqbBEirdNXUlnf/Q/bwzyeaWpSY4
GeHcpCm1B5rL1lj1gkfSomHJ6nEl5ta7Eo1aib+1qxRQWPGD+2o/6LPSc7kQSE+w
YudpbDX63W90WA/NoCZ8PqRkVLASlY79O5aRwR+Xn/9q55yh/WWiKeHGYuyuCkDR
IpTticwplTw95/LTyJOAaLhJnq/JJe4Mzyngd2gfK8gK9reBHhHSqydt75VXas+b
K7ZEiF7EoeRsAy8R8fE91iF+OBl/KnhQ7xW3m7DEzl/JhOqvsnfKzULX05Hj96ql
C1W8l9l3Nb9YMLEsbx6kYaX9Sg7RtQ1pVdid8pavJRIPRFAHHJo+hZQ/OrkQhSEh
hr8aB2DEpLAA+/qkeFhTZ0uImPKcav3csrHG25dJ0/zFd7zKnnPN0MNPnOT9Lq/J
AqMju8z6IG5c5a4QsO/Gpy/PoEvfVx3UN7+4fnZgmXhWgobF1e7bh4shw7e2PkUz
vSdAA251TSQ3npXNr9Z00w5MbdcXieQ3x0j7CMYD7NdPNdy21v3eqZUTCP/8eHmA
BGujliCzo9DnR9bmg82gumgOj/rwezuyI8X0zJRflknTluMctBvWNT4PPPdA3YF+
0IcgRbm/4LwL6ERBG/P4N9OVY6YasnU3kFML4AvNXjUADoMlDORxgflvWTA/p3tv
/d0dbehVmPVhKoKJdIDfbxLiH7HqmpnTB0vUBNxTMLZZ4KbPReyr4Zl08szVYlVb
WPc3tznlNdnK9WglyfoSwtm7X48bprmr3egUU7AeCbdva37+iY0ikRINbd0pxAGa
Uuat1GTE+2N3Ipsgm0nSfUSCIHRP+IK45kkinVtVq14JrDC4mhFkVye9RUmEdC66
v4Y8M5zwQyEe2Zg8JeA64res8v4K3c9rk/EjdHnCuMGQBCA3JiWVgyzOJK3mLxh0
w8PWHXJERUvSjMTN9QrGTezDtpN0yvPpMPAbkuKUvoch0RWPQTouU/J0R7TgoTAi
/GgwTqVoyMPfDBc1Gy0kox53x17EI1MvFpa2vWgBVr+1NBU5BhSgetdHPbOAgaMx
NMnwd1reBtAy5lK2JyW6mxYtuWQDsX9cmSH+Ia89NyOC4ZYYPZN4nO+j2FeWydq9
DnVxrwE9O8Tz7ANS+DEBrQaL4Q7wAmTYJ4FPXSsUpwVAG5kfzfyaZfwFQYfjJdXx
2hSojmDF8LZbnEvbv6LWznBWdcm/h1tfsebKak1qX8xyowWIAQx25nE6Y8FcUZH5
x4ANUG/mWmFg2bCUykKWcCQBeKw8EQFIeVQYg7D4TbDyEgWV1hFDX+eBwpo0NF+M
Atlyx9JPpHuOcbkn1hUMFtprisshRrdgwyuw+ChHhVPH3an61RL9yS/LCoQl5RiF
xG31In/1J6p8sCYkPfK8e0xzGBrRM1aITSYN8in501SyZ5bo/maSyDmg4jsX/tPa
fnGNXPyYhD8TYAIsH+ZHLC0O/TI3cnhZlxsS8wzxmCccYP8GEY26Y4wr066g8ymi
qyELku/02K3RF0mr30CMiVbYuiRvlRpeelT8GzBvZ5DSlovW0tYXgqNWIZKkq6Yd
qUqaOMvMB4lQuSGTo6qJ0En4d0nIwejxdi1/mmSAZyku6bgcmZzcFPmNfjR7aGcs
2gIGSX+J+QfUW7XUY61ySAwskLsqBuNraQ6dNkckUBleXpCMrJrEZqKjozmPNu0E
wcpuWIKGhU9tIfRcCF6RrtzbfOFFS1n+HbOrySil3g/tYTiWzmkAm+28KFDoY3t+
2YvWO9xJcmspmIVFLby3L7Tdetz70UtmokOOtrBMrtn4SlG6Pb9xVjO/p4zAFJYU
R3Z3inJxN7L4tBTiWPUv3HGIrEDJKxPXtwP8TGqPDOJOZDCw1B3rMIH0DP2htyTK
zimz9gZAtwRleGcteg0+cczy9ByMriloQR+HSLpf1C9lk7JPH/PNFEb3OhFwTSSZ
mSHyppbBsLk2rZlOPazlVffHVwdUhrS4P1pS5ytliqlzOLsTHIA7oLgO3GiOYHtF
/rlFhR4Bd1GII64zcOtb8eJePFakTM7Uuti9o7mLfzMDFX2QvZ53vabHdlKofQS/
JHIAYOIk9DbL94ZqqLXP7rv19Xjt5WX348/5IVMEbJTaHy4vpbtiA2ERC9HRzKj5
sh9rnMc41wGKq3rk7rVdVfXXmEPfWcjtRZ7PeC565XlVDmVIdMmej7Ip2WJWsBoY
k+GZlax95a0BPZ2yEmqyoby+qyQjI3ThiU31Gk+ga/bN9aFt1x5bxSI6sm28LnBu
/YPoD7aD2YKIF4K8lrVnXpeMjbxyfvxGc9DHdON5PBLpj2Tdzr88mUdaMoLtceSX
3XpTt1dYYAVbXI5XhzHbMGHXoiFF3JRUVH4I+XppU3KfP5W9rGIOGxsWN27cF3la
sDNBJ2IFA/w9jWg0eskTBBI6cGBmq5iczKbmDIiqR9J5B9MOYZ1oBPybRuCmlPkZ
2RxT+BmXFPyJ9yPISJGPUF5p04RYyOiOG8Yv3xf57eA52cttA1FR/ebmxCbmNIrq
1C/T1ydcy7rFIuiut/O5no1jqZ3IfbC4RGaWp+Ix1XAqVI/oNGJwgndiomlndl/9
eySXDrX7NRg730MjS4Gze/ZFxdNq8N7Jk5kEn791++ehC95MS55hldHEF8E2+QWQ
JyZom6mDG8Vp2Kw036PIrrP2Iq1f5R5y6LvlMpP1VltT32Jaz35OTuSTYdzxP4bz
TUKwG7g4UfFqNCN4T9WIbaWPnEKNAyIzg2kCNeBAFqiTLXFwifqgjj9YvXl6MvKP
otqMKM3dYQvTwMinHwllWavgfcJ3vvwaknEucUookgTSEM1Q5jw3nQ+aneZpGIsm
RNhUrclvIw1j4KtEhg8AXDhbC71/JN1LgjJMavJ17IX7RCzP8I9SxjM8TwavnvUj
lW9iuSYyFiZ2ttUijIVfrVY6zAWmaHJ8njqGwBnJaz0DB4+U12qxLWER7RsF7PB6
Mu2kWDOC9LLCX9q683BIgtqC2wvMTcqv2Oj5u8lSfs5H97wEm7uICAu42bX+8rfD
KcN8I7KJYIV8EiIe/KC0VOlfzi2l6i8u0rSX1l7JcxyfibgeMKoYDCjkvqTSamF3
5lr0S0vjthW885ztiz+rNkGi3mckRg+a5y0wp5xYIUILFF/sr80ltx+kFpKehA1U
nUETba9Ju5LL3vL/voU4vyUWVmB1xEy5pS7G0DlDaaU1Q1W+15dyEqgVi/mrTLr+
kjiyBCAg52GraRhFpeIi6ngwekW/dV+Wfj2/st1vw07pQnjU5Hr/vMy9HzoIKZGH
oHeyJNnKdvbtaiHzNJdWWl5+D5HbOpCKQ+kNKhlspGRe29hqZllAACIKuDdOYw8L
xTYbVKCMvn2keMFiJ2t7kzfgWqckmOpwySHqv5b9Y58Ffh0HNQ7BO5h4WUziZgdq
GAAq9CP4zJPht2cRp6De31MeLlDzu9KulGS6CST4luuGqNTua3ydyREL18FSUWbv
rjXHlzxWTBCSOIWpJfX/n0O0OrNQP/BsPvv/GTOtrgstrwBwYEWX3NfbO8/G6B5h
lUlr/6eqUDcUV1vS+9AOEjqrpdjjSTpVhQ/WSA51kbJXYrj8X1e2Ud7nYhdhykNu
DozHGa7w1N44unbg+cnGt6XRXxhiHWc12Szrf1bGoIezMDGvh+AvVEWAzVJ49Azo
8BeEIdPTstT5W7zEU80U/tBJ9rvZg2RbxndCmOZIEJRq8W3g1UnzFIvMT+EpxuKa
TKrNmMqDbhd+bLtNzAncY4Z+AekSXpHv4zXlM9e+L4T6/pqXwOqA0Q3H2+WsM2hc
ds8a8Ux1t9heO98lS5/Nvnpm8SeVMz4zDT4IJmckO0KdLVy/Bm29XVWSs95G4WNp
vekzdgkESt7keQ9esWR2jZzOilBi2X3eyagfleWD0xkLfaOwUfI3Xobo2Xe02Q6d
qUsti4GDzHcMBxUx1y4zn8AD/x5pJybcpnIxtMLbKbSO6n0udnC08kbqjk1piR+P
k05xqntMasU6NvRnoWsfMtFeK6fn1AEZGMXy0avxQjf1MCUTdcRAWZ9CzBHTrMA4
Asih18dyIflw0Ec8O72rJidCDEHm+QsBJqZHQGNXViI82BDULcFFXLkO7EfdMHIA
mqJfeb/aRGKwlk26BFwf5T5r9+JCpFiPlzwo4ggZ98VAzxMk7cgDbbkrtYaa8PUp
6Lc2wprwpW+djkTXvl5xf1HjKh/bl/pRld7yXfIKmQ3LFSWx8KyoF43zfbyhRcTt
0FtcCH7bVPf/N2oinUl3N98FD1lDjJvxm6Tl7AnDx9dJGft8pfn5caUWzDhqL+oL
CTJ9jRPE8yjIKImOEYi1gGsbNCKbeVIspSlhQ0LT/yWKJw+v6j+OUFpjkPCEN+BX
x/4KT/jTXa7rFtcypHvp+hmVJW0XESwjUUg5OmrYhpD67WTf9gnTH2VM9yqHFgB4
wPWVzLjWzd+YGQDETZqngehTdZkjaUbEOYEDatEB43+W1f4tcpSe+3Jy3C/9Ze/Z
SF9LBimeL0lzdIyxq7YbFjfW0fJFIYYG5lHOBRHHNtj5hN2XlAeekjPSmiCcg7pY
MQgwYJOO3Ndlrn51X2fgXFpcKxzZPISVxiQMR4YZ8JrLdfDlDPaFX6yp8RWtzNvZ
UDZmfRcEJLN/ItbLxtgrR1LFAgauaXf1l4XCsot4bLSeDwhjXHg4ueOywC+G7emu
7kc9K5H+ctjsV/UdOerC6hVFuSoREy/Z1XJA1frI2x43Ih/dmqxh+9k0syPA+345
5IcQSXmdfrMC0lnb2ZPNMw7CnxedOhBSfIZuGOqaRluVXJv68HY9sh5UEuIzNuJp
EdNXOX3q6w13aNVAJ6KPEx/q4mpDNl+eJ7Y4Zk+0u7BNZNmyGcXTmTMfmvXvCiY9
31BGI40c/R8+yaMZj7HMWGPpDtnXwMahKctzP0ygT4x/tBrC+zwDzETlxmpWC6vV
2SI8UruAB241Xpfs5cf8mSHhGTwb1v45h10AUBq9fQ4xS7xyEKn9noOlfIpeNBwE
F8ZrmF7vENu8oSHErp/yWTypbfRHg7pJBhqXhtqgKRqOziYyB96Urg36UhZMHBsa
6y1hgzN5lY5gZtB2adBNthQQFVMtjkJgIDFqkYjaESeNn74Y3WwGFZk670CANQOL
hma5KQNLHTxEeO6SKqXG6vlzofNrOzSkJP60H8Ko8Cp9rgFzLPPf+SgfzYvZ3yNw
82FVdq+twVtA/h79QLsDy19f6qNOJN+pkmpCtq/wYEJsokRtbH0W+D64h4TjzHQJ
i1FRNM5P7afpiOB5/b17Yyq0geXgHSdwJPCw6Q6Sah2YtG4+yhQ7EsskG/Nn9Vr3
sYehILwNS3weZcWwuQ14q2mlmX5We98DXFjh/qfIFPA8ZFypFdhFz6ka4g+awb1c
mk5Ga6Mx5SbW9p/Gzy2yIKGFghzyrms5GcTHSRdJSvnIynbLLtyOmy+xQ52EnFWS
SZhe0xFvgra+1L+rnGZQWHMVAJJ5A10f2i/72bq66MKznf+HvSw2ZqvzUz1N2JK5
3z5/pQhKOZ+a96S5twDhMn4p6oAoekeV/iZFG5svyzD79ANpJJfIv/vdTcN2C0tt
TilXJPgxy2yLsI/xdTftV28Nez3mK25CwQuUFTana3chgD257YNQvEwUdN+d2kmS
T33DqbHecDa61IeqKxyAMiOVOCpVOyH8A40dNfBd4ukPeKGQpQ7+cTM4Aso4ECfB
zrQ6YnvVy4kjp+YJBFdEcie8WpRrJL9eyRM/v1bcnHnI3Zd50SMOYAP8VhW7fGhH
DLgPaU7EbFeV1ygoT5BSAL3sS+qnv6wX4QksCJwKvISQlj/wznYyUxoe/LOttjet
fZOCbIzv/oTeylepnlLfgE6wVqq1AU+LlT4ul7U8qzE5hCw634e+2czom0dq7QcP
LJIcbP0/uMZhbCNaXXrxTBqJGT2TbqYzS4ktLOH9nfZR0xrgrg8gRypqESRDFZ6e
Dh7tj21ThGqczKEs5yY7DOW0M8dy0KtSs4tXLWKMFbQG+DFXmp829JsnVq7s5m0U
1AbwslI8qBa/jBVn1CKQ4ZTrWBR8t6Un2/eaw7u51zeSsDVFb7Tvwahjiaq8uI0y
xqRRDFuicvXn/t+s1/C5h4o/VQlAGX8EXC/FYpPVP2Aj94xaJ3KOw//HFweURTSZ
5iWgbumjpIJBCUtc3SrYky56oQNBmzdYu3X6VjSASC8cYaIBY9L3yCEfBVs03pMm
G1KxkNiNMetaxYFKJCtuCb/59Pt4XDaXl71d135vUKPLZrpmnxo97LGy0SQVjFJp
GDLJgtOsmGPYTSvuf2qtyxmGM50uF712c90SlKnjIM4dqBU/8XLwhAHydCMQrToT
eQ7DV/nBNiFMiav1NYcdaaMkezZPILjtcIY80InVls6GOucq549xmWIwMAZX9KHh
6VH16AMZclanP88iKeD74N8tu4myrSSfzy/+2j8zpxKs9hxLnKPnMT8CP6K29Qt8
mpXSL6KaNXWsfR9Nnu7TA8HWtf0+7CxjPIgzebXk2uwzyCQxnbcy/7i3wBzai0K/
AaGk4cA2mrCTKaGue1AVoakOqlBI5fihcMgB8Z4k/SsYPH8Euby/UGU349cGGK2g
CF8/ndSOpaBdZzfirkdWK/PoB6ugYDynA1fI+fxrGTNWWgyt/BuQkyWTU+eiIT6X
1Y+umm7HlsZKrVPQ8y1hypcRR5XnRe0LEly+om6wdqBdTy7EQCbHHnNAP7q3iCsr
HPloSNgR6rYZZfj2qratFrFWc5JVjrx3OFTWwuHONODKLxuOXj+6JrJpTQy5L6Cn
2C9YXiYqFrhpEkF53BlajgpRf6AcxEJwho/NJTu1gsVv3ZPpMb9jvvQpnrXkVvoU
RqysFi1j+zbyyk8AX6Htg2r96hqo+dgSjpLfutM6jjHe17s5QbR0U+2K53ceeiit
WuSBt/Qb4yCgtzT7XM7PpshmBJRROYrpfNt7ppORmIf16EmKZS7JEa3qi2Ih3t8/
/eVq1yjErOtgv3CRfs8bmztC/KLzQbRq4v9UnQprBMzfS9gRFYVvxRDE3Hu9llnB
NlscEsg1wIKHoSHawmOk9du/v/oaP+v8d8lT8teygNpqjWfmdjzwpGQGc4JQLftY
OSLXsA8KikDe4rqBriorJD9+Q0p6qgtc+Ni0F4r01RCKTeK8dcHvdODpDmAQDxSw
GfucoEngYbjenLBLXDVELxNVao5BoH6Q84qwhpYNT70YsbsfzP1MKqtLMeOVKLbT
dLeapoySTPcFsGtLwdUB3LJa+/UOmmIsjvKhiYcPWOaZi7EgHY6oKEFptA9pyiA/
USEgkRm6gnTNq0vomWjD2cenHXV9AthNK4TKC4cVDoB+Wfe68nia4XD52DzBbdrV
l9IYt/tchaq6IZPn6ANpCrOdoKJH/kaRMBEqmxfF937jgDb1RuHrwhfyXN0tPgsl
Of6ewh/MwK169jLKie5Z+MYUV8p86E/LCU55JcTh/vbqv/5CsnDBm7pdwxLIqszD
a1YR8p0uD/Zfnpag/ndNV6y+RGRg6Bwz35vxo+qK9Z3+8YJd3rMHQVMjfVJtTRBK
8C3FwoGy3dwAIFtjQo7717AsU+CmRebhdOb24aAF1q12nyiYpwqZyu0TmyfTfEIk
um6cAmYxWQgd6sYJEzDFL6lFCV5YUO0FmsKlB1B/3+AJxVlhgRKaFaqnlIDYpvHW
hPiE4OUveu30n5MhEt3iFWtCoCVVcEmH4QMWsN4E2avGpPfVOH/qSTB+h5ju89G3
SKfL2M4a3DC/j/nSk+SlwBvqj6OxZsCH7D+duzpnd5GLh9/BWu5p6G6tAl6ZET2M
ElLhQbPHyc8YE+gkG3M1dypyC+OCskN168JWDXcUVK6IXhtTFg1Bawz44M2dcRaf
S9YnmGORtvsrpQ444/ZILQc0g+9bktDkzKwXWPjtEYobQaPe4WIvOfyFm+8joESz
dFC2cjeuxZxuzKnKAFy0ED/LnYUOD7xqHf0advh/kkmuE+wF2Xueyv6yZOjDTpjd
pG9UM6ae/3lQenUZTNGORY9pZFyUTebN3Z/WhHPkxGoceRb0WLFcliE+92owzm+z
jgDnRQs74T31dpA+RyLZQN2mw2UErh3vKla9yk+5NVDwlmSP1zpLSwfMIXAmUZkS
fGBv1vGtQPr5LIXmEtcIDzkG5RLwP4/YI38EmqCJE2Vekt98q03HafgoIyHNe/k1
CJ/Hy3XZYNAN1SiFEQOKzd/mMBV8otjC3s0UmU52feigA3PeUA4KQ2f7Ux6RjOGw
DbkYzjOCTpCJQmID7NgPhyYNE3OnrbokerZgGLr4oqlE/0yOOfKtgZD9ikdpu/lV
GZGOcqh/+yuMm8XZxFxnzJ48HuMitKeLAuxiAi5TQKawflniVi7dbjIGoSkkt0D1
pGXoOUAgXPe1XebyO4B+VjtBNLdKnGfseD21YoTI8XCDt8ST+q8jD7KPQ4eM+QpA
8vRlWH3IcAE0gPjYtQ7hK3BI1nE9BUgPd7kDrpRy+KqYoZxPNjgfI39QBW8eNFoC
1Caojkg5nN8YRutfC3FgpdMZxGJ5cqp+T4Kw099JOAB59cJBP/5p+tHJkTMi8ZkE
NvgkDwScOxC7w+OYovOI5hy4yqsrc2pNwMtqf6OHK9EHs5F3myA2RcmPGROMV8Cx
25l8CieNyPHZ2UPAnpG8I2J77Ln7XZkFRMlkAgmbOH48xmtJrX23pTTObtYGBEO2
YNxQh8rYMKcSl82MdV6sbJnoebzh5bk0A+zIA7nWD5GtLFhMq1KDsR7AO3MI2TYp
D526EnfdAqz2qx+PVS1RHXOHGWgUpMc3j8+t5D/sR5pjz4kmfTC/MBHslBkqRCjd
TP1j7Rnk9BiyszAL0HIj4RY/O5MwaO9RIjuP4bLQk9Ajr4gonRT8qJqJITQ77mMY
YhL78aB2wetPV0Dvt0L+Esc+sKJoWrEOP9bfIyQKrPDHiP86H9V2ZpgXof/0SVwQ
XAnA10uTovvE//AVxfzJvG6lpMCCoByEdV4zmHnaXUx0IIi6aQwhorkCoBiX5Fpm
WM9tN/KE0AglrUbF57s/hcWYrHZQPT3qMkvW4hed1fb5hkB9Mm4M7OiYs68RzAGU
d0u6KJqi6Z3K8aU4Z8LAg4VuNi12+A5SK16qV1OAPeECOQnF8OWbfS8LV+8/qR9U
UBZdZj6l4578ZWZ0K25RxoqCUO+hKUO4j4aeJBYtk6zgO9MoHKd9yzpCJMR7DM33
AHvOQD/ht3xDLSJ4XHNcP5ZTbqi3Q6zLSgqjTMlCZkF+/Y0xFTJdctDJ9pUPHPHa
LOjpBv+sp41Gf2OxlmbaA8ktti0S9ah7ZPCyr+8oLnObxePnufZK+o73x2UdlCLP
m6gksaR+sYITMND4FT9n1CICqgWRhpwORja6khZMfUnNTwh/E/sucP+ZgUvmA5RV
0sWACDB3j8s79JznTRcdqEShMGTNZ/HG5n3Cxp+GpCmGerzTGsqeL/dkQNHwvuks
RMyQ0qcX4EHK/VkOKdouUYnYLfHoruzEJma5oUj0R19hLWrcLdRH1jKGSveiBfyG
SHILOwUNLSBoFms+/njSse72M8IS0lwZsW4oP4K9DDsuzYEsV6/HkBE8CfpKUwgv
LtfnvFARNp5lY1mpidd/hAIitBOGjiSE8+xaR06KQ5hWWmhlQ8kx7CXtmHTIe4Ha
NS8gf1tn2Jor2Sphsi2iZdVcICOGPloY5rfWH6En3veP6m9E1tgAughMw3N8KXDQ
Pkc6MB/yf6Cvc2T+Hf7g7IsS1qX135DZUnttgj+8Lu3SkbMsFsX4jeRgV7YZ3iPA
FrhJc5DegCkQAYuqn0YRDamW/GA5iALGACYoC8UDkl3qFNGhg+6zh4o/qVpmWvCE
ZJVTxruANDSvpUApu2V8QOHZ/7oC2dft54Jer6uYLts0KqKl6MY/uCuRxfsJxp90
ziUq6D/mWM1ME3wgxSjg0FqObZREPm/U6GAxAEWjiDH4M4cMsqXFkJ3VGo+Ovp1t
DQ7g2bMMBflUZICT8yGPBPfcJ3W0f1oJXfAKBbQDfVAh9sxlahTTd2xSIwoCGt8i
wvIV/CPr115txT/sAB90fZ/zaiNhQLrcjCVBOLKVNDTAMIUT5+wFBTb3RBAyp4w/
sbdlQJd+Pe7BJSsDhiGRHEFjYh88255QKQVKtseFHXlz9BqgmAVZTE6FSFKoc+8d
/uyr70CkhWVl3dRHZtDk8x4h0JsBPSSDGBgpmSI51vF5iXb2MESmrbcdz7pT86aS
BrU5dSgdHn30vTNLrJjlm+nM0vbmBuVwQsV1kjXDbWLcq6RTiCgORWi1pZz6fkaP
kVmZAVCzrw+/Y9QUkHgZNM0bBedpvFzCitdo1Q+Z7W9XsyiixdUd13RWySFPk2zB
Hye4e9SAh8vSOOpeAY6lnp5F0VjD8z2LRlTZF/9v+RPOu7WnTeA8SZev/rv+dTgF
o2of1KJ+yUqeSm2m+khtVIaWATs3OCzEnYISeghPV9xRmDv36aYM4sFcEI7FDeXT
bgKaCdqSvFUX5GF2Lagp8zVwliG6ptWrXN3ybNu7iBdoh8luEn3KiuCBRARBOFXD
RLCEJJN0YhcXpM58mX51eJh7/lwtbEJ4+J6IUDB8PIhX0fg5yi63/PAIMpbDdlkI
kadIeRRfhO+tmfWNfrwVQJPqFExi0nM9m8gtrPXBbpQpBb49M3T8scKQ0wgGJy1j
zYbKcjI9jcDSURmJAK+XK/Jry5FRQd0bzEuoH9AZb42ShRUTt6rIWW7+GMdoGo2V
GaLSkktb/HWeFre+uj8Ep4emvyc5Bebd/0q1z8nIr9c1STVxfKJ+fsDDOSuKnFdO
wOaj1jT3j9YOtCnv0r0GpfN7Eb5oAL+A5PltAEQ90o3SUbnwRcNnKt9Ru6iBluiY
0m6wRkMVjwq/DFtZf7PLQqSllGEmkqS2xdJQJT5ouUBEjDBEh8i0pIBFEolJae3/
iHIc+iLTkL5YpgCiB8miQF4g8S2N2wTjfNYyeYI4Pfb4peMWzIdLJXn5v4erSsoF
q484pcctf0Vt19alEuh+4hoWs4myPYGKTbXMWCEd64T11MVtyt0tJgUQYhYZwr9u
6g+qVJbaqaxVFL1aJkmKL4hAY9d4TcFwIC53kqgU8G09GD0pgnVXCsaiLMxhbxC+
Czol/vY8RXs7FgNSZKI0p61/nLJRZDKrJ4bGoDOdV0KUbxTBVnmyXZrpYhB+752U
rWFj+OyDrqbISkGu7RxHAuN9mY/jzMD9TakVHQ20c4HPd2jt8OHb6dgDDCgq4FND
8kQ+MJY+DvsqF+QpVzogN+NW5VMguDq/NgR+3lvPOEJcre3R35GRxnUzoJxt8zhn
yN4nIRQgxjvuNd2BO5rT/RG3tR7Ar3RVCPFbRXdLZF+ZX1lyHzBpT8igdO2iRqkC
XCHscWO7ZJyjHhtfiA8eWQWpheLprkO9UM+UBd1F6vodml9mfgUXmHm+8RnQEM4X
OfWeLJkD7ARtxSkb89bLQ5DIrXO55xI6yCfJhCFnw7obomHhnxMA+PWX/F1cQSZF
r3QOVOJj3IhB4945XUkCBymZH/GHsq3pc7eF8cDkac2VW/L7SkZaREiHWzPU56dW
Gei5ddsCiGDE9p6bB2Sna+IJHpDETbtA6JFP5GyPr3rm5Ut1UuxukftCeNQBYZ8l
d8Dzbx7UkMA/XTmvml4WnGCoZZcuAVUukVgqyDV4w3Ctj/Wn3jCZac6gX/WDnybs
XDj0nXNp5xmj6vRCt1QbqHJOD8cfn1SkHld4qyDKop/xmDWce1e2L/FzZ2aUDtTf
70x9pcBCeccO7x4x9hJ54Fnhicya8/TE694sSwdw53/ZxFLP1OiPVfT5iT4TBtKa
gp34lvlbrcxVNS5npuC6QlFtWssM2GNeGY6wi6ItK8hlIxEb8ggSk5AA4vQzna8/
jRH08ZDABhLDV9/+b/rUo0EwgG0jmXMJ8DlNzfTVHCv0Tzp5SGFFhEexap9rz6pE
hscmp1ahEVgE07g+aorGjPKfQLvIPQ4onVsJbqccA5HQr3HKpLZ/NS9NuROREvlw
emZ1LPcjOxvuxZYoQSnigzmYAZ+GZ9G1OGGYlarFzXCcS9BgKF4hYN1UtcXjJ+yQ
09lvBNHn3Eq38qvWWmcSMQ3RD5+fZ1gBf59LkO82WfCbSKsPMOwZBCQIxL65oQ2j
mE/AThV7JBUdnIHWsGicbjXU0zGBTSaVyyd3xRHfrtuMLK40PjnZFiNbHOOZnpRu
CgiJM3pF2Zx+JgxvGBTbMxUPA6HXj94A/93y8lz8TeUcYKPlta29DFiIsg5OAMCi
5x687jtUMDxz6j4CK5DcCnmFWlEjnMH946hX7hUU2asbQa+yWtzsy6FUK1Kbb2jO
cT4vBuTQ5M7yyIXkrKJsefBi/ka2o/+ZZzgzK9kh+PVpBCfmpexRjwf5Zcw4EtGy
Bap62Zjpn5V+GaYaY8FtKAn8OLq9SsyLsD2wjtPHpDv2XWSxjE+0QcS9DFm12Gkw
SWq5umBuQRkiXTSRGD0PIpC7dqTscQU6O9t++ocwTwAu5N5Mcfx7AWsfZjosn1wJ
6NCN50BOEBRT8OO/9tTcL9NWpNM/QAqyzNVd8J28cnjo06Ovc6b2ybk/uKqI1oK+
BwTOoUFA4q/adVKMK5FRFuZnw51bOxYwsLWoznFCd0cND1mrT5vKP1yDJL2yVRKM
AVxHDcy46KGFsRE7C82qRWFOZR7qv2fi2VP0EH3oVVV00cdBxGuJvmyju0SaFIib
FrgZcuc1X0LaiHxr/jlw5dfsTgKyIjJEJjOa2HZhWfstFfjsae176y5rVdgWYMvj
NWsa6pbavJl0v18BUvpVjUnmMQ+gnfgNEHqdvkhARK+BnSuFzXCO5MmG26pRzis0
ql41i8dtqw6++wOg/5LAM3qgUfKdqaByJFPGsdidjQoIRjxp4LtPfl2zIBazoaMz
OyTKFlwGOxn8rVo+PbwV4Pwjvpo1PGG9hCyCVBG8QSM5l0cORP/25B0LoeB+scdc
YhJfj1lqla0HkU0SKXzAOxv1LMa2D/FEmi0XiGA7vsXxpJvbZ3HDuQuRqdkQwYeS
e4VrwK3S8Yr1vbSObu51UTTOeetbjfiZpL58DemXX6PHsbONKO9JgbY7Wl5ixXF7
mg59HBS7HFr0DsJdtSPsS8CN6OMDKo2QXPBEJremxbKzPwrqvg2XxWb6UCxoANS1
ksLV6lc1oKIQ6Cxg9T/lz39eIlxwO9dXm0nNYpeV8qZ3bylIx2JrIpa9Xgw0UCZe
D7n58zVHCl+lr8MQ5fE7l2kECHhbOtcAGkW6bqOxKTI3DE0mDMp4K5og1KT/T8Vc
bEzc+b/2Dax6B6arKcleavM4jANK+stXjA9BvC2ONRQXSJRfwjMzcSPJAR0Q7jSR
5t6I8q/OMvJADC2CS2ygObUlEDpvHnA8GZqNGUvUK2Dp7cs2LWLHVAP4pOrAGzwk
B4vohB2CDBHTs/9gCx0SW30j095NDIw6VSeATlm34C6TrydNdwUN5iejaIoBHGAX
1ytbkUpGwhlM5G8OaqBm+pA/nmN4JRb0MkCqHbQb885lVubDXHiYHN2NblqfxGh7
F+FxqPrVNvLAaimm9BzkqCcDBxj0UcAi62z29rhz51gknc6pzFm9ToccfLD9L5sc
a4YfIByoshtfw2sEYKPUE5ZbG5ynt7N71fkE907mByAg2a/X/nxI2OlPLb1JQLbO
RkXEMjX+cwvGEUgIZPoPUfphQbGZBv9PIUcZD0IKIl2sLottn028lPvY371nf8K+
JaShbfoNBwqdt9DG1j7gxoJQrN0/N1UyAtqgYaSG0D1r7VAQjK0GKXSXewVbiMbV
OawTPGRnrGxfRqRawEZPBLtvSSVIdnAPW9mFyzcGXgEaHfzvSJPOUXAvt6H2zrTz
W9RXUWLan5WnL8e7YHbuKDvA/k59pmxwWNAbqmoBdXCSxTnNjQJedg1wL1s1xZe1
KI0WGKsSFQenJz0xzosVKQ0V+x3ALQZEYLFZHk9xhJBDYOEXAWWlG0B6PnTFAKLZ
jO1O3ykb2lSc1H7URZCI3RsASuD1iP3MplqUjePL/PZeLKJ8dSeR1d0z1uwYBVUv
PwPij4+Z9QGn1dfnHheqs+NIrSCaiCtb3P1IXCY5zP0N5mN9Dh8ZoD9i/ckho+Pl
uMEyu4BC7g2U161gmjT/EMbf9mu2PHPem9RW+Ff/XSEEl24VpWr+Uo5H95SRbI2f
LlMIFUo9I9sBhjWztQvJJz8tXUb0kD3hg7IAGF9zMAJLTM/x0UjI2+Cp/U141Cs6
HZ72MIOeUAgj1K3l+4ZFcAnzg8gKxgqBXZ7EacwoEe0YMF8uHMbqyoAYTMFAN7NA
ntkexsbHV003ZnqLpWLazi/fG0fkC9HscOG9PwCTHE+vROU8DdEXJL8xkh60n7vk
tdMzqSv2BLDsWnxnXxre9/gQTXPgjh/cZK2YKretvPJMMNgXyVla6y2vrCsSq+sb
KVaz4Jg2qZOqcPCka5FsfJ4XkxQDiRdM9uATIaQdYT2+XeIN5yW5+bI12v3+gFkw
eDv+BIE4QVU3bhVpnDdx0Pvcvx23khlAPkp/4k8EuxVQJ1xtQKdPfB8OAGVrQQAa
70bcYUrZZWEx5zHgMLZD7xn6HzOdWYCDJj1Vqtn2IXWLIX3+AmD/4C1/Qb+pND7f
MdRjPf7LP2zGN07Zsi+kq4tW3b8Sy2UFRNjGElGjuTF5CK703NEQWf6b2xfKK6Ze
OY9Q+mCRzImfoRL4W36uQdCMIq+rhxKoZS49K9tf4/oN+QhYGl7FuLKprge4RK42
eujlArX79nUYMmWjFRE9Y8sjPrcXKORJ/Ya8hhqEWhFUdMH/y4G0qS+AEOuyQ6Sk
Y/D96SdPSEkCAviQ/ezhfOgryqwx92ipGSTKebhBzEm+gqd3alDZQIaJ0xoD+Qm8
LzL6K3jGDZ+W/aBpPdLDT30qmEv/085zcji8xMx1mVt6L7JryYs4Xe2hnHhOdmwe
KM7+20MOJ+3eAxfTCgYOxlXTa3197yLCCTLG2LOai4goNNNXlNH7t76G3cLUO1h/
PlvL9NlQ2TwqEkrn/dMUoMxntfnR/yNd3RcKAnkwyvjBcBFbtNg0VakOBH3AGXgS
Qyn4wz14gGvPT97XOfz+fupgYIVsXOHY5sQN9IB+Ofol6gL2+SydlpTx4R2jDoAg
4L4xx/piUc+HfRPg1Eknxpp+oqx4HSU5yocJ0WZVIRSHBg6G4Jl7T3Yvu6FzhH6Q
GlyT2efIdeM+KHANNj8SpqwhnSKws0R/zyfdE/E97tKzaoO1VVg3nNUVgwegT0wY
NBolmyrAUOzXfLclsofTK2aw9ghPCPnbz+0rZQj2IzMwgWry9SpTczjUdfTDCPkK
+JPmabW2vMQyeXurlEHJZpkJSbmo8tUq4+kwC6hrLxN+6w1kKByRyKaW3N86iPHf
ZHklrILcNyXdQUjEFhXzO6vm3HmMqjhThORuAJvp1QVF3GWjfETcYk+zEU52U47u
/erC+U3WaSeDYnj8Qm521YVCzXCxKFy5+HPaQwN1wtc0k6fESY6990rqPKbBAE3A
rFy9PTpBA/OQmEMlghGc4o45M9V6XbnlVgOmuojmT3KHRG9lLhRKUQG0cAZ5ZVyB
gp4nYegh31j4BjjK4c5qaPl9OTxkuVGLtx1GEiV8wLernWfwAXjgnkoC06o0uM58
gv1RwdyFlRTroctzJoHiz36Fcj2JkAVTVr4jE/Ia2EpmNqk/ZfiFwBi7guizzqcg
YnBY6xA2lC9VTLgjp1EQnXdrDb7vB+/xydkEP5E+89D2DgHWhG79LzZMKv3xA6qA
ResLLfCtr+JBJCj0HZyG6q6SZN/Af48bzg4+uPTsw3NqfbSklggDRIpm1E6Ja0nm
CHZrPj4tFv5z09ER36SZMDB++M6GhasbBJ7FZXE7682aZj9g8mxTXkYTTDoCCvrx
uAqiYvLKY8ugac/aPAd2SwgpgBu6k9sYY7N8MaJY3kYh55TFpSmCqkSCCpFgUsRN
wSJdPumUTiw6c4i2T684xpXByIdPVgHfHriO0JFxTCqsvrCJJx6UoJwISnbJSh/k
wSOtsdGqivHjrlJti3uMbFhvHdgXe37sS0K71LABIL8pZmI5xpiE7XhMRYUFWili
1wJLcYYdOHaCM6NJGbyBnNQExcyiYCrmLeteDARkQXId7tT5dtoqz3UXsaaRUAQg
xfrSCIQm9FcPbk/ia3C0F1idTQtM5SWGGRm4XYhGsyqsMKdUJqQVwHp0tICdTgnG
Pl6+Z7OzNB0R2yPWgp3b5NT/f3mkKBm5xaZbkLyKe76R1d2BhDp+5G9Q+aM5nk71
Qf4cRB0ygh9BDg+XgJQH8DOlvAUi1Z3aS33WIPc2IOqkEUZXTTuflIrRPPTOrCRt
eAr4nUWLtgBF21AxoLOBDOputMHBAieyTcUVewZbGLcmGUvYIjqpk195csyoPfHt
x7et5MQVPfCuiZyxk0s43riyt/u/wffvC3zrAieIXGDIJ2tWwwC+xBMicuVeiWrO
lB9rjNVHyrCF7Ap5s4HaQSlWfPdjRjqdlRDztnyRxMaaUzJwCGY7WRX54zlErN8d
/64z/hG8jaA6aKUFaUiztprWsDRqjo8+vBzuyd9W0SVp2PVltFQwvP/wgM3wC6fS
9IivXX8jFQxpiYVVUAJKtfTRCqWeRYP7pUe6+aDDD4b1vP5kxl7hwZ1ecara/6GB
9z76SfgQgN9Uf9UisTm+HmPd7Wz5YN3p1Ftsw+vy5YrDjDouQJS5fndb20v1ACIG
dTUA+lJn/bMcyV0P9ywfA5KFCifSyemP2cGE/EWDsCHGI2Br+rVom4q2J/9qWvu/
KMPpfdAP2dgXaWSTIBpejbzpfmxVx9BL4IUNOvSfK43StCbkvEcB1EgUHIy8vZPl
1hS3Htx/0MVhLSd3iJeZHQ38tRZZ8c5Q+lnVC5X4HvGzbknuz7LMg86+L9Xf4fCJ
CMDzy6q9iwE58zqI1PEsXaT3Z65/sScv9MPWESDwUug1xsZIWkKtsJpvTBVkyjYs
1S7+0HYDB5LXAgfQ71E49Ze578PLKR3k8sq4ncA8uYvxAWd1ae84KSj5TR/W0/Cw
bLD2Wjz3kG1nNUYOspLTPB/L6UakLA1os3pUW9gpgFTAPjmlI3Q6jZmcCuFZUsRp
baebY+eJQgxBL4cj+795oB2kK0R/mTqQhmj6OV64KPekagJz+NcI5dRm6F9+JdtW
K2oKQgermoj//HzCuCfXnlNVuV2eZHKT6jEf0yhQRVCkPzBlYwywyujkuDECeh34
Mx6BCtO0KD+PFGm2Td1mm/iZ4UjSznadPciMFYrbIxLXHYcgU6fZo2ONgoBvmwvt
OvENhiVuG2U/NkGVgBV4Kn1MnexhYthQZL07IDTC5ICj3UMMSSBnHRSve7AsscT/
Imi0GObzi2U54vx6do3TOXlo7bXfKERxlp6XiAhDP2SzH6rpfob5jSME9kBozfJN
58uEqh3sWoSQro/fA19W2/uH9Lq9ghVX7+rWzs8ReFOh4BkVpx9O9j+xm9pBGLRm
LeShU385uI1FvLksD60BEKcAC5yNgEklxcnU0/3X2THKXd2tr+eyssqPJsjh8xTJ
E9m1TklvVxqZOwm9AcVNqfMh7H4UIRUv6U2XEZH1knAzDphEC2ok6j2hkmM670rR
QftxV9aHao3lIFpw3+CuikI4/q7+1Q4cNGkeSua5EoE48NKMYQMD0t71RMJvLb/v
ffHX9a+ELPggxLLtNpgtW52NFJQHaXZT1ekVBfWynsS0Q0UJC6dLftnsDMtmu0In
vi/KmGqWW+B5DABIFhN/j2FQM6SH2HXEAPiR7abUL0JTIf74JIshAd006EUa9/Rw
SVNaN7XmDZCCIdCDjAyn0X/fZkMuY26yl19Osn5oHDPkYQxLOxRdjZKgWVplD/uv
5aVlttffnGheNX8XkgviTBsA4IPQgMZrrHEL3Cr4bIYLeoqas1L9+FpLHxZ4X2Kf
yR3ig+HYfkTTyuU8hXTM5NHsIQi+A0Vk5E1yFJ4WwU80044lciBsQ40XbW40LVDo
0f+7VgfKiK9kYErdBRWrgsjQ5Ycm8vzaXRJaHxn6+UmGTOQ2KmCoqh2W/gDsG38E
+kaPXAD6D5QNGexU+f+v+y68P/HI/LB014SfNue8Ab+uKTGBTY5HyOeA46f/ifyt
VbkqWZ2EbwNldUn28n3KuCOn7oSdJnCiHUhEJuoZD4Tq2hZcEalWm7uaM7sACAsr
uTSFNyvJW8i9EGiWqMj8AOmnsVkOea3PmY0kYQx2uHdRvF96E0zORUIEnGr6+fxG
SoSscrc4NnBMYfgPKdV5NQ3F1lrC9kX9GNV1fm1T0VB13lMBgbnYeVefjX4dCr2p
YslE+VzDjZhR0bOMjcldMDZ/7WlhNgH6k5Lq/Oq+9O1KbQPQ4DqOge70WghkL+q9
11R1/HxozJ4IQjZOdVfC+EQGfxKRFMODW8KMEPxXtMv8CeLgFxHbncL4zHN6ZOPP
u7gQfwmteVkCdr9HeHvLnHqfxRFLppVZ6e1KPjWtZ1QXJxaveyrm8v3iumoTsNCB
cWaXgANpCKqKJ9cRVo5fIT2djBQYDYhPCp8fqLl4uAUgO1KGggGQMps30sSM83BE
4Se8iQJ0H+oHgtgEvp9ct+cIrlLkAgSvEqGlogR7tBTOGwCMbndzpHJ6GXOZURkl
M4oI/F+HJBgyJtnQKryMq77Gh+3z3Pc8MPuef4uNO0Uv5LP/deny0l/AK0d967p8
oUy04wM46mciQTksZ7SSTB1EdKiOw60PHzWHQRSMeTIBKG0OpK11lSJMgjLMXyKR
HkJuABIb++OUdJmRvKVveVRyCf/2SxZCNslXlP4bi5xRROW/RVZc4yoClnrfgze/
iwl+EB4u6o9KOx/pcL5mLfm4FpD/dQcW52Dqo+OdSstRELmwflIrmQ3acIEu8wQ5
2efaMAyjEsVklUU6QmFB/PLfdtGncmdmBZzahH0XD5ldA0y5mVrPJf1yFvgUAqFh
jF55vpHb5UfL8IkhmrRmSzAtYDlKi9ZnI8YO0FmyHpzPslKS2PGy474d39vpFz9Z
KAkcBtTiy03MX2m5m0JlblTPQaM4fvDzrxBhr8sk6a8NESZfe8Fm4ANX0/3MPihr
UZ4lqJipKQS7oAwwpj8XGAwDVkny3at+SsFoUDgVGCGjRKwE8++Uzd0ZL12K7xmy
4ctFvvkZUAKJo9/hrDKwlicw6KCrHUxVNtadDOIUeyndal2qQlQqbYDCJ5givD7P
K1Z4WRDTgWzLXNjAfovyhFbuV0ewaPnoWqP5PNdOuLY15OTpTAgtH5xBVTkeb4ru
NT3zhr71KnrY1K0yiRT4A4SPWry6DB+4mt6ovR3ayjP3hdlbYQwD8SC3VJxs7eUM
dTcxcH7YLWIDl6J5Og3URkBQFRxHdjy4HUhT+o0zR79FtHbGJD4sGlcdkFnJqq8o
9/uTqIKr3w/a6i4cg0+XMLvYgMOSvJBX68+oxCRFKyarvycDQCtPfF8qhtTfyllh
2/rLAN9QjaCvYcxJqTUK935tED72ZwAiMU6CHiGcwPMipImY2ODw85GvaSChZfeU
X5WubIa1npZfyg0NgbHK/LZw9T8iz9cnTsATbFudwae+XSarimPBhk0UGfnzMdRj
+Sjr5MXhC3JRKJIlaRuw5KyH0/X80DXSXLpe5NDKWTwD7BcxVh/o1qA5t82WVVEO
mkOZ51kkWWNUD3OIk/oqvFVPZhGTFOsFxwEkmgQB/WCnq9rzNyE0KtqrTeB+tZaa
6y8UdnIMUdGobpv0nvtceeXjHFdf1wm32rfEhRF/2y0mWzLs4ylsyM7qu9CuZnVE
2oUHtAHdF9/pOJECH9XCY82csmavloTANEmxqPCaeXNhtgPNH/i60c85cPvNeTjP
6kuQ06Uax4bHk6GMrzkjdRPOAdUeiTJzCNoRCNMrn0nh/QBG1xZAGxkjBoYVaG07
9n7Xfl4VnPdBwKuQ2cqcq74hV9Nm0iWWBnbZx+lcbWshyZF9YPO9sUWr5V5bqp2W
JoZua2Ll3ku2riHq8Dnp+/yHdt+tiSsbuMIXLF0u5Enm7YaX7qSBB9Xa82OgMlwV
WypvP/WuXqnZ/dxvKoAagBtgYBagJeCtrz7JzH83pY/UmDN+dYx3nEAPd5hijwqE
26xiskLvVf39F+h8ZPJ3y+hks2kjTQCcQ74re0pRlCc/M/Per4Zx487KoWzUt4ll
BCdzsC8U7vIRy1jzkz+/AjuQjNX1iRP+4pFmG4tjaCqnOljvTeDUoP2zXOs1DPqi
t7GjrSjZG4Iwp7/FKQkxbKKgtWceezBQblvJughb6Yrk4HRlKnQaGw2PutzaxLgy
/R3A7z8QrBNfhyoO2bIRfa3YRl2nFG1M3tHEwh+lRzpvNG9VkAMDPXeXBBWX9UNM
HL8lSW5MEA4VOTpdctOQQtV78ZpZOWd44+uQT3L9lGe0dv0fZAahK8VPRiOJ7ULB
AWHIQ28gGoUkpYAEt2D4IyBBd1vYcdz7MRFEXGSpWy36Gn2bwXdZjuY/A5fW/izW
ARn7ZLL8sYaa2+TwGHR0tDH5EU2Q3wNTbZ7xPNyvEcha4KP9SYqAN3xzEePH21e5
n3nJDYuIhGDSqIaxLj+UjU9N1PXPOYqjJVXMx9bgo0ige2fHfCeUso6WuScbKNz/
Sug1Brsu1zPOUotW9p5SkQsGa34XukHFsiazdTkssQ71nHRjluDnRVQxfaEl3i5+
qrKzR4F/v0xMzbZqEd8iGRXPk7qMN0X7CYwjpswNo1GLQIgvUHxJ8PedDszE83vz
n8wv6HNWu3f46/gAs0DFIYDy5TNzFRg12PFpGlfUoahtGLD0ZazqrLhlwyzzyJ4+
8NgHBJIOsFWU8bcZv2d/D+Qm1jmuTbTtPwMESxQqETcGa/CNgJZPLlXaFIK7AVjw
M6790XCpPW8apFbFRbQQtNotpA5/VWmW/hfY69xu5dxEoeWxPlb/hBBO+bgsQpcI
oXWE1qICSKg7nvJVd3mVo04osj2tCrzDgjM/vIbCnm3M9W9X9c7v7qeRA9N++Zsb
Y7Q28fFpWl0UUcoUOMoE1g/ae9lHh2ZvqMnFcAtlZxUakMdI9vc4jrqgLJU8xYpH
lBHeeghGYLSfv/R5BJKe4y62IR8uGcKxK1iBDkSijWRAsxs5AmBgmF77l/kczgMh
GqAOCWpUiD883WriowcrOCGxdeSGd3dmwbXeQrf+z7jUXEBXN+sU+3mEb8gdW/SS
g3GOzN1IKflxcG1ju+Fslcjsvn4fzOfHXqSoGScU0QccEbtENeBQhJ4mhWg3Z9Nt
uM0xf12El0yort9naJ21/usYlKzrxu3IfSKkaNCy5/QVq477l98foh12nR5iZbds
d5zQJHoDnw7tNydTJy13m5jYoC8vkQ8UpLR4CJ0fkSLyyNDKcZXn+151jEPc+2y2
1TFq9QQ8MIwSTOvZ6fgw4iAcL9Fs4CQ3sZhvbtbNanLHl1MGHRFhpeqL6n1moFBr
e1jtFeMbuRTEFvjBFhcvAizKxTfSjJBfmlEBZfdCNmtIeRxEkUwR+NuOX+DQHg8k
micSeWcau+f4i8lXLfR4VIMVnEifqx4tBxeTSyfXPPcGs5uTI2MKB6ZWLfMyfGMK
91wNarC+4Aa0AeJdqqrUlXfyr+g7dgGVsa/6ZjjtXLqdFub2UeYbVUXsD/zVFmAP
0ydK2ZWYLvxsqkZZSdiKoeIMFOzpHOOMdaDw5i7R9B5ip4cQd50qi5GpxiHn++JR
r1VoZwa7kg5SQj4GG/5yiaGbG13ylM6Qv0fks9aXF1KktdSPvOiyoXcbv6ckJk9R
sg/A33Y630atbOgwToCnFvWVbvYsH2waVwq1w09yPJ2A+3zRTc3ZmJOS1ka7RedK
d8Q7aQH9OvL4Sx4ybkBIP7zxv0XWs8FWRLo8SFrJthGXxPdzMJQ1BbFq46AKk0Ja
2ych4gKf7kdh/IrB/pblCNvSTM0ixgq5Ef1R/OwoSC71Qf9d1AEs6jws3MFmaWDn
p8vNLKf/YH2HSIgzOvtVLenlcHsgZtOlzAifZeA0IS2quUhLlb8rXphYXUUALPBo
pf5z+PkKmOFPZ5rDXlHpXabZhkyURZysiPvAdYWDynnqcNX+dQinmiZX+5T3p6MC
yrNuU91fMS6Yow2bljyOKNOvFttvRM+RWTF6pvkFpCeme06jWmvpJj5bOnAZPkjU
axBhgUma5JBRF+Pw+CXp+jRWLe2W3mPY6knFcW9Yf/UUYK/ohzzDQ5YgvqtKxF4p
ym26/+IyMp4YVJEQbzzcgvUKce8WRDLtVWZd+N3+kqx+KLTxd41SfqA7+96IdIBx
YM6rkcMgedG0r1bd248oLCDgLwMelLZJwmyL+Fv5csvWF98IabOCstPNNVo8NaP6
1ki0oRm64jb1wZFGUfZrgKYmC+chaYSxt2vjgXhilM2FUhF7Yn4YhSvuBexF/NLF
jVUdydVfStyYyEA+wCBwpVsOjO05w7VPtBVxWRGL7UYxW36plIvoXibbxkr9KHQB
ddCUJ0loZ+QrN8yttjccofgq7wWKsJ+6mcDmQnW7qieuBgjAbwb1pnEEC1QkY18G
5dBIbQYtoeR80eOo6tDbZll3PusiVpCZDIliBVRh3aAim7fN0wTCNX0hu2g1ZSVd
+mJVu08ZoAB7FLvSSnCAtN7i/QOPOvaZuIbziVrlsx+e4ioofpy8XKe3LV0bonVP
qlh0ufnAAhiqMJ0tN51vXAzcR7h6qecKp4mE+ue+15zI+VsJ9zY/437TmegkNhOL
SUee1g5T+RVnsHtQ3n2OrDPLBj34CUTo6WwMceT+U/C3eWmvCYAC+x5vecsb4C1n
hJ+XZtfCFp36KNcHhDqXMejsJxFif8kQP+URtxpQkY4YBnqs9TQI4wpf9aAqXS8W
PXI5QDwAHMq+QpCuFHetCK90/ruqJZiDcVZVJcF9ghfJX6fcDvtUA8Wne4OwaLQO
oIzZD7vMB93HXH/McrmzxE1agHZ0afaLsHnTwMcy+tdC6Om36gByvDRzVdN3ebfl
2APhojw1JXEjFwy/9kJMEls5meaQ+XX7lW4UYZzRbsXkbmCl+B4TiV2zDnr50fBZ
R+H9NCUDu1PBl8VbGlzT2sEmSGbRP6W1GUnyrNfy0zjglnjlNj/wJtPWbG5AXEub
ig3O86IvikIsRq0ooC5hqhjEC80iivd3ZmZ2tjLfdOiBOdlLsXSN6hvSmNMJY6E8
yjJ5Xev0oGmPchq4Ewm3BaPuzRkg0c4Ab4ElbeVdfzZHLOhcjclbq2z4GQgTp4L3
bcjQQ3wKxScG0YC4fD35uy7oeV3mz52NcefIqPQekjsbEj97R0+g1qZgNc5AFhtm
jHPKZY54TXe/JM2SxXoC7G/bhBSrrwZTRoVVotBh1yeZ1elGCkPTnlznGZO7k3AI
RqEhdEPOtIZoPmThpkw5jf5yCbWx2RXeW6bVZ1dImfc9757vZb/Ne7F5s6DWaD7i
JcwNXxM+bIxG5eOLdR6eLvcm4LGidUO48u4aMT5P/Ythzqk1VJW7kk+2ap08skIl
iDzz5pe7nOrBCCAdXeJzG+ahv6agpyxmtWdb36lni5glrYvft6lfRUZFV1IzOCNJ
tmFT4qtjwiPXP7dzDwNvh5G2VEbqXYbj2O4nfpauyJvgGH0zKs1/U+VXJvAI/YYG
s7Th0QHWpxGJWny5VW5avM3zrJROCe0nG42TCb2cmXBHAIn+4dRKypgrKQyytzMB
ZjKm+Ck1qWH7YNHU4660NPkGPzA6Cs5Zu/RLDC3cnEyLU0v7d8cILS7bQyKmCq8m
48TlSjHvxq1pgsaBLGqBHjb2JY4U7bvd4fNNCBSxRG0u2DIYkgStMVMHwyZNTFEU
6IMG4fIp0MMFqWoJslyWZuYucXqHLGshNIkI/1wqVg0f3sCDmMkUPz+Rx5xH7Y53
/7ZdKhHwuL2zruIDV+cV9vSh2Nf39BKp2Smhip9PX9DNDHmCvCGHZ/SzQ/VRDJ4D
HzsPqg3ZIWNNg1PJOPlkpJyzH3oJRfXhfyxFjok8/SAZz6tqWHgPmyqemdIohzCe
zrppzpkLSBzRv7UuSoRmpw+19DqmY46fWx+bssGCuCOx9xpY5gCiTxjA5tkiRZ0m
dhokRq+CKQvvL2ZTHOQxS+RxBkAbegAEfeK/7L7hhrqqD3ZCUypzyRV0QTiDdhsO
trbNpi25dcoRq27EUbS8S2KzWnH8N3DkHF1fUzgnZuEWT7gkw6E7PvUyRt1wAwZT
iwbA6Glg//CfxPBFxwyOWFlU91L36Bmo3q6SEekuhnWjMEYjdUnRxnPNbCvVwj3B
JPk8+xSkVcEvOh2e2l3xPE1yBptsXKFeK0bEvN/bkQKSLb53nCOW/c+vWNIFnhGq
KAYScqqRFX6cfYlRpPb3CdxQj2YWJDqhpWpDS3lE07cefwNEL8o/A1fdUlTACOj7
xaezDMRyXEZ1OK+H8CQJUqVta3EGTJa3GMxKX7n0rJ6kubZaxL/78AM3svwcCo4B
F6tEcexlaj+Ap7S1kBy8WwGyyLpg5OwttzU28OObX/AtzKY4GdfmQzNMPbXAG9we
2uwqnt49NkYN8N5kN9AkfPjsBDsxsBmoXbJwwZwexIXtlJh+k+B3eUjXT5nvXifz
PYIhFE4+TyJro1XmMP4aMku5SIz5M1tuXFdnNksyY47hNyf80UAQWr8fKAY7Iht3
Zz9g8Jco9bX2y8isYOxp89cxczwd6zOlaigB2kH/9srPYi+fsFELVkNj3lgeaB0X
U9Ll4sajdQIqbpkC6TOOR/jXVKMaYX3AsD/06g1LTISK3LEXJGv+ACyUnqk2DrKB
pyQnEMr0hPUXoobsAq4MGPwMhmle2Z/4jB2TMw+dHuZIMl68a6mLWYpJQxdL8s0p
zHeS+IAB8D+kpx39Ys/HPaDaUoCp2qKqOAw5SHCXLsT1mAxwFG2cV5YKp2UmC28t
WMbj34s5xw87oY6ifZygAEWLSTKyjkRdP/ZwhkeZT6RtUDS17XQnRw8tcC/xtye7
E7kgWNShWlxzROJc0hP8dn6dUSCAFc/J5Vn9qmNryXnNKx575FKZuPzp8lVEj06x
3BtxSYGOhfiBYNlHMaZxv+BTOiAhVS4TuJthlUKENa7pS8X0EDQrvie3Pdq0xTD4
PbkeKSlvV4PtJZwKgn0yTUQsGPUcPYDEmMrl3+OyY2Ga4aEDd8+at5wJvo+WOnOA
GBJEwpUpwgeecEq+xPZG7pUb5EvJo982BiAr7cNV+AGCM5y4qnh73/huIvs1bD+Z
xt2wRpbSN5U4u7aGFRAsZiG+15zx2ZaJ2tgDoXHqKWiKGDuD3sAtpNwtd4+wZcuC
hh1+jdvba9JtsCnN4rFCfchI10AHc7rN7gQmMn/1DWORPWGWWf/VB7WqR8TrV67/
FHT8Q3SuXtnRNJhT/J0K1Sc1XVga+sxYHSrmpz7JG/KlMkoTvYSf5bLyO1OCKXx7
dfVChYn2t7V+hjUsXOIUIG/TuD5bKZHwJo8W0c7xTGsugmiARwtbLt7i88p70P/r
zAhpQGUh2dKrjVsyakUKcKGBrCU+EuUNafWVQGAGFpdSeP2Zwl0KGVn8S5yu2ayt
FZ1eLX1aUC6u3cyHjqVMZ/6Y1lRmjXZ5G3rdgxS7kdrrRxP7OiFk/pylRABKPQme
FiIu5Uvc6GPJ+m7qP0R5NE5M8t0UQGBQ9eFxTEM6pNZ1xzIGzDLKct4f6p0v9DTZ
yFgn7AY1zIsFl3tYqX6AGfObeudOa9go0yi9dwlJWzKt+2a7z7jTOtVXt6mSQTT9
fkHxFZ5pnMLcvbMUvOBN7OnjHgnwV23XU7WXmqv0XlWesrImJkGoZkXZ07utNqKL
LZm72gymaD/Y6j1L7ZYdhahSon8hU2nWQbXd4OJjAN5zqdZTGh9/QP21xaQl9+se
0I0LVNBB0oKjXYQaby3KmyHRxGJvw4U16X0RMd+JlLw0nQnvSHfVAqJMHqs9GOlU
MMJaOZyc7JBDaY1Dg8rv5i1AU2dyOVRVYype7MdnHcGULC1PpvcFtMpktBba5WF1
Qo8f2EPoABUrKibh4mYHTQKZT0Y9uK25a8SiS6C3yqCD11Uq9RrMf9F4esJol2X5
wHOSXAVEAzqJxd7YrchEFTrtYPIm+tntVUufC8Og2O/CSYA+BxvGR5fGd+6MjQGh
/E8makQ9X+LGNyO9eHEuzaM8cbXJvZ5mB3fw8C5Jjlhgi7xrdyyO4vZ9ZcvOpvue
GGm19I2NBz4KHQwU+ioh1XbNEsfOq/+MgzUH6BQdSKITNjXTeqoytGmWQ+scsqqU
dkitOMmXtKBXpSdNXIwSdLu2HF/4TPVNyWl9Zfd5yHzS+sDAnV7ItF9i8hBJTIrX
++CngL9y+DAyjAJXMfID5UJEsyajvkpzzPuf87qrNzgJ9AS2nZP9x5c7K1RkOo6T
NIt3wKFZC2ujiCORgYyARxksZwcj6DbjKBJL7YF71KDDIN25hqBwmquvm9Al8Q/Y
SSccyCBzunmdTjJsr46bw3j7JoHxQS0TyQdzE1lQO6XtatmyBXra5Os8R4jT2y1I
xCyhQ9Lu4OailY/iOO6A9XHXKyo+zjWsw8+h6JRHeoWuJKSTHBvPgJYfO9UzAdVF
2OPJFsGfeAE0sGnf0gCsrPNHAY8hOMHB33bkRWpNhdZyOBR7q42F3iYVPnf5tVuT
4U36cL1N2lQar3qlHc5XEA7lLo0YA0AVi/8E1G9cjYdh2TFjpV5S55M0uAf1EVBN
TIanVCESKC56ac5NRzaXItIQyEf9MDoQJim+njMEmHPx/FpEjNcVaGuA90AymPGC
42UzirRvO/lMvpRnBCVwGhhRpk58xfRqMm0aCVPsPHdrsQt2EjFpmToWc6rXFB0w
1+6dJWlK71QgBpVV2DKHIPpUl8nF9tjG5U60DC6J6yLaiUBYLJsoloP78vg2yohm
ksQggM9gjxDh7o6MJv6BHUQ1gxHZ8e5u0IHtjcv9taD+ovPCxa59EgkdZYeXTxuM
KPQtY3d8ZK2V6WXJMBmyOml3VhRpXnuj+QNm6yzw6VZbgKM0LeDmO/7RC/uHMH4u
npKCWnnAu5Be4IR8yAJhh0rsR7/7xwygcr522USWqSUZxIDBVk5aXi+ooW8aiQeU
fd/c0couPL5OcYybp3NO4bLWbwDVqDtibdGV1xfgi+hh6C2I9+BKJuz58ktWg3Fm
4jrzbandV/+vubCoZOjS4MgR5au+pzCd0OnF1N55JmFYJs3j2TUzArcyeqDUjZ4L
sVjP64V+fav5JGkybr22FmbczcscDdCigorncqTycJXVkrCOeYa8lAw2vLGhWo3n
i1Kaltp6TV9fTD/8Sok1PYO01l+ygZqydI3lCo2ssk2wFOB7MpsAyTELv+7UO5Gr
APEeq2ZxfTQsqDFQA/koBUw92cvwivABMn5E+mI00RniIPryPfAXr1FZ4CRDqRGC
E3dRHcPCCuSsgbO7g0/28a4eiKBow+RI1IzUC5NnkDroyPOx0nKYDGYVU5+u4jpW
7ETNUwxPrg47ubRWwKOBBdDbLfx9Lq/HVK/PN/RoRMw1R0GnShhXLMgQmikwEAXi
10sPHPcBd2vHpFf9FAlCCa1OAWMF/KwjFQ/kF8ueh783B+NFmSNB7AEdmx74sKUQ
rWV0P48r9J+iA7+/rLgR5WqsLMnkiQyp1MAG7+HUUve8O8CWtkYGtadm2I8SjxVU
gwTfypdcp7I3wxWUVjem+fAh6x2aFd735sRixJwpPz2CMgfKUP2U+8q3QWfkx4+H
5enRbBQfnlk69y5faW2p1BjGJVAHb3bxviNrujux9WB5I0JavQkBKyKrRM/h5x36
O/l9X1laQyvFOWhg0X4Y206SPldxtUD5P8rAYGHV6Hwfmmt/6xxHfScDzwyB4GU9
HQhNWc5GMnaEceQ4ZPd28C/jebf0wmem0bvUbVrUzw+UiZL06RZnJYz4ALKi9dBF
i1TaR7D6z0CfLqZthODuHhtYVC4gm3zIGA9WhtfFHao1MtIDiPoMorHZs+F7YJzJ
dJhx4IHIwyS+rzmwuFFDAUKv+8m3mcj4TIX1yVcVMSUdZajCe09HTe8RQ5LGAFoc
DSvyT3zaCGBgUN71vuk+pueLQVdyMZ/pWYuEIrmiqXxK+JcTttQxCLpLk7xZtu+i
32cBVuKXTSXVeQkIGWJGSDvmjuLcbyCGyJWCqvrsDMrFhdar53rfc9rrlaDNJk4R
/k9XvdyFP/hWaU41cBk71AIPexXNDFg8W5JCEnt6ZOg8QiI2IPE6QP7HoX1oaylY
S1pVLq6aW0PQjWO7fxb9LpjK243/3uCeD7K5DjZftzvOBmHO28WMRcLNLQoVHwoC
Ot1K7GX7ltd53oQPzgFJr7LY9okgLu9GgE5Sox1pGGhIX7f05Y8e4pcXoiaHMfMD
qK3Vlw2cCGt/W1Q67Y6YCjVUY255xJK/NOKFhtRoxtSLEQJdYjhUZ9dJQCAeKTDy
6HN2jKpZQRTBmi4tBLnD0C3jmrZ3mFs2QI/GMM829T1F5KtvrAbR0wsFi2UAt0uV
I+RfKhGkw9+J8Wv+BBLXpVyIpESUhhulMFVdmNPO4/qs+xw3m+psSHSfJ0+BpoYe
RaJU9yo/V+6NIBkgtIT/f2gef8BC1+oIf2XGWeCHmzdDhxeSVVtykAsC+DIYKrj4
tQwM6ABzFK/QqwMyuHsJeSDB4CY3MoYRtHABHFPhTdr8L6reUMdQDX9lcz/ifEAg
3VAmGiawClVt6D7cgd+MZy7h0AGXL8t+DDDp8BeIU6/04bzEcCpfosB+deLukifY
cCHnJgh39xS6eJNxS+vYs/I8WWJiBj5SbHG8j8300jhwS4ZUJwT+7mFcBQA1kGwd
5G7gEPIU6hIOm1GXsd63fiU8m5lsrQqgjeNnw0gUpFPjvEHTxxi9ufsArQZXJ4cm
eylWvRKuckjuLmQGNZT74TczyIc/ezAM/7tKx0Rhd3zeqyG3WkH9Ib4pVY/y5Jsl
kn3ig9AaMbWG5h2kGecyP3QZQEBYVDe3bigmY+I9j8eJXUjNOTuLWTUEG71Y5Hw4
Ib/iOAH+ZcI8V0+jJ2z2VWtLwsO9EdhtLBXHOL0qTT9t7S76Xy1YEJ1r/fzSDwV/
WADmCf4XlCX+8z88BPc+dLPuXzX5xUD8WhTl6+WNxEgKd4rXk8WkFVv7+/aOONgQ
gEWzbpuVJ8q6sh/QujdLWz141s/zg5VR68GADfVXERwa0DxjjjsGTZErjhiwFzOA
JNkFd0tBx7UReMRDLiihV4wfZ37FJ7D9wOA5YkJrtJD1M53xaMi+t6TaKxkQEUmQ
lOnTNAtLC5X8JZtQH6rSjCnhSUdTjZyJBKPpILBBZwDzhRsneQMAEWLs5Ck+QvNz
oy9nLiWyxckI6X+CidBvDH+FdkQB5BMLqmV+qv0YYlWpkSCT8/hOK1mgC30OCBOg
h+utS1GPEAX48nb8OhVta2fkD6t53Z20+TeapgXDxOFbyTLupMn1eZaxyzVXImQ5
Qikc8daNf21higughUY+LamAqfI+86jlNS5VBBKMnsGIboBxWF8ZQl3g5dsEQOtD
mz0ND5gWN6ycbAlkQo0jHGCFzstwWWK05QnPZ9bht22pICPereV97PN0uyzr+S7/
3CCCuoKIGAJmrXW5hPEE+lxoSWH2IVeGiCQ6OSgUoLoStcD5smgpu6l71BvqcMAq
gEEfpK1/n34D6o+TPxw4kmv1OzBG65R03YwO9hU1dwNZjSZYJAyI/gFR1FBDIOa5
wERHdU/TzL2777ew2/MAw/J2kgXCcoAAndK/Zh+qAwsSD9j4geIa6OQ2wlQLw9RE
IYGi4hMv4Jm+zVIZkt/O8tgI9N29QR1z9pvTP1Rpd9oDRnZKhy4J2FAMAa+lgueD
LU1z9iczHaWMHFXTDdM04Tz29U21DRomCvhoX/+xOKoC38n4J6GL++VNQB2G0JV9
YUIw6H4/X6P4BpM+G0OSeajLKf59GKerdvlZxIh+y3vx58j89DkjaPHq+rU2eEpt
TY2aKoCFHzLXqEjllCMVYXF7Ey8LMUssJ3QCAItGKArG2KUYOOITHyLYLZ5KCk1g
i+DiOwKb6c5jV41huyPstASKu05UA7wpBIBV3ZuaKNwZrQlabS11yXAyobEHYUYJ
hqo4X1oTgeRz6zta0lsUV0TdA6YujHiW8cP8l9CveFm/sMpw98+Eaaanl1IlDhKM
ydpubAjc8FpS3m3/x07Q9QVOGWsSZHn19JE/IlBS2QhZoIbPr/X3aYiHoyb0hhCq
Y1WyRi7A9f3R8LPCNa5AGciAhtuZEv+4lpRaaA15uRz7mN6pUEtmPaM/XP+v4tL6
njd1A9hTdJoC4QfMV1DwAWgRDTVK/KZoR4z9Bk06l10hJgvvk4l2t9c/l35xNgqQ
k8e5aMjaQ6t8JgRQiFz3DY7bTbLLCBsBr4MIMb9rMIp3mHyiv3H03cSboQS27uag
A67B6D//U24I0VjBQ2T4gkm36NN2n/pqBC+3meBz8Pf6sml0dAfFBbRaRFJHh8ps
1CBFZp9Ztz45PfZsuzVVcK8oVxMJUFDd1cGLG+6LHXQ1Ch4r41wdujGWRFrvM10l
T2JYXpFB4n+9paCMYlzaiYsNJoejBmYebUXc1H53fJ+7wwl1bCp+8rxFFcTR+TfX
sWALfOLOMaFanbuQt/2hN74vx0STceiNJgKVCiDal0vLy9WCbhm6DWkya69BX8se
WTfKFdkmZwbFIYmKFsj/nu6CdugTTIDx9s7Rhm+4UlX/gfuPPkkIhl98C3jlZTyk
dfD8CZ+pQxmjB3Ba/sc0l1JgT/o7IvA9e7rOrosHt5Gftg6uCo90bnWKKOvMdcD9
XdfUixQur+vMDnnsfIJ6RsMHpXEsY/mA0nBbLFB0dhT18LHk/14LH7jCb7DAlIOV
nfaXCl1CqCCBPCY3MBhgSyMkLs0Chy9ILGV3ZkXIMbjyuhvClVmmLvk1rT4kJVRa
AsLh69ZiZhjshOQywHRt5YxSBKXuktAxg/e2rk7fJDyHE9CazdlLvd3ajATKaBH6
GYADLEtSR23BGPAOK9mzFgruMPETE1XRJwvD9OT9sZ6/6RaMEsq/BCgJEfxkLtV8
yArRMgUGg6bvB+FgWknSX3IFL1HoUvI9/nQGkeaFORR3aLBhUSvGhc4baaKLAQky
8DN0xvNOnwUVmV3PzRiJimg/v4H3lMwZOZZN9rPWvAvpLOtkxNFmIOWon+k1sriN
d+7ua/XLKCjUEjniD5wjvjuZq4EZdYIEU5cWZc465B0nUdyn7t19K5ipe96clO+/
ZPHV/2CDZmzFzGpRpJNxgKbz8c2lu3HHGgZ2Gcm10tbWDO8X/hyloIjV9GOIln4y
1eRBDuLOU67kSLZ5WE/0J/b3wFZaFS120J/AM5gRBlKPAeVK+TZyN840UCIe6Tgj
Oc3/QG6nT3BGoXUJE73x63XTDwFmCgjZWI88IY3BxgRf+tsMS+SdbdkoRnGaCYvy
0NpIFgP7fbG1lH+D1IvSOi40QvjYqY8Mbx83X4nhcP4iUfGTojIeLiS6bnU5MkLX
yLxCrkReKWMhgqrfY23XKNsJUNpzktEilWZQHF4C2/4oPZQB1vPddmrRLPu4QNuH
+gZoR5tRoA+qgRorJIUQEmUsToATU3OfMGoslinNQellNnJvLMMB8/ii+xcZHvEh
PMnUGM05Mjl0ZpJd/ckkOn8AZq3fN/hjR+lFpbFdE3h1G0KOJKBNHuErsQJxrcsa
a+fykWDBxm4jdL0QiPYmBZumnS1WG8UL7ciuNiN1DTs2ThFYBhvFGw15aKBrneJu
2TTkI1E/v8kNfn48yaSOWgpWz96VJg9YfuotiYhayq2BJZ1VjoE8rzv3g7Y0sYfp
rcHIR3Y/MlQBJGLre9t4Js1mjHpzkq02Nq+BhPlN2Bm+mssafTNasejEhwzdsa28
yOsJx5Z/4h3wLSXZDb/j9Wy6jpNnS8opqs/X64jgCj+DXQuLx6ny7WrJdI+0pXW1
+yuKsxBeWTmbLFURHFv/5A31z3mejS51QwYk4EbndZ3BUB6gBjaFtCBkba45MBqp
/aYeuxn2nVNaT5XyZqpz6XgzzJQNj3kqC/Zscp80M3AJnsniRdfoNFIH4xuhEIHZ
B7C/eRdokfL152TnHm5GFIpKYa0fW2L8SNqD1lM2bFRfI1U3gqUR2pIPSznKdzC1
wjB8GgAFjGJ4DT4pLU122tEzl+p+S/NL32xMjt3wAWKbimUJZlOFRbwQA5i1hNuf
KExyMYKL71zSu3e4WR836yUeK7CTkn7lpCwtXeggK3EKpPC/IEDBWiZRlKGy3/L4
1+j2CIAHrarNtKD15vmHw4gcbhg21FQ6MYSU1FoAl4ki+Q3pt0Kb5zUWYtdYDVUN
VsHOf3hhJc8TYOF/w/KlhVx6XndUxuVZo4Lu1BkIxp/wTgSoSP38hQWMqUNYc4p+
t74QyOQ8ftkmUWMLC9Z1HGCm6Y5a7kcoNp1aIj3woXlv27yyv3S4gtjxUbG3gbuo
D4LOL+I24epr5Z7rfbGXv7WEFP9LegLvJYLaDAZ5ePfXgsl0E4gUhItnX0Jfq/3b
fHRjVURcMxSJH3rT6Avb+T4hpC+2FdWtpvvBh8bB1twBX7t9Ge07DwWtvki0PqG4
HlPwjdinZKxJp+k1Xdq8dWn48D8iUMYOu9F65AGvvuP1hZvela24WaDahMLsOBDb
h2BGrsOzRPG6GYdmQQpJDLFBkYiOBeccD/K2wcpWlBc2+/dGNA8FRjKgC7aENMU3
+oenbwbayEVr9oF7Uhg6RviiLpKUrGilQpFHGcD2+FFtgp5PhjHERfU0cSgQF3ZU
GDw7q5NAlP5DB6sM/f2Zt3cYTErOUCXhdtk7K561zed2spl0dOXrr5/CLlz6grrA
jTlzfFaJ/ek+zY7l2nPvmSch/yObGXiHDsKjuSYw5bMpMpptMME6yfrjPhfpONsb
hNnyj3gm5OytFNSsyA5qRQ2MRRvBaJyDgQwkw45zzjS40luKOZlgFkJt+qDO+Jmd
WRPoVBD0PFjv7JrTMujNmBOyY3ipkL2RqikZmR9t3IfadBoqAnTBAqw0dQ5duust
suLBltZ/z2KwQquBWTENwsR9lAUMNJkiO/QtD8iXzG7CSoepF2eXb9DX7YmbP89O
YFXlX0bWLw22sf8wj0POG81m0KqSXZyAkCGvA8ZsHXNRBO1M3jKqKA5XVCz8MO5P
o5bPW+P1TjEHD1xhf/u/53+j6pfpsy443cvkz9Y5oTJsV3A59y5TgelaUKMkc7PO
cJtJAC+yeIC2yoE9rGRfu0VJOHPCx8XCyaZZArxOqQoN2hh1+2mdspGACKUqb6Tk
T7CBxyZMqdmI9EjYbHKpYAK9wL5DOesjJWRVtABwDvI8rpvRhc0r+HgSENMYi07P
iQRpapF/SwWEk0fgx7GKSznHkjXCoeHY6DMZY/4zvFUArifJPPS1D70gM6/lAm0d
l6M9ZFJv3HA42k5JFhaAbg3D8bzrot5jrYHyNEvm/x6J7dwwsHf7SeLynhvgw6we
qvjRHLrjvqMwEbi7EbwsUHeTNnznJ27AD3A0DwIPl1t+1H5EAAeCUAvvSJTx+EEM
t/flCpqE5WtN5vPqj1bA1KCRmad9C6j62Kna0pjcXRxd/LSjM5MEdi7eN0nYOE6K
xpst5sAgTw7s4nTYaW/SkzyzfWX+HPLMpTl6A4OXLl6CXqYvqSdQCdiKazhL8w/q
BbpkbZ8dvH85MnlNH9J8APZ0BuG7SL5DX01+WWp1byM5eBIFPOk5MRGvZ4ZQCy9V
sMzSN+ylHtg/fkqSi8vbb8FpuzGf+7OOmbpsRXZLiKAe7HEnahfPonbqXJzp/R/q
NQbDA1kKuvgBAfGgxryJyRk/n2ojmxmdfYcvt84vNDB2/5p9iJ6xxnTwP/PWxtt/
7dlVXnAvdcNgYXf9Z/uxSzSII7P03wfXVQ6YtlUapFSKmk5A+Area1bAesoIg6TB
Cw9ANPBXV/cklrlHT6j5P9Hg2+favdQ4y3o9Pw8Y+DRKTH04LW56/A8gYAbNrgbz
twMDSedph3HgomZ172PFUH/3vZ38bydjEDOhzz/vh9Px5TUMoyq/CoQUGB/PmNIs
bVL+TBb02ZrozcQnLtCfj3gvJameif8oBSckwh42FejFdbIaWBrTW0lpAmacbErT
v2USNCF7vF/xU2PHJHUfeuscnC8wsbU8Du5dkvPFF1abPQM7HyqGLAgK96Zrbf4V
Hxb0o1Kae1dBIbiuUG+qyYHPLY7beaO/YwWkHMaUUoUebf04DZuo9ZLhMWG+Ovg6
ENQ5qE2ZU+VHK5HzyRi62IEWL4kfEYxeo1PLu5eGql8su8t7kl9bH9IeLNN8RKVe
sOopgc+J+q7hwJJ2qXQ0agPp9SA7ejaFmXLaMpsMD+UBneDGDWwS3DrDI4F5/Ygy
gGRTKqIx5f23O1s2GfGMPd6gFELXCLE0gAbqWwopRCAqK5sQBizqs96TEzXd+cJz
h2LU7539GO2remwWpZ6rNANSiQmuxlUNiT/ocS8EhLS/QIqkcXMkKUcvETaIiYQm
xdAo4hPyx2da8rByEB0dpl+Et6urZ4iQBSN8UeoFqsGEjflTBTuvNJiWuwFHwpax
4m9hvsHbzKfDN1any/UkWJsxhnxgk81MfpkqLlrhauX/golpSCtxKgn79eOmDrBf
Iz1YQSW/7Z6spzo3YGcsa3mrWO8TZojJYAWR8gK/LA0loQCXXiCccjjuiYK3ZXxH
wJR9cdMYvcVWqssYAqVPMOggdy961eXhOymcsCHyA94OLBuL2MpvUhHE0qKLQDcL
bitylN2ZuAuLYmwQIEB6u9I9ZMboeZnDoKbiC4RphzGFj54ylVnnWt2FtBgLgHQB
+iotUBIGTgiWF9heqsbhG7kYbtifOYwUO/iIN9Gc+UnZCCbB31Sxs7pWudsnywpS
7r6vJFewT9Tsu0D2/uSIm3ltEtDxLUARAU3UkdEv4r4QnSbQkkDaWgt7rLlqZ9lC
I2TRROMZqtxnqOJvHMg9/H6xUbuuTEE4GPraLemoJeP3xn5S+mTNH7e3It/e6qCU
5KdoG1ECSkZ/2xJy7dWvjsWls8W2UQDTsVL0QAipQgTEldg/koSaRNA6lKoBGj8h
92EzryVCMm8WfHq23TFfiGJ8wIWA8E+8YpWm2d0l1p4SjREftWTVdRlXyA6MA8tw
cRmc5iyFj9aLuLM0k6Giqvl8YYt9DbItiQdWQbSZKol0w2tfxQ7gJrEifNYNiLjr
kDih2HvUOt3jwnXtyKFS1a5FecFYT/0bUPKWToMkzxaeoQv1/VBk/K+rzlF+rk/3
/2Z9q3SJa1DYWu+NE8LRZLK6jSM1M0Hf89P5RlxlYUmuhY53QXxuymFk7bjBFcgc
Z+Njg3essZIJBclxciO94VkBxIZBULJh2s7THdYDzMmO1zq+YrHY9Io5MBg477KV
6Nnf26M9SEfAZ3FIDCobg3nYUUUjfmO6vGLJ/rAE3W2T/tjWpN/+0bVcS4Sneztu
4ut1OAU3WbyK3FZM5nh4Ff2DTWIHiOS9fZypI7FeL1rWC2V5eDDB+kPy4Q5DmbdX
jIyp5BenwM3NrueyRGDOUqsdmivpPlQjoOclY/fh1HTfllPt7e6dQQqltHm3B0gS
DuRK3oAsMkPcX4wIePO5V1ATsUBuKM7g9Yj2YN0l1JVYTo3vr2r46+6EvBhMaumo
QfcrRdlB8n19Vlz3xaL89z2GSOrc2GkyrCfGL5RD8qTkz+M+5OHfX0yt8rcXSQQ7
/+Gbnf8N2Lt1GPQvsWnoMWS42Z4AezpD0DLmDeS3yo36kf4WA5+HIo0Y9WLRTJhK
rQgz/dcumLuoVkpfBkFsAPk2N/6h/j4KzfO98+ssBrGm65emuT+cWksjmXsIT9PU
Bd56+slJtTyRT3n/78MlCXKlpYHuOW6Z2mKJEuj3stFLUgOCL8n9yX6np1PEavtC
uu18Qx0Dx8Y54uxB6lEt/a4UCEap+7NVhFv0XNgSTwspCC7QDCv5LZD/efpPhonA
pbxXpJWFUIasbrt3w7zQBuqolsDSgwdqaqJljXg/n/QH42sIH3/zRE8z6Pehm3cU
fVswN3GaQ/6W2hS3IN3vVWkFQstaNKKMljPq08IScqc7QFzJUxJB75ApEe0SWXya
RKQbc4nd6nopM5khcHMms3MPkMNCOkLw9QIe3Slbz8DD9HnJIQD3AU8tJdpw3DCE
aFUrhehzAdvUfChVKGPJsBIHNFdufBpfvPJb6/nn22QhyaYjYHWQ31fu9niivPqd
hpAWXdTIX3Co44bbQoZkDIrX1zauKJjh4c3QxPeD0WQjrV+HNcoSswzmOD2O9isu
qibWKXU+F9YGFGf38RPVhCLP2XGkMRITyJZ6S8yUDpImh39y47dMA5vLsV5+NMH4
fAKcEmxJrrNht08VaVdMoXeixeb3v/2+ZijoB63xn6emnoOwkNGuS0TB5ywMbCQ+
iCN86hVUQtwthhp8hsHJ7vUWEeRz4B2D134Rd71ter7Vdo1P1qxxqWu/V2lkQ4Bb
X27NkhcGBwtpoJWpmaYNM4WdexPyUZd0SpiGqrSvLn4u3vOGjGMqeLNAYGTg+YqI
VcT4JNCY82vYK/fCQ9WrFfYcWzcEr11rZyIK/eVSDfs2oO+TFpIQgkXZiagdjMfX
pcSSP/mDNpNLNItMgIegRLtGYFK/uqBNZ1ptAX4chWSsMHjqN541xUyGTUu2x6jm
RYqH8MNfkOOnfXFnCdrqfyqfRSs+QTjPKU1Ch0EsBwiXx+Dx7KBFt5tv/LW93PLe
eGsnAdxBN7Q0DjgYXIhjpQNhg6fAfb8jEzhySnxe7dEb6RMslfVDYOk/MXkQaB7C
/IuqM3gS6LB/JwgdesL76pnCl/3xX/2p4LSlSSg2dRpeG9ecR9Yw8OXf3YJle9od
O8nL1coCMZmq0nhjyTh7z4B9jDSA7K+vnEYffdFyjfVPQhJ5L/ercOf6uoROuU0g
z0h26OeByrm+XtUHbGMM4OcJXhknOoSBpyIJ1V7IKUA8p8zX2aZHk7uYsdAMVdls
F6xtuAUPEsLn/DccAnt8UxqF8d8KHpS3q2A+4WjxPXA2ES5RkeHJVk+of68iwcBG
SpoOWqMJGuL6eqIx3x5Ndv/gJnqcCwfzDAw1cQlHRLMr/wEEAznRtnXC7bnzcdHO
Yu0TkIeUrQsxabYZuoG6LvNJW4Lj5bbBxS6fT4msX4JHimFZ0lQU1LEWWDftDmvW
RWYvzfyswbzUup7jlr5UAn0JKDHVPR7L1U0awB/SRHlZxl1Mk7qhtaFo6N2c90hB
beYW1BZ/RXR6SLkMrdaGmbxxDf7CtaYhgO8izij6PyxUDwzl9DN+0kk/j//z4Pa4
VyXxvVStu89c96qVLw2VMbc+d7NrLyLxXSJivqQI6wYRb6r73a5hXMmoz41c4fub
nnTsybmExQSOYjwedTpHMzqBVWmRnkloRUo+tZjw7VyZ/+BuZ6tJLvrShs+tH365
oykkR+o3ad1+JbZSSDHuohKTBQQz9vn3EtLDFMIsSm0hOOefp4XHpLDrQRyuDQvw
OrNb+zab1ZRdO/1qXPfdqi7oib8Y3J5nP5QD8Nh1p6TmOOSB1AhNZ2sIaPsVoNdc
c+z5dNEaQHrkbl5IFZTxa07ClkVuwC8b+CgEi3yUFIBBBYe+wbLZSpVczYod8Axv
vtc2jId3EfXeyPPVpxPver54r3sVm7EFHCFMeW2L+DrhWz2o8KxWLteq0T+DtKDu
s9lTu6NbskCKXPOwAgSnLUzOIqVWaaykGrM0Ub356uJ4qLEj/CDsORcLjms3PY0u
XWBVXNmQn26mxbROpE7iL+PYD5e66V3GttI7+zhxL/H40n03wwj17dExavTf7Sf0
UvNYu14M49MQFqoTKANipgjbhg54keDIa3DbHecRjhjuSzDYEt4aKzxm6znDj4q4
pPnnURhQiGQ6ieFrdLF2pIzplPtUEsVoNwc0xB+X9DUrijcI42gLt9V1DAkV3wFK
NIc7GcEIm12gDV1byuWKHg06kACEIu+yDYjFWcjgNeaSkHr9/650S1am8UpHaYU4
RAqz80gSIL93I0V/dSnI4Fpu2zH3vj13p1ShquNX7lnlb4ClxuDfQCg72MdQjtse
DEA5jUghS/42ooa5mG2dPNPwSIeDslNDDv0Of9TAsTeMisg3hO5H4qjrJnked/Z2
c3bb7YgbZhgGlHYl18/MQwVFrct9IBVYY5clVJy6PfmYsvAVTZF08WXKc4Fs0cPa
8rVOASWLAs+9M0vizMg/sKvFZJh5tUd8NIh11BMDepNCGpHAIvfPKCY/XXRU0OVB
ZiAP5+dUkXGIDxFMGSMpGZthdq0uUrxorZrpZBAeQRRa/X7bBF++885ye8i65/S0
cp1/AA1I/eUYXCN8r65ksyyt5BdXjok7Z1CP/bKr7HbioddQoqjuqPrcKzLhquOd
m9kIsAZrronKGEovp2bOZYhUOtYL6fApT4KtxuusuHQ8z0mzIXoBMCwDJkDeVKOK
tBmYUQLAw1fwRMQJYTMkMsZgl11p6WlG/JWKy0L44t7E3pzar9UPJHkOBeqJi+fq
Ud2IEnPUTR+QoGiYy437pJ7wkE+mU9dYu2XPcXE1chbX3+DY+wTHzBHgB4cazE8I
1NhjydKnmTAm3NCUFarsWt1gietWnYGaaFenhB6RUlzxWJKa8F+r2XyPpWmdJfAa
dasJfTIT0ofJPmDGNPlbF4v9i+Zwkhk2IPhqf74c8M1p8aXBhpzoKhqUP1JUCec/
Sh4CGkPf9U5u8F4+IEdZ+8CvtoqOyj2DIF6zpOfDJt1ajrEmYamhpIRS0+NRya8Z
sjQT8o7jNqeOJBWOD/+WX6utJ1S/S5iLKI1M6QeV8wD7lYsfUPVqYr0QrTxiXq9o
2S3Eg2+RLS/wWPjTPNp+NWPyVQv0bd/eCQTwYjOHI3DuQbKyx7JgN3kPyv6leEG5
NgS7kn/mmwKYNLphGLrpxw2TD0BBeHUDXCpKF0nu9LhNtkK6Z+6hE+lbV9yU1MEh
gT1YLRVpeC3nQ7lk8cDj1doaeKOWbxDGtD51ciNQ4/eIZnVVck0rjRPu7tBOBl7w
SnYTMVZ+fJv/soWjubRpatQABIx6wlQvIJnxeBiFhWcN2mt1f+MHuoGjS5veI0Eh
8mBXQ1hlJ7Fs33OD8o2Hx1X5HhfpIdda5T5HCMnsM93b4wDdA7VZFwHVMlhAz+dz
Dpa8vkonKVRkGUYmJAic9v65MFEUUCWojBkIqcaCvv4FDodWaOb6jP54QhHlc5ih
h7QCOynhg4ENaiYz7X9+AM2eZdSFrYi8tQddyFxIduOtxzfVsdq7ssST+qSS0vAa
QK6FfV71BBPa9OXRbo4TuFP5liv6VHIsltGqlFd2QP8859uXkkCLfDZ3NDCGup1t
wePyEM/ou1Ba1XZWFVWxLCHd2A1+JeIMRKBMTbSPMGRN/xGArfkFWAoG6XnLlMGs
6T3FC7Srxx0v3mIWNm2lYSkTDIDZeArguFcELylCLZR/WDce7toQtajmEuvAvc7B
YMft/RsNRkMj51/YHz6DRyg+S8YrfS5uKkdwHlrZvqKvsqkOUVbJb2fT/KEOvPv5
Rhwkg9UuiNHnxYBlP/nTXE6ytdY83GqAs6far8mFAEza8QFha4eDj2FZVVcaYkXK
bGZHbZSMH+u9hlrr2UmmuPbL+DohvQD4wtaBS66Ooc2b6YO3EK+vi4Niq3wfgTlK
7sAwr3hVGFESjzUe5ak51n8r1HtuD0PvW5HXb1dNEwUy1S9Tfy4gfKvLPwmCPoW8
orCtboB7m2eH7mBpPQqHZsk1lu6r4QCC/ulbV3JWF5D7j1OfxZpMFN/BMgAyhfkD
Na3ONKM0LTEbbBA5z+afmOEr9wLvq9cCYPbbz9vdQhGtwp432zDpyI9rs3meZzBk
jECJ1JA3wDWAary4jH7AnGpX0ugTsz6VYNk0JKaFMWRmUZQM1dhIHdD2O90rFz9Z
bjsLQ8Bpd5gzRqAXTF5DIadSORAT8aC+APSTyTxOHTj+4I2aPee2FBEmXTpvQANR
LjvKOX+xdM4pxaBaYEq8//mG5Pd6AVvbx2FJT+pO1+v44/b3jSUfNSHqk1CRWVBd
qMspvQy3/+WIz0q/EqpfHStXvoFAo5eBOO0uMt4tf5fNI5C0XjhnhVj/NPBFK3Be
hDSzkTH7nD55xsO+blCtWQ5XG9+4mn0w5bivQinwnGJ2EY1KkOY+M98dQHjrQtRQ
uMElnz+7Ecg8a9DFLjxZslqEatlUoK/Yli8Y7+Z430WogMI2lBFNu3uk3c10G2hV
uFdJv4cbSqBHUy11+NG0sXk3E36dxsdtdRtl1V4Oc1uMPLUNLRun1bnL3Yaz0flh
diNF/y/4eJVGCHlfGce3KmqARyIrKZ6K6omqLqsHKCfG2DyF2BZ/UBao+rVN4VMX
OZDArG6AASK3YqEW7LSQBdh9W2eZ6iGmszMeawv1Xurj5nn5lSAysU6cAioJlRtu
uW4gLXq2H4kgr8NJ2BUv2ilUW4RGmBcZVas+0Ppo+hOBWvbcG8azdf2it0DwWsSL
G6K++kEy8QQ2MNGXhXqU188QhvEanN8D0UqUxtKjysJ19rXJbJD+61TKpOVJBDur
I3OxXka11Z8KqO30BuWoVt5RumbZt7lUJEax59JuQj96EGZoTSgK00CWedG9Rzft
ySHXtyOFhbuZWROxONd48b9HzIaMhKmQZS/k3zHE1bI+jTeOfd7NQszlRNJvZJgK
w39Ay5/9CV05Ioo47WTx/yQ3139FiFt7RZpfnoSFm4Tcm6uv/OEcxNzckOGbtDY8
vo14565y+l9z6ioAhek/SEipYNGEaC+8nIiPy8nUOumI/ZgsAesilD6BLtrA8Gor
GZWbssG9fCv5FUOeRMtqpcqDzqnxx0DDSNZuhROg0DE1dUi0Hga2nHLM1ncwqmiV
ERn5u9U3VnCx2TnnZ8BaaBZkaAGDhzzwqGgf31vFlGODZ1Oa+OBmAztk295ODFrl
azxhrEQraPkdZOQhYUYmsin4s+X4jqxPFd4pbEWSnmmbwiuo5qdZKyLkZCfUkMra
LGhDqr76Uk4Qen7wZAKo1HwChopyV2huLAXymb8vTDJ+1dh9PFsqI9dnMVo3bFsB
mh3BJ6mr6LMa0KiDbin4BLl2LQTmCKI9gQ1fN2bmxj1yrs6PxP1B4oIYCo7e9Fze
Ue2K5e+bPQm6iS8DDObbeCPJyTbyS4SLFvJHsBsQr6OMadloriCYO0b2M4raGQLL
jsOMnqZbqa6NHOkmE1jFPj+eAjMh9bY0KHJQ7Lx1txTqxleSevURzsgAr/n6DW1Z
MJW4rJoQ6WgvJGi2ycLQ7e1bHz3MZFFHkFC9qnYawEq5wSV7sCatTVaGbzzWTS08
5flENFVBHLh1Bfzzhs3Bw7w0FCLSbaXF1HmS8halogBsJyX0TovraRaYL3TQuXKA
JeSG3mimJLwIHj2PagkvPyfOzxbCkrmG+ZdyDj/rQMlFr5CPzrcHvtSRzaqQqJ47
wqPeQc4xIkyiHjq/sPPdwIehMRnikm0TYxI+tbkFeXAsN+BHdVE9AoBF74EYe36Y
d7GebSSu0ET4Cky8Hybzdmm9UIZMnbljJOcgjObqqZyL0wZkpJzvJCYz8qSiQ4mq
o0FaXy0wt7PkEOy32wgcuDECOAaiuRhc6FpxK+aUWRVbGz1UXWSOuWRJg7FLXFcB
ZIzT30jFtK+V7Xm0PcEKxcX0yCU0aWxSam+CX9c0EACD67OdKvF1KNIx1zxiGqQM
N4NYHdGWxRJxP3YUK3GhypKh0vXclvQvOhlrahIauJ71SJ+uf7CGGGnrPJS9tjAV
y01AeA6DQMIAGf5n46XHZqWHCTBroYgECNUxjSOvQJoxkOCVuxQkij4LTbmfjfeC
SR0q4rznxiyiDblDGqqYn6lcS4R1GJqI34X/vSlOS2SoEAX3hZlTQCVlX+5RxfpV
FiNNUSgzRo/xW5uVMgvhFwcUBrWgeTJJK7nlOZqVO0+PEsd+Tbd7vzMqhaFaKzG7
eI43na/HrteNkT6H1XI6EJ0+hQrP+pYCNSHzLT45CxmsiVFrfH7OxlkSJUQAOoL7
COF5itBFPCbJMZAfYNUOvDk9XnKhJGMkr6Q6uBzUFUStUR56/5tfJh95uAAKpbbO
lW9rqI0tctMA6hMcbNBRTDN0IrNP9+KqjXoSxrBoObvMOuWgKkUIh2PCza4BYC2x
53Op158qmnJqe+osPOvj4jG+JiYIxtgfyeC9vNhTqGV3MoUyBuobfFC/SKQYJO0O
ab2xMAvtyb/cL0sMi5wpFCRTvW/r0+ArAow1HXUCBAzduoPTyZ3az0rwNGOjshMw
ic5CsNAr4mIE/+IQbwPrvohYwL2ScdCvLMyjYohcgS8aSCWoG8I5AT+fIPFPgBS5
jZx3whwMDMhBOV1+NS9mLTxkWH5NK3dZt14vW15UQ2Ik921MLVjrJGIDJJXWlUJq
YKYcjWkOvkSkBSynKBaruGWv5+bSvTWUjM0DDaJRUtKb2tDvnZHUI2xpqNgRo1Yc
UWjre8RSuDQ4ejpDl8GO6ISXBcroVDFb2orx7ZzI3iprm4I3dmy7suoYEIvp+jyB
bAiq/A95F/YID/Jr6dx0kCQ2KLknlznANpsX9IRFa/aI0AbvnGq9UeOBIpPxNwLB
DfEa/VNLXHri5H9slYuoLN7WZLcUw43cYwYpRfPbm1ht7fzc0mDkdLUrZ4crmAFn
U4NmEBJ2qR7CO4j6mdtYRl3rgn9DDJrxPzl9BC52XNKo4cfzItqVczwFy8DIgvNN
WDsH4nf8HwJxQCSwjHcbmrKOYI2sU6ZPCDXYN62ae2MC18ZhvtCZWTU+DxkLYKXD
fLPdsP/DMWh2No2mmTLk37GKnBvvJ+rgoDEVeM2CkI6f+npORH6ABQxwRtEaowcJ
aCU85MLQC9d6cOCYnoZ4NH/OKDphWqJ5mk5VsxG7kyMeMgI3SuXKs7DitnXNT7AK
oYyiKR4QoYU+6wWhdYtna6mGJWAGmnZUormyNwJLKCU28x7E+3qJvaPrFG0cXJvm
6KIsGKKzTB5TVgZNLq/j4RaAj8ntBxnklcUVAHpj2/COC2PuO86ALbZKyDDIn6tI
4WeR5s+UrsdcO1vVWlm9Vr2wmUOFtT8yl5IB0rqZsynjtcHO/FaG+/KHqzQBhOv9
IgtmpJYCEt7OSxXE7oJNMV1ub0fcfSTy4T3cp3I44CoOSg0pgMMCyxqU4Zgar5qh
DXASIl1AxzZ8T3jnEYrKdq3je8KthnE1jOIELJ/veTCGn/57n5+QFw6lnuxNoT2s
PI8+qQzWLAwJOe07evARUIbCyJRhaYPPDrHG2bj9CTEzyiXIFsrkH2tPKu6vRUsP
o2SDsReRO8S11EBGoT/uQ81tsnK6DLi5BUh9tE9ki3cr85zTetJIGBQAUf2oJStE
Gys+YEeM/xe/BRrY2Excjsu64952ceL1jwSWSfJmTziRqRM8oEjGHRs0h+xXVIi+
cqbO4EWxn6/v1SfSau0wzwP5kSfp+CGTA5j4frIJdA6TbhwkEhM6dipQl8bs51Ro
imeghHPwbQTpFvFaqVgKy8gff1H5ghBoB4fEftLDTXnxagUDQWJbWtuAkT2N6coo
naEiGkbp/LHHt/oAZ0dIO5fckHHjw20BavSdfW6nmZCqkT6lxFbkePIUtsaFg6Yu
97nNfedpFKxYHk6EO+50Z32Qomyh98TQ0yHoDgU1x/Jy5bTq0XHQtQOS1XZxznb1
cSqCatWixXXU6ztJyIrJJuEtYZm1YgLcIypkC7oNXzw5mWmLvYAY+c0cRWiF9rDU
RiJxIwSBear6axjiP0bqV434JUO6+D4DxHsypQ4jKZsKw/ZQ54MPYotgDhMUkV8u
gjyrypb/j0EdRBpXdhV/ois9QtK7zFawp+UoOvx6tnGr9qKd+8Q6OERyaSZVzWZK
or+2ubBQDB2IG3sQH26SQql3F/0XOf5xNoFqVReekWjkDeOeMhoome1/6qZrH90E
mSAuDGS0DDqohRvCHoMl0rCCuMv83eeRYUnisi9Bs1sJbuZqnhp9x7VEQSZ8spLf
TLCoWSFhoFyFGhSVmoCvKAOqmLc/YogOZJndDDjiDRn9OQ6l+rJETLmsuRIyfZ22
B7KVGqMvsT/LvRpXA5+qty7opWljB11veAATFYBWC1Oq5IUIXPn49Dr8EnvaTQef
DpoS+ldRAT4jCr0yMRM2hGO10w7JaMbjmGKhh9offIaBln69kUDFzS7XvzvYwoJk
liayAyYV4g6zFGawp2fl9KALBNkNQUgsHheUweLoj3gIJUMayQ+BFMzFJRVK00uv
eOEArFB2D6d+/a9dyP8rsZbv+BVd24sDAmNxSz1ElrIgPJ0+FI3Dckya1AaOgQVa
v2zNX7Coy9/zdlgR1PWshxEBGms7aiXaKdjowu+wuR8Y/t7Wcv9JA24XvKYqwF1G
ZRwHiQChZbfZoY4mCugv7RZMiQu0H91r/mOPShWXvlHqgAfrHkA+WlHikko697Y/
qvIKqV4eX/IqMmR95pQiFG9SPi+/9gFmFlm1+1gSfLpGuGIwqi/J0s/4LcC6Gm6q
iol9Gbl6tlg0VAU32VXutjh9z9QuCa0jf1mh3B/5sf+WoEkHuyozvX8bex7HyKQw
hMwnONXVMSeq5qmKu1lzOrzsqP7lx5M59d39gpr79NLIhVf3ecs/+HeFmWn5lRno
N3onT+eDKArCeC2gxuj8Un9cxdFHMVezlL+Vyb8JzRCD/kLde8EXun3t9rJQmdbt
/0mI4nlfDyxbLBhr4ewuhE3BY9lt0pB/ycW6PVSif6jE1g0bg6A9zmG43o0J8xOq
g0QMyA/3T+kjbj/4Tg7rBM+KrMyHKf3oo5yz3kQdm1334hrgdDV6GM2LIR7pKQ86
bO/ZoLBfXCJA09ku1kdkKSgWMSmcS9rGogxwOYCt3qKrhggZV/i0S+ckCYMbnLWM
I5ZqyABWETd9Sep4ejPL21JeaWAj8ChQz7dg/ijQQxVEIE/LrHfK0MUl//fa4pcD
AdEB356ZbGDF5CQkrUhYHPEemR/P736byM38xD7etOcqwPhnbEDMIuN3PtiUW4NJ
CvtDZoWtpvGpTNMnSyE1KmAEIgBwTfb3l0wk42/7lqlWU7bcjZXDhlzetPSouSEH
IUcVm5R0RqTg78NbldVV7HVhuvx29Ont3bZ1HHPrVEUsq4AzQwssxMvnnzL+7QtI
D6wvFgHb3Dq8Rj181IQWZ0/epWeCD4iva5GC1bB7XqfJsVSiE2XlF1/3KdTfCxlE
A8V21Pmkm2dSQsrvsjutMASWZkND5tnZE84cguwcKv/9797lmzSvYb2Kt+oNPVKV
6beaW1RllOVJ7tjolOe8SUCiTIfV66rR4+qphJRzyC27wNgbQSZhPgvJiUebvIF8
EG6/9GHtOLF7YJTqVcMj1rX+Z+sQIQcsk2Q9nVJc7pHlUJ2guidyT+2PQeD+bjI3
qrFistHRJFIdvqoweUvB0LOvf11hp1jk6HbPBjCx8gaLqwtkbQP/G+03EezX36T4
mW1cjKVgcrVoeleKJ8WhgHa7Be9fSNqsGAaWRrFn8NRbP4Lf34sEiTj/7Wc3ILa3
cA/Ip8zixA58zDlbuF4B0CtJeFbBDc39OIIzJNiFFEHVw0XMrjjw+eHvqVKvbxIy
xXvYSLBPqksCjiRaPIoWGhfWPsyniHhBe1a/sxr+kZ5t9sRDYVo433Rmrq4BoGWt
iq95Lk2h+uwieotd+W1zsiLA4Sba5DI/udSkZv1FgS+Vm1j3TrDraA0CoBZ7/2RM
hy/mBQ+KTRqY6sxUSxV4cXJhAFOnDERaX7StHvsszp6TG6Jfuw0FhexQklnVHdRF
UCae+IO/+TCOBhsDzrU/oYSI1Qd7DcGAsypC28xxlN7U9EoVRsbFOr6hO7XDX+cr
ZlqIvzKoLQw2QTyqtsmirQnkDF2q8HfdTcB4l+hRoIoIdk5Tcl19g7ik8aniIc1I
KxQrWM+iwy9TjzygkkE/vFcNsgD2QIfWIy3om4StLCogSpc86YYGtX2XahmeNLms
lMemZH3ZmGhJNZroGrrB61azYbVWVLGu7je7ZosOgp2d60QbpTF3pDN2bdKtt41u
jRWClp3LZkjDUQ0K6dpumcRnCjAbjf89jtwLG9OpSC2p1Thmzf27E9ZHECooQ9o3
laSalx5pfQlls12Y7pS8q5yJpeYpOEbsYP7z8o9EzphPlFWsGC68uSA9D2BOFMal
+KEM54eSb/o+xd0eAC/Bs/EtoiTSsxYGAXOCmcve2l83roR3abNQTrUrZiV+A6SF
XwejIeSAJqEzB4ayCjx7G9zITxofsxnrTTkdhQMB0vi1Y3ZQZiHAumySUsni+0yj
tE7on/7mWCfEwVe8gZW4zIlhiHD7sPLWvjE7Jv2ZPbNe8dnz9f7L9Nfpg2+K1oT4
tKj0OZGKP8yULNOJ3o3QN5jC9RPGjXdFwvUhCMuv2QixrhuTCddbY5KzsWbUkTtF
pgtL+gOMntl97g9u3w9T16QCN6QtkyiLLducgBvWbs4Uzmxtw/C/naB61MlQmx0t
XqaFa2CSKZge0SJz29E8U/4RjyraxMv7lclhi4RdUkc2jfzu4axe8ArpetXd/9Fg
uJVPT5zEKA6+uuUtvmImxd42fBT2tnwh3ptCOjkadbRP0hsR8w2o7TDfmEtIjkZ+
apHrQGMsKF6iIEfzns/h4GclZ46Bub1I1cxFZvXTQtQEvvuvMKOaaQ6RmyUm5skM
jSryWcWCZtILdZ2H28bbh3I5lg6ylp8CCP+FP3cROKffi7M+lptleeYcTq7MCNMF
L+XwCVOUVgRBvnNJepOeYqfXHUZcI43mbGrbkr5QcgCDysLuqJqwB9MQW7eFJnCi
UnHmm98XO5UdW+4UlsJrooTQE/9Fsn6dp05BinwmQM9kAWhYHX+dRX55LEAb3Cr2
Zg/qqE+MJnkpk/QCurUIQy9MEI1084PK9fgJnAbrzvev4jNobquCObDfTnnor2Lc
3UI6R2Eoy3+EjhqdK9Hk6c3TOxEgNobh2GtHKfEaUSH4V0L6Hen76XG9ZsGQa/2r
BBAQQc7rYoNJKSCAmOjWQGw3pZztCpCcKEiFLri1Za8lAxN87SmzPmkagYjalqb9
PWf5E2Ce8mojk5mx5AFaEw883oo+/67dcMQTvjW7C+9oH0SCfVErSmdwlVBDpAIC
o0wRxImnU2dlya5BL6uut08wG8ZvRJ5to8gjbspTzMpAtEz1Vk0MdufovBB8Z+1L
w6520dgn9rPqguXDOXkPPemzChkpwon9g646WpBOSc+MmRjDP4/nd1FftEIRxnTP
WnDEwTm3RyEevg1Y3w7CeEpTtFbyBi6KXGB1Mk3VADsOilK8g2JfDQnoz2PhbjQR
iv4njP958JNONYz5qoT+BsftIAS76xEeNOtD0peF06tTN2ti2eJLvZOdN6nHz9s8
Ui/TdJonaIljUsVMp2lVpO4WQ19YBUysGbNyJllUmew3rftgoFAD8sXyFa4eT1iV
QY/aXBSwe1cv+ur1vpfba9U31l7+BScKXzreG6mJY2YXKQttLp3cc4JeaNVkScoq
c/AgGF5aIYNEQ7Z3xQErMbA7vRB1S/sLu0yCEWLaL3F0ciDc+H/Ajz7JlfejaU8n
ZDTP8rXyENGWIqxCaXzQzrfpZZX+okMmx5SFo3/IpeBv52g8q+vHo4/lGUZCHdO6
qu04Kno3ZLFMKX2142bYdq4lllh6BcKtlJVNpwhHCcG0NkLXlYohwiwoWNvYonQC
PZSI0Z7Kap/6+6fwEuX6gtaFeYIlAol8vDHY1zmQiN1TF9nAqW5LpZGY+STGmBZN
k0C4bT3mHp3N2R0beztvtE+Ug5w2bdPAniofz6Z4PKa5lE/WsRdFfCt3sN3+ngpZ
U3tuolWxBRnsxp2Kq5oLidgWQjnT1gjXCIB4WEc5GFU/GU2xzX+1XtbPeW4GUqmJ
9eWsVptZwK6kN2nXGh9ir0BVCRf1RJx+LDMm29E+vO2Ewd9D54jMbgBPZYVF5RUq
mONwrwl7FIxIdSRF1WKyVznJiOcju5RVEHLKOuWha9YH5Kq2lM/9iM4alZIaSd0i
emSITaEuqzUcYRsH4dn3PSrq80EcGqqF6mobtZgKOrG3/aZ7pwwpGtJ+/LoGea9m
gG94DpP15THzbk4TU1QSSBEtBjZ9IDkiJpklQUAbCe3AZpEeHuTD12vDKPaeLj11
8Vop32q4ECL1i4rmCumEG8gjxDLlkaVjazutirgdh+ATNhESQqWdBp6Lz8sSHAAc
FENhpeU/NY22JCRY7qlCi5WDvwqMXlKF9cm5QQqGC+Sa2dN2R8O9djQXx9jnHHXo
z5X92gjNdgYRnX1SC0hpO/NQ8B/w6wJyz67MQLIvBUiP4gPVhSlAnyjbACJZCZGM
nWFlOCHUowgVjtu33yFvU0i76lSAaWBpVcPmBWUDZGGc6G1hb6pqXgBSiXS4yN9h
Ua0p+aWPkR73szw00JgTzAj50qJ05TkiG8K9EqLsrOUvd3qHW2+zJ8RrzrCB25Nv
NHOB8rGLkflMYftyhQFpJv/PclmxFLXsMJLIjBzwoBOLGpvIgvR2NlcCPGCcBeZX
jwza0+ElHcYNCX6qsdlnrvFS697kW0Vyrmafh7dDZZnNnEEpN05cZrP4wtTd9qtA
haLzhnynQMg+GR7Nc+J/FdIjs0JCJzvEGsExdU0yGUoo7D2f+uxINgSl4ff6E+w9
kxYdjzTBFIw9zV4J+kIPn2mIgIMpok9L7WAx2r8C4RXycug4IF4QjwDuL4laq1/F
88MZBn+McCWcgTTq5HF+PKPqF/oI+4l8NycEWq2BqlNtFcruYg4voW4tt46EC5FE
lXQFWDGvwGU9q7Tr8Y/ARmGfZ20J0zgBsidf4Db/1glf5RuRBAkuvrlDB4BFETzA
YNJ2JBlueQMvOF5uo2PDhOf8+pJ7FAEPcbQ4+xcEHDzfVjzna2/Lhhf/JI6/MimM
cdhge6/x4BDV2B93BRs6S4Ln+P1FUK995iaeOEKqVR6jKuUfue4cXXuCrXXyU738
oPeUPnsmBVd2Mtcx2oLWQ9G0dYBmN1OQhQTRR5nLsr2b0utar+O6RJIxXUN6y2Qm
qqyWoBs/DGrae69Qmv/UfDSifF0sF0L0fYcYjl0U6gb7+i2dlEzbVr4l8ERlGF67
mu5WvgB0npAMvv+XVikGO35GGiGfzuOKWGQD14eDi6x72+jnuK04z8rtmQUMe9qn
rI5nNRyEDfUpzRbytjjSnAn1Fhs/7ZvZoVPodD1vT2sxeRRdAdGDsWcuzmGmYbJ8
UK9eUYW2+uVdDD+7Q2UOYe6bnz7twVIEz9FdMrpRMzat83FlSj/PPgLCILgNqnAf
X0LV4W+2uOedFpbSUmToIGAxjU9hf+nUBAUY6Q3cFQEd6/ZBMwafWt/biJy8COdR
AF6q3ClzVsJgIsFaeERhs5hI5woa/ilyDVCt+uTas7WbQCmbIcvwoGAUEwFcjtxk
977eM5QTbkTqWIaGnZEiuk0ZtBzlp6iRe/sZQqflc8oWaDvWksMIllqrSrWAp0K+
mDiBtr9CJE+4wbel7HO5iGfmTsXkPgrj0aE8Rny7ytVnwt2vJIe/gHDS3siG3Rrc
HTSdhI6iXPhhCNTpeFEJHlf3VyxZgA3CyEZ/4sbxb5ZWQvKefNhRQoCADwVPmMuZ
/DnepaBZ5NF3IB8JM48odrPB67mquvWvli7TC2YO5hyx4pY3ImUeTJh1ThP05bWY
9QV8IR9U7qmHUCcJtGVVFW2f+j9u8NV2bGeuONUXzfqazYPBhVqlhAykVbRjgQ2n
YNbMcgmSA2eNYVe8xTCLJ6Dji7BEb9GPOL/x+TlN0Z+BhfafZ5tqGwwiy0ZCetvi
UsxNjZzI3WmFBgGfML8hyqf+tVKcJ4ayQdwAcbIO09bQ2/JTsDfdJf4AsLsia8O1
xoLLR9txmbKkvXTr3KU2jSuLDYV3+RJH0ouQ1aBZAQkQkxakNx3K6TzSTudGutXm
7AhqgO/7z6WaFstY8Shx5cks1nPjiqE8BvTYPEugRVYrk2xj7Nfr4bC6mfASVkpp
sNUEe8bK5gGq5XiuijTlebfX5sN/MnpmET3dZwpOEea0mm+3RgeWuQ1HozWMGulh
AAY7gs3Q0Hiyw9miE4t5RmKtDyHhmcOGQVg7B4TbpA+vIG4cPrgnnl6dlQZwOj7N
H8pue2v07lOfOzf5bD9FOkKWL+f0Thp6mZRr6BMh+vjN5e1g4cpWScXLtlwT8Pw5
j12r99BRHEBfqYKu1kboGrX+GvToR9uE3mRIvAgq/j9KSiRAFWd02fuo4l/pGSjs
SdQF7ioMCgcat0VllVhPRWDTODJIBvP3uFWGT02+RWeLjoUWUmSbPttX6eKkf9Bf
Bc1/E7oJ/xu5uuct1qxLqObEqq1Y2wlLrD03vYYWjOVhyanWCBRxx4b9K2EuEnUt
Y6kjit/wf6bkvjUqwHjTF9aLD1jp+3f6oh/gmP/HhaMYc5LLc52JfwC0y2RRcVXu
VLYNx4W2xk/7w4PxTNZm7exDOfW4yHJc2cEFVUl6W1+CJQmfN1MnYE1ekQXtG9Oc
qlD1IPLo9v0N+xFC9oA2BcvlybJjuRqtiFl+nJxygNm5F1ZY7CB/6cv6i7X8eLGT
Fdxecq0Jr3GjLxo2YhSqPRk7sdKpUfpSTXaPUbK8/epnSHagyrJBeV8iW8H8K/6P
f7n/bI01ff+ILq3JhVt+l1gLbfIa9YzzDtxhCBy4Cc0K8tXR3ZL3Nv6VAksuzugL
4vGdLLIlUey89wTyPVdzqCWs07wR1y3264JoYQbYGeHYz0wTb5dJNjKIXahdW6JI
TiVj6LGNpbxult8EeJ8g7KsCTYwvBg3h7Lz0RDlOY55m+5zUlLKnSwHWJQC5lx9Y
Fkd6QKZOZUrA41JgtOghMtIXAwvRLjQFdohGOfUk/PJ2IclKcomwZOi+uxajxveR
bNImVFtJ5DnP0UC47mK2nhfXu/+B84U4uirIfp92Vi2CE+nrG8nQ/ZLkFi9uvrlI
vOZkx2KYPdJhVsL7m11wI+r0917u+M5QsGh5UnbL5mZZD8NeCSjZlo5+djpn9bem
MgWJ23vykYE1ToBaBJ/H/IE0ITR51YpyXfcRO5f7VPLI6hc7J2tZ/A/POAAUWXwz
sWnFhXMBNEmkrpcZeEHwaQt6qOPvuYSJDq83s8VCHyzaY0BS7BtGUYsHuIfAsb7Q
z/52wFz/byiWLPBmGxZi2R2CaeXp3uCqwjzAEWWv8lQcnlt9PGop9VC7AGlJP5HX
FQzFCM21FOnuFN/h9lOl+G9G4KUE1iWQrQLPOlSd/aDMtTkn6SN00mLacurCdKD+
HsleXIXVejqlaP1tpNA+wbp/gp4SNmXRr4JDzGIQzEzCHas6b/D0xaU1ZcyZ1/sh
dOq3RjtTHCsulDO4x2q6GGA0axFm2tAbPxdO0Km66PJ4co3wwDVM5qtE+JjU2U1K
4C8Z4sJ2ia3U6W37/O0i/tsrlvdX308chL9hy8WuXFm9I6M2XCX+BcLljeGWFpDj
yHNJ9tz7gjnIfpSU69vCmxQJWLNOW7J1npgPO2G1RASnvDrYK2Xk/6yT8wx5egz2
tM0k3AV82w26BYAOAZa1iQse2UEzHRSdrb49B/fcNiwmoBnU4q0rr+GOfYPYiZQ1
4Fcgcqu3GTv305hjArXkqclPZ6gBrjzOJTqJV5wSPo53c1HnR6L/W3ZuxZsoHkm9
tI01/MvorYPyf7kgGx6QOqBkaV249cTayoukpAJ+dNL0GgkNH8DBpiyszGijdaEz
kQyPGduLfFx+nL9kR1PBnAAoyBydlghsKMZFC3SzVo4gQp6WBfYu8pVwDdA5StM9
EEJXHkb/Gx/3abrnxrqS8kkJNfVoBjgoLHp/najI3Fh59ldDIt/bhEGVDjohyu55
h+U8A2NReVshtggoTatDlaDJ93SLCKwgrlXyt5E4AvlutCV/EmNUi4MZCGibM6UJ
+A/MztCypc04QlpUk2nEbR5UJg1iudQH8v7q/+JVB/U0vKeQaH3pIIh+o9oUqffL
QhvXO/jXkgA1Wm/DGMMyUuUcf+t/h3cvFNbvXFXkDH6mTh+gSYAgIdlzmFG/r47Y
FfPJ91nMCZuSDshz3NLEpJ941gC4ekGGKUbAHqxgvtkZ9y4p7BDb1/N8MHqqPwZl
z0WBgKOtHFilCf60tLg1PkyrPN3eunubib8dEF5P3uH5Qh2hjVoHzBqiLgbFlVNf
Fc3TVUipqwEo57LIGMq4H0yhRMY/vcKrEFcfRTpWSZyB6uT7QjIHYsuPWLW7tK0d
et9z2+C1nsE2a2Z+hY/2xZHqvKNJFUsvZT6j0RL2K5v2slxcvtcjvdFbTNMyDxYE
GBY7Iwj1uylDBlfq8IAvU9KZACL72R7mQDnKVJzB7qs5Jy6Rcg+vPRnu827VrrKd
/B+DLJriBIKnHzvZWZg9nedRJL5nGB2Qxei8MyjWFcynlmYLaA3tuMtoJKsRzK7k
Z9VO441ZpyhJmWiwIwJpl9YuTkIwHPX4jGa525A/OdvdqL0HLiX3XWLkf5nCdkG/
G8Q5QC4l6o1dJ0FT71bpBA8rji5Np20uldOGjFluRk7yoWTfq5V3EORN6zjHhaZJ
GbilmOwq03VJj10yPJZbiGjCyTnua7kFIFlbG9aTrPdg/3qlenOO5OghnLzG1tE4
0PSPeYrFS7sJNwV6yPSzlFxv4Ki4I7Pc60bIdJHPE07bn039i0J8bSsj6twCKuK5
4c2Z7XhAHmPcHwLyWzHFF6xv966qZXjqGfpiF9Zc+IY0rpwQ72jBtcbJr0fKtuMs
ncT1d7j2468kljx3kT7N/kmUPhCPhTnNpsvNU2HBWtBaJukORPz5aTOrEs5nrOlr
ukC7BjxasgUnd8bRfOxGCIY/sOFOdsmwn5Uz+Rh2X5MSfIi7ijSeEzHW3J+FaYFb
6vdu+YZm7u4KCM1t1IOm0rzK0Oaa63xwreq4I5igwP3fi2k2BzhqtOxWuhOGdPfc
ht7ChF1FWbUD1VqFXDLmtzGGHjogCdNtIKwEmvJlV1/NaHnIOvzxMajxV3diFFDO
j6dBRatXruujI3Fg6bnufIoIIc/ZuWYcEmqOWuaM8YMBFayyTNlHCg56OklTj3Td
2L/AYpDG65l4jnUFXMj/CN9hqBHUphl79Cc1poDPpWzAWeJN7i+ZvSrVD/r2bSa0
sfPtZaKh9c9+hZSsHvSSYx2/w8MIfULKrw3wRaZ+kA6cxd5Ltp0Gbi3Gnna1ingG
yzBGnNlEmJNBzCL6CPSo+0m4dUjcbITFVFVgU0mqwOgtkKvM2AnvgiFjcBrudhfE
uhhtfSxKtNZ+5RKmAI963Z85azjl8oJyQksiObpg0iIznF8xTWldDX2+f9NoFOdN
tJb0sYsDDhzixFijNVYdbZD06r8J598nk5r+P3WbqTvbLVvpmFrNWp0od7trpwBH
tl0ed/P8jADki6I6UrgszhPeBiG0mNllOcLfjoROIoZSbEOeijWjkEXHM+cyxOBP
7UvDC5hfVVWjjlERklGfnuve0+RFHoUGloOs51/9ZMLGb65+NfSVoKqmxVcqcshL
hcKZZPr3NxYZ/hs061kbsmDEdJnAGUk2X92kNO79NYGxjgyf0qtupJMuS2H1sqCd
jC211jC77uoKDpII1WPlftAZslAOswi9d92mvNDe3c0fB1Dl7a1J5+w//PFjG3U7
MedQKOKP9gGWT+yMCVReflnnBrYl1F67DsZD6u+Fuk5CDCfZVLQ9LUFxUw33auQs
FpCGCHnbnb/A3MW6pkxlq5/CY21K4s2iDOzBIWDedbp13XxsAnPD302X5wJST1sk
bjadj4tCznX+kiMk0wdPE9ZdNCICoLQkDoSxcvHUj9HTxWn/ikyxP7/1ReEBkn40
WnIPw/rTemQWpwKtqUs73xC1qbG3eHuDtYdHZCpjVXWKnmiqA7Eq84LIJcslPNVB
kagXyVtrK6oO77pa1bTHliStvC/udgPyFgnq4jxKM2W64IFptnZLwIeEEC2JV9hf
jSZg3uW0jWB95ZhWSU8q+eJI4jBUTySKyVt1spmppKpXaLzBw2HKPGL0tiDwdkZw
Qp7Bbyt1NpROGWAcloSNL5Pr1+72XnHq+hIPtbWvILtJ1z5gbUXwBwlBWK8qGrsZ
/Z43yRg8/fRrTVpmJS4BGoAn7L3abE0+IOUgawr//nyDE71Rj673JGosbtTKl+ok
PX6lriL57ESt1Z0A4mXnOLEbfimwg5nuYNKuMNtiUlwwELu7GGHoVtawW7p9lPb4
yHzgfjMk2oyKq4xIm0FzGS5+RF3qpq1sAIuRLdZ+wKB8cDpyK0udoB2Elqg5s95m
YIY5KcLdXYrh+g1GsME0Aw1Db4BjVDCJEAy5Bz+wSu6wmr8u6RkCV4vY93xKoxEh
4rE3ue95F4rRbLS6koDnYyHvh5IkZoWjx6Bbtcpdwfep5kFAc8kqT+h6kUa7y1Oo
5Zcg8akxwjLdzF5RHUnXnanyMB56G4FASDJJTLvGP+lnwZY188a72rB4Cpu0ERJA
/165SbYzui9E404vLddqpkIZc8cC0HaZ/7S1dSATPd+23iVGF4cpD/dmKsdV73kt
B4luP+S3NeGjXL0ZwEbUhyUciIy3Pgp1+Jk9xon3iBR8LIpSpNK4scFurlPL/Z1l
GG8c116dK86y+RuR227wZTDrF3GRdi0xqiDsq8YvItpv8wjfEXn3YmsDEUv2qwxi
VyKA+tdgv2f7J6++cwjLiXP74yDfPYdFhuUB52aVlCpNBw0IJBPVKVKkkqLP3pvn
MzRDP/iqmm6w7Di4asXpn5AaflR6jXjyBHmdPg6dY0bN6zLmgwsQiBTYfiNu5/lx
LDytXVhRCrOzdy9d76yyKATnYHzH3kZestInV15flRiUy6YnmQQEzVe4yY5NeIbM
cavQpc8hjWXODfIa4zYjXvV1RNRUbFm0uzpncrnKsSaM/8oQMf+NKFa3SFxzq01r
/R9LqFFIhkm72Xtk2VCdM8w0c3J5rRXqzclx3dxa8oR+xxhpfLAHBJrmi7kSgG6g
q1i1IYzq1WoueYSVUesbyPYSMjm5OVmWRPrRY7BqlrIe+wDQ7gOWpTxnFc4BDanX
b1Kp3P0Z3g7pXlBFKYSA55kW37yBOiB3WozgchmFJaXUUm6DOd2IBpylJdUQ1n/w
Wvf7EV9g6VmndI0nmMtW6bpkaIH68u6UaNtcai8D4uvvxJh3IW77bpBiCxO6YCEM
RN3cXgCaFhQk6TOgeKbijQTRaO6Ut7zy9u1oyygyEjplsxrd3AMUYf8b+1OguD5G
6Q1fe5vBfC/oCSiK3S6FaXXjo8TPeOQcojr8bHy7eBuwTtq1EsK9kc6gCZXURl2X
0GJd9gdzzrjNFh/7AApfWwpI4rhRTO80wzZVODhsm/yu5KryqoNWLwffsscpWT/e
2cK43vIsI/RC5G2DVRvIfLaZOPWup0O9rBTTn59kzpyk09eg9RjM+pmIxCB606gK
4BDdAzKYFJ9tQus3HG8/YYw5JSn9H6+LQU30DH7LfVpHsmAr1lT/LDKf2gGMKX48
hxpxfvDod3y2B9p/QeFy3+29THw0N9ohVCuji5zvvz1ydykbfxjvy9y0oKV4N12E
/GTXOyRBw4S7YeH7m7ajv8djuB3Bn300wSmBOvOYCGdWkrh1MilNkj0pqBD8/Juo
2z7Ol3gx/momLBU9aCT+KsI61MYm/MOxK09TDPtW5RIzU6bR3fOB0ceKwLU/5VrO
rsPSJzNm/Q+yt0LK61CuwG6LONZsksFRoEeYbAj1fT1wXvmzgAW4iO0+0xZGKhAp
xNsT+ZCJEhU7Ic3d5EmUil97R8R4Zu4nJREIEUQgqxHb2gjLqNKHFgUCcTFJWvj9
MhaE+BRb4NyC1xfTHhGF+K0oMYlPf2X23nYqWPo6bWD9H7kWGcjbeFPAf0x7/krE
bcuL7BUTxdPwEKjictIkh28rEyy1brIAuRIyprY3MHS4+Kb7q7ipRfLJ9B9Kn5W/
Epc4dBk3BVWAGTKzMNHfWOjZuqK80EM3XSBab8AEsDG6Mbbd/ffWwkv2EZUgFMwe
UZ/tfZ2Td6UqpqHbnzs0byDw+VUJfLl4kayoQVTaHRSIaQKsJh2qaFKkZz4jG61E
oOan6YYUAHlEQXmLwJ8KOqHIldBSGQj/4JG+jnBgk69UQUv1gFPdeHF9rOQk/Msh
u+1fULpD7ydDR0Du6Y1sXJ1i7n91oQFEhh6WVgZVL+FIkhy+5xBm+7nk+uo1/spf
854Sdc87Ew5l7oD6JIRKrP2srvNjtDDBULXWCLp33dMR9ciML0IOsbwSBYwFeC/E
T6NfqmBHpjZw/GhBvpRfV6FnIMskYj8vw1NlE++AD62r1qPXBg7uoBAiFTYJM9rv
0k+Vzdof61RFCNfjejATUx1P4JpC3rlcS1X9Ajp4xjSeUVDU8U4kgew3hcDgCfrt
DO3LApA7SPOwqmdkr8GtNOK04TaKimyFOYvCJa+uq22LCTWAcpydIv3yL2kej5PV
j8A4DJyH7R1F/U04l2JY8UxvV2B9lGlv+uZrhPg66ICIGFM31AHRz1etkphsPhmM
UPCfMxVv7XkxCUgxRFBqbzzVu576NvPiRRl/QFZuSjsv+k0/kNIqEtqNZy1ROA+i
2M4kuEhLftXwsm5aINtOxSN1fqc5LebUZzfAeRt2XePFugIGDZZzPf9SutBhwPca
jAkV13m5ANGVQysLuXkN5KbhKUaeb5mhGgFv1oXtlIElERE9dR/sVX97M32LWuQB
EdXAk+zmybgG7ZuQSwdf4Ok19ueWiPiTvD3ic2/uExwRwyu4ytDk6He0/Li6u4fq
+y2tVmauFave/GwDSp/zYFRs+8IBWsu1xXcF/mfjkFBD0/i8CYQfY0w1WveCiht4
Gws63Ff0bWfXb3xwKaodFti87yGXZC5lSf/EXcLAV1hc2M0tAEv5rh0SLdSh68FH
V4rNSCA8x4tEUiIsqHBS5wawzwrYDO/AUaGpFrY8w2eyESZVuwqpfCPcu7NVPShN
cpjgDLJwA5bTQdtL0Ux/Tb0F7dlAMueJA43E6rg1eCAtbwf54BMq/bZ278V/6Hz9
zA4COyBk7+7VkaHKkqmm2o2v1QTo+iL8Ha0VNjDEsQV0S1skmPu19GASG9Hs/Lu/
os0ytZie3l2aJUDGA0Cm088ug2WGG31GGBVWicUPSw16uj6LiYGQ9gwQqgFXBPQj
z8TbyneVBQlAZ3djvv46qoLUDgeRHpjm/d3GsOxM5m7fSunENgzi8ujL2mSEhata
gZzLeWNfxgC3XNLYinyU4Q6mPSKCAGHA+xtnYeZK+HsoaGMxtFYdFhe2F+JxIabq
sQfErzeUMU+W0ETeELnHFRfosg3sAD4VZrtj/3F3TSq3w2r/C6t+ToYRekw4ThcF
Gu7eg/Rd06hbngZLTl05FqlboVhbNuv5eekmEMzlKirmn7r0xgTIsysiFTapRio8
VDgr/N7B0CKGpBAbfztrzzf79rwAiEVeZBLbnaFoHeWMLHK2jxveEYF8ABPc39FU
R7aENkWgqQIvkxPT3suNkUGLl3SIt1a0ccBAUbG5gLqnxTwKy10LDl+uSFyWmEHj
qg9I/2Aao1Zlx4PLyJrZeNVOGYs8XzCWHb8pz+0UAPwJZVMG/UAw2AQjkS+TynkX
A5mH8djI2AFwSrMrABXu7AxPTCRC/GTTmVyLk83PFADD8swQlISlgibQhx6oYhGQ
JtwnWBZ7Jp3L70en/W8HMoM/o7OsNWJAekwlbpREQUqYgmLi70qnZpxyq1PnT5fI
ar8PB8ElQQVApGCn8cCFlF2tTfIcN6huYbVR3/txz0DqU7vKIB2s41qiRsv2XY+d
zFTI2kE8dNi+E60nSv/Nwl7KorChXnnx4Nh7J8YFt/EKPuFtWkI2srlGAALzKgTI
EwJhf+Z8ilYGpyQly3lyCN5eR4EHwnO6ekO468LdYrDVmMb5aaoMGmnVyfXSSIWN
e5torYxOaEY62Fq2sZfOIG5f6sX0C6CAiAL5mwxwpiggbvl1mjhPRg+SjsMZJIua
hIm5QHTeezQo8RZ+vIAjFKFPYB+v6gs8E03v5xDWCPeSBtaBIgTl2McsAawvw8LI
mwy/cietWRcLhe/cJ/yrPBSr+TsZG68yQMXF+nkmZrPf4lr6sN/2t8I0IRIKAG1I
xuYv1syVNGFmtTzC28AXnVDyQgH/5PwFKW7hFBdqvdt/hHn2nYVArf3w0GiQcjKK
m17GlZdB4hzUIruG0glQTfCEk0SKjRuiP1xoPmDONteMExM/E1uAY700gQln5X84
9uPrWtzqeqy+53pJIp9xfQTRGUvU26Pyzmkut3UOmsekpe8OcCL5QdFCmnDNpmLC
39D3PlVlVTwfci3TYOUZjR4jfb7dU3NZ6QH6KqYC4/bHUEL6Afk0a0hviZ9mDfAp
gGqEV0AdEP4i80g1nGGGgFPFMZmxNCzCMj1zBVh+jtvg/hMhJRmDr4PxzJ3EOu7N
skIYbE05NjiPh8Z60XUzV/jhdXe3x/yZnBDiCX7dVQPh6aV8J+z0EfN/HHlw0gpz
6kjKFlGqLx/D8N4+NJ5/djavT52nUk33y7xc1FBhBHCtNkjY8f8q/AiyOCadwiJV
XKmngoqqyuABs27B2/WV1N6HYV16OJaXwMVJ8eFdMWTORzmEQstNUKCR/7vp4qw4
v1e8o7HeodXXhMmNy+/z0whLBmAnHa/B0JSvBKejYY4iArWq8tzH3q83wyOf5YHY
EFcjutpjRLerWS+U1vv9QIcnSULURRedqfZLH1jIQvJdY58c1wexIowFPsJzGc0s
s0Hkkev9n0DGxW7vePXmGnxQ5sIUoTnkig6L49ZIO5u2UAbMewIqIixb8b8gVLve
j5lu2vsQnKLOEqlgZYkPRlT8XhM0eszYgtdzb58svWH6WHpLBRLAEYD8e216Vf/b
ycebvJi5cOD4XZ8uH+6TdOvOwHtyy06H7TgDXaVRZbAfPJgTDjtWQ7CV5Kf0Jkfd
oDSRtihRmwjnTuljpTJCTbO8H60iYHJGxE1lw3fhoY2pjaswlvxHuk+z3iWehC6E
uf6IAfa+8MZR4pKFemUzx5tz71wmBaTofS0uDW9Look2U4ZKIVQ23sHqidCkPOJP
pjGnH68JbkQSwkVq66FhAAdZMrzGXa2tnl0n6S+EHdgStwFdNM3XiCXDOyg7UcZT
OFThW7gjDLnu3NHTcLZIHm7DhQlKem9xrDK5h6F0gvZBMhRH17yc8JiMmcZXJJb9
713mtF34W0+/nzGm87ZerB/9F3RvZQOOsOMZQyqNuXGfo5jZaAR0zoPCvtB+WCbW
3Xw9jB+tb0yzHzH86rzO0r/UQfdNvuQQfwUHMUnt1wn2Btw7fzxhKhdIyZGJdyqv
LgM6MNTE5/unusdQCLmeiUP553S1qs0lZ+4Y7RjFy3I5E012oB1OjjX37PiSST7W
ztfk7mYGc2JPUQ4sVoPsM1xBwEFkRKInJJYQdcLuHPik/zhcXlPiGJQLxpziVKhA
VPEoaznI6Kq9VRJeyKt7mZ2Q5v+5KXdZ9fRlLAKTES0OgcY2Xnk9KSZk9AtPc3r2
reyOF5Uxvk7rx4LaHl62q9sk1N5AYHuuXNHj7re3ANHG5FI9rPZ/C9IXuc9661LA
B5anXlYOMTpx5XvqJgCVAkxn0j4OGWNpM7feMBmtCCap9KxfKk+5XAySwcIkxAFb
vfc6Bz2IomIcqwopG87PEjSFiB21b/NRhxZHyzOoKLLNTsquEaQbgi/tvKOLriT3
yPXfWCG3NA/xfT4sc/eiJXQwetPkiMwliLBcTkYfTb10gawqSOuRUxB+x8nm9FeN
eDEmqgpfdtRFjURRac+ZwlJYWD+IzqXG9acA8L4uTcVQikf7ydbXVcuds4FByPSs
8+LDWN4I3yvfLeEnfTdwycCb+6e/3bMo3hA3NTi6O4BvkovalEhhDs9YpbxlD3T9
05I8PB9cwi77vt08ok2Cd1NqfShELoPOUTwO8UdVodZ7rOa3P8uyVRyBrcGKicre
o8Qy6cxJsRo9VDIPDPK7VaG17UhnrkEr3XeUZBe4BgNYMN88Xbzwy0mWiJ0eAWGW
J5zhTsoN/h4CX+usVtO/2hhpPYVOGWg1EMjgFCqHJdYMsyXPcZiTYfR6Rd8LvFUW
l2kWFP1Rxz3nMeDPWb4VDzjy/+CHROmIaReK3uG0sn3zHXGkZOGpL6XtWVqrjkOF
tF195o1NxXoWUBFZg9SQN8IVV2dEXav8Cg5mHl8JQA7yih6kYarrYhWQdOjyMqpD
HcPxByJtVqw+t7nZsItrdLRmNTz4sCR9tTUPZaXRL56fcfjOMMeZkwUGVmF5UY3w
3ZUXn3woqhtqjpVwd+f0F09ADstF5M34vhU9+2ln6d7Cev8zDG5jikt8j9eZBg3G
pVw/kbt/VB+y9LRsxMKffnrL+DSpa9pR2iHihjyetdKg71ul2sNYwftRTaie0D2f
iB+SeCNPcmHsCqUcV5yvaGooEWblLgB5VI3cYVMSwiydLirzk6Vq3wPjbSN/WhH4
cScdWUzy9owIYSkKVQ2wZDnemfvAcNl2FoG6KWzZLCELGLEWwplLBl2KGruEWEHy
yGQJNHrsAZ3fEjMlYyU22Y4LEe0kssrYIQpBtZdogMXdvozFW1IhUTmuyljE2Wl9
VALov1uLPBD48/UqRSB8ryaVb+QT/LIuhF2hJcuKQsXgAbwKEBwj4TbTPSyZsFcf
g54eG5iaaj48oumAJODoiJdXyw/j5pXN+4RkceqJRDyoTtwcvJ2tJZFZx5IcsaKJ
kyGmg5blyPfSSm5s0jpEEPj+OoVSBPjXm/Sd273FgSPujKN/lG9ulDTxtVhxfM4V
Nc/dkyEA0aTpZljRUD1l1QwvW/hVDTjbwy8cjqWK2OZdXgDxGZkZ5Dy9ZaNYcuRS
ZsKGPVNB+377vi9BYwQa9vQwMbvHul50pgJxD30FtlzO9e/DvsX9W9JhV3en5Sfk
uhQ9sCXwatR5wNvkpO1evYgJoCpZho8IIjuOAocQjADox3VBssfymmjW5RtZ9+ES
jfQZLotVY8kpjcJiNxTVpBiGE9cxpzYqPUd7b4L5K3tFgqClbTPvjvvGnFJ8F/6U
oUD4ueMoYsuJ0zxF5t6QgM7/MkeyxKRunRI5npF8H1Y7eG+CSRYynUuV1sykIawU
Q5SkcueBBiu2EiuWuzxz1H2yCM43nzA2+knbKDTq7Vjlryy8QqRPdLu42MJYPetd
k5jXoldz+i15SCv2zIS40VfxLMNVlgzxHHFYJJZ9dDKEfUgX/PXv1SK8fX9EOrRm
Av+b52xvbPspQl5YwOkIvN+jBIl9dQ0Y1m/jCS6PKA4FhstgavEIoL9cYEwZAlXZ
yfaeZDYPGLRstyZLTijieyIkMxykEihtCrV3PZPxUFIWOeQW2f6REjAehGdrko8y
5Gd8Hu8+tbP7Sou6ncP4z+IBW6pi6Tb4xmTLpniW27/8LpooDozCT/vE2LupStZt
GuTx3YXgOQjbRjc1IUa2DnWhSh/gbac4x4Oaqe9+r3EP5ibDkZ5r+eeQfaaDqiKf
1Wwvq4v5uRFEXgNy5JtHDDkoUR1yovODK2KjJCDfPfozUkbwazmRcOkuHR4GmTQm
+aKM+WMi6Wn1YtidJ6wHOlvP2ndh5Dp5dP1rVHx3N7EqbDIWrNoNDmEbiMJtxPhx
wLmqZ7dmovBo22svYntibTKqnxWKXvOpvXHJiaLRi053HoYa/lA3WfOH5NWW9B1n
MbIHnuGq8acMG4vjN3DkMGZ3FFp3P9fHZLSivtdRSRKScnsiqOZON5meP/TTLyU9
YEjcFGUprKeZTOOC7VnR/wI11CFUrPK4cpraa3lLGrp6xWaIxDBRj9pcX4xXAhTC
3RhqiAbI8Rk8stMyUx/9f5AbD7/r2QvEsh3/6uXVTpN1r7GbxE/riTqYFkFJFfCB
hiHgnTEpZs9frF+d++LIjFi9tiz6Nn3gQ0RvbU7I8KGC9GjdP7nc+n4C7snFw4CH
0MFyOhhURkS9WgtGQV4UJE9rrdU7jq4jB564flOb4jrCWtAd6iz3PlW3V2+YRMPD
WJDRgLd2yn9hi3+B84Q4/jf3dm9wa0wz5ji5SuFqEk5wznV9l/IEhZh5aP38AsEn
MSVZQk3mUdllAu4GHe37JhMkiqxeYKNuDZp4l0JgLX+s49RJ5F0fh8YtS88Faccz
r0XyWusn59Kjhi6AAm1J8rpGnI0K4rWHohYdBYwpYCmdLuhSu72EaUpe3ZcLZNND
4Anpzvsm0Bz5vAxt2wGyM3RGzh92lHia5iG/XHjIVBokvHlhwXnHjBPTRUh7OWwA
GprFoYsvE7hki50t0xrOsqiCnnmtWzjyUp5Ke+e2+uWeneTSUJTJ/uCLaHNMm78t
QjPNNgMPw+W/VzoLuToopgBP7cQ+k3pdGOB0ga0yUlWn5YmTQIOthvmZg5uOovbM
yY4BdNSsLTqipkYXYKZuTl+xYBZWjEpF+O1AlANTPzCMb7XIzhmc7wwJ9mbme+uG
I1gOND1cdRxB1a4Tnj6oYr5Z572RdNGLfpNBh7J2YMcz4Gt87Cqt56ferLtQf2KS
wOPiYknGhiHKnj820gdTe7M8BkS3ltZ+6nT9aS1iAeRJPgTFJlOKQpk22ei32nPi
9gkcZkVNKtOEHnRAhL5lJ2e53VA6VCNlxezw8X43xJO+T/2+qdlv0KNYatqbgSS4
TGWH5eFYdV1VjPKdx6Zsls5Jy5GwuLlnCcgr+IisihpgSANZ6Jm+QQXBF67MJOsb
SQJYoJsKk0ZsVGK9a2QLD08wQJArxrgwJr+JIzNZSUPadjxnrEwsk+rsJeWXPkcl
XjDKYTP7t34VAwKmTypPwr3NUEFI/LZ+HozzPuaWBMtHkDyKdQ3QX3QOvo6gSkWu
1fSOC9BjxpK1H5rvF4uhWQzTBcpeB/mRkA0wKrsKiNXmWnyIEAXRObNsbDfJm05L
3puJrE8i0ex01ByXXw3RuzL4SFZ/kiggJwHmRhS/VPt9ce1+rfqUpS/Hlst0DCjL
p5SLSCmouU1YKJRduFhhaqNeTAGLSPU51GVwDtdZXiOy+oPmz9F3bCrC8zSe/+bF
lOkLj9lUDNSFu+olPsyjdtcg7diiKDIrmTDbiHtpuQ6zXjbIv/imyFTOi6O4Bvnd
RNvIVPoAL2Og5fx8wylvShCleqDUC5XsB9T5yopu86fjcKarvEFcIXWhJEoOpGTA
NDr0bF1Q5mW0JE0xwx9qabOoYsaawcBigJbrWjFAxLZTcO0fNrJaM/6+sJ3/6XMm
qRL+vgF/Cq7m/TwlhTc/ocrtCZjxMba8JC8jbmafDfs0eJO/FKaw0WtzGIfJC/H1
oq5zeF2Xki59XcNRf+ycUIZwtExCbiIG/xMWwhGpNfk0IwV6XlPOcHfjVa81VDrg
d0dHVG6pXT6XFRwIGk+YEWGbdP2/OX/wQ6tBCidLBiz0MmBd+1fWWxZ/oCKY++/h
qA3/Y6pMF0bCjBEpVn61vAsC/Au2PnfGo+GCxfCKaG6ODIUgpznptaS10RR9U2KQ
zRdidTXANzn3gr/1I52MnqBzveDExlz5AJMCAZnahaNsR0A1tLGXwORMbJZlMsEp
y2qGCvsh50aAevbSePQBTPE51nXv/d5mIgyXmWzN4DKwG7jsWY8rW7izaaje2uAo
VCSUcaIVRTD8+JAGq5AfM661KGnnwGtVLc4XIcXQKsFbKNp5hONxVBZbk85So0b7
B9SVEO/4Bk6kFtYkEWPxBhIB4ck1SP0fdQxRPQcHi2aK8FIFicJBIzaFWxX8NYiO
l2gZY12QxL71mg+R1mtXIwdWYPU+1YHnt0Djs0IK8jmjZhEK7hH9r9JOolQg1fiN
3iCgeR0gFSOfHg2iIF+FY7bVEorPvqbsiM+Z1S7ajDP6CHMFJCn97c875MU4ozqm
Z1jMsu1UydpnvmkDi86hKRfKo10q3XNTW5u/crx0e0DCfSoCw2Y/lXHRvSOgXE+B
sdtmGAREcjzwPmZzXOXuTJ+TX5gRJ+gUmOWsP4UM9RW/Nhqolf71VFxBAgmRSP97
2TWss1XUGXlFTz9pRfZfpGE42wgirwkEJ+7Aw1SQXT/B/dhIQ/CakqqFby0/+7CS
9YHJBgoXYb7Tj1xUXXj6v6tqXxpwp+MRsQkOT3bc1YY5k6XKhvPRZQQHYAMyxwNB
60BRukeOl4OdMARrU48CSaF8iciJA/WWIzq2W1lLJ5MuRzC6wrju6aoboXh4nocf
mFVbGF9Bn9Yzre/1F70DLUcH30e0y2KIhwOJyxu4G42mggMUU09CzS8WuPpz/+R7
TUUAb8UrVm8T7RpYH7IdB42mepS0GWiAuKFmdisLZx4A2E4zBH/bsbmyyuSVBisr
aWzGDSy114Ee9eJbk53RLoBZDrppmE0VEGQL50oZfbQhO6RiYBQytrqVmzNvMYw7
z5or0bMZ4S4xPZuzi4d4bkBOVPwfZGVGDkg1wV4oPQ89c9eWC+gIaIA+1E722VKB
4FVfnVgHybXxRm0fsHhpEP7JwRscQkTHygoUNxRY+ITQKSMm1acQktgThbTCOQek
8IjatoHL/1stiBloVd/dKgh5MyfLFAH0h7cdo9hSGz6kCJb2TCTaaWDvrhQ0yKEY
CGHvtKcmZ5X2mSKmrFoNrA0pdbqAiO2TxLTI+mLwdCy2pJ/N/+ndteS8V0TvBe7v
DAVQbvWcx9RZ0nEJvTB6E0v5B3Vj3bE95wb0o8Zax5J5reP29haWSy52e+FZoMVx
4Ne3gtEhe6UxRIO/8hYSW0USyJsU8jRhRxmd9OUklw2SrdMRLLIMfYVRIiUKIwEm
qoV2om+quyVIfGoc9VtzY/yxHhnfxI66dsN67+v9BEdkONtX8yL22O/KgR+Ap9vs
jPSxZvIJomAB5ge06o0OM+tszwt6ACcIu6adMGUbAgb+w0wcfUpVaMpbCdtqpJDe
YoNSrvf7td1buBv91XbyKY137EoIEzmr0m1axe21SMCUy/xtttD6sm7457D0aVIa
FdD/QLnitYD7plI6RYjrOTu+laQ5D/+LRaJKfrqSXzJgGGiew+0OPp96B3PCkfB6
sTTlTXnf+F7gLh4tWLEs9g3j1+ZgpKiCTOtSZ32B3C/xYe/zpsPHeVw0Pmt4uBd7
j5DtQa8xd36NRDuuZhBTBMD2nGx7CNY7OSZGBaBvpfU0dEFODSikApyjFi7snBvS
gyk9o8P5rDG4lRkJj7qj0eF9Qx6EebB0xm97onP3Ak8T8Deq3CqDQXOpEBzQI5Ya
czH8e0UD1YIQFFpMwPpw2hAEjoBzf5JvCGaT77OdA4X5P+Kr8Y4f9mKiVcMIz2fX
IBvoTKAF9ERrw14var1YGKg8ocnGFKUBRNOcYOxu5vWEqiKCjgtv1rcQUizoAlP6
bawReLDqukJ+wnoyPTBCMlxyn7q25nbLHQOlcENyTnpx6ar+tv2l+TTh8QLb7a37
xHlW4Yr6apWNuM2oie2KLqlJsaAeXac4RBGdh9su2Sr6XIfCKaJpd4j80YE/rzd1
xll2IkdThqpMa2I23mlSbDei99n3WyJdFjw2EmokfC+ySpgU24IOcR4v3lpLjG6n
TM+IJ9VEYsXDnSvd35Kw1vdxv2gYfHpIlpHcx1r4H8znP7LJ1Fs262xcq3i++vQn
wpYXgOHIb734Vx5PijChbxNC0Z/kLV+wbgV2rFazTWGb8TySv31guoP/dXekLQAh
a4JjCvs+/OGC2koyUenuPJLcEKzlLms+DOHnoDO/hMz0QRDv/MVXaCzzATroAUo5
A8ylgHA6GAdh/gBVQTV/39GjaKBOzhXUxRpbmnyQjRhkVgjzkjaBCiawemRq12qP
l1boS8LXOcpqc7s9jMrqoRvLibSfXwzOgjWvPlUD33qalm1EvWcon6Rga/U4gVf2
8a5vDqUuh0yPkRzXqPhbJpOfTt0Zmnchz/imnio9b9oViEmlHhxUoS0kjHE70eQS
l88k+Gb2xptGg3QDa/zDSyQdrQaGzVYrlD9n8yrDri5SXEH+gTEMpRtTzmFTnTnS
A0lEbfBH/Dp3fSGsH2T+Kuvb7lE7GUHVNu5ue8BFlC1xNiSkv6jYAwdRDn0hZFr5
dpCV/2WpFi5/XP3m/0N5Gl/UTOFBVtEBPH61TBQJoqZzmPynsXD3XivN0NDGIbRu
iMNz8Oikiu50EH6x8Ws56TOeneI9+IedrxWmihWsStk/5sCZxo42xDR8Q+8eHj1c
9SUB8t0YQcBivWhY3yt5JzxZ/MRbCKVL/zXXo62a3HTzFxVwgp4Jh4PirlPxFcUY
QXudxNZ1/4NKdePcuPUc1o8NaJUQmggPjC8bXFyB+Uou4/IuC5hLbNuC01JpNyFg
oRMe0bH3rne3bDeZeLWJRvIpLT+fkmaspAijvOSg4To6aM7Z6W/O4qhR5tea2x5C
Y6nh9WJuE5ljR0KctPBJFOPLcFnsPyRk8FdH+/WBxBjgVnL6XKYjJd1PK6XjitlR
2Cyn0BlZiCj2ZRIIf5HwJssDvUPx7gJPdJsw3rz4odGT+s5Vzy7jpMJnIV+bGwlW
mj6Wh9UbVGB2t4CFdx2VGL7bsE/WnCZZbcRZijDNQYTFhilN1gjC0s2HVtDBUnOG
IzUmM8YsYGPPzGOK+Le91NMaKAP1vRxdYtr+NOhuqpM4iAraNKhmcA9QPDiUVr+g
xM0W91+r9VSOLgLrhyY1GlJo+9NYLxTvyBRaubJMq8kUxzEht1kwZJ5nRS6MlCc+
erwiyM8s74zT96qBIJWjf/xyN4lgitXwBrATHQCKifMUCWecO9W15rxZV0wICsL/
XJ4bfYfxD9rRbMCOLpBqF2/v0wVzHd89615N+XB2Jyph6e/+vmBlvigUZE9UbQJQ
Arcb6xp0Ms/ySIdvYYwAL0fA4TmhKkWQV2BV4/NGYnuTNRZJ2FK+NoXEtUWXIUEd
4TsTlYSDSqVH0/pyyQDGgQhK+DC2topfYVTZQQ8u81s1dvpWvh63sqQJ7G+aEVR6
sNhJFxlEsZf45H60XAIVQze6XYAhjFtAc2ZRmO1Hvq6o1aqSNyebJdf1x9kNmPr8
3rD4G/QFk1SIWGNSIT5zKkh6RTkkhtcPZ6CU4aDfxdAjvd6ShEeBOdTZ0Vm5BP2r
LYIPXrGdIeH99mHb+ZbnbOJPWJVpBo79OhjTwq6EG4rS8lOiqDfZ9L/yn2qJ4mhE
UN8GnKebeYVdtRLem8oU9WwiqiaChTclyGrH0TiyX9rYDRJjTqS9jf5Lz96ImRme
8IiP0bWsAFqYk8TZLwT5vH0SW3cxLAfg+2E+tqEkjHcczHdf2Yw4PjyifHpiuXwV
Hj/PkoPGU4/q+zs/MMxrzkYXz804pCO0vMbteilxF9Mwb74mLodUKIE9J7GFMCaY
9Uftbpp+5y8KcqHaxljmdmuz37Nsqn3X/ZNJnFr2wYF+1z6j3mM4ckFFph2bgIcy
JrG7UlQYHDgRaepsaj/Kl7nnqCM/EOR9MG9QoyZvB7wrNOuCBailD9U53cekmmE3
XvD4LB25Xs8B7hJuXhPkCfBTyLeq2sJggZ1NGXcGOkmAwS64FplbnHVS4Kv9OdOd
YEKxVnd2Jv9NnxBM/cZg404LrX4o5RjJV1gmBdH60TuwBXlUVxLNXxdgIGPs2kd/
VswzWItS3nPSjxc3cuISt13hVPWxkMItwrjmvvtvue5q6QKrzzsY5hm2KWfXIZUy
3fa/UJxEankmlQYAS72vT2DpjckD3wifcdnbP0VT7KF2n2Lfxw4tfc/yOG9OZ8tL
vGYCWzXBl+ZFPnzhQT99xq4MSYCNKEPkJicYA3/RJ59C6vRQFvzlRqcmfZHZZe8A
dTDnryUqbRX3bDE+gZ6gRWkm6eeLzhmq+3zyS11iptlBrt7rmv7YnOth26pP5Vvw
2QXSuO/dRp5F3klZyx6r78CNjiKQh4no5uVqLMhm+lYJmEJN81iNkPAhHS8hhR/j
q/RY+Lzo3aZzf39QHAjda+3LLGFvJDMaKcr1bIioP5d5t/q+T8LVuTWCI4LmdYhs
cg7BwK62z91OL6fANo87gSIVvqgkAXBa3AFCb9TnTqiCtFvTaBxdXBxtNoButBBi
yWDugJ7BBoMjOD888rjm7vCn5i8Y+5vMywPsxWXx1gXqQ6rvnEIDWdq+XY+RMGVS
oAqJ3V3T7IZ2HBO9+Hk0EFLWGPyTu5wb2+/zfg4rUHHkEAtaWdIqq+/TyOMYM4nb
LjWrYmJ5HxukLvMdBK1GI+KzbSE4U+l0RCire9NcmpfxjVyl0AVOGCdipgZkZ/fl
Jk4yqmqAA9xQp1A+m8IiUYe7trD+UcNK/FrKS/t1eiILMyLy/oPTj8U/6yXeyBNE
U4LtylvwrWytIO+34lKqnXfnVK1oWJgA8wKN03KG1B4StNfAAYfAlwYsuyI5g3Mf
HRG2l7ZcRfIzH9x0oLMCeKBJFGwoqMhWHlvGsK+//SlsFymJX5expzroEdEi5K7t
JbqDu5xG2i5DN71PtQ3fVgsNhQSVBRwuBsmJALC2Sr3HKUtQELRKA8I5OImcWIOr
HLlbm4VEcRDsZLfgwFg5Hs6OtYcSooBf0IOPD03wSeA/wJgbS0D2Hvg0PBm2o/P8
alLyvnKcFyI2NIoNW99qvVLizCsz3sFA8SUThYqzpVTINQwZSFIOS33GO/E5vezM
8aCCCgMCxc9TwoSopWyYrf1i5voN6yS16MA9NRH1OgLqvTFGbaIEjolWSvLc3Yy5
cgQ8gELQsbiPCJ0d5yH+ALwtl+GP7TeXf8R3bfKKv11xnxxu+nVMEBezKNTvUlId
lAti0BWstutVi4BHYcEyZHrpYtmwOHPWrF66dtlgkN2KT+Zxs0GSkEOdfjMw7HBT
4n8H2ouxRg9riDMEgFkd9JAR4n3FbuBSFRMZP08UmLtBGPWGg51G3BxM6szMhDdv
pxqEOHnxSPtfOISl/JnE2K2zWYH5i9G/Sz+WE/NkGujKOhmGv36vYiUOI45JpGIO
ZX4sP9A+91X1VjbeqNPvu//kxrA/7PVlg5loIQounFg2X3fE5OQXxOqergaBjGSS
q8k/pXUYWbSAS6BL5dPDYi1DJfgptXhF9XiyXRh0RLoYe8+IwPPJKn3Dx9C+UYax
YfROSNziNOFMt71rhzw+cpD4oHmgOg5mk43W3tOhafWyj0IrX5Go806LIzA5Ias0
iZRrtQyMxY+EelfRvr05k5YCBNayEyFeqJmpy2brWk7gT8zdqQ+yXL6lw1hhvRWA
EugFcL5WkmdQeMiSq7Ml/LaOPEZz6SpoZTD0rNqlOASHzU+tsXm3R1Pb/n20MQDn
XeEPxClassgXUXdqD/LXzIcALDhuFoUlug/j2CeGMqTmlyHHVI2DSKDEeYSUkd85
lYJnosH2gp/m7FIEM/B5PGUiOF0dbnT83cSeW6f/Wpy09NghYjdgLV29sePIn4kT
V7TYoaQuaVAOZ3zFL3Zv57zpIz2GXFkWnVxVC1gL4Aw8IHLg5CXdmEtaWzWbhLgU
NTQm6OEUHULoP2WbRGr+GAHTn7u/Dj8bS3UV1gdztYWccwhYzhs3Xxqf8eZxdbLC
Sb1NYQJ//DIOWMuB/B2fR/INItSHW7L+izY8tZFBeN8GKNmUerF5iPZ3b3k7bZOs
QgCiOSYGzXDEb/mjrTiXje1xFIpMTfPuk+Z7kNmZevj8PANTpXzJZXJ92DlmjNGO
SpgoSz+WpXfWt/vd4ROOg3/VouxhWVNDiKMucOyKw7k9zvQlZsMr8bpTyK9iqI5J
31XJJjzuh6TYbyCmIWCoA7Cx2iQH/d4crmePNU1seAHuxdGZKLhajWJGYxpq75Ky
YXQOt8oNCHh3KjCVK5o0E7gobYEq4qXUqOjzScLWalSiNEJKNMvOqnJdYFGtzLac
NYduX8Va3rQLS9ki37JD2BXbu+5H64X+zb8cg4XV9dUSLssd6g4ED34QVQz4xfNm
0hIUBNqSiacQ25GV8uct3zlaOtzUqf+8uUsRuWgnwF1Tsw+EPrFaVfgIZmKUVF4+
8f5V7kcK4DaJwZ0VijWeMSob4x9bymTqNxW726F9oDtWpE931ZKvAm/dZq+dG4pP
3pBC8IRz+5hdj/VzxwK06jKszOTd8X6LJJLYlbh0HSEn95w3Abg18gWMUUUZYVA3
Okt2afwahJEQmY+fbio8nlMywXnBLfwiiOydzo+phMy9ajqKsOtEveRXdCnXorWO
+H4bB4aFyJqaBMZiSbaCFkfxMYhfvDMPDT5TIk3GMoe7fH2Lk2fx6bV8STMfZ/4g
G/Yu7nqXXqnn0DJ4L0TIpSewwXwo6WiA526uh+807+DxvRa9GLl6C9KLlZVNq/Hx
8dhMZKK5jRoRtLcucPuZW+gwqiD2Sbb+tN6IJ3e5FnNj/cwCG7ZvLi0QjcID4LqZ
BagFuhWp3h8G0CllugJBr5kLDMUq2DJWDVwt7c2z/GAehIDud3RFIb3XrfhCcM+f
z0jnjoUavu0Z8z1Zlk5fKeY8hBTuO0k84K9EtVH03kz4/7LN5nUvc16JV/rJeHz9
0CKAZp8vCv9NhK+vXW7fsqKoW20jgvKxDrKs3ZNJMr0sdVxRUENmgMX3cVwB7cfP
jU/ybDVJWChcy3L/SEv32PeavvfswPfoLWSbnCN+GgbVBxeQoYrQEYmhc/hvOEMO
FttSbRsVoT5KV6yz7Iv6ZrtVbBD5E1v9TGsM+neuGnuhy3GuVlqQwBaRENU4E6Wq
yNPgXIAcPXKXkdJXMthNr351ljAGsZ+QFyryd1yHN2MRpC7PFxnt6G0ebTxWbK+s
l1eHrMasw66evqJOuP1q3xGcVIpMoW0rWzw4ADxlwc5mqlm+ELuUoSwBH2IvdYcn
vVLq7xDY2BFwixyL41p9Jz4S/ulKjKjWfC4v0GQAP5XA563+mi/8Qj0ms7up4r+P
oQMlqxv3YpgJTb8YP0KTsL8b+0cR6EOYL2YqGKyviYosDOda3ObFbBnkud5u2Vok
QDqCvKpa2tQs9IKvzwSYh7or8SiCdk6y6hFpTVM/MjM+JuvOBS7rloJg8ic8RMZ9
/SB5NgGba2n7OHawo79+ZzWbuE05UHKHi0JN2LtyJfL6k6mVko5lBEX4E4w0s7p5
kqOGoKguAzW0r9hwkGbWetRWrUYfrzRJm7MJvR10XqjqLffSFYI40xZqhpqKiDov
xXUN8RYH30+ClM7tBs6wspdO9Ahnco0h+gcjLTUXIYd9qR147J8/Pv4vAHmQYAEy
DflumkIqsb6n2SqkLJk2D5y4RO1SU/rR+wyLy7Hl4zlWXU2tJKc0p76lDYlpzB5g
yrnOtvu4QZ18yNqY4I8QTnGq037c+OybNkz6sA5jnA1VwvASzh/WlT0tOA5GmYCf
5kPThcUi/X9/wPUtisBkiKZgHu2I83GViGT9CdddGTvcJBCVFhGuQ438FkP7bNlC
IMrcfNqtNO7mZodqVQnn19YYKC7okhfq/zNOrgyqld5dgC9et2Xh6hvZS67GVkk7
uFpP+TGaTsuYwAOrw9yGU+74BRq3AHf7g+E7ZRVZdQDN7SKpAS9eJ5iqp+JNVvzz
LOaiXcVwVH0c/H1wp5fDvlK51MUvzSLjOkRn1J7tc+eBQjAYHZFhq+EFG/ReHMel
uCZeEenM0z9mmCijZxJpviEee+fu/RYEAxViseFCgyoF2E/nHj8zj6hre8Z9Hudh
gERwayvJKWQwrd/LP7r3lUhdPv03sHK1h0DGNK1cn0qi7V3eUCd8bNoBj7EQFxkH
vYmb4O4Vp9w25q/k6d/5hdWoRqNtB986lqY/yt5mtltBpD/AgSVeUfhGpagL5wdR
cWE9hWLFCiCElFQpE9ypdp5VBIffmL/PbhGn0SkWYYGUp0QXzJxlzUHGsj1U/dK/
KYSCAEoHQeU/KRaQm7KsIIHdxeaSRKH0YSJXkcqPM2SWOR8E5JqmHxOT0Tj+IsUM
2wx9p5JsGFFRAkvoDSMiPg2t260eRASZYNVViCIBvbIYphiWPfCFhywvXlIBBglJ
XeRTyWDXnTsonJ4axenjBQsDw5QhH/d4Z8tftSgT+R8KG9CFN/y3/9B7kJkF+Lub
JIuBtSEPgeUDeeVetggzlcXRaH+BXnxE9nOdJpNSUZxm8Vh3NNM7TRhSI/qGqC3N
NxDhJQWEpV6ARI0HXTzBKAfn4NjeEu3X7HNwTDLluagvFYCME5ImLCJ7+kiM9J9h
eBVEpDmwbOSRzXmlH7Jx9lbBVGRqHk4zZe/BpUptHLeK0bDZ4CrxdHr6QA6fbX44
zVenDcdiJbxjhw6Zp9c/7D05FZ6mPxeMYYtzgY4FOuVE3GyP3L5KPhVrhHLkBxBM
aSmcihV0OUrvYW5dkSCpiwKl4UqPVfOpvRsZq5uEVLVZMTA5fmn63ppsTSkV6e6g
VrC5zsgRzgqQcEb0lr6TF0Gwv5MUwvJ09dHNZs9z0P3SveYGmp75fVwcRjIpI6DH
LEtB7rxaPdZBrfCZOVnyRHmoNj3tKKQJicc+NDXckt56l6MxoinvK5PBxHeEkC1Z
2jWyCBQgK71ixcqKoIR2BG4TBerZX77nGQWcGFwqmisBZLqMZKR/J+zk+5+hnypk
hARwD1hAF9CkOAX1L9R+jmlOJ355Cuut9SGMJQ45HgrEImVJqatRIXDTTxmkXBFH
RJpTTUjucbKHlGY5BUkcorBhTJORWvRxFu5YEgR8sAW45ftGc6EWfnMtRH7hrmpd
f6mkA+BmtWd8i1t7lDZOiMn9Vu81xtVuXkgpRDXUGT9R1w/rUQm8YCJMAsAyAumR
GvGFeEKLTSCbKu2R8r1kHG+iWKj9Wr9Yxrtm+vHl/6IGsV97UfY3EK/w5acROUXg
BSmM04WywiEnm8yv7ga3Ae3brna2T6OhH+skaVlNOPlmvZYmb+XGhr96mjo+Qo96
3zRWeMImFHGVx3KgT6/8eAnCK3KTYq0XizPIMm6WyD7PtCgfuFMq+YpM9o363CH3
LQPWdDeyKtGYh3apDsMLa+dcGVxR/rhBaWTAC3KTUlISyNMd2NFGOCUFcPQejZsX
ZwNhkHGe/ojP+qL2X1NU+u5wpOAIC/LGHArnQmTqtvNeDk3dzNsj0iz5h+Gk7Ofy
P0qJ8NnMlMtr7OMILtlIskSdsJozv8hoCQct8lV9gSvHN/UXE6Xtg0ivAf6mJqGd
GljJKMqKGTj26c9GEMUs54by5uWAZ8Yadbvdas9ywcg+xM2kzaCVbPswmvt472F1
4wuBdf4mxN9pFvKMfw6Wklehu2A5eWThr0IUFO0Y4oqxV7HYHdNQMp5mF7oqI0B9
0P9RhKZZVMCgo9TL5MP6FibrFfQwOK8kCCSasBteo8cAto7INSAvADDcV9N2ghKt
Gx7uShNfyj+bDYOxjcONU+u1wWQeBSdqK//XH9e2Tsw4TcunHuqmUHuy6aifKaJM
Hj6JWYDJBim/tS/1R4v8dxJbgfmNuHhyRzYfafTiTWXCOQPpsnEm0KeGRg7jc3H6
7W8nd4dzDwvfO85mpt1jxPejw6fj0Izofz4XjhgGxJ4yG6HutytNFj+zkCIvr3yT
gf/jW65B0ympMc3EY+vDZPE+GwpIwAuA2/OlG5pGT+o80mqIFBCgmkp+/Ybp1IBJ
ymycMF3Dn/jS4rnI93qBJZ0qQ5KKkZVs34YIOyF8FQrepH8aUfA3nW9Pyv0AJwJd
NrsUdb9KY+9lRF8z1vEGf2WcuvTODgVDifg6BHtsyVl+MHztsVQV4UgKy9PGwlFa
GHubPZEOqJVj0RiD0fQN556zzHewRFbaxps1jYLARa4DGk0YWwi57kJhf6qgwzH6
0GmdRQ98Elqzkf5XCNccvlFcCreBrmpu2jyBkZT8Rkb3rk8ke+S933WNyeeJlik8
pTuqqUXBPL0uZczrtnb0+RzHzg9T2Hz7HidwKdm7t+Bk6mseErjH1DazumJNYtSw
5XYhHRJW7S7i3hn892j+bk4hB9x2TJuQ1ntrXcxET4ZVXj5UEP+TlWO8dJ3HrTM/
pUyKOMImt/cq68tUYjFPBbKin3N/LmJoGj698oLKSjZUp4rXEQhah17wlrmtAbDf
KLJjPLNdTgUOr1UEEGccVrUiO+b18L8AiGwTJr0EPk68JBAIGnvC5+LJFiVlbzBF
i7Ru5XB2vkaN2CMteho89GTAZfacj6nFJDCQyafcT8PJ2ZRKB8m60+YGml2bKDgX
8EqZEWUqOvxtZU2Do0wWU8A628FmKnEf5H+dB4CCRPeunKFFR2v4HbtTvO23PAKR
6wkXRPr+npCgsophxXSR0HK9mSJvKETfY2+T8kBcFtP2Zd/Xrgvguz9Yiintl0Di
mdXEeWxul7roKMg1vZKbSP41Hvc+poqAk9nqamO9DQn2PbafwoTyM2wf4yr9NIsj
5v14wD0jTvBISrUKJwbpWdhDwNkznPDgDe9F+dKSK89mPSBpE1N07mc0yvPKrJE8
aLQ3U7UytrMLQj7Yzq8l/gD/XXtqcirdzwlj3KZMXwDr1YMPrRC54kWsOSC/D+Nm
aDzWWWzH+VrEEgFXKwsKY0dnoSK+MHbmrNYgDYNDRWpmniO0WaZuF0yCQl0u6zPi
8BIF5dD0QFNmrK8/3eni5P/50kJWe5Obd6iNMfVzuDCdr457xDXAz7tWyqYfmPOK
i1fc5eEkeCcFYSzX9cpGv6MOcyUj3glKUdBiVBEhvI3oLSE+ZDOvVf//bx2449OE
9bEpuvcgo6OEK1xm7k5jQwgd0PPJEyZeLzfp4Oxm+1arcIhpC0mJPsTCcOIgD+Lb
tCNtH5ianYs/HPKGs8ADDyQDcZafg8HEO3p/x1L2v6I75/MJ63Hrwp1rFL6G9mYV
P5Pel5m3480Lbo3FiD1NuqD9bzmP13ozfyb0BuYBq7H4OWvBmBUyjY6l7wMvetnp
MzNaQ2ExcSc1TN8gH9VjpSgsJAXQYcWgpJGBduCr2l6mdcxZs89Yf6nSzJLiUQ0w
BEhVeKIlNhJ42IBTM/GNFuf0lxlPxJpvtqN8a3kHK/5aNcFR+sHogjvspEO7qO2u
yRXa/R105l+B4P/47x3+fRNQv2byCkt0/4KnVuD4gfoL+F7S023WBmUCMqFbUwiu
yUwkbnmIxBhZ+D8mLao7HBMfkU9GaLO2vuWldpa5XxTqnT78UrII65VR1mK1gdaC
Swi0sIoARglpulG10n0+4Mx8Wt6PjHlMPuGvxK6ShhPWz7Arj2Cgl4MTOIJvzLWS
WV91L9tBf1sdpzQ7BWSmCFB5f3ZwlOtPIZkjCRFX7UjD8UQGsyMRvCX1ZpuFHZjn
jaH5ndeNAwgSnEq39OH7Hrx+GvKD+XJijgzhX1De/EliYi+e3i4JqhH9X0jjbcjy
ZX4OIh+sVkOMnsxphUBCJS2EXoRGVWLJ/Pt8b5NI500O7nTH47xp2YyTbuLOTGOv
37g2jAB7aSR3KSw3Es2y6SzTbPAYqj/brDopPiQ3eEOlljh6FYUvYEOh5IGF4dDJ
+Iozzo4d5Z1QHCkr+v6nGhGio/np45fIP34dotSGKPQGD6zxuEtu3+u1HQNFC2ll
GDkLW4PbNdQfm36ehPorsonjj8unCZzFhDNf53vGbgsIsZRV0OSTI1S4BdBjTx2/
ZTExAN56HyJH/4qwhD/L6y8r9ybQqCYzkA/EGKpogkvLY8z3f1an799SzUmqTLJf
EiHGS5nwEjnbBxRcqU5Nl2MwHY1JrQznuWuJ19EkMWXeEB1wKcfKZEj5sZ/NsUIM
O9a10pEMVvkgelsdMhdnA6wIQGS5sObjFofjUvny15L2n1/8HoDDiVx4l4gr2zc5
KFMlwMhcjTU0YjBpPMJh3oRR9dmsC1clFwohJn2L1QXS4M5Y4ZO0ivmSMK0YRmU5
rfhXTZ37w//1prDwu1uGuGsqXlFgErEbenvEEXEJpYWdskoRXSkKhQLgF+05InSW
BNixrlV9lBZ6U6e0JIPnne+tOftxf/N/pJqx6czggiGdT50spRRbSokM1RzrQWVg
wuyUq+6c9pXP5X5eW9ksqGQyyglIpZ0zdC7EHlUTKU9tuA4rNW96aH9LiPyQyL3m
hn9FqWPtjytguj/Tyl3YJ33zPqiOo/5IMuk/LB/hgOsyjDOuMns3ITxsYUzNPcc1
YjZR7qnZkOQVqHGWV5fcGi36uAmCfrPaETw6neWOMR/6w9JnwlasCedGnTmP3pUD
Xi4Rly0V1Vk4EW9uMdEb2Lk/uM6mW/8/SMb7joPMHJAMsCT9u507dv2dHyq6DlsX
hKcKuue2U1OypTMbeebZPYiARwbop+4nZXwNWEKyw6/0w5K455boQ7frS5pxEOCp
nwDeDuor74Xo5eQ5YcbYvD5t9jGzCd8R/7F+LPIApoxiSbZWcGObuY7acK3wNUcg
MipR15pDh4yANoBcOr9dysu57SJLOd9H1dETrJQBGZKboOUC4wb0iW7Uo8966GTX
gQoRkK+xuuict19Ym051j2GV4uapV21aGp9mbCIUp2uY2/oClyCok3OJzpLGag6z
tUt8uh02GFe7G0DLfA4i04ktb9qhSTDkrhy3sEIwdSnBcQiaaEkbnYQtCD7HrhTD
WZVC1NGQwiQqVS/H83FVQZPRTH2pYFQF+Hqzzci/t07m1WbdlgWs7RxRePcBxFJN
nF3WDITfrrQfme8ksLR6NqyQKtrgVb2bfxgXrO1YleEqMRE4pisYfTEZNYZipiIA
5NI9YAjg81MQxeKOjEU3yTPVCZQ6Jkt02UK6fbqkTULDyRJbMq2Ec5n9tMu5THLP
f5mPQu+9hy2hqhVWlcLJK97kI46fOXx7f5/KzvlFS2MytLQGGv7Kx9XJC4ZU2SUY
0wZcf0Y6cBD4kFv73tDwIUTfVWKN3tFYNqEdiWPEx3tf9OguhLQmpKFoCRGcUKJk
ektk94VO+u2ta5hYPkJI8NfeP8Q/nJKdQ/RwuBtWbLec0MRllNHgqFl7vvgbPrlj
n7XUTDXvoxwAM/dQwqJ3zdsfpoIYAaCdGNjrFeqq6xqMjwH4+46XWOTKbmwVj1vw
hNUxdy+PA1lwhavRRBi3Qu0kLkcP5qE4/jUYV4VjNi0N1ljD/rY8LklAZ+TMkdnr
RiUhDyxw8d4LNohWx9t9CQdzJYpVXoNAecN+H5WoOXOMxpXBUZfX0gJRxWJy8i3W
lJTmJz11mvELg4+Re2mrl+2xG+723BcXYVi2D89Xgi24YR/IAOQJ7CIBM/oMg2Ht
i9Sn1HKpS7XMpSTyn578d+39AdWPPGk81/6kOsoGzketrdhuaWuj6Ya4B7iPmReM
GSITRE3fgf89TEfhsdYVy+pX3EpAeJrhSIYwbNKjYvGfGl5t+9I70KQjTaUJnQ/7
OuNBPSbG275x/1fha8UO87UpZQji3hjEBKf/6VPvm2tIxGgI1W5I7lAeBgzpOExO
QsA/dZAtwq7RV3hKPd6PkmXds/b8/LTK0SesSObCMXmRdY0TXB+3ZAswIg3yWK/x
1j7KuuHY80qmGJZ6Sz+Z41DEdPGU4/5YN6apSPjVz2bfXtrqIuZd2PD7/RmKWJjY
2wEO6ekimTtFU5mkkvcsm53XIFPk9HZH6Jdaq5+zhD5IIc3CHWfGIqax+bVJvuqr
6Rry5KB3d9LtCnEzFh2sZrZaW24b/gZLWISBmK9NIq3kkPUNIrs/6vgf4Nx2SZoB
N5z3ynLhd/L7W0z2nYqmGSCYPhE4rWJYsaK0Fa+irm791XE5OfxcF188eCNnyZNX
mAailiUAI+W82SV05HswPy2WAgGVv+74aQGLy63TWlHgj/WYt+oI5GwraGPbbUut
LKo62+l47yheuaqXVNcA0HJJeggDX8wjFm8LXPZ5O5mFlMgQrC2vqTOOnFl2BKl/
sCNAF91Colty6nooQJbQF7MPjLLX2rtxoqQnT6Welnh6JuzpTsdEnEc3gt9yQlsS
SRAhzwwOjHeXtzHtGuk+HkQFjLaq5JLUaXuqNoPTrNsLLHZMFhr+HB68wlWjt3g0
Dz6SVrrNS24CwjICzT8ujyGLWkan52E0PAC6/D38x1uqZUrNeIrMi92lPzx4ndPd
obbaiJlqpFITVAbZvOOposNTEP/siIWyfeB0KMUzCCDxfhaXc7MHcD8wtP0beQ2r
VJXW7eIeRJtC9KU+XEdH3aKRDFxMAUCyjV6t4XtIghImkoEv8XUhzm3ogoG54Y5p
wZOFERL4+nWMAvn6HvltFROAEyJXlaMFu5HIK2WphsKIN6kJb31sucf6W0qlo2z8
HTtHPLUsFPDptUg04p0+jeQ5WX6fsnQ1TJ4X0wnrZ0x7i/4DYA8UFC+8Lx/jBDW0
ua3tkuKiFnxiPXSgc4lSdzTstbyR24GucV2wrsFuo8nfqI/WnNvp7ma9amdhjBVJ
e6gd9HeX7j9pe6mD2MV+eu3iuf10Rhlyt+fylN4xILkd3xX5sb179/Jqrnl4gYyx
DlcPfoOPlT4Deo4LbHl7pednvp/37OgCyooBSu9jlyRQ8tK2EkQwhJdzGOEulonl
+RA6YUwUx+0ZydpZrPdLDUuZdW2gmyYoLa4OF6U6kJlrN6jbdptp7POdUbYHE7e7
gkqs1X6qzLbqSPzY6B+fJdGx27UZI47aW58CwGNae6HigKpQVLvnTmjkCiyiM5nf
7LepAqiapiIBgr3qcZI+GD+bxoOzlq/ZI6Y/apdHJjgxqW17VdNvkN32PhDRALLO
HOBupPn3kORgogBcG3MropG/q/gy6VEfyGBfllGXSXkeGjXrwwAYO/sXzDuT6K+w
NA8cwB56LlflbR4DZbEv0x0Hk8aqD6Ttia/zBkB8Qd4JNMg1tsVCs33YbrbRIEDR
aLc9w6CjfYul2ZIQWjGNAG8VHrmqpyy7NkL4Cwd07omi7hC4/Y7OY9Gkz0nKvoTh
5lqow33Cbe8+nR1o9XosBmbnyPva/Ck0iFF8tyaweKwQfUjporczTEeMXBBgWLEj
qk2lu4rbVzZMjNhL7t8YNuqBv4Gq84kFLpTuNVZwrhdCQ0inWbUXjVPWZdmZGOEa
+Y0bXE31lY3VfDNM5EiexYbSL2j2dOvvJ0HMcQIlQNPKz9+YZIoTE7sZjnHEP2YU
HInD4vQKg2gvYOjF39xGV+yA/CwYmLw3N4nMsj9R9EQaRZMQl3oegWRAWm7ACDZP
MWS1c1biGOymJyMftj4mBL2gxoTzj8guW7+1z66zT29N2/BwJQKG+gMcImH/ks2x
J1u36alHJbKfVdFGuCy2ESQiPmXd/p3fHTMx8xZcfqtSmovcbY9XbtcLLBTDDIr3
oS5LzAQb2ZejGRBkaMbhGHvo9Th2h02O2JWumkfijfeF1KoPdAvhd24G15u6osQ/
eFRFTHgsU2DCKKX/oTVTWIzOHrqwDRUDDj5ZliTrWdQxAwtzeezONwY49HgP/1dQ
8f2UJAb3z47U5nYYUVqtxgYYBWp+VoKEpPvnJiDntcX6EHPYOIR1/B5jhnHT3wju
6Ddo9nnse9LFletx3+tJ8Qb1Tj6Y3D+GZ8YMphy3sHqH9Okh34TZq9zxRknRT2d0
7aHSzaZ+DlqERqBJFkpzq45ojNAGHjpg7G5hRIHMbR91xM4ZMFs0ukuNFJzjkrZw
UhQUiyg7BBc3UyBsQw1ZeV6Kvr7He7ULLfOB253kcqizOxkkFT2LOneqFN7p7qb6
j9ZmwjK+drANQZMPTn/GRO1Bq0/hWdDJR+PbiNzMkLAVpfZnR5oxa+T8wOYyPd0u
fEwKT5gHGZYwIbC/D98ir8MiEdPOGREIA7dTuOtaV440xGdy56FRRSz47nnr2vhB
SoVFdGIlanqqDaKz/Z9yNrMCh9wdGA8qRm/JmppPNzyNt2CoI1ioCye8SG9kMlxo
aGdgl4d6o0+uSSv9/vWACyQUXCOZWmi/hWS5yZAsYcMgQfsvNyiCfd8izfOItaSC
p7DC2eVjxrbhC5gHCOcxvKy4i0KuDhzuhmKqU/iFQ2lxIEe1AEZiQlzf0lvVelRH
C+er0o581ZrA1IDXCzbcXGTrRG9FtDlbKCgaB6DQmkW5mhzh1f9AF66snHlSnaFt
2kRX1XnVB+FWpMQv+0jsqAY+WFxmVebFrLfc1eDMySv+Za++PShs81YzVBgbK/NW
X5YDRQPiydZcypLFJcoRsnVH61b9nAu88nckzt8HmozY6D4BAvqZ6Nv96Y+vg948
1VVadT5qqGSsXybcZx5ktlfmbjKW9FNRYkuLANcmnNAB7Jd/j2RZBRTh47JfTCFK
P0wtJdvVqgmjNuU3CsXrr+TEhoIKkpuRc9Kb7VnQfRxeEY1dlGF2s1Or3gHgA09Q
jLs2ZgHzzc16ZRd8F7CZ3IhfKrmfCscqs1NoZx7a8UjdYTS1aYdzTVO3KBcnkjPk
8snNXEtgWbuNqF46vuqAl/+wqSuinnQCa02+w8tP41SJ0YIDv7Di2+rHHGApv18F
ZIVZSmmXyhn9yvJRhyQf2hoUwmLR9ezGVaMy3DWkZdl2RhYZWFxvzGv+1kdKmx+0
CNvllTHVLxDUEmnWAONxuZEHvx+VxDAHuZbGfzqakOA5WJLs1RIz5jOM3xLT31iK
CACbQyBOrtYQRczAnRRyqjn7YXkAeApZnpfBXsKlc9OmRHCG4sWHxhgflgSiQn8y
afNH3dG+nn/+LxhRoEfbjboxdapV0qCJ/bO2wJ/tfztiXbf62AkrpodNRTcvtnik
TC4RxDbPwpoXpSdoRoyvL/WwdhQARYDPEdg3aD+ccZQBmQ2UFij353DDry+cLRR7
AbYL1CMdi9+aG2fXqWAaImCQYNtz0RLxXu0rR4OylZxiQPJxLKcJQd914dfoq6v1
5s/EjVTJHqM5f8m/e7pdDcSxv3Vmi3JtJqpUIthqc0eS+2+RXo5+HsCLnnrO2c4/
Go4fTbhFRkCxNJ+itJyLrrro3xn2Ju+V6sFxhKe1G65kIYUNSZlNanGiLY2DMid4
8KTbKRDo75khYNpA4ducnSsAk0dEQYN7Id8PGXwNp+1FEquPXF6ATloIIL9TC5yn
k8t827mqIQ3zhrlCol2QUr3QF6Xe1Azn/rcy1bK+BYcpLGtzRJxVhDQlJyFIPCBr
TS3GwdpI9oPouT8N05VI2CYQIEMUuhbNj2R46y0pMEjT695Pfh5SbXtht5pFUXMg
fSyrZ6ZJGAykR0sdaDlmzpTQtW+dju9C5fhh7R03bBixdotQGsr6b2MyeYU6FAdn
NtDspss5Fpw8WQEsCW/WdksZDozbXZF9V7gO83hm3WQ6hRQzUfDfwdBfk6LF/iW5
qcF4pjw+APJncq43rHGSQsqVL2op10HysIvCTxLZx91RGjHAm9bLFOgYFj6IEDd4
2BD/N57mr0qP/dt0/iSOztfyHkZ/wEpQR1IuvAdLsCi5KQnjdxjYbXr1HR14PzOy
hx0BpGWPUz118A66Ky09T5MmEltuPWbK8FFRtaZVlhQvskWK0aijcwEppCc0xmyR
JZDyogHg93HiM1of1pvtLfYEPrKN1TlB2oG7NJy5w9hzrgvPiJiiJEELk+/SbOzt
Y9xQk02EaT4hqJKp33P5GaRl0HpXdYNhEgpjUECtXGySSqWfeIIsZP3XkEE/QbYx
27Yz7c/IIwgk3tAu/oy3J1Lb129R2YsBLiswISRDDJo/cPm/6zA7ClzXTLER00PE
MQJ8OX7o3D+OgE3T2V33KgJ7/ZLN/Ts6jqpgSSW9li8/YpEj/M8dqE2oSv4ubD6C
usQPtH6w0aAkGWqgxrqUD0LDKrXBl7l58Md1GSQLewHmYKc+9xQFzwQ3pWMe7Woi
QlH7LnLhX9pn5qpieVRym1mnw85Jm1K+cubDUsfih3vHgjdB85CjYHlRg4gYA2TA
f7n3IXrEv4J31nz8gY5YehfmPVldgHR17rFNtva8UeteZCxSQPwdNfKyg7b5dWdy
uugDeCzllj0QvXLHQqZP9Uua4aCmmkqJtdy6dFk0XcZ9EjrIl0BKPpXTAkGoaoAu
6LQODX973nDxg6HyhufLmUyKvPdc7c4lO0XWhaTz0uipNSG6YHn9xe2cLP6LWDLn
4GP8Nn9LINvXkJL/gSTsBHa79FoYyTlIu2SIC+9DZvKlgiF2wHrwAn0stN1rZlg+
mz5id3BmxdWIJ8CAw6+xliX+7TdrZM7YbL8+GL0JqxNDr4+H32KeT5uFaYMkS3bt
vYlcY/gh04TBvy+sOeXQHXvTDTJe1NX7v4KfHCs8+2am5ZQ/C4JWYzznZ8+C+gDo
9qZ0n8I8VzWcRkIG08Y7pOylCg6ThLufZJANsMYGOZanSnJsn4/fn6qPOSoBsCzz
Ay3vJ3h8XDASLfVEUBL3R2LHs83ZDPkWryo1YoWF5qBZexzJICoLuFCZdA5uKcLn
pGPuOiqReNKHbl9aHAzs7SEbOsEfqoRS62ozwHpHmL3l1qBRDWz5jvNsYbP+dXTS
JUoWcqYF/E/E+xCyfIK4a9rZaRIiurlTtzbIShfkOq7AcViAoIvqF5e74BheB6+I
hY+on25PirActpGoG+p7e+UsBr0p4RN/mahea93scMH3we+spYA3rRl9w1mWznA9
K+qhBzxQhWvL6ODX7JxfdScR1jXQvQ65ae6tvZXZwq8nVx/ZwqIjcu4/ICKN9bL6
65vJQaAE22q8/aRvk81PVMvKGqkm0BvANOGlEioTC6dwaOaJ+2i4mjd6xJ7RQRCT
myLkoHcT45tKUnu+gX7gB2BpRCrqc5njB4IYO9rmfBMX68J+DgfpAvLnQ2ynZqf7
vDyt9iosYzHrhXxwjAiNIrFqQl0W5rwQbENcTjVDP0SFKaBAlxI+9NANQiRkBxTE
LKxSLAlUVOSXTkHg1S7Zw+BHTeoApoAKE/eLf4gr7XsKaOZ6+3Ro20F6Q2XJZBmT
xmq7yG6VciwUtl5ckbShN/uyOPVU5xGjMDQsJAyatxXRJxGWgB1e0w0d4Qw8nAHe
Z9G9WSqPz/BWXieKNtIL06PGQYuQDXbRCgu9lESod3Hmn3rD+GqsSPFELVfrlLh4
/DtRHA4X6F4ji8808wLy2OPFGNMugAC9jaoQ5OAAabugCqWqd2DGjXrnTroDCHhX
WlANTLt1fSzPlIHRnzK4P3YG6QNabaHgSNDqS6Zacu8Q3EXO9lsy04FNHbzqty+7
NQZKLgjw8H7DdtNIPqi56E81sBxkTNQ4sTMxcJG2UTDAw1D/6j4EqpPqhNIbRTvc
ZPtowPxn8YBKxXPkHlNib94lz7p6c52iCmkZ2e42o0xHe1FstfjTx+9u8M13PBVj
x5nP4AucTNxD1xyNbg+KS2nuBwHhX3zZo6wbxGnnmGp4aQAf7BnnuA3Wpo4LVzFD
dkqVArwZ3DjcU1ptynsL1mpeuRGPvSkHciWxqcKA9TRtXnuSY0jkFcwfpLSiozLW
ubnXxoUpp4ULxWoRdQZYlr+u5iQEHD5xIsve5IaM4eC2cpW07t18XMqgnC5v9W0O
U/sJBYCDJJJ/GBzHwk3+L4Vmjs/JYoYzeEi04gHgu5GrwRokSWViL8ftoIs2PbSO
r6+GwUhNe69qq99rz6PSHE2Ux8MrxtpFkX6WQWSL/HqYGh8nNKRg8Ar0hKZ3vwai
HjBHaiY2FbAobKRQpl9CjeFwwPY527CyX2mgUxjMO1dj+XJrAyz4rbKJri5t1ylk
gENjMdiy9KV4HWtQy/hwiEEVmfdIENWy9SnNhUg2kyqbw1HOrA4CRmdLDuO8Q6Lm
iFs0CZDZq+84105Qs5o52DzYMQ4hbOogufmd1FpHufr+400hizw/Tedh2lr3Nf7y
OYGmj0TzDzFMRf3kD4EroRe7yuaTAhsuKLGOWGOCb2wqYSzNDzBiUYmNGcMvi3fn
u1tanVz48167sRwCHdHJarYx5FyKwYOZTJ6YKW8CsTuGP+wi5FTLAB/IEr2+SFft
ATVdu6AU743/70mkKROfjm7xj+pBhdcPlt7KirCbuKP/7VyvIaywvZfA9KX8pW7X
OQdi9DPFxQMij4BoMyP5flUCKDMyS37WbGZXepsuPKZA4qd1kdhJJZ+6V72/CwnK
TSQE5aE9GOGk1ErbtKKclFSvbn36HYkfD/fVRLA/0x0/s9f6ipirR9kwDMJf1lK3
E7MHrBFWT5IG9uAsgSqKd+Ee3U0746DTdKWetlsp7HX/qNIOy6mIiEd+YRwbpPGd
7VogSNPTXx3Zx7/+/W/LqAh49P5+i9ttiMGcjLFnhoiXAOX9u8t3orT53Bav5vQg
Al7TsIvgVhVNSPbhruw24Q7xiWFBVz1NOBAABw6hVm1BdM7EkmTk1Vbxp2Jd/f7L
bQteEnEaX9ANGtoMcIIWD/FLejyLu6DGiHCwbn0GwH9LZ9Yd+YKdvyLjEzDhDzOp
1wv1H8TcJkjsBbmFurfQMQSR8lEGDDVIc5gXO3EF1stmXRuzNX36XLXveL4Ibb2q
x6rAM2XKt5pe2GfNkXI2gbwr4fT3zexeh5UK7vs+s6K6NPmU7X+bXDa4OHAkGQ0A
8/XXTHFFICowyqC/R7mwJJYLd13x4hWntEgnFbcy5RevKgBXbar2+DFnaI01u1OB
OuX0XRpZ33ixbtU6+h9OVDPiNc5mmjw8CwlaNZSbFFpKoUgHn2FsOORWKvT+J5Ub
8+INgqPZiyCN/1TL+XUWs0EtZkMa3Va3myIoAFT38/d/HlV3WBCxLO8fkcjDBKst
8DxIf0S5+9+PqEXYCzYoQm64AfFZ0wzQRDxlwHMdQIf1TyQBivz37CbXwj4LaM1Y
6vvxxM4wmYohsvcZnExLCbq+39ddR0eGURaFjaHcC0/nI9B9vYg+N+JDHocjGz4t
I/4bvPyAhTyjjnjKv0jxu38msyYGYFBDkW7ww4i7rSd9EMxTGFhhjpcJdLMehS5J
KKGX8KK3xBH5Jse5HhrtvrhwENN37ji+T2pjii6dGN8+O7oh/jby1jSTxbAWx69s
/j4QhE5sX+cHuzlz3fiIaoNdwnv19iur4MlpsvdhDaEuRIMj4ROV7xHZQflNG3q8
iH9+VCuVxamh4rhfYQ9FiNcBXRvgf+LhIRUxVxVgwCvrtYoG648x5F6koLgEvD1h
AHoT5KmIgPRgiB2NhOPU1n7Pjm/lIoLT9/RyLoLLYv/sqeGYUBUwVCWxWOGA4DH9
AHVMqfnp5z2qK69kEOFc5xr2Bx3DkkqNsOKxbnnf4zi1hGlUuhDq1IDf35DptgPJ
5JBg4v6LxfvedZy7zsNqbwWS5ovIT9I+ZI79Fqf5kkv06oA+nFZhItfqLnw15UKS
4PWGqKP8LqYCajrMOs6XYLkNJsyR5EqeukJaE8e6Z6UdNRoGiCCQNHFLTKBuX16Y
MUUpyqYkz91e3lxYEIZsiX+B3hF4hfnvW1SR+/HT1mAojKvL5yGu9HEyuuRlRy0Z
G5wABtsK2Y1pfqy2KCM31vqZkgCHqiMaxV+hmSqMH/ZoUKD/6Cm9kfRmzG/yHg3M
z2QagMa436XgtG95dZ/isq7dJjB8evtl3bZsZ1+EybpiLaUyedyvZCiX/P89Vpvm
Q15cRcNjh7CJwhEbpMuRzVnCMV3YtVaV2d/WZ/HESudAjI9Hh8E0SS1jwvktH9lo
ERZpELgaSE3o5ShB/ES1gdn4Cm2lqRFCtiKAhBNSGqFCMhtuEBCfNGrDycSYZ2er
enZ9qA3lkbXIH28/OUA8s7UQqtNeS3Id06lg2v/NcBSUyd/WAQguRlSNLk1ROAsA
4U4rfvy/x9qjqpQfXbzPpW6rGK+mkIR47vyAjPTzeYywIjj+ZaNjQ4EPYk3xnKEG
drE3NPOVv3Rn6WpfzBRt4MUVKNNOvjhSjnPCoThgdi3vYGnXKbTYuwYTTD5fWRFs
rEmU0tqNH6+I7kWthKGFMIT/DcZSJeWSDrmQSAGiiokAWvhqMkqPTUz5uBj8eg1W
CTcnjLeGfMVnXp12PyNhXOs5AA6ojOSDbnyvE05r7AbGv8pIyBt1D758xYkcpO5Y
t0YqVrqyPOSKJFJL0HA+ug2lQt7Ckl1bJIC02Iw4uLmm2/o8tykeSNZ2dk4ZqVLO
PcGo7nrtFPgT1C3pURLxhoWxSafUqk+aeaHlXq/p7yomeRFmwLBTIcarURxue7cF
ADX/peN39q7QsnPyt1QVJiSrSdWpOTCrsKF3uN9himRYSgK/+WPM7Zm8fnZ6MDJP
cjJn6EzA8hCFG9H/T88XjrwFAVyzrLphJFQ2kPY6H2iNmYE/M4YVBIrL+aO8MLpV
DU4cVJTtewWkIJpx0RJPrrJ5uK3IdazE9cOE4fa/W5SuWd5oX215CUoJhZdGMdoU
XJ6u1jKGfOwXQ8oz3E9xjeA6RtSof6PjLOKSQWEhAc0mtrNaqfJW7a6p+7QmwopC
hmJZY/9GHlEpg3yuUoqf57PFOhNQlFA9aT5yOtE/YqvvyufkchQ8qanCrCz0H+/a
mEhhOO3/NOmB8wdB9AZwJC5eEQA80Ai7D5pBjInBraPUjVplsxqEvu199Hbum8Zi
cWGXvZEQdUSLNiUmDR/GISVs6TGQStRTJY+gEaEJXg1md+FXxpDS2+fFJ/+aZ/Xr
irdggeREUa8DUUmqZ9natMq2yO5H3uG0ImCVc+qUowrh+nW9qk2poYlU8RaTNjDW
KyoZ6RzUNRbv2z+5qsvHX0bMpOTLESuK3hTauqP8Nhxez2mw1rQ/9oPijlii+hej
2hVEGUT+c3pwMYzanvQ2dSPTv0h97VXkOFwtkqeEn5nQSM8fyGEo5Lk7+rLqSOIs
OqYijn1eNc/oFP6qghicBavyo4n61j8sgxNJJOy64SKuCDejskmSbSQgXjuYFDQ+
ts5u28TiVUQGRbf42nfFILiu2GpVJeNAaGcDjoHgMQ+Dfp65jo2nGWXpSzqiytRo
NGEVo9QsEwZ77kuMPJOsIuOUpgqsjcurp6EF5IlFxpHw/f+DLYOzyGstNvDu4Yr4
Z7TqLacZuUqXcHmTuDsObXZeSInj3vwiM828N9GAfAIY0tUozxJF7fugfJ3eHIRl
NsCBmTVQi9V+Z3YMWOErhzUZNGL1S7rJ3oLBF6L0atlwDjkmuiXjcguPgQCQepo/
vbGFJqyMQODOUevZ3UX8zDKZKL9/fQRVnTFtqyOC0tnGSCLt7mH06Axs4seJF6cn
WcpJI9zYFuz4HwI0jZrbQ1Yzvgzr58xVcAQKUI+ftAb1eZR67+tdFvvdsd2npILU
DB40GCeEwlvoTsf6y667mtdsKyRiVDkVHd6RwQ06xte990bwpScmItwcDp/EzOgT
EukRYKfFpul9NE0HJ2NbEz12kxpRaaCJX09OQ1YyjFfOSJN411jpqS92PzAoEgMw
boRJTRmbLiTI7j5tT1ym9I7RdlWuqF1UisgGJt7YnJKY47p2LxSCPjZG2uZPUkyx
pAbtbKJAaRYitcIDTgP4AN2YEU7jdPBqzknBG2tyXcCY1l02T9A2oDgVVNbrX5wS
KklTtmclmoAsDWJtMGEwjjkGpNXMzy8FI3WfX/FxZko7BbBqU7m7T4zylzq52nbF
YXNPCJJhxZ/pBiKq/kQLzuwGNRsS5Q71cK5106wKP/HiYf/ObJA3/GqulcEEI4Xy
Ng7uysVsBRV61mIEHL2EB1xYmEBEdczEW7TQ9ZT5UkUJvLXMW8ZB57OPlAkc493V
btGblZEO7JPBtM6nDkg/+4msiZYf4xDblsoZe4Y8qNJjLXd4ugp46LPrPeJzJfUU
jLIJFO00cH1st+12Cx31ysthGVlhw1UUZMfSfk6D91iKlV+2vdDT/We00miq9kKg
eWDIgEA+enfy64paws9oeSQ5eb8Zj/mQndg93tpb6nuO+/Oub/igaZRmznXxa83z
QbqYcv0LBCnBLWSVmhWF+iOChiclAf8Q4JWxUPm0Vt+PMldr2Xr7xsa60Xi2H8LM
mSJ5WKHGcxdtOtMu3L9ByYIIcnN8gbFhH+uPD1aJnv5UMKO3qJNjeci4iHsYhOMh
azwuuz1P3IsqHqJlR2BJ5yzkax8L3Aqjaa4fJVBGTxhcuyVPyzPXwnvfvktW5Ch/
8LOXnVssNzM/sVBBG2v4//PWO4Z9Gb/wkS7qqP7Y0b4yrio1bsrbM+swXGa4OEEW
Y/A6AtWMvoB/a26eWgNOnH28YaYEauhXNh7z1tFnva/jUv77if3Zi4QuLdnGZ/xY
laFNugaG0gxkvg5Vhx6HMuHfPU6KjhKdsaEg0l8Cg6Sl/wOwNq3thZ0aX3fOn59R
c/VQT5UP/KYMXSTDINcq0gh8YBbYQR5MoufNj/m9K3mhhzl3fJHK1L8fRO4dC7lD
CKPBdUUdTQif8N57IK7foB8exwdKXwstTeWcp8rnT+Kno3TT2peOPDbA+fbHbClT
zs+oOtaQnnTY/jBQMGwLu9JWFTEMIvvTxVyuOyNiZVr/sSQrP33pGLkTNlHU0aBf
B6gfuNnakAFvub0SoFm4XNYom7mjyH8TrAA5Qdu5DX/VAxvzAok9cSDG+L30JHi+
Hvp+hvCZ9b6AMo+9y5Sfah+9WKXGTlQMTRHZ0wsnxrRsPyz6QhMgLyUyP+rIqYby
MhgIuqJCb1uUSv0mbAKu4yECrp9osZXJuEqWRPgBcx+a3bmx/IlaQ+3iU18h+buU
sT2l/UR9XdEA6yj27pOdem3djBoxpJ/s6qNk0rhPqu/1t/CbSpjTQFM1q7DgZkpw
NrNGLFo1zghLrKpLk4ioHzicJaoP8uRQJAP3tG3lc2I3ZKTAT9TgVDXyIFbU0GrO
LAwV98Kf/W7oNEK1F8IvUS7DCFAwv5HO/mUF2MhhI54E5CgqFsRr10bkhnz183iG
r9V6isYI5sV6/L99SNnXkELZbzIDMAZ7qKd4y7qnvxlbcWNM3+8Ee1VYC/JRijdf
swkiSjw/FgtMTsQRlbBlVNGcyGbjV7Zl3Rf44qQUy6uyNhCAeU68U1B63tl2XjRd
meVWOla8f2I70c96JaCZObrK/+e7IGMKKvAsXje+jJcigA/pGeTk+lnPLb6qapmy
ra+oGqNCSvLYgiekCNaNlD9LiLJIJ+i4kXPK3ffXTwbdqX/Pot6YHrAHrDeRM7/f
uQSj6TKL1tclufmzoj6p1QCTpqA89e0aznuirEjY0GmU9o0DDEbtm5PWgZMdCLvy
LzErgmtxHi4ysR8gQsDOL89EH2AA3LxgdPbWFas9Ui2tMUTN6pcWPBL4YrwiCmmZ
rTHci50uurAMnia0Zq5iIPm/o5+bw5FJRLAN+j7UjF+w1i6ep9+a72wMc/vr0qQS
wlsNCDyXaeTUU6EFKsL5M/duUDOUCCPogtJPetpqeofgmJNivyqN3wcmaAvIFnjC
WhKbnTBOlRht8JOLYbt6z+dKaxOxh6rsLCeYVMLqxs2Ct72x4qgo8kKDfklPSczN
7YH+X0LYZXKUASTNUabyKhInlv0k0EaJo3YHY+WVBI7lf3NEG6W7Bg3T+1FGGO0u
HamYyjiRlyG4UKc2DYY1jvMKtbBVpo7+4kEbEqXVNdiXHG+Qi4uQGRvDx8XZFJeB
ApKKmpNGudKXMwjAKSRPl0R9SZi1ZK8RphRSJvKbpyZxyMg9i+9MFwzwwA7t0j2+
xoMXriFFItSrzUJXXs6cO+TFgqmovS1UFUyU8d390DeatnxGi4eU+xUlVv4nQ9b4
QSvIN6+4/LsHK5TBagn+/5jriJyB5wUIo+71b3jHPoXjSXiKaNVzkKMMxwhJadfn
8wtbc+psrXp0aiKGpdX8zT3pOPzeRPSmVJ0Bcmq9D5RNykQw+4UyXMpxXaDqjVpH
c2hbTJK60XhmCXSgWPLpdhU/8Al/ntBsA8UHd64ATST32m1wWSS4o7431XBdkRvy
6jeGfcMMlFrp70gR12kYTA3PVYKD+ylYrVD/T72UWBHFG9inWMUKDEa0k8W50wTc
i+YzsPPd9JJ21twxfWP9jWkOeVr4VDa+ewNstoATT4LH7Rc5uxNBvPLO/BgE2mlQ
feI6l2y5V9M2Z6pA9fHJCiUxRkoVPUv9Bzz5U4EF+yFymOUl/XDAonMi0Zep8u7X
GQs5aAYbf2pEYMxnsNiHDcdQw8x9eO9SYBzhSLnBx0XOw29+JxmLOXFyeJ6HyqMP
+Ts3jq3Mc20T9Fp92732QWK22t8q0meS0PmP7vYhBRlmWDg3YH6Zk5Xrnl6T9Dgk
bAziZJtqGntpqXKTKVv881tKa9CHHCbV7Eynqiz+aQn0Xbcns25Fg0G5JBO4KbCq
Y2bXwMemz+JCC5a+kRkhTKBLhZju0JXwdeHEfl1GZ//0yGb2hHqvxK+ALgNAjgcB
uiQE3wLPL/2ZMR+Gl4UDJnMFZ1HWbty8fg95sQt5c/oYo8Mcm1q2j/wG3m8nrgGJ
ScOjrVT9PZxi+1Vn9voEEpQDWmTO9Q5w7Fpl6Y01dHJs8VnMZEKt821kM7gBrvge
Ax26jFfK23NnA5GUoa8Q/iCy704PxtKBXYtkfNfn+LKWThTxxRCYaIPwdgqOmixz
6W+g+5ArYUXx0g98YPN9lJpwkCTO7XoyzWnSStFKpFOqUgBIUl93z7s47ihY6/d0
A8SemUQqcwrvKXbfjsLa3rznV0uWwS9Fjzc/fEC1tIlSwSQp8ksc5WrTJ6H858tr
XuTx+136/AfB8Ma6HIIn4WY/glOJLKrFD+qsL6XxOVwAE8Y8eLCq3cvA9gscyLwa
N74l2LNsY9d8fSaf4OroPQVZ/DaTMFvCs5iF8kP3BjRBiJfZQmqtCFTWcosijPxP
/uLFQZmUq3Sogxg3/IVRBFceSo8xlHEgvOTfLIo74AaDBzznPegNq1gcpmyNDvk/
1U/kXiymAZS6AUM/fuH5FhaJ3GnBxg6/rj6Bthr7K5hYozzEpvotE3EnQbslJfHf
OCfNK4LvOOFIE436OdkkT2g78Vg/xtDhpGVT4nulXn8LvueOBaPluTzysnlQ5tVv
5CrjShyRGQXMNddG9RpFUnDiEdgMbXYEMfZqKRyyVyI9UiT6CCymJcjwsu5XgIGG
FmXdCW9r7F0RKrw8NmwydaCYQfFtu1INHrUUq+WV0zAyj2PjNC8/YubN3xaUQvKP
6ZDZ2+oD+xcR/2/qRlF6TEvtY1FMN4s8CbqIYzCPqlHwhFuW8XUsyVhWbLm0oHEU
35CF8Gl/twG6c04vkHxgR6vv3x2i5FPZU64vQ0zex7bhzZ3KeGN13zOBAMhP/f9j
9pMgAY34a2/3O0O+ghc4XG6SDBvVFT/CcuDZMNyfi1QjzX3kG+ZD53L1bhtiT40v
VRThFGT4B7M6pmMSvLoWy/k1C3PoB72QAecY0pcrgIuuP+xLx4WdtDuqi/LYmuN9
db8I0tepZAULge9Ur97ZvnTt+OqcHw9TxlNXNSk9FrQrIP/CEhOLe479I0OjNZwD
hrdWtx5i9uIh+b3xvT5hLkMp25zj7PPB438UM6qUrYh+oMMi/waqpfarFYXJTbfF
xNJAmaHXIx/ZrO8BGnscg3YjhqgrNADLiXQMtsRHBZrg355vom1fnqVD3UmQGk2/
7GAPkMlkcBUGmU4ezyNFpKrsnB0LK1cF0ioqcX//y3x6E6xEXiIG0slxEjxcEzrk
KUn/YUuhZiOEDUPOoL3a77jEoS5vq5AhPi8nSy/brpmLqcZZIYKiyhpGehQgRt/i
DdlfK0gbUV4ggnzVOHRe/RvLMcurIB1bzj+hnW9MxtorCznUzQObwfQM6onPFylj
McxDF400F0ACHuys8kwrem3sD7lXUtC2O7QQdHLKHwxow/MWl0NyyQ45+O6aecSM
kf5psMvHE8g8GjZceOTS/A566bBnNGWdyc4WywDq2G28a7soPEVLbhFhqKah/lxR
9cvR/PMglWtKp/MgrkU3/+vyiShp7Z/tYWN/JECIzfuYX58MdjdRm6tWiodl5amM
ppcWHU0cCUV3kbFwTFstEXMV6tEVowFzEUr/cZvtiGgJs3bJGjAJ60gUob5Nskmx
Km3dJtFmi9MeoN1QJIY80IVY1Gn6jIjsQnagyxkSuKSWVn3Rx/uZygrLcw+9jHn+
zFSnWgHFn+Ilx169xUQ+lfInqktlDw8FTfDGmJYMoH59vCapFhmn63l/GnDCDLBa
LXVxz+B40VKCT1QcFUeuKFPQItGLcy6WAE2XH725lGOmunnSdNBFnUd/LzDPRt+p
eFvm49JtAfoz5C1z72bFb5DTorxZBugCclmxLOJ0bt7D5Ml52weVHKspP/Osg7N4
3fYhRukFPOQyqJL8yAqxbMFvCWECd7AywjBkItfeu7EKYm9dyQpuzrFcaJ4jPU/C
AUUlIFUwkzRKadjL9l0zPLRq69WMm47QxMse6eP3dI4QM75emAHo7PNeSeFutbwA
OGiOSCOYC5LEdZQEHQfvTroi0A0HZvCZsI/d20hYWcoPdeiiQL3X/6kysQwzJ6XV
2OlKcsaUhGLTwe+PWfDJthAWaXrxz0ckkIHrGoWpKeDy0TwT5gnrlZo4NrekUWb/
QG3QwcXBDxskYN3jf4Ow0OMNLVWr2C0hG1Y+lrsMdFkXcnGcNkT67rcnvl/pr+UW
w3Mip2q0xMrwxvWkM0HSa0NX2syPS1ixwZovD4kAlgMHjCpEgJDQjixEo3NyE8Ly
PMU/ORV+onN65lZNkH0PjRSLGYSih1fcNfXGRTa0o5ETqPzwkTAehOtArl8kUuRa
En3OPnKip8J/CYWORnxOtSE/iCdqCBumwvlNfaIp+hfB80n+X/8lnIu6L63CR4R9
vi7HxhvwhelMnmf10o0RIzqGdtNkA5plXktK9mOPe5vTgNgSAstjbQozCI/F7r0K
acLT+wsE7g4qQAM2nHknq+oBL/aXKPRxS7nI3C5MB22SuDa1DA+nfpsacd3P5uv6
Y0cEgs3Sxmx1HZanBzowpAEpTv/+S16K6PYaG9/gLNr4sATKEMTAjYrA6phsMGdm
QxAPTpBoicO1SfJHVkYz2F5yBcN0sqYKRppM+PBMzppSBjqAKWhwKUEUfqLvp4Sa
tNxzF/t/VwDg612UEw15N6vNc/jXg/7EusPMlPiOmuMlRQ+CeEBV30MtGEyO7hhX
FEpI9VliqFqnUUf8AGn1LhODgnnJvg70/kjsuY372giGUBI3WYda+sUqvPgX9QAm
QKywCN9Y2csIPAN/wcXUybey/vZPkulgwmUJuMlMYBDGmIlUGE6hYXiWrfM2KL3U
QaoUVEtPflTJnA6DDeUHpQHT/hW+2YICXWt5jFinOjRPIPyT4Rjgr/JuqwVcpwXB
gzX7zdQUDxM45J3NyvkvjJkV6HPv8ZlWpfWJViFYqrRY5FSFyRakaQLpJ9iRE4I5
753g6xt8NJcm5+/PvFggplIRWrNjwgcIu/7XfRI2nnk0sKoGKTkOcplVlpOY9r1z
H4OPtEEeH6vV3NmCWk8weme/vwKK8xgzrR2Pzjq7BVgDYc+Zwfxr5GCk8QQhJmMJ
Y3ZKFiVus2XgpcUVWQ1sFdEuTZUhp3dFViOJJPusENRBkLPxxCsqRKWy3r5srpJ+
mUwezN+1yOWCCNDR11ijqfuZrS3AshkTrcU6jObiDpEeMuWKA8uPyDqwIT2GBR6N
cV+X9Qha5kQ0r+16QKtyE4jYN74M3PfAAYD/syx26GOLZopZAMVvM5P7WfeggPNM
A6VRS9dhqpYDuzEaK3jd4VdT0bBMIynWJiveaKdQjUNlTHSJTHFgy9D4Lk3lHjHJ
Ise1qxpPb+EFIE7/+25o0tz9AkQRI9W/lojeebLzozLvWRmHm5eQc4rjQvPXter5
RZlowN7st00IpNyiCqChTL1wSBEmWk19MAPpzDFUnD+BAXKUYfw/k2No02a5Q+0S
IyYqdypIGuJlOCCt6DLTUkyw9uTzTdZYbrHpTULGPE2T9YXnR4sWFiacs4HMfE7w
+Jvvo+5yhgre4mXnEMmLfrWTpF1t8thiXDTeVhXVitmqriH4d8q80MiPuG0FHNiZ
s3OCHVtN1kYAbwaq+TCsKTKDuBfrKV8iRH/3vINqX91Ahq1C9FDAtWqf6tWZTqtG
hRj3KlIL61gYrtm+qnfAmGnWqrS4IPfUAGY/8qKtWtc0RRc93ZX7IWFGwvbqAaT/
e4bogoUxjFaNPJPA+l42J6YblzzjuBK7k4/UlrcmEdESj5I+4NshxDzCgk81mqV3
rBXCC5UI4asz4/lK2J3mZW7ac3l02hZzs2tA3TtNEyPfkWQxo1rioFNMMTUg3y/f
wgcSQvoT1ueTfARwZqKolODsf3Kc8PGY0NqdHgjY8UFEgUvU430hPVdc2DLR5ihn
PLnjMYs0m2E3xuw6rzZ3N21Au9aEl19laxdPJVJ8zRUo5vRgR6zEzcAj9oWFkgAk
ftR90C4yX4SESks8mDmir43Xww5oJlF7Lh31my9JMhNKNNvcW/A8n8zjlE4/846y
PcnSM5dm7FXtGJXHvTg1ZTPB1p2GErff4TXZr64ik5wNS2Y3G1bsM+IrS3C2rLgP
K/uomprwtSuXjx9BecQ2aEsJW5xCbecSZtSkgfT28UpLet49yOho15cYJSpEipry
1VMBVBet7wFM6ANQLwj23LVbTCbmP3CCluKCGPlaS5u736H37xFo5/hDyxnAhVC/
vcdIPhrhX1Pl5bprirdB0TMHAk3vE1vCp4CB68u2p5cPPx6W3W1Kf8fBba0pRECq
kc3nKgcJiVj5xbciaNXgISXXCPcZLCWNL3b6VlEO/Wee9oBXnr/bIIE4yVheu1p7
hG+9yiirBdv8yXb3JvAbig9IubsMAZfR4cusYjG0uJ/me6sSHzj0VzpYZ23h8YGY
y4TKM07usHABOTIzy2rp3s5yYcS4VXGVcBZhyxKTPWMPYUGR0ythO45HH+nlQe/0
jhnuNiM/yryuzqItoEcElR7JIYqLd1rkT0HsByrRJfowbfZXB7KZQyC7hcppn+Vr
AZIfGx+rpsyLt4V3uAigGsF2ZI7KA7G/2YT9zSRpnLSuSZfci/EC2bltrfteMsUv
b2cyOFdTlmpzEW/95cKnUxLOm0RpypqEDWIGiVb00ERzNd7OE1qeRVPCirWAcElX
g82pQBaey+FoN/BtftVafdq2DZ1PoRJu4L6vLHbFFFvS24KoOPYUoTLWbLa8W8pA
ilRMmJBK8H+zozwr5zBRh5b0kp30JmKzcIhr4sGCw5qukxe89uDOLqMFWHttWQLi
8N98GRYre53rVrQX1IpsvxRY16u+abIyjzb16DT05tjiSj5XSX220UtMLWQEo/hm
brT20D9f9dDCwUy0c/z3fjzRTyx5waP55A646HCKa6ucQekgyS8jiU9rucuRA/Qy
Gjvp7fBM4LAIlPocEWbyU03P/URC0Tbv/K2/OKeLkZi3hkzgiX0vMheQhhdOEpq4
9y2istHzM4y2+h8NA67TV3Skiy4SmNo+sQuQbZ/EEhM4cUbMsjJUd0xMLUKQb/lo
mYsUREgmAR+LIO8JYzt5R3Bc8db5Fs6MVHuJ9rJZpgVsMxIr4RYJPVxMuBQL+vCf
5p5AhQWHuTMJS0WvTzU41A+07ZnHIcBk+kz95ziBVPcLi6ej2OPNZBRZSmUsLycR
H+A6fOZ9GQ7bkXj4J1INGW6XCKmIBag5urriz1PxycYV9nYNM/p7U3GTK0I/HwFS
Lu+lstg9OhTg2LGipDriXiVcYK11yW/cWBaBEhrODR/jlv/T/KgPgsFK65cPwHmd
U1AHrddHtInzcIIqHwcJGRipvc1pqPn+gYEQuvD7wtHbqrh52VFikZFzEpgx85qJ
2LCuufUrG5Vev4yHmX3PA5zHkaItUsP0ZaBlUcukbW2jQq2ctJ7/d4jPKWMYexgX
4k+CJER/zC2UzE6JSgqFLoccFetUcN5Q7G6gFh/64f7fxXp6YCnniGjhQbW5GZeQ
ByXD39xGINhHVla8mj7Sl7y9RLlklLgZ/spyyC3Ct7wVpubGC9/oX87zTL01oWEb
5vElaylhknBLvOp5DvW9ZCL3eIDoksKY+94SlIv/RMfm+CLeTpq24oCGtmO+mhu4
4RNMfpVfCzFgJa3n+MdHNiEUXIkxuiZ70OO8jnOJHOZrcxAlPaIyxVZ9HmIdDcoR
VD8DstPvP6jlmZbh6lfhu29eChZHIY4c+FZvyI3e8d0c0o6DssbpNpMCFB1rECjv
s6t094Xitcuuh7UHVI3HQzhHXBCEWPu8jsdczemjo2ejg7unLvio6HLelbNBtJTv
T6+tK00d79OhlGtQbn4ptL3VElsnjAzhX7h2PUFdF3LJmZyCrD3SmpVU/NBtdJFW
9xAm/M3eJiRrpigIsvugi2BIE7w21yTYlEwyXQk1OZrlPxZzPbU1Dahl0axMBy+I
DCN8ee3pKjXrn2/OctCPysGxlNUPXKV1dvHqbcyP9j5KKnw8h6qvmGPGRuaZMJcf
8QJygSvZC0YAP+Ee+YCudN/YM8iFNssfTiK4fGRKfP1mBJkInYFl+vymwNxnrT8J
X7lBPsWJl8I2o98EQHPcjimvNPONU83j6d6/xq7WBSgQV9MbHlT1YNHSHrVDUJ8T
359Cb64ykyMyfwybdQX0ACeAuorQDFo8I25M3W6P2+2CbLFhPK9smAlLLTzInM+D
g1jiyG8JHoyq+R1vhyxahBonxYr29pwpM7AYlw6hYjzpiQuj/bU+pwDepyJcSyT0
C/k5Vfo2r4EWQQnktzfJCyeetwCUxM93Npr3n57gDavAYaSvgdHTPTc6O1qVPN16
4WAB6D8H1wknCZIhYXb5KfMAG5WAIiXG9IhJOyqTecdPU6MPtw/8JFxxBN2FwijI
4z5nSD6fjDmnLTAAjM4z3k9ZTqVrl1h5ivQZk6UBLpJQ4xrK5TCaJ7qcGfX9IyRR
eiWn33twBlaeTedv0ps+RIgBpmGlKDKgxWzL8CvgK+xxC9SwZPZJBuNalo0pJzfd
2h6oFunjxZx6HN2jy25Kiag9iAUfHnL1wje5eFDeoqQKHxqbsRE685JkCZtdCV8o
Hig/5trIB+tfbHSuLc3it748YLKtBo8CwrbJiXpybm08Nql/GWbyk6l6o+zPh//L
031LriyyldRyGa2JMQfXEjvf6gfSWynb+PySeAnqmnicHxCDCwhjI44O2Mi/dvmv
F/d7e2qonLAPGfribFdWXEU0YoIeRntmlDxmRDK7fvB8Db9P+Vp+Ff3aaFYyPbuI
wZaQpqud/ZTouYub+Xc1Q0p/t/89iNMpF0go430nBBrwIHY+dB3qjW2304Rmpiig
Z9a6ggNKORCdp67ZYNVEmbGxMCMlM7D/UGpyfv9ebKTaZgEuw0IM08C1YC4f5vKt
Ej8/CToWGrVn+oMWAopALKGLxsgU9lml1znzb7IFuS4bXb1fRKHE8E4hjqzBJxN8
lrVnRZGZFxmyZNLgEPc9yyYjx9jVIZqoF+LtXbJ1j0Jsdo5dOmZ+o35a17dqoKUt
fBb7NfLaMv+6SX20i+9UzpfywENC/Of5F0TwqFcftMrhVAbf7YOSYBZcOx+tLEvx
bSCBatIn0sGODKDcCvxfRNStP14q34W6xEuKWNoKoVWowtwsDnqnkrJ3s+c3u8xZ
KbvMpFQ8YoU6RgC0pWnh4g7y67pvx/jJZ5ERJCujj/DG99PJNDTdxkoil+VK8SUV
dMMIiUd8Z1hIWUDWl+1I8O6jXUIsdMUwa44cMaeHCn0RnKOSFUmSpLczijyZohZz
N57xieA9slr8Hhw+b3l0W3EqUQpXRfNquHJpDekYGT1sqXFQm41Zvktaf62DXYbY
hJL2Te12RLiBJtSV0443eAdXkm6ook+BfVIopC87XYFt7evwKJrnXsxyrVqYlpcp
9LOjD0wbUHj31cwyFcSO5ZcsF8t6tvt4qx3cD0ERkGTy7EmKNdlil8r1CMBh2k3g
H7K3U61O1zxvcaVXh4BMagEQGIEEZA3RZqbbFF12Gqf03aFsT1PbxoTYd9tFIFbI
ckDq3Z41nFvnvlzwWn5gdoVyqb3I2/SGpzwT7GaP6BPot0IJ3kSj2ny7Snxs6XVS
yg92+8ILicpIwuGET70J5g0dK+6+2TBUywDCtIipeSkKA9FfeIxQoHwqUBVaPEbQ
vk6MjvZh79OWjYv9bM0t/DdmcwAqQhrA+J5iOoFpMwcohbv7IbFmYxWfvi3/4gTI
mKYo4wN4UCmNiuZKBmpYrG5dA2o844QgrLEQnWbDUk7IpNmZUQl7c0WZB7Xr6c5g
6LQ3Z7V21/AgshBxSzVfV6Zniw/K2DiBpjAdAYgVoboRkV795qFljpI5+xDMuED7
TwXBC6e+53QDd4/mu1JYv5DnbYnTugrA20KulwFyfkxKnG/Fg3wpbRocoBeHnNtl
Bh+CPVirzJld0TdwOuDgnNNcN+9YBk9iPXmrnfp/nNh6Jd/dQT31oYrwevjDWKlZ
FdpxqpwTYYW+y9W+JkXHpTce5eCiosdTGo7OfIW0g+8NDzwi0j1A30+hl5dW5ljn
gFlIlKPtjwdOF6p/JpufSmZtZ8/S6VjHlJtnriEuWYYc0WZPXDGDEN0u8vH0lu3f
3UbYotmD7FLTZQqLoUHzVcW39o8gimTnE63oi5aBZbrjMBOgGmVUtibAhYo2AcnR
OuLT1AFISz3Tp9yFUro2V0rqRopwExeu9hKefbrhf68SMXoOtYH6Klw5VqA3R4aR
XJT3pHjskaMAaRvtijhX3Y6SsgeAGXqmTnifRNFfpl1eTHhhnfmUMoUS4n7yvJq7
29xjTZcd7+LsvrIvu2Xfvfg4UrfTnJ1FuGdiuufMtQTAPdqg5E3ErcjT5Ch5V/C7
qX5brnOv+x+STGpoC0Bv7FEfw8FBK8LDQ/p9ayK78BFqhddThHAP2/U1W+5wqq26
uxPFqYGpWXF13Z7fg8EwwVCTyTfta9pASsTafaiJ4Cw3gXz6YA3N4LiIRoP0fNYF
gc+LCnB3W1+Kn8xBVnk2j3cVHtYY4dIWCbK/dCwP667KTIdk/cfw8K7qws6/Rskw
csUJJiac/p0Q11Y28UKK67j/FI19weiwX0wrKT1yMFPJJZJhvyE/BmVd0/s2zSsc
b1kGCHWDkmECl77ccbmgXFHbr8dXyZXeTBDnpQyPP/lMICD2RmUefjsbtNIP7skG
ZsCWCq+fVfN801Y3SZIV5ccr39vIQVTCEeHYiesZasOZVlzTJbDsPfEzcgy7t4jR
GMbfBEbw1k2MeDg22vSuTUxDC3MWsrkFHItT8oL3gkeXeKZl4ON1wDRYJjiLET8j
+yWv+6A+OpPeurHrVBEseBfjDiXQiM3GptwLbpE0k4A2HpiMhD4hUBsJhyx0AGdD
W1HLVvLGooisQXVSc7unIfIkRe7fzEHgQkXt/O5+VD4/2efzNyW3g8K/QRTsHlXA
gwXfgTvqUtQ2AqBycXEdBhotmIvKHQfWhQRYC2ggQBRh0y5F2/urgHysubt15Buw
uF1saR++9EaARcdug/xJbFTDJ1edKas3IUaNHn8DSd0ps3PpsSc16yrmDJwTiZtr
QpGQpnDWlG/Y5L4T7SqehSyFDKK6hPywofnGF3/7l4vyUWegJH5aOkBivpLwDLP5
PPUllBmobonYxWolrfVFYiKPOiBsBSj2aFd8DcjEPU7LGb1EQ/XrksDCmpC7ehlM
r0cqWtXLvCYCNxhGVWx3Y8medeM9imxuQK++uZlaz43PE91jCDOcTDDwEEQXkHZt
PI2ZSlX2Xyxz+H+JJJCZDX4wGf5vsl3onqQKyMys1GWKOXXdXCrlyfzUEurHKvlw
pjdtWrXzfPxn4ivTPsaWgfAd1Wyn+iQLMNYxQGqpb0TVlL3Fk9Q8ql4bGrvLhfgx
fCQTX9LfmadcXVB4zf53TpNDEBe2Fst0fl2zDkTvk/pcGJ4ZLcEIgfNttvSBmVA0
8wCvxATyyGoDT9sH6J7TqEN5v0V6FPjvBhLS5kbjbCnTz0/xJnrBe4U4wt3UK527
96e8jjfkEC1gLewHy2MVfCGidkUvRx7ON8KDuqnoOOo3YSftTtcHQ31RvF/QPDDp
VEQt+negtu6mnE/XC9PsLZn5v5XHGS9ePqRLth+Xw5oGiwj0QEiZO0j3eD5eoVcC
opxPXT4/4RYve9WNwxTa/lb4XyJOCEuLZlaheex6GcrmsyC490MueVjADJb52cMU
eIgKRTpJIhpzDKxJuHHSB/Hy6HBl4uPENAn3kYld5/KII5sfXg5pwsmag1dvjlUf
yTFicA3pNiQ4ABVYAEkPcWsriuBxcRlXna4YB+avbB8xkCFcXgStHtdJ53dItkh3
sYww/Bi5RJp7F4hlFsR7tFfQWRA4sk0r+lrPeYRMSIQniMvY18Q6zezfJVLqbC7+
v/BAmUxOTHBUgCV+cTPU6eIIPAwhwmYv8ujs4Av5tsG2nCCLlBnDE33xS03CXV5r
POlrta2AqsM1Ls0A+Kkbomy3aUXBF7kHe0y47Gdtd/nwfbdXEwN87DRxjdTw6rIA
nBIc51ODAYjejnJZrr8ljHNdRCCHQYdpsCyVJ9kQj971YWpr2ine6jj9nDEFo08r
PirB0tAxRyC6nscoO4slGYm2oiZ9qBBDPPtRDmzlVLOAZmATV0Fdgar/M9GqH6NM
1/p9Y5tlGIis4yGDW6Xgn+FFS+CLQn4Hpi/IMQUuidQMnyv87Bt+QJGwfEL+O1wk
aU/097n3/pbrtam3JYE4fAY4wYe0Ug2qle1JhdqH6I85lRwKeEd8tI7ZE13nYWA5
VDwUp+WRnzvcEfeq9gPbRXXfZN/etbmCsh6rI/0JuS0VKxw6vgDkAVEbKVPqLoLB
n6UMTSKYDu9CCPsZzyV0hcoXqO8F6Nj9/M4Aa9U862rkfZ6HMVECCqQ+CzwAJgs3
RBoyoVKUew5AWbqSbWFn00uceHNJ/C/USuYoiYE8+ZdW4PXla8HuyPCJKheW4ksB
ZZD/VeliSnuGC8bBHYvgLlQBZiyf3/n82CuyTR4tsox4wkannv6zDQwO7r4oKLdy
2UWwlKzd9s9bA4NhuTreTAIBTzc7GCaM42XRt0fvWvL4CSpa5v5gf7waqCn4tA7g
2nXG5eB1L1UVrOaClZ+xa3pt9EE/PKNVHwwJvstPh9mUA/RhthCeRKRCy/+hFJeJ
roVhQpH6rAW/N55vumJuw+GPWlNIl016IRZPM/w5Ur/pZ0xkrlVzcZlcSM5NoHRo
JgeS2DGOtt17gD0GdbyCjB69RZh9FgBTtsWnLiz97Q2LI9HWOJYkMWRcKERZEu14
wlBTtwgJp26DXumvyPKRL8EwKjQaC6H/MIqO6SKaYuD1uSzRee1UfycWzyTh6+qe
E0KX2Z8fzWD1w9f379N55k2BC+s64yX7HVJo1Fqvyu1VHwFspqIkveybXc7ttYtz
T8lC3sMXLuWOPbEh5cKhz3u6Zr5a3H8YKgvdSmbPdy6fe5GCdXkVISIQg03B04s3
U3t9K966tE1cCgApGj7p4Xk6iakz90F9vgS27yOgXS7JeOaJxZIe12fMW/Op+GCu
gT17m9bo1tVO4tzRKm5VwlEuPaY5BU4plXh644IPxalAi04CdVwmtJHsJ5YtHTB6
wm/q8KRKTZE9ep1zY6fD/8y0EhEyteZdIbE4tAlMygcrT2nrUHFHgUPKIdkDNgVi
quEjXPnBQA5IwNRTYJV/AYyTcBG8iT6ICZvUCeqYLtZBw+L7wQow7r6j+m3Lkwtg
UrRcMFtJ1CxhuaaiP1zUpvfpmIbLiWySOzbAaiJXInfI5rQtSJx7NIx5BMckpsyJ
6IKsrU0dBKw2L2KXKRpPedm0I2Vsx8eIX59mLLMg6e01gX8siwQ2F1rYZ38mowZb
1+Dw0pGcBXRnmfgnZjKT0qypu2TPcQwp2C6mwfhqczaXMZY/b0iLtmccmhR1I8aK
SLf+tCLSYbty3AGi5GqwKbA8tXDWyE3aUszPd41R8JwMJWYVc6Wx5pfDGCkOr9/0
UET9+nvLsl8EaN79uKcx1wJmF+9UMQZi18lFqPUkw4zzdfehPMCXfOMvqi1cqPB/
avKfBiHy/ztEspr76samZBnNNhBiXyZLIgyywzUi7kYNseGF9M1md2bdShmfWl+1
VGwB1Gv9XUD9n7xnA5vBOBp4KO9lU6JJcHxQy4cwR6PyGRRuAFvVS6r4JbBNw4l3
/CT9DmE3XcAwvU9Bgp82cuDc3LA0hUSUzXPI83nfKMPUtjXl5p0Tbl96iGjRSpGT
G7oeYMsMmSlNYthj+O7Cx7nNsOukFkkT54ld8cAoKg1gv+Z6q9aGCNl4s3J2vZrC
0CAn23jxUr9fqi83ONYfdCNxA4guowAYJDAPmKSIrFqlUjJv/w3PiL68aM8yYEpm
gLx6qPJQXLZHeLci8WQECQARylMvogJGWVkrgOSAllu4vtnN+8VNfwM5lax2ZXYw
TCzEIIay1j5HkOLB9mWVBHcVWxopYoc//wBys9+8wvgjmNDbE7Xq6xBgJ/0IRae+
23toQD4VssB02RYdDMQfW9xgB4FEbqziz+cLmcWTad+jAFekGM4bg7Hdyx8WC3sV
E9lMyVH5S5C9IWLeTa2a2lEyvo3UZre/2Ze5HUzH75m8i8BgWxCBZLhJwhhbB3ih
YFafHCyFakNQG4qk9OxZiWC0SnM9l6hkhrlHask0aTdWBc7fObgCFeLCnK8m40SG
sND7fF2+ScroskjmZ7I/SGyc7hS9cwTAOh5pe7j0tacExgi/Fs2yHI0BKAoyHBTT
0j9rPq2WAOIu4e0i6589jjsk6WbG9ak++Loju3cCami+gIFFcMGbvxYERw5jalgJ
BgVYxYdG9kzembhZlP97UL70CyhYE8l603p+z/aMd/l1ltPZDqyIGRnL6/VPPs3M
Q1eMr5w+eh9hr07w5wl76ziBvj3rvmSk+r3sFe5P7wc76MJkXtvGsbkMtCd0G52t
LpYKwICRYDwaSQYQ4ppunJXVigxV3AgUtJMpccAebvsbQ4JoT/hW4rvSbk4uORDf
VdRKMnnMeaaG8vKJs3Wo6oG6GX5b4D3j6bqfgMIZXR/5cB1jV5/mxrKYjmPVdXTv
3TogXBdSiE1IvHIf13FC117RmlmNH2lAPr2zyhF7hv1szdU+F7fYIIPEEk+e5Q0t
oUkZIowQJwWW42OKT/EpZYwQdcFnbAJQGbDrAkKlLmDEHPGLybbP1JFZBm5ywh8L
Ywek3YwFwObQ6nF55WPhEOp1OT6cxdQYs1erPqW+sZMwfTc5q8KCKhIat4rVhhEY
7kwMO/3QhxTTYGKkJ1CZMaa6F/cd4yiL9Xf6XMVzFDYoSeyv/Mee+pz83van0uiI
8qC1JBdJHZA7N2Ym0dWCwIW9Bfng2fY+NUAFLW3aixMnqkHENkIe6E9kCXk/lbuw
APOZK3kq2IHy+XnoAeGEzmgXEMNHCbvRI4l0vwUbg7SRyDgkGSKhg8oikrpUNdFT
eU8bNyPBy/NDELtPgc5a3Bj80dL3WRc3awdaqBushhhh1ZM+ZFs2Son/8m8TKq3e
9J+XQurM/1QlWIQ7RJn2LJQKnQ5aSapD/1dkZ9g08WQoLLDT91oB6r5JyQhJZOc9
2sBfsi45hE9C/jN/7xcq5SprIp83e56yw94hk85mIMIbsjoRAL1DUDtczF6wWYKO
rtj/H49LPAz/BmIJQYtVig6kHa/COCSHAUT9TArdU1JolW2UKI8DAzbAEUJUmzy6
c3sp/SFbsb4qqnMAGrqzgoWl2/SfuQuHRaC7cPva0rWeU5skuYorn7Q3bKzUvQCS
TxwB1abDVBSJ6kCs9fRhloZeIIYEyJXlQFKyE2z5LnU1165Db/RKyCRyH4ThGSC3
cJbOvhzAT7NxzpeUuwqmuFO2QiOhch83M3gkxQPEE8SIfYNwSP+XlcmDGBN6bxDY
wq1HDBP3DNd4maC3enU4vz7yYHkJ49zJMTEk6WBzzRWNUT447CcPHZtYKd+1yhBW
N0VTVzWmVSwmzNen+8d/HJSF+80TySUfC9Deq1/G1+NJmeNQp5PymfvjAFc1yQCz
sU2GdeBEDldEo/CaA4+8vNg+NXkmu4/WPUdqKkVNH/KHHwqTF09/GFC2bABbwqqC
egJZ5eg2EibwJhGpETfxvUV38INtFVT/WfKYVLEpJv7YVKAyExPMH3b8B3tseQKD
c51PVneqjaSambCHvtuCgDENJFj8SfZTki5dsie01J5e9RxBf7TyPxRbYuCqVYwY
S8jTewDGzhfNTdgvpSZ5JbDgvouyw80ztd2mWMFL/ZZ8trSQVWVG5r//5enlR64T
sHuPNJ15OcJqFd4Nnp33+/M3HVqoFXp4qydGD3q/HlRpCn5Jhcx1d12QooX0WoY3
U6CAqwAfNVgWdzBz4VFu8PrcYQdf5cxZ8wXYZ5TVoYVnyOIJ4g4FVxTivjVEt6ww
DuodMbxIBt+I9+jpB5nW67ZMW0ipoCFHxWn9wXkfxanZvomUDiv4wKJCaGJCplmr
5cDAbGVB7vCGGtYZvEFhJa+o0xVihMiqnV9jUlozL3Myw688g6+dxHzOHqaSZO6+
0JQnMil1iQTyIFHT0Qz0FDdxJui2ZqsswHUrDeRkYvqaxT42JyW6HxTneI16RNE3
WEaMCgIRzbeTjK8tMpUfCssHvX3dMnODYiufEjSEym4qrG2tiL5Y5v5FS9mqDmHL
jA/mUou3D1y4/T5wiP/q+Tyhylae/OAJhfqlCb6qkwR1GBk+k8sOg22iCGJ7PzK8
uXArHV36NCw+dPsoZdNgOBUAyHNyea4NIZbr/6P9L+/9PBNcGPfNbJUr2vSDvCP8
RAE+mwrCdVjRXrqTYhFMT7vFZ0cst9/0cp/VKH2RLi3x0GM2oXr5FJm11YkiytY8
XWhnF2eDFb/e7FwHBgf0TdAGug6qr4d7nO5snxEAXb20j8REu0M0si+gFfSJdX5A
uj//05eZRH4TWgpT2hPHBiaUn2DwElknPOa8hexK3Fee4gcUpo7+h9XZ0rgf2azw
euO615Qt2/84N7PoYlSwKpHRWt+xxbK/9w6CpkeIIgvQN2YUxXDujRwiCVMjT4h9
UsOyCm62AO1jOq/U33YhGXJW19ejXnHOkA2mho9OcbqGpU6Xk+CS2GXz5anLPFyF
AQEmaaVeovLs6aaYGWZNXGmMa4aHMPNl3OU7AJ7cCSS/4O/M2R0USr4gXhD31emV
Yt+fYFtsH3yjmeSJMq9NgUkCEtVk5bNCxHxCqK320C2WGVtHu6w+75WdzigUjVYU
NW73XiGDQAoNdL4hW66bICuI/YTUvEcIUnzZvk02KEXgB+KgkYi46+LkYrXBhYiY
zvVY6xTKgTZ3+mvySsSVb6ri5bYjc9bXELFYL2S3KK2E6+VRIfYtA8K1oRR9ufu1
sNnZx3ce4zc3wVWjGaedj2ZK3TS4rlJ7QSeHzznmCnv+npKw2yL8uIXyALlQ7x9A
bdZSYRU6+StXEfmlcVMJSixA6v6ljrdpOhrXsHi6zs/sgsoSAEm4o76/oO30Q+gv
+TctdaX/6KjXUKvNgFNxpiDi9QLt17jSSO4ofJt8wgqRInhjHBqbzFcjZzWV5Qxo
PNe2mbAPxFx3gXoWzrTFKVltyp2eaVI6PTFqia+GGdVe2xErYj6OcE+omD4ST7on
bOpppVp9XYb32qUJTxpS+Tlxvn7DDpRBC/e3UTl+fAxA9v+/KXiU4cfVo2v2YFTM
Uk477d4/mtAGvp55mOtq9WjnEvavnRqW2WZdMFGmMuKfKnU/EFdIDwBzjElwbzmU
DyuE2nIM84J7+ZlCZ7PsFB7bQUOHdTbQR9mGRrKptNMZLAL9Rq0Wg3PGYKwA3ysd
EZXPhDIs9wGd2yZC5dF1kbscF7pZ9mXS+RLRtWvjBtMNsF1iC+MI20ahzqJDbjsZ
tW1KQOrONat+gKIIe3atQjZHh0qq9LOLppqIV/SK+U02AUG3MMIYPakyHklMH3T+
qQDNVAR1uIdW3LlwnjGs51TMkIs3nEYAG9glVkKLojRf2TqM1bZiBqiMlh29Jm/d
yiR1HiaUnFkI9VNcTb4K42gRfxiUVtpsum66eeUFSyqL5iHGX5UU1p+ywsKMcq26
y+ih5vM6yHs0AAE+KUT3P4a/D8Wu1RXv1rMRT7AIQvh41vpVKknTk6AkEaWN6rEL
RpZ8UBfR5PIRNrx1VjGO57dYsvA9k0A09gvEcXJRD7AKC1U7zmd3GYAVrLQnFHGq
g7hbISuWM7Zvy/WIBFqKHBcaKEAguke2qQBAUJ/Z4ehxBufl52eb4mYmd39XRmyf
Uv6hSfRIhPazw13aeorpRnOS+39zbIoU0tXCbOebhkK1CrqWbjCcaWbb/MBvo6FU
w/P2eqHKeOgLv99pJ8jcfj6zrcG4FtwbpTgTVdu36lhCF/CMTvVamV7mgt/75SpX
yedtBRUifM/KDnpX9o7qU8x1vI+WHgFJ8DbqbeO6NoaxkdgqVESy+Lfg15k0PYFc
P/zSpqGyj2bVdcRZFUqdwPGmAO9yGstgVhRn3oH+6bAyJrE+cAcouW0I+MgDrj3n
tjX5jMQXiYwBTkGFCpKcdZtt6uK9cn/F4Su+Q9jzdLan5kBqkxe3UHUSBjd0cFlb
FtYXWNAQO9VQo2/ZGUUUgkPIw8V6T14UQ0MBKyEcGEKLB894lK5kG9NKJNpoMUuQ
UR9WoKnVE91/yewjjdXO1rkQInYFvOR0f47vcQHn+83GFt2x+MyHa5bP2bRcvuOc
YDzpIj9QKs3kL+7+owuMiQHgKJy4jc1HMRyC1huJ/aCDwOhs2E9gt7F7OOvL3JdD
1ZP6ys2hZxousjBF3hGZQgBG8g3gH5dIKi0NthH8oxdvmUIH5EShmcVhvqyohXaH
VLxvEoPomDgGnRMEdYZjVGnUlLCyKGqMtgF5xnRW1EXQEVKhjRPgdUWbojVFIPZ0
jw1Sgda1EkyUTheB/G7oOOuNKp7hN1vBheWZwPSZc/I+F1UKUm4P7Ibpm0VqGFLd
ifzgwEwXjCEDpSnf+hHzkgF3LFd7zwCwRF6klpkKM/Lovrk/eL07tYGvMFZ1bSa8
N5PWDlyIJsxf21bJENXhMaL85Mt4ZNa26KNFeDyiePsk6+ncuc4eoKL3ckkY7G0/
lBTyjjuvByPsPQTioWyo7GbsqyUCHalwJB1QuEF4SdxXsdnLGjhE6mSiluZ5rY8q
P/SyXt7knZiVb8aMgyrRP/1vF2PqBUh1HD/9hrFGOe6eB4DBb4N/36q27DWKG14W
7wPJrAobD0wZE2+zgmLxSWVbjEb6mZZ23rPl7TS0/uTwhCkK+HQ7FdyDajNZJtVP
155KxD3UAPaNUBP1B6JVNFtUq3NX8mrdZ5h1LsIek04oHHAhqWOpHaXhQ1NL4rn7
zDCJlIRefnG+UWOHTtMw1qcz1ZfxAXPUirT4HNU41R+Kr3Ip9pRRL6LDOwKIWMNP
UzUY9pXEs5aiUAuNjFc4Ab4qBvmiDGugmlORUbr5KbZZ1X+//8cRAc7uVfqNSC5+
Dp03Nv8/IWd61+duVdtOHeTcZ2LH24RkHgXymX2Nz7FrnBnTSYe8GF+fNRCYzRBE
FIDsrEL5jbRR+LSP6MnEJFgyW4aWN1NSdfCmtTO6ZrYcKfvs6ObA7w96Rv654PQL
XqKt6qhs0iL6dpSDGtYVua/6KwA/Terwq344vndG59loiI5ooRV9ykzeLnTK1p9a
QVriUZQznLUmwygjT3vYq6dkbktgjNAwP9phkOClWa6O2hKC9O2YjB6PHjObLMco
HDCFAsI991/F+C1fsAeQUeBVt1YKPscil+3eHF3aTX3qqOk6GEtGaFVLqbPDN357
35ATCHk8ycLYNmEhKoibvr9/Tpxmru0VSPtRgN+myuvjJc1UkSJEhphNT481cPZI
gwibxKlHuMyKaB5QlA3eOs++DvgqDk7UnyEdgExlO//6q8sYrPxQ3LnQIvwtSsw1
sk3VLOtO4lWffGQAva4qwfA1vQUUPpgqaitUsSbexZnONAfu9odm86D05ji+piWT
ClL1g0VusN+cf49ccYHjilzxR/vm1snjKapiVv/DDa++Xn+JQ9AXx+pmzvfW/abq
w8zWy4aS7gwqf6685MgA9i/bDzOkL/tEyZgepHEo8oHk3sG984YX0/PpqrR+C7sQ
PXHrYHTJ/hrSYF2EcAmNBuYIVEv1/NJePpbE7hAThMRcuV00bJ3sEA5Hz4DYt9qI
+JZlr4PRRTYvZzZ1IRyWn+FlTW4mvmtgHpUigmWEF0G3XauWtVIk9BNiCIV0uHiz
yWyRuIXv3hfmm5JakBPoHGsVWLPLAXXvl+lIwGaetJcyxO34LIaAJiX1GFE4iRJC
HvmsxCN7uVMkhVNb9l49JGXs1mNpql3DYMo2tIIUiKXcsD/pCgFGQJwKb/vKCdEe
Rl5dV+Bgp7MH+J6dMxzQKJO0jRUQrZTMbG/gVB6EVz0/z1lfmJMahhkPwf0wS1IA
IbT2Qj/ET7yC4tKQU6Tg/2GZquZSfcpfUNH+vtOngtJ/l1nhZWX1YVJJ5KAU5xRq
4bQ7wTVXcefoj/8Dh4RIPDiL2jQdiRdyL4Jxh+MjsBORpyIiMXLyk7tT4QC/C/Mb
vUpXyEmtNTGFTPhm3twdSjaGL4pbxfwPR2RKtf477HUku5M6VDDqKaP0iIG/9oXV
wswO82BFeGMmP2iMQkEpFhumAPdn2NyjSST6czCXOoziZe3WNKEAw0CG/1Foq0jJ
1QvTQ10DEIBDmVjaTsMCy5chaor6d9Qh3jUfEIEEyw+LjJlT2Jp1GGM4K1cEO3Mz
6+9/l9YufDDc/oAG3+EaCbtZnWlU+lE4FWTdby03T/KRefxgwnDB7sHLQMG2aCSn
YqMCcxc68O6rRx3jagdWaYLpaAK2eooZXAWvVG4YEIsd7fMs2BSklizMeRRB8e7I
A5p+zuR1gtlOGWSZYfV28ki8MDf6xRl/QpZRZCQarUD4ikA3qaWzdOtb59xWnMvZ
gRZoio+owLJl1OG74AhQ2lXHYSWrhL0NVVme257Q6iyQk7CIiR5v0vSC6RCrJ5DE
NIdq8I/ZxvGJg01dLd1OL+5SmwG4jNTm8z+LONwM9X5yG7O0QgW9CaTybMwXNgjO
foJeP8ha7AHjsUyNyrr/0TJ98y/bFkw9e9KeCjx2LVm4ChLA1X6siWnIzW7JJQzB
24mYhjaWUilZHrnUG86c1IzBluS4BYV1KAzw43sN8NWRhpo2Xu/Utbt9TYGmie6i
SJk7/wJGhKTlkG3iAmVfRzXV7BrAoVx5dVTjg5CNo9MCDVRwBLPQg18DQvIgB4o2
AFQmpmasWTBmfLSj68L8YEuQpoFPyDZcQCzsGRNvqR958QNyk8NKkMrY5l11ASwm
YPSgD3GcKYxL3VshjtWkFU/t4Zo9TR/Lg9On0ByR+6LwsmhoP5oIuJxpLDlodbhz
I5ByUVGUGfXiJSMhtOnR5Ewmj/BVVtg+uAj2fvoD2gUoS4j8phHa51scO3hhIr2s
IXkHTv04+4EPW2o1PSzfRrNCwyTz1Zw5qHiuHfV+oTnewVhZvd+AiDl+Bb8NjV4Y
eEJvTSrKmoWbGuZ6ksVpWbAgUpf0QskSOv4Pv4NnvwC0qu8b4YapBSC6qxDLJUJl
1i3FLeFdnC44HngkdP5lU5B5xjtK7M+XLEiRvoH/Okcn/0LETfNw8MUBr7j/C9Ww
w4+MiHzIFqoEg48w68K6dpn9ecgXytJC+8A/ZHF68efE35cmFQPr+IGTynNhYQtu
wJrzcKn8dial9xxNdBvcajfwU382wAvIo48NCsaUNYlqLyV7ve5ZZzliJqfEBG+4
QzX3C1p94PTTeoz9IPilscLLtDHO1Mt6WPMupPp3F0JOyPZ5UVRNedDviNiPWszz
vBDwfJXYAhHRy717jCRcYZFY4Ji0F9xc1/26s6qEpfL0kZZNbZsoAHTC8YocynH1
71hWC8ji8fB+9pX3E/bHUHW/aFed1UnNcFXTNnU8HGaXAU8YUCkdvl5ieF3nKzZT
UNSRBQbf6fsQg1VPa/ZvX46irwshxBTTRyvIEO8ZuTu5ud6+9U+N5TlKFs7PGgo1
40jtTPsHNuJuAS+YNPC0nBf/RzZmuLlUg7F6HRgHcvYhtUp0LMGOCu2QKmnwCJBp
YG8hSrpPGJ9CAnqhMHPazGyxhT45lPRhSSWjgCCLcUsYgmq+Rw/yfGELOCVdCszR
+nb0bKBaZb6mbdzKiyt5076sFMAblBlku6ObEtd4UViKRh2zpHx4IKKbThC/fX0n
7/bN1krTP8+6o3jujIrFJA34xVK88p4yqoDBIMJ3cr6Rk7q90lR8Z49cvYO+YmZV
MP5QuLXf12aJa6o3qB2I8Jzkwo3ftKHMHZ22Yq0PjJRobjwD53pNieQwshOn/7XB
zI1kSMprXnW/t9sVRpZHMFZbN42jPwD9ilEPXmirKv+B6bvArqJaA16BLmO0ZuM4
ypkP/B+A1ZOacrDQmVyti4wsYEWKF5YQ/g8leLOcgxoS4dqw5VMUxVg1ZxY1asty
6wVeYP8yh8M2w2uGVJc3ip8NTH+yATw3r0IjAgsuMusiwXReOrEBIXF9I0OIucki
I66sjxz6f+PXDzJ7LoxajbDvBuyggL6JnJNyOy5/v0tygsb7TafwiU4C+YThzYcF
sKNfLF4QRO7PDt7Uurxa5Wu/npX3j4UPMfw38o+D0LGTK6lxP49NsPK03iaLVEYD
SshrOmqr+hvEKWm0FavMVLfHEI/tsAFwAmlGr9g2qc4zSDe80oj+8fu2/vD9FAOc
2a4lErcBxpkaQwxztF+CINmDLvl6sHQ/OnzXx+ZCn8wMJs6BaMNw+jCDQL53ah29
bG2OkPyyrbjwZnEhFzQvee1L2NSia3qnKovMTkRY0yijbd4Q0h/71g2sCV+BvXk7
HWxVBEwwQGXigfYqn9DNIglaf3xfy2SVSEehrJiYtH+797+LFrIcJnquzfzFeAvs
TVZReCV4fhN+/8qm7CbGNuqonUyFpuBSzw8fmg0oUEnXgJye/X+QLncsspxU6pik
fz3FwgvHjoIXHD2WU/7X+1D0VDhTaLKfJfGSzJXHYnUu1ZYRDK8q2ZP80v+5XRYY
upxQwhYIWgJiAoKL13aVPVgYnUSPWMhAcRFdSwcMyf+j7DA3iahd2ZvMYKNtelx0
KW8Q48Q0o2/dwJLxQDyj66AgEyt1LEZi7lXPKyagdo6HdYaMmBCz7uZCb+xKEkU8
PQndjU1vB1mkPpdatXXmam8V/n4h1nxWbcdWNKdO4+j6tgXkyEUKodWjlmK+EyfR
BJ0ikSJ5Ia4VHqMiOgEiDQygU6ONZhCKeDr8JdwtJGLV3tX2Vg6m+NecNs8goEsF
FovaCO6N/+1BSkf+UELRSOAL//rK4iwF0uBKHRfVf1v/NVAk6DLvkSPZViYpE/QZ
y6eVLB+d+Xzu3IV1Q58lZ5M3WcHd0xNGaojGA+yiX6Qb/J9fJvT46WjdVcfSW/YK
hXyaQ/X/cQZujniAF7tMhwLWnoi7LBe6k3ynJesw6tS03Vwoyho0evWH9XLdv+dD
yzalVdVcxAjxG4Ix8DuYFoWnawq38vWWlMy1k+IWfVmQnArwox2rNvhcO6Ts5TzB
UM2w5x4i6CFnMrD2RZYME96G8RPN1+eAF6JvE54zvy1BGlUpqXBgq4qpu6XO3U2w
5PBWW9ihFILLPjNEKeBBx9SK1j5q1DX9nhQabSMV/3IfojoYDs/fPEv0aSxuOtiJ
IW5W4rezYJfoQPaNcdcwaRCAi+KWs3Rqli5u9l9JKz41yELkBmCoBAoeYcULm4eo
1Zb9XpoPSUFCKmmgimGhHRtBUO0LyodovC/Wz6k/L7HjCVKk66gbwY3pLhVAyeGI
aorOLXbmgSnpnWbaWHkiHJgC9zE1H+8XY3if88zHi7oXd41CKFJPYxfoK1wpRz2+
A5qyJXJ9oZDYfVcUq3aAza/pL/Uy/QSiq6UsA/ETJfP6yJxvw1ZecplE/BDh0/aJ
qZkyEq/YkLEp4qohO5o4+W8Pr/bqvndcurVxbrM7HUp5Yh4z90PfiOd8rNqR82fx
pgyAKrvpdITs6ksiXSrGUAz0lESJ0SDpM9LIQJ/d4I51Bu28oGgGx7n/xx2JCsFU
TqtYpBDdMP+gP/orJtu3l83fMChHjalfoIOwXkWBO4TjJpOY0glbcAnfX1Ln+7g4
LyivY7cESTA2fBo2qL/IgcDG5lg7O+jmpiKDUv/CKgwEFTuJ+mp9ovTu9pT27iNn
dsyGLFNxCTgzDubHmdMrQNFBEiVwKqAehyNrFsUTfdGYHId86KEUTPIaqeYBYrwX
0am7+OE8Rvwc8uwS4W8+ToqZWvpGQiXttxKC73uaVgU8defDH2UUiJBsOf+fZ6i3
71H+oMUXy07v69Z66SssJiE8cCKiKiBZIJ2MVKLG1DvpHADdDC67FUsMH546XVhF
huenFgjaI04aCw8E4zWNxRi8Dc8yTA1aAZ5srw/+vu4GYlOlZFq/kYoCcCgC7VgA
GjcZdS3ooU7hjPiPeSWn4qc0iEkgytezlog1ia8PRRTYww6Z4YKCWzXG2RuiOSby
Mb7rcXUOHvDdEEjdI+m3wOeiwHS2f9NVul2grsaBBtLRa+DY5ExqBiaSxUEu+6DS
mJEE0M8JqkkX8d5YfII92TUIuwoH42EZzkURmerArSIhNVcEo5PbtckasEZvHRlB
h/u75p56OQr+JqbOGOa2kQ0tHA24BxENU1/tBquurTg4ubQfu1/N5+F1iNiIs5+1
pK5TQrdf0lxKjr9AKmuZAe9vhda3nxDxLhgwXUqM98vTtbbb1Dz5JP3GbYx5nXsZ
IZVSVv4H3f2vzKCFqv9oo+JMKaJl5LjPEwH2V9GsL59roRtIuxoAziadRKhZ9sR8
X8LjN5FnXsH+igx8FZq/3g5riyFvNJssTIVpBN5wRbnDZm5Sja7k92sMtG9IBpK7
9aKbJxFppdM4ckRnlsb2LOQ+1RdKjwh627hzMJZhX3FXC1DULJ7Vmlt9pBpkLQmU
joPffy0qnI7HZU7v/W1/OMCHx9FLwNmPk5nFG98vZOA8PoTroBVvXSG7dzVAvVSY
7pciPPFveUNPIaeqLo4Z6xF1A6e+Zcz0ViWIndIvDo1vicqgjPg0FmJuG+So6HcT
iYvkVoKjOKUOUf5yKA5HX0NFEhapFY53COwuNIrW+qTkcbVW7Aco3lsm1HdSk0ie
h9tpO1ZwovNNlgo76TG5ctqsfP8PhqwGDnIENCoxOUWV1DV2NG8M0jIBTH2nB4nL
tlXaZjErxjuI9Om78J/Ih59Gr6XwLnT72fKieVEkbdxKVTMlaIMcWDw7LD68yzIc
spB0+MiQ/wNoNDN39KqeVXEZt+eSCIi95KAlEZrqPQ1rX2uJlUm4iO6H8W+nr9py
rc6oMPHwwRsFDM+nHh5dcXygU65JSgUnYEh76jut6lhrqMm7AbkR43Q/+DWxmmj1
S7O3WGLY2JmhVW8tijFp1mjV+cOnQOxXgl5BrBEbWZGcsGKowe0YuOWXnHiHZR6e
agybtdPKrtPqH1yGrUG4glI1TXnQ3QQ/iSK9zK/g83w8GkKaClMWSfR+hkbOHuBL
wNY+bSvkjznV3bKo7+Pu2swQYaXMLD8bki5u3ADO1/v2AbG8HfS1K2uvBIBZGj6P
nnVdH4gS41hYoxvIfrI1gDeItbPOGX4YgBLVFydWjiCNA7gyYLAJ7d4lPdf9L1fc
HNBz0lOOm0cfcjJOJEyl9a+V+9mgjOrIF9XVrA2IBAu0vn2tGBYUkrnTYDULK4iF
czUEAg5YOk2Xx8/bpftIXy7RwmcuUjbpmvWWw29q1Cdibl7GCSSAPewU9se6xNJv
Zh9fp1W2IXNokq/40+gdHBFL88JtDzc5OwVtal3xG8emPTTAJQcx1vTe1+0hmP0+
/8uUO1iwyU4eUcNBXJ7DFOzOETdTL7zWyyMy3XQviOXPuqhriwGLoRAmtQfE0D2C
L4g17lvsmKDgi7+hx+IeXpXSPL/vhtMnXjnVP7PFkHYFx86YL5/C2mcgobj0Inuk
Djfv+EuHhCdt7n8+pmRaHC3+W+Rwrs41xLmhPcXgdAczrNp0kpjxv4lzaQgqm8/A
rk112vhajuQb73zyv0AEf7NbEqaJsCIGml8ng81SThnB1KEq5t7nuspip92uwHKf
AiA+rZFD2/undN+GRg6QG2sEqM3Ros8rETLPYTfeP+AtE5QyQVFDH680+bl7qku2
h0sraOOWDWlPY4eYzlmESaecKpr2XYidHyMNw/nI5Oi5JtFkgmSWaNV4KKFhdlbW
SeQ/e+MjUpJqqj7V5wo0R7N7p48wN/fpOUIXJWaDqYOeWFGNKC9gWbg51EfuyMZK
coByEnURGAOsBpD/pXEDL9fllL7+EonxGmDLdJq7igd6dI3+WFy3PpqokdnezYJo
WZm9oqEDFK5BnjLnYWkoTpGk0E7bMOUzGjMFu7SE1t/vJfHD32m/FOdpHzF/gQcO
BIfLAbLJXrqia+Uk9U7l88WIFkSx43IX3vlWOXXXLrV98Vtf4ajJJLSqcSr8qoGp
zSvliwA6ECVVJU9dlaDsUoIcUOlvnfXSnt/qnbx1ims51swkV5b2hfHcCWu3aOUG
IVFATtloUf7yvLNA16ko9yLzfi0lKJwtSrcxP0YFLNS7IyHurv0WUDbeyCIY/lVO
WG+F553SA+r7JU9fGLDqRiXzPnFyjWXO93V91J5Dacdu5UjcMWI0pEfZlr3Ra7yL
EMz0+HKwIMF80Jd4kn15Mb3eVnpNNHAa0N+i5vbKriVXkF0nIKKL2J41JZEKJIa6
dtHMLwD1r1vFinyzaoU+cgUvPUAB+ZaFS/zVTQ284EpirracfnyY5GqFYHywShQw
XmK5/T6iC4atOWggMVIsLp1/7YJeQmDUwG2aGsKvycLsNmNacirBPLnYnoa8I/nT
h3N3vByqtXqHo6kEDoBrfG2wna0hD9GrYcnUvrHrK28UiszhB/eOejBTlmC1W0Dl
LwLJCYvMVN61lBfhUvC+eFE4CzKllEup0EXIAoQR3XjjCajUoL/OTR7cdGJzNQ7r
04eOIqVoDEZYSz/8Aljv6Yh02EMFeriJSl/OgruXNFiyK1JpF17z4tRpTV5WMajU
k5G7FadThAp6pPqOTMP1VBWVZnAXDB8OSFVeifwoO9gtsCpGU5w/reugs61M9NJy
ocKWiDyFEUhptDHWqVBUY4mdXWoHJUxXb9+U2tNtk+f8y1y4rUFxUwzkZL7TcWT9
S1L+wyT1r+az16unFbx9oFUMQwvO+bQ7UuGNZaUPHKi4kWsop7qJ5lmYJGdSJSG7
8FXAAxHH0FKgIjJHv7Ivdet3pBYhm8EpNmFkb6z9RdcPAIEK0aTA87X8cVwkuAMS
BZ4FwTN0lgo76vlczGNDZ0DQnpNM2TI5s2woogyC8tsXVi99S//R8soYMHhl8x4k
BOYt2Yrs8SUHf+NqIqQGWiGdZwjfh5A4EUDQ3zhfOzqNduJ/Kjyxj8wUTNy4Edjt
mfsBMJURSaPR7Kw+d9uv1cRydj9BrKHe32FaiCA0/MJNeHWjjQiK1VCXqWTf5h6U
tqrsq0Apog6zU32IzqYw65sjtvBreZ2enDQmuSG09PLJIErar2/JMC/K2H6kB//G
3+bhiD5Qv90o+TwjSH6pz9wgCHYdpmpmWp6LYJFCqa//JDDoBDvFJ2XJRj5gntjm
FKGIoNULDy07PlUZ8hieZcBXps+NkEdNJvGgG+lkE9G4ld6UYrl65Dl1eBYTKPRu
FN00DvhTG7NzfseBnUYdiHGIQHPhhMh89l61v9YMb/s9S9dFT/oBrrJDWOSYlkTT
dKZ8SR9/HzwPZpUOYzXGsLIeS7jWXRMY41+5YJg3DJRJW2lXRfcT1tfQHAj07pvq
9wA/+K0OinESEJdsRnWd/XdgHW0pXXgVE0hwPYuWMZ57lBuWUJcb0Weop2EjRVGU
PVdnS3ceUY5Ls18gu5NxtzeFiQ11zj86Gcz/TGnXbRo/tw/dCsiMLoMwjveASC1S
7sFp8vkp559Q66mIPjeR8fKjdpaBkW+9y56lLBJUgp/D4d5vGvWjdQK/wCTVAxum
PQCESb8iryxN+gLwDNjGv0EE4NyBF1TGqq2g5xjRZqBT8/9UilyBmL4mPgQTUpww
0ezqgKrG3sylPi1oHaEa+zRpcefzrcW2scIsFaxStIW1MVNurzvBa7aEgQ+etIvh
0ldtkzyFiaz79+ZLbMcAFecajOmVuGj+CCn1kZAUdJX8fV4Gs3X9idVyFxNwp8V1
1D8sVkCgtXfdWz7d/JCVi5f7rcjCQufCZB0u6wYJLqRR/9aYW1pwQbqcfVUjXyJl
dINXRXA0KHn8/yrymewHdw669LOgFtUY1K0wOHY5r90DAVJBT8Q32Bf0DaMjGVwF
oAW/+RO4w444p3D8xQPjgLvlWS3jy2lRxgvnhXonWhUUjLSZNMrQSjt1Wwytmiqe
pb+DddEA+qQr4zDY1We0o5A2l//VqwW3+A3aNts35CtMrE461unfhazhETwyEy15
0GBL2mlFWWCV7vWk67T7EWgvYO+HbT+WfX+erLPp+KMXx66Dib0l+geKMhUt6Lwd
Pory9d1IdynTqY7WAb1q+pX3VJKDdtXZQZRGym2wSQKzalpH219fq62JGEGEkfJX
Y28hj/2U2cv7imgjn8tliC+ZdAIrHNPRf4swiOx8Ny10jhLdjFRFQ4+y0kJm0oP1
kMnMtMNgCJS7LSOnAjA4U3nsbUrGUD0fV6ZxuyurbZOS0JKpv7qCMV54PHrnaXZu
qfyAXph0cYUSwYQ1M5QcRIr7s8ENEJSsOaNxDPyAtmamVzIv0M9tEbSPG3jjVPx2
S4ns8GO0WWJZYAF7vaX6Sp2qXslE7MnbBbdeSKuJzDL3I1I171tuvXpMPcNltc+f
ITJszOjvE3DsQXB3f4sbFcNQKuK3RuDreINEPqnJ3N44LitjyR1CXltTR8g9n/dN
9ffouanFQWyr6+JrKDxSUo7x9gW4K94hRkioiRCSfb8It7UL2Jeo5UFqki3oELMT
2bl+DUaSdTr8NFHuMiwRi9vFDJ9/IoDTJUxP7BGqybkPUQxHDXljzmLVg0UgdGon
MKlBmJ8ocdB8PKmCqsm2Sml9UsIfFfq/dqyt4Gu/vtV2sgVL1utTjoC12nJ9F2xQ
zo+HkiYZMwhDPbZI3nqlYHXHxYLLJhDFTFDdALYHmI9TasLIXia8fJ7VNhGmwDtn
uJWjcs9DCiF1nZx7aQKS7Jp8aGrMPFCJR8EZrfjE3cSqMam9O04iczkHCD/5+wsb
bX6ZKbBUXISLt4UGnoisSJyLIhSIuZZBxyBrMR5H0QQHFCJf8CMYVS1qz6jRP/Jp
9MamTq+oqjvTPX7m4fcOZC8pla95XBxtDlLui2p08aWv7djZ8cAGQtSDN1TRixvO
24RW5cus5zHnLdMHa1T1jdkz7aSwleCACoayH1gUjsPZSQFiSYirROb08zDmKyNe
KqWKsX+NzgUrxl977BilJzbh9Qv28POcfwGx4rNgV4DvUpFUEESFlielSktz9v2j
1yHbJS3SrpVgXi4fKg61lHyb3bPWAgJbaPHabjAe7z6cfGKWJjAG7oNSzkuBkONg
qLzZONANikXOpuAojRbYVMNLmwAFTzchn/HI9pe7McsRNWfG75mg3CwzSMClsnwC
PZid+P/nJl+oNLfTzkn4WZ/HpPKB84w1DU49rYd7jORzXarLOJAFvp+lJgVvGTQa
w0OlNu66vQDivH2TZe6fR60OrPl6b3GYZJfX44kbzv9YFzDp3Nk/rHLlfWxTDXkP
O+XrJQYtBrPhR6pCPCsG5hFpu7OqUCZDgzqRe3sG4yk73NHCCEFHfpEZmrAOooVQ
1jhZ5z+6F779nkU7D4TteluKtBmtg5m5JQkZAWAzQ+0mETmQF1lXM+ncf5Oj5zIF
xTtwWMo0tXfYZo8Cbx1MZzItMx64gNHJ1n13XYT2we1EO8w8HDf7lHMlqFwiW619
dSDUdkS6C+MTdcW3VX8q4DIQFb+kqWRtNxLCouEKVcPrFdGnmnGSEhWL19+j0iVP
0YA5sOdsD7Maf/TJvzwZAr5UgSomZ+7v5+Azo4I6w7/Myb7fM8XKBvvS4aguJ4vO
wd9WtWQ+ADY11IihpPMCF3TMSE5qTK9X2i3P/1CE8Q7Q3iS556PqOr+q6jjKjIHE
1/fjne/ocWXonglhoXepT63NTg1AwwTOEQ+jk9C4+mi7fFSIncrjj+OsXIQrJut1
ZXxKI8pk+kUYLmsokkurej88l8vLIYXJkYHpNhIWQvzrMsOaatyqbVzqCKumjFpR
G41wRaWsoNQhip4WX0iAXNG4uYVXstVmyVRqjlfIynGWBknG5ag8MjLcTHZhdhpc
G3x9Kc75Ap3oAWcgwYqEF71ZHJkrMynswaGvvAwt4zGRHF8ixwmijm4LFnBUMIUs
z13zmk3kJvFqzijumS6HokEhe9x+NDL2GHQYXEJ3/ueEGk6hIWjO/RCfRuMcjn0k
d/Aj9DY6xJsNj2TcDZYvpD40e41FPWgv7sDqzPsUI6zKSkibEheTOnixCg2c+gh7
RxxFIIvJH4f7stz+sWTPkMIRwZ2/4Y/T1kVI9qQjcn1SOBTuEb3eI1YnSuQqJrvZ
9hM+wGUOyJLOzHFq1r3mLx+2XbW2UJlrLDKxz0zmej2/gYO/Jqmsq6sgUNL/FtWu
oELdCg/GfyDVtEL5pv6lYi2ZZ34YOdVAaQpMn/5qT8iTug6tquBspuvHZEbd/dVl
cX1V+7Tqqgw869nNYlCALULZwdSC4VyBvsGRVmn9kMuvhaFA5gEy0kuBlZ9a3JRe
euY8/x26kLo6mX5H7dC+gjAKLr6OAF3R0hJoTzxVFRfPBbKrphMX+ZVw1+IrQQV9
A36e8bp0lMwrfetKZifYehMi3d4HbQ1c1TDsjttwYPnIDSd23KCyTJYVnA/4axfg
7tJM590Qx8AmyDhv3OwGd1aBQw4zBKHAllF32N01MoVAx6gdiB3Vs8SJSog7hJy7
/keR3tTnQyjz6rY91gnRolOsruSs5ojqOiMdZIYg1CSx8goq2l5bs075PaSG0Y1x
lO0rJ3hAeMOWEwNI7Ohri9PylphJv2BBBrcmo5nWxN0w9Qg6aal33NNOv8rBlEN2
92vfclyEDzVfz/nGmOBeClmyIL435j471+8dbWHHKQvxGrbeAUvM0TgR8TfGWfJY
xABHf5SdEovmSoc9GeVDXKmI1IdYdGIg4p+RO4BS/wcn6dyZRW4SV11PfLg/iTIz
jy+vjpR+59S1LLWjsc+8MocrHb1NJHpqlEO7/etvVgHNdgV6MNNNaKmtOIjOfEdC
I1yTKgv4fseiCM/WlMAx+GBeLacaRY9llg1F1jTFzi+wjZF+OxArPunwkDWpfeuh
CEML+y8QTVnwNxqsZkNipTdnrnFEtQcFWRcQrnfACOFlgXNrIl8dpONnEJVG/msL
7R+4nTO/WiahqeYp3WuJErsr7kQZAv578E6oE75bsp4LfgEqgTJVxyNt5awwTvN/
WTQYmJYAM48u8aQ1iz0dWS/Dw2DAZk/V8JauWqCXTlaz3/ImKavIBPug9jOEUrt6
8MQqTwmtb/Ix78GfNGNXYh7rPolnRgGSDBirV9mz5h1Sy/EO2zdUwNvod2HmWi9k
Q+eH3O/c9wZ8SPphgokPttRXWTr0NYUWv1uQ2dfKkIvS3hIRfV9ZgjqxXDio/I3h
vp6zA+ZnuNS0iyou4yCnJE8PGmjES81O0jNAs4bsYPZvSPMNoGUrdGXCtXWWlgqu
ot18mCM9Rn9Kuw1LBjnNvGuNjV4krMfaRcyJSC5Rvc1UcadREy8hqMP9IpKRKKfz
DOjpnx/qiHghsbQlnCK5pj0qKwn4YTMI4mTukJqq8n3tu4Dp6PWAtqzN2NewX362
QlmE3nE6F3JsiLAB60dnO254WP0WzvX7LqDgt2AI/ofuZ5Wic8GXJjJg7Hgekd2h
WsH2T3hXwfo0cBTtUrrifxh7Y5ZY2Dn7vh6ZNdR9LZ8QQjwqhOVH/3qp+gjBFtyE
SNItvKRkPiWKI0HOaZHtFi019EbWsdKZpVZy582ArLErLkREa7uLf1KiwR7Hx3ja
YmpdgrXThLqWCEqhU6rWdXYsvQt+9mt4FzwSu1/oDGSy6XOBdDDgQ+k/mljkRgT+
g7Ooj8kWhbTWk4Ql/yFAYO8XM01YDsVWIi8fhjHuX+9CMAQqIlXTqcZHtiaZFxS8
4/gKTFvcnC1/Vi1/Sr6PKDQmKXRKqvsXRRWT0nRVX6f6GtBq0ui+O73q5T6ph4/v
kHwFRbH+E50BNt2nyRyrqFrn7s1qw1kDwO4eorO6/2i8GWU+lZLYhkrlLi/FXZgh
C+9p0w6nXVY+jdsgfNRTE4j3LPr6DgZi9hDkk1ue2r8kFsaG7FMuIBcWISvlVIG4
ypMzT/apmp8nREY5ghLZ7CTqdsY5kZk4yU0xYjW6XNBfbQ/aJaRCy2wSAkHGKlbs
H69p2Y/vswN5+3RpV8sKmW2VoohpL7CttvfG/CIuxlkQnoTCIqSZPgOh0bVzuMx/
h+YnOgjrRCvqgAi6EWRIc8AoVRDlWo6vhAwFVndhkolCpt75OMI8FcZO8Bl8wHt5
zrOpGw3dakm6LBOUwRUq5c2YND2MjINxqa1ykBxYfVFtAD3/UexjXT/M2VLdhs9f
ldz6OQL+0NLZIaZBrX1SzNxDJDFKT21kdm10cm1Eb/2GLMzXtFAImyYarEHsqBfT
Bh0gkneE3C2E6ZtplHy/FXBezf/EjqFlR04X4OH1ID2j2NjLOOzz3IY6qNGAJq7r
1BpNMEAF0mPdLefvSQzJtmXorzdp4wvOYRv+wjcHNtzyK09xsirLAX5DWHgkKe0d
qEAr+NA8wUBCN00xL0povaH8MnNEAg8AS8PSeAyHFm8H756qDyXojycRNiPuiWtL
V5Gelt8mlHApR1oTK/OU6or+nCUQCosVtiYdylz1DsMw45z+G6aWe1HOaI78zjP2
+B/PC4IdNb/gKHhfYWWBmgZMlMt0ez9e+eDTZKvOpQmU3L2nP8wBNpLFZRENBNdw
KNDsTgxwVgfb4IgsWD1rCtGPHl/lqGJ7La1zzetwF7NSX2Y0gUXJz51eYYbrAdlt
uT+LWrKxQP1mDjvUWEoLUySfpNBUHhR+hMvWzY3qZ7bZk2nIagXE4YXvUdBaAoIY
LYmNQwbxfWWac4nw18KAPyg2miKWs6rgzAw56BkZXxGMvRetrmHKkShGv+VdtzMV
fU+PtaPBVdXZYKxK01C5q/+t7W+WXkpqIXSWnK6PpODHlzZ9uBhHCfY2W6ObZ5ML
6jpedVj+js41cvEwdp6h4j+CehY8vxV45nccAoFryJzJSnQKXxOHIHla1plbbZ6p
dqfAalKTsZ0/5/pwtd/OWLzYEomzaEMexq5rZh/+otWr8jM1gwNQRBHLSFCswkJw
gr4Iy7qZr8oRbuhlYddcHuM577pTb77tLhzU4LE0snWwduwIGhxy+DjLVcy9qq+F
38k3TyLbohkPuwUbt8hO/Pq7GRTPLu+XX/TGK3CtDQ1rt1o5n1MiO0JGvgBpNc1K
joKcGv33iULj00UCKpPX3UYqE0R0Nd01FcA4EKVaCmJTC0rL8vvqyVY/syYqOsCO
i9AgukykDNe6Co50H1foVjWO+KlKKtKp/GuJqLFES6HbCzJ2NDOEmJQs1qtmkItD
Y59pQYtUYWSryjzDQrueBB9u1aZnKrp7o97dX+ZtlGTy8AKcZAbSJsjNvbYKFGez
Mqke5zu8FDtHTjikkD7iCiggvqjc8itqcyfhWUSht+9yU/u8+44uo2DN8NBoCtqp
9cTSid/hqmsChHeA4BnHFGrdVYfmGRNOhuMAOSGslrgdTPXq0+sAuPLY5jMS8B+s
uyaPi/4Fbz4uniZpvp5OFzHoqTMHCWLpBvbouJQ+4tKUa+UzeUApvsfraqdPx6ec
ORABd7lhVpCOege2mYb77ZRbCpPrPq0DoKfrEEyDSm0k26i/z+qK93yPC3fyUrYB
PcG37ZkRwcHzq2MkJaNQfp4eQ1HMi5ejxDgWI1z/Ox+Ccqhbe+mQGWTYAu1Cjzz2
OgCn6EthUVDQWpHNZ4lSoCIpEa7GHBp11D1QZdcOhH0+lcNUVN/F6gDfUdYscZok
bPRA7Qr+6hlaEEOj83uqiJUm1iXhWUIlOEmHTA1w3mQ1rU3GCmRPAXYPybRxeISA
1Kf/zE8NjiH0RuVoXvE+X6g9ZZdhfNQLGEKAPMw8rim0GNoziek051Xrn3eJn7rD
m6igqIfVGBa4weFXFuwwbXYW3x4DU9ufnvasG5ZtPpRA5tDYQMh9xDA43JXiQ+W+
KDQNAzAxNp07S7w+X0sGWNa4dGMAcmOK6mdFBjEYh9QogKAnrTh1HysImwbc/pc6
9GE7MsXezzaoByCes2NgmLyHHTC8Zx8AJV/y0GJOeWgupVwWIYBcBy1ygdv/VFRy
q92ZO3AtozTTdeEUDzUhLhsFftwdnJK8q0vqUMbgH68GPw5DMmtn5m6tARVdNMQE
cxKWr2YkDSNa5Q6MrVZMrnPdfd5U6UxXWCd6rtIuvuLhaW7FdUfcEMCmSxHlLnuh
bZ8plkJfIeRFkuIhYWvpcFNBnu/R/WVEysAokOJvuV9z60yLp/bAngd3ON1fp/BX
l5GvFYP56IJ2utgpSHX1XW9nGMPixMq85mTTKd5aKdZ2SoMV00shpY6cSLdTmuu8
llW/vpRtquOMJD8XeZF/r0xjEmFnF7W55effBUpzhTJ9Hzh8dgaRYPfirQWM5bj8
dkSNJ1qDsG5+Y73JAGi26Iri6f85+40QqMcflCOF2DfFkKoe8QpiLCQyptbcCRjb
cm6lpRKM6ZeK+BBdxm/9opEZxZ6i/8TQNpnr+2gC3z/W2sTmQ7G9te1I0KL9YIzV
q4K13WZ29UGZ0C1sX40nj3mYTMt58xHLqnv/6Ok4Yx2orPhKGNgZbMMw6vP+N2j9
g5aBfsLb82JSZ9ehwzR6t9LdqgmrJr1HoHxLkoHdIHNs2f1ym8XtbJIvf7lDR76E
kIqvSeJemliZ8pGBF99d8wQ0RUQ0Vw8Wn11rycG11oEXcJzLcI7IDqin9PHszDre
Rf3hjgfwipvYi/VyOqCnohftfzDDaRdvwp4C+bcAGnifW4Iw7burXWne37FmQREI
q82ybp8oDIcjGMQ4WE1tH3SYrMAYK50ItrXoXRamGwhYF75XBStlgEW0sXCmklBz
m1xM/w5v35Xsolu6m0C3bsPUA+4kMjz6eEcsXpT5wc8aPGPlkaoarJhugvsBqQEQ
y+CZWb4JzrTFQ9LFnAH/xAXr6Ha/QsbrtSYi4q9huK+tczikiQ3Nvagf2w9HIA6k
9MuQ9vJWQucbg0QpgiBBPW5YCDiD9mj9E90AhgIQqKfvkPJL2iUBKZheAktSm0xQ
dikKZrFJdtQpCVZtHuHGHe9+BDW6zFJPs61c2PMn+4K08rbFIWTe5H/Lu1igA5Vn
JByqI/hvtFgsvHK5Dhpbx73HygwhU/dFgdD4VJxM0guddk9SrC7zhrQSOLp5MBxo
0MLhlmvpg/cJooNe5qpgNP6RrojihJ+ECi9LgONR9k3mde9RssCVueIsoZE+T8Lr
TXL0k2thby2N1C37JrBJRVA9YEroPZVuOQqdRSN4/0x8iLrpPJpI95R1b9XM2K/0
sXAkts3udvHxVYzmKi7PkoC2+1tUoj0IRJ5KZt0YfBQS/1oJVZIlr7ovql2+ZqZ9
3yJwwOPA6je5MxNcd8wHYQg/BsjtHJ9x8pHRyBNfulHF/rUI89Pm+ZZ30Avh9M2j
a3+ZQenx3us7FH8BYrZE2DpXwhIbLWJilNTLUykcfFjhkuAFGziW5b30n8qq84g7
WdNAUazW90Ut9rawu2rdob9aA/+lPUUaQkYgYlxVS7ZYJFVHg6s5E5TnahHV1SlC
DOpl8E1lOyYiZu5kyikTNXB6X6Js3/CaHtFWRLhDo58U2pUz7TZMgNs8Ggl9o3ts
zj7I4pOVB4+8qO6RcYt/h2LxKTAePc0Io7itPpS4fNPtt43mvexN78g2JGmVztQF
fR6a0HEgBp7hk4NYcnZIVqzLSF4pCusQwpKDkfGrfzg4+KsoQOX/z0fRTkhl1RGu
C+9IcRgVgny1TntIlQcs1lt3o+G/nIfjVlQEV1jOnFqrYvwvkpVoWsensMAkCkjT
GI+6p+uW83lMwkakoOPtc4kQlTumoNJQlMW6VMYJQ78jptTmBTLthgVxqhuX8/FT
NIdfKfA1vrqRQS+0k/hWsmUy0ifQPAgG+IRp2nhvlNR4LdDyyy1A9FCJl5gAdjoE
H5ifJ9AQa5kIoxynbgRZIMfHjWgYrPKST+pQD+dBo6YXXZKtdSitx89vSqz1VvXX
grpbjA7tqVCOR1HeKNmJnBYhZy9/kfiE3lwq8hJ065ZytegxWibLW2hvUM74A+Zo
jI515AqugIBU/cRdTtpzqiuqsOC21oGWpzh3dXDsmAib9P5/NOf84Ynonp0B+WIp
97T06aF8OJXId+u9rWHUz+Ye86+nyCp4fcBqPUu8yz9JLYJMZFXf1T2Kt54YeGGi
T6ewKKGWuOORG5q9YS3NbHXoOoWqlQ3IsYRT8q9T7NG0fdyfADhV3uZ8hHdrtltQ
GCDgqqIWA8WAztxv33CSmroIIy9tL3BJJQxYw4TxRlXkyu2/D2Eez7Qvt1o3wa/4
oe4s6rkQyuq3s+3WMW1gdT+sazF1ZAPgpsIEL6zpR2B4W+PvYLGGPrWNJNCwAl5g
W3u49rk42mBVpGgtD3J3BE4mKTGrU6nmekbP9wcaHX3x1d3uyxuP6yoJfMYcTIXb
02WwveaHQQUFmUYjpGlQN8qejIVqtn1CkxF5MEPPSSYpjyi8cRJEUv8WoWw450j5
eBC/kET5CJqPm+kyK3xAmzOY471Z0jOGMySTzQxd/p7DYYgqIQWOUKFIY8wwMcvA
Gek8TCyGlL/qV2BOWRLijg1NiYzlsQ40aSwkWOUWfJ1aPw+1LzESpCOboQtXKpto
fqcRj4OtYtfjn7F9jxGq+hGRHf/rcJ+Onqa9AL2jXoAoqVZToFkV0Jn6E85OQmW3
5dzxeHBP7MeqoBX2Z9YrmA5Zrz6cjuVA5LKv/rGMINsK7YQjhZUGffy4+6CSi+ON
od7aQPJIOOexFdx6b330QyAKVZcxD5V0r2SNdx2mTUg0E/XKZxLZK0eXNpSn8IaH
2+55M0wWhXbR4OkAWtrWtVle/KoIn6vyQuaO2Wwzj1lbE6c+R8ocBEL3tXdhkCn4
Yp7vcE2gEz8J2rNQSGiV1/dbU/ebjDzwLjENSqqoEqqYZzJe9Bh5V951XUlUO2zV
qyHPlYj5zaq5hxXz8waKd7UXC/f9q8Sr5E0KFD6DoqTwBYukMXLXMLp9Zn+NrCUG
xJlUqst3X8G8Xt0N3etW5tNIYFi5b/HF2UQmeQZCqmiMHNGkhOcxTby++wIjpL9X
fxRa31DegINB8hNxlqKXRgNT2gJqTBvULOos9QFk99Atq/bb3jnhGLpsvuKaCbDG
Dq6Z34nlLE4B8DiKb3tG1NOGSRx0PhAqg8rI3hkQMzWMptbHP/6a8PMlhFNAve2f
yP88Wz56UQKiO2Vpv6oJmbs29gjhffG3AYa173I3O+xmFlaPgpbo3Y5R8uNj2wMF
kt7NiOlw1IAgR7ZOjtDkzXW9V4jfFYhoFh7CY2pe5XFhie5zgoBH6SGDPwsyWRzo
vI1UjiJHZ8+DkvmH5yahkj4W8WUzdvXyVupvk0nQNXZYaSjrAimH+C2nfHxgtV4R
IxPmThxVcA0T3yjx4lWXt5+bl/9KeysksnY6eOICVJGXOix/adMlg+O3IBJNpqxu
4GJy7ndAjBSd1qiCG/w82vDDkvoR8OejczZSWv5hrmB289FKvdJ0vjMTZ5ELLV6M
VSjA82tFQ5EziwAqKIBA48S5zLtxkZra1lBm/0UgmNMFTrkYTg6OP/ooFYSNC8iI
HbvRT2moPfybiNMmVRCNLNZPZEUiE2MT0IS+OWvNHxtFladwoynL8wYDvv+SQ91b
K2HcF6LXixzgLVjzqh/Al4dXs534shulVi7y2I57H/8dD0HNzfSZPUYzgwzrglFF
NRiIn7c1gqjzBbbbj1/ef0GFykv43kQfiyYeNOTzb2hwHsjqdTkoGiTPZ6Al0ken
NwoiF4ufSRgZzqIpuhE1b52l4WBT4ynAYo3LxGDY3F4+ncpmMJSIsCkcrRobPAMb
LWTF0kQEPziuF88JjaJECJzxE+V2JWVeIkkr1risnntPq4QALtZjstVhW1AvOm49
zN5T9sf+hQBe3jt9xnzgRY9dipK4AmWGSdpIcmC2qGx2LldwkkzMQB4QFzeEUn2w
ySKk9BFLvVYLqeuz/y9tJvPFefVPMkggQcQVwclgGDGX+W3ujh6XdjMkD7l3zBdX
AXW52HYUIGPFJ9+upNMan7P+1+DK+AVJQOTH488LBXEWddZuEU+YTNr1wZUXQi2y
cCJulgaVRxDxKAgH91gKOt5Ef7X/NmikdMezizWInLMU0B17cxbxB6VRcsDYBQLn
Hxg3vzYZq9rxgUJNRRRhdgX1IxR8K130R/ydljLJx3/s1ET0I29wO56Cwdzjosff
dLo4pCxAxhgX/Ro1af6mCF/RB68G9+ku7R9x8w1/szCMrsvASX+TilmnatRHS0uQ
RptLCA/HWjLokHwmlp46EHpF+T0Dz4dEzoGr2aGt9IlYnxBojwI3Btj/QH68zlzy
JblBU/b0eKaaBm0xHv4ndqyDn6+tK55Gsp3jHWm8Uu9VloP/sq3J1sAWEFCzEZhC
FPG7UWsEgk81iQq6zM571tcBq8Euib5UGCBR6f11wvf9usnUhy3xXzbS+drJMDjs
Cjri2+t2OOR23U8AYFn5HPUGXoMpH5v3kqVGUJsTIdVH1OfmSrwNR5HNc0fQ9XfW
oJ7yhvtJXeZPz1x6Iul15Wn+a1s1JrtkmbFCQbIutVdHt7TyK5OnoZ7OVIgsswXz
vZvvU8gmCdhDwOqFWZ1+yCs1CgxHtH2GkQJH5MZzmYLkGEEA38HGG4nFvD4dTKKK
gNoM6VmWpwca3z1VHtXOTFSEuAm+krV1a4/lia/aWueOvqZUn5cJEHEGBDnT+CeZ
AhfJVSi5zqSGWmqkQv5calWFryg4rPtb9nGOO7Abs+fLh0WzvpdFbiWx34mdtghF
EDwOGFJbPLlvFfoa6+qhKtsIJhC0VArPCIenr2mkyhzb9EV4/JzwYjrvYEpTplwu
wx2prElCaJs0udVO19DFZN4jCMpfIuJjMD4hrFoOx5bic13HJElYlwd6AF/P6Jht
DekcjGD5Ww6NOYCbd/hrqPjVU+Z6htonIIu9qddssh6ejdA0Pm0gVXISUdRumarT
GRJp6Ur3t1O3OlZnJx+JbWkyO2htYtoi8vFTRKPYxxEpB1s13+SPR9oRpCmTq7Bt
TkMpQjGZm+jLxhkVQ+Rpp8ZcN8mnG2mKA4ELsWftlcZnmwT0xYYi/ecS/hH208eO
0kLOXyKLFJbXn8Pg/lLe1q2d72iKajDXt/Av6pAcgm5iv5BI2sVEDUiJQHC6xqgW
/QgbWNxAEPOAzfTazlHb4+pJxBSzVLAplF9HcG2u6XVEjuyeBoFdJjjPk2gplBwP
zRR8aNY50ehkfJsWZTjcrfYTM3xh8n2jCTYxCX5yQ5cgsumQ+Ir9Wfhd+BBeXGo0
AbVfaVMc6qvpVr574jAXXR6Zn6Phs9xo/mOzP4dGnjnBrWGe8GbALhaJlI+pLmo2
zKLaA1DkkcPuQ3TsLqsecWBsLxqCXeVcD9XcxYW8z4ObpbbH1fUG3NKsCIGQ2h2H
wolsQ3Ipi0BQDNMtuH7MnBwGEnlKhQuMkS0xfGBxnRcBM2xcuOR852cSPBFr+lZc
j1JeuOjldOBSdaxZY5Zww4OCf973OQxm880OxR7Tt+FjO1kStfD6z4gAAkgegFDs
etgy6V1zJC9+sBAvMuBKJF9nC86ryQ+zc1KoyFzy9q/MUheg1HQkhRvLjNW2/Kyg
YUtwAmet/8Jrkl9D/2UfGiDhfu06M3xrlUaFyswNeLh2kn7jdgoBE76tr8rmNzxU
VUMUppKonLyj9Ytwa+/MMmCncTC/2+T9cRmQdzhLBjf4zYKGQf+PmnkGUm4LM5Ig
hekDig4npuZCRVsSO4WRUyXnV2GkGpoBm/ZAzYdD1wqEW0+NKkp3kvGoInhzWWbL
+B2oxHQ390GGl8VxwP8rHjpJ9kEWP2UJ3oyRI+lWRcppzZFjT3hT0QASEkbYN3Kq
VbrKo4CuNN99u0xvK9Kt7sPLggR5uc6CZCFxumZryLeydeO0wt89KSadncugXdyj
kRukvfojPFqM2Wa8VayyiSzsTEMTeIfjMjOVUykes+1220OW33TZ9c30rrtFXZqY
tzzZcdtwNZSofTxGxs1Ua4wNHpVLQZwFHIWkMvgkkMeJoFwDnJQwB67U8Wp4jlrN
fCQE3D9Y7BJ2/qw1uZiSAphS+P8BEpjKJ2pS+dUzzxK5F9JjMZbBbt9iuLn1mnxF
HU/sXPLBUI2SwAWshlUTt+6Xb6q2jXnBOhlnOU5ncrs38B7FZagNhMbhWWUDtwQm
gkWFvYf4PgGwTIfsEeSlZ6D/01oSpDlwJtizw690Yiz9t9wV6x36ujWfROdDDVKW
DTyObq524e1OnrVraSd5+0IY9y858sccZ0tNJRTa9fnae9Qwuey8XvDXZzmR6Y0l
EVdaVTy18MVqDHFJ8Jor7dDQdZSvVr8AsXPbbmwGkEjJ93lTzE+qieO2ruBNkDLR
uuk/IMh+s8JbsNNfyvC5TKsQPzyIL4abY/9wGCvDrtEWICI7Tw+Ctz40Wh5X/Gcz
eXCVuDLfJLCdTr2ib7FBogLiOmAO1NRinKaN20XEImtozX+RWsTPBiSwLb02OBKG
VGegq+bD/mOoIelH0nO0fguNszsXJw0IS9O6p1SNtBY6s7/ilHN0AFOdkULFjmkg
PQYUesyi4g6RGOJ+3FKBxA6RiXhbGa+gfWgNrsqQYyNL60nQwTgj5GEaJHbyOrLW
dfA1Ga9Cgdc1EXgUzyoIk59KD7/qcXPlfICHGU9gmpTiOfc/oYLZRDrfkbMuZMqq
Hs0t7vCK+K8oVB+fiBJJdIr90BmiWEABUDEPZD+Wky10EoFxqGUpZWG0MbyCtHpV
u+IfIFHd7lmwyd66veM/Jlz0+2OJeXqLgozCNnA0s/2TTSyjpGV9BAh9vwyPvU2H
qnymfTSMoM84lTnrVudMI1v/XRqfDfGEEmpkIinAD1Dlf7qOig0K06wxOIVTkOc+
MzxwklI/htWJN01zusyL0QTMX5C4Y5vqIAuJv4q4z1slhguuJ4/HYJ+/l1kfc4Uq
pPlOciLxN6CIl5uhUuJxS3FHbPukYEVwnFvV8rWgF99K+udwFeTdrwQ81lkbDMuS
OP8KrK0Fvnp9FmF1e0f42jxvvgiWFe6pjH3IKKQ87LyCVdON9ihkK934HArsPfsd
88YC1rT/t2O1kuOWFrFEdN2SJG17qDrBNXEWjaUb0It1SsjhW4JyWWIqH3yMUbI7
yfOSTrQAYwH4QO6ZOTEpjh2r5hY3DKPvPwvAV8zOVL2fi2KrK8VLy5oT4XMHQlLY
9JnvtDb0V5CWmo88PbdD1thNyRucm27m7khRNgE4yACCU7A/QhVxcCe+Xm8VVdGW
ipu036OESe+pvD9F9ctQhNliy9ENwYgNrld2d3aUswVlax09zIZJAFI035WU3Fcs
j5CEoftbg4m66kpJlp5mP6MRO/FcpVOEpLy2CTSZ8GIzfNfH6kbS98bZnVZyBq2V
8kgCK+MroWSSCx3CZNFrorWY3DVTk22EPTyMeWUm97wRBCH/qK/zYwWLk2BK86np
yLx/A3gob1jaoX4Ol+dutgTRWjfrMmcdre2nIqKpdFJSMfRXwXKs2U6AqOUawt3+
OwTPJRowiNo/pMddMRYjXPBCNnZdA081Mc8StnVP87Js+CJo4D5tRc4Tulm/6y0A
ra0J+qC5IudmtCzzqWe/tvvxwVPvcW9UEUC08UDbVdgCLHnm6F/7toK3X88OT3xh
DR3ZF6JlWV26bYm0JugMKvDx7CA5qo0H/bRcnlpmjDlDlM1SEbtJDot/FPKQlxcZ
xZm4fisGzzOsMR6eU93EQ30YghaJgkhyz669XG/wss3F7BQBCE/2DggKLZrK7CX/
7Supl5P/JpOicDQ+8KgeGnPuB7fj+OE6mnYNsEdwFF6wHNl+Y+Dz2dT0WexPIJTy
R02YgDKbbaI5mQD39cE9mSH00jt6pclbkZV3bvxMhsCVVE03MgUn/YghkBS1u3AU
WCE2ERbtW9FY1gI/I33xAc2UU7PscrwKXM89VWBY350uLsFFR5UYOE2TTZJMM5yS
6szpkS2ngqXskJNUqAN5v/5Vo3BZmcNJowmOoTY1+/ENKVkEhXasDcFlYWCwvH3L
KQLA44exgjmFBr3i4vYqaM8VVDjOwbxnKVkZVVVctmqpQ6qBpXuwbDy5Hw+WZfvx
pMO5ra06Cw7fHL+nAKqt7SAkpP4ABf7ciVufsmsIVeEBdggHhhNSpdQJ5OB9zun5
uMGV+0zliod/uelJYV/6tCjKz8QPQ631MR/ypwrtwENPKhX3w+7W31j47Kl8jQbL
Mme1TTqZjyQUCaK8udaHhfqysS2NReHR+k4S4XNAdftyTrOR0ZfZWnWPObklRhYr
Y2hQBmxtEwj3k1NpijK7HmnnQR8w2qb1+G4ZklnjjKtQbwCYiYxMFGLi70+w8a9n
RZ+6Cn3xX6UBCDqzMQ3bOqbDc/lteLi2mUVJCa2r9Hd2KNY8EGncQutyj8QqksWb
8gBwv+fHl5WrdD3AzJzNrZ01J4HZLyjHLRIMLr3nc8EYbM2IAuL0YXRLnsNmms0F
+Vei4Hsv15QAjzdcmtSNzgMYFtCejlU1QwlZFzfQJrEDSRhIF2LfwP14MUdnt+2r
I1Vz5/e8TbEHJ0ZAs5z0LEpD/3Oc37R3Gx/JdXepfI2iVmSrh8tnWYAXsOjebr0Z
kiChLcZQh5nRtmoYHf/lN3YTWd32cHvh3ddjQ5I0iZqb7mCKRv9Qj7D9I6Awg8+w
csN79xGCoWQ7KsNKS4Vl5OC2ZlRSLnMwsg98lQ+Zvh9TK+6eVxNE6BLV/uNYa7W1
vTaVIFuVf30crpmDvLjidQ2gZHt14Cry22HlGPiIqj9hQtMMUVxMBbuhqmHJO9NR
86FG55/VxdXClJf/vSVp4vnasKYd4t+HIkqmmvCFfrmIAxpWqXJP8LFl5mVbcpL/
58ZgEpXFb2bIimU4VDpcl85X08fhXDxEc1yhpJeJ+7nHkHfD6ccn+tAHazPNhKbg
FQLDXmMljlmRgnEq7rvyhkB2Viyiu/dQPQQWzw0ivuWaoe6A2n9Yofs+06iclHFp
bH162M3qFfX86uGtvS76aY9xQk649h3CnL2KD2wo7IULfvBAw2evr9vricCBhPt4
XvxrF4i/Tzjrg25ngAsXC74Q2mUC2NVYNKvwDCtgZIKUGDru1znckCG6VyF8JckD
ZVLsvv7DWsBcqr1FgaHjA9xN/6sQMCccRjsa/5RKsQg4nd8V5oE8NxRX5P/+PenL
O4QCXdTDuSG1tYp1ibVaTRNlkBk72hCHz1MhrdZw5JJTqZkFa3fcsgmDR9BHvcQK
DNVQomTaJwFGHh+GmK9D9iae06xCD8EU5WkM7QX4Km31E8l/InM3K+Q8DtuOU1L2
R85ig8Uw1axJZ1pk5koaPZUuArFmGr3hkt6As3/JIN7ha0yVHIDUBL3LYP/dB3WF
eEfx5ym7OAuYHs1ZygZpJDnCSlQdNBtI3cHvCgm/xJRIRjrhRhccgmAarSBTbtvf
35fonYjBcjyLxumGd4f8oOfbeyWMOzUwSiRdZSNz1eOyxkN4fW41DRJKx0xrAJG2
dnBNrYzM4hITik/C9g4fgNvAvYXAaeCnCJ57uFFG0fVg7EiTn4NOzjNT8MfUa/6f
5UjOU8B7GF/yP2U6mDQyR5ND/DzLZVy3iE9XbfMyhGUadTB2e5Z44PF/7XzGtQ7o
xmwxhgfzk6vSPw+8XwGUxf6b6d+gNXmHOtftZcXCIs0YXsw878gmzubNi2o7JGow
jbiNsXZk6+QFoCkPvoCsEhpkyg/UoVIfSjzmKPNcFZzxDvdROGOKa8qKXrVCT6qf
gKdZ9A+BltuipADIRwZJiezyjgSD4Ptrj58zFebMareiQZWWKMA+t3FkLjtWZAcv
1fN2wZk92AdD3HT+nckCDhZ0xGYkQWtAl/IPYJzVci9rJiTXENVn5OT+ihgL59ak
PD44HOYFWBAXfPr6GxdOW34PFrxy7Br1oFRY4YCC/HnubYdiRfWkF3omI9v+2ahx
OKEr1YL1bEhWw5kYni6QFJ/wPzj0VZgSpcCowuRVgqY+EuA3NkYbgLgmT6YuDF+U
PHAtEE5aZVqZuczqpnBPypYoVXnt8hmJRYXlNodqEKNSiCVuK0J+ZMdf00drrFij
zTUzrkY1zOYyxP/nzVhG1rQOS4/T1E7UA5y8eRxfM6iLTY2G7/nltD170LD/uRY/
1Sr1d6dNw9RO0XdFiN0W5JJK6C9FF31PxOXohMbCNVEzvynkUiK4MlfyjG3usW3c
vHFRbXZkyWU5mi/11dw8IjbL1YQmIYd+SN9ePe8hidWUpuHez9cnjvUjchxM1BJn
ZT1tmVH03pkSGVfXiEZZkig5Ywv/QkUXXRCkmvN+xTPS3NGdd0XGpPl0gkCCH5Z8
BrfW23s80MwC5xVFmxA9O67AG/BeTKtUvnKYrkRFUyviHXjwadHcGKk6Bww8idn0
pi1wvOE6EVZ+X66FuqidRYbEpf36FkcWM7z+cDOyi+WeqiLORLS++CU7LhEBuS9c
y5QnkFJDIn3rKnb3+KHnJXqFDJ50U1DHJfTMXoj3rVYQWxCM58dMN/TTtP205D5Y
YXBzQmov/HMIRlKDalzdANyV1Z5hnCtKxE7naE27CvleRoXnCDIILCSL507B4Xp9
jnxDrSHf+T+/YkfpSePY9mATRa9fPrmshkN/uVlA+MM5Elyvm3YzVrNhUUgcd7gk
PszzPAxhi0P6VQAih/Hie6rNBvWjr2pm90b0I66HKIjdSKFQ2X6cI+XDhQmj3MW0
S1t4NxZ3h/P4wUKAVdXaHfSRL9PaajEnGuJs1eu08DMFqIY53ScRfkqY2fbVL3HB
GP0Wv10m2hlAkThKX4lfmJv24byrzZb353kVrqPuL8xHLiBcRuG9db51AsEYwaqM
V2enz6yqHk4GLqhQLDSG1kYd0fxC0lQmOB59j5f4IK5tPkjIq5AKy7pUXiOu6hVd
1bCOZdA/OJGHxlhyg7fKzPZTxw+hx96Xvd+4TE77Lg2rKOk1NTYqnLPFCavkgRa2
VwcbdO7b7OqbnNV+/J2kVZB24+pH9Lf1687SlAQYnrqNbfNilFu5Cy1Vz8VNyQIh
CpQEjVlWsrK6ghrTP596ceui5glhLHx45JxfRfHKmm/0R8oXK9622CWOX3yhuFtZ
cZWxZ7vvPGmjdJ5WqMRsu8bh3KL7zCqHohgxYQvDdpzXebP2pNCKNqkYeaWzeI/+
T2dWdxTdcFAAQXaW0Pj7283hl4WhjhaQRTqL/ATbge9i7ZKYKr8LiLJDS9if1N96
gWSXWJm4yg+wfBsppYSAkPVt3vickENMHCE1iig/+64jmY8mnFLu7TzIg2nb3iLo
hmY8lRTt5n0KBSTd6ETJNzJp/b6E1f4Zv9OB1sIMWtw4chD01ww1u6Ulhgd1/ZXk
x7XozxhAparonPj/4xQmZmfY1uekPF+70coxmYgYNJqueQfikTPG6S8g70v9U9wD
rX82uOemkbf32/a/vrluaas3xR68wpJg/gVXl1GMmM8QT2wcbIBoYk0expOi8oCH
Bp1ZfiHZZTElp4bhL55QR1O6NdIr5ZlkSPkapYDmhMbVB21/jkcYUkwchY7GwIWs
WrgKsT+uBjYIPwb1pzn5pNMpIpNq3eGSe6z5Y9RFM5j9Jy0Pnhdv6D4dVKZh6mic
tSY15yDZAG/eh0Ky5UtwZ1LC1VnPu0eMZH9myR/5R+vjjSkH5sljknuTD2sbmy0a
jaYS+VK6zgNL2cuDSoKT77zU4dnLBM8q3W+jP3i7u/pDqCqwr2DYer6llroDlKpU
Mecjt8F5xKNXBqYXYGTNITZiZxkoxBQBcpEGFw9NzYsuCf2vJ0tqtWg2vsx7Uyuk
Ghz44y8t+r4TgROdRH62NE2JCfcZfXy5hOeTmzOlMH2yTz2xMBpqf63EkOHMH5i3
IT8waWlca1L0DUxko00ebhWOlOYhMF5diRw4SyLZuGF1LC5qJjHfYIgXjVYuFiXh
9Wfli5ktYaFkQY/k2CO5W5bUGtH5hBkhaV3TB15mNr9HDxZV+0P24WyvOgwzbjKs
bdR+dXdBe5QKh6zxtspN5e7HJ5zsMjVeRVQIR9b4Wkh4Bh8xHacKpwvzmqLmhkPm
K/GiDHGwjHZqmC8JLVmJX8/Cp47dL7gQQzRRg5obzTUMWhOJ7yHU0BSDqrpcRoW9
OQb7Fq16a0wqHJRKgXntpsBJgAZDdWEJZVrgd9y1dB001LeS4uYdLvimmx94d2xe
QprRcnih17pvWTQPvQ4LlTXF27ZBz8O/NP2rPJg2F+IAWo7YwiNox8R8C8PCT7On
qP7IlqX4T4GVsm12stBO/+MD39283RFhMsPiIgnw2wmFlGlKIl8NpmjbrbV/kBw7
LxKoH57bd1Yn7XCvWol4xS57nYKEs+VOF6UppBZtR0uZ4ZrXkjd68iKoie4enUk5
IEYADbFtsT3AakETnzETYSwQKj/jPSQCKpPV0d0MnLsTOJXfxUPCNgE1/7eSrE7I
Db4bDjm+GA1CLlj3U57EyPmgkap971qKMvhAmh8K40I0NOtLV6vB/H1tsvZjKhBs
XGJ8zelU6pBdm0Z+vc5FIndUS7MdjiAJYgUoyedosWrUV/zPmmbhIkbOnFtho5dZ
jcMICauNcNdIeAkl6ODwO9E621B6w4o7Wueb+Abgnrn4BdN6RCJKPTWn/gJWX9Cn
nn27cvmvk0FqOeHjVEUe3freCwflIxpN5jjXyzCtw+K9ZM/tptrBg/JqACN5y1o/
CaHdaqGj4fBhmesvnWvdJtgDGQe6vLOPwfSp/fseH2V5TMNbA7PFXLPXE2Ea6Gwz
CpwFrv77r3R2MZshLpz7DeAdlCnVzDrlq652ucAO2NdpCB9ll7cpZzY6tZ77kDDX
5bcBSaArRRd4XFQlHOGlr3Y8zQas7DMygIBSH3Ih1ciY4rjEZPFSLz3D3xID1pMJ
L934lK92eyH5YjN3vd6761hHucDlupxIRNCSLk7oKJUonxgFglyW+w6GuxsS4bJj
R/rVzK0TpK0sss6fQudiHHDPQiK074r+xVMOAZKi69A4HB4whJL5iq3ApdyEySRu
93CdwENf6vKIZBqkaxRDfzQbWBFSO8SZS2dNxFQL6DaPXAKl28iibrJxAUCMniQ9
hUM2JSVwsdQDoXoyR4Oa1oeodd9T3xteRWnVhzgU1T+0apfEWLAK0Lnr4VBoNL9L
f5Gb/DWQmECj3iUn5Etwzn4kCnOdfPcY7pZOj8aRNiS9DmNEO8Vtevn47stoaVR3
pNh268lhMzorZ9DPNA5PnHrKLlx9P4MoksAB4P38gPlHl9aOxeU7lWhKMHXVd1ww
y4gdPDPOSrrwy8WkBZD34KFVdHCO4jLxCSf/0AetECHvI5Anni1O2wJVWWYpoWT/
gUjYSG1/X+lSL6kyqsQrPCkaiDcRuHzAtzhFuXpgqYVL1zDjWxiu6KXKibDVRFTR
T+MFpSfvEbSHxplDiDIAufLqpR+V2LwRkbx93iVXEEJWCd3jgIFM+VWDwR2767ys
O6fq0CnywYxPB5VUYICQqvze8EFXWUgy3xW3ybtcWApk9q4OHjribLLX702GRRas
C5H2xOpugdGDps0OD8Xui5r+76Wd8K3ZL4qidA7Ir9C9IXE7WjZS/a4f57Drk8+e
44KUH3hiY9kmQSznHxzFd7f/NzH0rBwNvb3DcYN1E5Z0laRYxFX2VmW0bjlfTAPn
K7jFixVcrz8eeYIMpSbtJeXsZYsoq353xUWjAnZywcHRw7tR9Sq75rz90H3aqXBS
GyPmCeTR1wPtIA736dUS7QHyBBr7Z61fgxxxgMLg71nJ2x7/Oyh/IQTptxrQADFQ
8svCTqPVbPfamW02xj3pP0qful8sY6aH37FdWO8ArWZzBdFJardUF5nIRVGeSqbc
dJaZk2u122oZueio72cvBbPOlw6zNKRcoEmavdWZpafbmTff+T9XSU6fYAaSSua8
FRSvRkZc+CasvN4RkehUXcrz/5CrrywJuDMWf/Wxu297Q/ssT7D3K91kKvjIr6tH
JlFHsz0Xmgtaz6aGCjBZctfzv4bXMnF1ciMlb3BS6USRYh67d85vR0Bk2A+fiSX4
sL15P7VFaFzcXKwv+CkQ1BIIah14J1c0dCPaMOnNKw3iGwRXLnieVM7V9UHP1xM2
C6cIBQMKFHtbsYzRajzOzwVDgiZH39XnZsBLeNZPCut1gmuG43LRAE1uVOe7euCh
BNn7GjpvGorhM6tV+NC6cEsFb2ljeL684amrxwf+PKGO2uiCaEep29zyj9UMGEZk
4LlbQ1E33TgMty1QLREz46ULLpq8E1Jc17doGkNtGSzpSnAYp+lTV/AJd8l+gfSS
df0ejLzQX9/3q6C9bM8ek3+UDbBrXMSmT/4RM2u5UUtKnkGSbZdo1GRPIzjW2f38
eVA7AIuZRGIBSiwd0IbvRM/4hWvqgoCJFYuFf6cJmqkRfuSvMPHIWCdG98G9GRck
Oqo8iWG+4C+0dwvrCYid6NM8mbTJ5Y3NaWu9OGV4tZauDa/MMuJip3dIHoDCZ1MV
YZoduznMcZOQN9fPsnc8wq8BksH4fXsxCPGMusspg+xzRayZ6bY2+fS43vjNQMaK
RMZX0YngC7/J+io47iBjxCr8fXzcz1J36XWiuWpxN6y1b6rdIt0nQE3zLP/qy8U9
kCX3QPk+mTmqyvHvjfY4Z7L5jOmvElHPK/IzvFWsKgOS1YKTihhoE5V7GHbrhHCn
BSerIP7K+3gq4f8iSob9+LnnOC0ZlM2RbdvV10GfUlZ83ZEibuE/nnhXOgzWdI+r
fgYKxp6TOmUNEQbV+J9qTk7Hz3fEuGE7SLdcKrE51rUV5yps4D3nP5cYx33txA9K
rJI+lDz0vXrW7amgMRXln3iVfp24fymN5K+QWiUDo7bcjXH1KXWoYDOxp/PC4qmC
dHTwARnNYgIDMYn7eIDJOjXVng5IWeOQmBgNBmy6Scvj7NsaOr3cAv+kYlAwZMld
y0JeQuYdU7WEvyOnjZpqsm0Ak6o6HDFlB6iTLFNgHMq8aaJCZOQbuqWm4NCFod17
WW0E7uS9xx//u17r1wRpxsC650K3lsMg205cT6vAXxb0h0+9SGEr/V7CZKPOU/BN
/EkVcET5V3GMa9wuBXtWXQShJRBjseB1/WIyXJ8s2AWzuvRbm9hp+m6DSbOhG53U
3BM3Bg08gp2/RaoPrB+z4HQ98LzPY0IzVvvIGzuJKuycoQy/P1LGJM7XVYW3dF/h
yIRS1Zkqy1tiHoggPiTLxiUcfpjnY03BFD3AKGT/hr9Q2UcV5iJ6ejkrpeXo1wjF
7XeLvPothz0XhIY21eUb7PwT3jADj4zJslaTeC0XgpSC10qtAY56tR4AT3MVRFBj
2ysqbSCtC/YQX41iD+Lt5JC4uWfcD1+N7WPiEEOruQduwGUxKgP/Eo7xUBNUOKXu
2LFqX3XQ2BPobEnyv50qoZg5mg8Mp1+iB2FH30kDZ+AyNdUn64iM4D6CTZDj/J46
BClYusFlBgCYB9psjdCQsydg33S4+UXYf7KGaCSvvKFVGducOrl+POpJuBp8BnTY
IUOsC1M7uh+qYATDX5p672WJkPP2o4kliLo+4FanSid6YzHNTc/nKg3a860S7D7U
e7HXyH1XcFTOSIqXqGa306Xdl7/187D+dFV0MyzOjBiltt1T7unGz0enrJA/TdHo
m8OFFlwnzDUO4h26+YMpmFC59pCqoc2pzyB/bN+vremocvZrUyYkVVV4riOEfSez
qU8nMkXAwaCqYUbidUo2oYkaEww33KDXsXHJlzxkPSUHT4sDiZmNzBWiLPApcnip
dkgkFaKfbK8mjLP5Wuar7jtmcWDBIziakuMx6UJYZn347cvzajelxU2MV3E+mhrT
n19PNBv9HMBqZ+8UThFbh2iDxZOpFrxRkQRF7zD0KQxtFzbKz85Mh0amALiSot3e
Dys1zvuR4W91znj/r3ORJulI669RIzpXS4jqFfwsh6lS9r8ByPbtZ+pAVrXgl+B6
T+EfUC7etCCJ0S57G/9w2uxw9o2840RMx9Cf6TZDz7+Bn3ofVJfiPpAQBxFZehdF
lW1Q3Ap9+beouXzvbDHwxUKceDjeIwcJWJccZ2XY36NQ5BIzHYveDOkTdx9dZ7lz
l3hhSDYWkqMctPzfBkI0KZaqhqDBrFgYm1fZuTb7mDf4D80EUxPTour4YkyAyn2w
6MBtHtljvSaM7Bid0h3KZbNa2C3yiaRNMelG4UC0hALSO6hm+k3Lsar2XzaK+Tn6
Chha0wY5K8mqBLxJKcLrrKg1A/B/AkfVkn0LJchsPlXwFCpSlruIUFnQuGyFlz/+
zIJVQH8cfRCoq5xFpy34W0CoPThNiyX/qnk6ErsKM3msgCPbtw2cTjqhd4SEfg4w
fP5YSRxX1uLqB0UnT3KHKM4u/2K4d+xkI/ZC1B2oSEtXfnNb2cuRDVCXhkReEzPo
IjRJbsubZrfjWiltGAaJH/XnQ29UF3NDKARYB1tILs/SXwmH81TBWl4FCsImVOV7
EXsTfsJ0YYLAGNeLjryxE//TxUD+QMcSshXp8e/Bq3AUwbiI3PoWWcneEIKKcTsD
FhznOMlL8vdHmYt77w3YTU1EB8gbBLjvpJlCKeCUrjIDebwcDklqAOlL9RZLuh4I
fnyyD4zCuSXGvFFvy2aEc4MNSt0V8J1g112klxia+ck5c2xqkTGMPuweqCwjXw09
3zHxp+lL8nIYPItHQ4V4JLMy3JWvdE4X4FbRUnMB/XxYFKzFqUTxwOg8wbWYuKFq
vpoX/ZxZs5o2ay5y7cxfXaBxhoMxc4iR5T19KmcI3F4nARppaX4zl1/iP00NhaSZ
6ucYH5vZB2hgvcSmjJVH8n9FIyGo+Tzmij731JYGWJJCPU9QYpHSer6xvV3axYV6
GXfPjBZ4YlOJYc1NPtmyklNjGq0yVjvyzUnNaOef8YkG4vLvWwzMYXhmfFyU06Gl
RyYZy/CNnJ7O/3ui5xs0z31fD8Nfy5loGnBzEa7Zn+XWy7bS20A6+T+Y9dJiren+
jLY/WaGVehHPsTd3kkuaifRumrvdwtaxB/noEllSFKeKdSpB7hmpC5fUxD9Rziks
PcCMSOnPEFapFTpgosg9XKVUTdcjeHJM0t6VFgRyAQ4EWEJgv2YcfAZItf07rwHk
2r2MFKIWuDC2ZV8seq0UFMnQc7i3x/XJj3A3kgu45FH9br1X9QJ2queq7pmoIPGi
8FKB2xLmrbce/7QChQuxuwvW5g1ycA66jFw/ZGQ+d/aWP+75pGW309UvYlhvNAQ2
LvAopqmymBt/YlMX/QUBGY1v35wGFxNdXWbkGHqgT+SjV0rJ0NRY6NV4tgf3qYVE
XnZpEMPkngmoZHzKVAmcTBx0v+G4mhcw1M7y/wqakaZtY3W9AsMKbkTLS/LxA3NL
kUUNetM400CNinUXFUmFUVRObiVeb97VqLTDomXiWCnbZJ4hs2KVhcSoWG2sEcvN
sI2mXpFhb5k21PemNalfdHzVeq8St8Ba1cUaIIrEoI3957OTQCrIJe/hiY4KEG8l
IyGMNfX0aKfRtQjN2eLIBTgL/yXPNa+Q+ZSBLofmTnTYySS/ss80ctMjR0VIMDkf
z3Va4E63h7OwXV5JD9lcH8Ukb0CRCYQQIm8zT8NIQTCnW2nlsqY8HUhpyQ+W2k4o
bbBWkB95ij8dmoAP1Szc1bzrmXETeS8EdkYtd4awMYgbqE0o9jIiUwTfHvnJ/BsP
P4oQwWJqHD8pTdURvUrQ/ZBqJ4b+uVCdt4h4E4NeAMEQ/8O+i95LylCzA1ELszDJ
L8JQ37T1Te9SybeLZWcg1dgZvbTfgsV20wDj4NGnmPMi7VWPZOFU1AAeRMgHLXxI
BOjRmbffVtbx0oG3zHr0XbRcaQv3c8KT+ZCYoF/OZyeEcR2vX4YVSZFwSJ/ClG9e
70J3XdWb/tTZfy/p3WuS/nBJC46HNrw0J3MZX95oUn3DGFZQOmi8ykBz799kKSNU
uou/PqhU9DCv0sc18kBL6Oa8pDrZ1ZP3Ik0gQ3Tmn3529hA9jZRntBJMp1cP4FQt
kirx1U210Xgi09le/y3k8NiqtRvIeG76K86lvujFdYhE1C8A9SBJxuLFJfg8j071
o5XTETsgj5Yr97RWXvvVfj9mvwOdJ7WcY/Ikrqv3+5O0fJI19vnieyUmRWhcsRj1
qM957iA2jAf3xhEu9hHOZp5O0sUZQQolCAMJXtlH3ZEcPIxlpDVswE55W5lYvlxr
6hQYkgGqn74yiyS8D2ot5JdEQjyznC4jiBVZeqd2BJOLDDjeeORNoflSzoYHjO46
0EoMMe+dxbEqzLsy+yIi847cauK8GYJoeNIZjsYvqAf0T7F57pjpbqewWFfhh2rF
Si4RW70Ghe/dyPymt2EypM5AF4j5W9kpA4baADC6FZcUXbICS/KhPibpbSvaJ/Zu
gPqGs8jJN3qdnEGIlmFaXKs8yZ8t5dcHxk35EQCzvObgoyYfYhrRfzbkO1N9Ludb
5Qh0tWCBQlsi6bGNaRzq20gvcEW+CwZMUPPclFtWnqYLFOkqv+RMjjvU0HcOXVd5
VIknN5xncM9wwgmFfi5cNN3M0JN2W61UXp6xCnq9Lo8Z4kJ3dQIJbSCQEupjnOSj
FBBOTL+4XrhTSLxZ/rDKC5mzy/nFJODR0x/ha9nQbzG3xV2ShFg+oMX5xypCXeY5
Tr4ZpXCeTwU9IXE1jC25J+9NSX5yIrimYqdjrJhaw8Ajj6CZLDh48Xl5fSafvU9g
wEkW/uuRXiQ95fBhODO1qmEB5z5Vb42U7OXqQyoJUeDlCAMfGi4bTPuPTadVhBf4
1WF9jLiSMevsKNy2i44guZ5T6/j7gid2wweU7EyZp5JPdyjmDxav0lPerJhvCGcs
zCToE8yB6ZpGBVGnWzLgWSr6qtkDCHvxRGbVqgZeHo+yVedQcsiQc3Qe9MGpvhp4
rWMQAEazKjJhvetqQtpQ+/ZJ/56R8KR5+FjD40kU8Wp1vMUXWCSvDzhuIEwXBbE9
HuDdS/bjxVuUtB1OKkfFkNrf79dv8MTTVMaagr67wU/Ncrle4UZL5rUeB9f1WRig
B9Cjs2zA9RDzVmXzgIZ/9gxzsIJqNFbW4rqwb30JeN9LbdP5bQkkrAL6dD/g83p+
EXIN1IVMbB2RddD+/OSzBr+/x42wov4XaxLzPqSXKTCBNTtTtiyW/unNyAGO7kXb
krc8f4iMxaDw3IFb+IPZC2omCugwThdtxbzF5KyNvARMvjVMab/VtOSoqXNGKqnr
YFTiUREO80L2Ud3sZosuboAdoVwLV9owOloecZWuQXAA3BE5RBWu5ThgtlMXBQLP
n9rYl7pBsL2Hd5mA0jDnfINxvYb7FbF+M6WDuCptAn/B0rmCsQ/i0fdSFLbSlVyC
EHFEaRGYBd1Of6JZrSb3VdWE1OedYea3cWus/3Lnbww+DlBIDKzlXosSaMwyNQtv
MH+1acOKipVSoKvbWRYG33gmIINOL3TNceuPcgL4dgY8WM+mTV49Vpr/VY7w6D9r
KqeN4lT7fXkzrs/i45s7Idd32o5TW14xn9O2LovZF9rK/bZ+odXMtl7XpFYT9HnC
5MvpRKusavQDc64aql5ur77ziXInOuPHQTkRcjS//1ck4skaK29+IV5Mr1aXPlbv
OKHl/rh9uss/siwG2YKmPlIChVVW29vPeTHjdB2p0DMCJC3DGwDrL9+tXgRFdGwb
QdqX87R8DSVTRuV8j8OgADqDGRfqPXPuQ7yas4FPjkjNG1jhPY7fC4XDRCNknUvl
MFhnE6gfU8lpFP/s1mnTB93qBdxmtOV8Rq5XeKQcaozhu4uHleHXpvwuV+3Tm0Xi
W/hRRNVXI8nrj0Fnx37EcRe7AKiK4x3lsDwEVKomE8/98Xch6akDQcylF5T0CG36
d4PTBIFqGk/ar8olAasRacwUXDZWEze9xKBZLO5i9FSCoppsf2tQYXVFKlCYsFZN
0N4Eqs4CuTqliWcROqc+J5IfNOHVuMDQZgw8LodALHU6uMxvwFxA02sA4jQrl71M
8TLY7/pLdmLWn5Z3xvRuRVDLCTbjx2Pe5Y2WERirT5fn3oicYZo7Y5L3G0lXoeiA
9zxXq3g76uz3VfsryZPB9gTLBqc6QAq5vdfPEft/rcaIutv06L9CexJPwKb6obN+
YGNq4D1ddN77GHrAVTwcrsh8q140zghr0Ywy8xnZCK6YiEeBYXmgkCED2jCwJLd9
lEM71lmTtbTMERFYfDQ4kJ6oUsUAmssd+WZEhqFvq3TLfJJx71SW2O+D2BTBYOCA
t6iSWSGhu4PvX7MfPgkJbkjRlZEUnYpAk7+WgAgBL6qbfYFy55DErpKeh7C0xQCk
qmWoJ4OUe+tdnVtsriNAdIUAjJi9Q2r5edyNsRwvTRwfN/4YxyDg1eF8Odq8vYnm
ydsH0XpwQNyqmrUTfiouIc3DOMeM8UGnhmyPzFLew+zzi2q0L+Ffvp9Rltna+PHl
mh92g00TmyIQJDdzOx3GHCgSecluKuPvySh/NosXtjVexo6mlocQkQmwFu0uh9LG
xs3J5tIAWEBwj7ks3cBVDMgT9jpXomyfJdMHvPU9s4aBs+tj4XLdqwUlr/xm8jZx
XYivPH8655qwKgLKgXjDKnlEw2xYs+rhWoOG7ptB8WJgl07zgXg5Jgr6GZA5upeu
q7vSMMUDkp1v/nIowdsvySb7EnMe2pfjqjmrG0cXUqYkQFYlcYNSF2Fq7S3qG4LI
P6YTMFvzaseXvHSqtf11+Zm+KEhm2bE+nEMXQhFD/vEwVnKOzlUOOPb+6mX/IC41
H1owUwkXCZwhlfw/BCxGPotrt0cWU5t77qqd1KJNzy6MBDYGTV9ZQad4Y1Du6eww
HWNt3zdEZrKrxN4K5i03Fwhd50XxJHt9yQuLfAz5bKMqEpsQe/raoQ0Nxc4W9clF
3EThOr1qQXFwIutGn4TJEtE1A1blcgITG0pAB6nTtkAbXEpTsAgjZYo+NdKBN3Uf
aTIhA0tyLzggcgild7Rptkta03thYu7zEaC5FAjlD12HBmkai52WfyLsapjovRnt
mnDRbYXDR2W7MKv18LXkLqDK14D90RSSZkBy2E2gSvxNp5Gzr4/AwvAGum8lAsG2
5EfS7hPpVyzmoejadrSwC0Jfzz1W/fj7ozQTRnNm6D+yFTjYWxx4FvVa/gBmw9l0
q/o09xkFxwJUDfRPfCkFKd8samrxJiurZHqdkJ1uQy/ObogzJHfCDYWipSKndzt4
jrHkL6jq1JCBroHV3c04f9GRNCXaUa/CUDQoVJ8Bg56L+05BBVI+oix98vO0dwu7
qVTgdoDPQAomc7ZBJZAWbuy9+gw2sZLYGWFENOKCsrOagk1jjjnZDBY0SfGGuEMD
va66ClPoYpDdtpmiw9wRfAOLYRHm9DYTisDOesI2P5/Byb0RIXLDSdq1UNppawek
0l31BzTHLSLUzIZFx23Wx+8wNJtToG+USLP8fQ35Ku0dhQsYmrsbZl5wmf9e0fU6
3WCXkc0qFGWrRUCAlJUQSCBR287InxQy+aX+n+lu5j2dYHxRDZX1sCamR0W8ECtY
cYTpi8MmksFfE8wqea90DfjemVFM2PI5J5YmxEtEjACMK+OjcGYW2NUSt4U0ngZw
KbDUm00SBoYVepaQFMKFklRfZb14gEyRSTQxjtIkHWYDXl0p2oQiJktHjm32PqYg
nZiSuzEG1OZYssuK53oJDFQZLwQeujey3rPb+hfBCtcWsXTODNO2Z3B6V8freU3+
mN6s81LW6Se1ybPPoWeUrRpoRfEq6oK3S0toGDZURQktQ2RpUliN87zNWntwizI7
JVyu62aSPMN+KolBdasYA4m/n+NV9jnbnMfMYly4QWVOElRpHUAR/luTm6p/RsuB
3auyaa2z8JNK8OgnzPO4tNNbnxsogDd2FOeo5KpEZtTnME/SpFBw5dJzQoWfXFkW
yQYu+RNTbGxUceA9pkJ678656QBwywQFawdG652UPB1U43r3bIp+Cldae7KU6y/U
zwHd19xqOTK/VKId25oVKTe4qWjUlTl3j5F8hvql/22v2jE1XHZv9psAPka/Seui
4SClaU5RYgheKGGDQNhntqGugnZoCizdTKqhNk6zlKCiPmNn3Fqyb3kXkwPTQ4qv
nH0MHXyhEt0pqLDkkjS+UM7LNi773k0KrCy0iP+t8HO62WHHeZbXinI+2WGtasG1
4hiDxqs5yEcOcvMo+uFRsuLWdUGYRmRXhuFyS7FcrHs/t01lBLmn8etVAmQVDcYL
bMQp4NulKgS59hPOlA+8DzkP8MW6Pm8gtu+3QUK5+w2bp7TPQkYAq+70YSGvAsMe
aR9+zvvom5Sn3sZXc9fLs3fpLbxYLsk3HoDXPTp0fIVLygTBsNH6hUNk2i+2PsEZ
r2ww6eDpT5Uj052gFbBxo53ZUsXRn3lJG4SwNVQXqK80zDVsUfR9W6hIKAvlGk3v
gIgP0MY+1mXYW4pUREb7sSLOWbJyTx8GH+FXtm5Bb2bfcakeTPnPK2JFWW73SiZE
WKZhVJZmxPq5FKdZaxKqVxEcuLIUnCTjvFwUVNlOqEgP1P6Sbjf4xbqf/hmh6A1G
6TSsw3QklSsyFPv+GQLRhtwnGmSIk+cQlHKDkuHT4jujdJACyHXHL3bM+OY5FJqI
dLnSN7BYrKWwu1LqvnUgtuEmSiYiUengumE71gb9zTj4KxfObA+D/EhO/Ic1b8KV
QOsR5e2roORINt7naHcQJMQmEVhvcKpjlpdujKFrMuc+eMq65bqx+qmN7kan5af0
Ds9fNPkaXjU8cOdcfNfyT+DyuExopmtdpTz1mngqynS02fgy1CHxooV7uNRkLJbE
NF6RpC6HQFpgt6DoA9kOD4OQU5crPP9hk6NYBX8A8v0kuhDut3CkD0Mf8MeWX8Au
nBpX9sDPgf3wDzsjbqHu48tozMoGeM0BYApdMMdmw3IK4M9r3slNHeo+7Q9UNBgg
v99erVTIPEo4aJwL1NA7dTzCbPfHuEAym0WbLYqBfi1uCNstPCj7r8MIOnEeTlwQ
8GFB2P1iN6HIHoHu34awWrMjlqByrR9lPgffkSGx27TdxGRF+x1m7ECqTeoURO1e
bMEzUZ2eGFtzU93MG+RkUr7JmKsORsCUWgA6tyUzl7zBfxSyQSmnxOmNuprAszGr
YplKwv12LZ+8nLtwe9DD9o3aiUHWow2PvHLumRJlWCxgwSu2Hyb2i3kbaYSpaoJC
X+fsOB5bnt4ub8eNsFLif2eUeE8nfk5LlyD/eIbWvYfu9BHKIjColFYWisru/xdL
bIS1fWXsgVwxVha6JyqkWCi5tAukLeTFfpjmdS7XM6AYoKIbsPR8mhf8kqjhAxqN
fGzQE/6pzmzbUftqn6A4I2EDTpIZBj0BjLVW4xOqdazjKe0PAyGBRaU2ncT0DCNE
F5JLs0sEThjXEDdfLrStpSCj5VRU1DwwK2J2HUC77EbaU/nXgNwJHIJfiATjWChN
yOOfunX35gnljVC3qPcy6rgKHsqQgcKwmtJrlWz+rtJZ0r62STMCF4gKcfG/Mrly
05pSqjp7GwpOOYJxPDAuxTayCC+IOmdYXFsZGNdFTI/hzu3PdUzoW4F6N4X/L/HC
nIyYUB6Rt+PwaVZ/4PetV5wwPKUe/YsVMe6g1ObDNGS5IViHfF0+KsSX5WwFnFFq
VfL8xjJtv7+NGqevFhMbtV5z/3gdE+zcMDBZQdkHUNe70xxH0VI7/Xg6pgzaoUNo
Az8VGsKDuZCnmxUrI8ZNVPkhe2hVVNCrlMKhPspcX0zjCBaHQlB9oGnlJL5+KF/l
1LRuC1sWu6frWOM1u4p/hme5ueSKHTZUUkJLBnwHlLAdg54OPIG5dK8c+WLLVyUf
vEZRZLcgZoMPqTXeYOrKWiEtrNI7YL8Gg+CIAORZqncAYXVzyy1tRicgu/fnoyCZ
wIMe6KAZi/P9YIeyucjmtLQJI7MRSm0acFcGiTYLP12f/wXKXaJ1cSsCIbBDQd3O
JzXR4q6rAVCiMhox+e0UBD9qDr0PVkbDCqIIiwfjyy4yuAWYepfyXSZ+toFcDOVm
7VYQtH7b0oAZBpWK1KGMeHVofdxxpintMkzeMDDg+ipvLQnSKom5GlT+AV+qllyZ
3j26edxctw6o+S+GhmNqNX/2NT4MvYQsf3Ce76xwmj66lVRZ7rrQcycKE9EdXwwL
SEFqdSWuyWtApC042F357taTZ0JR45IL6E2+4wsMrI4VYz4/9k+0lNyD1HIR+uv2
EJb+rdZKWwwxgd9W8CeNyPuyvB5Fxw3RiPMDDheIYMxzJmv5JDNE/HHX+QVVr40T
UWCEwcZq7ZqFYZQNIW3hu/li51UqDTYMV2LOv7wtmoBJRfNrYoZVASCsu7ubX+oO
QuL+b4MmPJPW7CjaanbbnsE4lEMubY3jXbgtBdasZOnIgHvr2sVt5TUKupbxEGc/
4LhL6Enhp9vs093gjwjBMGU3cvczPo9g+WOh5IK+0hmHHT6skgWxy73YJRreb3a/
cmGgefFaFn2poE7cuWb0Raos6YOzYEybyoUv5j7/L0mSh3uBr6RzsEmzZYWTmFij
wDX4Cn0YvdbDBdP8FpK6DjGKhtUvfPdTFFB9SInoYzu02yOkQQIyP9irKuF7Bjv5
oKyaIXK4rPSHHAWPDJuxedxy0TWbvUzbFWtrA0LjdKm3BPk0SO+ABKMNNoXJjzgc
MTYbCxM1+FOQYVxplb4Z9E4HzaUma8UX2c4kSF5aA8MN3pXAAvokGy/Z9H9AuxhQ
rSBf8oW72xzMyEJgL8FUNJN27+WYIRRhw1tPx9hs/BoxZl5I4e+lXfyYTAyE5Dgh
3AJgDD5Zu6Tz5LvTgKk4EwOENsEdzhif15QC0FBvRZXyGpB6BNLp82OLpbGZSZPC
RNh0VUXvUfp5VaGQEdpSIvg9GANH26B/Ba+V3CJBD9wznHy3OYV/dDziAFGe7gZs
pKf8wLWTFjVxomDhpHzCbuA5GU9orrWFLaxK7E/3TqMH4IwV3W444IXHcnD2oSIk
NRseC/ByjuCbKgxjsmgy7SUnaG+Yd61dIZRMZ0DM/KvFXaYg4hbeNxQvH4j4Hm+2
mHlg9RS11IurMb6FiLDIVwGUkWe3jBiD9H8T8s3CurFxK+71ZTfDBSJbfHb4thbE
X4SEs/0SUfLDD+KB3NFh3N9OY7z0JSGv9oko24VH+2XPUA1ZgRpnNuZFks1dChsd
NsC5KnbuEt7h7mzEza0Av5EQOEBYF+sdiKPr8fQ2/t+VklaCf4zgKtFsLg89YhmV
bSyot7TTCTiySgq/1d12w9sSkOznsNKCY8onWkzXeJsxJl/lcdHIjp4wAJdqZVFw
nop+wyDnKMyffPl7wGjDzQPj4+YoN7monnmHPhNN4xdE1PXbR6C38PtD28cBNFOP
sxUvLh/MMHVYYawYm4zMagakRkD5sza6fEzFwGirZe79JgiTODNETSHZ3MdH8a+H
LeCD0hA8AE6o0OsWqAyzAMhUg9/SW7g5ITpHTAY/Vyz3wBcemHrmSIyKJdlaYWcz
AF6YL/VvMpTHnap4BXA7I8hkNBlbK5kFVfCk8EZKAcZ1k/N3381een8K0yRzTEBG
G2Imy82xEn//2QXXHyQEOU7EldaytN5smLZUnJvdeJRPEr1nSsP3dAikYVjDX5Ep
sGuMLsG+OlLOelBPeAsvaObL2bNjQKlg2PX275fL/3Dp/jFM1LtSdSXIUM1b7r0X
NuVU3p4RY/VsoGRgkmHrkhT9HrRYEIWeqhia6lvIjyW0Ul64Rws2pO+xfGEWOj2R
8i58qiAs0V33iW4JA6SuTWvaUZjUOPQ93Ps3o4SYAGLbJ8JvBom4UOobznS1BQrQ
kudW1agnqpXkbSah+16I6sXzOnfSx+SvdyIY8cX/QcQGYFrDQQOECRi4h43YJWxd
LNq83lzSEmz9nKL9xwloirq2LUBmVjd3f63dAeH4S2IrqXU0wY0G4HmgCegL+z2I
Ag8rUi8BO5+Avms7wbunokolwEjq0TNP7pyBMvIKThTGy0dSeBCpR2oZgqf9Xmyo
PLfmjfYc7vN49EnfzvSAZLGHSEQdW+V7V0uu1TUEm5fqHO3fhFXFWNpSBj0MH4Od
IxybO433fzNwedIwDb64dfGGtdIowiPvKqHcWpnmJaoWs/mbc3ftpGn3vkEoqtEB
tR+H9HAlerVVVLUwBT3tmYRebVSyIOFyZoDXJ6cc63bndkZZMfEkiBYHg8MNfe3+
ZCeQ+FrNdU7FXjmR7JGjONUYanZfTY2SqXAvLuj0MRUbENOLPRLdRndxZ+P84uOK
4y261uKBOqfVtx4CGbRrU2ocRcTHHahEQBb2f/nb9xdZYrCDFgBkyRKqkGUzhUge
ay/3yOfmyYDJkiG+hb+uZyvnFJbTofxR1s1rI55+fdsT9EU3Br3YuZ7QdX3kgXGy
lvXilJnMPa3w4D1wQhmCYKme+dJHJ9lpp3H6p32eWnkbklVO9S5bqfiyA1FRQlF3
OIAc4lao79c/6YuzwS+J3JIcADba6CXu0/cugppxtLjhgBW+KcHui7tuUxf44s1m
d6F53KCd1M/bFdiCbiUk8kjDzF0JCfniBO2elR3g/4CkED5UBR06T/zCOKl94kq0
SSnbGKAEKtXfkK4OJbdVPOQJIl1hL/QaPk/Mxg3T5DrDQj1hfOIbpV3nOgvJXsOc
7fP7+VPnZQv9tGr3iIU/vKQQyOyAnDCU5cNI71Jd9IGaUoA8BrM0mKLQFTxBBekU
5yIEUcbHmWmWN9bFDRjMtYKEoHaObVPeY5Lld28h9V3FOwDwBu6MG9Gwnx51cLfm
kJhP6SyNMLGHWqr1VnLmu7j9acPeTgdtH8U1gYb4pTvAwZw8bH6FiZijuZCdu0K6
U2nKY0rp+ZGCFojgRKBmIMt8rT9TH1muBDkN1QrYfLu4RB4B/y7zYsANtSf5OiI8
bn+U8RS3pFOBAzPS8RiGtaVZ/mlvR7lt9SpwTPwqcaaklUNpAxxUREeDZ/LejWKZ
/DjK241Wq7NVwBdXzJjZZ7y1qTx3CQvmbLGxa78TwwHA0eax7Qaul1vSJRrGsn7R
G+Px+0yHKqCVnAOKQAxSFLOx/xULFCg3zr4a4D0bsAyHQVgLP/seHtr5n0usOsqG
zL34Gv9bAOpX+6FD+QR8ibZ5oQRLizMwjZR6l97oS774nH76gi/8sR9/Rb2X7Scf
0tWcXIxGn/DHoqrCk8b3g1hofOIMjYsbKJMOPE8lrnn8YU3KaF2iI/O98LCQkH5O
7riZWYO/X4KKhgbI8nuvJARaD7xMst6hoTEOiE9+sByVcJzo6n78TJjqoCia2ea+
1ku7ubBgRFBBTdPl/YBu36PbJ3FAxmZgbex1laumxLGeFeQZ+0agci9/Qu9sXGvG
v/3GLvBdowXgA1XFMvr47xGgEuhM4r5HoBlT2ySYHPnAMpc7jGd4M3dkl4Qnpytu
fr0MpGOvGtfJIW10h4qFFc7OalKtjP3R9uGlwWYOO2sDhtpLn0pqFiuWmsa7Buk7
vZtXdD6zPa8S1AKZcWjyjyb/NknFPJs4rUgrBgB2cWE0Xlm4nzCsL1RTSi+x5+zL
CJRdS4cRUg+nbt7gZNQ0KKvNgfXwSiD+sjen/lt+6QE/b3oGxHNw2JXgD1HmDF5q
Ggs49FQd5xlAqIMaou9ejpy6VkSpZXElyKkNpYp9pz8swlZLBECB4lXg8kqsKy+8
Don412Xs5Y/TkGoqmtb/R1Inpk/kp9L2J7dbSq5+W8WGsAUM0BOuOdcP8Dt4Qc3k
Hezi8jYTM3J8bKJmtlXrYmtYSkOsRCCMCFCWi02xqmDlj910Fqe+arraiJixBvg6
Sb/WFg/Ao4z1LOI4VPaT3x3XlF2cdFdto7vQZEUUSEwzj/Dy/zMVggWhj5Ph6dSE
Tu12JHDB6RJrWpHEwW2oOFCX2+1CaEJcJ+tm5XTzkD/gsLKPW9btxPXu2r1bPexh
3uC8FUTNHoUp4Rp5oMAbUVtKzrx1wMylTnxpgmVUoc93ySjp/Zh22MHkzNfeqZ9+
WAdQd8c9A9Tp5tlZXip0ovpviwVOcjaJgBWEWPiv1xqBpFeUpqHBsNEZm6S8kGjt
0jCxr5PI87BvyMjVv1EOWbcJEj+fE3gnTmFH1QoWwvgDpeHXPQ9kdUFV7lfgH9yS
7yzxUa3QIw7D4kXA8E/l8cEBsVOkjRyiqA1O34cVSMOjOuUzYLGJS2XPv/Qk2jb0
2/Hix+9eCUDgSGrN4l8MqSkYvQyX2FuQvNvOJJNzGUxjGh6yzVHzEJWCtOF2epLb
xyFStrb2pLBgQm1mNGgqQG2v1s9q07hmVTugADdF/laivyw9jcBG5J2vDWwgo1FU
tEIH5Ifq/0fhK+oXEcmGAeUTN/Oc46w1QDiQu6eirB/RgLtAR7yT2nl1Fng+ND6j
0HPa1szZpTo/VEiQBmJNKjuTn8tooDu4OFQnsJFuYCdP2V2+kn5O4fP97SUM35xZ
KK7r9ZYla4rVFNo/JDqckoFgAvU2VfQid3ScUkriOGny0ew4o3B85ckbG37OUnwN
steRhNyTSanu+QFHMAtHuYgaBbaQ1eBrCv7YwFRGWfd3QRAQYnpWOVqWvtT6APjy
nQ2MTXT+Adoy+GMHZzpcVeU4F0I4C4LxqqboYAiJiiG/zIgXs3LjkppvnlZE/cEh
4eMISM2JRPwzI5FCrDg87WifV/NlmJLWPNZByaEQmxoUdLdTicrtUJD4w1fHwCl2
3MZLJf2ZKGUEuTPJ0mRrCnIAJ80t2Jo8Av2K6f/kJA1BGakDMxrozpIYfDYNqjrY
r1AurNsOevLp2jTjyygOHyQrBoAbZ7RzLPKpjumkqe2oYSIYTGVgkqneCTDyiEI3
ifxGNA43Rx/8ZH23MZQ1zNUWp0PyWsXN/KX0S3TUaMfmKD491nhdxgkyo/Hj1wC9
pyTVW6fK+wwMvSmu141Ub2w+EkJprjpF4y3j6/2xWurK50/6tHykokRIhpLoCjja
9gbn4R6kE7X/refKLZAEB1JYJ4A6ykKRMDrc3N044NUU2NcQfGPzMbeAfS4i/B7M
zmDBEl7z/u0tH/yQ9vq28e877Hk9HM99dP6I+f4SajKbUgOxe+4mADrHTvJOQHcL
fcniyHJBOytSriG2LOZ/PBn9SkglVBv+APURQ0nssoU8UgWs7BTof5f2lRbHIXRP
2NEpGM/KBIJK6LOl/UAkh6WVsMtDxdUjPdclYmOxVPnvM0C6BdJnKD87AayrwXJg
a9T899svICYP1wGuXHEKkfndlqJMg840fj89mGX+/S5z997BjIpwuBuhfS9TZY+F
YWqfP6o/+5OpncA+L1T49+JPUhFZXLnsX1Vh3fO9om57unl0VYU+Yzj6usi9A8t6
wJNw7e+pFoy2rv94RSkWLtnFXlIEnOHjqsNZtYkk92e3PV19IMo7I8GPrLpgbtbR
aBGmjwZjBLn5eezY9r/Ok+uTjmgVsojfYBAqxeNCSCcLabh9aWZmDcfID4I6K6Qx
Go4CtIJs6PMBaTe8vNOrUoItqdAcU36u+fwVBnqYP5k2o6t47jclpeFikt7rC95o
Ezx0yzCzR5nHXvzCLqKINodHPSl9Lx+bD9rNtYJZrfUL6LYlN6U1NQLqGh2IgOul
k/iqA/VPYgrKz4whal9CsG4ZXzD5OVjnuYhFdjiWE+hf+wZR55eLZd9+IsC6BWXQ
zfYIBugOXMJkykog+vSkfILTkUUL5/DPADYlyJejgXSi70xXK5iffbAONz0QTJ7F
pjNCvqUrTm/2yn8K6PHKmD08HSZK/RLf9DWSm+wvOagPv0fgiSsgSPV8HKmcgpO/
IxcvXz+88jrX+qOj0O53yh1uo/b3Zo9VRyfLFbRcE8wSgN0E2H/AErspdch4HAqT
ZgR0rC6xkjPmqHVOXAu17ufVO0JLXtVMUuUo7bH8Glsnjxva52j3N7ViVD57tthM
isCb7u1T7tP78ErDg3D/77iApAiVNt9c2s9snYHwqiwb4W/9HejfzLN1/xDFF3Mt
G9acrDA91WN39eLJS1Cw1tUBoA+qgTweUK1L9HGGwbecQ7+jX5MhsdeT1iHgpxie
qnoUkDj2OrFBYVMixx8tKfV0PBneKzSOl08FALKKNtn01N9rQAwUcuBf7+xURC4B
WCgkTblhs9ikp5wT9CWQ6cgch/LK2hFygiqyu28JA5NrOwcvoX2IAqUJJylbmsnA
NxQLnU5ic+4CHjhQrynSO6SLKfaqdAqhM0L3sHFOca/AeiO+BZmHrdm4O/WQhg0w
L6tvIkS8N5ADTtHp60lsEeDTZnD6XUBlktp2/FbDWdCbZEqwtGZJ8i1WQA84cWUx
MHFuLydIkYGqYRKyYTo95PYacANHdxOfxkcZxRj0b5JGhfQNfoV1NpKGkrAY+QNZ
/V+S3EWbNyHfQVgrEF0JYkujiK0MYNm3wpsc9APSsZ+TyZdjn+09gJvCR8kkMfjl
Mrk6+/6q3reNRoikEoZqQd/RP05JDey2BlQ93ms8Zg0btw7C5nZ3K7LkUj+Jybx/
87lFZ8VmeBkXWTC/Uu6S6WWM4vYK9Qoati5g9hAcvXDXDZxaSunCNYJ4rcFLo9O4
HQIapTn9Z+vvVQwJ94yATjYR/P1kHP4U00matHTF1pNbbmWpDcq9SZcOi27WrCwM
boSynR7Rdp2q8ki72tyeIxIQGaL+I1jdQyB27D2qlrNxTF4wewQmp6F+lG9EacZX
XnVkZL+oa0j15VrJb7pa2i3P4nt05Iayj0OSTOvfh8wRpghhk6xN2kmYSCxaPdmI
OH9nedJ7ahiFgUikkkOBHXx2s0P+vuAOogQ2KcMbqBH7kAVv420grTrjjitG+zbf
xfx3WaOfbTvixDvCtbKtZg+nGA+0rqNG9sC6JeTDK2mAbuRmx4Tyi+4C/yDmSilq
IvuJXbXBD+Us7vItrAtp+tbxIMFMaQpXGgO+9RyWe37/azx7PY0MMHulCoG1WoUx
TJNsSWp5v01FKtQS72ci2fA49jkvw8FvJib+4tZPydtaP4C24cIRnw6ZaqEYPcFm
lw1fFrPubfiUq28coZi+GrHqyLnjSBzThaVORZofNi6My4/4cBR9hgIxadj1eEkG
8X9PyicgfjmppS1+Nly68U4bEP7VqpyKyhYWnVnE8JUqzoHseJsLuZS1zmgq+oaq
UWBulCxplym061vtp8Kl2UAfH05ousTi93wj+DZt5ZKHbZQwSKDD6qTYLp7ZWyVR
HD11sxT+ex99HLwKt5Tyi17XULPf3vLd1yjN1gm276LRWpeieeyPUtJejoyUnXFF
+/sLu6bL9m5/IhkFa9UOmQEfSGNS8FyIsLpZ2O1hHmWxJ6LR79CpPxjm6tCvya/F
dugo7gP4C3+xFO/oBnf4EPHYF8gUZd/CsK2/FAWC9J4nQCCzzwEf7QzSi91qAJub
7RbBXDAjXqZRMPltpMQUuqLlvjUdSoNVjqK41DKwx1i150ybkAfTCZ3KcHe/u6Q6
oGaP3F0g2e+qyHeQuqn1EDQ193wqEQTFMYReoKBVrf1n1Qk12IBEc2KHmZw56Kae
CjTsVihQ/QfxL3sWLz5z6kTDRM71VG75hTq5pYhEOJPtu9afVlN5qgButlN+CXYk
PKzgiLUYMJtsgmU42M2MvIibU5ElJpHw/o5BC3l0PzK8FCaU0U8lX2tIrKakoHqs
1GnRyo8eDDQ3zuNUtK9hk/C5FQWjYKWSF7F3Sf0Ao86Ml8tAoDDuT0gl66d7MleD
0JurADE8w8X2IRSL9lriNGgsXXL0ODMm3ZBMYhXY0mxFNlAPKCPK3dA0kwvFi630
m8FDLzZHoFOAKLVyIsS9TdyIARi1ZSSdYO+n9tTJw4sOjPCuS4/VJ9JwL0K8QNaO
z2spSQPLZ7bPEAFwq6S6HmMmlldyCjQ3ML7fCX0KvR9jwLTLpTNQXwkYFE5sPJqG
Pqj8AEv7KDDlhcqE7jWMv15kmE4hDs+Dm/0seAJii/vRK+YyojZGkPKa/9Im1TfO
olgP0IZXFG6RS7NidyXJwyY+MtOyrRCKo5hf0EVRvveSvDKrHqArKfhloHuzkrg3
sz/Rx9Y75lRPI4pG5Es7ITSJH5w5pLyImRN7iHx6zPiB/CHXG6X2c6EmZpYcvzZJ
pOkL2c6iu3OjUFkjXU9Q1oEpIyiwkJe+/iZ3prELo+uHCv41pWodB0DrsfoXFRW2
j/V9eX8FRf2L8Oa9z45Gk2qBQCa++o/Kv4RewlIX+fjHd5+hiMVL8lDFelJNs6Lz
mv2i4guFMme081SswyxWjnw7zUTiu5y8d0+V0EaB9CIScPmxxPAptjxw0XjKEqCO
aODBEClYz0BwRVjapFzZUOpdM3FKQlsRn1NyB+lI5QJs8Cdkxzgid6Q0YJ2PaPUl
soTDiS3MA4T71xTLFB9DNFQjYDzk8Nyvk+UHgAQdPff+FxxHmKi1DF+823acInXL
wZu1SXL6uKAvg1HS3D6V4aio++OvKZ4VAq7R5AwxPep3OSk41OzbcAVWb0BTpMnh
zCY+Swe58e4EQ0QUwNDn52GwxsM6Tzq23a1DZGMlSeS5QmZ7czJPrr6/yxLTuXpq
wCn3q2X/i9eF9Pt+U4fOUS8Tk2lMshv+zQ5+0Yed5Bypv3EmZmHoKomVQ/lE65e9
E0Wxx5ARNS3Q6GRP1k08GeG8s1hvhdN2IRuBl8JTTJgg7dFZY/7aeagS21orB9Oe
Aw/b7Pj5VQUPSgqyKxtszrGI/bLlzn/xbpuIKUAb0XzvNeafG1ezVXLPodx18dc+
Bp5KksE6FCKPDG6boIuwK4ros+IRjdVjQguSeIX319C264Q0lkmtDPC4IKqOsabf
LbKjM9d0yoKPFfVgkVz0BN156T5WsgQEZuiBiKBGypZAznmNb+KYIV+paBaotL03
izCLQ5dTopWuuxlqAQaYKoGnS63VIn60HL6zc7YyxJ0HaexLKb9IoFA0kmx8nh+2
yVGZm+C78jkB94Bagpt80/CN0CByyKnH4Y5JCG+c/cm8dlUzL6Y9fDO+OS6iuplH
m15ByGqebDx/MIPitnqXFNhz91AS7ONUFEuscATaAVKXOvlWAGDv2TESl4oU0Hxj
Vv/vqF4Rn1ZF9980iJuy6+Mx32fEuyi2XhuLxD7+E2bFaLWMYBIU9ZW7KkKO5pkR
JxDQxMXHp4omvFwr1of7dvp8+RZg3LLXPVmlNcsPqJIPMuRGtHqOFUzlYAdqBeM3
rhlrHRYAdsZESf1KgGlLTGnc2Eod0H0DQ80k/kTT7FY3eLBqnCyDLkOWdgTWAKo6
v+R6PMl+rK6rv9aoqyDUIIAbzjNIzDsSWtAyZQcLTLGpI47T4dOOIThzsjfd+11c
HQCGQTKJcbSL7/MseuAQbEbMPMwOyYrkXVjodNuxtM75DXZu99LUzFgc8IouvRDA
QeG4BqSwKACuZUryNnfwDJpHw1wbrh18+eKva33BU7hw4fVIjwdk56uDA8qMIa3g
LyI2RwjlgkmhdfW/6+ZwJwF4upo9Chpw+QjfdTEGSws88Nnyj9Ys3uHeXf19sgfJ
mPZ0K9zZwh0ZZKxpOD55yMQkjLyK+wbm1ifApPHM/GvMv6sukA2pqOPVfiCfg64C
kvvi7itFkY2j8meEPTO9Sdd+7wXuE8FTD9V/JTTlAqEcdWwLEO3/LmVZ1GdLZPWE
3i44i21ZTjGzodS+yZhmLsPgOxRK5XrBuywx+BXUAnN1N0TQuyT0LrZo7EPljtvl
REfLmi0wGjNttwlIObzR1xXpAtHYqwfHQayfSeVLWKJRFS7EuY9mCuy0ciWv6mEk
L1W5yS2rGVbTtFLNq794YFlwQC8rM0zHu5hQadd+diY4c48SjmI5lpnY9zAiNaAp
4NPu+11ElnH3megXpUL+VgSph8SVKgEaWppHBsZMKTpSYPtgUq3bRsjmgrFHOyQp
Yept1/CLF02PGn5u+iSCBVAZ6+t2Egng+sR6sDzVpxpSYB55FeMyu8Vuaa+Nz+js
5iCf6upKRLVMWp/k6hzUp1e91AKLAiXpjk4+GiVkHg2i6rrqBlynpAQoyYD3N0QE
zrFKWO7TJjDNEAKDZAk1JzjA8naZAIzR+fFdHZwmaXOetUutcJjlAjEb8qvZB4zS
5hH9P0iLFcXX90ZEAfDkeicJ28OIdMbACOXKfZ3tpQia5unXa6byrVtwCuWLUaJB
IouHRkf/6qG1itMsY75f9M4DqwuJt7OOV9tOD3rSJMno9xlUmVUSTu8XuzB1jyo0
qjxBdhWUiSkM6+t2RzAaXliRgQhohc0+K9XK34Wa1jrGYZ7xD9KgBRHLjVrnqHAu
/ro9WxDHZSWH+J7E7NCTz5ManBl59z+7smeXK4cIBvpBW6x6fr+zxMyQiQ9nQl2V
CBPqKuZ2Bo0osos4bjAemB5QFiUjjOi6Fgrx12PBPnaY6PDmGZwlIsnnCHUGuL3V
6loNZh9CxRcPCYLDQz7DL/K2dnyDGH04O8XmtBv+XCs7vtvI7SpfUMWhZUNeKoIN
+Im9eyq8UA7Z7Pn7uD1Tgm0oaUbusO2exASjY5OlYtf85JwSopaQgIVLhJhGNkqT
1u1YVdrVBoH/FAo3aWIhYb6n/7fVztRNo/IzdgoTtxPV0+fk65U6p2/N1nFxcDlJ
+LA3K41aHZu0OsR+u0dpYDJCs7HTlSr+Kv+M7iTxEqQR2hhS4UJviatTovo5meXx
x5MAM5TP7x47R8UIj+jsBAyTgV1T8bdrl5VG1IUZcAcDvQD1CyFs7Iao4BJ5g4bZ
WAFrufwiB6aVPXkX0V7hn+nldGUTpE/sen2cfoAdcJRfKy8s0kuPQ5xDpT/5Ie+K
2yT9U8iqDW2jankEOKWPlRn1dXBov8iDp/YOPh7nFMZxO7lrlfVqXrGKoyZ3vsnm
KlSfb4L1WLLwccfaPHbdFYChMzkcg87FHJmDkguRB2MMbzxXCe+GhJZLVg7iqsHM
GTMYd0s8T4CiDhgJuRDZxSe5iaWGGKNjKlUuL8f2ysI22YEefUr1ckWvWz1BHLeS
6ILrLDOuUkQ01tqFxEq0YngdsJPnhK0q0Y9Cuj1gsG5Mku/h2JHz0bO81xGN58Fs
qTOIS5JUe47Xz6XpBUBuHTc42iqJhJ6BTLa1hwB4VphgfkUmMq/VITnk526B6tEE
CsYqASkjiZOAIX+0Aui6lWjgDvNeTN7zfL5My2ahThkRftIf9wh0peSNtucjjEsL
jPixptJgSDhZLVM6UD3c1s+MqS049ZYp1rxsOuUa6VNcG2PWW838rGEKmxAtgliY
J7dM+XELKthXn7jYhqSFU+EfrtAHzfoQ8roUkqp9+9mDwOKfHKBtoivoPtIhPeWv
CrJdgmPkQKNUPthEXJUSzEPxWNNzg3fqvi+gqvC1mmxJwSeJhWrLCVCCPYGWxKaR
TT/yBPrdlwh57wt5gLpgRw8m86f0zEvZXfUUM/ly/lgTBF7sJiY2mHItTy/UfhwB
OThly4dpEAtelxWWz7MQlrWfd8Zt2PeV8W/pR7pfqV6Vb8GUg0NUdKJB2XKoQIfk
OzfTjDfjSfTxKmosxkRxKrvH3DQMjNGB6Ha8bejyvVYhzzRURf/jO0Ap6jBrdVSI
xulVNAi9rEtRDI/GUMUTA/WLpVLV5UpdZpiBAEETeSSrRSi27UzaIXSp4Lq20NKp
5ckHKx2QoIBrQ9et8czBP596tqZfkNjFHmG2k5nplmzypNPDlm64AeqyE2Cweegy
1Wf5XnDQOMzYHxxnXMiHt6OEj0MwtMyEzoKYWk9Jic1xavgc1BT4V0o5+T8WjYXp
7RaeFUuIEz5t8VfzxLOZrTwzxRtyqAIjM7LegaELBW4KJVtisDIEcq/kdIqMfmw1
CimxuGwUd+EduxK21hvHWvYJ4FOTn51QXvKqjidsksj+gWbzv59qYHNjsaIMMABZ
GyQbR08NltRYiCKkdTmgV2mcngSYcrd2Oh3rju879SPY67ba5PZMFAFWciTkQ9PW
7Thf2G30mvQVpP46DLG2e68NFQRXSE8u6XlfVuP0Mj1RLxP5IwIgVPtGAvIx7fwR
3/JosmbFCkLr2rnf0KQFw0wIm+gI9QWkgXPzGQnlC2uCQFX5klzTwW8Ef/unfvzE
tOk0WhrrI//BD6cLOU9JxqPxUgv/7sADH0gAHGwptdNAz7Y5VQMX5PL0DCEQuuWu
d6yEaMuNUtLi1Z55GTpAQ8l516M/6IAVuox7JYYfFoLOmywKRF2PbbcusbrilhEX
p2apXJe5d7hHAzYMu8pT6kQ1QBhXavfqLqL4al56goTs8YlCG+G4xJh5oRAktJJo
liOmQkxF8jHD+V8iAwLQnWlLaE6HWhA1pFg5cTLTOruQ5qoYYo4Qcnf5KQuAcK0z
+ikDa/0mgQvid+s6lVGWsC83dBlvQ5VeUns0p5vsMaX8k9JAb1WRtb+aGOfjVqXy
CSYLDT0VoDqF513GPt5tPounH+7pgcg5DFRH6C5DTlz5wF22wxcolYQq5DO3+viT
+TxBhbeagQlainkxfU7+hkN2g3WGUrXoLm0aCExE9YSx2lxu3C87bJp5UErGSfid
0jk6xPW2C9ULfx3z2jevLYhXmj73MPoRkQCzcQXY/qnAWi6vmbCIMirHwqOq33pi
D8p8Gdc9k/3jXT47jzu8VZVlihon8GSSuSimK2eBkRsvnSg8FWOUe3mhW2ERwpBA
Ikz4sMTnSB8E9pAckcw5iWQi+/0I5QTZpB97xJIhJNuIyyeFyRsPm2eCsicg1qbi
s7yC2d3f2TrLvBzPgsrAE2g0bdRZB7VNeIWHwYHtyd4CtxoL19Lp17tvX2BdAK1H
aXa5VpGTvs6yvqmxUlSwbBsJo6GwfJOR/7B+c1GWSJdb+sNXppD6c9T+6qj8IQm0
EONGZv+483/ZBNPV/Vc+wFOrOYmr1ptbHbQbW8IDH0p/Va/hv0XAhO7K0tY82zZ9
mHoc8OS5J+DUYu3cyakvAhP/sPCLwAaxAMEbFt+wCLiFY4WR8+MtFgsl1bMdDVLe
gG5efWnfJm1uH+Ft6Wea1ug2dLJPNMHKG4IGAnYSsgFRIQLtk5k1aXVLWgLdgJLd
P0TOBP2/7bvm1bkclhL31zhhvNPp9UKpSC7fQiSAHuy6LHgdiQfQeqYml+4dpQCi
LxPPiq98AfiY3l0cUv2+uBVIlW/lT/UCw7B4O//9ooC6difO6awWWesA1G9h7ooi
pGpOv0SlQBWd16QdV+J/zyaUN5glJh2u+cZz9JSQ2mYVt2UjZeu3NbDsa3xyx0MD
aA6re5R3anR5i7nOH2J6zgo06U95B/fKK2rbyJMaU/XBtiSLsq3V86zGWoIZKdhG
PbBhmb04Aab/Q81yMkAm+5D3avgJ4KysjuU6BgOw+j1TlgiEpqbNP1LHEMQHOOO+
bvHEXW4MVUJ+VAZLO2pOV3np5ETvHlDTTT2oP3IQJQY/NQgbETc8knlhVPTokGM2
3qdq7ujh0HdMoBV/94QMM6O76ZY9TSLFfu/O+HHXSeBub2mswEkS87bOaxKt71iu
Db7DsOsJme85P1WaLpk8b3Z3Hpd512y33o+rXhJ6SmR5rCcwv8MWzGkrvH8RPn31
HEoaOBkmTkuJEQspiiHLecFYXHTghcUOEbvL+/ieWbfnqBb6oZbY5pzf2EuPi9PM
IVtidr1ZzaLQoYRmhIxXH4YfOVA5X7NB0e5mIbE9CUvin3nt75qSHfEIju2BUT1/
TQ0aEhv2K9MFIQ9MwXNBWWS8CQ/gKMjnPl8TjMuD1pbuN9XSbsf2vds3hT3cCtr2
/mxN4lmPZ5wKtBuLVmzO/QPBzpnYLDL5we1I5XysTWsGDmK23j/0CrrGZ0EvnWWe
OMTc59oNcm9iQn6P6scWVudZ4xzowxDp/P+9uJdhuisafx68MUDGXkr0jm8yjpis
aeOJiVRgc3bDG1zIrGcaycspJuppcnpSarpsI99ABOtjZgjtyiq+JK3QGTFPRdEN
jUczgafrZYMuh0oWt0CW6Dj+99mKRZwF3LTidwC0qBdWdwIaZXZ7tHD3wIVAvLHs
n4Bh2Kz+hS3vTiuu1S6xQbDD0+IsrCftd2nEDvmC11iR27SOMC+ZySRh/TE9vR4O
yZj1yvz/o4+G0IQiWN8uNo+AfgAry+GxWVRqxREscwKR60glUMldbYRFDLGqPhGv
2ZGyChKrc0egX5wxPj4aSjaplxdibIFd2JjpBRi+Kv4ZK8AtvLYRAwQDhLTRI922
99iqecG/yeFloWULiNQW1f4KZ9/DmR1fDKhlAq9Pj2oKs8niskctj5Ibjh2lBXkM
ckA0JeCg/0Ce96h9sSUiDfP7L1JI6z8HEx0pnZatuaMI94XBb8CKSXVRveFEmPbS
dTzN+ATs7xEfDe+PnltDHS8uYiRm0EAx0Yu4ZYGyDKY5pgrQJVZJZ8y/ZiUw1Ccr
0zurSh40N2Qq0SO3occdPCELGulcd/Kv1MvQEgA0uYhq+83R6eBrDLTBGd1T6Oip
zTjWfDg/USrlsU/5bC7Eel0HW11lmLLs6MHu3nj54K0gPg4eX60GH1W1K3Gr01vF
+mH2wU2LvZfw+5CrHHMSEUxXoqLSjhI9CMGNotPIzdSjcAv+kj5olDduoMzph7Ys
ekxVEK5vqL9MpbuhA+r6fVMmJUxzQbO9CAWH5wJjzvdvuVllNF8qg/sZ9H3rWQ2W
A5NUvjqK2daHERj44TLoqzZipKeKXsvQRgH49/FgqcHMU8IOclxGYE+segiRQJVy
qJ6vPj6QIKjwwh86710UrSdJhqU5pweSUoluEOyp/2OWhf07/Rnhm/s/XRcJNvBd
AYwlPpuIEhf54BpVIh4bRBOg5j8ukup61vgp7GmlntysBDpfLvga3QsX9gSMpoEq
F/HyyqYM+lv0DLYTY6QDm4ahIxLAWCfS+VSNgCSnAi7sULCZ4D7gTvTweSzlmqPF
bOey0La0xwUrrjbTI1l6mTYLHDd5OzPs3AH3x93PeyK4vKSJpgRXsNobN1UT7p0y
LSd28DOCMHesFNL4+4oek32JhBkTEYAtX1Ney7kS5T3CIWmvfx/2LRD4bKcdkUNQ
3sc79zDYsGlVl0L8DbaeVYEerDddWtpdC6CAmz8I69MQLrtZ+W0TQTCJmMk42f0Y
5AXAc2bH4dE/aaEjW5JlQc753S95yU6wqfLzw0FpQxayVxeon+5duEpwmh6L3nLL
TzyNklIicrbU7/2vi2ZF5M9BzbbnsewUr0fRiLXYOIgwZlRDf8zqIRdUTpMTS6uw
n4Mhd28l+d8SOl77RtSmbNlXjsPvZI3s5PMa0B2VaV77xHnObw3sqGS3/6+UT7Zw
L53qlZ57dA6qTxJQ0SKj++lD9H812521HEo1NqbxhdKRrn+4ENryvPJxCJS612EF
KjqC+xijnzb3qU8FXmWGewTP0jLLjVlYxed9aOkw7jgVM5vzSN+t4Eh2pP1L1e/e
dq5ytp9BHBXYJ0lQIlp4c54Cs4IkPFs1RkoQTjfcbTsrQzlThDQrYNqMNM83o8ya
R1KrtcGNgXNz9DfHJvVRkBxAhyRMzToJDabX7HdGNmX/tfmtJHcswem5gMMB/E6T
F4YJ9SBDrg4FcO/c++gsNRldQ4NUYdskCHT0n4IaC0AXEaOMdVJh0mFOuXts2y90
0F5NIbJbs7OJrP85APUVd0COW5BwHwGbG4nXcKuCnxrJhwJ0+igyu9lamCuIIcVA
552/ZNHoO89wPj7lJosk4uu+j3V209H7C8xv7Gp2KHc1DstGGv6ZplV/qPvlJwT6
f30xCUJRVmYCZWQoOfb6qQjxDYWFoUi0604uud3fFF1uLLQPAdLF0yMh+hi3M3+n
KC1+upIv1lYd3NK3UYgRKpkQIFNOVGL99fWXlEtLH98l1i0dM8d2SXJJ1sSxQtrx
3EJQU8ScYuQ6eCfh+yd4mvsTlk54Ky03eILA+KZ52gQljzoPA7htjbZvs3aJsq4R
oepWHHK/vMhGgo+HICnr4M1Kj53zcpZ2Tj6TD/E/V6XQmHbA5WGF3lmev+a4dABi
J9fUczFEK6RmxsohWqcgfE721wCSFKA8LXCrYTK5jAFvjaYOqr7Ch2kcGMuGUQ+q
0+aqgtGdK/wl5RdWNhT+3XroN0Xugd/Y0s462iyRndtfUGGw/rhth4qMz0uRJ6W/
4XBFHKXQCiln72MxeXcgtXRt7PL2TbAEAeTliPGuBeBdo+PlNH2Trz/elxvBchon
EvGNjpUU83zEKb82S4tQJvwU2h4eqfqsLZi1t1Jn8wGEL2tYt7BXiW0zEd51M5oR
ZcJFm0ew6Wo6YZZazgtJoUbWOIa5jn87OzCcsHN9vgBSWtRWzCTRB1Q79tI/cTuK
g9HRocwEjKgOTgg81mIJVB/q61He/1dIHtludUSviqmt7jnZscipTQ7+Yt3ZgPCF
jyD+6Sq83/LqcYXAyYvSsFaNTW0fw7zUEAQVwljwgpXg9CUmAmZDAP3j17GA2EWA
rl60MeF4+RaIEqjVftW7nHzdRFuMwfBdANbpxYu5bhxij/nZihg21uSDu7Ei1ju3
9ApSJduvHPsJlbnMNScvlEIX0PbGSBLoCizT4gp6jiB3kXEMNdUGLt6cYFI+ivVQ
0HeDY/z/qT0QYQ4fWouqkL3GYjr3HWLlw2Rn3s/sRZ2viW+xlLUfy1q9WamEyFXb
4Wg0QJl63n1uEC5v2cHvYpiARIJXTlWmuIoIWpk069VpVIwxGJ+y/H+kprM4y0c7
l8p5p4agajemZwTyPRwOQqdALB2Bzgw0tsGtArKnr3zlTa9BcAGzmhGTDOGS1ByX
Ao7j8SSHcDhxG2hc1hFVkN4wPb/CdO6/ZzGrxxqQUQ3pgDww51ypSYI+ysX4Cpin
mU+xOpffOpfxBZZ+lhE1d72o7EZ7qHNU8EadFpnywNGXSBBZTKMujrbDT4ECMHcu
6rUkdDumzXa7Qk05AVBqX53mZ4npN2nruJJ3+yCDJjFO3bU1QBgtr/RkaisBurEM
g08U2CSwmaikH3m5QQG1elZxyb4xh/5FOKhEs1Md2V045JBv0pw/u3DIUgmEA0M6
dI8+QwxAloxCyg/jtRlVoeJLmXR+I6zQL+ooEdLagcH61nwqz8YKoqx6TxgZ0lKX
66U6P5B7qcjb9nB1Wrce4iV00cpHntEsVtDqBGPuTzkGa+q12fzI6uMWScEZN85W
TiRBNmpL1jULff4tx+IVQ0/I1RVr0M92+2o8YOSFTUSBKJtBhIK8fRILkxfz8Ur7
jJ748ZHClIwhaZpJwJMhwA7xIDKzyVO47s/NXRHOwY/tu+qXPjD7t/4qJiEmFVxk
PvDKWGRrFXFIuITyjiW1i43zz+K4CgpFUadCzQ5zEt0Ki4dcyAYcE0tKBgbaFQsB
dJjyhUS8PJEGa1BidQsBFiUGXDzCBbU59gHjcw0OV/qwF3n6R0+pMCMouS2rfK4R
AceoqBn0Kw5FvvwOA72ean9l3kylvk1H7kwcRaTfO/EMAsqNAKkbdhDn2ACQWVF7
ioilh5Zh7FtOOzgoKzrOPI8LNr9IhAXTCbaCPzy+7CYyYO0pYES9eNK0ig3ciE3P
IPhX+HF0uItWsa9+xsz+sHSrmAXfml+zwlEzTH3egMrX0rvVC5hWb8B2Bwl4R+dD
Nz5PE2eK7Er40c6wJEtu6jxBh6sEkkDHRYuM72jF160dZiqvXw/NHWflUMhFNWX0
f9IDtwIVhS/45V3gkoRL6JBL3ancy4QmXDk8U/dZB1IZVRvtRnVOLaCuoTPnxrcn
Cf7bbSoZjOlgJ+ucTg9UZvq1N2GTFqDr29lQYsX/1S75evc6QNLcehjSsx0T10qm
NncBAC9O34VFXdenSZQ+xr81KkQ5lggMDKhyGeobsciW+LeHZR+wNvWIatPA84E8
wi5jJXwy73nhjUVvanUJBLGuVeEsmwBZ2igEbg73F8HMTfsm4ss6lLRtdiiPE/E1
wPHDPoOB2ZwO/lhrlVTEwOzeocu9rVNGaVOfcfREdMNBg9gW4xfNCf8XV+oho4mz
uv0nsJsOcVXrkmXciu4NvnyZsiym7CMEbe6jbPm1FHVhWwRr1T6KYAVYpnoh5pHW
ftmHMN/UcNLBsXQ46ecFOhz09VuN7CxUhNR5Shb4WaME9QW6WfEVRnRUQqVBZHPq
9GQi/3Xovvb//pp8Hy8Kxg/0/cIyMdGowDUO9ALCW1E5dONFY3bPMEZ/nX0W/pmt
RqBEQBdWGliCZI2wh51PSNosCECiIiy+SHU8bJoN6OBGGJZW9gO55I5zOOSpqolG
kZt+QZMmm+8DB1issU/Sps6eGXbOtbQ9Jn8TD8Dw9XK1/Hep5eNbPqKcvXnTvCnI
NPoCwC4oW0WLqrA2twmDI2odE3ZRXT8n7SJLKh6J/G2XXqTR2JqYIC69XbsJgMCB
5brUnH6FeyNWodloNFt1Z1V1rGiY7FD6h6vWXN3jQNE2ztbzv5G5LADYwO81wdZr
KE+xdyjvrINOqMzcsGx0Iis9wUDwghIh2e0a3LGE1jbUEWpJIY7gLZf94gmtFyLZ
mHf2U5cCdr0eVkdCxZilMDGXHxZ53anSias9kIJ4qcPvFqSpW/B7oJ6MTD2Uamr+
hRl8wXvnTkJ9tsie1cBQPsRa3PNgMvCv8dJxfKxm8IuTt6jznHJaNAPG9sYoInjh
6wCJSGL52P413Ovm1+sFlAZi5I74vdCUAFtrwk3lugN4U1M9biIX0VAt3SWWIOcc
udZCLR75dzRbxLJYwV4gzkdhc5I8Vu+nA23k9J+yBXYyciwVxdUEnhS3hnF2ssxP
vi/afMtiuixpqJthMdHyfHStQunDl12ctIs/DB7Yx/cMQaTVlcYEY3UnUnOLnxT+
57UGSffJzmEisZcEFpxs7gC/zFnu5heY2jc0btW0yXjMlLkUwFa+oeUHgRoLyKqX
zAr1o7GXsh5XSXLQ/d5AHAJl2lzGTVUzmdhzc64QPAGZR1kgbACM7r3fpYa2Dq+D
L77aqn9DuhvoNGsYtR4TLs+HbusWBVJk8oYrpPVVZmrHOytHMimV5SeEhxAiOo9k
r+vfeiUKVGZWvIlXHr07AshUCprUuP8NyjGMxOELDFSjDl0g7vv+o2EDLpPTeh0R
ulNwkh9G5KVEwMHTvCFgVs7xkW8OBcfTI/d1E85UqYLdgJhON+BGohja/sxEH/9Z
pirjFP0Fos9f1+nY8VJ/S1Mv3ShAeCnugLL0F04HLqp4cv2YH9cihn45RqFYouNz
2J2aqCQyg7+l3MALBHQ2NP52a2+MReJUJQUmljEfIZjSqN5kFcdMnpRTQUcyd74e
5BFy06blTTNKilFVPXh/8+1lIUSyP+5kzh0NraG4VlxsuLxX/nmJtPNE0xzL+ZOn
0bNG11RvFhUcQA2wCZK6mVE9pN381dEiZ8Hm9mCO4pKQLia0/cqOCWJJnRe2QF6j
oHQ0nV2bzAW1trrQAdDKNXLW+hthhkanWGLUkTA/fQJ6hNQgACq9zBKo5jD4IXff
KY9FHOIB+3Bvmy+XYZ6V1lWSzaAr2QWFy2moW8T8MozvN3oX5XAb8eg02RX4bRcC
UE1so5/BzePe6tWqKhv6iztnzviw1/yHUY95P2deqjCzLPVa7pmmJm1VRkhhcW6O
liJa7AL1lP+emVRmb/obYU1MRx8cCb2zQcvEKAmy3Dzbn62rC1YU5LoNbjIUXiCU
9n6z1QG02FGPFdfd/pp0dApxUh4ZQkva9uJ3L29WB7maG8K+C3R+HZ2YzaG8kehs
2Hfn+2ye5RO5+kqCIguILFD97xsbKYTwPxiQ24LJcs06I5LZt05ag4E26HSgUGtO
/QzSP1ABTJsUYQS9rqSHnSyQB/7ZhmCI5z62WoFhdQb8r7pIwhJpjgDz4iV0DeFk
d5Q/2EDymsUBGYM9xVh4+zaRSXvbmMFupy6oCFIHoipIIuEh/6A1kVl9sQPx+B6o
yHY5aA1bNztAKhJGuhfWWawbDtKH2mvqkdIan6fJoxRpUiuCSYLFSYu6Vyer8kbU
LbugYy1iQoD6MF3/oohJfIKpLd6zki55K9sAwQlwU5wDwlfIRQdfNhqw5ocUVmgB
S8L7xNW8rjkDkVcfvtqVkkk7LBG62iH0JOXN5MaPu4431GXZgPHcz3bNMiGImnbn
Y8qS2eUOBrYTTVwhZbtKknu7DjHkoQ4w2wgIa4X/YWV+97UcgPaYulHoXqk3+Upc
LL4sSzK/eRntm2/2nVEosSq87QTAM/SyzZh12KYg4qnLcfAKRnABJc75Q7Ohuesd
emBMTc/1xt+RqCoPUGeNcoW2qAPcMz1sHyNfI2cPI0I+KliTjgFygM/aP9TpgdM+
g2cO87eNPS7lSFAzszOn6ZRxYTVBzDQDiEEr6T7Rznla1KxJXAQPb96RM4v+PFeN
IE6DF5jy8lfFkAh+bGUEDRUhZkegMyeUR1+m7mVWUl32eutpxINqfZpJonwYlzOG
4+VcNkOwQwjtt+FgFc2YOhjV/toffOdUJVfWNYLmiULg8vJhjxBqmBSzZt4fbp26
vjEc0zuZ9xZOJbjWGDpG1WM1W0cOssIB4GpIirWP/y53PzeQo6LU02SxQ9naErhW
/zPnd8j9YG2D6AiYukkt19mBgyuIqqI/G7Q3rEuXPUH1YhS7roo0CtzWywWLIX2U
7L2yknN5PDqJuDiRMY2XyQ3hQyin/n51B+E1XHMRXKVdPNSYars8BtqwXexfmbcV
dV4vVtAAiRndiM5qN0TcJU9KwJyAPO2+YTneO0XZpYBmyCeby5bcBog3h1Jv+Mir
7xMSLInrpABx06skhHK9+BfHUIE/YqzK87hcFaejeWk6tLwxL2d1FJj/FHN6rPv3
YqD0nUo8i8ql08Z6OuNxGVL7R6ir9HPNwS0wli/QX5RiRVpXf7Tl8wuexQbKgbFm
FpRrNyTwJ0f48kAC5sJ1fVPvN2oLnEszPa6uXFbMWzDNg2KSQAR1KoME7IahNRwt
E2GLV/3tc3kuaUDF0msQuae6HFhvgBlXMiaUa+A93i3tY5u0NtndIy20IUXg0K2y
Q0l4VCfjTRonJqTVe/Z5eesZntXvRd8rSZ4hi1RYF6qAh0pGUa1jpSffKxDJjuCI
Xs5O8ZZa7GJ4hHn+JnkMDe47ozSICJ7XYumT0keJlQPYZwhK4+zy6HAkJbMcIfbD
2oTipLpTdIleaXLWRpnNRHp3WvKlhcVMb+pZ4/VZDaIdf05+nIjHPudvUZuV3W72
MrzIjZBFvJOU478T6+4rYas1CkO51Exdpg7Ww+ZvZ+/7Fgx/HbBbtG8etXUQLaSp
cixt7eztl/DzSB3usdf6cMa8hcIcE0mQeheYDr1XU3DZrNjueZ+RdcJ6d28Quup0
ZMBuL8qAaIzJy0Kmf22S0q5pae6kVwEa8foobcgZqiqthu26PxLItLr97StqS2UP
XRnMsHWtwO7Rd+kLKq+/447oCEgMlj4Z2mmd9hIp2ToB9e/DzSFj+/56/HTBlJv+
pAAkupX2mk8ya2tI84PCwvdk6Cl94Ai0NGw4jaSftRyjBNpCimEKKPcQ1Mo1UYOB
xlLrOxyUzSJ/ff9KyISObeIxFbarg/U3G/mTJTuewxlNxPLeclVZM4dtL89Of/4I
AMFi7cUiCdoEaTd8cqmxhOwjM6DVK6AzCWXAKdbF9ny6jxvxUk0R+quUpqlJIOBZ
3SJQZdz/rKlB9fQz7dTvFr7Fs5FJUSGUKe7HGaLZ/TiIWsGmshFFlpoD2ykcDbhl
sjBYajgPESWa6HO/lOmV2uVN2dNuo7wz0lAm5kSm0PBxf0NoxogAyCRJYxoRg4xB
YVddsLWqAaAEbH6sBEpUxmb7rFVkR/6jC52wAAIZF2Alpki+a2NBStpV3yUf0M/t
DIFHKUg0W9QE8PZ0vJ4ocA2KqTE+qs/R8vzciuH4G4XZ+J4jneouZ9qAp1PojCRb
60FcGfmYxw6nS27mZ1fFBt/8BZ9/i8Jj35zaOSKoJBgvSGkYmg5sl7ko7XAwy60J
qQOGKEG6NSNIpS+6TxJRjjDao60G85e2cYdhUkhsxZaFeVWPes++Xe7ES0XPxISf
9BE7+915mSFFR5gdYmQ/Dl3bhLdULjL231/QUwP8R9WwNlmrd7r7hpuNaa4J4Z4q
LCg2sn+1wtIIMYpc+gtVxmvPsjnS5o0Lg6b7vLWvqmOGuwLexvO5/+0KcOXLQ/Hk
2t0U7z415BRZnxlfg42aH8kUsOmbYCy6jAkxlQxGVtf6sm7+Rpr1uMrKdreH9+Ny
ey9hjjJHF0cdihoz66Ww+MDKAoREpkJbhBgqsvyyW2Ry23tvx9u/i4KkmZIXikat
+BX2k2D8DSeYNsRtJWzi1GWtaNKEhDDJaNaeKKHL/VWyKcBPrEyh71DmSySckScH
ZZex6oNzVescI79snJUf5mh7CtLuf3ezQaYpCyO+zG/vYVBw/NteV13JSXJx6/xw
0MNJP70S3Bm0Q0Q8w0VCnstvUiUSawufxh23FSoxVjqxMHwqxAjKEmmph770Cutg
PrHptSPGlmTlDdLXqgK9LDBUzJbPdXD3IwVuV4O6hNn44PQocKqqSTyY3oNed5mc
Cu7OrO54brODlo4OiLLq5+3D/037KotWhuc5/xWHVKjLFed2tPw5pye+7l14I6pH
4fyLhe0IBDI4bAy8RQkK3GSqpfzPSfIIlTflKk5uI4r3MJegAM0ucK2v8/WOnR2z
QpwiIJQnlO0udWjSJ6HeU19CV4/CvGK9h1wAUEerpTM8Bo2cT3DYzXaCr82ujt7E
MhJBsgJTcM8Bzl8ezL2XF0OwSLNvkAwLp5UxHw+v/3a/GcN+0YahTHlf6LefIWCM
VXWaTOQTle3ELR1JW8tOSV+V8sYXs0fvPLxNoZA5Vu/LAomkW/4XPvE8ceVurY+A
sZjiDa1SEAiCDkm7l0t2c7rZU5pBpJbPOA/xobcZMNCKZVgJp6Fqp6Nes3dfezA2
BlvGzHA5zzHPml3fyzwyZj5dSOzIu3YDjBhppsOywerfi7Dy4TU9N1UjXNRrR/CM
xCGr/N8iS2z+wIdmfLRViwBxsnlZuxVMqM5ruexLajeU1Cd4qWL3imHAIksdrVEa
/GISNnwNmMbuQmOZdbBbCBZDozFNWW8KGVDyZuE/hij+HRq1MLPl3HH15XLqdWxA
qM6cksbLV98YUi8e805T22pNqAKrO+kT5B2cFkWINq2TGm0nWEgBhHX8I/aRWwOr
8kPn5NFAW+c4CaJXaFz1MD2SUoBZM1HRoFGSO43nWGPl1thVLt+MV/zwgKb0N6UA
YsSV1DkUYb/lDMxo4dpyRcsr6nWPWPt7UHvO7g6EqDwrTZQBncbEfa+Gen7NO0Cs
muic38YaJck+14O1X36p3ENcqcQXD83WP9DWfj3HfD9OroQY4Ly5jbYKnisVhL9v
CqlxUCLVN+5DXvTCiNQ/uAhXaurqceCq/fE8ALTEXUPBCJTXm0q4jIiNoCjiImke
UKkC7cVdPpSiWSlcD+Tw/8x4IQqqUEaznOh/wVayj893Kcc59k+PuTD/CCAlOZrZ
8xMfHpwx5Iabp1oDZU+AUdWo/SsZ2bVksIyn4s0+R2HupklmxwkcmBB7vDqbgKFG
K4dJ2CawYT0iPreD868NDEZB9zp/7RBn4hZ4SuUj4CzYee9vk9HdME6DFglZSQ4T
c5bulhKm2FwRjcdtftlDfNl075VfMW8tCpsbY+0iK+m8jSwxPajFWvdZ5xiJoDpS
TTtSrXIkj0PFdqkFMn9eA30SuBJLpnbUTKIClCIMxPqRI8Elxmm7Z2pgdSnm4Y5J
gyULO/tEt9cwdbeOzmjtMulq3bMVcIxE/fJAZBeVLUVvwDUewLHDWD+APK1jIsUe
ymFKo2qLZ3QSvSYuDvkJ5kaw83pEpAPM2D//x0ng3nQZYro8v+Zjov3jr8Tu4kuc
kCJBdGvtTIfcv23oq0vrtsKpq70dr964CC1UJbzBziDnAv4QUjjIh3KGhcDuCn5B
yvdb39sq+edIaVByDwwyLoYcuIhgJlgfR/Nrh0kdwdSS+ZGXwZrn0aMJNaUnr3hB
DhqjKQ3DuGPKHpcxhQ+RqwRfQkdegxCNnTVRo/O4qWDUV262iSAwXGOE44S+rCqz
L6fcbzob1gV/Uo2YlekjixNniknE+Xz+u+FnFmy2le6Y3RZw7K2nyvM0kZ009lUa
IMVPYHOW8ihd0opoi3t2ClmS7MOr3jCJ8tvS5o2i/Q0e8KCNfpEBd1iPaRB0YDLi
rDk1qQDrg1KwnhbunjUvRKcVdG2YczSynYOIsZQIOR/rOwyxhUXZJMWHabkgcAGV
Q+oP1mnhdDsC4RQx1+0fwVY8U7DSjFQ3Ri6bUeKwsoPCqDHHKUN5/4oXeFSQOC33
mInFLP/IViMkEMmcp5ZXZsUonQ/m3LHQMesjXOsFncwUBO+vADgdLMdz2/IvHUSc
wWo7lVg6NCaagkBfOFMlpzq/S3AoIVTzoa9EJuktB9MgBSuB31FOHdGzGrJ2HZuN
+8fG1tOrfCjlKO/VV0Npii+iGPbLRSJHYMcyLw7ksXgZ+SSkpGfD6bp0jNAVLwwP
0souf8gKS3NMycx12HlxKjYNFvbijuymXPPxF1m5px+Qa4m4s729pyqb1PbchXEy
tebCbQ0QT/8r0urvpubJnNhma/y7u07J0r74HjmQIqFu+0XQxjYa1kfZdDl25k/D
Qz5x+3jrlZDBMpp+lHyKm28otqzh36eyq0AvdyA/fq5x7RtWLcqE1SCou0ZzAg5E
9Gnv7IJPE3thg+iYHPpUQ21z5Lo7fXwOTqSCSV6m2d2p77hRJTBkC3Xc6mMIu6zL
aV0fQCTTYIqiTRvdr3qkqqcuEQUW3dIObR19QlXvJwuNVM3oXC2VTDNJgHIvAcfD
Myub8P2es81Yu66dQ6Uh70+1kJjDojOHJqveY5byCexQ3QodGUXOw6x+6E7lu5KQ
DA4d/lf03WVsHn6mJaoeVGhkb2s06B0TeP3CFKxu1/+/1FeBWb5CC9JnWCQEE2Zy
26MBROxR9i70ZF4jQbGzrs70Azjin+k/XNB7PRO62/RF7YJUpbOwz0pTVP+GxNY+
bKgY+RT/EGzlhZS9W7vCiNci1NVj1LmuxZm1OK/i7JrIJnoi5MV1P+9uqFQfbuJH
aE201KpgLoPlg+3YHN6wX3raquh2XTy3YIqj0uGFfMPF+bt/IY3fu50YuKYD8BA5
wbFCPhw5+zCI1HPosAg3UhugJsMd9GDfmlR4XZYR6XpaSs2xGhQBOOE/N7HEfgrW
hP9m8ExWd230mrlk40z6EVxcuQRqsqI8t/pr0ZGmo+kip39DAFUvE1EG8+MEj1aC
UXA2gtJdH+E3Y/mDVQzS6mlt8xN6FGgKuNUtbfqx2odf0XUx9TwswAeGl75SwZTq
lzvtVNGPmwpKJCWh+jw7GCWWPAXdjfu17D0c2VLVtmNAapxf3EQP/Ij1Im3hUIf2
GeDU6zJ0x7W+wsVuY48xy92CtEttHYPno2KOfmj7xwYByDikUw8nk/S+gzxgnJsh
FD17Mb/LIrRJqpcTFxxi8KuYShEjplwB1gtxb1Czx4gX0MrYnFm+6uyHme816/7Z
2fYHKAVQkSx9+2nBnY1j8pqQA1oGtsySJmgeF4LRf4RQeINFYHyjEeGUucxzE2xm
1rksVg9pNLeBuchU5VxlPKFaWb7sQqxHDrl2vG27nVVpUGcuK9Y6eI/8xGKwl55a
OoTOLGYVMXKh7HMsl+iRDvqP32HWpb2Iy+nSDsKR/eyKTMuWRygf8Kfv7KlUETCJ
VuVnTs1qjaI5Nk7kujl5o8A+A8GrL/5cvet0LvRklEpt0bbXxXRqLEkDMmV7fXpi
ikDH4A7W4uzwKTfj0/UBsn6okmdyBjwpghbcqDWEhR/7t/EHp3h2OWhRY6r6B1x+
ebShSK8csZGR13IRzBeIxbrrrKuX/bGixo4qs5H2gzWOvuck/8qQfCzkOtZl7Qzw
hXOlnHEzpwaxRkrRCAu4+qIsVSK1A5gwmNaZnsWNlg2dagd1CyNzPUrxmm+srlHB
Fk8Aj0bOZLGX4DEpm+OPo5G7D6Rg923w/usuvAEMmM3axJ0MjJstsIJ2NgoqAwlg
B6/2Oy9uOoWaO17xLj44J3EijxS9cLkhvSq4sc9buzA1AcT4/pTux0HkgaeLld9Q
brKWwrZUZlPvIJu4mPLfXKBwm8GkllhZM1Ip3Va/1Xq/dftUCYS8mkQfvp0hElli
X7pbA8KX6qoPWhAYd/2V+s+P90Ih3jQuh/7cWukIk4LhcxMCCS/1Q/rCmlrLIXgW
LIqmMXsINASgF4YJeWFmrGDel8wv0VekQVC7qNVK/1NO74zQPa7huRrAbdMsz19A
wA/az77zVaxuqoCD1LJswDCni28oS595UGzAMZd0eJt0+RY7T/RYN34gJAZWW9rQ
Ao7DFFyvjZkTOJRexb8a4sV+h0CvZnQ4m8AbyRpcGCu3qBdxG0QttYSnYxzZoSH+
AsxMj4BFRSP7+PnCRmZPjAhu/veAgldNDNxCLktricRlVRMf/9Th6aIw30x83tpd
x/l4Fyv3029hngfGzyl/RBlAEXXvga2oVePHTGZ17lwVU5RYhV6RC832wYj9/GbK
FRL+uSKL8lNPkSiylhiRhPAWdj/KpCmuiy7uUVIzBR0R6NibUTkGU4IqO43p5mqU
MdJnir/AZEDWxjELWd7vM3wKw+kycrg3CcY4nW7dfbCJNc1Cou3dAa+md1z+eL2Z
gpFc9rBFj0XKnoCf/JhHB7K/z/uylIkZ5+NCORtmaJnB3LYNoLdpc9HTKeQpXWcE
0fe3jxkgb0941+MWrq0Z+vjAf92lV2oEcR8kV8DmszobE2OTTGusOoakVnsxnYU7
hg+XQV/2KGyDGgQOMPbU0n2gxlUWAip8vBBsudfICiAqVXeTTpY54KIQCo7OvXQR
Y2WE+5qysy6Pp0PfYy9uzh5eXbQxwrJ7bHqlMRfn64BQDUYfW5rW6NACbFkKZSQt
8g9OX0CrTNxmPeENIG+1RmBW3EbCgnUn5mu7x3UxPpO0278/voxRZDUgSd6fdOmD
6B4PXUnKGuSexZ1IJzqao/PDz4Fd7juI1lL6UWfRTK2EJd4CKgpxY2hUsT+R/Z3F
qij72mpIfBmBafbzqu7fNhekI3aq5yziObnqxTWt6sv9EHtoikRGGB3bct6VWx4a
tCXRKP3FIB3U+XO9t+wrnWc4tSkqP+qczfDqGGd/8DRfNbiz/1tgXyXjHDJaCeds
rwc71nbuVyYRHXqzg8L9QEz0mM/jx7g51DAAP36lJwEyUvQLY0kP1p676bUXYnux
DhqRfLHWU4dhzSNBu5tXwrg92tAEdMIds+oWdFDrxDBTx/9Fo1YEVmjLaFm/qQVX
Cf5HU25qEL7eh31NKhySNxKCwRcScngQl0KxlRLrIyw8Ivb3RVOzKyhhwhBVqMZo
HZmeuxfDiA6ZtyCqehWkzQCTfz1WguSH+Z0Wptyb9UZ926OMTJW7IEhMwwIg2lvL
4TQeF4p1kbq3Gyl4SNSj+1vQcRZzmoN4R9OPZ37WsCN4kvabjcibYhHl6e3n+Y8v
udpmm9STcAVB3aqhTHiwuLbWPDaCBGtT6Xu5PC43RtbLKmtf/skxdXWajh0XIGLM
0IYzb4GoSrMykDuQ/6F+5fejnVcbjIMPIKOiwrkAcKOjJP6U3q/B2uAAQc0Q+qks
XEJB7DlDhTvPOqB8MIH4qSX194MtXrn7EayYwuzA3NsJKGpIxPC6qOMj4yGnFJpF
/xH4HqfaIOHh15y/9P+Jv3uBa31kAD0B/6pzQ5c/lAdDjB+2qoq8L48k6Twj77Zu
QS94EYmHuLWzgGh3wIGenMIvkyHXkB1pyvRFLpbVaZYhbjdoBHx4PPNP44kLXlE4
jSICp2xnIUqCI4M9YBNfVOpPDXFMoDp7SBkpLPrEuiYypBLdwFnghuWWGNjMRszo
e/XYiTEdoBcrZjXY7soav05JbkE2Av9GG/uTlh+uxScIToL0XB2ieou+dMzTHySh
73I6ztipif79HucSXpKxpl/T/o1JnReEdJolQAddXQqJ8EHG8wB226uhJ2qcEPus
GUTX2Ud77qg9quWQeREc6+NS3TiqHRdzFkxzvqScYmdHQNxhuwh6LKyrWaPF/Qqe
Tj4tn3YppMfbSR4T6WGes1kpSF78iNUUfpzcwpyGMlLKlaRrhBpoziL1TvghYaDX
ux/L2DSCIdm/1v+hjAn6PAYfq0d7a7sHdoy7AqWtLNuXMoEqJ9Gm+aTer0C9ibbY
CMFcDHN44SlWfdfs9w6hcZqSrzFgyQf9lzWu6/Q2v6XDUtzZ5f6KwMEvAQPAl3/r
06VxgXbp/6SKUIlkyFZ//1vns2QouU6g+34ELDMTAdWSIgHvxCVggxJrRlHHqgEg
USSZoRbR39Mu885iuDNLkXEZLQv1gNbURVMNErdvrFXur4EK8sX892NoygsnLHsf
STQJT/7rUIdzS6Od844jIv2eDamJv2Ed+xeINIF/GE4qdPPxWr5FWD2DoYJrP+cM
jDGGG8dJOgMRpktfLurk+/TeLMo3FckIYqcVnFQMHGgXzDu/lHe+kD+lfD9JTLVy
lTS9ynCaM9AccebsefAUxzeVaIcnoF8UZcw9uJ98c27Ku1HLEntMkN+3zqZ8Mr7Y
kom/nWpM7tyX/ecA3sygSZnqIz0hTj4A8Tp1XiD7mHWUOrtVXudYaGtwbBP1A3Ag
8X0rnR7qAb87CyS2YngDe38g51Rby0pObGPYGEIwwVmOwHH+iCbiOMw6rEqNpsAI
YiNANKzc4HbST8o7OiHBlmjiI9HeZG70wVq/aWP4uZ8psz+dKO6yhEbAjytEXs9t
uwiiyGhBVMYCmKuy76w7m2ey1uQ8Op5CIF+3++6LS26JzuUxYCzrb8U1plZY00Sx
Ibu/YJTN5YrInEzc62WF/PniDWv/4UnjmCrKUjq7fQCbebnEzvAPrDnImOsjTUOu
EvzoSMHt+D661Sx2BzWYm+WqW1e7luCuon2Ty4Y55rmthewTUUd7hLUo0De11GIl
SQuUc7tvzjqTaG08apJhDX6wXBHRgr7oP/Y7gHgxMGi9CgvORmzGhpCKDJpHOHwV
RRszSNrT5ZcShNVMhdXsErgi5S3wTd/2Kt+cDAb2kUvujSylZjLfHQBeRl2QRLEd
Qa1p1dtEbTbezArF8axjqUTHFU7ORbqDYWAL9J8IybE62Vvo7YQeldzcbvuyDNt3
0Y7nArfgdWkcXTGVhH44ca9BKSBguG9VwPXnqCmrPxuINKPwTDzFcgjAKrFn+/Q8
oUIsdq/44uZ0x7TjFkgEIHrt6FosNbiwO7Wc6U/vGyrz7bB5F8ifoFLtTG00CizY
w9CYviqrPwZogAUjI8AhAEs9hDZM1RoKh/gCv0czMCvRczIiAm5JYY97hFTrH/+6
rA5aorYx8Qgmq1cETwenw+KHDhyp9QEYp30qrg+VlzHgvd7woL5JE4aZd0jjMbIr
cVC0Hht7mWEi7rPvUje3SH6G/GYA025GUL9WnFOkMzbpbvEhEA/GP3DmBFeiZfYg
l4L8/pSkZI/u4wIUO/7PwLpAZr0h0XNbdxFWvgu/z9DSI5eZSgmHtWOffWeoi53c
CUMzVzDPIZgyloI3LA1ra+fUX0WSze6xaSOLGDstp5cthcSPXl4cGwxwr+RzOD3X
0Gzub1jwkUwEbXwYS3UaJUdfKxf7mteJFI+h1Q8gxgQxVdcvVLCjF57EM0xYveHs
9xXeVKtS5KLqdTO78us3G1k+wdVEFlsNt0pPuYy81rtb0YGISlCfur2vF2LPTojG
B4nl+99+OYtpxV0dA0XbJnPpDR6cTxBKmpOIcPpQ+dC0p3JUJYWpOQSNF0lkYJBi
R9/cb8GqIFl5Ma5nN9TXI4eAMFpp2jKEyK6vsHyDsUaVJlkoz4/APmGnIZHGKxfs
/36BCDE5ac00lRvntLkZVgCfnXzDOPl+CHhBYQ/lRML+7XIbK6PwlDHDqvtB04nU
vBg/EB9q6tw/2hM809DxBCrZz7WRzmbbCaHFLVdrVCmmh60QS17OPGyOIxb80FOr
Ld5hKe0Fg8jys5JIrNQUYH0oMIF8MNV5WlYkq8KEQFYfkRo+FgXnItp8s8re8Yol
cANdp+1tg2D7JdQCRBP0lhYN0oeVz6lGug7i5Awa32saR5g8/Rq61QWdcuDRRlTE
rlClWuxCpx788hVN+ME+RvVjrmwyClc/nTFHGcpWcwPIA8odarpJmbkR3Ozjt2EC
OQlqcASgtgdmqArlgVG0ukUXRSJZ6z4lW/Lp8fLq4DKZpAKTU9xM2/AyU6k2Wc+M
5u3J8Sc5T50IzvK+hkCTao7j6QrwZN82t+4V8/72T3ioQLGKeDeLedn/U+Jx/Fn/
dMpuOhfuiB2Pvw2luOUkF3rI7+YaGBrewKVxA0ADyJzm1i20tZys4pTtb21zmMU9
bcFsL3PHzO9n9Dl1p21pxMwQ2IRh09A+/NJTti+O+fFqTEB4lI/Oau7o0jqxWnDm
psdYpNSmHVN4WxuNxCBH9mNVEEnxLjiY/7C0nlPxJV8sdDb+G7APxc/zZbwmuNLt
F8DJxZ6r5VWLK8qG2zpCfijGPRF4T/BWNVHhOqo5SHKKOTN4EVWwLt8hoAv9eas6
cHyfdlZ0XwV3tUWZmLgKmR7DJ+HrvXp3VONTp0EvRgMH40f6IWilD0UeMdqWpZn/
pxf2FBWH5X/nkVZaxT1WUb+yQkU3/K7biLCFrAnYLRH0rpcYg0oFEpkKx3OyQsQF
nQCrziv3IcHXfbTUBSYevZ8ox6A0lT9bnhoIc5Bb6Xel1/vmDaaoAvpw/OTphf2o
t/crelYuUkd15uM2GvLgzsa/6QkdV7V96/1qauxDtEw1p7qHfNzSj40EiqMHlCVq
eJGh4hbo1Bf5yV1S1w6xWjS51BINGURXQV1GAPMp1FF47fYY8JKSMPnBiUWOXazM
6cQHB0W8aQgxWT/BMYxMOtzOfEcW78J13x2B0snGedtNnpXbdV9LqjdJv66326u5
/uSQACViuIN4SyZG6xBT7ZUo1yKnFiMyX7hpgJryUrAiXq4lzm79Y5ytmrRHgD/y
NQlm99B8j0TYipI1jG9l0/lM/FRwe194IKIGh2qIBgfd8nsaxTBJbjhKmxQMyKd7
i1o309V0WLdiAJiLI+Bw1knAPElYCeWIKukONTDlF7BnlQ3QjufxuqhaUrPWtAht
DpTiRjohofG/kAqkBczqgBdZvzk4VuHKelgwzZoJt8SlmrX2GZNdiBEEnFCTgjR5
X/S1kEnk1tRf4HHGbwefMAmgWtyEUvZHKGN6OF5zfJnE61IRzJEJTfvO3ePfCokC
S7koxeOhwCG34OoNylGmtlL/pw6h59JCAXTp+qYx06W86bX5kof91YrQ3U53kyG2
vNYN1huXPauBhjlx2LDMvBACe6Du9Uc5hnfBAKeuR1hSKz5eXcTyLboXQEAJmsOh
aV5qDZpP1oT+AVtdnew+ZTV/tpYT6tC1NK7vjFoy9C48ca5lNHX7dCpyX2sl8nc+
Ss9TMQRJTL4uNFE+fYGV1ErbpmA2qBhKxmahF5NAPsh1lYnebyjqreO+UlsVJraw
u+3/WnBxBvy0H6CuZsgmGMpYdHL+/+/87wGIgiZWQjGfRyL9LvIhQXKhbhrj9KBe
ELMKYbY7qpoz86H7jT0s7/uFxN9wFKZnt516XvHnw2rM70rZZRPjHAwF4bYVGFVA
h+3POoZmILKJKRgXBjcEEt+JHJDfAno4XBJhEJ+sIk2OOIbIpFRkQQVYCqLNOtji
/ekyEA32fZ0BeVUR88ZkVHXQPv2mcj1tl6iOSzyuxQoFS71jLr1MD0DF0WBRWl3n
miOx0lDGCcInat8NSumv8+HbkF3FX2yruF3GSIxKkQf3a6c7UnaufDWiM2sXgkIL
JOQysLPMfH/ZsLlrRpiDn1ftObamgLd78Xq/+ODut1wJBuLAhzRFSA34pPjFHEGb
a0n5ChU5uHZBWo7O3xz1A003NAKhn9aCfU4w2+gkB0RzS7nrshlAH+2smKHJvguq
IJnt77nSQwXuQo/oOiCdoc3hH1PjsUc8DEOCO3fi3s3cJsNdNGXGqj/7Qm1fmyle
zgWupKJG89FfTINzuJBtGDF5ZH7FAd5e4JSbhi+bx7v2SkhzxsU9KU3JS29qGmBO
TskFBv//y/WkFrwijLTg4TIAtb0cQIW1HDHwpLwr79FDe/EvcU3d+VZ96bDQI0qv
04tAuSrJBMvaa0nf1BK4MNpUUqUeGNs/lneH8aMdHbiFRvEnVmd41UQh/aG3lSKZ
M2uTknW3T7WZx/LiclswdT/Q0tKJ8FSVF07vkt2PuJJWjXx3WAGC5z162jFD69xN
VT61rSAbWtkRsaDMrdKOBmB8FFFnUxZeNNKmc/iz50rDPgVM/V/2Fg21bonq+pNe
EBxiWM0tcVfSo7N0EiVcfPocUnv1YAe3ZGd9fQWRQhPTF5uabBiks/hromg3KE/E
xTdUWazJUdLbQrbR8ccYDUs1WoT2lU9wcvcjk++nvjtYvaPy/RMDJqrPAtlaEtGL
BiusSZENz4wSOdhFS6IrLqoK4FoWTjCenm1rEiIcSJSmw1aljS5/yWuOrw3t6vJp
EKbZD6Hx6qrkmWg0yLWhy8fd3PWMf/GD71d1xvqGh9d6XEe7id/O+BDo/5TfLEN9
yNxhH5lwFHIFVjWcFX/ZDDSOm/JofQxr4a8Lm9ZPCgZfT+gZ0iSfPzRO6VG7+NqQ
vaaZmLDaUEHgS895nOV03u3w3BIIngRjBEo45jUUQvgN7nXnaY5YDLGW/wf1g81l
l08So4B4mffgLjltNWN5hYIsZ1Aa+WUs+8/3d93v5q7tb/8ZIJ64St6YWHXDbvFK
AsmbP5UAUpO0acqCD2+UgHZTBm/nU7qNukYgtkbhmEKZnZ+4IsRToLY2MdvBtcgC
Sgty/Q0sdSSac0i3yCXxm9/6tAtYHE13Sb6D0J4TzTnhC3Iz/AYzGfxHATSMlxH2
1qLypQ4VuD0PgRSY6ftskR0N2jpH64/1mTdX+FqQCh0gO8IgItvgmir2Ca2cHlpD
5D+A34Ag6pu2Yahn1Yr0f0GAyA1ulwQvWxXDeSpuKYq/Q/1Q0lpa1ooDhSMY8owI
5/ayXRJU7CdeEj0eAYc98Ui/vST7ZHAIY9I11Hlji+UUWjILu6uu3KFBLOSntACg
v1umNugBhuceluBqv9nxVf1hQ00rrPkkB8QTAtrVYD1A6wBCiAGNCYv+/amONkDU
JqpoL9u2M5kjSuUFrb7NeNY3T2ami/4Rt+AzKS9fgT7Du9t3JLgVOhOyn7XPSAEs
D5GjCCNgqCt1myEi7zFJx0j4+VYkpvTtN/hyeQ8dZhrZEexQ9Rf0238uAp8RYqIE
3z46ezGWtDr69xKPcQEc89oqmJmveGC/ifaillQVwRuOOL3ojCOM8ChE5BwiOHvC
2brzKU3oiUcyqwfpVL3Y+cqVzwvQLWah5Ku0PAoL3IdR/zIbB/SdnACFlGyd/UCl
UUfqgQO37XdprB8U5TCuRK77nithul3El98f6T2h3kkVKt2WZmdDfX/aQ5Kr6OAP
4OVdT66nKRlSfFbA1x2uEv5+BugIWh50esZxEY8v13+/WxS5SpXwXqzF9aatj0VD
jvRHMKnEmw3FcudaPHWz3OSOcJ011wP3GRta0Pnu75mQj57+6ZRA/lc/MEbEVxPH
R8HqUKmDj22pbsAIH+YTtrnttCHtqIQH3CK7KCRM4qglDXS/4Ij34qci0qRMVDA5
TPoLYGcIJFyGuUVQGk8E6pyahKgRkbWVx7SRLtjkQABeGujowZdu0aZ76l244Mt7
7a3R3AskJHzzsSFyzoohH5ThJgNXKszhdbi2PcSxNlVz7LZktvaassATiVmAJoD8
+8EnHp+Nvcq8sS4tl8lsX2kah59hdyqpIFtxIztT9QXV5HYk9zIS7znDpOnDGKJq
mutXool1cop/larTD9lW7FLEsM4nGCEZmqpaevDQwhgcYsa8MrcAaBZa6REKpPSo
wUJiYAeTpCBoNh4Nvtk3sK1vxgMJRONwcyHZFWfHgWa5eW2UVfjti6Lk4HhSEzBP
rqnXNHhioyUv0wK/iJ3PLcaeaAZ0ldpJAKSV1pnB7URDQEnOQhSlujE6Pc5u7PL9
DrCOcrOlxGx3U5Nuh34DaudOqP5rFsGOKzOa68ytlcwiGUZAUxYcUT1hWDyiXX+l
mCKuevdW58DV2KJ7avH4+Xx0HYBLhZoCAdzZfWJcug+yilIHrFmFjgo1G8SiDlFN
clsozcVMT414/JXrJXZKu0iq+WERUuiZiLos0sXKWGZZ6xXT9k20DIY15O2nALLI
2yNBiikywdYXLTYoqbd+a532Rb3GTMrO3WrGfkCHA1X4ZmwrEJyxxBqT1chRpN9e
NiPEtt/g7+Gw26UmgSOZLu3TGSAnIiiCaV/T1hjKqNt/1Wi0j2IBOkSA+DGFGVax
m0aNOIOzddZslp3D21EkR9Bt42FjWP7149Ao4oJZWLKp1v6NtsrJS2tTza7Qxo2m
5bck6DU4rIy9lnjPVSgpFSxQ/oAI6Cs3QFWXB+7Umxe4kAJxFxXYzTDWkdnr2gDU
HlUmcgvV6BNosVWNjOpARMzT2HVJj97X55woDncHwGzHICsVo+gvdEJhM/hyLxmv
hMom3r1XmSDC14/96srkcjJV0G/zZrkaNdtF2wA1+kMXHixRb4y+yV5/RPmMGpM/
AYeNnasRVzh/GFffALV7ZZZOnnBu22T0PKv2prp+v3eXvG2cJQEQ0Atd6guBzRNf
prVg9+U0gdfK64OhfgfXTuik2UEIeM2b/EwitUkO4klOAT6elUQOyzZp3EzqOuv3
inIFTn4sjnYjjszr+m8/q61YlpqYT/KwReRpg09eIpd6JHQNaXHMu0RaUC22XCuO
9vnrpuWqFKalsePORjsXo7HCV0qM3XuI63XAgLhZy7kxPUB+82eMd+Ae+mKxCgRr
tlxAcwaUU8uWlUEcTH8z6sDkvYb3BBk9boSFbNkoeBz+hgV8ov+Mivi28VAb5hLY
OGAXxK3NZGO6i+7b4WA0Gt5vovI5xBoI1wYGOvx41WwHSGTAj2QdxU59XTNHSzCh
z2geyGLdtfk9Z4TGVytttUjZhfZBTH2767VsLmtuqXhlWDyQnDC92FA6bZUFp2KX
AgM2/AFyD0taNo+7oh6A18su/dYDwE8zzMmQr8qF/ka8nbGIidGBjp6AekkrRpnE
LNV4p+SbRNVVmeTSVsc6mw/ZZIEptUFiC6sAogGzv5EQYm11OawkRI2F9XZK7Skg
tSHSW9ywJ5BkOs4lhC4KQXy+6KEAFi6sziNUCWw2N1/eiDXV4I4ynX9eVMhi0Xi9
4EMU8vu3/mNmSxcIZjYP43ZTltMssREkS1tUwJdyby8bvdGV2326fthwlNBnKMnX
rKeDPnw0SiO1i1MIu67Gxyw5Uj8UAkataM8zoLvLkNbJu5Wov2VlqYU19IjX8Vpe
jiHJ3+HipxopMPOYnSg5t0pW78iY61EwzoGrzt3e+I/ek9FLDAviySiwt9XsD2A3
z//oB7HC0BAiwy2roZ5iU51AVhX4eLxHJ3FZ3zUMEnM1YI4j+cR4XB3HEJzSqFmX
aotfgKykMicLuJeYuLgSwQMvFo0msCiy5ajYb77alLK90dG5gOKSpTHBw8/rG2DG
V/K4EvKwILC/UW0wBn718MWmrLNdd0OwcvmUmWjnZSILuH80Yl9UIQQHg6nagxoK
pudD3nkwLFB33jfIVKNnNmkGPHWGFSqgpkUGPHNtPDxUhzFomqpskND5ZNBl2q/w
W376bg/ZUMVuAac6Bqx8uZOEy6UH8K5MXK+repTO26ZiuHqxTXy/kmYyFqZwRLAm
xwN6F2oShfR+lD1Pv65V91Cl3Fu1Kz5+izJPACUPDt1sfWD7kCc/CBTp1+O/w408
vobnA5djdDyOjMl/qYfcDbURTP/H0IrKAHCXGQue3oTYFxa2C+Uu6LPlEdIExmT6
tfPVbelJHb4PdrVCso7A96eG4XHx6se5adkfrwRQ6imqMk7YOrdGeoJvzPDvM4dL
LtxpkPkmYzq/UYA4Qgpvzj9wHHBfwsPjXiHXrYnOa7vHPYDAO9E7qzMVafwLmXGq
VQBad2EEFNk/Z27Ctdyi2lcv3cijGpFii/amQ9IrkbZtShzJVlmRFHjwPhOiuhkW
m98kyV7IQnLPpm63C7DwTQ3l/MsUpXrgyhbhG9ijbjSk117ZQHtZGTXpSijiLPEq
guNY28QQa+9vHanAdouLGVeLY1ZBfNLC/eb4WiRoHLHwxSbBsxUYPzcwEUfZ/E2m
h1nHuIPejKzYlLNT6I6mPyR1YKcu+jlTOni3g/9+xL/DMVjZDM4p+O3ZGO8ybCL2
dl8eV+9nO9agBqn3b/EePX17uaS2TWgGTDvI+q7O0S6+B3q3MRDFVQ4BoFlsgHs9
24J6rlxw7xZR2DhIemabNn3mHKAhYtpoNJNtIChL//GhvoA/CPTMQpdthmAMGzGo
wmtVwl9KbXJ/K1e2QXwonqQAXU7+QvQ7D/dwOGoKco8ZyjaC7YU/4h+UzXgYLCob
aYj/Gi4o7sJltvaawfFdkGIiVQK5N6JgDEQbd4IKagE6aAab3lEwRDKePAih66x1
fhGgBImWNO+4koZ8WRKSDC+yyr/ni+1Joah5PMXKAHWq2t1ptbArJuvGxwaBYHIb
WCogeijVLhxPGPUHlQrRjyqDpy6PniGuobLAeuIMOkWw2gQvNUeXyBw6aGdbO4Fk
f/7RGq0+rsYJLT5upQ9rxN5LgC2De87BCSDOEuRzloFV5iDoA2EBgfMxEH/RMQmA
PD2TZ2Cg5VkEprrf8n8VGNt0iiPAmMwW5qQZAX5fD7m9VAR2z6Ls+qyBJCMAF04s
OlOOBbzLr3Dv4TwSQlISaKpw1f+9pqRDBYgpDCWBVoyz7Zg3C6Y4oCd5begemc9p
9vY2OaQXGSbvcGFxVh/CHzoeUxpkzI/2PRMOsAcw4vNA5dqpbkfZTtRkwMYdouHg
gOQFn7+6iHB7G1L6qkOaC5F96zx47dC4ksW/bpql4jHFYOB4Q4VK4rIA1wI52ufv
Iofu8oVam2BGTdXbhBp8Rzk2ROHHLOZev8Z4skOt3YUyU1vnCz7Wl/TCn+vvUvoS
9gwoJqiGX53taQ0Yz/qq/PrSAw62wM13ruqTaguSz+oC9goWWxZ8SVLtClzHkTqq
YuI+9HomThGth42fYs+5ixdUzPElqit1MZv/CF4aPiCClN7cmrEM5ikWuyjHmajA
MJuFbvrHztPX22+x/+Vi2r41yZ9SuxxZEqXmtwLRgCf9HyiqhE/0VOd1dSXtf/Cc
dVpjdIaQUteFfUizeFz4hEls5ubPyL31/bQkqpGiOrTGbVmz1tSS0kbihYzi2dQi
cu1NcErt4t8sOFliLVtBzY6kzs2S2qc7n2KDanzdXYZ55wWmztb5loNjt0D3+QHQ
p6QT8OEX45aLa3fbnrntUJWC3d5WaroJCz0v3sPFREKn++r0/SYlHLglerecv6ww
QeYGAoaqUp2xk1Ojs0n7FuopkkzqJKcSmEg/XdaDZWuk/ospDKPoucQM+tYNlrOu
zERdETb84XWENN343zV0WotYSTUEsEuTK+cZM72a0n/W08slTFHKR8kiWpx7Elz5
rA1WVYVX1THZ63VUeojW2GPivbn+So45LPw8LLv9SA9tJDACHB046/eVfkztKQc1
qQgRwuemVS6NODbKI4LYC7wfow4JpL/3aPrLaDgpwCTq8QTL2+p91k6niIVCmOMV
aEYvgaU2tUv5rJF2blVsjVGUmEW5Pe5j2/y/IOYOpQznCrGbI801umOVyk80OCwu
aRz/2vk7tNZY5KkSbVVrU8cn6jnuyHlrTPG2lNXjjF1oX4y/lhCwGMV2URtUCy1H
A3jboK33MgggohRW6cI79BNrlVlYCRUzNTo2XBzvOIM0UdoXjRxlrs448zxQHYfx
akeiZevmR7TRmmGGJjAXlTAxV8YKH7RqlEWh/XDo8uaG4OFQuIsbpXGn5kJe2yd3
wq7oAGSp5e91sbAHkQRWRrrGoksZj0w4gKx+BxvXrAFDNRtapP+CwFB1+qUrq6Cj
1dxVMglMjX79Vj9AC0c7ErU/ifw8WtvpeeyGCJgTm1NmumrkQX/ffOPYoNtV1Xcz
on0RfRdK2YoqNEUrNDpJnVpu0w9k/3nRRaiiImBgAHe8fryqpeP74ndlY5ofBCYg
d7bX+GpCzUAm7Mps2HNavOu8hxZUCTxjvLdRvtQAzjpWXWA6kS9PHeRA4+7QTKZq
FXoUo8Z/oayN1AYDyLWf+cTUdZPn+1ezEUnUMj6+KMO1CUAIj29TctoufTsvR6/D
NRQxGv66QD6EA0fxEo5WP5Nbmw1J//6wyMYBFhrUz3kubfETKCqvQzw12pg1amp/
f6N9jpwS8Ex0LGPSLGEaVHbc6U0Q08xRBjHXchqJPbSzHbO34JDbtD4Ad7AkYNrr
AFGBwgdjJ/KBJtHqrnD7hTSqdeq5m5I88vFu8m2oA/dwkb2XssiECljuLS8+tIro
yrat3zAfuKjovvrfradgMdmVxQ8t0UL0KiD9jF3qlsm1IIayBdYjiqlc8ZpnMVIG
19k6Q1+Zb3DHrx98BM/FtYx9MEErJXBYIvn7QgqR93m9hViV15BhZ62GxXphdL5e
NmYhIUzKYD1TT4GwtjKb5pwJ2JwskUaNQqiYO6uGkfxTSsk5sYchV6ctSYvPVnbM
tjN3It62gPG+RePbkmkse8Xhr9gRQsAYWBOI/zaVG7oeDD9asQD4dWrrxR0f30QH
xwkn+/ECGxouUFwhEU/z6MfgeBwZZFi+xvBMF7XMlfkU7E7pl9hvWRCCdf3r4ya4
g4JX0FAv01Ym9dfJVQT68BZlgq3OIZTXtzw8RsmI68qKC09J8t9mldBa6opoP9Ek
oUjCBUztPA17TbGMY2qqygfKHu9VOhy3REeZDnhfwtAZgiU/UMTgB2hFmaiQYzKI
38VI5Dl/hqHIySFhilNfihtRYOXA3rSA64384WNAkMIJCJ9XI4lUHzo5ZcZWycPi
NgL2F4t/o4HCfBD9ZfkBSPj1SuHeQp8MWA0qJs9l1qd7+raMJmJVBv0gBiMwnLsX
YbTDDQBkMIfJ3Q4M8mhSHsF9evK/kRCVihAt64nRR6uprIRMB8TWROGLt8eHVla8
IeAzRXF1oThDesaLUT8l4ccDs0rJV02KvEurK5C3Dbke1pTGNfNmYYBa19ha1pQ6
YTXtCJz0vpU708eLOs+RYiM8ZzUXtzHqUrj9S5JJslYYwoLcqxDMgdp/Bib3qRvS
JvVfkbk+8d9/qBH0ATOzrUn4xYsjhVWp3SR2LR7KtZLU5SVT21Kefiid2lKq8bnE
FUt5SzzzsVMC3OSEhn0Lp9xhQgrq8uO8jKHuBHc+fIGzY/ujM62bzqwfjhaffRC6
oXoR0onFh6yMmrAKJSsGXf6+aY7oppkkILrSTj23J3t/UtmoSCz3IYGaKrawlxxs
baTBwFTKm9LKxlJokiuo6MmwaDktBBDqBgRV5+OvRIbstQSsd1jKZ2xnWa+Wwb47
uu7359R75X6Q4rr7d+BoFHK6x7uw0jHIeYt/t1JWPFAGNg8IS814A6RAflNypjvK
5uHvVBZlIUS3uDSGdI6OxuDOGwmK2wcCYiclxSjpFEoLcwARezlj41YXRZhhJl2g
XDMasObVklScCr6xeeG709WHMFsLiFHOjKlMXxRFfLx4K/E8nDVxlNdD3RfIY4Ee
KePLDkJZZzivijYb7c9c034YRFevjJCKcsO0YMFH3nJCATn9ZyB9pbjRZ+zrn3hB
5UMRzGNJpxq6Xdvtu1Mp91as/TKh3bkbMoBO8V2tMa2+3HQj9pjn9I/SbGSX6iPq
ML/q4rSkg2s0JURnRvu1q5vQwmRdmGXa1DMahcr+/6v6m4nChmQUC2KNbxgg9+PQ
sIshQtAqPkcgKjyK5ynar/LVbecyuA6grB3XQ9PSTH9zxkkNnN7xWU1F3E7KJIEg
xqFT867hX6TmLlUCVrbd0gSZCV7D1QGBj4cLlKB+D+lMBbKSYznbJc13kXE5saAT
s7/Z41SO4gIyXpwq5BC5vv0JdP8+bMrSHYqtbdbl7KthU674hMIhN3YwLB51OgFA
zS8h+v+ZIzo+v/6W9raGm4rh8c65dDLcyK9sddnGyNv2LmF8AMq9OQfAiAFKvehn
FSh6umTEhnHbvEIsG1v6gHXaOpASXQT5d+FtKJcxBuL+/LdIFOPxdUJaiAcNgcN3
RjshpaTcClpr3nOfuDxpkbpLhSXAz3dVfqShmP6swNVcmGs0AKngXEqfe6ecm+Yi
x5MmX7+/RwVy/TjgijZkp+rPQ6q9N6sxrna0wts9dK+QciD9/WubzkrVh0TeD1nV
dwR43mtw1aEoRBx1gyIfAl7824HnWSG9dGPLD+oRUrcWqOuf0uhJv9PJP5F1de31
LW1B/73ttUjKmbpGvVVRej/MNjdxtXf1E2D0Dhwy6ZKJirHA7iphsejhK7VKKAIe
GZOvCXS1KZKRqcIKa+jhgklNxe2y8pjwpfPSwtbys63pgSpLtDPi/RPlMP8s+efJ
zXrr3To+Tjeygs3oHZltE0rs48VKqReb69vwpZAi80bTT55IJjgnlwUc0kMoQEk1
+aOx6Uz2LppyA4ZfAUu0joVcE5XfXZH3+DyWW7mCRragibh40nWrHndDWa8BJ+By
PIq9RQULNBic6NRipxAh7rBsLpBbX9S6PFbP5xqGbq2RpuCKvLSBovFaIF6ZtpSi
AnR2AxKFfD6hRgHQPH+Wt1zZ3Ce/zH6o7g107fmJ0CM/pabL8EkO16LD4RTi4uL9
dXhBrUZeBk44m3wdA89+XedFjT9gUfzMIapYKjqJ/gc5lRzL19bqYavCtCshAZ1P
9hnbVl8/2OcuFi01owisBnUyL7MqGHuVm2TyBnh5q3VJ6W4wjfFGb9EIiHwcWbmA
gcWSWwk/qzbbpKQzLTmmpybe6Aool3KnL7W1dg7y/bVCfZ2dmlwJJXyy6tO5oNK9
srCSE5BEElasw3RCoL0ORcRspLu0c6OXGGj3E6CyB5ld1MK3wjm5h96L+SpUHmv6
UBkZneuebx9I3zrB6fLzQM/TCpU68N8np4ypOVZb33nrh8/RhSm2UhQHGgdBjTuJ
sex77Pkn53UZuQLYqk69mxR9UvkgPS9Pcdcf/coDLxz6ddBPpPm/zcIdedcdyWSY
nbofiJRe7x64ShlDZmKhylxddObuFKCDNVUWVRBGEUojk5YFbXAHhGWNH7HlqCKa
Ucp73g4fZyHozXEV8pU/sgsk0SrKGcwW7XIvZJY/ebTWdZQ50yiTdo/jdkcDrAM2
SgBLBe+jMaMQQI6cj54CkRxmvyf1hWx9SJu+AsDYhtTsKZx7tgo3vcpEkOiRZ8yE
BjKxJAwMHn/npFrozHt0CA7+cNvwaNP7k2qgFH7Sm/9V7vnGM2ALjdbCX5HQRY6l
CGwwqDNT6nJS4wn4La1W8Xo+UsFgtDFOXDmNm4zx6hOXKwTaPW3jZtQ9oWmOpOY1
uI15m9hPe0PeoCmUZTvR2eVKyK7yNQip/CwFLXET1QyWCJL8KS2QDTXaHKwzsJCT
u3MwXv6vVLvWxViNq1KWhKNe7PynSKmdFnZRGV7h7NS0FaEbSY53uj2N1U8hYQnd
f5+HGzWgkBASGKSENS/PnjjsHuj/7k3QXc5q/rQIQZt0E0F3tJnWkNnyLORglK36
VeS98dIRZbMkRrZ8/4bYiN/HXnNIJhXLjaE9AdjmXMyqftzhPq6OC+a5RhSyHp+G
XrH3iCYVLvScTeHofnvUZgya8vM1XrbRWToXSO+Y4gWJoLhnQ5ji72jK4RvLsD34
qKcntPX1/mUo+0BGWPoWEgfh1yzWHcB6jRebbkp7d8jokihS6+OS/suR3zi1j0ZW
CxrBr4+mA8qJPhnV9GAxlr4q6GfdiPIWJ6rJlMZ3RyY4lWiMCe644oh1p+unCZJy
QaQUeaHuh+/rRTEf8VhGTS1zOs9Wa7xGzkjGt5GOASgIL1s1QQ0UTdZfGmOvoDTw
c/UD/shjNlNMgPDYkdhzoFSTvEn0uInv5M7Pd/xj6p4Ms+Fk0PYmNdsq/eMHhPAf
qJ14jLWsrN1pl2oreQJFvjGrIf0pgv+DeGGF7Qs2vmcTkVSTdu/nFBeVfcp8j4ZA
2nEXiwSEhVQAKXSJQWytvwIyoMkQtdzo9QV/BVvvfLeZGVywdftCrAd/i9q870Mc
2xm52SQNfI7s3dTNAMVkzqtg22a/PEd/lfOQ/iEH48ApJaltKGxzRMkqPbBvLsgC
H9n7czlcftGc212dP2jII7EZiRi4Grt6ookIaVBf5DSrqes9hRzDEqnaAxoltATK
QGWOqntrmHxvvs9ctv7XvOJIM/hRhT3m0TDMgub6tPzw2d0/z6wsHQl+2bX3ad+m
KCL57cnwxtRc2hCLWoF4OQIesPSaoDnplBFliN/t4Zqumu7/rdcrQsXeuTCfrUgW
e7cqXt+1/MSp6BJDa8q/102BK7T629NAx+0QMbiGuO2qOC4Woz7SL/tape7tkHDs
nRR6t2Rqciljnp3Cd6ZvLvvID/+bhOutugsjQtp7Ba+TTAy3m/emWSCR4nYIXPVl
9u++9U/5B4LGGOz2Ku1J6QyvOhhMpMuNkKye0pagNRRW5ypzzc9FlXqopegPMWrY
UknohUawkHGFy8VetVAEBh7AyBHUWoHvdnjbmMdkhf6MLjzg2zJLVoMPx8F1jxRb
OR5jkg8IIggfWtnGZPGbKBBR0CviJ+PNIItBooI0JOibjfK2XbJze9x5xsL1396j
YLJZu7b/jHY7V+DHV4AmLcWSrYzcXIb9VVl3tPbHbjJcFz4Wll4KBsrkCSCSeljm
UwRNB3bTIMfiK21pbCtsZ+l1yHxzJpRB56nsHFepvfljjmwheEqM38ijxMLwv0An
Y2qJSaa36NnfwOCFLd7Gd5EtI28ID3iPvA5+9eeNNLaVc2Vji2XlGUhW+lb01CSG
7Yt5SJth9bEUl5M3iNoh2AVM9LRGVn+bVu7CHC8BjvuhlI4qQv88C6WAu4G39gZQ
VsOscTcn3dtfZDDH0VR24nbtPLk6QQzJbOYiKyZ5sqnyzA9ZK5ONzts1uovIU3WW
+rZUYo12QwU3gK5zhMZL0aD+Xw2gsr5w4fytpOZhGaF3dt4sfKw/lnkNGd2nli61
8Fmeuqq/KXZI1o0HRhex3vtRlnlZqKhsgKWZUmazcJmAQxM6+xx8U1DpVGAn/AZn
tooFs/VyReLVDYabFya3neQ4KyuHriZ3l//8XRkpWVBR8AcJmQdu5RoC+F/+jAlD
4jib1VjfHrnIzyQ9bUNWatnmHnU35tg4LkBavuihc57h2G3wgL/qNBdGegz7ybYj
++zyE2NXcoyW7a8k7pJRehYFuhwpzxpQ3ENPG6mMTWR54ZdxTsmHrhmjmRJT4j+Z
nPSRJitAzmzD7pc7sBJjuv+1rBm9FvADy41vO/H4iGkTJz0vaty8lxxVsp55xAEL
jWT/YsfxAG7ozx5QSZiw9JaKtHzQjW6OJPsj8B0ehpy1w9o/fZhksGHb8kkDp+wr
iq3uUELZB2/kKoD6lTcV1oYhu2UKPZzZhf1crbdisxTqVuO9U1nMG+OQU8PlgfJB
9ALmTc/Q07Hg6GsaSyuJVATSvgzCgaI8n1zmQF47W9A/fyYYHDMFAP7xfCHUac7V
AePhkKnAm94Zv2RI2ntuarf8U1jF0XSNh1XAt81T+1C8+0I3TUs0mFR9+6Y81K61
gwjIqZFCFBkmxhDcMNa5E3C0BSdnMYQyB2OsXqILVz3Vw1I85ALTYShkORHBQrqQ
2VAw2K4zXPMwiUNsSKkbyHpjV3KiSVm1emjKJw/IrTeY3HVfadArOYUmOy1NK0jx
mDAXOL1DdRHODzGcmMlFOTR9zHuaBdpu5FYggIi3nsJGf8PlFQrMZqr1iK3gsqzk
rVVQkxDm3+jj5B5Db04Cn9rPKJMm5q6rCsb1YAbf9jYLuUGcTTLlQxWe+YDJGZEI
FLPxglW9wST+SeP1vfQXxKUaT4UK8GcOU46Cqm3XIMgr/QBEtoaXt4oDxRazrN2l
oUkuGs+tRlnRTWP3+3fjoaf+hT52BXtM1Hn+e3WL8eyKyzmgvPoTHjNrSRrZM4Wd
xdYQjA2ov0qJDmin0TOasK9Nz6y3XhijNAMi1IR0bIkEgqSfBNCkU2GYietcUWuN
U0MEtademNbYvjCF6xVd/YEhNXjtXSh1N94q4FKliGC8P9xJIiD4oS386XQPBWRH
VaQPhGibQepSbNq0+MiBp3/sdQw6JBipwPhLfOY8KZMKxmWOL4IVFyEDAH3hZ9wK
YhtKhWkKC0rnNd9wNpgGn8EIwxk/U1Dk6KkW1vVqE2RRcSxGUETzDib6Rx7F/xXt
UHGgsLUf8ThH8MFo4+W722uV374LPdbLj1AX3SFelXi3zA9LPCZkP+hDQT9QAG58
ZfLLsQPGscEJe+sJivcB3l/lVgREID8a8zlQTElG0AdVuPkObdmihxRbktGvXKgD
zZIicybzG69uvEmG5DQq0sSrforOKhAHn5DtjdLcA09DFy3/ehhIjFAmCAi0keJU
TRjtr94EDqkn8s6qETr97GcvjDed6hQJHQ7Hf86w8d3rUsii/AdnhyM/OJ6Are6K
zrO3hcu/6+U20W7HpN/HkLg5u5cYM+N6etY0amkr1yUWkFyUi5xNSPKr38Drvn7v
3B/Oa1q4YVmMU6bv5kDw4hq1fvYLDilYwNkkGb189DsgiaA50xpfIj9WAdmSEZ6T
pZ7SUXZSVFBfcTty4Jp3FmdYnjkTwKS1C3ZETVwoxIJ4IvJHllbRPTZLP8LaAd9j
5Taee65yrsyVQM+ERfWEqS+8FQaIW3I3a9J707aWx0PgoL7seehDMaQSZ3jO7Zp4
gtATcxMsmIgDBfbx+x37/DhknZV+C07mV0YLs/WjrNgHvJnlRiEAftJafG1oSNq8
yMrIwYx1Fd0UD53uMVN8OpRFYue2bdqKcimfSNnc68AUyeke5+rlCcxGu+zYMztS
wYovwrCoAT6WItS2VXTIG/LXLn/M0u2fQfjRLbCv+hcI6yf1PDuxFXE3RYnSLrpL
BPFSvrkoY+ZnB0UQVaEz3PsLPDwCyrtwMpFWabqFm5Pqgbk0rngIoauOuEUSMQ1j
0DLB3bK1JBGvp6r/K0pfaLGmj8agq7vbDV+r0Vv40ko1earGoAnRRN7J1cw0bh9F
s1+DnCq1eZUO/nc25DHvs8h2Llb2d+679miKVQ+6X+8K4PUiXJIRVqFybQnEAkU5
f7Fb09B+XNmFswfkswDquVTqgMacSQpWnuEx1OC0CtCvHjUDTAU6ytLXl7BWGf1I
3UTNSfzf8/AnhItd33P0k9Q/QItiKiFiVzvXaKGLbW7STvq9TeaJG5V9wXKCVzpp
tyotKWRgH+QqsjYPXU5eWQ5eInuocypodLhQACSriqHAo2kUH3mFOP2zIJs+0jz+
xdRjl3Ewmcf/aiWUsBlN4UQBhjAcLncPc7dldR8+fjJiHav+LONBvzvyWRqYemE1
YP2/kn1TsyM3ypCqXHAZwUblyo1+4ohQ0ALIlTCVy5R53KhSbzi0xtQje4kSbS4V
Q4S7VjORjfhO7vFWtdPpxjVuwJPlMd9kmA7ccKibzuWBquoUYjaYfyeDJE1FgIO0
z72FfNWA+a/1sKvroB38ZjQWiWliqdPv40yCem+KGcm6ndr8MQdP8c6Tv3WjL+tr
2r7zxp9IVOsNq/A5R9P80/50M70oeksP2GIvM0NcKmu90FbwXM6/2mSF6Z+FyfU7
2xFUtxUXWGAbbQD9JW536S7UZC6KAvVfjSQRJXXRWpYq5BVm9JoQCx9DKOE032KG
1kNfgej51A0XaCqlCPfdU+nMKt3Nf7CL2/pkYjRbph1Ujfi71YWwgDix8got6gaB
extf+s56U1EQhKdq85+pevyHXKQZn87BJVEXJyh7NMVqBXYw17mLVyHiI+kJu//k
Xrn/0c3oURYTkJnYQ6U+JcKWXHTSx1rqQllt8Lr1daudppFFENQrxj/9Cubh/jXZ
2eYBgYGRRQs+eUIBjA9FPH4KL/5ZUcg7rsjtQjZn/kRtfIin8vufkyOg/dCTU6Df
BTVIz4T0g5KBcsoe0HG/4HA4+lB6lgkM0y13+w/sxHDqJ2WXTivMJ9FrxS+mC3rg
qCrrZH7tEGwW93ZmhREsTnbXvLdJosfHOe4sHApplHTdAVftNqmtdCnsemjyoslj
mfsIXSZ5yT7M5e7yjg+tZZE4XTcQ5TWYRtr4MSXTiytJlj3evFHngvuwq5OClHaC
M2X2CrZBP4mdcNS33mxsU0WYHZZ5Zk7SY0IfK5VZlHB5x3PP5dIsGE7yInXIIehW
ADScOTYgN1G98tgstNLRZ116sZsVUU8P27Wze/j6Dkz2EOQOiFDVdcKek+5KIuCx
nVajH0WpKm9G1QgR9kE+hVUJSTyG32PMXudj+8w+CnNA5XoYRYLdpMw4DY/owpI/
YUSVVVWXZl3QWJaeMTK5MIpTcCcVR6qLgKiQnWDMzl9PD78bNuv5xv8Q/6suqG2K
CpFdQwjJ84zQR/57KSwHZp4HRUmaiddGkcnMEYmoEASWFGTQNT4tHkFWboH/aqFe
qDKdYflc8xjXRbvUP9ebMy1u9RpP0GpgzFdd112r2WldDA0GbrpRXQDsFBC0zRWa
Rb54bGawNBEK9QMPWwe9pE8ojLvOFe2tT9FtwWgxRrUxx6O4of3wM5M7Yxpuaf8T
6KxOCCHLDQ4u1FC6LPzXl0f9EepIZlfUaIPI+WNZXKpGPFiTOKx5CcqAehfwIyMw
3jH7+SDhT7dLbGqbLEDI4Uhb+N23qW3d4BKqfDy9Wp/KveOFR8sEFb0Zu9JhKApr
UNykAx96nYRjhpACJ2Vf55G3h5IWkq8QHAQuNdNj6v/gET5UQjX4IjjWRTZzZ5f4
oJDQT+c+KTFrUu/9BKCypmpqZxvBxV+Tsn82uzeOk+wmyRrAVIiWTCkSSfY5Bj/Y
x2ljswL/oHhvCBuhw91dG3ucvjPvII8oQu6TBvpO6+nHo0qlb2pXfW9IYnw+PZu0
NxJ0FbkhTOmQg902ho8RNc0bQ7Wf/fUW50nWk38m72pIDAXjyRXkmlEL7UoLrtJU
WzR4vEQ1dk46OpxHcJ078xxJNa6mJBvCjOcMWsYHxh19zHSxgln2cWMGR7CpoFd1
Uq+hnuQkllpw7ibfku0xt4gwD7Jqb6lS3fDJGZvM5OH1P5wJSubdNAjFDVCCTAtd
3ILPgkEWEvrpNRR2IbhfPKVIZN9+85wvlwYHB8lscOvowRpYPgwcqsiGFnpHMmDv
3MYJsX+GRxJ73DUktLU6Iz/RtHDEYVhsIemKiutKsj8eeeNRCBbl9s03hkQDViYg
N0qrrdcX6X2I+bNmJCUYeGD6xhoxO9LlTqqmIUtcxEsmfWxb1e8oCAWMayr8F4/w
whIzH/rd6o1w0W3WRoS/5h+1ibVf0ANfhC9AFANAa8X2APPS768irCM1S8nCbpNn
XsCDUl2wnmflufSe416fT1/huIVfAS9lLix4LuysmuwmZUhJSmICJK51OBLwo6f4
sGAa3iXITxq959QZqSEFna/0TxJRgeNMbdSBDD1YMzzQUjLmZSNozwZnFsRjiIF1
SFvjQIZaFTmiRq1crk4bDWeQvZczMNI2x548W30Dliefyle99gsaqRk3ORm+R7qa
Qx5nZccnx3GD28hGD31xjGK9YxkH9eZHFJk7KTrDLLuDJRvSN60MYn0Q1H2chViL
szsYGhEfWtqmbxixVEni+eWEGLA4woU9hX5QIwuNd4fTlNOu+FKSCY/KrmWjMFF4
8X9bDI6quXj8Bjduw+vlkw+3jtfvZuzY5fwCmEyTGBzf9OGMmLaSb1YyW2FZqJvJ
J4qoFiXHlma1PTYac5YoPMxJabq/2yviCwyjduezbqDsEcxjqKpU1VLkegvjfxVI
o/vKsfe7+I1daIOSzup/DWox7+rSQcg7zM+dw5I+rraLeg9TDbxDgx4GA4m3NKvt
t5DlB0bNVM7TudSCQw6I9FXLlVKHng9OJkWtjT6Zu9zZ//3uy1jM0q3u8wYei3XE
NpsYpgfUsQavyAyK3HB5U4AFHK9NG0pVZa7xbBiBbGTYWKrMIdyAUKn1XDWBSaEO
sJxOICb0pMMXKigcfKKCeCyBw9RJheiu0M/3HIARwu54rWuyAr24trzxxXrxO5xe
0U5alZMKpO59HeH2yDneH7wlKlSKURViinp6Pma+zkGYge87wfNTnZt2ukPNiASA
+xF3IUCq4OyV6H20oekZWnba2QtaBzyPrDCSKO2vgNa2Ae9Ex/IiKqkHlWm6FFsc
YY05eYTwWZvEnoYBRKK+gLtdjR9hLqP7PN5uMXzmWXg2HHvGnnIC4bajQT1ItnLR
U68bAC28PXSWP7E1dd8cgCvDIGsXfuXciuS/NB180VA0MZHE6Mc0pB1cOcaWZvA8
SVY+on5RzsFGae03ewTrTIPHrbjAUjo8ksQNBPX6JmCK+9y8GuSp/DZB0Zqhd5v/
1I6QpXMINjw+I2aiqfWl93MZL6dfIFgjkZSf/jxkOIfJwFrtG5iHWEx+VvijUkEy
1KfQrJUU+OknJyqbFIr/NQFXAK2Td5NqO7UiC2ypXxllvGR6s683QTmMjdNdNMuf
rgEfylHoGShPJnQrqz1tUXTSDF/N8nUYAn1JRIqhL1KTmpCsqBEr8umJe8+XRidT
iXiPgpDaa988xohak0lxo4SH/TVLDx2x8tSjK4vBPqy2CHv5DOacAx76gh2eufHk
s4thDu6BKuuzHcWl55j3Pr23wSGy+f+THL6gXHlScUIlEZW6WLcYMStGLgGuXDNA
WXYFD2K2N4wwkbhffosAraOZO+NQxHMueIgpl2ozryOsyATE7LZIIEyh2biG/MVl
WSCxR/FvbeTv+5yKS8w2ZMIlAzZD0EcW2gbwh5rDMEscATn8XAvMuxdAU+OpsdV/
D7T/0fEPPZtkfNX5DzGPpAmNimZMvM6mRntfW7HVc9YBjOww62emE+0SAV7r2Y0R
cWhcgXHivtjKCmxpxygem3Sp24gt2pF7VZLWFbF3aWcx4oirwrn/yzQfKN9IXfK1
C5FCO23hXh3xNq9/DDAHD+MBdqdId0qHqNdMRY7fMVfpTlbCBG9+bEo6AKnaCalQ
qOnNcAp5JRXQNsO8GPT+4xlF7z8iRNh8mHg/FccV631kQJH5kkmf4jNMZIEyEjRL
fOIp0MEEJh6q/HwPFmWLjAbRuVnyIXKhK0I8Lnfre7um76wLJhB0QHaaKDIw41ov
DyDjcBj483QcdZ1NhRrh/TgDYqQDef3dKPZpcY2pw9Dw7TyiDi+8pV56suLs7fZ9
hWi6cA4+CubeRAIb/3I7SqXt72MPo/qD2uMSRBdUDpaA3xdzRMABmlBd+uWckU7h
OeVtluAP9H4770rWApQdGhEFkI5I22w0kczJKtR8b+cMKQL3JU25JYUPHpy4cAj4
TS1KBp7Mu/bM3I/3WyrydAG5JYSWfcri8zjp77AgOe4BlLcCEk7tIJyFOxcRzDRw
XJzXlU8sIU2erj4NzHSa2+5G7FR1E7txSA1/Hg//8OwU1tlhzJ+S1UZ8qxQUp0l2
SyV7DamSYLKj+O/WRTw2XPX8ZHrejgvJHnOAZFOdhgjxlzn1VIpnSX4rTmT8yCXw
ajbPWgVlMus1qqpZdWmzeIyB2a1FWkTZh0chhxvOtM3wuLzXLcOANQUdYTzVjurR
WXHTbwaPSdpSwBpdqJFeK8089bGiNia65OEFiFaA2kFkjGKxccDMR2TgQ+KnGlbc
PBao6T8IecSlpsACTp6wF+wmlLhxbgOVTSv/b3njU1dgNpV+uBhsalkhn2JfKYVO
n1qKQUN/q2yF8xCwk3YCA8ivYW+1i2QWEFvzmHxmW8X7Gx4LRNOY4G1GSPVDki0M
1AO6WvFIOu+6+p/h6f7IAC4HT1NgsQG/Rh/vLQp3k1L0pJKmtz1AFlcsVKr344LX
IZF/rB1RPn9g0Ft4yG/P4o2g1PNAhdiJQTpg14Zv+8Qt7w8RREnaKPlRHIBmXpTG
189Jp4b/R3BRDuRggnLB5NBAdBwpzpKUVPfAgOmxi6kujtiBjlmMEZCJoH6c05Rn
NV8f0imBLR5oQIPAd78hZTyUS0gVn+LThnnoH6MeUTSx7JIUcFThSAXNo2VhN6Sj
GT3o+OFAG/az1z4GW7cVYuxZmcvIDzok/wMgya2O+lNuWGks/YqHqOVPmO2ItPDN
9EtK7/+IUduLOyuiM7tyX/5wnNnImTwGuuw0dO+zVSisFSD5URI+USjhRidZRCSb
UqshNTmhWqmI4zNVZ31wA/XGYaAyGI7ckruoR2Y0GqsIS9v4JLjhx9oJf5hkGyDY
2FfFybrqgf5FW+Ii2RFz3zri8Qqv0qKvZ1p93uk+Qaxz1PLVbS1tlUh2gxiH6u4O
OmKDXfMeU1T9HZgGG2qAGQb4eMNpRRGXCarfcMbokp6GdsyWorNa+Tddr41AW6Vt
xSRuo05fBHJ8KJMNlbdoqdxbcqtnvRghUxWJQDgNDPytl2nGBILjYhs+OtU22BUu
JBN+n5Mvo2Kc0BjkTm36OIE0XtmXSI7MdydCCMj/R5OWVc75U0gM2TLoFEhSedRL
gTlJltT8nM2f5VqEhDyArONbjVpCxwwUUfK6VF8glGeQZvweWbnD8RqGhjYBfSr2
1PD5kQeMb99Rk9GT8iOjuwyKMkvS+UWL/50N5DdWuyome0mbD1ZY7sMQc1VcKxw2
aOcNQDTfzzRN+uelyMvDR7sbwXJRShnJ7wdpdeKdK6wdELDcIgUElqjvuVOT3xZc
8TuTnzNF8yJuymN/gAWNKq3Em8tLOfDCXTWzB03aw6GDCg06tDm/cUbavPFOYj0z
O2a4wbqNoRQNEGlwY+UVpic7dspkHJHnks6bphaMVHcopftvDnZwNnOddY2qz9MG
W0xenoYP4okayJSlbZFDd1bgWbWWEQlzuCdJtq6rbQeLN8MCAlL4Ks9Cmu6Tm2Sw
EzyyTaViz9vlOiqbajqmmWJQZipWEinFhbdguM593CGpWWK0UKJKXsuSNWKReWBy
rC2+xCtNTzmt4Ksok+AoFRCiXVKuF9kgDgpbH3LYgffo5ZxMaH/k+FPMcob0YQBe
/aGIgIoFcapRLvpFzoEsi19QjftN90j99/8jglQwTIOm97d6rc6LtFu97YqVVgIs
0jb2qyMTeTUiIr0/sVtBDco8aG/xYSVn0TXJinZMSOFH7ScwAbITpbm9AaGJ1Kcb
ID9sq15c1k6yBGniRIQyKJkFZgsLX08cqWZ8gWxVIcYThyFqdx1EUfCo2X5xzC89
66SU1/HfvXlvF73QGiGmNE0MwPP01Cx03hDF38BAwzrVX+VvcrHV2SNDxO6xWtmY
oM2nlLILzbhVxiLuzElM1UOWEFxRTmwSDznU+CFNvJI2HOhtBv0GTDWDBY79XXvT
wHd882VmeJxBQP1X1cSgp/uLKNSz95g/8Ib969knOoDdRozKe4hid8ExcTXSSR20
AOnIAfDQieewPOuSSWFapPjHguLtKA7vN8/yyEPZPd/g2ilzeTqkCPbT3spoZLSx
FmzjcIqMeTUEXLs+WTSRg01D5PUjLlgNu4bUYuOBRVN04NBI/mmcmhAcP2aAjNnj
+CXQSV7WPd3+hUvMa6mu55UWW9ZS8rOvdqJwy+Cbm5bqN3IpR2ZJMy0fnSOwQ9Zc
6+XI/zoK++ZviZFlPkkQ3Ug+ou0SeCzQyk7uN4BinmCmIVmjpGhZNZrTDAcLhzki
MJeA7u0Jmx2RekYZu6exVt7k5bG/yZv5a5f8LOymE8o7m6QVzIATVASC8gxyrK/S
sH9JNWpSaAUhjE9wpMhZ/9X4a5FvTjujGMzPv2361vLLdWSelMmi11qlmIPheCQR
7ycnxBY6t6cj2L0ow+7IgfZ0fvzfPyjVWbhM2U04SusHJPjB/Fe7MuMA1jM4q1At
kQyCqO5rSk2mL7hwf8bUQkoLRqKtVKUYsUGBywQ96HnkUfRMRVMDk6rVpBmNGc9a
FFS/X4EuHBdb7HNciVvMhHFd7JeZSh6lNP5y3Uq7ewXx1CaziusJzOC8GWJW/+kL
V4RgWPCgLYMM1ee61UA0Kh0OQzdWY9xk4Jt64V8i+hp4Yyg4LSPM+WOFuqivQGEv
u+di/YnukILJo5878DQPiMDO00SHdIMyDfnWIR1q2y42Zwx+B1jFcwSRbL9n84B5
QFdVgSWWfJVAUlxECrpuyg+4c/ALSqRZS+36AXJnUNmiv6DkCvTqOKzP87zmcQNA
F8eO47cV3dAiR/gZFPvTANg3j10TvWnbeT8URPk2LQ0uc7uFaPJVeUlEPFUfSqpS
AHQogX+fe4HRg7PH/vSwMmdJo/4Eow1ZFll/A9O+1ysnhW910lkh454dUha2ezIX
ehL8aJagL/uq5J9q7UIpSQJOwLdw2Fcohfn+29sF9oBF5aNZ/5CdW4edIUUWmcYj
rTx2qJdtYapP7LGzSSCF8tsGuZ+SHP3zE9RHkH7cw6ewEc99Be1jyF4joWqiypcY
15srCoXs4qnJ/8sKL9NVAfVMVU2vagK0VqN0sn9Y9dyOOyT01zmSyHwA16lCwn88
MmhO13GgLkeVuNsLOG9JNrr5rTpzZUxWdPqU4ERupN6/J388JEStFlRvPhMbBHve
GZz/M1ihCaGHIxxv1Bkbth4g8DTdrIebOiwqNKnivw4kUFX4Q69RgMLFTzywzLrJ
LDPvG38VqxlObmgQwtDF2bFpG6cZtpUKKheX/yTQbxGNxYR+LhzIXptkm6L8k1zo
cE9MmZ62nYrcgOUlnSzXtu/1BaOlNsiuzMUoKLgy/PeeSvChc2bYBKCOxi/5+ydX
tOLUGgQlBGnhyYWmHLfFi51ClhvSXJmTXix9c7RvgpuKlwomFjpta9bBkb3ekwpk
fN8deAbsJ3mPF6aS0nHkk9CvW54wnOcSY7MtOdA8W1gGxcYLXS9AeV0x1P81t+gm
K22BcyfHHhKGyrDzLTfov1NtG4qVdN5sBZq3Pjll5iIYlapV7KRaiXBtZZ+5vC6y
VG0xT9fvdtAzV/xLfYvpJpj8QQhGGwiIdveYM77N5+iZwdUSG5R7a44D0vRmWV4U
Z0/KLLcttqJxauJChnr8o4C7b7Zf92nfBdjxSPkg+h/4erZT5Oq10N8dAIB6HgpV
uAGEzIPZwpA+yHLPP7TyBNgeAIUbscY+f8cWC8z8mED8xrrA2pR+PLHqlC93dQiA
TktrTKxuMvJziWdoDb+KsaqyN0HqAX4noHH1O/ZqJmwh2R32XE3BpyyafvbB6/JW
9jyBdMo+Gj1ZoLG6MqFia13aBvl2Qk2ToEfRZScJgssjnw4VcEXWGhHNnt/rto9o
Mb2yzb2prOVCUqjfftliM72zN647P0lp4wzyFbR6FM41QK3huCakjYALcMSrP2ph
C2PrytoRok5RSgFlMJ/T/oNXhjqML1T2P9qiXYwZgaVz8Wxkts2WjMS8BMnkPPN1
2QtDbTrWAD0fnAX0J9cs8xD0FWw/KsiUtIfBU1Bf3MokFQwawb6Ovi+jR3HtX/f/
eFcy5nlTU/lYZdgS5me4kywwJtRP57S4vkS69G1e3CbgL2IdFT1H9ZDxrG35zzPY
5L4Goful/5hCewvD4eTfDZ9HP2yUZhs1k+fHyXcmkeuFvy8QubNiNCj9U4dJLJwN
R3m+wwOm4EOUww4Foyfz9zztNfIAWZfyvKmH50rHrBfuaCXI80wukLJVbQKnsuP2
vbP/ajCqrMWv0gsAry64JTHM/qGkjG67co80xB9h9Jx2qyk3j3PSIi3mg9bxuLi9
3ztQ3ewfruNNFYG09/a8kVyrcxqqL1LEW9LqI14H5NXImARWuMxW/pwDZ8ImHncR
+xEO/lcWSP73JdH6ChuXHh+TPr3RXhDnHXaXIdMm2UKMOHzvsfLcs3XoWD+F05lS
1DlDEHKjeht1cN1lYKXzm4muuu8TJnTgYTbdBbisrzAaoSlLYGgw43/CmW+sDb1X
DLED8IWQ9W2DsgukXgEde0sv0Rb3cHs2b58zoRjCxQTBrFKHGIGW3QeWdPHVjJSH
lzjrGTQh3twRw+jbTSZPYnk2tKrOMJZbB8CSX8TlRFoxnU5cVTvqhQMcDZDlshL4
X0pFqBgci36f/lArq6ZAPsmht8/xO2hJaBQ0XVfh3Ro2lGvxY2V7Fa6Z9oROmf58
KxLpQPpbz6ehfvwsQYO6nCr+9aQomt4WzQ0u8TP1FGY3U25z+1MjxA8zJXrhfK+1
frjrxNc7k4CXhYde5MZirVrja+Gf6bdAz1YuSfv2JzHj290UkKKDx4rVjJpndiSI
GMae5a+4i3Dk/NQV+DdMQZMW7eMbS5bVE54MOuhK2YH5Dhc/KtboxSV0oPRP9u/W
Js1+tGrEHa2oNcR0Tlo03h45x7NigLI9n8DNBKpcUa8KFOAIs2ObDFaV5snip0/N
glG4Sc7ZMr9k1KV9BPHAuQlUFf7URHPlltx3K9OHYnLWasFrKwFo2I0pnHqtYWEt
+yoL+gdDs9MucZCnAkh7vlF0r4Kje8nVHh4bxW0ibc2Mzfz+uzXU1qRGYPLp6zvt
Xw2t1VrYGefE+7dVix55VkFdSQmlRXg8ls1yif0+nSJa2vm+wsTaFU1ZSbUVk9em
zYpyVE8xLJCMg3jnlydQpMknMK5DlmqXOJ5tbtp21HIIGtbsZvhjIvtJD22o+1bp
QaPypEs8WIJOg33GTimy95uk72Ghg6HNEVJKC5IeKBhgwKFq/w4Flvfdj+gj1vfF
nQWPVPqfnkEzhqE0sjzEc41m7MMTmkGWMrxDDcMIPabpwPCSBUxSH5HBLR6LhDNZ
TPdb1LWYlwoD0ft/DOJh0nCPVnHTygfvIUSsxmAM5BHB5iJdBLkqKL+9N7NDdgwi
Kj0U88imEoVoWkshiFADXpMzps45Ev9YK9oI2Z2oFnFwkqiqOtCdwzCrMc5zIQ5c
g0Pg7RcpILtxxODqbtgTFzp422t9krOZhDix7o4sDo5d+2FPSN1QSoNND1DEBHdv
w5PO0H2W0u5q1XOQiLUjW2VTFnSMbhnxlzsBgkeQE1mLtpNuzwkBCFWKQUzW9ubJ
uDgrmDeVD8oICwmESI4NGjgMVC0UWOlK52Vs2ohBYY5HyaHsOSKsVwpWtlH5dkPv
pfcyQ25Qw5U89VgLFnJHsp49jojFRBfR1u0b4C4fY24fnnCeCoSKAlzTEhVLUaoK
Fl5WzSHEDCqMrNGChipCJ7xjhTlPpPWuJavv4WpUqhgKotxtyLhqV4LUnxWzUdw/
h2n2uoPjvuTGTjApRY/iyJykfcRLrNhLbozx6a1gOEQ4tipUDlYpuAZT7b5086Dw
XUAZf73uu963B4ERZ1fV0PE8lUSDCvQnvRL3+Wy3nI4+fZsQzzxZEkljNx9ZBIh4
TYIY1IHi3mks575ZX853MxuIY6vKQhjcjkbfgf+7NQd802TWH0GQ3TNza9Ef4GQC
9e26KQ6VQwufOshBk5oM7N4vf6puWr9RYDRcA4nbkh3mCRvbZd15EemkDFGvvMrc
XOLFc+Rvl3HGxDN44sRvQ11CuDyHOjM5e867PUpr7Us3Cmoip4XbEwaqfc8ss26T
ndqBQX1cqUksTNoCzEcrqoV6J7OtVtkyLR2Sp4cPsK/DCINt3BhIQrEZfQSeOlkg
PVAwRhiNkWU5GtgbUM6evVD4xsxgDFVVda47bS783qTMx/wbXg35h1BwGybW5e06
SYelbaoJAma/iu8NnYmDjp7OWvTYhmwhWyzqQ3Sp68Ik4Wt4L1Onw13UxjbDJd2i
pxaKYQRV10PuJGCrOmMxoTdBfWwngHFUiJbdgK+lKhdVupE9knuHj61yhageQ6yd
bg4OW42q986oB1eCHrni9VSwMWhdYLem/4gpgT63dv3NubpQ6gVEC9K3eeK0uMTD
Yojk7XEeKxDD/P3/gyK0FqcMm3ECDzkzGZUzbMdkYygazBQAW32szHIPliDSJhQe
0qYZMfCGX345FWgW0jghkw06ecxRMDBlWIrurRuEKuG/yjjHGvpkmRSYTPHwpIOC
PXiUZjRya2MBTUrk7MysNs7WukdbURvZqgc3TT3vApg61Q1yzfARvxos5DhNyieo
0L858EatXXeZScD5qdR4DmcMk/88JLSPZxF2sedutJayTNw/qzqQ11tTDYwDF5n5
aL/DVqO1So/LbR+GLLUorCcN763cNCO3htaBkEzlKrTmRhYfJsJBUX+N2fgSfDLs
svZe8L4A8SFhPulPGiJ6tX1sywhx/AvL3Q/sbNOjQnUscAw7EXG3RRrPiNqcruDo
fqBQuhMW9KeaHHK7t25RAsMJp/tkBEfhaC5ZqKcvuCscc6V8CnlxGkqoXnvaHkx0
0JXfHSV227E90zL12TQ9YWDVCR4m1ugy6sYbov37yA05wpyJlP7ReHxqPNI4IIcY
VCU5mIsfTRrL59+e+kLJLYo4tMfUrd79Wr2/92wec1f9pXuekX3sEJAyXfSRg8ch
kE/2D7vFPV7yUbXEHDe8rsBAkmk9o75yWJLNerrIKhrZQ6ffvyWrtksqRMAlGHXu
pRhhbj9JNuJ6jno2umvX8+UwoA5bVWoA38XE5ysdr/l/GBtyru3dTUCmKUD02dBZ
Pry5/c3i4oEdbuV2bUN+LuGEO57onUsQ1yJRhpIcK+lrZj+mOJwDhDT1n8bAQAss
Aq67pxnGJ1DeOpnOLZw7pEawVfC891xcdcBB5BdHsQZcyPp2yqxMegsSJ9X6ygOW
1OD8WVuJAeCyaJGFbijzPlHLQLrV2gTkU/wSiNUDRShat6QNnqwuSgnwhUrMYd1C
Ezc673a4W0g7VBkA8dsDesS5OHtA4WY6mJics2JVBM8hv7/omNKBrDqwrxevshp5
3uQjf5WVn6+lKS0HHwG768ywLDDs7UfEBVjLqKqKWYI5u/4j5CSV9FMgxuRq1zvO
oPRErx/cbrNKSJFfTJHHq2FZIWXQm1LzIlun1eJFnTAlyUssGLNDm2KLU83tkqOO
+MzPF26hboAJ9ZeRUp0G01/9XVYIiYEtruiLgdlvxAsyah2Ub3U4bk1zp9BFaHm/
dW0+32I75hCI9N3W2DHYRtHp7e1cEFa5mcC4/S5he6h/VqlRnexlSgfXnXQ4DYtR
CADVzw5PTx+0as6VBC5O0QUHOoZaX3sUKv40mAWfX+koKlOVjwU1bQqdzOEJg0UM
2BXLyjiVeMEZAKvq5DLCiH+Xnhq8l6oJcDuPhOK5WEsc8g3kI6b93FgCzvcH/fYs
s2tPCQuqtALz7iJpQ3OaGCSuxnKaqWC++N1+KX7sSzEkB4LJjbEtzgzJy3Ija3hd
OPUrgUB1sKQgVcpQmxTuxrQcpR3PclMp5Imj+43WHOymFIjLUi+yFVVk8D7t7yip
O8qfZ28HZSrfoqMNXGjpRYfpo+CBGJyQ7qrVesurf+1JOre8SzGzM/QFsGcoAIyD
GYPAXqfyIUARkbdbjfm4WCsWK7U/1dnBvGPUMZW/cuLDFRcL0F9Ss5VFD1K7/W20
wU0dp4nfPv/DrFpWemO+NiYq5g6903X+8/DAmE3FkOZvY66ikAfXUkLah9D2Ikl3
KaVC4eW45N/do2Y1j8S0FGu9Hz1xs5z0k4XiNB3eRFhkqy8vD0RczesoViCUsrQr
BxDLqE86FBHo+RIbzneFvB1mEPbJotJM6h5AOp3RNMgGYQJFgf3YIWlikDcZH2ah
JFsiCkoKpGltEcjN66Z9Oep4iXUw8xkF4nl+M8YG8XQSAiqy922w/cKQep5DKA1j
/8YwSIIM5SjG6BxCbU/ofUQKgmr+TQL5f+8znamqdigyKxmOYmNqN0rwb/oTnPHR
lk0lZgwwE9OZ/On6U5RpARziBr/e5NOY2tWzoKJYKw2CnZnUjcKd+1nQ6H9dexMX
PzxZEUUFcPUvfBIyN2+vd8qd/8723N6NUW/xAaIyFg1XfBq/6s2eU0rL3vmHeban
DwRjfrBli1aNIRCNqqPkZbIG8LOAmd3ofd7LgGe4e3snGWFN8WNt2ITkhe1YxZZ/
mEQ4jcPXzIiVKSG9yHhTNdAFxyPpsNtVSYeKwnjqQEJ98NwGKegmU3nkSlsA4+26
yohh6Xmr8e75ZxDOJWPO6C9g14p1lz4d4cbewJTiRmIOwAl7Dg/NngHlCKSaZDVS
Tp3folBhC8Luc4hShaIlp7wMNYoFcIBUN6P1Mzbyip40+aTS/x711LDkz7Xnl8H3
OC5IrzlP2Ash49yQ1eFkhl+Ulf/HJ6F/u63Fv6WHKX8mzvpmWNbCpZ0WMGCon4jq
wrqsfTELNcG2EWA7okeubrmt+vZ8Of9zxrROjNlzAwIijiN1mR/xJwFKkbkp0you
Kwnojm55cB29hKzNAK7FZTmBpgW9Q2+J0fTDjJajBgk7DMyS3971U8FPOIJTYzu9
FD2dvuCoKcT83FUZZS/A5oMBEphE47Y7o6oVEfwAszX2AsquX+kB10B9QI/80OcA
i1hJ3eahPZdcbhmXyolLRQCLXq9jIHJbTerljrRFZT0gOzmdo4mpAQSPTBXuf6Oi
h0XKePYUhXHoP+mvOn24DOW4T8lIaWJbIHtb463iFsPBhBu7xDn1dNszVvoXuAg9
XNyG3fijI7uyHma9NSuj/1k0nYPHiLbpGjeKPGU/KtadCu8fttS3IUwNJrErfl4M
ACsv7kMusWU0txkxJT4qVh+588ceMZssYuMu9HkfaFSy7uIlldf1WzQxiiGS1kyD
pD7CzF+Fdly7ynuZluHaJ+JOe6mB0wwpu5vs8mNO/exyya+uTK0YawLFwWPgS0We
yO/sH5OGwSDN1PkqGBh2vLNedpLD/YgIXEAhiLi1v/L2iS/8faHDIJWMjoKIX1Aa
rNAFVL4/JTzoJcruBKUqf+JSdufVSog3Z0wWjVqE6F9H18PL7ndpCZ7kqf3N5806
uNlZpdWUTPbsWmgQHid0PADCTncgQGbLMe1dFKSEArT8LBHHeL9VlHQdnOAEcsHW
uhOyeUGotLMYiwZSbjuQBhrwtkpzbz60j+CT7geik2AATjEaQ8e13wzKnER1AkeP
ruhRgQlx1yntb2nCD1L/PE3ZO1ND1ueMi3kpP6oYuKR/p24ez87oaqgokoophDxR
rIKfNOy2uNYqSx2tupY0U22ftyNTQEatvfLcsVlrSl0WZCNDkf5Fl5cbbOkGcmZn
/b/l4XF7sDV7R0nYhxhLyk0n0L9N8uNSWviJIxMB4/CBZrmK5yakPzUBUXiNGmKd
t8tP0ldAjYu3X/W7mS1rEOBL9PuugvOdATqsHLNbVgk1n3AVrQ/4021VnzGt98E2
XhayWuzq9k/+EPAz7XmOoiGAiH0WHYroUbBYe9SGy9TfeC9fvhAKRxUxTRwsPUxq
A7aAUeTxRWJtXMeqHXOymwDbTkdhd/3rARWj1x5hSGxeCdTYUqSn5f1XYq0mAm7N
OAlKRdfpVl4H9/2Xdvc26qJQ25Xlb+IJulawPKwb26W6RGKo3KGLszNfTsnJJ1NW
FVRtSY8950I9YfKOVsvS3bUxUC9fk9NHBYWTiCckWrAM3INQC1v+NhU3j2Vgav8R
sk0qrn1yR4MsoLpG9Ta7+RDFYXWwHw4sdzFzyy1tHMPsIRLCTFiDSY2ijbcwtmT0
h37AKzwAVGkOWyKvY1oHAYj6tQtBmke6BNiNsJRM8QPYBuStdYCHbJ1nR+ngdR7X
1ORTp2w7vz+4Y2MiuNRfAaS3krIdcz/dzSBd9fRBhGolAYqc0l2QRiTpXs/z4/1d
snodCE2Lal5BqKi6Dtpq65kIfmbi1aRahGevJ07beBW6sOAJXRhMRyy+E+7FK3yM
JWJqVcVkWFJW+LooDrz0esB6MODU87AQUYPZgOP7wEBzrg8EC1e4V02+zsf8yRs/
ms3OwnsVRPCWEK9hGSPeCJ6NO4Ck05XC2kjT+fvwA8CwPtNVvHQenUHwaITGhnGB
u0biIALnzq3vyh76Y0PI4J8s2SLojIUqlWt9+UDnvM7iEAsIqZuAdYyi1bKTak7T
LghzGfN0Hd6Sr5QX6S+NByzwPkYDf6SNnFad7Zl8E77OmUvIoBEW/4zeaKzSwPQ2
e4IbbiG21SekyN0gvjBenAP2HiIOB2sTVP5S78Kjio+EGZ8Drd9EouV34PHPqMUG
kKTesnvwB6Z6HDKaNq+7Scv7NSnlWYoeobd46eGLLgo4b3DZXZwMWBg2CF9IiDNw
NYXO3iYNA0RsH2MLSC8OmLCljWLNhIPnYfWvzDVy3Ij76pA1HIRgKrepH+pX435C
Hz6A1TXZ2gZz488qUmUZCyUCWGn7Hb3QVNqUDimvA3C/mSgzcp2WkoLT+1d0exnC
MPAGYGEyVpDddhNcjOuQ7e0VHwcjtLRyUt4pyfrDBakzRyEtmEl5O/mmwpYtt0vl
kYZ/QjXkPL/18e8M9bh254+eC6U7O5e6jszB/EPhEkGrrOu5VCiKe4LRp91bVH8k
vnNwJTkYsAx56bE7MQLegRZlj2fH66RO/Lu448IYniBvq0U1XtwacNSNT6ZEhxd2
eNUFNd4zOepz8njWKLvAcnuJBorVbUjD5Ge7vLhAhOm8ZEMN5Pt0whHYC5k7d/3O
2pVYE2hmErVVpcmnag9/FOUXHECUKcgYRfEvRwyE0bfYiY8Qd+nY2Yzgr+Pr4E8z
IHAi6+ddFkTEjEmNKyzySiDGwtuGJ2umllKid3+jaWulBHgSiVPS93r8uOJg+3jx
qYYmvhdgAe6ZVLV/Y7zQmCSW5oqtxbJ3u1y7Vh7ZCmEbxX/vcSqndZQah/gNLRXv
G0LsIG757kWFbNUPVE+sya/RaJZ4S33creshXoP4mC885kA1NWO3A4ZcaqXw0D5s
eB0AGr740QCUrmlbM5E1WgEnrRAkAdN3mjdPr94ZbagRjHIoODcU9huiHWA7dkIx
Wn9D/lYOtNza2HGnYcbAKwkTUgGjiFZLEzjYybapO4+GgtbwaKuzvhsgu9NGZis2
fGOhvM2++a1uhEztT/er0zkS5FFtA2QRhd3oOrgab/4jK//4KTnzoM4EXFA5gPH5
UoMFF85/WemecFr6muPilLMLf06f8wtE6R9C+D8YtxRyuRcLdjkGqY57AQgZz8Fr
XkRr0Z1uaDvCgbAHHVGqW31seeNrH2ouudGrFrxwxgDPh7zwmWrtxtkeVGakaCOS
tO+VZr6j5Qxk21xSn5cp3BulPxEoifdS6pvr4k/XMpOUgwd7cE/AkyDG0pczEjYZ
yy8tUE/81w5ygEaWwUW4WUAAviO2purkjOllIiwCD/fyKUcs10FZSb8it0EfJ7fI
jrsMz6gzgj1IxWoZQCU1PUbwsVWYlYa3d8zQqG5vXIUGOV3kFb0cyMXjr/wTPiUm
WbXRdvb6DDsejtRbYzUg2ypsKTaJrSamW5RtYY0TvSfdVWiWzP9ZzgoB55Y9YFom
dDIN0yvZuZCvL+coirCfMWMnXw4YuYtv+VPsLelvU4cJKomA+10BBdLJBFL/0lZc
Dqg6jLORa6JMd6BCLyNzpWtUVGFn1S44it5zPA6glpuNabSb6g+6i4AJRjAeAkuQ
xYRLt6740GjSOEbz7rF3I2OLfwAvqeKjq4hHYBuZQ8G90n+3eBeyhZhp9TXsviUn
4DrgIuBXsN++TRoxMBF0e2xnDBjOw0f9iKgIFYg3sjSubSnURB/7Mk9c8B0pX8f1
nc/ihcwxO56Lo5QQTM3tBVC8aPneHEYnSPEitgEDvvGEpXcq61d3uyPIwcYVSKX/
mv5mpOaib+GNDtYNN9SA75s8g3RFewakAFSMf5PMa99TElZz8EgxdKu2aR4pEq4X
kgz5SGqpOH4R85zs1bNGC60RnBf9cswwA7b1GcE69i4L9I3Tzt7yibLQOsgLCwCQ
O8uHklzWt3On+X20owF/ZP49z6ycd+LsYdttQw3uyHylxQYGjNao/wZZdlgFEstl
FqNZVk8nbkV0OqmK4MARmg==
`pragma protect end_protected
