// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 01:23:56 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SsLXST4Q289jHG0PCioTciBaVJQ8Rfs4HRIyxAIyZmMEMHQQYTNv7tjzfpgqr381
7h1TIwPXOO1KQjJegli+V7kuD4KB76BNVXgWK/WQFYtTTfhHuOjRuLBAU4eHeaOa
FqB3VbAqaob/LfnqJc3Ifnpsptzjfw1hTvcNjYvyraw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10528)
rECjUTiIZL/GsQ+UJvvw9MxTUrJDEZsZ1EJjFFk3WEqfaKymD+zcYzmVKbq9q8ej
yHx5Z7yPFWoRLuaNWfkFyoRlt6nUq5MuSTGrjVqIlQwIflnoD7ch5DLXG/oxFxLp
G8+p8/h0iVKHyS1Wva9fVY5S8D+jLxkLD3O0roDqWBJ4kv5ZW5ikbfwtoubdTwV9
tBJI5YHv1yXZ6tjbl3a0aC+OBXqygRRPk1uLFzQ7gFJsCadGt5StyCTIwoNuJHDH
x4onVmsEMylAYhTtMy27YESvAbTklEy83zHObY6wcItnb0dGZV1VpC/k/5JJkes9
1dOrBp3U2MdqYGczFBGgJNba8A9i36Pxh6zbwE3oKQngPi6WX+QWLZr5nNy4jdoi
F2+A8syz4rbo/pg27ZcqeBs+lJVSrV0XoJdM2CIkFJu34ldb+eCyl6CBUDzIF8UW
xyeKr4iicEaLe/Hpd1KnoWeJl3aln45clcS02MPIRhgPOGgBxr3sioP9uoBfyCtA
LhxV71rzPZ4Dexww5wMQnWntfP7fwiNA5af14wYTm4POeCLU4wMZZcGq8y8H0Wj5
zNcWNrVSy5xwbWiIIF7pzvkYGYQVpfcPniNUOQ0jy9cZuwgOchId3w72GPg3PQul
aA6KjDfU5O3Gg8EX2tNVH6OaCT6XYLLyjaBtd1C2Ge4LiZN/5SWT6egW7mIA+v0R
sWpn715JGk+rsxy7+h+wU9lFfslnIMqHVDBTXnpX3RliqDWVUopwpnGh6Z8hu9/L
VfzOZHCDLC9Wwq6l6T+ozMe7qh/qyRk2+Z7A1/HO9p87XjKUjwysaeoHscyi9vjX
cL8pi5F8nj3Obh4iGRAG9Ayb88OaEQfBLBPfcxVJqq3QyYgFXm3CDIC68O+HC7MQ
++KCFqUgIN1bSgvlNVFp6HVs+RhNe5qkZEHzf6Fls6dE2IYAzQ+xJvsA8cIbURDb
HHinj6LnPWVKyDWYK48920eg6xq3iZCFFSVK+VLSemryoH15D/kzXrrl95y0n2QL
cUBgREzq7/avKzITIxNvBVA5jG4AnF7EQoiaD698L806eIjI21lVykn5MTsDqm+I
LRTc3fKd+PQEqmzHq+w7YZwMNA+XJx71o398UhE/ce7hb809nT9Azo0ZmFmh7b4S
F/1kc+uEkBYRweNeo2b9MHoQsk8CzRun0GtfXqAqLlpnPIrCS9vZFgpxZmC6hE3f
i9FLCLHQ1Ab6S6mUR/ZBedaXS+XlYwSQP3BNUcHF1daB/qb2qk1fPPJCYQ2GglVa
f0BtpJ8MWAb24UKu+wcz7nFiHfvJ+6NZ3+hp8lCWbKEczlqhCd/PSejKCMVXc9DY
dZrSPHTkD9v8lUCF4gXPbDJEfGfsP/Ca9cIg6mbPtvljJZTesrmyYQti6J4tHGne
Bt+S2PYIoOu/UsltU0SAfQahjZ4YQS8B4lFuheQMcHdN/OMLKKxOkeS4iZ2N1ETP
EdgcVLWMCryDSRY5Pm6F3cNpAUdqvPTMXFn6HGb3L9oRTolDq5Z6Q23Incyz762B
GqgTkQt6p8Q9KODYzMxpiTvfyeebwMxtsJY4LoWfzjMbXNzdJKN3ll2RSV8KkCE0
WaomX5zbIm114eS0FJDFygXghJJTcCEOfBghSZL6PEB9tNO3+e6zgy3rzR1f+9Lv
K8kzJv4O8MihAJgt4dVRYnh7RbGgob+42dmni3++o4kPYKk/oGBF9NOr7CjRdzN2
j+OQR/BMIAj7JkRYBwdPC4HiogdUoD7ulrwCOTr2n1qOejJyBaTB0iQlM1lna4Co
H4voau68Zr68StRrHvRhGBL+NwtlfQwaX0y2NJ2+hjI30gmrjzo04mRchcBq6Ri8
T+3LrKdw4mAEIJVBaBx+R0aN++vyTQWQV9LJcD8Oga9zfd7fwnAaGKRnewCpzdQy
4phlJplFuipQogrHPiCFUPmBNO2pAFQC6K4eU64C2vqebz7irp64WFYq6YEjega4
MBLWq3PTKfsoqYTL+E16PwYtS7p7u7uFvQKGkDcTsILTmqwBddUimioon+ntJeJh
Ssrx2hLLOySQZtjDVWjzkB1u4qn3XN2FupzK8s5bIs1AVp2+H7y6zVZDcIaMl5SV
4CWnymBK2TSKKLydT0KZNztbolVUP4uSSLkWwD+YIwwxxF40ztP08uGcSnERHv7L
Rbz7l3qHbWLKHSTC6LfjfayA02C/vtJKFaCfPKiTpmekxcRbLbuksi5mGP87B6iw
3V6FFURBF5DkIQH6Gjr4HMtPLe9//kGP7SDyOXn7K6VRpHum0lIzDajeNYOVmDug
bu6GLe5ph3/7aBMy4kSaPs0C3DSurk9UhQ7mXRwQR3gV8H/QfOM7Chb0ud9VVmtk
Un1lAmuMCVy8ND7SS4ctO/XEn/TDgMF3nLRiUm8pwC4d+1jqIUsOprMeFDbsy0D9
s7X+tHrrY9wuf2rR2mLu5V84t2AWOSWcJ8ci8qV/z0WjcPS1BmhfSkB1Jcd3mYq0
hKvSCInyrhIcOG/jso5dd8YqsBfe2lKOEs5alNmt4HMzM7TxAn25lrGlP39wMWeL
Drb/urI1J4aMMxaY8zYOjV+GC5AmqkZ+a0g9X2qiXvvG03Lyx8SBd3EYGfOFanIZ
/Um2ptIWxSmbgQgWqhlhGB12x7eHTnkuDhdd3jExAEx/kyUGl3M5DUnzs2zYt5b6
c48FVtk+r9uwgw4DiuxK+dAWYUCc1sipfx0rnAzQtBjq/OiPiYyYuUwI1CBzbXRi
ANYY4Uqorr6TTMv14LboQGSfK3fHz3chACunikAvzCOAIolg7fwDFDxhIJZtPm/u
ba2tOU0iW+xHTY/aNbBuHnk7Ww8/qj9pCw+KfQD8l0zwr4tIwoVONu+eZbShjVTu
oUsLKeGkScJHeL0n6Tc+poSb4ImOXdxfRaQMQQKVO6FQBpZHvm0HYkHDajRwy9IS
EbYm81qNytrh0r/HX+esIuijOd2oD/flqGxNxhqZ4Jb4xmQugpfHenPguvR4tcAs
Fe/DrSNTTNv2dfcAbiUB+TvE6GVRAumaYySSXqGgTYjer1YuGfs+Isgg/GHuAeVw
bFL6O2y2IwSQ81ctZkVCt0couxnKCQEfYf+xjuTl5L2aqm5Ztp65dPEa1X1B7VZ9
oOkHT19qgmTckw3Drq/2SLKioKv3A08ot24f3x0B5OtwjFxauRYSbg8xYZ3F5RCc
ePyF5lHdhm8bFZmNnhkDqz03dMwEwzm73Vsr0lpEP8nPc6Ye1KEyasGv0sZbAAYP
oPLHqUuxS260+zFOl3AT500pVPChxBVSrpLV05jSV0ToWCrZBveNAD0hpP3yEfEU
FC8+MuDD1G1a897foyssSYFugoY2oo1ozFGdI5xU2K9Y52BDeVx9vfwgX4UQB7Ti
BEZqSTyCSEq+QJnYi4/wUsPqAk5udzzAYgcEwes0gX2AMCzQyzjVwWiui3KEiH+H
5R5p8Mp0chBVw9nRqxxuGRq76bsYNs6oWq+jJm6dwoy0Hffu0LeUdecnnQ49XcI0
SzOC4e53JBwJiyoZsVfmiEiiSo2m16G9Egj6i9hnn9P0J35z3NtvNoO0JQO9/246
EbkWfSa2ZrJMXH1gI4nVkRcDQG1fv/iOcU7d7wrvYeRQwYF5bQyaKnyfbfIsjWu7
LRL3ATLMkD808Jl4vJbp4yDAhxe+puShrr2woXwZLlpc0q5zmyHtoroTTLLavmPa
WXfluxfwQlwrflCPnccGkgOgag/0wVsKtFjaz2NR2Tvyk9OhIJogU5VijXx7UQg3
R5VCMrEJIMzIxdSKpV1CdATrDKh1wR9+xgddMWGz667drHqJtY/AGR4lsL08fchp
H7j0jB+8pssAu4pFPcPiNgzlSjoFAcy0MY/16cfXtzdFdEM2MEwjGSF9Oeb1m0bq
yWajgcQd0kBmcnm5o88d0c3dk7CQOLjY/EFLxfrZHMahYMEmhVOt0QBT9uWW5TZw
t2SWRKlKOdg4r8dPJdmlDjU+6z3stv/fP6J4PvE6k0Qj780ocL0pjrjK767LX4G+
q968zrHnykWtdQ7rxCvpvqmunGVAK6f67Etg9rx7P2Hy3I622Iq5XHyKIc1K7Bay
Rk0UpU+G2sN6o9nOOTlZ7SqThafwba6JE3qJs3CcbamO41TK7rR29bq8dqiN/LIV
uDxbQaknouFkgcrzbjd1UGr1Mjc68KHMM3z9Fqf/aks7R+7rLwpKCV+2mVr9Bfqt
xZJnUJqPiZYplOp+6y8ztjhfr4I2kwftyrwT1l4E4vxpxvxhot8nTfvPm3Ox8KhT
t2UOfKnLFEL3M9FhzfnSgCiGcZ2+zT3UJrprsmWWXIeakXsPuIiXh60perY4uCYk
ud+hgXjssWKAPpmF00BEJ/2q3WevOAIE67SsccfVnwjKsEB4lhWW6iBwafsEuvOw
XvUJBAbNBt/YPY2tMHqWJijdKFHnBGP3mJs7CqUnsY0RQ1cM8rvShMQi+2nFc6F9
EIUoZKoddWVbsMglYns7x71KDh0IPSJbRZQQDn+mraKfouSvYN9dcd67Mmz+x03l
GDMiVr+6VT4BHXf+AttIHsMlTkGruk1JsfVC5ZlFaN59J61QfUSoOzRdNL2OWIUp
Do0xZdEQUsVi5qlSJ6lXcVMTk3Wbsc4+mqR+VwMP9S6wZuiHl4Z/um8P9GUrA45l
A+6SBnofs9fpOCfFDW1CWi1GqWYYH61kt0wmXVdcKhfR8RrtFAJpDK3bksdxE+wQ
80aGLlnroVXg0BuJu5bOYcgUkawf3Y3TyvvoDe9hUt0JJihxeluHQvsLyuZ29/M/
yG5THyt+P1E2xcq9lhbLbORcOIfRaKuop4Plby6TUqgYgJvgCQRb8o3b/qayTzNP
1nmlELTSoSsblaY8cALHo5P0paK44YAaOm1iLZ5BTXkQa3OKyPcvoE2L5s+pzO/+
hLJJgSlv3CgOv8GTqToiQHc3hmHxcOsA/WohHoLE7gYwTqBE5TA8x5FXnKWrGufh
sQOAMVDTynSJq6GgqCRNtBFf7VdOlKKEynSmZNY/rFs7xwlco5qes/M6b4u5vIs3
v4As10Py+OOgo6FyqlmOPoxfoEd+mnmmDUNpuW5RVyZoY3KZARD77Xji/34DWKIl
TKayxkmDDygTCGBRxvdABg8KTpk5jUX+vW8/mFK3oQDho0L3uE5jXzJADJ6CV31d
W6LihaKsIW/iKfsnB7XNlVn7zLEMsyZEzttYpZLBA8TATBWmWqvBfL/s+GHp6n1z
bA/CZIG7lk8KzuXq2sn8/KRP4qEWQ1P/lkS3UqOszJCIeQT1Lpov9eEJna1Q/RhZ
r5hMVE9PHTtUg8VdfETf2Gst5KDSbeA1QQN45XTlNYb3QKSZfChlHzLHPIC0iFvY
K1X9o3YwnPwJlpljKvBn/T2ElkOjLw0AVoHAIOYA9ECH/8MGomYoUrMYSBezbSrX
Re5HAL3u0EfdJCJyMHTiVLbefQFoyuh0QqlJyj8fjcxfk5pb63fgo1xt2DCdVWGz
Czxfoq2Icgeo1fsF3sOptJA+E9s1KiPCSDEG18YjyQqPei8cZqFrycrGBRopgZeZ
QVEu3+xlEwlNz7TgZS/d7OdqXP1i0ueCbPiHKLjHCvzeGjZQTsIcgYN4Q5R/GepN
IsKguW5IjztLC9Iy6wAO6Hv6RYR7r5kUDxYruerJ2GImR9RTgjEcqI/53Wz+GcQv
fS59Q+xBbNZTqpiJsliShZ8jg1SJHeGlvdB3u446GAxwXbZZCAWnGDuHOmiDJxh8
/aKvufOLYwGlVs4W51bMyt0bBLGMRCyucNyRS2/NlFutUQTqa6QGqJe7JX0/KR+C
nbttZl+g7JLVG8oyu96z2C+GewPAEpcqJYPZBVApmh6MVYEDhBZ3VxW0m5+ZmrRQ
Ogq1PaSQp1+DFvRtpiI1eGI/ROCCcglnLiQsjizC18EbgUBaNxEuN/PvQg3SCT2x
FOnNSZmoI26A+uthZYMpPaZzZjLnM5hGk3q4V9kGd+guR1+nPBnEtQQuQLb1BHc0
wkKfRqUMlTjczU8Lt1kgpUH8OtmHxM2lfRaqH/+BnrF84/aa3pZR+oEwMXt9Tog4
gaTYMwqWW7JRIITDlXWL8sJq4yLfKJwwSzLDSt5NyQVvicb/bAdAWnth8tbbQ6IO
sq6F0o6yabtXsyqRh9Pg8elM6HhuQXBLam9wCHeRSNgOlMP+WkvkoAJdW9cr5JAu
VT6cDRQlD92BO2/epXbai3w8X6v8YOAAK7yI8PSQS4EpkUzo9xmrMstoF4bS4pVZ
GLn5d87jap92m7DkmlLkDkGtAa+iBzw7ZCyxoqy0iyrudZZdX/SsYtxSDNPBbD7N
t1dxrJUEhCawfYSfzY2nrSj1QQ802+HvBrh0DQ0HYCGKU6ztScShyCtafP47kjZ1
jpIekTr/F+kWA3662eIQxBz1QKcC2v4v104g7ZLheqNqpw9mu6zGOPMdS5EE9Pp2
zdp7MO9Z9rJ7w1Zik5P+fG0vJiyCsFIfPS59Lu1ZeXj406E1LgPT++3pt6nmX6nj
BgQhyOldFSsKLLeM6nmVZupZUtPMTUXoA9lTSh7OEvHJWdEawRiUO4OgRF3wCDz6
8/vyPmDqEBEACciCQzAUuyFTL9o/BJI7ThxDE7AV0mfIjk08h+nyuc6zj83L7TUN
MMybvYueU6KnvgZgLF6XN22sJ23hIMEL+0N9EV1pdhNvAlUDMEzNI2uifZS9EhhY
bC3Uf5p8Yf2vQ/OSS0hMGmqByd8eYv+gZaV1bYkBRFlN7iYeVPFPeioVEsAIh5vJ
MxPENqbVzEBVNxyHzmy3LycSY8A54Dac1ptZg859RjyNRLrz8cY1RZhaTJHCs3lo
VvlIaGm7ApXVj2ISVT54hjKRo/x0DS8m4nXObG4WqIM5m3MldLjFKJQ9KcWhurEl
6isMZxQl82MxMbneGfnPjkZWF4zsQBsZwGGS6lKHIuu6hiEbJpeiJnSMfgw5qXh0
PxSF++eDcXkpVbE+Bqx4VEa4CzUqQUkV7zWFoDrhyK+dfNqjmru8S030wGZ444Za
cEHLJFOMg9PNxfQAfQDngLbJgC0Hnm8QheDO7gDuIL2tI8bMpmRib4cVyEKsdX3q
VuDzqZPwLENKT+5y6XFeoUa7JRflL8yOqPO7rjKIaYljkgRBihZHiY76ihOUkJJ8
C1bJWbEgCigDD0mlm5f5xe7EgQ1NdwG3p27MpoU3BOAy/bH0J/188X9QQn6NdGU5
Hdul1y1jl+dWtW7f47vCzqQsMoQzgNiGWYiIqr1Kl3/nKC+lojxz/Xsj4gu0MpxO
1Soaj2LSVQTQdFv1iqhyhExzPcqI0VzD+trnCsNGjA6NUH1NSCkQhF8cOWOTv6dd
KxV209lIsv9RaTDpSHJisGVM4U9i8CI+qP5Itc6sAmlsZJcbHvwKIxHyWh0iVCHc
jicyy5DF6eN10WkQ0WFqpvOtmoFr2X3M147JbWP2U0UEXCDLYPyHCcP8Rx7Qj0oB
CI0z3Emf5jRc/mVw2wsaW1FI4P0hzO0ijgKwdAcMLEpFPpi2fB7PShPntcZAPEES
OGYaTJbmEBC3z/QDgxAW+0DiOiNabO0BmBmWmAE70MFVcYKCMdMQhVfqpru7I/gS
Ix13bzvWoSguFwBPVZdsdn5/bGWrmMC/bHE4AXCLgZNpwDwl88r9rYkBLdtWNDUC
+fJu9WvzKQzo2IVGQO0jotj5XskPGeszebO+25JbsL9fRhD5WgIObjo9bC5v9HGd
H5YEvwG17YueJxY35CDS0lMcNLVq8m/S3sMextD0MA7a5xgmLBy9X8JsrUCdzzXi
NQL14Nl8FUzst7IRToFmFNomhmkDRvwT3PJAYdgysr71mZnR3MvZ69dteDdtmPEP
JPg+OXWpA6WnPzC/ck5h/bBtJFpS60vQpTBZtvBaztlhkVJFbzcnoDjLmQNLhgmL
cbpc7bacJn+Np58AdChRk4lz3jNcD5qmVQTlptLYHpiVIdbAD+j5FdYhDxkPw4so
uaxZGevaoOg2/krwPgisQETMfSG0kMUPWJEICJk+WD9EvMeutgofN4dCBGPcbAUP
9KV7EGpv/3fdKuSQvdfMe9k4YBG0BCTfic+kZW0YtlcWLmua71WtO1UuWYfj/MgM
+bkS2LO0AnzA7ajjvu+tkPxt88VQ/AlTf3lVutDQwHXJcXiPg9/oG6kGCQOXVVyg
AElE4FquR4hWWGySUoRvOzzJXVlN60e3MsrqwBIo4UQRE78d0pPUVQdGgevSvWTT
4ejCr8S7Xxsvsx8Pe3hqjZPOhSmAiEb03e7ZaVVOMaJCrWVpwYUim6VjM9S8kOVT
eZxUsbhhr2bfYIKRJPk3JGcekiAXyiaw7FJOh9s6fbHOZvPTbkezP5ylV81iRPrc
6k6ZQVT/z0GgrNoCuzO4Yau17DlnXpe5AAOKOQIt8mlMAmSVVwcDCZjtJ2nzjQyW
ibdaXktO3QntbWaq/HHAT4WlFk9OKOyCriSIeDQ9Y5Yp36Mx3vq/vuNvZtUhDtiO
X7blxusy7i0D0XbbdgaWxLp1qMnUod+OUDVL+FJ1lBnzP7CsKEtN2/q0WdTILUt2
3pnVSZJ2e5+vZc5z9HOTDague6uNjeEE+Hw49+MKUxpm5ERSxieEDRKiHPTnTeYe
lwt0+lrqt+4w6Jyq4vfuS/ux9mevrRdaeLzlTZe9I3cz0PfVdse5Uj6zfzH9w8dl
Vi3nyw1xJXPA7d9Bok1KmmhWBRI9DrXkIVAHK7kK1DlubpeAbP9zIGDyo8CrbLiY
aUreY7lpvNDGQlzwl2KLfYKEQvZ+hVFB8fAXLVdF/0TPoMEW1kC5KzxU6cTBbNue
gwhJcUvobQ7HpZ53vTDqlTFoBiRgq+Wc30aR5aVnrOLqnSyrx3rkSrNF//J+MvZL
T7QXCKEroKEnKrn0wwmLs44ZBiObT/qyqmZhdyne3WImY8if5xllBKRbwLmpjxmW
2WctAlAWQxSKEQRTI5Mt35AowEk6d6QjiOcS/zU8j5EaVAxXi2X60s46pW3TBbGn
QQ+hIi2lGbf7GZ2NIIDl0X6PIJNqpdfBkUbyFcnLEYNsmz7Ha8fpILugU242moS5
LGIYX6sM6C+avycJ9ANwD5xjJJreP++4cP+JdKSL2LdA/x0PzUc5B5oqqj2C3UBt
WVeZ1py+75N61DJ0H71rSu6ZdfmWLeh6KY6/gzHSG2O8ZiIWQq8mpNmXUV6EXF/4
yNvPh3QDVFDhmtbXd3g96ucK6aFtrc5TlMfDX1xpRP9e8nGRQN9fvS9zKg2RYOuh
7GIr+Akld3sPyQrJ1kycEW6w8/YsoT3FJgqsQTlYdoC41k133rVwAEOJlIkeN7rx
Ozd1KhNowBbqLazkjYlbmRl313nqkj5uBuVYJOtvAknUpVN/Iz19Dnra8SiOSS4i
TrS3IW8IWP8AZ9VH2nMIAm/VvpL5RiSX4/0vwJojqppCYYlSqryq9e4rc8oGPg0K
FQ3J3AYibPRQssOAOK/2s5SYw3F7DBfuNFPbWbBIarDGBqxG6qkP/bVhgrK6XOwn
KEdnXzwr4HdARGSinU0vUsiyUOgu+iflok/5KxEFJzNSvuW0tEwdEwQv5Vpv9aw5
0fPbBuc8M0cEcqkxE4Ct/DS1HhTvc3TrmcpuVvrDNoicGqo5d+vPs2NxELBi9bwL
/HbPQNAcIxSXZH0jsEB/oRYN9QKI9ivrrK4PPIXgd3E23rRrLeEKXqFyUIBTAfxK
x6KiFBrhO30N2ASoMZx3f7YPw5ZxFtyO9TgwAz1P3dYCANa9kLsUjD31s8daoT4r
EiVJ3y1BikXfCMset+MJMHO7JlrhChwNBLCMuOqQExWzBnOYjUhDeCmcH87VaTKb
ucsHTzCgSypiCEjYZ3GXmRoRzv7w2Y9EXGVQo3bijwaWEs9sUtGPsGSRsFmIuDCa
jrgruowIg/m4LpyjqJMg7bg4qS2A4P0zodqZkRhD3NKXeTdo26cclYQ+rkUU55PD
SFTHWLR4QNq0x+GJaV5muiSTkiORiywLAB57ievaANjBuvWrhIGWcQhRzBHZ56A9
zmTeh3alxSRAF6XdnYLP3mI5E/cD0mF7U2gEq2ZhfmHR/B66s7bXkRQFRIkZY9sa
ggkaTucl7a6AlIRIulWEvsFTcTLkQuXTFbKhc1LnSqowbaZg/4Dx+SOlyGJt93EA
BDHO6JbuDTJE6d6Q8m7htwG0T9rpIZ9vfs2hSmdZrfSiDOgA7TCZ2tjPwQ4mQ2oC
DGE69OchsvuuDhkuv8LT62EJYXf0ox9I8A7yx//zuDbLzw01M3Ht3bKgJOj7lTsO
Jj68+im0ziTQbYHCDxSA+Q1Qyuii7sJXRHtar7mcmQmHIqXactBBr6E/35chI8pq
ox/p+tFDFA1gUxrq7pVoegZqXRiiKxXbYDLkQUwDcF6u42LZ51S7DibITOzf1QQk
VTxiANYyIUuPDauIPgRwq6XdFVJJ64To8brULhPKYK7bXbL50eAcY83e9jhyFf3R
LRTbdi+yseEWLNaiMT01n05CdhfgseM7h7FHowiTty/aI673zj/YynmLraeyJmLe
5B44KGEaboqLOpg+eXh20YE6n13FYN2Zl20huLgqmQ1nKv1dI9Gu7/+cwKbgiuVe
07lZva1+huhDgsuUlft60xZzC1Rt1Tl7aMq8+/XzcB5hTocTnaIePG6RgCuu8NOo
FMBekPJ2e7Gdkr/22HXsNl+NT/SXDFY2gyZTlMgoH11e8XXSPL8OyYsJq5N4SS/g
GiQ4RcEvGnt1pM651KkkppFtqEWep9DgNU03DAltXDYjasbUxcpKaymHrFblo/MG
fIkC+Tnpbt24gwuU0Te24raIS8jYpTH6mzoB7fiK2nNJGLq69U8vlGvbp4ctGSf2
6qNEFiKS6NdLmR4llYDCRuMAFc4vWR7KSIR3+POaafnCKB9VCrsBAHwy6Qvk6IrN
/j1xgS/HJJzF2pyyDuo6lKFX7+WZhsYg7vFrSWMd021LwuWhYSaVhpdjrg1CSEfW
hi0xeZLO7H0UqYXO7hQiT0VVmfg0LeVobbbhU5dxRVNBvidzFBPnF7YG58CZ0fcU
xAOBcWu1hYXoavYVaEqU69eaZeDTDqo5eMGEBJy+EASwwGlXAF1an1SxhvKyY+Py
uxFB97Cl1IbBJILKihJfqiPcZ24V3Yld8ukCGKAcOAHz3J4vutpsgFoIcTWgCYKl
FFAE8taT3znBpYZyjU8bjo+zs16Dt3bw4A0R5kTDrAL4FPrZRLeqv5unl/kpzzsx
nCkYGR1USr02rGxW6ngoNpYYKZHqxGu9PHzEcphPyupDnSc0aaYLKQ2DrUKw1ygJ
Oyy7fEHlMXenpIPiezL2wpxiZNe8d/pNrBTlwG+NNvMRE3T+JOjis6G/DUNT5h3y
TGLQtx+zsAMBSzgPjoFYlwp2hs8CMXBhD63EHXeu7APCPyJzmn+jBvPY63B9lQO2
WG2YaCAVyzPGwU2wae7ib33QWUoHKNTKRCP/Z4Lh3GQF2S0qLj8k+5PfLGV4uM7U
Ztc6MvCYolZK83FDUABrBKj812OI9jEyqM1+Itu4CNau8wVJJ/+0kYv5jp9paHTy
Xv0w7n30AeTXoOsZm1Iwk7qzJmwnZxziB57UGmBUkLJbQkcgwfjRzX+0ig5F9J8Q
nXArBEnkNcQl3c3QFkRizggghnUYp+/J4nZ8WpZNn038U/5i3NwLnVN8dbzlrwJd
c4ohdHaGJehJzjTYFBxpr7Tmqcz3E2VvN6d9Rem9/HpBoCcawfEJXsJ/H2SPCK3u
bv5sHabvWbp+sLsre9EYs4y3UfI1LnPNo+oMAxmVGCAdzEi/kFehfE6Q6XGqL/VH
/KPXG/hcsra1pDA3Q7yQz81ZTj4bBmTit1y/Nac+Ho9Yk5z7oKgVtSSxiwjXApiE
RC94RK4BubkebZZIgLX1xIMzQ3mR0xba3jQNu4HbnDh9RYj2w2VSv4FnPaFAwwpC
p+FNTO9SnBWySAsSXbbYff91akyTK1oqC2vn10IoQdI0sM8M++Tb4usjGLKY/Lda
ASfkFQK3WAYP1Nah6pmIQkelGw6Gh6I5gYoQBiNk/riiUNlcGrNW9PTUquYgkzlK
+05zAhwgSHyxPfa6yCl1qdTEVGFVQxOEQWsLXZKrqWXJkFQ4lKPUQfY35Us5Fb/9
lfs73MZUK39g52VrxWeqvxBhTB6tulPp+Qcg+EC3z8HJ7hy3o5KCPTuCWAqRq7Bl
2pT5haz5WIDYatxNePEfmBf9e0//XWToLdV+9Kt5/08rFIc99soZM06LqZ+H30T3
TDwkP13D2WzzrJk1Xy2WumgCObpuivbyGWgW1CVCyOr9swTLXQyF7v5V8u2fj+gt
JOeByXY/80WsXY750+P0i1PUhR0UmdBq5LoU0YaL/Gxz5doINCWgXUeK2/cHmahc
DG8p19zh9hxG5bLekCPqOpynEXliYiyVch4L8BAGqk8K533rbp06kvyVa1XGGBCa
+oSAK7w+lYsGMyjTBvsCtiJ2UOKqvK15oEs1gxyU3gium1EetC5GciAKL7VBHrFz
NdIqcaIFBHpUiy1N9PbpWSdMh8OgcxmXpPFja6SPndkCrpea1HTgy2hUcA76VskG
4H9CCjbDV3PexW84BtpevTsjE3eZaBo8Qim5iRe9zELpYBo9/HKIcuXB4O79yZeo
n0tYXDnKsONJhKrUb97NwIZ709jxRu8MeH+PRpO7WHygM0xwlKOEbnNFwzxVE9CM
WL12JA9axKzJkI5b6T6lwO8Bb2LYrlij18r2EYF1l4f7fccyylhWigwgO34hN77Y
q6APFxFznArZwTjGY+u4iT1RrQAzl+KHUm4xYUnfGWlBB+TBp4nJPsbWTYpa7SNr
rbycoUar9XeXU4WLBqoikMASvEXRPoLNWglesKTiejeFr1ff2qfDvIXypDGSnkSq
Uwr0D5WCL7D2Xj4d2DqHKo5l32DQo432o+goik+DojXsvsq51+O9A7VaSqUiA/dR
a++xpgMQaCH2Y2Wlq20ew4carb039yRmlgkrjPGNg/klrB+bpbPP85WETUa9D6HH
i/QDaP0Y5SeDOL7oJhiHERLa/906oxSLyWtb5oAmE7JVgu4PD6dr07YMkpDM/kEf
T6R/OhBCMJzBx0R4fV7o7GZVpsApyX6aq7kPvB7rOFYjnZ9+erxAzTMXhoUok9Yp
r1PkBoc5zBJiMnFiQR2Tp5/70CO71fcbwpSlWGhvzYUDnbdfUelJ8rI9svL/k5wj
XWeV3mJZbyhnwq2z8hVkdaJfhDlC9ZsiNNtEGCou+X/t6hwoISn9Ka4cBht+g32b
lhXBK7UNUA4Hh2GXSttgrD1O2hqHkuuurMm6U13I6wuWhX5oyj9db+pC1Uj4zaxw
cGNeT+cePW6pyVaVHuAmwoCN6VS673X3C0rqn/KwwJ8/ZIX+REN+tFtEa0b0pQAw
yH9VQCfZ+XzVUe1Sh7YzCTp0k1hmXhu6V6Zta4z2SHehWfEHpYYJMplsiihta2b+
O/OV5P54POtj/vzJ8U7dPGx4XgSlcd8feGGRy8C+qn44f7jpHS7pOVGa4XJ8leVh
LjIsMJYxc3XMJH2DT3zp58JVaPxjWnr7vcnLMXqhImaqAOy64l43BIZ1U/KqEMZ0
54Qr5XUxdze4Mn4AzJF3NC/q6nTPxLzuPQgDhIKYo0CSbuZ7PaGCE+LVIuDHJjPe
ZsQMFdrek5OlcTs3bmqRwfq/15a2LwkHf1Y9tENIJcbnkvzUZTixKEbJQJn63PER
dNXOuqE85PcSglgdgCKN4f1mrkxzmsgtAzxDFHqJOhT+u+ADHYteCfbUTzBAa8FD
ygDXrCHdW3FAKCllnFUbvxawazPKAIdcWhvisj7Az5dudTNzubVJv8bEnupQBXKd
AM/N7k7CEpsvE+65ULjGlzugJkiTY4eiPMvRFuMmNeLhFRNLwFOTQ2zFJoMxOvq0
I9oO0T2MdFq7R337qdWwmqf/YnySuABYFat1JjnnKbfeFwL5bP/lL3Ykhx42XrIc
kpvZ/jSGMEcyaQhKgIpzBQ==
`pragma protect end_protected
