// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 01:23:58 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZhgwrTnqWpYPCNyakr5ESHwD9gF3XF186Iy9OE/aR0zrllzZyDlLcqT07ZASBS9P
uLvapTSnONp0R3CS1e1klqFZ2RoLyFPvCS0+U/UiWhx5NBi7ZNT3xPZXgc4kLkSj
hE8DMFdk6p3ft9Dvirq0vVz3SLtZ2Ujvro4N9KCtE/8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2976)
QMRR9T1ob6omQ8WGqrtd2Ee25AwaLRih8FwIsbxiXkuvlV+Pn9TW0sBAh+yKM2Jo
FVsOKAfCkJ0jkfIrVcvZ1Rnv5QXPU6370z1k8EsHSeCrKKMLgi27ogSlDZr+bwWE
gtlIlCB2ng5V16TdV01ZtHwuHa1p6RGDTgAubRliYFQIheH+eu9VycIHfrVWBa3/
TSzwpPX9JE8jbSloYfWY81gYntg2W6fP+gwseD8QY2PbWkWtMDFAUv1tBXtV+jVW
S5S9/5uF6eq+x70aYjl32rbumtLHkthk2D6z+OTlYuebWE8udiYzWkwINPea+SHg
8xWqgpiPXvh6i1tiFl+Mi1jNor1utggUKtRs7wu3Y7lZLtpE6Xjxs00ZcE3xkxeI
WgTgdFqXFYabuleNMbavugffdewpWaCs3OoVLdO4ZOWjnG9Iw8KjTYB2/vohHpRL
i0CscUE1Ma5gCrWZRgR70VUUsW64BT6XjnGeP0nOvXzwZLA9cJEKmh5ZN9/+xzeW
iC+3ZUJvZW+eMvd6g/leY3dHojQAKlbwiH2ipcNsEKJSI6LY8lLHPJGlXfUv/ajO
aiZE3efMIu3JVKmQIdmHn1+kWExS2jptS+I4DOa9eVde9mJmyj1RPWZJfG8iTyf6
QfVUsb0w3+FMvaRdIOIWKP+09Fv/cJMDGTHemYwbUK/U+d4O/OC2zLFW7rydz7jN
T5KtOiereFgqpjC/9YpucDxgoifWDCYIptk9ANPHqYo217E6sNqxfzZB1TySNgr2
xuB/4AcdgiSgyXoGLoiRvppCPx3rQ8dh6unf1/djrW/k7/f+/UCg4iYw/OqL/SOo
ipacgpXHYlIWtNZ4LFuiE/IrcKj9SeJKYf7xur7ctLrbcO0XChfgmjGCa1n1QiY8
tBG39cdKoQ1VnerhfX53K6PkNqjWyE+h9fR/N8GG/jc42IIzKzu4nL/7h7udhHoa
jzBdrVM4TRi1ENbz8UWkF+RBFEkcDKJTkAgt4lRMBtZxmdDXEHPGf2+ZTa7qv5x8
7R4/uH9VMJm81kqic5O/9Z1yfEniXAYmBOf9rmFx0zqZE/mxS67tRpnnZ7hwlhUR
s7lwfwnDjvGs4pPvMTAwwSHTW6BJPHG7ZqTRbSpGYDpKcJuf3Mt6GJ0GXF1VMBph
+f2Q7NmDN1lVlOqketq7EgJnJxVdCf2Im94Jsl1T8PaIxJbGDcdma9wBJ4ausguP
4j+eGOSIyOQmp4nAJ7hXOVRlVESOJ4Dlnq+Y15R/TKgWYf4eTLAfh78SPZdVdjwf
ycrtq/ASvIGx1qR6dykraSEZ9zbSTprgZGxGDNhuGRClesCWDjItyC9SsPkq7YhM
RG8IQ7ZdESoVit1aMKjrqNtl83zzaKzpsOkU3yWUYfDSzPXWLc32h5sREBoOEd6/
Vz1amv4sPI1yPTQKHMYMkvkD7KgIWO0b+0JHTpElE/LHrIlAuw2/k8vBdeUPywHp
zsf8lTEWOd4u1egfuQhNeh1/4M9vTq4kyLOfVhGjXT+LOvDhkh6+uo67+KHtwU/U
DLVBbE2h2NALHOLjPl0C9wDJ6v/vxJ5bj6KnWdtZR20Vxm8mFMqsC3idsXHMNMw2
NoQXBpyNAaURiVZa2NUbsJLs56qnXcBil+r4MsKkfGp3iUwwCPkJFOxZj1xTCR8J
qJitTaGj2laLl3+7FalcWI+AkXm890uCAuZOTxpD6iRqTF7d/lUq3FcsJ8qi+UfC
vMJF6WkqPr34fudC9FoLVkperYDzjmEtIVvtxx9/dcEy06Rfc2E2IAJr507UByxK
TesZ0T9+qP3hzI2Mj5n8EU5h3tl5luSXWXt94BVN0JcOF50GLw/qzH8slhCVkkGx
6n5WMZTZDrIuCR/u9UDm3QhIj9Zr7aTLZw/l7onmPKs/wKH8zhdr9mSHExgmiqyr
uTRGVHh0NBdXAK4Ord+Eo3y3hmIdaqa5FrCbmxkSzHxNFu3Lq5OU5ZGvbWVlPqRm
RIudE7s8Hk0Vw5SQSsHeZ09I5yeO9oj1JVrAi0TbLiI/4g6MIsmG87lhE/Gal/qW
41WjNnWnhfJjEx+Wp5rx9gCllyP7yOfTSlw6TxIo8mzMzQLvhORL9ujk4EmKhmC5
BaW/9Z6LTkF6JoIeysXx4y0xyRbnGxqzXIm59hzDEEOSdk5kak5F+x6Tyq4IOGrh
UmaseIKpz484JXpj0pfXfJEEdmRXLG2EAKw4IXoFy3Ek1DWq5V/38snQIfz/3cGN
EbVNvHsDGtOyANYKOJX1EvGWMyDXWozVP/TZYZSjUv0t3cQnEZpwxMwbuyfzxoIa
VV/xdf/wXFkeejk7TOrMMyOzmSBXaRg+LfYYsGXMvmNj+X6H95QH4WS6LMvjr0v3
Mt6JMfqSmTaGgodvk6xngsTa22q9hxeI4sbcKb+0hj/YiLGVKRevw2mqvEqdYH/9
urXnqSLjF8pf4bQInQNOoHJGOOadyOpe+vy66EsiHHM0fl3Cszb4L8ZoF78sZ6mE
A8pHAtaTEkYVLVYkac15/5RPtEEqD73/0bW594Cy1hW+Re6gqlXxIbkbsOkm0VkE
gOCinXo8r8CuHXRA8fHI5A9pqJdtRT6B3svnEXZUVfJAsHd+a/S2iZ4faeMVnC7s
3Chjw0YBa3mc6ytrmgfJqEq7LHbbFbDW9Uq2vLciU++doDFSeynPEokZyotcYvgE
9VY8y6K+YUtp+HQIHrczw5DZUdbQGCMmAg/GUqVD5bHmeSorwNDo8F5RnTXK9vmq
IRNxItnKLJwj2eloflgHorpCagmKJ6qlqdGJK+VLUVorNEcGCNRKjbIsqVOWWUSN
JFWWsqLhAF6LJtq8owtaqRFpvvc/6Hrbea97O/DO/VO/5Ec6l7yw3qyXNJ7utPEA
7h+eD9/laK9uNZDcTLyXoYJa0HT/EhXqa+ZWe3+MHshPR6YrmuepZl09QzJ4AtCX
rtfnZBPnvKJZ3AEODyhk3YbYVic+6qTkUTUaUYziq81it+Z1SO3FrsQh8DLd52sW
JTG6vB1z9WnQSVPc3NE8EOo3XQw18KEBtSuXLyGo6PGped7xFhQIpJOc45bCDyi5
MpfOL8/RQmVeb1SQf5xMx1Sm4U3YvqbaSCrfXJEqybEyUT8Jti1Gh1Htr2Dh5uVt
FYy9Q8QOOD/YTjGlmzw1z7VIQNPSxfOBtu3xq1MnBPvSsP8fYoWrLSnEAWkjsyHN
gSYDB5uYwJFMqHFnWzNFNJxyCUy7v3CZJreV9Xiqfl9svF6KzN1JMUSUht+jmGIE
gHEFjtGIL/e/ty92U3NUxCPL9gpyutkYVafEPz6v6eS8ODhlQo0mtDhOYD6VDJFl
FoJHIJDYSxQ5mSVL4r7GhqGqzmkfjBn8U/zkzANwqUqUckGJE3PwLIB6/1RmAZ8b
/pH9pnLfzYAhrs3lLGE9NFJTo6ACdpWRu9cs1+pN9CB7uuExYZB7+tEIkP10Hxaz
bKwt5B/i5X5GA9yFWsy7m6Dx0xPeZQOdgBW9BLwO0Uy7UTv6bY2I2Wi9O7CW8bSv
Z4B7nLhGJ6LIC/DiUF7+zrymtwLzBM1kAGVhrwaycKY3TLJVj5NhOORUPnOw1dpP
aznCVIYM0rkzKmCzTX7E404yobJd2ZY3PX37doeG55Jbrylc+V82UxKgk6Xod5TA
EYxbtigMOkjVOUPnlwltohY/4TlG9/0O5KwNbAnZOH7QxFHlcP85tH2PjBDSpmqT
wyymeZzVUGgMgQXqrlKnJOMKfrEQ6F8wtFMVJBHU8IMMLDijTV9aYsl6JrgNFB1P
a3MhtDZkgg4Hjhv9UJNtZOyExbJ9BAsyE8tmdEDP5J0m7E3XS/fYmeB+y4SFQDLj
D1XS9Tcv7ztkwBUpX1OrpmPGjCop8CN9lx20EuP3rJ9wQsiZWbOjGGpP/Bj11Uo5
uiOD13O5JRBJeRlNffqCB/Ef3mp7AK/k+FfAkH7RlYL0W6+Ba5MTCk8nigFt+rs0
`pragma protect end_protected
