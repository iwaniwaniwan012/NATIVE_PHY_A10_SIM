// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 01:23:56 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
apNU9tLEC6pbKQ+VsWtZyoY+9FSLMMbZMfu9VPjZ3go7k5mIDxWtaz5b+/pabr3G
MnS9gLIRcWKWOd3Pf/y8USSD76OvP5OpLCmGvOEW5PQI+s4/Xss2bSSszOvJhD8u
pNZ4ux4rXI0Y66yUUUMQGksrLwLbrAYsBIbfmwshvHo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 36496)
EOjnysHA+mkprv0esqcK83pCeYg9IyLpZABNuA0AxnP3TJrKoA7w4KNVGwZaQ+pG
6Li7LjrkIdf0fp1Skoik+3IdtTKXQAj/7+G373uGCyDIZ9kNnJ/zTMsNLuSZnGgd
R1NkZMcw5VXk5eSFzmBqYX9ALCeUe8qX7oOv5Mkmi+iVvBPriH3UrTU5PPZKve+9
bW8iqe8FSRIM7OQNyA5v2DcwXPdN+Cf4W03G87SF2hKMfQCMeZiVwzMAqE38qjgK
2NMczIvneyUhO3na09NfcgE7oKijYgsAUGLHQZPKuckrlWZTCJwWsXAgSEds/hQt
Uf0E5W7jCX3fZT+xPNFvQ1+x5U1DHRTmVBpcmnqZ4AS1jcwIB41BDa+M+HRqG3Ri
jlwVFY2TxsIbw/7fEk7FvN1kG6u3wKGrDrs09/tRgWhOCwOdsfmsmjeTAdMICwsl
R8RHQE/mPuK36f9qcg1/e2pZhNwX9zXh1eM4gjXKN8z5WPvDWLfWIxltAYNGEwHf
2t6NboMqEMDPKWokL9tKIoGn+yJrzYND6HTT01J/i2k0LokkPUJeoFfu2MZFQUdr
CdR4/eTv5xS8R6MtxKL2IO31pN9JDEmmASB6eo3pT75/xw7rY3VT0V9EqCTnHk1h
mybfE6u0m+cO1PsqdN57SE2AV34tjDjaOTCIT/TYC2y09aCMEufd5pRVFcsJTzDO
d81+Q6GmrOJU9863utwMlts/2WDJdKFqOftW28iO/lIDiZDCY6ZbZ0kZTXOCdABs
rI+vxBFkLTRahiqDR67SKhjoetLu2SM915DmRG40D1LHJfEA/OsIZ7e2MmSenq4F
zRryK/Pyg/K4csgGpwIoZk0Qhw8dAh1yez4hcxigzAzicRYSl3ADQG8ftbTUlKzX
xO9Tz70CFgpXJiJstUspf17u0PVwyPOeNX9holohWQwftIflNPykmFGtASPc5hor
HN6o/Is84JAJmhZvBVOw2XvfPc2kxUEtSPPdOD9Rqu4S1ueNEZp00OtpOkotmqI/
sF8m7VNh7DJNqgwzExRSp7og9WdVyBGuefqNq1WECwq4yrh1zbVUvJGHlkfmcSGn
3ia4EygATpLoXKytNqgfniclyQ0F2kfB80hCBXMCh61CSkSf7tTOZaOPG/jn1HmY
cdFeMNb6CLMAojqVbkEoqAeIDJjCm8gRXzAped/0ymygRkX3fOo1P275WrJm18RM
ylzTGTDuUQt+k8a0YZ+zK5vL/VPd6N1i39U3//vLEu1s0EoVGHMIO1s667RPV0hQ
gXw2/NpaKZNgEEOfXiJ8Y6Ck0wSnSUur4FoK4I7GwK4qWFoxG+948wYODxq/nBFF
/wcHAfHWR4f1TKtvVFSxljz1ff+jrEU3doKtSJeYDgmeBTVxi9r7ILuXvrMM65y1
edtI9aYbUXcahd8Tn2zKnkJwSvZBwl+CYQogKhGHrvBn7iLNZSEXRq32zyQUiOZw
wUJerzrSfUV5Rt+kykOar4aXjYl/+LEAKsqkJOesPWKUV6dYJcpcFtnsccibscM1
IyD0Bu9TLQjXaG94PBfsr8D4RrWrYF2Mod+50SxkrwommeiwFdTuRQpLUoibxwA4
LFslDT1zPwNko9KxMZ0MVsobcJpZH/1RRQ80DtMlvz74UrhwaV0kKD6uFMhAdSx1
eEZ/hMD/Krg7W+JOviIiY3nFdvcR/NiPbh8qRJR/W+pMTPu7nFYOMXytXYfH2q1G
OXqm+01rJuw05LP0VViEz+qhKklipUs2m/F6jze14jkt4n4eOzi6A44ipufXb9Jc
2YjzSvqU60b1LfrpoXlL95mLbqVJ0LBC5q5smzsF/ptP9D5Swq0IVJOhwbgTqzbv
Q6p1jY9RaAsPr3zRnou96B5/Gr9Q2NQEhVXnKFpNecJgYiMm/BFa0fh2ti9rEX3w
maYgsKm9FuONH97o8Pbd7XSmaHVyJx8wRS6jdUnaO1OPIWp6OWKgHhLZcH95ieD5
RelKPlG+0G62TyuhvuZJT9vGgiVSBL38hjh3cyUsqRmYLjYItIXNhKQFm2InT6EO
BpTByiftu6mr/roXLxRpEN2WaTgy0RYPZTaplXNlOz/+rUaanLCExGO3g6jeSGEW
uDzb4IDk7pla3cF46HofrXYJEz2MJl82ysrvrYeawxpNjZ14XjGAUOObFpmqmH4q
3fT1fDz7mqUvACPCliqgtzubYVcl2hyU9xR/cLCoudubUkJMa0Fhrt1siQBaXwyp
7b+Z8IW4Tlx4SECJOdpQGPGCHp66jC62FUaFMavRagnLiXg4m+ucfZ023Io+GiWH
823Ix0P5OQcMm5kGAt32U20+RyWJct7cjMlzvIejU3Bbvwgr9Ch2GT9yNHMPWctv
MVLM9iB7kFSwKgaf89XEBfx9KbnzYUvKjobq4o7w2MZFP3PUpObsq4roXwKvC2rR
VLAtGhUCB/XR3Mfqu3xZNAu8VU6k5er88qbiZIxdFgWpfPrnGBo50XWafvcgZpGW
9mgkD0+FUZxNcpNeCgLLTN2x01BS83OUpy8G/nhh0vynxZ80xljwbRXMK9Vm82Kw
oyOp7giD4CTiXmzHLKTr7QAi1hNb0JZhgnrLzSBBxUDdCPks46i+Dt2NaHW0o8CH
0jSfDRvoUj9cp9vosXjmHt9fVoVpSRSH0jiD3uJZoZTHVOEOp9J0re80mBU1NEVb
38UgGoejJ57fWncxDZ39VuYcEKtCRq3UOf1+kuNqcNCvjCAe3+86RMD5Qr0yMx2F
8T8sP0lGhn4HsuEPg0zphtymAYoRIosS40H8EXQAveHi1Y70M3UX7d6lwmQvstYa
/vZlBQpWu04Rtpc2SNrIs8ZiXLyq20taK9DSZqMI0AZ/kS7aonDIt/IY4FfzH067
rV/sMpkp6cHGi9h6MNX5gSHzsaPS2mSRPd+dlXTGPQsPAMyykBWbPzoJDpOzlXCq
Ru9ysu4x0RxYHQ9GX1/FjEJE/N89lyNmD8V+20t2QoiaIpU+oVmqusdFls7aEDXy
nsW7IjwGnLWihhOSwZnouqoNXF3BTUWsGRhjLNUjz0JndalGWmaMLaw3LZs/9lgQ
bGlWy3J2AmHMJ3XObUbqoTUxef+g/yhun+jPBTirSh3/2UHY8Ck2B4ekeW9sZFi9
4uDxGg7fQeDgEU4jZD1L1fkpsXVV736JIx8txd8x+A3vMCQodfTuPltNlY5f5KPl
sXvt67eDJeZritamqKuPn/qN1R5NkGJHksy6BLak310/O9FJDUi5pnhva9uoBVQY
bh2Rq7/SVC+Au1t9Ok9N0kc2Dowye/EQ1Uf2odKhu36RKHIl7VxG5JiraORWZPSh
pJAZn8iAPS5ASEyPgqIWUYy4V4z+FGPslfbIWklblfB8LCA0cGVHrbD5Of7psi6Z
PuI7bnLkz8wyJa+o1ZpPzjGAujuZ6wSHksi9ChIcFrqC2D3iM/nSv0OUd9sCRuHp
AAEekuhtjf5WTKEImTiyocsIcIrEOiiKUVza7WIRaGTTeO29sMksc5BOHKUwRwtu
amsIG1RAoYWq7CbcK9q9ZhXn+UGiNWNP8nQ5iYYzHAyO6VGw3wYBin5V0OVU/3gE
JzQoMFrR0PUf+o0NI9neZS/QOkKcJAsfMv/Xkro7d041cp+KImXwBQhAAE3V3UPm
Pp0e2cpvBqCio0eRBVlX0ginKMljxLsB68Pzrraz9sDve0Fm2/FfGiUp439C/f4e
APLNpIXP9ykCWegLPOz9rjo1yWQURlUB5eMa4MrUlQ2N9LBolw55hHZOXdfhv5AF
7o190rGPxYdZ9tGI+9ypkgHUmKY4gIuuMGbQgUA4dwhMrLuoNf5jR/IvRJntmzIJ
/J94SdkelRICQQDNIqIbZF4181xmsFMPd++x7luFHhSkjNtxJjbzlk862g9Xt7mZ
ZavQjd25FJTCkoP9JWhVvkvemjMwkvqSSXJGISpfz3TrIP2RdOMUkN/SfKMnEGdh
JyU4FmNk+UnA+FXOELBHqeitwCB+iecK7Jko3q0pLJHBtkfFGgwx6EQBzm09Qg9X
2yAwAHn5QUqI6beU0J/SduPtkq8sN09N0O76mqDzeSLbt+O6gege9MG0F+98Fk6J
uMcN/ZuRE1PgctFlGkOQZBO3UxCm4J++Pv+zToOVwlLW0PWHu+lQC476sNz8ujbq
rAXlXJJ2VQ839r5K8PBf97Vo9fFq/BzE/9VsMxshGkLrcpixWpZIMAvZP8W2KfEn
dDaqx+/FPwmP259JN5Qog88NYWDVbxm79yAKYnEUtOzLwBeHXVfYau6RkLp9hj4X
m76Mc/8LqymwfqKm6e2uEzZbgHvfCcncwj8K8BveUDevWgIgfNxCJDPwWAzom8hT
KpkNE/4K44QiVt4w9/uIVO98NPfquMAmbCQfuA9gwGmryBg/iT086pek4Qq6qZe5
9McBKZ/7lf6y+ueVGpQZ6+i0Imiv380tUV8PJPvvcMjEloZp/IfOtTsAvGK3wL2w
qiiL5SENItQczJvZ4WJsQ0jLOIK9R3lBLv37Su0Q95DNqv0x/UTAISSUJ+5Ns3pB
LGH9D9gNIUB3Ygzxvg3vzqxSo2n29ooEKNWMrXo+Cw2rvv26cDsDR0vBCNf9uR17
cVr2mcPB2LKESlKmPQsm8DAc6HSwFL99WcxWFHUUyxPSnjMhot8mOriNOsvKGMs3
YzijVV/tUDCriDzstopk6uhMjDA57s7aV0DP1PiClF9gwdSwI9FvGaK4v6jRXugs
oerWLd+xBS5b8qwV/WcHaRJq0ETOQ5fBkywISNiSOsOmuNbG9MtPejBbtyej76JJ
GPNHeGCIWks7jjDUEZYNse6ihV+nnciwKZ7PmqK9CyPQn2IN1Y4coZ5NkzB4scR4
cZKWX9wlFq7dJJgl1Zbo7/JZGjCXEWGLHh3kQ13B2wQ9pqiPlY16qqlSAI5dylQj
rJ0RsQgW29m7wnATZUT9Yw4C/Le4w56xixxectho3a/4fQ5NnxMrJXwHK7PL0JWe
blvht2osNBAm3TZ+5mTrBL21DgI4OV0hM9klRR5DGt6DESwp/ihmeJoBAN0+yqco
6wpjX1+mfOTkAjPE/X/yv+QhBqEyNjKU8Lu/ACyDnPowbkLdznQjDTExx3ccE2A0
WqYeoTwgcAah358eEQkGgZbWDlHRP3/Eam1Ncnhe6Tk8wkynsZq0BX+n0aSQjIe6
qf4zHBReLR7IuNb2hkitNuWg2gmFOz4w4zbF2rFgyu9Y4V6u9b0kbjOq7lbqasbF
XEBBK50OiXv3mhR5A2Vkj3x/41VZMLFCJtNOw0QwwSaVmBZAReC2HLTDs7D7UMn9
NGgI3qAT9OmLlrnKNd6T1rniQypigoBJXA/cya0ee4EA/5/2UbdiTdOb8QFdO3me
0uTQnTBfWLyPtRfcDqJ5kIBJw6cv5UBD+wMs0d+ugRxBUJvT6lqNY6rL233x/eXl
qETzPy3HM3PWXaR8HVqeINMikggc5xXgq5fclO3DAyMDXCOpRPM5fgyQimGhQF/l
D+ZlplhaCdf6yLfagW4vKGDMvNmHi/Ia6pyheT1B3npdyGXtWDzUQh2wMb2z3ANK
HqMx1SsqrhN9UuHvyD3QATM5Th9OIXEzbVkkmiSlkxVLFDGG2YOXHk3Jsca3UuCd
Q/YCv2asqVm4DQavPI0Jjc+LDp57tGH4KyTkIPpZzeQMxe2W2Y61zFe3f/Oq1Ci/
87Kt00rnROC0DBcvGWf6T06/YgiK5YVrE8LqdS/86qlzCGwv/4LcIY3lIVBphuXT
PVvgXu7CdZZ/le9OLUWIB0gLikuQp1QhTrsZZ1xoaMe3O0D4p/SaJxYqvKN9/ZSX
HhHVxuvfwCcl4I0M7VzyVW2YHTE7mlFGmxNcKC4FBb35kotZ199/wv62V8I6V/V+
10EcidTkgZliYFADhaEdce4GwsTuuzjCK+NoacnO7NzPmqMmZ9vcHeiw9JO2X5fk
zVO/jkOfoEh1znBNJKCrfCPH4j7Lk4+D0wG1gxqgHW/wRXrNmqjIMWB+y48S1Kqu
7+SRJ680D/v+PLv+kOLtJH2NXBzB6BHwzhnh6Zfuqa00dhgIyXu0uVJL3qaQdQtO
JlcCdJUH1Qm1J7JqVz0S/diI1CIw95JRYjjyw3M61ZJe/KTs1CfMavLgK2ozJqq3
6X08HXiXCVS6FwZOgNIDlYN8/bBASBTsLEnDuee3KIy8+/cfoElS5AgTjDBa3Hb9
1rGG3FA+SYHvmiR9KXN0Txn31ia6m6Otn4L1xnLG5dqH1I8CD/Eh03Fg3qTa1GjY
ipqNfyNwhSS7wWfUrkKpAyNjl63Wf/ekFyZ6P3wV7QuE6ODgCo9KCsuf6J//FKZd
A+/fZD06XayM3jziuE/bYI2zVxQDKGlEtkjdgFClZEF3B2MPHH1WZDt8vH0Iw5IP
+lDRHay1yTNR7NZYY2zxEl2Sd38bJhJm4LdHP/KLjVIWuctqdGhsQrYqqlski4gk
9jOdhpnLExBn7reM2nohTHPyBT++QpsUB9OTPlw9q3aTY4UhbnE4kK+2d1m4Xr/N
JzQ5WbUiA62a7DSbcLqLo6n+KLV62Ts61ni4aLAId/pv+e6YTIgGAKRqKJAlL5H4
MoZolsnSfDwtGCbPoOSjw9JYbXiO/ddf3L2vL/ue/WAtGxYyn2oQiqaG1ZvfCEeF
NX+5rnX7h8uavJMT1n9xp6foL2He2LrpQjaPMES2BUYj2XY482y15sRoktb0Zunv
v/smF+iYlZcxeQ3unh1sxF1f7zU+VCVJOhqDumRnuU3DNVdNHbAhO/RWMuu+iK29
gtt0ENvmUzThqAB+SU7eXPHzJnVY1b2mla6ALF1q+nfmxifD3hnw4/05yR8NtswP
BuZN0wsSNmR+NZMUSFBhnK4wUHZEXpAenWQaEK15TYCIWyo4ipSbsusSBY7WR1Ar
I3byZ1zKPyNW2X7Wzrbmo+h/BcCZvhhUU2og09T+zZzssDURlO6VxCmfM/EtkpMr
6JRQ/G+nAedPRm7Ttpljf6owl0DQEQy7cpm/xLvH3Bb4XKh5qxfca1A5pEyaO4R6
Cmb2cmEQmZFcryFtRAaCxKXLn0wTQygwQ6zsulyge69BxBtLL+xS9xHdV28lCeU3
nZlvxtSXWD1U7VPVOHyBDHuUPhU0GYOh4K8/n4iMMmcJffqbf0p0qRy9te+hGdBT
gxQP8xtt5HDfWo463dFmi/f7cq9eCzSwPPnp9M9X1vAb2evnxkJ6HMyyiffF8sxy
rbFsXXpGnF4siKG/mT6kaGSBZs99Ad08thKU37LB4vtGvCdbD+gsnfZ3mLupahZd
U2Vtjw7U7B0PrjXP/kB9UxJXRjjw4txj2zsfHjKAwT6VFzQlf3fh864EaxC97aK5
ufIP0bpXftyFjLVKGm/QjA/9BxqQL+fTwKjHMTOZ8lh7YiyvuurIuBdfUsD4bhMs
CpHSIqwMHYx6d88qwzj6nVsFX5DwpMzEoc0QpLPOCZDFd2XN8ptDD5wYUUEBe9+7
FnUUoNZfr2D4gMpAptl3BlywUg6W9JAQbWgMaYo+8T25FMXAFYLuhkEEKGYvn1a1
FqeZ2xordzXwo/V1oo0/SvtatDo9IaHeQn934NskMiBgP8B989gHev1/7eo5bpfU
x11+zz9USMakJhFxkP5bi1laTFkz0jqSdiZUmrfqJOQ53++T/OFMF88X5g9FNbEe
xn9P+M64cQRPXGg6GDnbnruS5L/OXx2kzOp3fCQG6eGq00/fWgWSbmEN9FkLuo1w
u46Tl62N1Di4ODS0jpMVllfEUyvCkTA1qi9wGmwGvaz9uUfSojMpZU3xmW1YXVzv
3H9dmphH7lDmsX4x5h88PEj7p0TJ2s0cBGZ/iFaMJDaDmVoN09L3FixZxtLO/hvj
cAWQXXr9mDpL5Gs9T2uJshUg6Z8yPo8iaFmbZeRyb78MZEFeBxTr/4Gttlj9NufJ
BRe/E5AEIynnrZBfWURdOZB2ODUKTn7Bo7osjV+2AZShN+SXk26aU0mZeJyyIW/1
blqHsbejHSZmOsAYIkSGo14sAalLGX0ahcdJ08G9SfxLbPjNW5aTj3Cpwe1BYqBa
+kg9Im0t2tkg34m36MtsEkwejPHj7MdGvRTBn/2mk7QceQ6QC/Jntk0dAGGSnEYW
wtIPsxNEV9CzXyo/4Jz0TygI2rr9hDuo6FRyGCxAmzKHREZkYlPsFU6BjcH/UWsY
qJhk3Mpfpobj39cRlg3/PTipNYGQBpyEP/YSGK6pWNRlDzIId+xMnA0PUB6ukhAj
6WHMIqAaN/FxJzJpYR6c8uVeEsQRgiW6V4h6pkN5Q+0zx0/BLdYCsvPCNBYSNanf
tjErI96lR+N3zY6BtskwsYUtBVeB/wR1vPn+Q1RtaQ+WbRd90/uDvuL5jCtDDARf
5poXKf2o1I9OM0O8df3vIj2MkewgnQUg//TtwLGgBYHI49ZdcC8NU8A51SseULAh
yfVT0crJToJPdmV3IxHY/XGnb5MkUW3T0QdTHaRrG9R4ZhX7re1qddmwWiJFx0Qp
zf61RJpoPk8111OLvjkHm1kY8M2aV5kfliur8oPcfN55Xt5b6lvTzNGyZCGUT4ls
HEH/YCP7p8O7BMxCSY/cKWGk7lfg6uy9BwjKRa37g+cO4KKoq2XM5U4q6d/cjXV3
bc4KNyOZKqr08becKqz44mm3sHYaSonsr+FENU7mns5bUbX08KT8VWPNBwWh7HKJ
ALQGvP0rvPibf5HCE+y4NptV9SY7/0d062ONiUtd6x5loVe7MLNzUFeKmU+4/rKj
oILANUIcCAJzTltoPWuSu6rFA5F1CWykQCg17Bdi8jWPIW+9oJ4IumiiXykfDJt1
bcVv2zxHlXE//WMzXH27ddqtenZOdCDzRSsII8lSswUumQYe9mtB8A2PAI88iuk1
cPWRiggTx3ZDejRr/qnE+npX3/U6AHNXjSGpXDn6SePtEhjNg+AFwQMZzKPxh+U0
K6aXZoxfXhnDwsyJgoyCfj63EwzKnQAPuj8YX7e0I7s/poTr5o/WXqqFVXoCyuGN
BhfDNtkbvBviXwRAeZfbOIMupF0zd5waffi/4C9JESavsQz/IX/+XrBf8TZm32Xb
hPgrSPtrJ23oE24VIKRGVX26iqi7h/KNilNyp/mtDocNnSFSeU9+r7F4eDKQEHib
MVZhVvm/wJUoFaxMS+pTG4JfQpCD5I59EStk2C5D5TIz9v7kxj9KpMTJ6Shixe7Z
FacITPt30nWNkIM8oxJg5hSr+BbxEXe733yD1aVYHeleDuZ1njrdZjwsPabGgF0D
ViRXl2+YwsJNxkve/S+63rwvqk+Vq+/pzexBZ49doy159rQksTDINn8MJZRYECqG
zgnywT6OR9WF0gU34rrTdezQfhgSzjuJvyEH3NBYQN5ZPFxQEhB1dA6ik0w8wux3
bnsWC52fNGfe+puNwLSG9CIeyU1P101RpRAAxqLuHRXAopzVYp16xXHvn4AK54rl
4jDP++RiYghZLmgxNJBitbeUrCtjQfYzdbSrIH0IHwD/iEn05Zp2JsQmuW8E1Ilp
glGSy1+22XdBinfZqpoAXP3FoMKpbADlYuw1EzZIcTYpu4128xZZ7L5LBueLlQLo
fFDQ4JB+IgMxr48EIXS3su/cshju40PWUZnc7aVHn3VKNNa6E0hYnzHggiWbQl/D
Cf96+ekcFxkZLft2Fn/+mY+za7AjDVUVEdUD/M9JMf7lDhBHYES5im/3ZejqnjPi
gIWPuBiwKoukrFEukM7iwEphaOZx9TJMinhfW1vDzdR3Z+e91dda//I+S5rvI0uW
uu3hbixdR7RP0K6q3RIFIlwzaVWIDz8CxiVqZa6YWrTpwaZJ98zh6pp4lAdQWaSY
spcZzeniOlKC5BQsiijQnF0NKyRojkKDwQt6xGz3K1FmHMpbUUT33s/+9w/bpS/Y
Cph/vGVMOEY9HmavoSLjUnZk3z97S0mK/CXmXUmrzT9v8z0pgNOB6flQS63/5kGE
C+ICl3KrnreYNV8Y+ZSquszmzpmQDzyabU67YxKulMrVUPUowpfTDXarbgGNu3Ie
NK0oJADlopWY4AIz3kioAqf82A1ZUEyx4DBW57h7DEEIIA4+VmsUcgknlTkmj/9k
cOOFyWGOWanZ6//LBq3LatSXaGkerKLhLt7QQ8fY/HkEuPEHfhtTCC/5611YSwUL
G06form0Lqf2aPFkK/DvKnyIfAzJMgSeTTp6y8TgTexWYym1GeUVuLs30Usg35cs
wwbchn9B6ahsY6eSjDYJs5iNM6W09CyM69htE3AFHlplkIs26mHlYAlpB6kA0uqs
ghLpkupze5XnllIY+u1Mh8RZLi1s0RDGkv/s/N9dqea0ewUJj9zvfsGcA1K30EVd
nZumzTdKsNTua+JnahHZOyylJ6FYB3OkS9WoQG1VxpCTZrBJE0lz7J+JgLNdV21k
ghcQ9YRVy8EknAU+Wqm1QCdd+D64Gam9uoBz3DZt7pkMKwevqriPx45Tp9wPQXZ8
Oz9S1xnyldXYtBfMtodarFdE/sNV1/21ooCtFMZ10hTZZg5cUsk59VAXoAGeDM1s
O7qJmDmCS+N5zOpiAvDgWSfLzmLWZRn3zrgdgdM12EeGF3fmsVXRmooRtuH10Et1
YelIUbsojJe1Er/1G10E46XG8dlj4eI8EcqeEe91r8kN/bmqmCAv/pCx9FSgr0e2
UuBGHDD511PYPub6b0Gan/ySPrha1Kju91xr3b0sXo/KwugB9h/hAkac/x0jsb9l
hQFS0efOZZCpSPDGddqttYIYcAaVZTS5/DMNo9T2ymRihM8taceMTpEwuonVmdYn
QZ8gBGZwYGCqdgGyqm0Lqeovi4cv4ktPoqKdN+MI9I2LK6l9myTrOGUwibU+SROB
6dUgv9amha+jPQW0BG0VgaCFtKnZo+YjfhFPGTweH6Bloa0vGyBWOkAJpFONdS19
j8uL0G0hw7BkTTLuNWlE+NN7tEWiJYbFRz3dbMksfYl5fTzqebNMb6juqL6jBGGY
/vjpXT8Lhdu3AdI+cbQ6UlphQkM9KjaQnFrCMPq3eZC655KzSpZ3VAMR2V2PA5wI
RsgEIA+9IcNpnWQ1PTpBr7AQMQProKh16fZ2yoqnip4/peSxiiUbknIO9bzGlD4E
NcFjVr5xmUptUZD+Qf7QjwRMLaPVawYp6BFFIU2NpROUAyzEMD1R4NBmLZVkCCxz
x2rM5tmDxLbU1pFOt5/pAf049LDjMMmaj8r4es2nSdtKfJy07/sXpqaoWtIU4BLN
oheNedYSfhMRxBSQOynUAedY2F41viTEuCbbXwUUm6E8LIDX3Fe8j3wQuT4z753K
Ot4vSTpczxt4N4gcoqegWDUEwkf6TsaUWCSiLsoRSJj/KgcmNGOcP6ielLYv0ua4
D0H4B92Fhmw0F2WYSXeAXg33PzL2la4NU96v+kwWQ/qFSKdB+62E30U3nc+XaI/P
yxOWUOsM4GGq+eZntruyXgZRRIZj+uHv4TlYuJ6hz3oiKYgLX4/3HiyGaJDYtn0p
wX+hlOkvtZRJpySM8V0/dWpR4rPWgkTfzzyQgVGLKLLSPMSnoH6fIXsUx6ZxPvb5
Hsm84k2oRJe3vYBmoGYfPix4Uo+G3VOHSGmhMRSkD3SzhAm7mgCW6X2tRgY3Vs+D
AgHk5n8N3oRxtkOWjRZz1SB6GXX3ad38F6GivamDqZuZyAObn7X9YrUy1owU+3nT
e65JZqf+pPLcf35w9xXYwNic6uff9fwLTDtu7kcFQZzLnwnIJPzmVh0tmKWffqZw
Y/fm1ePwabdqLCNuhd4egngiqw4apquqY0wWowTn3LraoQFHy2vFbsKcV5fGQqGu
ioa8oY9I9qviffc0hxzodIUInP2OUsOsTXt8yEKbdAX7QWf8NIYxRTdQ7qKWD3aN
wVnCAEuIoMPj5QrdHlnw41c/Zo5N8NE36wW3ch7AyNm/jm77nRfC7mTlK4cXLCIy
j+pTZR3lIYY4Dlj4iDQ5ZyujGkhOCkGVm1twQ3gSW9VQnozZnBcXzTw2Lal5dLHj
kl80gTt3A+Jy3QrbPpuZL+A83vcqc1Cvvqyc7uZvLWVETIsLYjeyVAH6MGUiZ7hh
yEmJeEumk3C3g3eotcrjCQgDKwhQ8GULJhMYoLdqu51U6YLFSGzdTGgh7KmQDqU/
mMcfZZMo8CBg1pUeTiVqEABFA9jLAUjNVyA7dzOTvFDmUAdrw6SQhQCrAHzvr+yU
jFtBdvNfnt/nzoYFXkKdMVl1goZWHZxUt6ZgPD2yX9V7hYMbUKI0EyJyM3tu4YUK
9H/zyxNlDPOPPKDMtYEVqOVRMinQgJ6CKPJrBvtca2S/+Csfa26BdBax4w0i39Sf
F9axjGmZ9NX/4GClJ4NK42OlIBtvsaNjOEa6iBMklx/PO9hdHBAPICeo3AEhl9JC
L6ZWWo2Sa5251FtYQY1E6ZkXxGN1ME8F1P2VOC47Me7TP8w9AN/ijdpRK6TU9ZtJ
ZSSI+vtkkJtSoP341VB5SCWwch1chnO97Um6dHaBXKyUfQzzJUWs/E4Mi4BZ3t4o
3VTDX2mlhxsMuQer8egxBHG7yvwF+dII3M2d65BPewHQp1Nrevzx4lsagxcvp/T0
iAlomUIdR6xT8XEmFQRUsDnCbSNckUeYAHDvpJ+2ru5pQpjCNmf/wH5XidCP5pDv
E8kNCH5/sqUj39zy20Lww498kK6ZHRKLY12R3vtayc0QeqttrvYilmsmjxHovx11
by7bFSgwDOIYb68gJDdxWMz5c8DlzOV5aZrd+akWCGOXdapIQGwpfidYph5wIWF5
Ls/fwnha68gvjaIHhxhGMQVTl8b1RuBvrn7EfFYTfJqL2FCc1MM0dgCXDtj3yfvf
UL/v69r6wpvk09yvZN0bZjH+T0umaQtzHbHFzkFockPg8P5pmxz44EXwGMQyg5P0
ngTDFaxLQSs8wyfubJQkTsbLak1wSbBmEd8keqy5B+fi2Fo1m0BDP9E6XpWOhSQJ
xklkF8RPTBmLC7kYp+43e89y4+1cVkItgbGsDwl5rg6eSepX7j/7JFIvI2pV0Qwz
xMX3c9EUjYCXqunnSYAba3UBVb+Qxfvyusp9OKYz6vSG2cX/sC8/PXDMDzJI5PIg
NBQ/Fpc8ZteBj0nCcfvYjlRmX/4OEYMpmXhtehL8LX3GLaghOJHWg/hFitGCxh1O
gCaEK7x/mqILbs8SNONzxaH4aNNOo/TmRVYevbm29xeMrROln5dmQw3K9psmKvTB
65REaBANlN/LrC23EkgnW/YyjEx1s3syAvln9RH2mmnJimdh4J4mNuwwnLhWHqAZ
HS+0YB9sxskBWWedwXQ1/8DP8qd4JM3za6RC7sWMBVGy+T+CfO9XXFBFohZh56ex
VjZ9IgPK60MExF5JRmN98gfUpdUmbYRUgc37Zhzjb7CJRXJpFBhgxH+qeb0cw/7C
UYsGtHk18EQSfZiDDbxasuUZnkr2emcnZE1xN6SKLgnW5haQqaFZ1JHnXeNeY8rD
OLiwXiBo5Zv1EFutA+Kcf8RdVNtNJH0l+MYBjJMK19DcMwMeFx2bgcq0RiRxvmHW
VHJYf4Gg59vxDoTvmNWMW7SmmHMYctmi6E/U44D6PJmF8ZS4oZidlVHf9h2KD6rV
hXc/3uMRTZtiv38gwm6sGUNTqUscZufQKgPrM573FiE7guDBZxKM1h3iIbqVk/nW
uPQeCKH5nFTreRW6D6DGrGGrdx8WWrm4ZiiIT3pbItMieQ0M3YnCCzXTGY5trwxh
1b0FO7pM+qRuTzR/jg0sBI4KXL1Y4AmsGBk5M24msjgCX/CCcegb7ulahTIAz+8T
jRkhxTPiqSv/cLHLUptz8Xadlb4LpCuomXzRWUZP6jE6+t9aB6ocsbvQQ0eEH8TH
K/v1LgyEl7ZH8hwea1MvWN053F2GUwxB7b56XgLUIOJ7H/0YqlISg/R0oXEaabYK
fQu5mjMRhi5g4bGyOp7F+FumRsaSVdfEWlKNbcj6izqxADR4Bx3TZZSAa6gZ3kBh
5BhAl85gxjK0IA7PGjZbB7ifyVeGrU3wUUPi+yw+d+TaC4ggVZZBH4MCXCU/DLtW
w365LBEuHEbAiIxaItiVbVxc7v608x7ozjrnqpAc6jvYM3sE6KR3/h4lCw/IWIcj
iZbvX9c2lcoAoK9ZwMut16ZPcAFclJ0T5k1Zi9zgaeg0ZBJQXgG5GSlHDdJmlX7s
ReVP+ie0EJ0PzbDQ2zUETLeaD785ZtkQ+TJq0gGzgjQbkVZ1v1WxrfOaZHx2tBNS
Xwr8sKiTGX9sqkSYvyPQPRaxuyrV4uWcg18GoTFKvGyAF1x3ykl2PmqnpyRsYjqP
j//QHH04StV318V6c+ShiySMaSuDuyHvjPOSR2+WzsA48joWn6EyP/5gHT5sTOIi
uAdXZzzZYocZH7CzYABEzefqjJAyJTiNgAVrurxt6c6tBc2vEsaWTADCfQJ4WcT/
3aJ14a0O5Rws37o8HCDybtLYIHwmApIR9G/Xvi2OV52zVMbYVNssrJRF6QKxObXQ
744/lOL1ec06HuVCZ41ChFBnnGsXAnY3orDSnikx41HvShDLS1hq5YXXW66lFcvd
X0BIzn7IzEWv1Cyib9qkLD06WfVjadb0QIqBNXXrDMuTGSBYboqF1v91SWLhxie8
VGbZIsX7N89yKzwbh/ImwujXIYP2JmL56xuxblrE1yEBZk9t36aXILJce8NjhNQh
F6bB0aIPfiH3VTrXN8wSy9+BoY3VgtUBrPCelC0m/HWtz/dpcvrKbDFs2kwPpJz9
Jph3Ek79rJJzE/D3XGfZDutIe332UGBfY581a62qh/6l8qfuowquT7TOZ21Mq3CD
O6b3H0FalRdfpMFIBALOCIicwW21Q/hQTsfm3jve/KdP2jRfLAd4x2GI5PI4ps81
c6W/oRuDsDbdjBuHiSDmcYfUnHz0PZAA7dPfUvYv7fdCup0CXY7KtjJkqMhmWBi2
meREZVzq4A2wk2Bo6rH9yM80R8bul84Zcur/icJW7ryXuc9PrlQIpeRBhjlFpIMU
kICZhFK8BW0ZsTgOgcX+1okEshZAKVZ9qHXb8oj2Jh44Ga9XxNQ+LPMXaNr1ZxSI
ewDybvKRK/U5j0XJQPuDfzR7BOC7huXlSeKFwBnQgsUTLkPq0Kap0si2UqNza7LL
9o6E2LcsanmLfp1hpaAgDvMTTLbHrpn5cl2byxAnAUT6J+cT8Qxa1Z+y2wPYNVn0
IyIgQhX9gihyAIrrJ8cyXIB5djalPzfbQMIDvYFXyMPh51kYWFqCxKwtyfOaGdVE
us77R5X4k1UltsDZ1tlBjQiJHIaLfc8iQ2TBnN8bRUGKKTTlI8VVyklFv2LWX+Tj
2nP0UHVivJuT89WdGTvpXFCrFPyF2B9fHV+u1ecx7N1WziMLOnwGrhvvVGTbeptn
XuF7tFDN1PoJka2KRSw+NxRi22vY1dyY6GH3zC5SESqRocAo1bslUk33qiUs1k9g
WRT6s41nJtsKbyGw70q0xvPZMuU/2aP2cysiHMfw4LYK9wGL5OTA8h7VqseAJDjw
v+w9QeoB6J587XOqidE+Kno88Acq49tvzayWVeRycqnteJJaVfxP6FOo1QRUW938
p3WX5gJjauycSaUduOzIkSkMrBimqIqvwBBoXfllGwhxulGdAhq8VFgz1n8lCG2l
ELmGaa+cPXuvHK/j0kYJiwfYX+C8xbK6hZpmOVj+8syO0bBQ20v5vkwLZDqztq2L
YPlYzYeQ3QoFRapD3lgtOVtcgE5sXcYXto+AaugYgtXFiHP4OZhqnQfGnrncybCM
PrBTdr/pgOxFhNFhaAAXmCK5Q5xCRKNakKLYRPGnuYCHgtIi3NcoXEZH3hPR1HQc
2uFIMxEG1u0R5He17/uIZTMl5dvzXjLC4s5bZ1awpsdm9K1HbZHPcFHp/JLJ8NR+
BUDaeZL9F5JwtA/M8uwzR8NVI6XoXcLCdSi4qN42d67ZmVMpxiMk4J07U3KHYvVq
WHaYqM4JD5eRAmRpaCIhT1G9XANYhdAsyfoBzpXPDybId7DBKtoN/272YWVi+9U3
aDKNFdI0u6j9C4nKlOPZX3cgq03M6Fv1XUMgPvbZXldO+gdniiU7CvFQctUce339
4mnDfEGWXjUFbtSRNVQ/SRTNnODWdLDeq6ZblcLUwWncqndh6puudhCoYpJBqlw4
7nL8YaTo2PRu7EeT6kpNxArS1droAEPfdYBpKFgzvRvtYzmDY5ARd+tyNal7EI/F
9ciR271UrWTNtgF+LG4kpGtv7xsVdKYGaBY15ICZ1vzrSDvPOcUNbv62SefZFhS6
NGj++D+0S2gKEXgxBKU8V/RIS0FB4nrSuuGtaKez39BczfD0bqoTxpEZXulRiEtp
CtiJwmNXXmMIGE4fKJKA0xU4oeZYvr+vwi6732PI58Kgscrz+y1QzRa0i3ZSNmUj
V0fyoDvOuP4x42yveE0MR6lP0QRt/gfR6QyHtjt2lE1FD2F76sDlsRN6dl0FOoDm
nxf2bTzFL63Z2u1Z6GuKoSSVlZ6bQwAgvUqJZFqPTerza1QD+Neoq3tI0GKaDfkc
PvEZmBRnfdRZ1OHPVpWuNI001bjUwGa48NDKz+S6xykDJ/Wv/FgnG6QYGY4+aqyN
QPiF9vNNBwLW4Abx5pqr8iYZ2/6Ocz0ogS84KxnFAKSZ5/6kZ8wnU8/V2a2UUkWa
RniOvibf6kgOLXp44CuvxUht/4QQXUzv4m0vBJ+T9d47m7bysLfl4Mn8c9V//0dW
KQyQjHs+WKXx0MEgH+/3kiSDRt/ss3g5V52/Ckd1o1i4uVKOYQ78Fi9zha6/AY/q
IIozm+R9lp+1GAeGGzF3H6P3GguTVju++AYIZSJXQHv0YWri20SJtsKWePmigv1e
Z/cCNSXqFFnX/rWReACigaP8ASbksxzUosO3wZIBwzxAQZ8/mXweyvv8zV/YHXKL
zU6Bhpw3hu1FbzpaLo8oUMvO0+8WwRncdsN3gPZPAv/FeEeUk61zkK7W2bY2EjqV
g5neN4UKUPzq8532yLu9KdHIE9v22c4Ak51g3SNd3UApq+Dc60rgiFP1QQaZzrxJ
DGmY098P5Ti+x5/XktkhO2clpbQtPHU43/zUGcReeDGKP1rEaOGMNZLH8EhhUM3G
ZG2mhrVOWNZVH84lyZA1Hd9FL4R7Q2/LwQgAb9hA6OSErAQPKgC7ZM3iD7xjtO1P
23wGApW1D5b3g/zECdyLLtlaU9aPLscCIe81ae1J+kAb0/vjaqsvSXWchQCiYuGp
7mPCZSDv87Yq12oaGtTmF89C5MNVptfB2WpkmSvAuBAf8gHgdWoIRgfms0LIQLik
cK1AkMfGK+QaSsSK9owBRoFpuBdOlZ2khZT3jJ6vfVDn+EfMamTkHHQBM+V4emmF
ZVuYo+DvYtd9w3BZslGtLU+YaC5SqsxM39UZEpg3j/vwkzWFKh2kr6oyqir61OxL
nfQxfaRvtIPJgVE9Oxwoip4XXfOPCfvHOW68MUkkv/VLhv0OC473K+zujmyBtrrG
CKi4Iroj0MO5tgWKXvl6li2m/YhRBPnH/FFCUO6YDDh5+3ylhWoKCMr8DFLlorMR
pbHIstAcJ4PuHeVPLQcVA88a0jFQh7czTZoiBbHVrQiEHVUvSTRNkGlfyXSNaUO8
g3Vrc1xLImcr+OkDPVf+b39xwPGlY3y/YVjeBqPAJBkm1dRexUGBValKp1HdX2zU
yY2CsC2gSY6n2eAd9sZd2hJGf0xdUB5rAxfiO/2s72IQMsN9zZMc8pWqhacq/mTE
/6EFlg/jZRKeN+/EgM9Wji7PrHCAWGVYlSsmKYkg+GCEFa0Q5FCDT1xeEKU3ONq0
J4aRPSAMJ9VwvTPFYoSiLFSAaal8vy8hB6GacZnOr9zF7A2o/8TRxPGzEysMIz/N
NfTux8K7U0hO7z12rpmyoqEyqyxJozgnihpNlCZ9e14eVVXpTZHHoeyeHdzzP+p2
pJG7llxccVsWvQEqiF47qpzMqu9cmB3OYc+kFL5a9zFoekG8A2D/GPbvF5bV5kuD
pSaXofp1SWtbtefmoEvN8zo18WcoIFB8FWDAftsJUPviOVXQ4ucbW/+IcWBA8eYB
0xxR7oExyuYJukeCshB8LFpjzROlNYfFW0Mrt2p2h5UGaZxz4wjVuJynQaSqN6Q9
38kF76J3Dj4oy2Jpyff5PUocXgWRucNZ/vf1mU9P907My0pvT2sKxW13zMNY4R+O
PCOXQO6KewbKsJw0WtuCJbXTyTaWEU5IDWWaIjZH469IerdW1T7vM6MqVWqnmsd0
PlMgIJJ6NNOuvm7yV2nxAnNU+2/HM042hngjfgYlrcB4XuWh4XNBYHI++WyugTB6
X/RBDf8zMqVCaW1OqLsckKf3Zp5yxOpY7h0CYVTCNmqIJPLsOXqtamIn2eZ48bbu
KJWjyRE+6IiTkioFOQ8vBQUxdlYsZpQuU3xB7U6/IxbvXO87IqlIjeL17Fz0PkMW
Xk2q8d4glKZ5uIfWIOVL3PPddt4Nkhf+eV0E3nVtV4eomhm3yTNA/MttL8jsBdhp
CXf3VN8sJXKCqU9VPyt4KasEAdUQQ/mUo6qPNnfeQYg/5pIRuVfWopbR5MGaJZRh
WhdeuSHF5TvrpMniDt+S1OqV4vvN9HezfCW8jX4C33sOZWM6TjXF+by0oaH+xmSl
EFoEZt3TU2MercoMa+GCSzyHWT302WNInNoS8fmRceRQzf5V/SuuON65059NgHp9
bo9PVqBm5PL6XlDFVvK8Qs4P8MC/lU1dxfcrzpNAb3GMluQ8oeRa5TIC3RIWtkrt
bYP1Gj7kVNp7JY+RFqR0AMLI2/LtWB1bXXAqj56uUzOzCHhuBOrIL09/nhktqAZC
0ERII6N49VyuBeYc1g0iD+uQJpDy4lclAhCaFdQt3tHpBHJazwQ4/Xx8ShtTCkZ5
maTDU8kVEOJRcLY+3QxP/wB4Kvu5QxbMJXTKKRnvhfomIaBx6sxTyubuzOh9i4ff
vP1Vqn4hwp8CsD/3KCxzT7tmo/2A+6hRayhFwYcUTIQs6/+kCEc1Frg1W9QhZxKS
bHXvUUoE3O1vrMW1hZQqepRNvP4FQqWpNu0Bd1fiAbGHQUF3wnb1KyQT8FFH71yy
Sq/S7WuWOZ1P5nx8FLsnGXt8zimB+1eua7GL+SvH0ihxfIlPkjbWnlX9IRgGTW4K
0NMs8C0XXlaAEy5T0TJQZP2xhYRzvvZgqsW+CVfTfQfX3TwKa81tlsIMm4eH6rTv
ZDU1/UnNdIVIIuADW1lii/f8fY1gi4ytn3hThciXY6A67i0JUcko0aFNk/0dTtJi
zi7qI2E+Jp/L3aNkYxMhENcy8dB3P1BJXVqp9Ki0RgAvcsyTkppXicrIaYl34ofV
jBdS9BXFl1oeV92TAfNI9RIOt0S08Bo+iQEoDzEGjUP+puBe76dEpYQXPHGslL41
Vxn6jJc/agipUzihnW0zMJh909xPNLa+i5Wz8PPsxjiEXnsQQjl3fooHMnJivwkd
QpBYYziWaZZ06BUmq3yv8xnVE1iFOmPq9Qo9ycQfU+Zl2o0eDBTYyZciyMS3aKlp
w9G1xRz2HVI85j2uLRAFosdPyN1WLcYgBoNc1M7ATGhQTFLsICdoEtkqJb4Pjuha
tILEY4AJrVHPDpCJsBOOpnBxhPOUr1cEKWFhJL2X/q9sNyUCySfti3Zf4tJG/X/9
yQ9F+awbTvOFvdKm3oaL9bp94zx/kC2tmazMYGQ6JS8A5Aw+Wjrdv21slRq/g+Ch
GI4F48X8UUapfBWf/G3cAMrJ3IoPjtmj1ds43407GjD6ZkIHr4CDDHaVwaWuTodD
o03E6Qwn9Zd8a7EpOKVkoW+iqLWbMuUeIyOd2TKlu6SZvvsCFgnxQJQ8StCn8LfJ
p5X4boHuqufob9LwR94Yg3Pn9TLvfd8IlwiQQASPbp44NOMf2c/8cqDyZolk9/hx
qtvmBI4J9ztdE4K97tSNH02pxXd+obW4ycn3U66Q7OBGqoCgdGz5sovSOnWfKsYq
kZRJrwbb/PmYPM7FA8qE8UnR5hFIeW1TA7uLp0oH69g6mKUuydc41OPCcslBV8cc
Tnz0DAp/5yEsDuWDbpzdrpdl6C1KutxGAwBXe3Gk4ozU2OXbZ8dRhxe3qN/KDHSb
BNJJmSOgQ+tgZc3hYQQDXjaQSVwgYC7Xogv8EfDtrHkCYApzLq+NQzfl9C2ZEfF8
siJvK8WBRiCr4Z6JUlkxsEKGWpyL7Yr4byft4IjUuYTmZCP2dTA0jaXqILYc5AwN
fu6VT/vpXuOvTUcSgTnz3tjTEboH+n+CyxgfBh0RWN5wn3HRmjSdYT8BKmmmW8+V
opIje3MW9hHWfbN/BW1rq6JBDK3hbPVVx4c47DDJe+6O+LtzxmKeSQmodE6y64lP
wWacXG1FEzIw/0fYOZBKXoX8coEvtTff3QzNp50WqyyyIOxvs1gxq2m8cTcA5OOF
lBfhILx1iHjsiq7h//427FkBV/pcofRH9N85VfQ8tZ0NgMBDZ1RN67ywF1jJBNiY
g1DzFp8pAQvhdF4/4FKWjPZd2VS/o8ATv7+/qBojEiHU8sWN38jVZuZhAv1zx444
4gSHZZDenmGNBsp2MMR0rV0q3ParkUZfZJ60LzN1i97T06KYFUNrt1+/Je9lKWoi
Qjt1bPhuV/Hphqx1fZ8dScXp95iJqkr1lFPwqZT26FNdKRd5IEo7X3Ia8V7yOXZh
Q79v3s7XwRgMqXOobrsuMqu6cMPV2+Fsov6TlG+Zqsv1JgaqlKoyzBJaq5qV/Fbz
98/otf2NJKy95ooBirquiALOOVakZU+tgIh8rzhH9YkvcZ510cSv5SRFDn+QQ2yn
bIsyqnmQ4v4LvvaU8hxdF4wMcy2NynDmjs6TX7UJ7qawsOa14gOP9oa8aoeBWv8s
NCpURGOV2OeepBNW401h7Tubm58XWjPs/OYraTBu9WF15eNP3MrAAmBFCkw26q56
18vRPfQyK0nLl15OYFRbo/1z0eS5UikuCB385ICOa7E+oP277xKAGd2mozCvBmjb
W7pVJtiU3n/3RIED7WWCJgj6TJ13b5iXlL7rxqS6JBMqAXeuDRb5MxLil9aqhsE1
WywGYrmDyxdtrlPiX7OIJ8ipnYW1VzRbYjZaylItE6lnR1tIREWAhulLmVoBuDdC
AG4pHjS528UwBG2sB9R3n23HJ5VuTdkwhlffj30BQl1qvLLyoySMRjdgjeroVjHp
McciqtP/65kja7ZXZqgXfbG8uzXliEmt3UkcfWYfZfT2Jwke6PAHGUwiKybUDNrf
ZaEefjbQ1MWgJCqFCNoPXmU+Jl0P2QfoQvO0aP3mTycl112wYjDQxMrJ4btKyUQG
6Sxah4dFiztVzGroyQkAMhdkUkh0vzdlDw8XhFCM7FtO4xnA+5cNRkj9jU4OxjaQ
Us3OPsqeVyRTwzLZgbmjAlB65XnGvp4WCi+i3CA/QMtiJc7Pr3nUac/qadV0S2bs
Kba5P/OPbQ7qbczRW//f47jS1DxhwKVLs1TNwbqt4MLmZ6cTgRy97BPfwE5uf/s0
mC+4ZiBLyj954zfIVxknxVyZe9jG1LufN6Vl/gjFK2bYZ/HSbJsHEDEIcrIBV+Qn
jjhqUyQ6Kh92ejqZXPkX/Z1y53k043Uq2AHljtgPTYe16wol9YTPLd6gtBkYgKHv
Iuv/7MiB+oZwUtmJS0sYZw2Ov0+SbeeeR0QJZcpkt3qbT0EZ8MoccTMQKEXk5iZh
aeR9J0GFi0CNI3Tk55KiBImWAnlbHFBW5ZsugFzJ1wujeJfn47xEIuXwwK0wcBhU
6AtjG1cpQbjCwFX2PcnTkL5Je2ULgBMN/MjnB8zkQpXp3hEpBQNFTWF/nB7tydQd
DLSNPCmFeWd5eRxsdbWjp9Uvu2iE32JX/kHq0h9nNsTNjbW5zglC2MBnvMeynaJA
Wyia5E14vRfgzlkFBMxImq2ToHIOPffEBNrID8tM4fJzc+by4yCZoQZ8K/70WSgX
TzdU8pCzfBJNAImXXkP54BbwULjCFfoT60QZEkas1bG5PP5E+JCfQYTqNd9bI52z
p8yp2uTFZh1pal/4zrVQmh74DK9PdReZvpvgGwkZeTs6oM9eNdG9M29hHKrbvq1d
QJuRW5eUHTq/Ceu4JOEM4kPrVYSMpuoFzwbSaFsNJ2NF4GwBLSvO0+1cdgBQSctO
AuQJ5AjMykxMcOsuNeNhOsXrwahH35ZyBlt7l/bjXSWuue+bPnlgx/KP8cFvVwAA
IJ05B6vc7tz1wKpNlYcNwzAcOskKekhoOJwUJFoe4R+W96sY0s8tiuN0CUfdMBcx
5y5rsgNt55taGjF5Q0iRJvhsO/FcjJu4tN5nS4JZmBwTXNqOwYPOhs8ThxTMDM85
P7yK3cOffwZnddHMW4o0MXwFB6P8loxhxd5nEQnbHzO17GwZz/STagHIao3Qnjnm
bDM6C9/nWpphng2wPR84/ww7eOWhnrLdTZ+DSJZDonCTkHEGUpxAneLa3kqhMoPR
xj55iid/YXLFg6O9miCxVzH0nxUXjCeCOW/TLHeTKbpxnJk8wQW97TpS3cSvqf/Z
dECl8ND/K1R1xqjly2Jbp57uhCt1C5FhousE12U6YnmMsZWvmJV8UWkMUQr9TPc9
cGbqyKuBD6xmXtAKmSObfTwyrvZj3x1j8tbTLGE3YjEcok4nyOCpL4BDZQCwBI8Z
pMc6c4HVVR1zYNDaFuVU5Jk7hu85dn8hPd3hOGqr7gI+MSpASaJmsLhbtdM1+hfZ
e0ZSWX4L2rERWF7IhvkNxXtORORDzT31RTLKERAt52Uje6ZnOR7/Kxh3imJ9wMzI
U0JT9S86/NSNwAOhh9s/njZZRjALmkFI3qVbNr1btFB0c2B197Y7coSxhS/gHoXR
M94RtPlMWE0TOCBDEvr/UMkNW6jCGhNqX8SqZSTcCKOn9zKUYMFQHEsVN8Yh5gD8
W0LlnXnYEetj0W2LKY4flda4NaKTlNiCANKgadAyPB7VFiTisqmHSz7Eodx7UgL1
UMn/lj/5XjjnqG7+ZqUfET+eZ/hc8mLkw/EZnLJNhwpxOrKt1SN/ewQ9JDhe4l78
RWAX4oV+KQMxaPWMUxw9VSp3PXK9D4ISMKKggecucvy74spXiu6egFPKEl97JBJZ
laO+aJalEnfgGwNmZkfJo1GTdZWtdi+qAcGb9MShzXIJN3nTaXJHZ/Bh4NJJkvly
aikDTACAzT43ojBlVCHu7MO6Hcc2etyaPL8Uu3QT098MWVFnvvThgsYtAzKFtb+9
XdC9uQUmxWE05BApFEzkGf28+BKyWO4Mj78Ct/SXrsGY9wtFgU/aCLNZ//RSlu8r
1Hk3FxKh8pT7PnNrlwHEU0cy3PfaiR3NZcowu04C0Y0mz+OiJn2dzoyujHqif1vS
65shmI1+wS/mXL7lOS+N25eu3Hjserg7ifdumWMQ34tTRLv9BIfCvVZ+Mpi/oh+4
y/b3yyKSjlr4pQ9a7OT9x7ydDbwYzxj71XRkGKMZkkIcUGxyCsm7IkHGHnIHMc24
WLX+5EMyJWCwNG6eozLWQpvZMj1QtyQ+r1CdKUf6oPqCg0WHrdPJe1whO6ufFv2w
j/rcChodCxhBsLVV35RIabEXI7AwziVbRiesotPywR+aZnYQxlb6zXpnil8p3jFf
rK/1zh4G3CmjbWabdL5aKW79xr8VDFscDI2obA7SEjJH+baEkCzx3UhAw2PHDwtq
7v8Ntcm/zQg9IdT0kpXpCrYw00nHUh19Z/WRJ5VmqCeqFHFMZMYkV8qQhA/n+MhP
QyEDM7JZ45WRtUeSYFwxyAEHrGsTzPjd2pAAOSs9UYIforMuPZtdIovvG+cjcOIn
fF3ZNWnb5MzNQa2zDg0BY6pC/TDfNs5rg1G/e/Tr1uaYgK6qHulR+tDuiYMi6puz
JLsdeEIOf0HArHzDYm3yLhnvsxR7Gzj4UTKgKT1XIB0ql48kAuzd2yVUJp+58p5d
B33bjIhrT1BmgKdwSuza3GLOLZ05NafYIdKW6GYfbcCbqvjsUUKzGyAbHsf9KJTD
q3RMBdojVQMlz8mlIIEcODX0h/4depnWtL+Ko8VmiSjIXpZNH8e48hBMH+R/VPOf
Mhnn/qpqRN0Ev4igFryVrkANzTJUZFfHUkKIPk2buBT1hlncrsxJzM1c00skZC9O
dEWOeARMjzRIwP9gFeyWMgO1vfQezEr/PogXnITtKU3HqCwza3daccGhTJ0IW6mr
EWNeZjQwfrtAgIsBkmPiEJdnwZGIjcz3/j1nkybkjmPV6UAaj+PtCZOL8MYuoxg0
wj/wnAESFvxJuPhpTaWQT0PX+tnu4aUPxq/lorSZ2H70Rk99a2YHB6jMkHZHEnrs
S9sQYkohi0bqGONu/eGjpR6GXC/S79V1DguqD/6vCjfC9WQ38Z2Td6F8gAWBShyc
+KC2RIk0uA0WT3THKUHKJIhhGiEN+w5lpC/OsRtGn9MhZMRStyobLreiGqgD0QUf
L0tNUTpBcnZuJ1A1nonYEVPglt/NSLq9tXDOZ0rUPvNQIj9UUS4roIrVuIsaOrQg
L806YQvkD1uyo2Vg5xYNAhkpvv2Ga6IQrQwAdhtF7Tfso+vRiWWpcW/Unl1mUI33
KeQapPDKbUEjbo4606KlZf5eD4EOxcTdajiF98TyLRVTDxRHfiId2VJ/5+Da8J73
035f4evfA36KIXfWCVewN+X41qyBqktnrXfe+951GS2JIOpjaDbPcsWFmYkutu0y
G/i1ebkuGAHf2ykg5WlYJ6jn3RPmIu4t58o5VftpjWvMBX89l4YpTuXCTUKg9zE4
gUXHIR0jdtcMyY9IilKOogF0JaD/XKHlEm1M0Uz/HuakwBMRLF/lX3pBkBRrd1Cn
Qk385tPd/frdpVWZK1zlIZlVPR6BIByW6X0DD4Ca1YlQYkNdliqmlpqTHAgTfCcy
wemk9XoE9d8bu4WZ3jUqtCEu5kudwbHXmE/yCfjhMDvCgIC5SaW/YRodFwwNX2tM
WtuGsZkobZ5EWKvpiWt4b80F7xkLhXeEGSDTZtnEGgZiWM2XYUM1Q5hd//o2cTwZ
dPZxs+/qINt3VWstQQLODUWQkzieVGVHhP4P1337FBG1jCJ3HRN8FRltYPLdX6s9
BhQQVjJnAIGoL+7m1/NuEGqv8iW8qBD2qggPff7GLpQCkpIp1PLOR/xBAgj47Ks7
FrKbAvKhvS3CyDjsYcwKIcJUgplFD5HPC0xqmTuKF1iUZbx1pLhDBT3ohrV3BEWA
ryIjnk7fISnSHtr737DYM6CEOhr6/54Nnd8sknYdakthZmLigcoT/jfE7Q7+dQ+9
5Ng/KKiKdt1n4LWjlmpOeSYGutIAFu+Jlz0hgip1CUOSarDxycBk861EXza3ClS1
GzFCeApq9nCTNyM568x40EuibPlnEjBp47qj3+WVx0HrYO9GjxA6Rh3A07CVQAy2
Gb9JnyT2fSw0suLfXdcOokW9lMuOHLNOp6vqm2ZVbFJCTT6AMr2O3C9nUfyUGFG+
dPpXJJVb4RO3C8BPAoRzu1FXId5AwegnzJ5bweUVm9Q3AmdBVQNjN/pmzi21JMNB
OL4AUtNKTROG85CIrseBxRof51BDqZJI6t5cbwWk77secq7oPXG7tEnbxL3oJ+MW
Xawqn8He+b+KK7qjo4c4I5vI2lUfwJQhvx6e6uTxEFdxQV46V1u9BRMBHtQHxsF0
KhA0R6ObgtEhGmSn8Wf058k7Xv78CXoz2x0aoGXWmryEzpOpkx4ziHZ6KZO9kYkg
aL1/03HQJPQNQvucMueeAkdrOToRNtLgNStoI/UL6p+b8WP+GOhar77TckkDIRNH
vgG9C6Jvp6BNTyG3Ft6QPybqxNe41FURUfwGIfnYnaOnhp05/7G7whUMJXjQLUDJ
gyOITMp0m+Vr/eZUKT9Q8dm2H9xcg4h17qwcrX4kZMEqdD21IdZWvVbTfqTxJ6eh
gckN8hXuArFWg66kQ8jPwCEYwDu4/qQNlfo8rL1rep4YbjHBvoyJcVPYx0lu01GX
37jCX08en8DmD9fhugzyODFCYR5sUSHaRAu5b+eoNaroT+iOyov8npobfN4pn4ic
oA3kM9yLSAeOg0telQgsM17NfMLSVgCDUaecUXiBMExYz8cm81rSuVgzhWVlsLsH
EHGQbCr2XztwNNayr8dyPdmEDtyQzdAzhaoGoRdANYlMJPWBtKWRHWvy1D719jPu
Yw1tj74hiF7yyEshdNxUw2xflCg+Uh1+Pf97v6/3Ws2wQ3jRBRF8zcUdnb1o6EBy
RzSP97mm0avalYP5Sgspnds8Ys4rSPO9WDepUnLoQTF9zwxWH3oR3mTLvG0YXF13
onIX0bVyBjklndv6VEvKorZuQYhjDTtkmZx6eAS4OutmXBD1LJdxbVsIn6t67CIs
UQrq0Gba6s7JDTo+EYUBbZtz0+lSFTc8KrIN9UGyFMSviJuAAy9CEe9L7oVg0cvd
rHns1/2OnE7J52/cAI50mRbuwwud1Xu/RUHTJL1VQO8zOrG5wi5inFfWMtt9+Cb1
muaag0P+XKezi7cTpwfbKmR4y919dkejba2pVtumRk4H6uxp5IyUZiRqX4xjyJNx
+T8vNGmOl1EE3zBzalrBySlZzdCdG3WtX9n32pbeWUBKwVSJW73RHDG/mUL55QZ4
oQWFiq+bx3F4HetKbSvhrOIiBuLs/DHQ4KC+vduiGRjWlMCRng2bfq/LLAQLdrMf
lU0jaE3Alf4+3YozUjzXQVXjsKtN5M/05oq/sG3q2ijXTVocfLq3Lx8iYMSVscgI
H02bo2+b95bGUVe65DxARV/GXGT3HhEIDlbdAkPkZIW86XID0qWdBuUGpASFAu8H
rV/6SPDshtlXPKvP22K9ynTknAZ/pfcTd3CjuauGGtD9iKS9mNZ+cxoappGpiARO
2TnF6rwj84YP22pcSm5rVbwm9swoYd6vLFxDdkkOIVHH67zN8OOx3plY4Gq+qv8i
u5Jjz2nq8b733f5j0vg5YfMEIAi7Q7tsNn6gJr/rqCSiN2Zw/SAQkNk2hP3e0EIK
OUFPEMY/GMtTatHj2iqAFsDug61UOuVNovxd1TYF3RIHTiV8Bs76XamXCvWZ//wm
ib7d6+xHAbxUsGALop5UhLoU/aSzwUji7xGyuXt2uPD4WmW37T3JjEBC7Bla0NEx
dGu3Ju2toyAlrS1PQJklvOgxRidXArky1COJYXFGwSGUd7qHeGd7+D85WK99Qnyp
8gUy86t8by8MtcQz8obxn9vUJYWfCqUYQ7C8CzoKuiZTxXttKCnM3hbnkh9XO1Vq
PslNc/oeuPCzMPdiQ4HslXWF6XyWNOFrrd2iJoYfmoqq/hlV71eO3KayPr9Fm+lh
SdF8LFbY7DjNsvJtDL/cOX9ZewYNTDRbfG6qD57sNKDSumdZKqgHW+RJNuAgMSMj
btg2kR+6Mplleg2PeW51nDi6JBEt+rKpayuRmxWiHOxecsEyIh37bdt6n2bT7J+U
J/gzN8QPB2XQWIMRnlA283GtPpK/6n6kUMd7zYox+u2f+73dAfzBNBK3ErESC+D+
qn9pXFuMsZb/4cV5iOmuqNDwqUZe2htegtZYurGyaZzYgj/etXvyF7JRTP0tL61m
zku85HDVbifrTri75OKaK2iH0UkglvLDOP7jv57n4NEgnEt+oh+jH4X44Pm9myxC
i0OdJvSLESJgv+LV0cAqVCaRaW7a4Hs2g8ldyhf0FhQiavIMlYWvQY+YzYJVj8TR
s7wUgLBS7k+CXieTecQDkiBJO3+Fs74/SuG+qd1O55pLjnqlmZ0Hhsns5Aoy5wP1
kcHMSXp52tT3ecKaxO3l43NOJn7p1StpVxk7nVZor57VIVrQv0vrGdbdlWB5MMIf
wUcxu+sgbDJmwXee8qQguxHckXOtweGzxx+o0vt5sW3asHyvAMoM32vU2nKNmvrC
HfqA82kQEaqcV4OnZ7Rm1mXCzJYNy3sw5nCZkqCjp6A6Jxl1+xcoARR5c5A8AUs/
G8zpsiRdEUj9s4khpzcZyDEjSOEmTONzwxmaIsuMONxESscv197rBHfuubfKJhZ4
c52FLi2Smf/nOGrUtXuWOIt9Ej2rwh8dFypvg2LGv4DrH2Q+D92AjwhcU/TWXvBl
O1SV3EKBW6pCdQkzYMMPJjjapjKKT9qPiyjGViCb9MKUYFMcDeuZdA52mBSCE2UD
QghOA4huqz/WyKqEHEFKZM4e73GU9kfqXyhOstVpd91YzlAPU5b0EoGQHb36CaXw
yHrrFBAMN3CgIg7fQFsx7jS3GKf4evjYe1UUAnGV8s43PVPJOj5hFMt9ypEm5UuF
ZbEfJ6e4YQ/I9dh1uCyc+xIbgGJ56G5eVyqM7YOjS5MyZFHAxGRLDGa7G+M6ooYn
FNEwT3unotRp66j8VR8OPP0tjfCFYl1XamdRmNTdg44XPt5+v14iLSBjZ1PoYGjV
rxFa+HA7hI5OLy90+yTVqXFZ5vsijS2W9JYWePJlvjzAiBEk0AVeKKDo5WBlKG/Z
s3i8RbkXVpIzGm7kWa8g0anPUKMqHrmbWOf6zJHZLtX9d2tX95B/DaWd2Wz5RwF7
cPEPMdGJW972ZotomSt+qmIvX8ZyyyWlvDz1/iVVAkTe2N0bhh9Q8vvWIimxgh47
SBGKmT96ukQZR+G/oUOrOwiqHjI9jez1LGssU7puqpvPhqMhtLvEAK0uOfKCbIC8
2UlmRM3BMhLD2RjKrYTP9b5+AgNAM0WDJsMbCkh20UUdAPu/5iFefApRenAy3pKh
JahPRt7ptA1p/qXys1Rf/3nZW3XOMyCJoV4Syo5hC48KuoZJbbcbHRgA5ORpmg5m
bGiS8+kYRkixzZZSREwiP6jjZAIpZvwl6X26p+nfOLIHVB4znkhFbLwNXF5TL4K+
FMX3Owi7Aws0wsMGI2CbTVbF6/LZGj53obwr32U7ITrlZrPDyHZKfYkQgeEf7AEY
96ry78pdcoamzN6Kso9Sq2K47hlXRgwWwtef67UWJebPWS3L7LaggLy0YZsGpYsX
zZkwggRsdb8ON3+9cnes2pOKGEvR4uMUXmW5RHKRo+rYi1KJ4ylYuXkkjiEwArfr
JNzIVX6zyRhltz47sjhPRmQGzHbLDxVldW6B8X8SVA1NhK7++FMCjEtxicpOZ8gR
8b6kMNDA8tGDwdOt8iInQbIIuHYeud3ap6KwxDX88uMLhxxxJVtLT4hEGXGBGuSr
ahGPNPLyOgKVRGi50/c4eg6cu8ENJxo8hSEefgMFJ+Glhunxj/DYrA/2aAea1uMK
cUwZJgqGkifbohBUbcwL5OijayLg4BMQWjoitOMxAqs5+62D9lYhvh8MQUR3xgTV
JuuLXt09ehF76+qiM8Ozwi5lE7fnyvKmlIpJhcRDgF2GAXH9aoDU6fppSt6SQi23
OU7e7rGXqsByUkfQLER/j9GtWLwPgt7AaRdvi9AnB8wUIT1HmNkCcUt8LREgLl64
b+jcgOZOsduj0UW1Dzm3KqlkUUqIhqbGTyA5gxe1Wr6T11859/0bxVrV58VJ5nlH
oYNdVOK8YIU1tuhtU8T/+Rxk/zuIEPaVbMZ/dTApcYddh33gK9ikc20rIblPbKBZ
TuAAMLRcEjEMPXoACtV5mFZn2m6yQyzaS3wzz4eHte4gqHthVN1aHkzeeMCEqA3Z
9FKC0AigMTrKA45SHV+4DyqvESfMV+b9rCwGWiFgg4M1RH+r8hY/2+nOa5jAG4lX
tv6CeVH03CTT4dMMfuRaZgsEikxf7XQB9ZhaCm6dZk8hAomDD9EyPu/WL8uk5lGT
ff6h9xuU0GqKgZQhQ8IvREMdfMmaCVlhPKGfTc7+8TsEgCXDRYUFDB37s4awaN43
XCW9Kkfi+Y8W6NZKzIZMmO8dU3zmSeALMw/tnVQ0a0LcpuKbb9iSK8yajEtfXWfZ
oqm9x0/YeIEDiFS5RaDPJMgejoAfn3sOUW2YooaeZZRPP0B63TrvlHBqz81PnfPz
bVtd4A/mwUU4YgpakRhHQ0G1G3Fn2pk5SGxredlWo3WhJyl1ELr4muhnDwKCjIhq
dnyALmwNSnzVALuFUwEtdO3MDjxIEI1f0syj2cL67vK8dEGMwGOlrnI67rfX/MWO
xX+FbDdpz5aUX5czmi7ka4uBEdp5Kh4GU4RJmdq1jk5FXvubJvo3Tz3RJEr6KQbv
MNtDjSRINlyM6RC1cjTBjxeEPHlG2cHARLCdGX0zSKCj+D7cBgpudmUTfoTInTLG
vZLpGV5O1W2UEuZK5gDBlReLMeLVkYEbHKbhMaCCsmNvjoda4HkiEyiN+3ol0wfX
1veddlMAOyecGFtKCu9+hhe+UJx9170R3cAYRgYBT7hTuFejx664GNHuDgv+w5Pp
pk0nmp67zM7RoIkyIYdGwi/tV8YfriOojASSjn2rwdyznB8A/4xtPbJ8eguA3A/t
IzOq8KubeewayCDs5hQ+eF+KvkhApTK32X9oqXaSBMKGrgv+fmcrK5pDi28SMBAn
eL/fNf4lMSzVTCMbu3NeThQFmsUZGLM/c4VowwsVqgveYLOixzWad+Wt85rjvWWw
z3C46tpHzq7m41gPlCnGzMMnTzeird5MjSzgaeQbOWKlMMHryOpNAXBfclSnRPAg
bYqy6Lq3Yxx92a+d9aJoGjhPZC3/o4XV7QLo716X7I/QbKZ533DygQZgKxSI/aWk
+HlibGqXJAsGDi+kze5zFoi3eT0t1HDP7Ql4qMfv0U0se2G0wLaHd/38gCf8Fhaf
AcmTz+NeXfdDG+jq98TsZ62K25vnAt3yrATX2gajBLPdaA1NK/0yA3I8P7/RWGVX
bIps7FhMA80qswQMKwJxQyxPi+ZJkDO6poFradUh38KoHQ2kFmadxCqiwYA/9LUv
y33Ylq/mjVyP0/97ikSZdn+3uiCBGkl/37bqvdbbuN/5ztV4i/XV9cK3sDxMkVMm
7fR1mHbO5AeDpa2Q3t10StaHJrKsU9EJ97y8aehJKMmD96kF3Oic0W+1WxW7TIyQ
e+ps3S7H9CzDlplEIzCcap8Hg5r7rNkTaC71CBJ4tp68GA1PdsqA0aVvTgwwWOfw
j4dxR3G6+yp1OFL0brKmuW4rszCh4/BAqKWbX9Z1T9tmnEbEQ1unMGUkYVpct9gb
OWt47GT8m/4BPWa4jxaR4+CmzYh6PlQ9/tLCzyU+z5jj/uzoQZ20tiJ88W48QaGa
+rLXb676TXKUiiQKr2h1TMfvr8EqZ7MtRMSWtB4F8PotKi03VZfVkwBE/93GgG8G
A9/RZkikuNoBh+GlNemz5WEjg/1GNnbR54uY5KgClhBaF9MSXMS8vuv171n35Qgp
MsjF0630CnDRMZiMWmne2bQDB83Iv5+iOBYB5H2CR5WIg8f9/NSNtsfiXH3sx99S
EBA4FNRLNMRvkE2W5UxLoVW9B4JvwjW1XtEzlVts7cxQ8rZTnKoqPbAl1HRNxfNM
gtwBMrwV/ryA9i09S/GctWSPbNTAP72STjVT9gKYfDk7jtnXkLl306y9MohKKMVi
wccoE5bnQxyMrRMnsXqfS6amO0eX/BbaCzRRbpx+1mDqJR2YZvi28vt4IUE9LtaV
pDdzKWhTa3ErGOrXYCE9ocPJeFujpBjmAeLk8iUANPYU14XOObcsONYbkAvv6055
LV+b1g9pesTD4uEpwG2mrgT/8SNRISsKuEtlr8Q4pI+DZWJhHykqfR8xm7negeOB
qR7/dS5M2OCx74FYTATcQmT4AFdKLW/2BAwN2G6n/a23ISpdpqzrepchJqQeEz6P
5GioD6iIWB2ov59zOnidyyP2vs0U8/BZEdndiOzwjSqm2F/OSidWMDBKWqXACH+/
fLw6NHSM32EwZSl9S1/zPKWVmRzYx/D/IFQhFGaqhBNUgAXzTSEXARRA/d4kDC51
JVUDdCl9ZesN6JjTnVEcnFIShvcO3lOdCstoDK+wwydxCHl1+lsjZbf+b3ublY7j
t95U9ngcG79wbXWw5vCFieI5XH/CLdn5dN8tjs8kXIMUXwmCyoIVdM/Z+sn4vP0l
zKBndg3roNk5c0yzc0dMeCD7xdRRz6CoaV2qsdccgppKZxzPVVcFiycL4H/WmpF7
KcFf+BJTuhPZcGFZ7+wgt24/BtN70HgNNybtByO5Zwg2P4QAkPDrxNrhUDlquVpA
/aVqRM0Lla05U6jhZHbLbWaUD9C1cgC4HJXGHnPj0ZDxNKPZamDR3U0jIQ8foAS9
ns6pGGyF0gGGngtA9OCkkYmfFopVjNA+yDZh3MgZXEO/o8xJdpVb+BzprTzJ2TSY
wJawG9s0UBWmPrAdHAbCY/QrCHuekoPVe5N8gHZcYasofoPpRLo/3xX3TCt0G6hx
PDTEqzOZpT5z56dlDgpO80RcEUVHY5yKhpj5LCY3cBxd6I2GDqPUykUusoQvcPx0
u6SiE23AQC9OUIAv5xFC7pTHl6GAt1syMX/MBYsuBjmI+zLoBKh+9nGHg3bz5Pyz
O3qd8zVKsS+XhmOuKBhiQ0O7GCmtJN34g9LYgekRxX2y/35rgsvY321ghH+YWES9
GAlecbQsyxOskaw5rzwJy2ttaG4CPA7CnxOoHJ+SqwNqKMKRRqeIRaTxrVp3C86S
y0SxhmIoEf8GYbyr2Gvb/bS4ujd5SlWjDpHlPBiCFW5/64da/GtDOf4IaZ1HCigW
tfWtExM96jZlbqV6eLOV9YzRcFpvklMmKpTGZUHrESz2Y6uT/+c+7WOl3xhjIBiz
Ry9GISm4LtnX+qyoVFvqM5/PvFAfZEwL9BoIkEUb1Zvaeg+zXTnI/P6lD1ZGJoIt
4SWPM8TcdFGYXjCK7erxhulEcAtVTHU/Jl+X5h7AlcpJFWlwCh8qe6FOz61DnAx3
RX7YkIUbNDCIUzTma2JJHK/Aut7id+bbhzs/QuopxbxPB7OWs9HfSPJvfwWLrdw1
eTZu74I0O3VPrDsz9pPLXC1tR0GQz2XBRe463EB4Sy7tsq477OcmpswV988jXUHQ
W2TAsDdHL76jO3Q4ouxq1sQuCzltkCoXJyHSHCw6NPgEf6h8hPo6YKnHn57/mTd8
jgNZO2mzhlAM4spUmPgCD+LU7MFChMHAQR5JcHgHFX7iRaaAL/BrIec0Dbv4JwlL
r3Pce2JB15pYdCC6BUFLi7HRMx5S/EcqPJCpQohBazp1jrwQGcRkq1iOt/0COR9f
kUTwBAbxSUUywIfJPYSjb5TMzE0+qpLyhq4+d9QwVMrgTjP3Kd8P6Lr07Y6eOkOd
rrhrDo1BWfLb09xEyfJQV6q+fpOOcAf+257SFYSC+I3QPX6ROQc2UXEe2XOceWpq
wCFI1+Zy2dTgQU7L65IWdoKAjT7Dmuir2MvMK9EgHU4kyPTn84GxwDQDBYAYAOuU
wvb1/Yzq3ho3tt2TrKcY8FF2vEVA/ro4Eb0+ZR1sGr42XvpVlJlCS4qLflRkF7Ly
0kIv9OFhMis1Xa8gP1cZgmBv3J2eyS++znuNlRk0Gvcvno0x4cY3dynJsvFbLlJY
8s8ywgR/ApyCWNS7KR0gGacNJk7rzV/K7aQmdyMvbLQBH1eE1k3rsJbo8mPnBqxZ
ruauNwILFFiYWsDE6U9OwSL7gvAo+J2jpc903QvP4C8RormpYjvwtJT4SknS+DCN
+hVL1/jZkPe6pwV4IHoZBDUoefrKg2iqvtMjiOAnB6C5y8oVjxCHtpj1r4p808N5
Hwhly+X1Ru8jow67MiK3mpfaD5WxLLwa1ot0zIze2dYlCxhqNGd+yuVX2bzWiJoT
Rhq8IYJ2T0gtegJ8Aqv9XOGMBWfw69L0AdZZyLUvv9AVC0oDWXT7z1iBrbvYTpVw
FzCr3XC9dov/3BikRgpuY9+LiLdWIQaedKHzJ9w4MzF2hnzhIXzh6ITDtdRhFR3i
3ZBR9wMKjLVKqGziYp0nPZdnA2s1Ew6t0zTLTUWVu/y3hzvp9//s4aLR+xQHB336
q2CEhfCXIXhCXOkUV9yZkITi4eL+doMC9w+okxIkELf3ZT7n+oPbfvA8GHECE5ZK
tplgd96FyOw9aQtWFVq3zeIEDVvyXBWq4jAyigpQ/oEy4IbH6V2UO1lz+AiGKhh1
BS5ezAH19PVzR0yAXJvWIPrvC11csuNxYVt0pu5v/T6DjZE6+FQnDrCPo3zFJXDC
YHIloghQzZb/METofjXwhPY2RnsO9aFTdFcCc75lZl3XXPh/7AvVSJeh5EvMFB1u
ymE0Ts5VubcLlSuwyq5PniHi/RJViKn0YnqahxAP8eOV0U99LsYWno+KEdNQaee9
99F0UfZ5lWopmaA5t1QfNHPDIHjBJEBYOq8kngU1wtqxSmIejEltu8a4qnkxSjoT
oPJOUZsWoU06XsSm+K9O9dezssta06+W6b1Yj6IBUTKMincLHpaPNS2E6gqunlbb
zMMsiXOkiNDoil9Rw9tLfKPLKf/AO36TY78lz0V0czickNgMjMfGDIzqlyjZiMiz
TiZ6cL7H49f7xZ5KRBxs0m7Y301SkdVbGK4oJZL3GTd6b4cFMxHOF8IiRMRLQbrd
hHpWwzbDJY/bvGX2dhL0fsH5/psKIEnf/krDKkzKyeqWV/vWmyQrSY2ZbMcVOv8m
keQw7VmX4xZYIDtlEFNE9lYZex2/uUHSEcx4wBdhQ+L6lzUsYrIyQaiM6t3X5uXS
ZVLRdwLHwJ7cdvGznEFV/chvGMq2SdPfT+riND7EW5BDQGhyyBVWW1L6eaj+6ioa
b2BENk1UjTUBUYpEQafyhhV+MmXvNjwxHGuC/ZdCjCBJDgxIChlGL7bCCzqeEihu
dtWgYGk7Gqb1sX4+JG/v/v9OfQptsEud1cbpI/E1NB4dyAWOJHiArwfvWhJyb55q
P4mMyw2kJxJz49TlPm02CharxrgUk2eOmnYSIBa39QohDmOtxtb9/D6R5b+5QJsj
ozrRik1nRqUAqvVyM60hwZDon2Zw/61WjWmUKwdOl43+eNr/WLacMGrUUJVoWu0M
BCDZ6p6nhfI9007hYMQLCfGENkb+fJzJkLyPqAk7kXKb/k1Pk+4wckaHHA1OkxYM
+orPdQehllIsD5Jh4oepPAXKWOnpl4BhlUvXjrdP7D9CNF0a+yvC5M/M20KFeATU
1Huv3vfMcqoa+AY3P6TxEzIw1qZAbnIh6IOQ/fhQ85s3nkxvs5+qa4wjdO+sn72f
/C09v/adIEiLtRUS5lAw0fpMTbUYvXooFfUthPSYKafGlza7YbAjUYwb6F/4EFyY
ZVnk24FvTZ2REhpDfTMv6CowCHalxyDbMkqJhjaSobdpxZWlVZvPeepfyBXKCi5i
24whPrrQ34aHpT6pghII4PAV59Hugw96m+MQCW0b4qxqpvZURkjkY/HpbYbmiI2a
FSNTPGwUIyCxna9OvcUnZcug4w5mhCh2EoZX19FTbzxbpG0fb8rSNFATSJDrEZLt
RpEV1IT0vFX5HxQlTJbF9SZ5uiGjTp2o619GKeNxHErvkQBtMb/HP+cg3KuRWaWI
AMZq5vcy7Dl2gDm5Xpp/aMRu1Rr08pi8zoIB5TAugHf8lY9h1bAgHgkMmSgZyktw
u5XdfuSDEAc+5Zla0nQwstSTIJ1v8h7b47/aijhKtiIbhOipWMjTia8/UU9/YyM1
9Kxjj3VDlCcYBh4RXlQwl6ptX22s7IrLP91xLvSpxNTX01MlfCvx+IP57GONVHl6
wPXdu8fKG4NTLlkOM1brSqqC/sMLm6cQ8d+0kP0tL5YTp3QaIGWwWUaNPRVD7E7P
8ovLDB3ZCXDaMUQ8dTCYw4n08eHSuv13FIv6uyVGeN/IYHSi3aciAiQqA6QJxZkd
1BGPd/gGh0YcFdWzP2aTynUvNQJJ2pJcW5SuKotJy7R3mQoN7YPv0L7LnSEMacKT
55tQL7sAQ85Cu7DIZIFctiT65qDffsi5HWA+A7Ne2swIw/kFPNyH5HVA8eObheyR
xYq0GwAaamo02oIchcHN8lbhAh5UpSSkv8RO33KOdiAfQYBxkBF0/BmwBATqR5eZ
lLGFXabyxWoUvNSk2miy3xoCkaUkt4JEtFToWHztNqm+DluPjIXSc/jc2xB7/GZt
Wb39ujxiNxi+rZyzAXPadHxPPfeUz9wpmz7ykjk4yhVQUyK3IiX9ZFcBrkAvLl+/
Tee5PTDcw7C83FtXLewG5mFOFTZosz3fv/lAVONQWfcJp+DBRk0BxufRpGhZsMFd
5lQKDQq7KVfaZnz5R/qbBnMwRvcOL8VePvc/yHKe3MZzCBI/3OVejLYakc3/IDYN
sPmcnZ4n3M/wO3x+lLiCe4/MFAWVdpmhcvOhPDZ2KSgq1szXLPWdZFOfvqLaQxH/
9wCPR4xlBt02z/fyKAXsIHTTpnFfV8Vzf+w5DhHxE34zeUbkEMvbxT46s/jvt8Yt
vY7fm7ULyXstahc2uRUb5gYJgttjbjlsjz5Sup/wzea6O5dh5WozAN+t5B7D46yU
rgKFjQnTcTK6zOnN4Aliq68eVmQjOI8JUTrIdq1oR/SfZRgnEz1Mrn46GQ7S/yqL
jEQKEbgbEsdIN0uq95E1WOcN+aeiesvvSk3/E+5PrahqWffT7BUCFgL7OM3PMhZp
ZCoYk2YPu+uomJv0EGRzWkhX8tsNvMCPRxesINdIAWdvIF8FmkzYnxav9lRYjkhs
6ggQzO/AF6P6UGwiOPzKA77snC3Op6ip/LfKjKu0zRH/ga9UQxDt5id/TSvli+1k
2EZQYc17biFt3gbr161QELe3jAnY5EO9niSscrkivlJMHYQkGR2p0Q5OI7YCeW3D
YuwjxB98PD81mV64GxxkpceQQMTn3wAICdSAWOeOdFqv7bxcsuee6uRCpvGpCJYY
AlNJvodfry73bnUoA8/Dd42QvrhHIpZc8mIWa3tLdg+eiSg6BQA2aEWJ4SSuFurD
CM/lq+5SwVDKmzsflJAqKjk7BdxE9hHatugitzLilTqXiMYpiZeAtkLZm+pPgKuf
/s6l1yD5iz4mYH7Hjv7XhiFK5mjmMx++w0FeCtX79XQe9LQrENSXZT2JeYtHDn6c
NDj+NaCN+Rg6WRk30QT8zbdCXn0lFOoXiScXetK6As/6zhve95DrcGZAxE5aEiXH
qdGLn/NJTKwelleIUxiJfO1jsyjoimzcNKWOVUXvZ28MSXgdFd4AVjaDzGTifzKQ
KcAvgf1JUA8tmK8DJhCWIcnnpG7c4PjaJZKsyRyVLKQuvc0a++uLNJAfHke2SzjY
blEok5QWHjWKkzsmuWx++L1pIPgQo7L2AfM5V7bP5Kc6Ynf/8TjFU7bJnUXlMKm0
NeT4LkJb6j5F9bMzbMLy1vkd3K+T13/YcOaL98esybCOasMG2drH50ir/gg5LIuG
3N1tF5h7bF3yb3Crj+l82nVE0z8J1zIL0QNscFUeyrA3rGBUAtGAKEpEk4TFqARD
8oinwZ7HngWtgwzjOqzCW+6QjnLfUr/rLJQ0TRzpA6mXpLabwFqCCzhN9boR3oM3
oVJoor4SejI0k7iPY05hH1iO6IzQBssBo1XWTPRR/Ate3iSE6+THSjzCmrWLp4j7
z0/LE1HbPG6nKfn143djNqujz92Wit1eIucqqAk+fQIu70hnLfcYYsZB/3ME+/E9
+XcwUGFwHY3Iqs3y8gQaMTRNasC992LZ9B7adOscPUkr5IqOzzdNTTOx1rPuIaH0
Mxvb3ky8uToF3i66p1cPBG9iFn6Omt5Ptcu8zV2z103ps1FyInmvWlGFtdUVJwI/
EAhjetN/RHOXGLDkBw7W1MPM6Urlaj+Xwmk/PkucCdqoT0BDXZppdaEtu77jksdr
n3BcpfkDq3rZAJF0SITcJH/N2c+DNt9c2kLwtgS7H2kUcX/zKbvuRpNvOzgNUlsB
18oBa7a0eqNuNfURc5mEEXcaK9MbwyhIg/osdzoC4nsyqrcBu677Vk+GhWxd+PYP
0F76N1mr8cxOagXAq8eazDvryFb3Kf+6HU3VYrkY9ordJldVCCsq9x6V6cKE/YYA
jmnV9TSQ94MArs7F+Kfu6KH+mBO8g+yWTQnXcpqr8MM57A3G72lyhqbarZBOT1Vy
AChpqH9NvHFe9wkZCcNq5vjDl4epQlvOS16CXERxRTfX3e6U3n91gpemhonIj1X2
GhWkNS9MxqBDSuOyScFrz1/zRR9qmygprsAkHIUiU2XY6lLM5ZonTX5s4mHbE6es
FI4gybS568TCJz8HJY5Z1wrzdodnOOp0qOoGCWaoXrPQKAot+o8y7eLRq9EDCkab
D4NSeyNFfpfydfQBKQnY71sMtsGayDtjarYQ2QhWbDtjjtBSfaEwycJw7OwoLj9s
4cXZYT+Ah0hZckhCh431HGPMcGsBBRXDNyvfohlOr/2YDlMFaKzGovRIOnC0qtbh
91Py0TyX33611aiGtG9gyh45w8SlluMizdweYBu0QkkF0stFy6NdmgnwAxQzHWDr
WeX7mp2M158sRpsL6xf9OxoxhuvfzxI7EG5Q0dhVV6s70j33kSy1uoIVFE6Ka01T
n2xrDgdAEKyk7jzfAaYRo1h+UINEit9Nx8MdFHU1ysjqZaShY45N+jZPgkH1rJV7
xzmdsH2UnchHr7qpjB/heq1W977MSHjcjv+4ZyK0iqd5dz5PeFcKk2SQoc1SMhWH
6ae8O7co/8oyBOavO7RHMtGlF9kOcvclYzO/xji8LD0AiFmD2pG5LPSiPI/UXkl8
POsAj5eEIZlisnBqVazC8vAK8qQFRIbMCbUjU7MHIur2iKih7xMm5izcMmn9mWFd
Yxb7+M/ILJsJsci/CM3qF04ch93koYNEv/GT3y7qr+dR1dFNuXlNBMwkoU9HGG+i
QCSL6mCxX4fMnEWo15hVRL0n5AbKUas8Dz79EmHbsFq081s2dPLuikskQOAt0DU4
Ijs/PUvdq1mqDg3BtpCC2QIbNY6S4lW1RKhdnhMIpZXxABp+pxD9hrd1aerjJNDq
Kpxd62xNqHF2rdxokUGDDJRQBpeD++gCwmjmMfvh6VHktf2g8O0aSKSxTEN7+U2H
OMKy9dzjYBgPfdXrapPFrws+ozpgQPHv9kgKRhq6LcoU0KE82c8iYQfrxZ0revs/
GA7scPjXNAu20MeLvY20nUmP0XvzIz3C7inCGSRzRdA8VVwlaCzU/ZuEgF9EdRsQ
okchJ0O4hCNaI02UXvbXYJrtxmD9UNe6N1FOgM5wCHAW7WFyd2HVCrk2JM1c34Ja
8DeC8Wtu1iVmqygdPm9RZxc2vlH+T3tixtBaOGRxORDtS1kLyl647hCFIWOdNDP3
Lob438qpiy1cjcg3yEri9jPP5h2GXWIrMO4MAbKsVAkGOlV5/ZEcDsaOOBOZ9GA1
myZxJo6RSsQyWsBVp7ktTPuePzlYgZeo+H7rqn+oWipdvG/7t1C9aDdvmmtq+flJ
l/P5OIZQbdc6lIZpYC2r1Zr7i++IvNsF0IMk4op8WLM/5BnrJJ0Oe01lBr36C3td
9sS5B/QqU5i8kwSbGBQjRtctAgUQ2JwcOaHB/07Ig5ygQNph1hGP3N4QnfDc6GU5
Nq2nHEXXMqQMM8GdkzJFxBMIgNFP7c6oo/P1Gqjas56PNgPX0WapNA8/FabvgJTU
p7PIeoTtXlADAPfeQC4uUK/7j6k1ysEqt2atne9KqF8B84Wh3FYYMVbMJDAVicQa
NjWe+wT2mxO0vHSUcJzCxBTQiivyPMAJWCAerMUwkhgEeSpSR+TDPv598k4IY4Gw
yCT0r7GKG+lrk4BiDB7vrrJUfSXJEKdYvGudlDjySTgyYDX10jpC73wcP5l2uBUG
mNlyHCTj40xa+f40viTNhI2HOkuhvAlk5dX06sMlqb/xSo3btNTTQwjHa/Inx/3U
XhaSncbbW3vj0m/5vdJLvMQk1GlRjU4Gt5vxLYH+guQYeVZz5tyshYNW/PI9osYo
m0FhCs6sFCCfIGNXKDqZdf4YlBT2u44hd3CTbi+39Y6Yigy/rABBJby8pj35q69+
1gP9stRn08/zznvXRvSV+B4VC9uCUztQwflkQI1MTkaE6Z3Daa8AUN2lx104vLa/
Oouyd7p24Jvcpn/tfq/co/TEwKdtiJpQQbupzLcskpmrPo8JZrjqMsMs+6txru/6
JMHA6WSt2c0dFTT6KljufwTRdY4k0HxPDYJXbIBTqJZR3r2Vygly89TfGvIdVONY
KpPKmv9LgiLgvv8neOCgCAeeIzrCiC6o914Sg/sTVXYStC7/ga94BtCTYMtCYTFf
Fmq+F/ruVYsGry6jZg9hdLVVU7tj28knvzoHnKuCyrotDrAXnhe/wP7iZAc9ZULk
wzz/uPxIhKogdgwxZ3cCUGvrBF56Rt8GJ4RK9TLFTEeVpKSJEZAIpD8/t/++12Ww
O1XOLLijcoMxY+2CwLmRiFAmG2XCnCK2uJ3TTEeVNM2JwvK3Hg1TTssFD7+EGqc9
kKs7o1kBtUCBL+sO26fp3r24WAeGaPjWxEro+Yt7a9x6nvdAkR3pvwo39lHDA9vi
oPXa/Z+I9bN1mZU8E7qktuHSyqugl2IQTNLiO5b/MmRazfr3cfyRhbmYyFDmxoyr
X2T5nbV0CWwd0pzToXlqGQ6CoS2yyIILC6T0qFRZkr19YuJPIEle9GinNS+s+4Mx
qxIsFF8qpY06xklXMgFWNv9+h3+ZTwq12cYLGYwjSlOqhC7HYqi1BHfDoThLSu5P
7ogUIgYU3hSW1WySviZ194iWT0Jzt4jtynGGaGjEVPm0uGa2I06wvQal5RsU2D5D
16lFKCriayxrAIznhlg+GGCKFOIPOiofd+uMYegLwpCGwChsnkaevlfZpLZRpOyb
aVeIH5dxHxVFJeth8ZwtGVBQxKVjcAVWqGRWQ1mc3R3BQdoywRrVjf6g/2G+Y2bX
9IQUPQhNjp0uBEXjpmGC4J0CGN7TPKvXQM+eOHPOteJNCwc+1c6pZMAF6OXCeM46
+aVKwVUh6xJyCpBhKxExFfSdNQHL0ZItHInrv2CGXxatbo/V+J9HJDngrXDPQhLF
o+F5r/1nHaI90ktFIMTWxRe5m3+0txj9ULRN4Z1RugN4y44/1AaNq8NYv69ao0yF
0dGDZC7XxD9LxCJViMvk5yq5AWA2jYDgPx5ea86KlVqumbl7wXSmwRnWznOkWw85
S+CYDN6UqXgs6px77XuOG2vvs5QLpQ/1AnOiOTr+oUbZlrR8yYDOdpYxS4fajP70
vC30ZfEEyQpRpRxvJz/NNqeF6fg1Bpj1iCbYXaSUCI4RSDfyRJm5m78JBhEbwFQn
ecr6SEiOSIbUYSXTYXpgaSFdqQ/WeoHyvl0QLr5agGJfl2jRRExFmnMW4SxZT+oL
OQnEz8Ssj8WUORF7vS4dH2vsItCWJFYLvkcrazUaBwn0cepHvo2Fv2rANXRzQybA
WmV50FelRlKjv87SYMGR7qxWbn5ACBYGOUj8xExH9JVDo4Q7oVDZrEnM4Yzd+RTt
ZtR4xolPWz62RFHR/rAe5qgb+qiGs25egvhcPBaMUlw08sDfUMwvdN3bm0Y7XyfF
XkwkPXZ8Bj8nCEQirHi99WOwKJq7tRbM/zj3waVUQtUxZ/PWN9wRh4jOGatjec1V
IjNVxNZCpJWKHZU7tQzyCwc7ZbZbT8WhXBvrMg1TJfIRN5N2eNmQyOJEN8Ay3s4X
1V9RLyX5IxPuAF9w9t/mqEElqkwaHksviJiTyv+voLk6ZlsK1m/J1/6bsyijEmBo
QL6Aywu4URnlXW6uiETHMKFOa87BHr3E/7YUbrZD698enboUhyI2NMBqlFFyUwxu
69XdhhPIfZzIm4oomuu39tMPv8nyWG0MJx1eJXSMj8C+oAVsYrzoM9mG6Bt5T2yU
pg6ybk8ZYf8/uDlJlxyRKQrJK6bgQy95SI+muOCKH51RV5M1CdDRV2Yl8f8gK2FZ
j+JhLT2uOKWJy7cWN1R/5k/odbkdefrnKtCjU6xKgE4sA+GZi+2nRnfgiG8RkW9q
AzE3Jzb0oUANa77hXz2Qc7fjKwuKGMVOAMQzsH87e7YzOMvrRdC5qwPwIF4crRYP
1ip/050Gj45nRqzg+09Q6j/u35PeA5z2fJpJsv7guwtVuDlM4NsjfZSuaig0rHwi
a75sXJd/E3MUS6OgyHMjv3P/9besaPzP5aALxkk0O3JWokH4uMOHSNgy3Of+sY2T
DREGdaJUYH7xaH4G6r7KgvF89m70wL/jlA5Bu2/ARZejl7V6JsHS0loDK3Y7jLIe
UyMAwwybBn43lMQsDCpFt/3j71a8oaubElgs3RyTPzdjgfS2qOWdeuzXEK7TzM3m
pZkDM82xCz0ptkjYPsqMLfuNNHtOXRr26ayVqpsfK0VKwNrxiCQfKj/zex7OzFvb
/mpoxaQdLVjNM+lDVXn1plafOPhiD8pDyJ3ipNqAjcsZYc/O+gtXbAgXDmBk8O1e
wke2WfAXc7Fydv2SMC4CwhJe46o5w0y9imOzxuHRJvUvzho0haR+l32HZPb/+glJ
fD7ZopDwxq+DYDh8ajE//aYn01vjobSAhRQrtbPGeZtoxRoDyt8MvLLccYnJztq8
JoZM8gChj78gWIlaJlQ+/vt4vtQZdubcGzmtcxDkyv+MoXORI0rzuJJv7i4hDI41
l9Nt174c/TwHW9LnNwywkHvtuT458yTPJPqwpLtauUKKaNXfIPwjCv56rmM4UwNv
e5G3jbtFHynBZPmPE9EeMRyAiq6ZuIjkGuRj5SLK5eNG58SLrR0M362aEX4dPseI
XtrG/yFzG7bXZQ5IWZN/P8R9uB+LMufOsj6kntY8a085j5g+RY1djgwB/Af/j3cA
OI/qWxRMxQEWFFyARRpk7cxqmKLdmgnb2uxdlIW7XKSdnOmgib7d8YNfnal69GqX
7fBxU1elAMsP/CXIHOewt7DZ1B42A/3Ak4ehx3fHHA8maBxFAKDAuWJI1Mo45bki
5zzOqoFqwVENUf+L5AFf8QOLdrgebpWZnt/X4O2kgL3YdnmJcjhpJaP7dT6kiodt
Om/xyUkUMaKvgaLweCj0Xvhr0VWUoE9uFgGepn7fgNDl9Thk329kPc6uppjnbsxS
je6wpdG3fJfDXdqna6AQQiWiKqLb1domzH0DXxI2KdqCPBN4soOgkOUc5/3pIvF0
Yi+Tlsk5Su9FXGhoHwBeQK+QtCTtC4GwLv5yj0tHr4G489nh3Q2idN8VvdZ1ebZ8
CrdEXFeNi0zGf5AGbUaV0s1ZTN4K+1dUhE665LuX2nI6/0jfxg4cg/bmpczIoazh
0y2t17VHuW07/3XVzg8vykdE7laOvi41WBMU/WICNqWldYvA888GFEV6r7YCBf+s
e3tnB1AShPFP9/MPgTpINEAsE0OQBlLhLLWCc3EPN8oCkEAphMXlTW4N6mt6ngXk
lhclmOcbKLAIFRbGj9x+/Rivl59wI7+jOxemNN6NHJtIVZV3P55aNtC6SZS0Be5E
ICRj5ny3qi8LWvxwoCZkHJ6Ckh3utaGK9xI9FeLJ/3PBEoRB8aioboqksbWzjcpx
4UdmvoeJk9vZmaGMPF2gkZP7tp2HjvIwERyJMeMm3/IdfABleRwhS+h2GIsVN+G5
MXXSr+Aqs4AdZiyRoQKq3Q0mqb5A1S9RRS1DyysSkjSYYJlNgMgtFZOzjG2KHaN0
kJOGu9jZliHgkL8AOKes728eIp59Epn2IafJWpUvFTSXa3wdprMQqJehyVxh3Vox
fAKQBggipK8YNlM0ttNmag2ySpp1HGhJljliGtKNrEF0dSwkRVVc7U5JsInl4rf1
h8VPgMSJiZPzLa522GQge31kNTX5v1Ih5ihGUBVDRQF4yoA8PKExJkJam73fAvWE
Ij6SpBw8BoigTZmwj7NGmVaM20wftSk+vqiDH7uJDa97wQpoKWdpRbovrY5VmyqP
9kqmcX/td2KtylOF19n9FJ+qECxir2e0hBNBrjPceP4DwpDuX1/DeGNsby+Oa8P8
S7sPxdHq01XZhIOmVgXbyzBJ8vFgdrhH2NlGK8FP8rBC5o2LhU9oqzHI58ntY7Tx
EZYvHy4uPRhOyxnbg2m6uF62gVS5asEjz21uMR4LUruIUqlK7agLr+waFHwFHup6
WBXqPyhYzvSS2QjE7zBXeNraGyC/tZ9YFFll4/3K57iW4b5DDNom2qRMc/py+X4j
bA+0QL4fCKzM/O9C967T9PjhvGaGWt7joAZ13mHxPkdKzvBLMpdwDVDnHeNoxSwZ
fnssat3s0UJ4k/A5iScQZUK9HT27OIqWUkvkxb2QaCOFEaGhvRs5XKnaHypToJ64
99Wu8d/lpOmz8imB5eO3fJQtF6dgkruEQ/KdZumEoNbJtRwKdairTSEBPyI/2btf
hgvh5EDxKU1W7OoWDDzvRSLgvMPG9Vn427EAaWgEGRG+tL1D9i1Rew0E8c1ww/rD
gDEMdO6wawmHbY+Fz2ee7NnDn5OBHaZmKpFFZiHvmpyojJXhtT4uGtE3ulOwj6AQ
GsozkfY7nzkqajsJXJp+au4WTcEmL2mQpxFke8PVsCv2DDi79UDBDfjUPqDgsno5
/9FKApgSdC2o/ouZ2eBal3uK1Ei11eIFHblsemw+NtJGIe4BdYf60JyUYjynaa1/
61jQWIy9KaiOBdJdhHmE/2etaZsfLr7RnVIMt1rJpwDols3XiiunLZRsplN1XRuo
9OlDM1WFNMX7NgwRRK2pcAvHap37QwoU5P/vaKKgz/9e8hkkSNXDOSp1HtZBERGP
UoLj8ShvAt97+rIvt7JX2c8HGyqgBoXC3HDPRnQYNBjSt408ikghv2nr3kSvBshZ
DBc/LIluWVwH2xo02qdzuIZcA92fuKhlzcfsgx7CR2LTvnUqi6z+XIVBuPssMomv
QEMyjp5MVHkuu7O/Z09UEk9ph/ds1kA5kDe13b/49Ui8KHYs6qXRqUfcvjhlAYCG
+yRmVEyRKkmtzcbdZDMim7aC+e3PLzsM5/tm+6Mx5I+BCkCmA7sqeLHPaLT3dE0u
zx7QyYyKLJkZtetlVTCbj/ULeaIj24p8pQASKtYctbwRhsexsltt5jYY77mdZJgc
9Jg9Pk+BGxETxhnONvz/3/2kex+Bo+ViYx6C41TNbQaxnDTeuOf1Iy7N0Yb5qzjq
HiJ1pIeeTu1EdEXY0y+FqyEUTjrLfqYXFuNXoYwsF5o60Pd4nu64sS19ixcP+Oi4
1j1ZJ4ndDG6E4997T9wEXXmENgiJLKFKnRjXnPOJwSDnIZyM5NT26Aq9y+2mTcgc
5Eb365sffSZGsDW0iLKx6zXUjUTfTPQGjguOAaGWmKF/a+7Aqpo5OcOCrdiuw8xl
oW3KB8Z+mlnm6lDFTzBMqeXrVSgrHSmUJTpZzSUrrYj3t7EinvB4NjX4J+9/R2Ae
INAHyP8KcK3pkJ7p9MwUrc4gKWvg+Z4YpZYvGNbpgtkCi6C77r3Civh5VBbUcDTZ
pXYDyj79CkwTb/n1jMzpveCf7tc4RrrDUGhhvNtpeEJ1CHEDoonpp0aITb95fF/K
ZdBbsvQjZ2JaQMJ6+IbbaaZIpHcHh/r249flo8ziexoXs81ZIU4FnPeeKp2xk6RR
rST4UbRC/GZBfAndBryDcpZrBRz4C+HYahV0y8+PnNZ1DnaesTbLA/ZVndgfCMpx
xDy9/PER/cECFkX1jEDJ6EaYVmGcIjZVnNr1sZGNvoNeL7/qS+g19AbTIWM+Vr1A
nmOd3ksu9KPRcdLP0chS1fbWY7C8szYiNs1djGq4ZgNW/Mx8PWd9YHwJFFr+a/aM
Cyi1aEkZabwtiYwJHe9ZOn74zfbXMxagae1zAFYOhMgBGOIXcyk66fxHGw/iuLBi
bxh0RW5q8v/5vNbBkiKigXjdZ/VGOcyUVuO5g5IGQzxkbXmoOrfWenGAVjNjEBic
WICwIgpRjz7VO0slI0kf54dNWhl/S3EJioVGulCItIKTet4slHiQoYSVMwyEUiUv
2rk1yXmhQelhJrs/RwxNX9gVROi/xXrnz3yw1uzZTU/cIry09ilzBeaL68JFNOlL
xPjR2M6MNr+0NFBWMUoMIowAEgVXXj8oiJe8kkcIaUKEyJQlfIEmVhmLadXGZS3O
0CHamcddemcfV8vxtJCPVWFVDazslYFPXqI1zdSH8tHmlblr35UIyeBdoNylKc/t
1qeUYFdFDvoJ6997G4lgOvkI5Xunti29piOH8uGek/JIj1bD7lDZSt/uxh5Y5SkH
/uqI+nqImlWS7Le1PZQX2Uk4/+8TE6Q9de9lekWpW3p7TRi8UxTVMqOF5mxphsAp
NFXfaTqidn7CsxJokm/rp5Te+J3Eq8GfrQY3QTf4zWnBQczMKj3l8njvxc3KxdPU
5My8N8TmJqbvpdh0RKL56F/gMndZLmyg6q4YYpJBQjZPScsIyeuO19KetVclMxON
Ak80GdjYN6Z6FnZr091faB4p0nvcj5j1aIKk30OpF3qiTQ4GOUXRCgIFOwxRd2vp
FR5N6qUsJ3dHMZ01NZ7to01I2VdBK6SF2ntLNg7f1SiqJkE3Gj7G3ndiGK/i7C1+
yJYcVWuPquXVEWamCwcAa9udvx1Jhr7mwXiWa/5REj1Og8k8vJIeDooBGTYeWXdN
36ebU0Bqcz+ZMjCLZmCBsP+ot5AgmN2SkfjK3B1gAQogKgvQ3jR9/7uyW1y8i9wa
FuFYiRlkEMYdaIwOuJrjKLVdIwTojX0FLNViNwbeIA2ZKTLbTXurvFlalUWvj9MM
ydQp3Hmbk2tKTyAXfgz7Ln/HaDQaO/AkxagxMWLu0XXIZ5sq1eG1nmNOiNk05Obx
mvY2Ja71R8WJa9aTd1co00GP6066YpG7KQrnuNXFBa8aQQ4v6pg0YdZw9CAYviuQ
Alob2FXFzgNnI8zfOZCB+aPf0OBWywRWT+hi3VoLJNFg5RHjyNdXCJMFKLIK1XPY
mveeEPMqKM6e9rlZ71elxwFYef75yvXWW6M2FWa8kAC7Sm/MQ/swLRoGY0P/PQPG
gumHCszrfkzvZ0i9v5JEb1H4Wv23fVDZyf1GikRddBvF7cFtdqG9X6X2Yb9Jg6b+
9u25T7TC9B0uKp2mEg6xRkwauJdHuLmrKBwZ+hQOTC+x810bVnFcYO8y6V5gsDeY
itNwyyQCwGyrWOtBazvr0I086CTVy13+hUUaJqSqA79Xt5/cEm4eacl+r42tHMa2
JdJacHmsHg5QJL4eGiSrw6CdDyjKSiJUPJ3OaAy5Me2gVpRCo95nllhtg24Bzkzb
3Z3XJ1MAn6HNWo+C3t40cmvE/uV+rOuHPU/aU5F1E7EFcri2Jlomf+d1k+L3Snxf
aIZvNLr4726iJoCHSU+Jz6kXlQLyN/lrHJIC1/TdhLml+oLKGA1vmwEHqjtKbEDG
to0pC7tqWb6Bdj/p+6Zp2GkqHQBNDiVtWCZJNa3j5COoznsw0XxfA+GKHiBY1h0r
t4CaA3fWwOBkYBvKwleqocyvnnsc3qCE7Tp2JfPzBISeUn8C2JVqFj7xQIYz0B6X
jIkw0obbTaUMlSIe2zQtpf2kwP9ZGI6JN2nmAJql4VrvW3xy5SbYGW47VNGvRf1J
3mUxMFb7fZU4XKl1Syf50hyP7A3M2pbHeqAB3VzrNruMQNqnOUwn5swSY93ryRP1
eERoACpONGu8PHlXjC1fvJlr9t8S/blFjUYHdRjmeIpwmqUqkpi1JP0LnXRRaq/z
t9ToMYRdkWnBc/9+S1o+2OCbRomcEoLs8O/YJQMWlXcZ6pl/FicgQMZjTvqEiqMX
eETrLyq0RT0dOYN+QY0oA9+Bx2LcdW1u2f0SAq1s236s+CY3HsiIj8gKBpFqo6u3
Bx8NO3eBOrqnXN0Z9/nuEdxZG29HXEaTrrQTdQGa8J/lpfGdZgBOpxYQcE1BmRJB
vnxrCnYuHbOpO7aOR2suK/RRw7FRGCt3+wGVRbjHCEGxsznlGYHNGESE8NUg8JYI
3xwiGLZrqo3OgJpAlS94dmEvdIel0I1Rdc73Xnv9EczzqyS0M7fXt7GUdIqFTu6L
Z/le8Ic1SRdTfbmVg+Bqxy00U+GH4Bjh2Klz+SEr1ToEeODwPMruuSQ+jR+1ZUw5
u2gxEstcC6413r/t3fKC1rYhtnQEM3xIAQTLLDJh/tlTt1bhbcUsIGJzb8RLBOox
cdNMQkwLO7WBGMXwATO6ujAEnMd6FLKQyZdu8BIx+b1iG+Cw3txYCHIpYywIaiS7
agg7k1xlKuRbz4o50tMhPQIBPCj8ZUSUYIEs60UPjtoXAMgUy4Li1ZvKIO/+Gn5n
QD7JLDdQkwEBc6+DojkgWvbzzq/+nBmRpuy6m6Pq0VCxMEBBcRCaoQ70iojSQ6o+
qXkUUnxmfCPr3kl8te92YLDWomo97NMkDl7t9iBfhpET8AWiSMNolrpvA33saHdb
1JBvrKH8gE8Iwv47Yd7bpfyNRDsE/JoKhKDCRaoFjI0cMuq5kjO+L/eGX47LghXw
AOrT7/J+e2PM7m66lxTKuq7jv/ExnDtB4u8Qfh191i/zBSzh68UL+tV3D6Xr3qxQ
zaNCi5cYXhUNcC4+ptNGFzb9vt7+t4GfAtwa/geh8E/YJILM+kxd9OhhCmIDujDD
FaGLh0BO0uOmupxfmBx9cRw4E44X7H4THiPYEC+JaJ6lpdt5ixOWJjSwhoD0zSUa
k8v+F6caVzUVYRSyx6D+Gg==
`pragma protect end_protected
