// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 01:23:58 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qH9zXmr/qWLqrHQU3LMeHbN9gY5xvu4ScHzf91LfaVvO/7eToQ4w/ubjWSmitdbW
ncZA5pnGEH4Gzgvr1W0APJOwDZH+mYwum/d/cYEKIqtZJPLLcUm2kx6LebiO8rYx
K+icqRxZ+S+uVwwN2wwSLGN+ca3jjHOZpl5wwjEzeDg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 749616)
OecdOYOg7aUm21FnkoMPycZHVnj8U7iQVC9RtkrCFKns5G0gFTbRdEouqKZ6V2gV
0o7K4NeeCK9UZBHvkNr4iXkwyNsjR4qppWwDoLLFsJDe1h4GmwcTs2ET1tZ1nU2L
QwiGkh3x7opPL8txxsWUU1r5og5lsPAYtCnkppoLlpKKlCGHnYnPg8emDASTf/Xh
/AnAn/pR9qb+P/kds9cq/QjkNtWGSi02Jsm2HE3t+vZbyJY9t8k/wDnV4F2qs/Aj
7cio4xKvSGbChmXcR+wdC1J5BKmuhZ7X6Z68shQoGoJM24Dg4cDEA7UwYzek4nY4
36EGsCQWbrxo4uVVNcvPpXvmj5Q2Pe1bzObO8X8RwPXwF+86NcdE6vzLbpQ14PI0
3bSnL2Br6Oqssc1RuPeEM2Eb0JY+SBtJgeRM61sGuiXp/WX2W9+cQ7yIbo/MXy9a
16AJuJb2YwEefPgBtl1d0RwXDjG3wK1BnEZgnnwp6Xj/+5s7YiEKar03uJMsmcKG
rQTAL/dA6B4dY59Fw7mNsYLxf1EyLU7e+l9NJUI8hwzWv3oNPxjc+xZTcCUtNOfB
8VDDJgT9PcZyZ5AfbFYOFs8i5/w27A1+uuR4m/107/BCpfcVOiKc83Eo0jez9Evc
S+CQ/sy0ZbAjqxTeAaNYoOgR7JJW7qdpAURUbVwnnm2nCCQiVnliG3MfVMRwQkvo
U4JbG4UZ2tNFi3U5t4q2RvmOELh4nCKB5Wk4VQ/SqTp1efJqJ2YJFIW2w8t9sfsh
BDysi6dogF1KAnDcj1vMjI1At2BrrlSThPCIGp09D0/SHMvbDPSmMKzGZit2qkKA
DC2TNVs591XG3E8TmXKuYQFJ4mvdsSdwF7vLgm56PZvs1WZcHbu5nWdIqbtbopZ6
RRqhXCb9Oqd6g1t+ABp2MVqGe08J08PuAfDWRXYM4A5+ZZ/mjh2HfawlRjw80YXB
09K4hlTVyMFkdy6quH/RsD6RiVn0ywX9jM8/BBePo8netololTZdlCE5snRvDyr/
WdzS+vad0RH+WpV3yuWzc9gr3R/K5BH+QOtavkZn8YJ4p2yke1SODi1RhcPuOQDC
pWwX0gJXi+iKjWZArfeSCkdxItH1fN5t0weEUWKRuAxg9B11fh0Bt8NMyOt5X1el
IAbQfamUllptp6jbyZCsgC4F7+JeXSAsJIbVqnrF4oQjbIVE5KnQ5N0CG7LuZ1Br
lsgA4UuejJ39+FYfaV3XWxz2kWOOmgETLxtC0sZ986ZDc5uNgF4G9KVrBz7NOWmC
6GCOguIYmziBvsKSo2EXAiNOOJaFgiz6e0g6+c7Sc610yu4ootnTRnAMhq3Utv5U
hrIYSAtasu4uH8qbq1zeuerYfaJATocXGPJHhNNkRrEmFQlpOQtdOnIdA6ChX5xN
TVcjDeyXAnwrCNSPjsLFFqr7xMW5E2tPu4Mab15AnSNMiisgKwCwo9XFkmstWoLI
QUI/k++2x6H3ABrPZzXh3uBwwbdBVrVsMYyd+oZDJbIjYQxi0jtfjmfgAeRNCOPj
jTbaxiDPpZRGh1ILi+OJ42yMrG0x0Sia3dSF7NBCFsgzzqQH6ICV7r+db2nU4uMm
mca9ij1FF52Ryvw8A6yHOY2aMfQqKJgXrs/VREPjurldvolQWKJP8ICFreohHFWE
T6snjcNyKHbPVUI8SS3LcmpyfLjAMVLd94hu87LTfU8Ailepc+tXdRLe5dEJ+abf
p0STKWdy0+jYlGk75dN/hBB6h0aa3nEVOSphFrB/5hC001z//4eNWJ3akGmPwmi8
vkEatfuUogDcV6tRFf7vQCqWJcYXcNdIUzuDEaFrNxZR3Le5ER+2OwHlsyuKGO2O
H+Dg8cCeQ7PUcgUM2GQmO+XDHaQpE+ZMgvra3u1DMU2/v4UfmWTDEg9G7sdfGIGd
c0K0KwdOyVmeru9bg1eN+7MPz5+YQ6xtL5E3Kgf9wIQ9zIJ1Qdt6eLNd+z8j/5Nf
zb2CPaOW6SctDnG5s91DfNw29UUjNqIVe9pj7Nx0bOyfka4JI1aJ4HBZh28byb7I
vYM+GUS8Sr2yH0b5hn8fVMD4ajrf9LEgF+nIV6E+ZGmFJIwoVkrJl06Ngl4Ucggb
v+SsM12WlsfV+TDIjkRZE1vhDpjPpzAOkvPuDCFw7DLBSE9Jkc5onpVB4fKlCBaV
+vQAgfDWp5vscBbPdbWNe0jR2OowsrbKqGCQnqLhxRsH4fRba1o/hXKqWo69aLid
QkUiDmwBh4jiuHWOKAJyMqU0wqBZ2z5Ifk5hyv0Ba+R81M4cArJfR/c0n6tNsMkR
mVigVRb8YTWxEBzesWDT8gg4qKmdPPpyBApB4g8BA+QKVUaAYBlBft9dzrD0PmcX
3YMJjfGnBBzd68xQzbJiBoE7vPhrJhXR3g17ygFHVznhabWWWSX8Wqf7CxlJUn9W
9pVE727rwfpCphIAAIkC7cS7MXDc8lWA814Cbnm0CHIkKKAQZHFQUovhKfcUptDE
5hHFDKopfWZAg3jm2BOLnSrl69XkPK2enaWmxgedYOrnYKDHkknMiv2x4Ue7aZPW
pgPWQxxMn0zYWHlVmeFkMO/Hv0fE0LnJipD43PlU2gvPp0h3juy0GyN6+pKs7tyO
XMxh2ewRu4v6mJuToqMmNIDWOWmn6YvMJ8tcyE7DcybE2VqYFCz7k5hspTIOAFmK
n7gOaeI4WfVguzLkFt3RKB4SSGSacpRHkYOIZqjwEKK8fKP6dCEeJPkCFG+j1vbL
1XnTZfB5hdl0K5+8jS2H/Essrkygz7DrIvZO06EYcwj+HRNiXnpUuf2SUlGTGKFL
5yLxh31vzs6H9gzMKWH933TvgyXY0VdNPeApzK3jiBmSqt9SODYr1i+Q7oUEbTvp
cUudlAWwbe3Jws+6GciBxgu7hDICoj09Z/0DrjkaHwpfcHNbvAL+JAzDtVTg6vEN
x4soqu0UckKMfyqJ297Vn0rpNHMF5HF5GnVzsQJj2gTBsocIRb6aLzXB2coo8ksx
zad4pzUAIW99paG8BJ4t8PJdOQ45fkuR/snI6wOg2AVWHs6DYMvmSN0aX6dgMHov
xiBCkGVxnjxOJrN/brS4vNWt0MZejVB7xoZmdQQ053LUK4F/0t0TP/ankEPhG/qs
JsaRfP+ajED7HI+Bevkh0VDqnJ6K9tJ2oOfeIwIn8NPBhRjuNVy/1DNWN8Jyu1aR
ESgvBkuAoXpZGf47JdM4uPSE69t/1sQxmzMUbldnSMKn1zXYV8Oevy1oRADMxzv8
7eHiFQvCZs4XnGHQgOTxO/WEserdaEehBZcu7u4FFPiGtd4icgoJ2hdaK21MYMsd
nHLUyVyNPey184zwYcdjQEV+bGIe8lL6Mg6d2grrVnNaNth5s4VyNm0/rSidiy+V
OVTGeB05ujD9r43Tf9poW1aD2utUfyDJkz9TCpW/GzPIr1Nl402UqhpbVFY9IGIf
ybPSzt1S4WdmYEHrcGQlLKHHH4VgWxigg8FefejrHduKIDLhI8avuKTY1eiD17cD
1n9h5ZjqpJzuClxxCLiE4aZWBUBkVmd5KjjdBDqaLEA10CMaAgjZR51qHJQTHoFi
sTWFIj3chv7itFkkdMWGr3RzD0ERJ+F0ZNZsoGW5XuHjcFf1s/vL1T0GXOA3Whsc
l+t7JsepBqSPAhfNkmEwUjG98FJWcw1ZH2tUQ01HBcnc3Zkj3ATu9v81n7vgi3wA
P+5IpDA+Gb9sNYHC+w6UDDM8kcGw2zapH7tUlBc0Y/mvxoJah+CDgKGX/0JerSzQ
fDAWIV06nwv+gzHteBKCrppeBnKLuRmptkISRBqxsyGjPmTQPgI4XtOJi5oTu4Zg
Wxi6bHhbpPvrS4nrEtxGidBeXCCtYBg9omHY2dRFkYDgvzpOglCRKtJhsW3jpgPo
wrYJXX3hNDn++/tZjsALcokhU/5BBEjhkoT/WDyfhvCMvyWGjp4piYRRx6SNmQV1
R/1pz1Br6vIv17mLzJdm50P8zfv1FaP7ILm6SyNcZRRXPjbn29A4HlNmZoFXd1iC
LPC3Lefky6KgmvMQCs/1URr3UNI+oHqs2cj5cIB8VzrPeVmZj6QAK6riMa5ngTXZ
XneBadwRbRIbzKT05XIDxfEgVknKsoBhFfdOe9IV+T3f8Q/vsBKZCcOPDUMsPIr9
58ID8P5piQxd3QdsBbV4yUfDQooiV5r9LLBai0jPL+uOFwE+FOMNx1gvYRsnHPOt
iB8eR736euPGr5ByHORpjH4C3H4wrpAboTftGQf+b2IyUeSQ+bZnDYS51s62xK5I
lzn0ymU331E86E731PvPBQ99k5qS4nQVI0Lmb+83Qgi6/oFdyw3hlRL+jLB1NO9h
DImS1i/z5DCmqTez6u01lR03ClTfU7UuI3ldgxPrl1HIH4U0Rd/fH4h6xI81viZq
SUnvLa6CZrzmuRpxfE5r9JNPTU3XRw+wDkAYVZ0oyiobSEr4xVnA3c3XNYKQQ5bn
yh9FfRX2BNuZa+0v2gB8IuADV3bGxNIMuYlX7k2fMtNcbjlrjLn7yVeC+SwTrRQL
L4OY3LykF0U4a8e4apNhCuuoS9hLDGcVj4yA9kHrEZh89NU7DeiAb/j934J3fahG
Zsf49QV326bGkpD2jvGM/ofalswpH1nMyxhjaMQAE8SAfyDWNqmAqNcl5P7KYr/7
ZPBvSuQwXP6fhKGR02cS3fgdPQZEXuexX5b+Xo3cgnaw4Dovoh07Mgo6bSb/pOWL
jd13LuwzfbnO4piPL1aGUfQoP7eLcN/nHVzxhOYuav2P+0MeHec6ilfza66zeCcu
DfBenWwWTXM9nFw4pKvX1cOjDox1h4DTmAjMv8qSAnlEPh8RAd3dPE+k7hLsXehA
yd4x/dviFfuCq0I6M3cPoDgrqvtKu4aZkRxXTGWoWj//8y405rhnQ0StOOeXty8e
Ru+gUBYW0f4OIOFKvRLRzvTPqdGMzwjHrGWrbxqPyjgikKW9JtNPDM/z/LlRl6Mj
19V+dSceivM1tJOLIFlRyBqBe79xjOSHF5aRnYENgIW9EokR8vY1+H/gdVDfoh9g
GwyxPn6G+0yAu1S6pmMKXhUOtEcm0ZSLz0CSwlBiX/P4lCAkd5A3FH+Lyrl4DYw+
xJEuOdAKG8MU4u9f0RUmvWEy2RhtV2e1amK5CZQog8mFZf7bw1nJu/uRRgPpgVGJ
iRPNkLs7v2UqGwtYdr5Ke3wnb1zPuWSyY2MX1rycZiJWa9nmFlwU8+bVik6wnFBI
zj7HdsvzJYeTVJMV4c2gKx9K9Y1z+if7/ggR1PVfYvujaHPJZjP3C0qbMCbRF//6
7+BU1es2RyFP4ikE3wzP1lO8EYFYaQZ+Wjkd3kcVJaWas8iX3TXajzT3Zk8IlnYl
ovPXSDx1k52hszt1uNY7Y6KTPP6mxN+UKOi8D598CkpSnKLwWRb9lvo+7h+oAOVk
5ongbq22MMZthakrOg7bGSAVHgtDnPBffafTIPxAY4OHquvbibFAT/XnijrPvR23
e3jo5Pl3roMhfyAAPa4d3M2jzglcqI1SZCZkIqsHd/xQwKunJ24Wa6esEJgVFxYQ
VBeXBzLfk5QdVa0UPCGOVF4agRnY4VUUe7L2IgVCuVtOtpU95ARZru1M5jQxm0fA
AGe7BmRGGmo7//mJBcALkQaMmLzUq8Dh1FDAehi9kDg68C4FgSDzDe4EEI98dn3D
N+n7WFdeiQfriW8EX7+dAgBYd3n64ueHMZJy8WA+dK69FC6RpKDdkQN29Wlz31nD
fZJb9KS5Qyvi+AToctbRTeAbm3V4XjXcTykMrAf/NLeBRM4StYR1rKrAVKdqF36+
Uh8gqPkO+LPd0J0p/X/u0FiZ4SA3UsSM/qyYhQv7rGuFAn02ib9lKh1uwkKYFk7C
MfGz1g6D+5KXHOBj3LHwdAdlUl5boPf3LN1Jo4YBQ6H1m9CE1RENJhMR/k3uzr0W
BZtHvyCkmJO0JIm8oOXat74wH2zkwCReOzg1BnnPbEW0XMPE0gPzJIqop0/rM9YF
o+GeA+QOoCli6A9VAc1BX/Mnj6Z4L47p/7c2J43Lp4xoSoilh4CKAIoWcWWzXnib
3gircQkSJvdJBehmF4DBlfEWxrqYuxeuzm6Atux8/cpiMRsI5Pi0nD5jrRCty3iD
kfReXl0aNth1fMcTSbeMmBF3C8UC3c9NkvL8fiEdpNWElr4uMj59lCVvGv76BIww
AlNuS5vYeIIdY6GBt5c3x9s5J7QykGvn8pJ+TpkQGaw2lKL9I/flJzvP66WdKYBv
VhijBoaqnCrayK3tTcMLg21Rv3hgfTjYRZoPc4WybMx53uL/mDobXoyn7De0svJ1
Y0XEpv3ghjIwZ4Mke9feT/XfTD7pI378wGfFIMq9SJp1zWMqYJXi/NEwpZ4ulwmm
N9UNfBxY/BxvShRx7oYsyjcbi0vPdjHY1SJiG43QFFd8UojK0LgRsKHnPBeSQyHz
xEgdn8d0RpJTy/4lBFxkSfPiQ3wAH5C+4IABxgm4AdgxQo14GQPbLiPSUCtjG8SO
uaz6xaltMdLndoE8pl7W0qHX444dvtTPaXT2LFyZ9KZz/iaC/YcjkbzbZN87UB+4
sZ6k5Db2GbwZujKEi7y+8WhpHQp3d5fDlGX7IXBu2Gen0hu09Zgw5ypTrAZh0sqd
cZXWvbIf0jDC8DWFYmLv7Pip74g0zc0UUx7Js/jcZY0zJkQLJlqkdDEP7/jnr2L7
mB9TBUs1HSrxsHyo9fpPPQZuH5Jl3ZiUub9m9qsNSP2Z/X5RuyGduid6ZTxEpfcj
Rx5mCZvzbPbDyDkpPdf4PdMO00SD9BxMH6QbeCu+AIV7bQj3TNQm1u0H1KH6yYQU
yqRg9xc+w/v8i3GLkkcoDeZchaT9qcp9m9gQImWbcOglBeycRU0FekLnoknzxPei
9CPRG38Z5PUih5kvFh0vUxZerggz7pp8CN/o3i8nmwCI7hI3lanCOG3Ff0CHLKeB
YFCFdh0OEVsL4bYpDa6cdWRvsjzNXhsH/D2+JGz17CXUWX4D8Wcwldti1H8INXpb
ED52PfhqCkOjPr0RNYxl2Qu7FGo39I3Kzd1cdwugSKBn9t6Zz2WjNGFrbZ3dzCuB
zO7uzJa7JrM921NBx3K8RCbchfCKwe1CGq0QGigPWdgQClKruyqLoJ2RbEZbC+0d
KRh9jdAvCZ81xQVij0MRH800z9WDlxCdp4TvlMskk+A6n91CITQivgCUqdw/d6k7
X3/0UF7bjpGWabc71Me9PN4yM+oOHqVWiUnoW4ArTVmdeec648SbPMu+qPSLQLRl
lK2k6xXDXVdXb198g1M9//rhMIL9+SHfExJgrqagjCXi+Mhb1oMV2elvRmM4gsx9
Sw553GsNZHZhDXdNSb/wMeCZ9WhZbQKyHUdq+qN/zdmw1UUKT/zRozXAIyrpBymb
6VkZvYChTUpTe5XpWL0YaQdJe8e6GOH0NAPUcisKeO5a8+0Ojii1TfhfgfXzKaM7
Nr+kqOY/kZ0LxAlua/obvVvLBrz10IENP4BHDEY4+G6vGWYvWQ6soe3U74hYzHVP
tkuqY2SKID4/epVu5Q336a7bS1flPULKsNfNlbydEqR5qEp45p/OH1Xa75tFtHLu
f4qv/7u3g6AsmMfmtBhGr2H3BNP0XP/+gsbDN9r1TWUJap1aSyR0fWdXRQtnvOps
hNh9IbpB4EaxaeUNw0eDq6WMTGWiGWN7nvtuGWiNZHWW5d9i0DqvY3UZfIZgOwB+
Uvuit1kcECpJxrKoZKP6adC8aqQFijz/c73pFXKRRC5+FXME0ROUfpNZjELXTSz2
qSUzT11QNn7q5spCUDwij3tQ9fdQxQpDEi8XYQLiS1zouxb3SbEpMPkBw08YP5Gw
UGFXcM8tYXUZU2SZZd1cxmJQmQalESSZtghZLoYNdSOVLncFcZfTAKIrF9T+FnwB
/71sG8NShEgmQLkseZhzgIb/sg0ubhY914v7YbVHlQZPD4jJB4EeVXpRK1B0AnW8
sL1G0DGxvOoZ1CoWbieZSOLFGDM6IcZt8kooZIOGy4pdQ1Vy37kXaQRK5jy4hkAh
ACDw6nGcFvCuBUoi/5Ibj8YZXaB/aWJxbbdT55XSc8uv5eyo65Aadr6MSIVE6qZp
mPHWPyJ7syxCUREHgUXF/hleULsVZDBlRdxUKX7JiRJlsuXyLMfLMP4CSP2pI8m5
qK/AjA/vkPFdxReZS9szmPJvHNdT9dOWhUzNLtuGNOJRI3cH33fRx/d6IWwadS4B
H7seCE/Pi2OT4H5WPYRZ6+08ygWbiTqQYmsMlyoAXhTut/oWVhBk50At6sZtPrg8
lW0XcNnS8IOdZukCgaWpV2xwwuMy1bzoi8KVOrbCiI9Y99OBlCtE1I4jfSmxql+r
T7GhMiCgy0eJPzHRd4wTlROTW8RxPP5+rrJb+Zc6rH3aOGxGvoPq19LfyLdA3sWz
bA7uqTPHDK6JutvanUY3POk0fzqgVZ2XCXTLbD9NSX8YtEIw3OER4ow76uvusECx
tcRRj2NO12hQpxN2Fxl53tTDm5n4NAEz/6WolOiFkTL5rAkWOuc/cps1qligYhDy
Z7Peor3dD9e+tkM7O7QDU8413HhKTFWH21l8obm15AaqzcmYis5pe5holTjAtPEN
wqevIR0sa4jSqyI/v1ZdP8Xkoj8UWgDDavlLKPxFk+ZFZ5IGeIgUwJBU1LzFQh2i
mfP+VrHs0XhbJGjLc0oYe3RcXB7A0rl8AvD9wI8hOsJ4cmY33VAt9H/6ZATDxDDd
GaPRIcTHPhxxEf/hWG5+UR3CxFzkNn1vAN4EvPAjNF6UEjXZArDO1C4OSgv4RjYc
RU0JQXFAnANM0ia+VP9ywngztOJuo6t3pr9h9Q9DJo6g3jOMKwIIIBvsPrh75/sK
RyQbEsTG8fuAgBIm/oK0RWW2yJt/umSMbuWKTFiux6/ExLHUj+Y3Ko3Zf6GJl0MY
Au+Ym+Aka15LUwA/XXrZsAWdwpXcxEyFR/V9y32qjKc3arF0RA3HHhXPoqKyZnau
Rr2iKfK6J65fyPUzaP39QokwXxSb/KbHYUy4chrbuvPANl0VXjYEQi4tv72Vplsq
vVUMsJrspQ++WayZf90R9CUk3wlpfy7mv1fKy0XxfaxRrTZnvjAA/+pfhdpVpM7Y
+ZTnmyVcKsQ2KNi7cZSS/nyyurlYR1BOB3E1L+ZvkGGYU+e3BqtfpG5hJtYlscUq
NZ+OQ7cjJRdW04rvAf9bh26t5OIUXaIgCbUwf/UVPjcVqc/wEA8N81QsjGZByTDD
c1GIMVz0ZIi5e9jOR4PEn4AobntmTnbhsZ8UwlR8t+J2hFSQyfljvLpnveiDJ31t
43WquGYnQM9S9pOtglFz7l5tLA3oOYB/w+x4gwUpQyaNMleUhFF0QayxjLLKS7tp
n9aHLJGu5l45xEZwhes5eRMpwrhqhvs7ubuUXnEFlBLQQzGvrcKzv52/dHkxHx9z
Lg3s1fKVkR9mt1LBUCBB2vnhabBd15WWiEPhNWh0+jpBQDifZCZS8gYLeFAbW8I1
EvCNreSkIFx8364C1F+3NA9UvnDwku7ZOSoa1MnwXneRpN7GPyg7fuFr2hud6b+N
x1TB9al2Co55JPpB/PIISMczU5CP/qqfxWxZZMPTdlpG7N4T4bAKIyMVyIS9HsfO
UsbkTwCPjqfDVOfDi7SWugN3pZlU2svL/O0Mddhjh/ZVDZrriBVgy2njMEIhN6BC
svwt4/qmSpUkEB4maj6PnYwrJqcSTDK3gaSExUEMlcsQVvRi8GMtMQwgy5jDsV61
Wq4BMiW7mJShdWa82SykyTaIfYe8y6MIHY73TlmssYDLfbiY/Lbnr0m8gvCttF7D
YelGRiRUT5Fmh2EgQbb/XSWS9kDp5gOBUkK85UIY1Fwi/fAG3uYVtiCmAGE7u7wQ
acINRJDhDMDlPAtytZ/Gj4SvDh1SA0iWunZj9jDSyAWnByfFk9+KKKc4G76sPP4g
A4KtfzZH3Jext7yKfuIX5AqroSP1TOxNAb66KyuRi10EsdFdASr8NgmuR9aEvTY7
d427rvNkPRaL5tBuh8fVVxQ+culAWsCd1dTwvRynRZ4/NsAbLq0XLQaAa4xDHDsg
t+2+XvXlJ85SeStXhRTVaVO2it9P55dmG1gFJ/WYTJodHkjRLW01ASX8ZP8BW5Kg
j+TXDUJTGHTvR/a3yqVEJOxvJqZzO5xcREfdiOuM+VHZ8RA3OcdtUicktmhCrIvm
KTYF2vwHpjrVwqPZ8QrqGDOBWjH10K2umxBw3q5OhtJX8eoTxI3Wxgobed/EBoO6
kXBArBtcNgvWP2tgjJAKuXn9mZ278xZqdhCxwKOqwI5njSkK1oJsiQqjLD1DkP4F
b+hfBoTyEbAs82bPr2nOqjViFvg0E6KCs/QR+MUL9yWLaChDapdaHCeYUQu0fAFO
Qs5tR6R1wRDCzu4XgVw2t74q1jP6BYKs/ocv5D3VDNtOKwyZk+gT45PDZkXE7RCP
XwdRarF/jVT9xBX/fuuZw19GcsTmdwYNqnR0kna5AxLV3aGjxqVIK1/8XF+YjbA5
jrSl7wkFR2jYIUSqqJOZXbxX+iERfQJdDZXN1PpEqQvBOoTHTrzP1iuq3Gk8W6HC
3gS3ZUfHAX+xJ2E4HWXzZXS+sNLpB0j1q+hlJArOBb81tuocWJDNZ3JNxu/Pefwr
phuMVlfSGwTkvly9+T4LCu/Af+uPh7yIkBENFIKSDM7QSJU4xelmkypN4arJsfDk
dqLT7095gBjcN0/nLa/30gBXuZSjwBSgrcCqOkFyRq4I3YkP+U6J5a5UUK8r2LYu
gW4pGLc9LjUIbijghqDomShCsJXLe2nDg30cVgXGFtCJLNkDZhhyWA4hLNzbr5ln
w4vPfKxFx4EVzFgJHWxZBGWwSsKeVVsOeFPdFlLtBRuS+IBM0Pl8UdXciI/p8ZZv
bKn8wI4cxH8DDCoK/VT9V1UrxCXJ13c6L9liE9fL3xR5rqnvQPmMebVTrut+nuMC
LheFcHIDjXqk1TatWK2SgkLzOCYkkVTLUkfQLGgL1hxvCvh+ugOVnGBZd0B1t3wT
Rl5P4oJG7OeaqB8jzdIpp48gsKCZWbYpi13gRr19TPGcKoQ/2kmoDQK+VF5x5w+1
q78Eh/Jbt35187I2BfqY07v3wpV61FnCRZVdj5LQscxVxct58KRb/28z1PW1ifhq
v+CBvqu4a7c2PzgKtplSmWQxE2HBNPvkcO8M9wiekMjIyAQmXi4XZ0H9Pp4Hcqmu
oYC1u8uNpicT9SWGnjn+by2pSyolI5QhT57oFiEAbZRjGPrTzfF0/9cHSRQ1YOaE
ugfnCKJHpfnEvW6PrvuDsjWCGgFtCjhtrUxJUKUmFKdHbvfRt5G9r2UqH6aBC7jz
8+DGzlxmyIpwLkYfMUr6g1XLondHCFoXPlGpLLMlzdPyQThPT3XhJ3+Rh0do6Wza
CAzh0fu6fXskJrV5HXC0+GlfIq0+uaiV6xTD5w4YBHFclhBanGtUg4YeCtJD74LX
6utak4fQhLtG0OKZ742jsF6ueaUPo+9g/sEbp18kSreda9UwkiNLCREv404RqFsD
/0TLpvj8SK4faodDpdZujkaTwZ4gU9AhdzU3AOJWZ6+HQOP+X6IrpBwOXu/lblGN
rZix1fcPzSo0Sz9skKEiNP8fziCvsVRj/t4FStP1Jo4IWlpVarysJoumtUbjzTI1
+WRo7dt3l+ywho1AO95syPurdv4uEmaAPgU3itck9oiB5FVe6gv+21zsr8EtsrYI
rLyRJY80TO8lc5AZMr9sV5eLKTrebZGtCdNUi7ej+XjbCjpahTkAPULzrAJ9x2vA
uWv8SIUnFE/kh84wiMdoIXzzmfcTGnXK5CKHcR7Fk6G4Igt3SbWUDfAsuQaiMXio
rWUlXAwxIj9IAAzJ5ux7p19pgSlC+1b5oL4KYw7PvEES9uUqNVud+XkpE82O8uWL
/XF4V/yccOzDuJXwgBJpW+8YEGXWM4ER5UjOKwnAP8U+BfQiH7J3QlrRng4KLh44
1VXVxGsd8dizmCghNjQMGMIGUNTv4wXxbV2v4FRmSNZPwR0CIOAZINxbKEv+j7SI
HeiXsXZoeFOBcWWIGqPOEA8sWMAO6NT9Cfy9HQcCcjdP7uWD4pas8OiDUJM0tEts
zt9BNo18wx+Aa64F1m+4jzQl6MA0R9ATXx5CsFaXFST+sQU3kzJBLHec9CjNpor1
vg74vdcuxofj5PcGrlFTWJecu5TyTP1nLh0rp+nv2TO8x+LCXr5Qr/UEI+bwSCqv
z1/kVxho4YUfrvjW5PW4qal1YquNFEWYuY3NrYAtOTpCHn8z0Y8nVCgMTPrz4AwC
VdD57JzN1ORmVZ07w9IqvU0v4xbhuwyBSLEvgj7fXokgUAepNMf4jqnYWOxKSlX9
0gLDyaW0NURxpYSaRg2Duk26P0TCfF1iWBcx9TmwIpm3qKW7kNkcmqBNIu6RmXDh
BKB8UDSNDFw3bF6SFlYSf8v1I4iHP+qwrU12g95HX2vH47YGZ56ZcxAa2flg3yrr
zP0Daml5ksjFPzWLui0G4RMhrqMyDM6PZ1XZ4AZ9QokhzJzgimeSOq3hNKElc6LX
GNjTlacBoHROO3wjG+4Yon2yGnShbf7k91ZvtSf/McKYbu64/nxihJIevvczi68p
Om3HDtkdxTkJLATA0vXFEiemLUmhGbKkdfL423B0B4ycMW2gtrg14dgVuFYoe7qu
rrc8rZryrLeFORXQ1BaluvENnHYuIEJMPyUF6mfB8SGveS34IeOy6shm8Z8edSRt
12lppVFS1+LZ67abbnSldWzFd8titbnOewI5XCvcJmH9Df12R6s6YvrMlq8cJPYl
HES7ReWplFb//Ltun4GFNL2DexICMgSsg+yPDovs+RCCWNzddz+RU8Vkfy3Fah2O
+GMLsogLVqBdTWwEd7PLOsRmEx40dvVctak/P+3wXu8OFHTQCXOiXATlLQ4pyQdT
iJAltA1Gw1aX11s0t/k8KXUiaQA31KvFZiMcPEc4iJqgtb186WI3CoQOCW44vgkA
CxWnL9bRM2wYNtbgKLvEzowrkg2fI1dB/xUt1PvHLZNU39Z5kVn+qp0OmiX0DxEe
X5cbdYtd9Jvpj6HUc4gAiFX5CQqKVGvzkh/++1UopdTHEVh9/CPisk/ejb82giNF
YgSaStGG97NDzV8L4x4Szo03X8xftc4AhuXVWXuEVUiXW+SPm4lneYrQghBrPymD
WvmyR1o1EG6YNvkybFm0mpMeZ2ybILPHLpN9RV1tfKuylnGI5Gp5kf9PAjEGbvRJ
GjMHriGP9b/zoPPw6M5p7mD8ksw/Q+hO/Y3AHhimLBG8qLAGwT57SSgV9Qmyk6B6
CeXJIi5t3Xr1Gw6sWEe6/LLPYefh2k9d+MVjqndhY6FrOVcO/2XCiLaIJERg89wx
aLSDnhVPsBP7wuwoslz2GnrEPAVmCFgs7yBO3Watlcfuicjaox1cO7E++Pa/UubN
pntTAAVD6GNsoFC3Y3TrvUJABrUgYrVQ0RctUqIFXptxzzXrQR1Qug754LgWCXSu
GW6O06kYre2wN6w8MiSaLRfQVvl7/uyTBCSWn6G1frFT6VGbRQAhDq4oQWHbSKJW
MIAW8Y/IOQo496F3xbRqpl39KN/07fSD4g11xlJp07fwTFYsbTztWclzwXGRdJ7h
W9ugaLXquoEbMaack+cHYVAy/DaHkt1G4a+cYatMK5qRMdlkgdVzeHp4RTneKoQz
yOjCVMZUQh+PP6I1KtVXWm63rel1kLYLWo/BcJA/6B/UrUCTm8yg2w+D/K3K8RRw
rlNh2Mql45GYHfYBnNVYPLWWWH6d5plcy1oRlJao6BhDp8beeplNp/qRTpXPssEi
mWxx7MsBHhli/DhgEgKdS2Ln743l41/tx2Ih84E1NXSnRLN2Masu7/vt30ahhDPE
HNcoNRTBLaqtIMFrFhBBBkfySh/T/37aKIKb4TmnxJehpI8QJ1V78KhpnUmzeyIC
WrIAhrC0OgQCWIIPYiaNaw6SGDlnSa/4HRjqnW3aV6HKL9Ah/31eagCGTPzj320F
4nQDixLsd+BO8Tsgw5W23jYXsbiBlRx+QBiLK5EgSXXDJzVkfYnD+q/+agcGiea2
jBfrVDC63jaaUlWM7CEcmUmYn+Ege6d3/8Uuvr/IKLTo2q4erxLR4ycRUcHfmNf8
wabFntxH391Bg8xnvS5+lokION5KhdjqbabdGpG1Ebc14T7+vyRk/H0OWsK1lpN8
RUYRZJjevzaRtMOu8O7oqQvHH5yHj/AvIDBFLX2Ed7rHOewFSMaoUKUovq5FGj/F
Og2Z+Gxhddbl3r1lKF/LxXR+nssvZs085IhHS+j0c6d6GmAk+jnJ6aSggP1vdr6O
txKRnAd8VyBxVB+lJIw3ptiDTmpFKUQjIvMIh2ztt4ulWhV/76Ssr22aDy5kSpe0
8UQkLBp20HCJzUXO/tcBNerYa4ccOW/SICZvm7KmxcH8td4VtRSw9sabHDImpym7
EsuPnDqMByz7YTgzAOuEvakG63T4irx4IpwaIJKRnwaHTIeXmD0WNn+U/JtbLgWg
QC1h4R/5gOJ5V+VypiCCUdVTmW4F0URf+BNWHYzUEuLSzGEMmupJaZcaIaiwEeTt
O0PqhJfsEbeWZ0gBklRIxovAz3GSFz3P3FauyZFunTmAxmfT3/HyMZjzhnCsJaUM
2ZzaPB7BAJbH3ldSlzYZ9Lgvk6WoTpTdcBjlYY2PHjWra8eQ5uDCMk5TyA2/YSJg
6SFo3OSQr1q81wQnIaQsY1dbxUKBJ6/uyFlbMXLoDAN45lEL8aO1gLuqC9Zrb6tH
N2bM1QIPXkfVgu/t2IupxFpj/tWaNgLyW7oSnaB7k+/BEE9Ast21Trnz71fSeQB1
fbhptOlN2KxuN3MvAT6qIaabgHMrE/PflUQF490E+u6slxYtL6k3RJ5Ts4VCARVp
fW+xu+tftfna72iZ6qBy5ZlNfIYsKCNFTNKsGZQw+EHQPd8vkemsMkFpKaFBJz+r
xbX+wgOMhoxlTCd/YXTJctcPxCcv2dBEMBMcsui7LXeeUu7NRottOO55hL576A6S
JRAnKG3q/+1StHpbwtcVFyl67VvFKp0bD79g600m2MjTQmth80CjfDje7VODsWqP
gCH8Pv0bLluzYlfY8eWLtJpyKQtQsrvznwXvsDJHfXiEV9M/AcPBCcTsS8mShYMA
I+axgonSg32wwV6xSZldlW6uOwOOStxNrkU1haL/cfcq0+kXV0JMgx1s+49k85QY
+BwcrLm0UQQ6g3qfBM5EOSw2TBSPKPrMigQ4tAh4bXFQZ5bzCetfbexq/e0ujU8w
qFNRk3Al4Ff0DgapZ7TWvdzEfkcWVqOxIb5Nm82vHtGxmtW9QM93qcKTr7mqi4pm
RkQuiYrPlX5dw3srMLFSkSxKnaGGGY5rEXc4VeHcm9HsNEF4dczD4PJA0EXlvkSM
usikwyTT4Mgj2xFF+pJxl2JvDmpCVp7sEAZpGKCOA2vTJoK2GF4mavLTQ4UpjywL
bF03OMq4RaizD12M2HnNO/mCNLs3xqyBvjFvH68aEGfDI8txyVYRAVj5C+Tyf7wK
VTMshyUQAzm3KU1gpTptp/sb27VbAJT9ZEbtKJBN6abD66aJ9L5crImXE35IfBRQ
DxDWRcqZJZT7BSRF1U+O8NlmcRyjtadOjKSfWqAlbPxaLIUsfqwvv4tKvXP2j12J
zqo8eTxGbyGFZWQKUE0nbXEKc0srDHd15Hm9Gs6o0EADLYOPvQ4qm1TRV9PAa31/
9QKRE6USQf32Rr3PxVceS8GAPeS8/xX+N+sywyfUOP3asl/2G02YaFmf/sYnkOMc
a5OihZxBImYXKRymVkKo3d7AO2tuuzlwP1KRJW4mesT1JQ4fSfEKvntx8sMelv3o
eLdNiF6dfWm+KVrj7SjjWYgTqQWJh3M+2fHv4JEx7m3srY9fP0cuUfB5Y/6y8GvF
XLIyngffe8h6dgRZ1060ty9otbetu2ldxrBrg3vWPiKNmiBrTn6RtAm/omb7xGfj
vE/zkzxJPR78bhx/Lgun0MpMnXVHzM/bmELlrxTsOCSMXiSDz95aauI1YBsdAgkv
/IYVo5kpqkallGe4EBjLLUxMWaarev90wn2aw+BDHtAIZPtYXo8jPk4OxVqOIK+5
xmGZpmoBj+cqATp4ko6VC5tBCMNUNIEmEm0glym1fPvsEc4FS3AnMt3F+VR1Zt/y
Ajr73eYqbFrsubaJe6cO34K3GjMwqXWNcFE+6UxbvVUHX6UMf4K1TSbg4Sd1aLHN
bIP/ZTUlVhlbLoAyJVpu06g1ekf8N3PkBXs6Ga+acflZQ8eSJxwWUJ5VYRyvlfK1
Pi0SEcp6NED9BiCvEl3BetnEiL8p2jC5NP4TByjBUqEl64evwRaZz4Z04HHG7KH2
utE8Te+CkmB/x8lWdrv8OHxDC2MlOg1EXL1vY83ImJeJkjsqzB9Zs3oMe+JuVqpS
RUdTEJXD1LPdFtXEgC41R2Fd4joASQDMACQZQQnKVNRCQKCx3GXf5ObUuiVHQYlj
pvFBjZV7Tqx0aR/bQAqUcXkAj759f0DewAtgzXQnIpkpZ9LIiuXrOB0NYEkxy7/9
wqSIdd5yovie1Ym3452UvxQ0QO1Z5yAThsg993BqxBhs4+jg3U1pLUfBaV4hC9im
CNYNteU7fG8KX7VLPizMRr4KHv0X9goM8bh3eY16R+3OLkzHSuHgw38yL0XMos1d
2lTWCAJP6WIrJkrBz1U8/fe4Sxou1RBeqRnF3lA7xjBBcg/LAtTR2g5Hn3n1uqkz
94Cf1FtQJYsXcsyxBTHsxM/P38ZNY7Ir+H7XZT0f2VAa5gpHaLwTNmo9u2n5zSr+
XUs4D2z6Yz7icXFn1DRbaPDaCPjoNwb1HT4IlLhgpzdY5kqWboghEBoyP0O1RF6E
x2FG9+zvwljHNt3wfMiKCds0KroTc4EEvztl84w3bSQ5+4f8YifOgcPG7/YtdrAx
/rpt66PHyPgYtX1e/kV4AfyqYqIkN0lp1kWC5caEHB0b3+jITaq2f3h5/rjLvXdT
4al671z0iTu40tRTpIOeqTBw6w+gPHhZihmcWkn68whL4uhP/AUmvXTBol5+k7XH
WIWy4ZoVRlrBKRNCdHN4CEMA2leGvExFVcin0LLnuJtsNCpH7tl6OvDuBFpLrkd9
AKgFlTf7lTwlQBHHXHIUaBngUNFMbYfaIkhOmRRb2GtaRyxsF0sMvzMhuodwZW4Z
+K0STs9iupZYjAajZ1lL3ANOD7pu/1I54SjZsHp7AVuw8iGxpz0obpN7bXEEZDjL
iuk+lZ05LnfhVQ53VETz9Y5ws0ZQYBRBJzsf6HfWTSUxenz0T5KvaCFrbtg9mUt1
nI9Lnfmx8SPzhIadZSKnRXC3iXV9Np58DqiKtSkfta1m9riq7NxC3oUMMC6bufca
B7Om1Hgu9l5pwDMUp2EXEjHQ9O7CHTwh9hg2Hq3RgVdNPsHEpn37wqo+RztLyzKo
KMj9+f0yGAdXUIGIwIAe2AuemjBc9KRLDgC6EHvJc7qZzIhOQJyUDZtcNLQceCv+
9j5ZgqDxaWrfRH2behR7Bh4ATEyVSxz9zdqYQwTgW7CTY47r+VPcgoS2cAJxAlhL
aUT3W7Du6m3YzvEcomo1vzlMp7A2qehKC2la7RgkIowh9NmR9YrhtIceOkmsfuXA
tEPezoouwuVW8Gbtu65Hfm4JMLv2Py3QEy9Cw4517K6TcCTCXg7TTQm5DQ0NzLS4
tRBhMlm3lcLtIW9Nh9y/82fR95g8JSZNaAzG9oLxubUH+Lx+LOlz0bahyS9/JsKo
lIuNCLZO1UWiKiJoz3zsdCzjwP28n+42F4vwvoHgXgs7i+xepNOz0u25F08FARR5
gqiv2M2+voTPiMpFwoqGQWqvor8JSunIZn6yseXa93PWszyz5dfCiCphW2zm0/uO
UVp0rQdHpp44h5LxqqhRL14xAtsOWI3sM7mF0J/nu5zZtGkFlEiEy3GM6pDx6T9Z
R6xk3/b5XYHtwt5U2WJHfyEeDLxiXuL7ECEQnnqXsfNXNShc+RJCqu08O9FG7hV6
L09Os8EtgBcJxUs5n2/l9Tl7gT8DmLRt6hZ4Ktw7FZVcpT8iwbwN7AoysFsx3e+E
GetmeBcyDjiz+tnTuiBbyzglRuI+rrhfE78/fb3lI8xdE8c2cKY6DbH8FO0+AQnw
wiavOREwY7c4r7d+QHXQM1VvRrcXO44TzcvrNgtds0vc+Vfj9Dok9zSL/pkvV+DB
9W/9oXo/Iefye3RjUlljoKXW8YnsBG8vRQk2tdGFwI/zGlZLlQG4KOJNg0MA83d1
10Agp4jsox7NQt1+Wwpi4gC3u61Ozj5ch0XDefKzVB+SRztJUeu+mhpawbohLHux
hdgExM/z7VooVQMDArO5nEon78xqgP8HniWsI9O389goUR7pBMA7zczuiAsrNqcx
5otbbZbT3/1DmIqFHcpusBEZMtX/nv6l/rvugFgfJKe4UVJ+zrHENtMFd1XQVO9i
SWL0esqniOQt9eqXhtzWosE6FaIeCWYPsqWDM+BZlTcKxy9svdXLqicmOu8I6xM2
l5wVf4SUcyNk+Xe9r+gvLz8DtwjUsnD49MFm71b3y6TQAvtY9fNtQ0lB//du0oq9
us9sLopre72/bsYpwQJebhk/xH157vfnPGj5Fbb2Prm2vs9cYYm/x3YbcHYNQnlc
oDiPieSzcrjEwstoL0kx85p3cbEjZR4qQxxy74ChGod+9R/ig2tbqB6RKS27T+4j
GuDcRC/4eleccmtQU3VVHK6dAPL8frDHeGHfwRsH+M9kV9JQPWYmiafe3NmqndGx
+gHsS+Z76m5wxhid8rxklEJPv1E80KsJX76u13hPQ38YBR3tMXmyuLtR+xNnZZ6s
/frWCuve+hFslGpz97At1L2F1fVT1ov38JTF0JExaRvHX6dpt2OME0sxRg2PPF9V
bf1mA50QS4/uN+C5HduQokB8bucxzy2EBxGkFxV2luS0B9ekLpXuxEvoXvGzDTpq
9FBIgOx93mwfGXsSKnfLufl2QYA17DM0B4gekxRIjRd9EX45O/ieUvXNr8gFgYd3
LxricecghKSB/ZUfOMSdJNOxnZtedeY7UP5Nt+7k+a5cl6BeNYijrv77PhTImqKN
joPnsuFFzqI/bwOlq316U9EduovDr91i50Wfsyq+9/WYFcs4tdwYqIk/3oKCyAKX
Q8gtIUSsDbhTPJjeCVUUOuBpS+9pmWIHpdnEa6Yxe6Xg08NTP2swR/JZVUHQ3SaI
JEA6VJhDO8P0fX4ImQA/YEGnEn/HdaiHTkTF5C6Wt3gERl/Bj39D6zm++s01s/NS
pdq0K2BR8OtfAEpjyNC/CFzDoYbzCpa6guKol45QKcv3gRuUj7g77lJ7g6KXz+WX
nZBmBzksDDNDPXXaW9BXm9oFa03CjmSdwOsv52a9WUni6nNnpqXIsZkCcwsR6mcQ
/4067bZN2eFlQzXjNdiSLX46+gb+MGgW9gIpfRnpOemD/n7Ocu1GgiF+1D2mCTP8
CevzAN92y1AtoCM5XbkYBFrlkEV7cJh41Z8IVS/0Rdw8QgeIiIZdEklFA9CMDMsK
YiLfcZYCTiOHxjFD72IbeVTP2rFg21/8+3xajjmFkuclL57jKcaVdqNfJO4lTyTu
TJB8nyD6HMXfo1Uht6+dt3sy51rqEuCPY6mWjVQM/txugVP7cwtBU6+JQjrkcNzy
5zUB80tUAMi3g1/rkYjFbs6O0KJmpEP0j2a7341K5KozRSpjvd5iXgk+iQwOoRzy
4Cm3Q6O9Zvzphyh9cOYJ0N2D3KdgEdEVljixBWJsSFO41nrlXqfsaq4Zj03ybYBR
So+OKJyKBfue7MxilsHEHZoqwRVIqgn7KT4kvG4JuT0VN16REtTQNvx5QsPEw0rU
enWy33ozImja6D/5DuZ8k9xGdKintDZWxXwzdCsXc0pSwmUnljy9a1dQNjGd8fhO
Pc674gsH1DHw9po2PXeU5rSizxpiSAiZlhjUJU1X1tBTWnvGIsT4DE0QraHYt57B
NRWj+BH7jjBo+H+jbVJYnkBUp94CLQ2nJ8LAOf9hMqCTm5DwoKQavNrlOXE/iSfM
qebXBLzoklVo7uCmFmXqqL6IVWO7nmGx8p51ucy3LjjbRUrjjcRSSk3XW5pT6n6O
7XhWb9GliNlIIvxvZQ7JYrYQC5SuoLuJUNp1/2LH4IUbwws6SNQd5DUEcFSNMFhe
petMlDMD9H9cW7vY6W5bsjmckRn+yL5OOanWv3lZa8T0nBsE1/AQeAixTvcZeELf
e3SOTw/q1xLPKn+T1iTBXt/nc4Ku6VX9nccnOr4a8SnQXYgaNl1K1U8u1uL5aYps
g9AI0iJQkScHdNZlx5b55Lnixq/OtQ/oz1AF9Ci3B73Rk2uyUiPF9ib7pPDwGFIZ
5a6QepUN6IH4q/1Oma/Bdq2cV94bXABU3oI1ASrjBjNwzUYmkE+NJBzbT70qzDzj
5I/5tTiXXk3j7//5XLZ7tbw+eWSyS1EpCUct+kJjQYjUyN0p/hk9OHD3wk8sprQe
kYElMzULQnMwDx01LOCK54hY5mzVsUo/gFwVGfnYYvCsXGhyoOiH5LHbkuScnu1h
VeqYfu+/O610VCSVfKGYbJ/1tvqtQ9thG4IvB+7A0N58B2IB6Qs3F5Fkj3TQAiHV
iPNmImEcEQfwn8CIhqG+ZneqIt8A6shTy+JCLdP3y0/mDmddIW6b8qJuVXgKl2gP
kWfXRqPT66EqsQqFHlCsQW2RdhpWJUiCXBbwIWCeGeJtMIGHqlhLswziJfTHzX7q
cvDOP7uVL0grHXqS8Kwelu8MzEd/2nx8/+btRpRrri6o3p7PP8+Jy3rS5xWiAdU4
2X0N9ZmEiwhyEtEr+j2DEHmuWbzzBniWEE4W3OjYasHJchdSa2W0AYeaIX7bebuO
0AzgT3h/PUagj14rGfx88Iz+n+kTPvHszjFJt1xPimDAMvBk5TPpDxtrGKogfSlU
Vj7EYa8Rixmf6tKQorZaaru0v/9La7iWBia0mCJjfx4bi9V0B6P15nQe1K5/74Di
ejfjiR4MNhEjUOt6vA9AftyJpVNLdiS5h2xJOIKsu0wj1SRns/cxvHytELUpTieG
tV4OBWtQ0ahxDlWh4a6Q67OVmxMlCnBc25hIvT3uuGnSnvvDXus4oaaPg98xdjMp
kzAr30q6oNbJZ3BJBb5jKKq35FvVVBV1mAk9fKv37SZeI8cxwDvSAnNoE54xp21G
FGZlZRFzcMGzpbea1ShTD9vu+o6NaEcH3Vrhv1pod8qBw7bPe2bysPOmbyKcHcXE
ExdLRO6Z1A2FRAP20UIwOs5V82MFnjDtNrb9Yl5rg6zaETwyv2z2g6G0FLKmHpWk
/wG1PJgcU2+a+Mn7oVugwZ37lfv+KvMNK+KA/MCQ7flO4NMJiGTmEpxm3Gnd3lE1
l9ZnHqh4M/j3pKtcouMMfyKTKL9VvG3wun15qF/tUro9UrKteOr6hOqCtgeyW9PA
OwYdKigjUjd68upgB0xZLfrjsP1DhOljSF390Hhe0CLEdpwfTew4Ted8Htxk0hOw
f1eCmxgHIrwlK0+8u8+qXHtkqdTGrM7ALUs+pmCpN4lR+CUrqioo/f9/m2lg3CoF
e/uEFs/pfcEGYoiNJIvG/i+m1WhSJ5ekVu2Yr+Avxa0UHm88Jncz5U3FCrxBdX8z
qQPtsJkhNWHkNEM6OGLPuMrAVM0Gba3TEVg1eb5U4zNMpbvJymfVjX9dPvdE1Rwe
f9OeXgkRjcyaytLfl52ga4ZzDHNkMfaEBq70jPV4qm66ggCgKUv/IojTkshfW1Vg
/Y+hTKHOSvYujN4xUoy9sACfuGZsePEd33h3dBMIwtBr/jE5bsy7T1hEiK8oc4ZP
oMemcj+CdW+tq3IRe30iqh5g/iUJirVea9gL8Dz2dC4Srt18k3UY4lPd7OSbOiKj
ZapJgEG4mLi45JxC5VQrdrdtmTBcjpH0AlE8cUq4df83KOXnaDzm28uN9GtpoeaK
ulVsTDa0rBOjHv0RObesTN6wUEjj1bH+zhYOFxqHgkuT8hgLrxnuxZ9SUzZX0HFV
oIRd4tffQ0ZHCZFhIVykfSEcxdvBXReCmNP12fD+SC5b0VR+XeXbUOGYO1Qz9SES
bIVaqNA+VhuYDf8nbwjT50vlitF4WNZdPThG9R1sQg1zb7nbpU5qXRrZ/qL4d+cd
HL9yWVplqr9BWgNBDd70apJbdAhu8VNisTgahJEmuDXj7CDHyWXUMatbf66c/DaN
f3ShhkKCuzFPbN//j8iCz25mgK1WeaKfmTLroyrsIimgbjuFkdRCur63vEesXVkh
7fobOIPy7g/746V5WZx4wIt0eHGNuWSZLJq3Od8n3GH3jpCZu47k3xys5z+N259I
Jz9E6HGiJiSdosncGGRytYfT3t2w9znDDwJtJAdY2YiuU8LVwZwJP5l3J9D7bZqa
h7lrwIdSPVL0BkSER9iW54/LZ5YkRfjhqcO6UYuI4/RTOuxfikn+8rVd/7CR6XZJ
YegHJKG9aR4Oyi7iFMi3woeLzpzI7swPi4J2f2DJELlYYyhqk7QzYyLDCnruWUn4
yw+U/sw/XzRGWiaEu2qD0q9BWXAh5QiWE0EzOGkNKfdHUmS9qLz/F2719C8r6sF2
e3fsNyuCO8EGX9P4iow424u0vO+x37eQMbTUAvV/cyR2mw+9ABmI491sefvLHww9
RsSSNwmJu0nYGSQQ9CHt7+9/0Ho2K/wCg6pBi/o5t9b+Jlx7J/FHh2QAvZk5KPAC
49yNkifI8Nxt4fXjGkPpDxqXxbvwJVictl71zUSgLWChavcOJ+fmSCnoRKAOMrxX
YkfU8yv4BGCiLRdiaR73k9wplVE0WYsEaSq6YlUMIbWQWZKtWN/nWfWxTEySn2EM
qD8XGHQ99SDhH/o0Vg9tYDPel+fbw22eScEQBjiYeLDSblbl0eSSF5r4A20FBclq
pzUmKpvY4CDapFgiRgu27u2ahbypXLa6Bsm2/uJyismk4wMW5jSRcztvzLx1BUuu
RWmTG3YWnjKljfrLUzKvt5bxJ94Ltyg/H168P0hbEiE5BXEgqUD6HRAAvkOulUAI
QUyNj9sIYH0cRD8UUTtjkjECPgyV2XTI0q93lZBT2z0vhXEe/kXAXj13j2O0fys5
vbrlV4xdxvJLIGYvUUtFWYKJ4b9NAQcD92ZNyYrkbzRVkxsb8HpmTsPMLze1Ruop
LqWke/zPpLmaCs0C3A3AIT9EE4wE1QMZqEkCbPHnB13bUvW+83p81OgwmWe3yfI0
8/2J1EJQ/f6D3J5Gl2RlnyTR5eAc2Ht8ekAuSov15BxgZTdEYyoILRhAAvHT5Hy/
ZElJGvGHlrAAK/VS8I0hcP9c+UThis3jejPqEMboOT0gryrYKymJ7UdAtjL0rcsl
5Veky8cDt6vD6T0syZLhY+8v1p18g9fkeoyLXpCdQ2uPOxENQ3iu84TW64x+Q5ih
hVpa0IJJzeGtdgwAU386ibM1cd2pRtBozvH2okfSKqccmJH2nnzyZvS6skcTMiDq
/t0lG4f0oYdeGDyLvEfFx0ObCIN7D9BxoeltHY8dO9p7qXSUs1/WbSCLTaZfLqnr
Kck+ht9s5pnT0FUsY9KdgHn5u7otVZTdapGxwrMidYlYubvaHUdS1O/2fbHQAPw6
OL+kLruWihGjXX0OXhnNpVdGAJlrlAsDcK8yjLvWeTlq6+D2+F49p9Ohxi7USkTW
ZnrnXSzaF/dbab4iyzRLa7cYY6nlyVicNP+oml3okbS1kEwSOhAUZ8KtDKdZi2KZ
z9zHWT+1Ky9TsrGLbdv+vo80L4F5NCAMsxIBzOwIabw4Lrfiz9JvghmwSOXESkU/
BGytEPVQUVdcWkp/Yf4NQ94aN6VZU9v2ll/fr7j6d660DmPQ2dnk42OcaIBpHQrX
yjU0t4o9YjBvQj7/YuOnK3pPq2jpKSU3TYP0GvQhT36csKsHWbvF73gfw2LeUkDp
1H5O9ca4wYDdSYpESEfFfsRjEy7sBOBTln6j9GjgHQwFZYkTrl8+uSRV4iE3MLdK
xvM6Z0goP0OHI9Kr8OPJP2AXOovbMraOc0tMOv0aHmqZXTLGVk+OptRMoQJqIwSF
aToMn9GDYZnJnXPuGbP39kKi6eASv4R/ANbOhQFRPYkDl1wKgNsMkKRlhbKMP0ck
1pFPx2X6Sd4DpkiGTPNStLpCCSxYQ6wSkt0BYs7LoxgOzAHyYPWrawVMUxwbFWvP
6KKbE2TvNArN6gTbq25fgHlrWH2c69Y/S+H+ht5Z+kgxq6uy+l3zGVthV4jxhqjr
jIaiZH+DI0RQqelmpqo/D+cr7mqWDwKQ2yc7rf7tr4GxVREMOBC/6R2lIgQc6G58
N6Orcg9jqi7rG1/yVO4ihxoPPVGkBKT0GMSv89KJKsrDQjlRu+CW8OVibZ+UqHHQ
HdNBa1kU4kIoyk8pC6yV6ReTqakzQY1dF4tLYmebLUWHH8Yv0lJcu9XN8RJLUwyU
ZQlQn+ClvSSjTKrj0W5Ci6KgKM5M8/V0vQcIfvQNWMeiSU59Hi2VgJv3yxldTXyl
ysUH1uylCJFKo6f74Arg5nJIt3tDvMTlnYSEzKZ6qgZmqyEc1n8E5hNbVLfJDUMI
UQrwopQWTZcFKlNi7pG+TWHZPf2YjTHdHGcJsU7Haof6eAsGDVWNf2KDIejBZMOt
y5AZAvQectalMDqmBw95Axgeg+b68ZVLHBfJB6sQNZbXxiIyqMO225/KS1lO8j6U
CKwIMfu5TF467YEV4EYrLiOZ7WEBtrFrEB93DHHuEV/SsOM1Vg4nxLPX/HKpl+tl
ywEA/VbGVn5ASZGVx1aUnnuD/XPAWfVaGK5rId/80UeSqxcuZh7hefWzRt+MyBUO
MPggOZUpiNdSAbi94wnpVoZKbDjC5pWTzxRJEkTyHJ8AJqXMSxF/zdtsshavljJz
ZukZxKEQGUpqyvTaqVX6XVjN8Sms6hHjHucvWdQ4O/Lvtdrp3xMWGR8T1DHKoQpE
9dbmZk8su/zSBsrMiC62IVHMg6/oy92NpNY5gjzUsz/5L9vvYfw1sfymHmdWsGtT
BF2WuWT2N6EEP8ElvZn4kkSWSKxFJ8kX6hb3CZR5QbmmBuVnXAKKbSuLDuzueard
ECdHM62B6/JglRcPXqiU1T4yBWDCSNmWSL60wQc2lRDbyG1wBVBGSrrJaHNDDID3
3307AdSHg0Hcqjv4F8KEDDOWz9F7A3unQbb+JSYv0fzRW8qoa3UCTbVltIvVp8/A
qCtt8r1LJXO8RlY+M+1lq8651XjLyhkKPzeLtxl5OyRjTxPos5lnsESCF/VgfLAo
3ewlMVf6zbeycK31bBj5DCKqBRG0KTxRKMNF5bNrvrvVs/OtdkLmIoiPOvFkqKrY
RDdIZq5+7bci0gWN6ljokLCcUulb73fKYTRGK3LdCpJZh9SuLFGa9WfB6c3vqiP/
29Dyho5D1sIOutvW9hEBM6aMVzv0j6ICHm2s6yKeN/HHzx17M/ALRVU53T9ZlT98
UwlthX9vzD6yS4w7XLZEg1B6BdZ0I+lgP5jTtD7zL7h7gPfJkdSHYd0WJ8fzHv/F
MszS+Q0dQu8eMAOrhbz5X+/5/0xY0M3GgZlh+qYr1wkTnmZvjpCiD/Y7QvKVPeSD
I6YR61NtrskYY5VCfUIpcft10b9ZYwhUvd0eOTVacYo9L+JJu0iX2+047ivoCdPR
3oKF7/m9ZYpy4nmG4dc9dgFimnGlNBReCGzboTyP77LFFF3osVA9qxR12+WOsUpE
x1le20pAEgb7Y5Nrkm+N96ZR2NEBIxEs6XfJDJJPTR0L4Wclwou6VIhiQwHY6etk
zCZXH+rlHli0I1MY6aTxcxa3iB1yFo0APFSFSnLfWTZ9MWdDl4PGFnFhQrZ25eQI
oD2MgebZ/8YWeS/L/rEMJlLq/VDukQiLBjW6tz0F2kIl+Cvvsfudu1qiM5l71G32
sKuGTQ01BtzZL26fr4AhcHStX+mtuFLjY9ogzBNc3eXPWoQE2cc/pgqEkGAS+Kt6
q1kaLkLbyH+TWZmxRaGZxHJniGxC5TN2PiB7oFq/GO8GW9i0eb23pzVn8aYep37S
leUIVkZwg9eoxSW1KmeAvcwcWbVDN9xCRweK9RECCHEqmh1BXmY6qu31WFFsi7xi
r/UGeIdceJrrHwESpNRe9Sg9wFDyNvQlTHB1k+C/nhiwrBclxQdYzbyxPfvQzUR9
rBYwSrK2VkcdOpOStwLE9xqbmRIrdssBIvp7zdn7EboZR5dCg1C46aRaFMMqv1hY
PAX8u8eteQAXf0RFodWZlGYZdPKVZestEy64EiBwJdhO1V2SWZJAq9LwoXaLTeWX
JijHn/jWpTFbEMmsKTzDgtbhC3L3ha6fnSGxn02p/eyEAQUzchKN13d3e2ASCctk
XmJGB3xzxtI+pumqhCj21IJq+hfJVnX+qQr3ZaHI0vVgllRrLzOO5nL3zwbLPmPG
aDY4Hdp+x66mriFoA0yzcwWUsb2PIVZiH4J25Z6Qd2XPpDFwUtIw72SdYt0rb1Ff
7Vxgc4GDOfVnLxBQQCvR2XwfSSRSK6AlOamh8t5L9VcNOTf+b2d9micyU3tI/pSu
XZDMHm026qF5xN1o6O9iF/OgDvH8ci6hIoPQjMXyIZ5Ifh6AuFQ3X2XyW9ni/U96
ycCBURc75UACWGve8gx0ytI5UG6ATMEdVaZL84RijjpaZP54WRs8Fx8GcXBMifay
rSfpnUOWq/tHi3oLcoGGqYLYY2suoSpXUfBXQ3RL6TZquDnpthwJsSnq9TCZ9Ryn
bTrcEWCaFFogqOe3EsUVlNMRbF/5TThK/ciFz3wbqsVKZy68YBMG9xvD52eHJERL
ma0sdJAECkA5alFCXCR93kauhqH0G6Z7pMj8Wli1S+pZF1doCwdFUKUBIJcGjKfF
FdiEX3Hi+SKgs0dQYLzW0BPLcWoIve/ItsbZKJkTW+gVx5/WHVSVyRFeGDo+vcNQ
Xbh7ajT0IweOxnuPk75ZvAnJzLoX+rWMgMYodYU3h9oE/pfqvG2uAAzId+vGSG0w
XXcTP3CR9clTrzns4fetKYJCGgLsE8kVK6mHD+plGYoyUpUpZKvHmgCSsFJMKMD0
tha39SO4lhnCvfV+aLVqgjm59RxtBm5l1Fb5Z0CdgXY4Wf0Vk2m5M6dLQxw1yi8u
rqUJ76zKJ6N2Zvur+iBPJ6HV3zraNT2XiZN5MaprYFecs9BTwyI82iZRAtUs3tha
YebXIv0XwP9+Dr1ygKWuyQMRigI0IakGFTwDx1BigwG7P/qy0pToe6FhxrPcI36q
eZEm223kReQpAPreaDs69ZOyOJw0YrALC0ZpPtOqvQ2FHSybJhujCO9EFq2WMbeH
ETAKxcxVinh2zD5f4Pga8NkSlQ1pMLAldz3ZX4sKjsbn+kaRYPlrvP5ZmcgIyv35
flO9OVvbslNndH5kAJ6WZ4FurJLghi/8G+4KWkk/0CxHmELys9vqmOQo7m5e8Mys
6in0eXa3o7uPDQSoHgBm7Lm0eEgZGhRs+XPLc7/aTst7mTsL330lx3fQyeaq8JTm
XtbXdzTSsjszTjzhziwvnOpy3wm4lxsz4JIPV7JqCXCb8TjVWR9igSCVOVszxyE8
ED+f66MHgxMwND2K4IT7U6ssXROHhIqha/IxtJtpqDMwVwaE6Pw9lX7ZDWD6fF5+
cgVl8MYKUzJ2x4cU/L/M3HqheEVkBp0AI3096pJrUs4rNvNAfIG8nudMiA2mkYo5
TjzSP72aCPLXUfu3h9nAoKq0zDr7I4s6TdDX7W9512FtahV8NxJPmnj5FqnAYHwc
89TrFwff5V7MiNX/C35nqAyVCjxZAFKl6DID8cCULe63eq0Rpjs4rkabnyZy2+mR
5C8/2GTGDXDQpMzRebxHkmCJS9yiCVHwe5KtLLP442bdfo4cpZzT/vaHHK5156aV
XBjM3IJujc6Ypuyj1ssdqEGVazKK0wc2Gd0ljnPfoa4rc7fQIktCEJozAIl2qZU+
9iae28S5FcDnK1f9f+04Tz+elivNKNwBO0RRYtTCybQPSQO65dR24I3iA10o1rNB
zDBSykhc6EV56xLoBt9hxgJ1VpuSIvAQR2X/NoFUXml+HLCZzbJvLZFUsBhe56ic
AYMYlJqDp8bbVUte9+AHWtdA9avIFuuqgz1avNtODU6ySjOwr/qGgf2pYTODOoG2
e9uomA5M1OKf6zpXnE9Tj2phyaYn6wMnz7iRXOU1aOBVWDVJI5pif+uzB9l/TUYC
xsR1OLy2IzxY0kjOYJLtc5BlB447B4Kqe2UP+ink2Er7DkmHBVNO1yD7MiG/yARf
NvWogKcYzFDWTlQND7tsNzRuIBZn2gA0nOypXt5JbClxmOT0PlzB9+qUwlAs84r3
o5W4eKMNYaUK06/Wb5onPmtMd6Tqh/YnXs2fd6kujw5595/MuTS0q/SSHupQw4Qg
PSylsCDYOMHBMYvU3K2S0LEABwmreE29o/ErBg7zgyVzd9Aiie7Sy5PPytQC2lM2
wc5RUdI1mY1EyZm3184bASoMFfxQejt2PjL03Y8n+8Bl7ZSc6Nq4p8XaHsCsy0YW
Y7Ma5tttlqdWlzdA59Z0TD2zrRp1KRuEyeq8nmygyc4KEiSryxukEx0P/MCBUfW0
vYFAJY3OTrau60Pn02FePKcQDZj3bLPyIpKyshENkG4tMgYkrEsn67tQmiildXOT
fpBtvCD4O5P8TqZ9qgrOeNOEbu7hFmlq+pExLZSEK3y/IZ/QFqTHhbSl+m3e6AJ8
gwRSzwZ/d079hPkODoGANIizZl43Y6uHW5H3yIJet5KiVoRI8xXIcZzEK5ImG/q6
72ICfuK6T7+QC73y8/33ka9f0Eui39u61MIpleQovYFPRf8fa50LMXAnaoB7sGtd
noyyyafmg+FBKdwy6lhEP759uJf1vha9n8KVetrh6RNB8IVqpkF+xu1cyd9hOXtS
1L8nR2sXqMEJrJB7onSjihgjES3zPfN3L75P6POcCsaiSOaEUZuZQTaA/yQZsfVZ
1p2v+IR4C/RlnDBRyaYQ270KRjVLaqL+W8mEFX558vSYMPvZjtUUPLPUNa8o25ju
DPmkK+GPhWiym4KsxzShgEn8AnJ1lPHMEIRgvBCpur3MyYD+tPPfiYjOZNVc6wvp
X2Dq1vx3TO8bgpwXELUX6BN0wmUywacVxhfJsSHFtN+OpR+aBFkiJMHMussSNagy
OMx2avsrw8pg0JqKjlax5T7A50zRi6wtPb0iueqUd5zaL9u4Rwx9fef+nMGx0UPq
amidX7QOO1FZAX8Qof7GfAl0JKvHv6oM3DnFPcN5Ld4PNw21NyGG5UzNAPUvqMdU
JuvDgL6gXozXz11PFUyDJMtneqzEmwud0MzGuCxhIE5DRdZgCVm5Gz+Jqbol57zw
fAyRdjozd5LXYh2Enr7g2gAOHI5eappcCvQ5ep9Hu0Tvhbzed1+Xla2kAtNIAVW1
MrDqvWs4ydoCz36/Z1a6Y476q0AAKjaqVLsaMEAzZkvzZ0XIC91vadJudPbteNGD
H8zPocOIm0RqHSjNE1P8ONNJOfEki1timV9Pu6rhHm+VltWUVPt2ryXQgwTpx+Eb
tK8EXBefIzSKaTDTj9htTCfNymSnYcaga4otcqGPKRVWdxpRBxbS0iII6S1YsaOH
YW+fdbqQU//e/f63Cq2Zb6bovq5whmn2aoMYKAb2sMGmT2K8HKzybycB7yRIXR2t
Lo2PpGInFqdQjWvpkRE7a2mdcygeKIQVJqDjd+tSqTaLGztKk/K+RC+Dn0d9qS/G
GTsd4bR52vLDGrnogI3SU7cP34f2f9SuF8xtjq4Df7maIEfvcCyHX6zXhj8wyWAE
Uq7wMQ84BeKGoLRCyqcwW5IUeAFRYGr9xXgeSHh8NsU7Smhm9wUghYFParMFYnME
W0nbG8hVamz/VlCAgVXujugUFJt13DocPrY0LTlos2PIJTjjz6JmvRyK91xT5wsH
FA3geOG0Mk75K7Qnz4egVyYOosmJD8IJVVwB6Zz1cL6qjng1GJbxykn71ye4UCP3
TGuyuDlyKLphEp4ospKRjwSJZxFAhmjQ2ZJaRn1jJjMyXspBdVNWZr2mriE2wl86
MpBSQRxw35RacUN9wiRyu7bHyg3l9pLtyt4/SV8FaoVYexXNhW683tKq/cX4chkd
3NWDbFRjjC+ZgQO77qAaOVkme/8QyTNz4THpIa3JbcntA9Sy1FkdwJwfzjs7W8eq
FQTGrEaWZOvciekFcU31xdyg+4c/IbVxO8ObC7q+0EDMkf7dhyzEKBfbVUPQrcSe
QLdgKRxOmO17XotM/4Q3VCIZ520Pay0WgL48pNBqVDe/oEIIzZ+pYQDMi3AEdzGv
JKXQ+Kf2zG3DTXiCWWcgyRPed1juYdxJHQU9Jb9qEWNOkxAjwCdq8oOYAvRZAHhx
vPpvuSP8kg2ZPlzHXbUAxt0IztKx25Fj98kOP6aiQtPUX05RM163v0L8CKEGnhMA
Tl94Q20chKhtkgDyVGzdqRi5LsMKkYdinFrJeBtBtJCH/UrMOEqK9Ph0cRJF5rnS
FUEQhp73EGrndxzrc8duzahlUXFVbACSZ9qNZaZ0GywVcxCx7l2Lf/y0EA6EG/rW
L7jM6PwMXGPG/BT7ehLdVfi+aOc06QjEJ8JQjosLIIP4B+OpwzblCqbVPZ8yDgpg
GKg+KX8hs9Y9RdybdTsmvRc+oATVWfbT79PnpH1Gv/qopu1Vg/Y3deqghbQw2YCk
QLqZfzHk49AO5m3keN1gbC5K32D5o0DZTKBCSHKm4W9EvXP698yoo+DXR5+x5KG/
WIxHNxWg7cUczvUDlO9ENlDJQpe6L3oVK92uVpJV+YYh8mjM323f7CeCedSoUTKg
F8wIhP+sth9xzzu127KaXr8A2sqSNnBGFVEauZl3QB7lrSPgUzmNFmkKOIOret7G
6B8M+MIUeTB6RyXdRfiUqpJPIMSirb+WLur4mCTULxhSPgQI2JIVIKHzzwL5J3HS
AjaF/qGSwp8M+4xwSTUVJVtJC8KR4NxWm/v8jIb7VNYwuVAKYc9owUj+psGZHrqJ
uQxOnr3XoYaQGd4OMRbzr3PofAxZCMV5opQoFKJA99ua/Ic86mIa5xG9JeLQ1pAI
aNBlxbRcFzzTX/wEM01d3CLi3h+DIvDZ7JEhfMjk0/Txwk7TGT50jDO10jpUFZD/
bLFwi9SAYr5K6dR3cfoC+uPvodhs1ebjSY6jKIRK6VJUkRqfW+9+rmuI7HPg1usj
HIg9c+b+WygS3mMY3+nokcldS/fEfN/OtI6U2U2htX2Hjzbo2gUfLfnkjtluGSpo
lbJGTKEjQVq/Z6y8K0vhmnlQfYzh/H46PSGYfiKQxXuBlBa/V1bvBD+BibL6fbRk
f1K+c1W8o0ubY7K82ldf+WgZ77+nRz0qVPXUhJ3EH3Peh3AxlFTLRcPVUppQiTNW
AM3YKJmNQkQfPLRV6slkpbbo0qAG+a9MGZ+Z2o5sTCkLyUdeFNHIHDZMF5TFPa8z
QXrfH11Rjv2UQDnLsGxvWB3lV7CPYEBDLebFJ1uEYPmnYYh5yKj4wMC3pbOAGgWH
wRIqZM9s+EqHwLex83ip0DRRLNZOdrIQyqQIUxKc+vk2GgBluDGIQ6R+u3A4n3Za
UP5OHO8uPW8XoWGYkNZhuO7a4oNLTFSW6AgIrKUIxoCW1H6yrHFYivW5QNlUCRsD
62IcqOs1ZfxAAKy2n1RAP2SKx1RWg5NZQ5qiOwnP4bjak6e3XGDMo5funbsC7o2z
IIjARPHvZw/2QbySntYI7CjjyozE3aAahLE/Awog1n0C8pGXPiK8o6ebNZDYligy
NMd9g9cOuC+szPjjdMKzz2s4SCSL09thyDuXpzOTqxGRe++PQ/U2QYP2mm6Rl3Rp
jx58p9W26tFUePRA9/lrabs6KosV3QOfFyQR42C360c4PPloG5c6qbzQ4327v/sh
2a8jMFRQ23KGMNbl1V7GVrWyPJfTFWszwpGw6gBkQv80GvHkJLstv690jEaFVoQy
eyyaoHk3IMSgC6h6ahinEYO96YiJBszvlgkoz0XP9hKfU3N2X2miRpXZDMrsuGPy
Wa3ir//N/6TY2a+KR7e3xcmNd1URWAsyrqi7LMK/BnQp6c8zooX5/SE+5dM5WXR/
rcC3lWSpn4DUy596dLt9s8RS5hk1fyZfZtmvHS/I+gWLuAu3FGHbdutc3RH3MZyA
bp17hTFCJDA0rVPKMXS6W2QR6wwbCiqPaIm3lRWdlA/xl/H+rHrVTehHxgozfYpj
NbA8GLZyEecuxnbsLyu+6Oy1afwIcvnIbHk/HdM8U7qqSEqamwEXuijbrL8PmwCd
VUx3eBbx/8rdzMVh6HyqMBMxGzIOZ0mh5SJ2U7z37H9THwrZpEfbDQkFh57gY86z
DwwlDRqrwqyOzzC+Jrvx2/iVCLznbZNPymzJhCSOUgKvs8W2Y+J9+pzML7WXEQfl
+yyj9JBEnAfCFTNZ0usvg5cDIjqFWI7wdZ0cE1CXL1NYaUBXFsXlu6cpxSXB36V9
nBrVPgokIfspukvFxtQx0/YXPXX05SwUyampDEdvbErNkBc1WaKnJmhJp9FkLeV3
QOeRtU5XdIz/8J1elUpJORZdyPy37JN6g0W7wfT+qrIUwswRzQ+5Pq4Gb/yPgfCv
EQnoHCJwZCGtAyzodLPexyMZhOlaxI3ysWkvzflJMEgDNGxx9nzsM15ZRpR2/Pxe
PCVaM7RaNng2/PjHg9bfN3PJeG5+zS/F4UHMNa8HYiNlm4KDy82TA1e66e5TabtK
UWfGYRvJDVvYfm1sekONGYcNsckExH5Qv5r9kTu+QCHmsC+iSvVSIQI/gFvcLi22
PATlOOkWGUUHEyuDHzJDeUvXKUx91D3yPBb/q+cwRlDu9yD5qrbnIVARh03GjwsB
JuNzh2j4NA3bqy7YfpR1uOjIOyJX14X7JMAr2l9usHZ6K0bYc5yfvuM7NHMEhilD
CwWQ4N/2CWbi1SrOeyVQd7N8eh1y4Ur+irO4FmwV/RCophC0vbbpHyRu0RyZr2yq
47MJyS0JPJYzMe6BucO4SSUmXoYpgh88F6LqarMBRbKAIVl+fBOlnPRw7VjxV/C9
C9DjSp4cPGwoq0wV34RYT41kz8dFCaCQh8LfxdI1lr0UHL//H2pfgRex6+waiaZ2
8Vfa5hoYs4VIVp3ef9M9P7IhgM8YI1wGf/o3vnApzqHTesn1z/sC5P0aVGjVopzp
U9FdXMnjiYwRJVq+2g8x95Cb+YzpMBEJIUyaxVoAE737F5ldP6sCAX92NEm+5Tgw
+RLJMu/9D85S4XxXDBG1d2/yoVwTPeA0HnysUb4kuySx0EM/1QuowKgy0Ux/EMkQ
Izoic/wavocwWQfOOauFCp5uSn5Lr1pCEv5O47FdBgp3Y/9+YknQlVkYSslVWMv9
anVgiBfGq8Cg/H/ysiG9LMIbxTzc8v+OV9KMEgQKt+9aL2nEFM6EEXqJ8eMqIlfC
sYFQfrQJ9e+ka0f2FneTH8RnXgAGddC7kjkWMT09SoyH4yX1LrGtDteUVLTln88F
6FvyjNoDhGBXU7sp+nks/e1p0o++at/ieLg0xnFbSUT/oxsgb9Lp96wPWVn1MXWR
ZRO2nqdQbZv2FU+5Q2kGlfu5Ezkvm+cTQtitNModPcU+xtHcnltGH9XEag3DKZvG
UIaedCczXdiL1i0J1mN8mlCwTlB+bcCpAABY0NSnBMER7vm0TpHtZjaVgynxHpIS
HW9lQhzcIpUJ9SEOZJCQ5lmy5aZJuwZLOGLIw4XHZ7Lu2v1nVPvth6Q1Y4FuCq5a
63qWjXUdK99zkMY0wUA/xNtyB6CNwXFgKs7atf0VnOHFEFDXeWjXWlWnSpd6MoHB
F4VBsWCHOPQ+AZ2jPgAlQ28QQ/z9eR8SrRDIaVH0gLVaVlXOfksslDwSJEaxs01r
0TTSkhqnvDoFn0D3ecECRzLnDV+/29I7AP+bAcg7cHN54CO8iV1dZq+xpZu0KpgH
c0dF6U1Oouqclr4G6giR+gHAzCoZech7947OpNO6vAm5HL1Oxi2YyaKRjPfedPzI
MJzo2M9ZFiDqeBuPrSSM4dzpqgWgApigB8YEzwnQnDAqQk5KjMIs5ctgZVrcmy/L
OJ1bgOk7WcV4rPtv/sBpzFM8Alh67aeAlTYoKrKDIinOvgXXRmLtNRJVUTnwDau9
6URGzfBOHtPsGfZ+DgcLfjt7MG3lkgRnnamWmiGX9TiF1b3pM1rfSb7hj6I6XcRW
i9xEuUiPts5UYpMXSoRg1yihbBMNaRumoiiXMKZNOUOsXPYCoda4gljSWjraRqnK
UWTRyOdiMDhWK9g1miopAv5v0LDAmRrUGNzrXzleBKU4ciuAh9imUmbPI2A9Nczv
zHPBwB0DYWjLQagixRGkJkBNhbWgCKE8MeOmaYcGUPqAUZkQM7HY6gDpEC3kwaWZ
1GbVsncNhI5q02g/eCy25GXN8u3rhCdks+7WJfFiaASKaT1M8gLvJYBYCrw990+Y
GrtS0JfKK7MNw3ow3RtNzT1kiIFL2l4X0ZojpwTMZOLS1h5ybFQSkoSjo6d9zHzU
lEpcfceTfQO10rlaX9QV3QxyIdL4GsqqCAPIbSGDHKEjCHVrRchXIzBX64gaI9D1
0Q863F/VRpUkcVYB/bbbedPWVdyuMQoldPmuQ3+ZvSEzCZ+INsVWakQATrDfOPur
fizny2dv6l2Reuna05FTL9r71hWRLv76ctE47HHrbkK3zRsH+5usMQJrE7hLWIVB
vxYGWT4fkxvRlt7mqYC+KP9JFHv8angy9EXLU88v/RSeRig+N1zYnPD7/zF0aAK6
oj8ZVVzn7ohlrnzFMajG72mx03AQlWkuQ3y1SW3kHn7plg+9rlJcCOzG4SM7cWTR
oUQ/Lbl9ECi8Le1wJiYgaD2cZRkzdAsMH/IN0SBLVFWi3d9eHLYz/bxejUxksUmC
qjmFQyFZXUw538W5Qj4io0UNZlaIlsd32BkNLwXq5j5hgmoMf0TsELJmdwhUTF/k
80E+lEqjWSuvEjlhp8qtH/DdW4Rg9sD1/K7ygIF0YV3VvchkdC5rz7sWCVwHyJGv
H4S6x7N9LtU2kgaF5B0OYTSFcBGDZ0732uh2y983l1hv1nPdA5Sw0svSoYfRU5sr
e9fDqPHVsTvLZ9cQUa2y4M7/SFTyeCGLKZjKFABz7LlFURqVf7dpmGJPN+7a9GcK
ZdY1IM5rOUdN47iEWrqVzDm94m4MNzDmgmTd9TJuyoglNByaww6dS7h9PtxGcmA9
5QYiaYKJRGtaA/Cqk8N/wKhqVub2gxYj95qusMsqVwBzNhClIA/cCa7O9UpvzLDi
YgZdFaw2FgHRyuKVTuG4eBqTi4AXIF37cOa1MdEVLxJ6KsZnk51NBqN4yDmRTf+Z
Ll8t0rAfCf5PPXS9OHk3/wPFsMNbKxSkpAo1z8/EY5CEqKnSkcKMe4XurLLtdRG4
oyIqO0W0qlmIJMRReaoChB60455WYtDXdc5Rj/on3E/LLiG5zwm2FPcLRb1yWlT4
3jqh4kHNeW/RfdYblxa/cCstqdNagcoFMS/csZDcfALOkrJKmfZnHkeWk0xvEp21
ytwaB5Q+hCHwWfRcn68smeWE0nuJYHZ+gb+TDlYOphbiDjF94JJnpZw0V5IOPIby
tEFt6izLgVItkivKkDxncGok3fMRne6paY61WTUanqQvhZnUk632/t5CVPnRwwBy
0p5XkaBx95P4FrLbcI4bNEHv2Q1ewyZIcAb13w6tmAkCkU8JEOn+7TeY+2A2jIYK
O3HVG2a8SsdIHHz2xb5GbxBBFbGqUf+C6RvbW+u49ehIc+vC+QpnywZgp2y4XE69
F2fNkWTW2uJvnmhZynWDKM4nvfVdwnTMD1S/pSVzctu0woAb3jPTAf6QGtR5RIjF
TpXZsZvjINMRbVvALUIVy+pcTtJscqgHXI1VSG9Egqvw5kTUUTuCz2iPzdIzJ7GI
6pILDPQRss9DbU8zbFx2cRDHEs5SIQdyM8sysPC1jf+uYuqh0JdfJnAm3Ct0Hl15
hEqVl1yCKSMtrfYwWupX5ZL03/hKnrhjr+i7En4SEcIlbtn7FS002vA3SP4QaxuZ
YTRudpMXwvgummPfCAj2i7E6fPIJMmuXy2TRLmPsVchSbpUqcf+BBEXuRJrzUeRf
m/UGeBSJ4a8asHaJ1t6UxKqVyHQGfuzcLCVty1hpaM/qcnnlrALR2fkRXGiHz7EI
zfyd/yOW3ydcKdfC/85zP8ZNDD/B4NNY3TTIfZzJYBkl13qRYdp2+JptnHGsqbxQ
s5wB4bSLCGzQEJVk5HM8WRcPeDOew869HyWKenlo2ZWNWk1Jy0EHT0bcHTqm+Xof
XI2sD4e+qb7+UQndjHUQOMAiSDh9GNkLn3a6OmrQm0Lzpl4nrVES7OgvsydD+5VH
dTfQtJAKmDfTquuem2zL+e3Z0YVA2xXcpStBVuPTFR5JZdntJfQoMNbdG1HvGZir
xAeCGEbcwiEl2CsPecUguyHugFAeatzB1LennBaIkr2AbnqlYBCxZ0VgpKlMHw7w
x4h9jnEKIBRcfNwwqyG1L6UNHgRR2Lu2MklPffUg+UR8ISyozOFDOOWOWeDXVJAh
TUOkRtuDGmf5mT1EcMEmwHFVswMIjmtFI9YioSACrlKJuoScPxoXjUCTtRIDU6ZG
MHxN388jOQjzoRNO0T9e3D/6vQtdV4d2a8GCbj0t9dPrEAoww4FsdPxfifm/MxoU
XiySIHFJC6EE8JuVT7JS4XPBnJ0qMM2KTxCJOl77sU4sASNOQjC1+cLQF3AlMvvR
Q7lO3kmHygnjWCUyDB8UbRJAchKs4z28LyxxmF91P7CInD/iqDx18MpUhYr+E+iY
tgs1iEShWRUdauIBNfJTz2ab1vQc6skPEqUktCcqFJXwzUwalc97m4A7/nyP2Bud
NOZZG2nxBJBhj00DQWJdDHflszi9Er8C2luFdIAwABTje1rJ5+W+otPzK4EwAbu2
J0v8Hppk3FGVTynufIwqr/putWz0ivlQIKf8GjhWI9e7RNZZ7XRAbe4P3epKlOp2
jCB7+nrToG8DQ++EAZ/cJkX1qwWF8DFMeN0mLsgWnA65lk3mTWirg6AOXmucVYZ6
BAu7VqgyCWFGsxvQtySdJ4QIUQAS0OYoV+thPFE/39y9hUZwwgF9bjUwU5LgSssr
Jlj0Ks2GodKOqxIRimKTu00h9Y5cfG8hxVy3UZBJnN+13qjHEeC+wcfe8HDpf3nf
BXc3uBZWdicia7JOEQbMU9Gy++7KYrt0Bz08AX2ACI31+jJ5y24yphXZYaLj8TTk
ypR6w6VlDw6lY6Yg7c7ypxFikuczRTaCfmlpJpsm7gkijGnVPkHSw8RPdFne17+B
zIbHdIX1g9xRmzXKlKyph2T2sFGbifYNjNYVOpLtWU3Apbs6M1Pf3KHnDxTPgXeG
A0gNK9E8xc90G1W4KAZYffiWpPI2o7MfjjbgPtJgqs7s6s4PuTLOQ0PBPcoEfodm
HpGP+u57KellSJr7K0FhvtaqfEAtzaBYv+ZnitY3CwaPedM3cobV28SCVEyALDol
ruQywaoWaDtGz8qrhNNZP/LNaTrXlywXZl9dgcVu/5okp5TfiKotBLK5TLhGVMAV
MaxsApb4W5GglFunkL+1aaTDqCD2dLTMZj7FBtM1zA/YPMWL/BPMEbb4DBSPNdJ1
L8UdQDjHb6zzJZKgItciip+SLzDv3pMZ6BM2Jbi0pIaTQ4dE+Za4fccAHrMnCtVK
fNOVAgCCQ7imJAAaAOPk7c0PMX5NX43UeuzwehoS0JhQP2j/no2/enP6BFEiZJHv
nnbUDdaO1FrsFQ4w4KFfgZx0aiHzWePP/FuvviLgO3L7NdESG30PlgbiT0+LzDXR
vfHn3Xui5YI13Ntq9svI/qZ2KmT6PjyzQbY8ndb8YTcDz/bb097nxe8bi87busGF
miKYw0fqucfGpcwDrL0y3NohWq+WC1cHTpqg1TCFBkw5EbDImhsl9zFjzc5WlGoh
JH/4adQbMv29nNjl2Ebnltc9ya83OY871hygURvWlTQ/mUEH8SynQSy6X4glvtdq
tFUIC9rxPliT5Dd6yCnUbZS91eo2SgoBP+FTgV20Fqcfl6AOJ7j8GqcgbEi7txOv
X5YJ/q7T5ufJGZwpHj58tb47ewnvfSdv5D+f96NU0UC6sUeYNGEQad5zW5ymOImM
w8gB2ViUhdMLRr8g7em6uUcWwbropgIynCD8RV0PNWwl1PrP0JxcgC1BwrdbJPCK
KPbYntaKxaxkJ7Wfa4sgtqVG88IOz7EAgEaqDg/4wp5zFD5GpW4UGzb/4U8hvu0z
pR+0tLNh7BgTkP3MAe2U2WHzcvroHngoVwHnMyCVbpeRIEJYoJNYUxCctFt49bcn
l0acqMZLYLSVPb27+J8Ix8vJWRgLkfePSaJTwiHGfGpIjmjnPDxTG3NPb9OTYG2f
t7Nj1Z9kkKQR15W6GCZH+aR/bLZCZYcG6nYq+oVRa1MZVW3Q0imxnhqhF2vNy5xa
EqdUxBLhpREOuOXpVLcfVoeZ5pCe8L+HQ1KFqjskMfT7Le9RL23e9BS2zNqfsGw7
Uhi+wKbvmr6OOOrFZVbesFmCf+umR/Mj24OsXbwN2q7xz8SjY1Whuwq9ONNEmdb+
VksLc5cEyXSAFUb83jH3Kreez2MuV0jfIEj6n73QBN9pNTCu8FTyaBFFez0i7Hxb
w4zUkpirEOTmpG5gM/50Dyiu9FelchfXfuRBqSTx7txgoBytkC/xaAHjDEUOfh64
ukX4kF9sLQBuFdlJ4ktu8rk+QIDZNqYG25uEdqis+FaTcAP6w6WLFMf1N/bZrPtz
D3J4zERFm0kU15odOjtru5JsvgPCHQiASCG5qfFfslrq/7wotqYOtfbFML1HBoYD
znvY5x7NR6w7WNx803P3f1hw72N++yWG5qgI3G1vyYdN9mp0zIJ5WC66/2DqXCNH
l066LhtuRgkFVfgR4azsG0KFoY54u6s06GJQz9EDrikdcBXCVUzncArjLZyDt0Sl
H+5gdwma4LlSH3fYIzXnuPDwDizlwIbCTs7YhzpMXATiISWkVXHGrUkYelzlmJIC
1im2zcLwbzCzwH/Vcg90ejwsSSbWyVAdFkfjXmG05p3QkLMNe3OrfKFzpfdce4JI
eCXKs3YeJ3vVR891ogYA0gfWt70CJOY1tIHgwBuT4muhZ2u1LDQVp+jQ3LDkmCCx
diEpG5/UT/nvXIeohwypcZ6YZKDD5xem5HDkCfkfXLK5CgfiJLPUN4Z7OqEINO6p
amT8Af+SYFFVSXx6p/sK7M+ovvR+BvlDjkmCSIqRq3CQnJGOEovQkAKqXVqaApwN
bsL9oJzsO99OO11KI6iZ7loY/WS98c5jlguJKzKdlm5dspcWjx37gbZshjW5ICHt
OpKcnp1FD5rPpTHznz9ig4zU2BpI7nPwLp55q6WYGUBSeSyyG9SC1f631kJeUT7A
a9PZo6A35BqnHHRwLi9e/HByN/asyg+c2d8crJODAvIqiHO5gCuCY27rHZ7rlE7w
IYHw+hLR5G5rCogGeoKQI3OtIF0SlcvmH4f0CxXC8AWWvza3t6iCuXSguuOAxQPZ
ciCzEi88aMUGdS1oKHOOBTV87qoQiTEgDK4GPCeDK/jr+CEXYElESCAJoTtUqp9W
Mk4yAHB0RwJ2ETXLOWX1ZD925RX8v1785jin0Xsl4KE2nBww5ojQZc6jG1NAVtoL
yCeQpT7o9scrtOyw3/yJObh3nYxFXJ0jxYwGWddN2ljI2Hh2RI9T6aShqGqhvLtv
oLv5SmKVKV48ZQ755CgT6XA1wUVRpP6TB7/MaLijKyEitIA4QtwkefmbqGFnbZR6
ZQexj0hVZeQrz34sQSMw+XU5esIiDqOwl6FoicxVkWGEjlzM9QGPwk9QPc6RS7KU
6zBipGziB6kaedb7xC+9VHWmRe68LP0xlrcazldOBUBFqGJy3O3O+1DFqukESmnB
Q446+xE5Q+881CHS9XZTGc8zX1PMApcvniRaFTZ7sSFSZUgOBF+hqDBKxH8epV55
o2ZPWoxhSw+qFtKj+/n6O1TYW0dEFvxjx4AgNuC34SjoSs6XYsnmkz2Ri5YTFkkP
xZmpiqPbi1O4rJnO8lWOAyZgXa4q0FVs4Qg97YPp37CGAT2Ymdg5k6JMkDgVYMcR
2q2CanQeXNEpBPtSrjo6a5RUBMe/+kOUOrDi7w2tqgcYqZGv8GuznkXuZP7Xnsfy
NBNP5HXjo7jxuWl+xlBOpCchXqXcaMr9Ys4qSFdU5nr8T7gI5W9HcNmDOIxGwUNW
Gki7IpKmC7MjZAD/yQWwz1jrPk/xsmypmWgw+0a3HgIOkg5nrROqkKHJYg9NCOib
yjQzI6QQg7/Otcaxef8RGX/14KAYbGgXWX9lvruoDBqUTIpnv+84khLgGvmeujbd
hVC2CkHmUyvIt2s4OtQnj4qgAK8jjVGiDYXOOOIG2AL1nV2dGcSHJ/DvnZVmoWkZ
F7uGy3gCpzJTGR4l9QfcOJETn8tCKIOb9zH1wSvSwW9OuWsSHZ9Le3DwDJVrjp5r
kmV5bWjowT13rh1Ywlo0WttD+LSCfXN6vgkbR6StFxFx96wJjkvINdSNln/1Njox
MIcKURKXr73HujZxjl7MMICO+mc3MThB4JOFeaF7hBowieOIDFvcHuMlVSq33uZ3
59LTqqW5qMlXHxX1qpKrd95kgeJSoEZMVAdktfB3iKPwJE6IBNRoaKcxsmCs8egi
XLT7LHXvMyG5tqzEq5dfUh8Tmaj2TyG6mbMFXg88SzWKSbK54RhXqnsVayIBbWDS
/OIzXGonCmLXxk+S7/4ty2AkGrdJxhgHG1d/uPRZZQncUfTpa9rRyO4eygxTOo2a
0JnSVwWPKcFYodb0fHVHzfULUx/u4bGoWIvFL6ejW9hBtWyq8qpUV7eDx1hoJ+sR
mqF1A6lg3fJthJ3qwu8xXi59OvUP7GnU3y6A2iL8hyK21XwM2naucOydXeNZShYg
3YbLYPvgw5rzP9b+ZRPS6f/bRh8TSIFiiGIxPIYbZv9pQy1U8hR56TN4HdKOHNqT
/SVgu9q7HiuNGndT17TVW+saRUT6uKAXfYpW9UgksawpTD9gppmMHWVJ/9Bv+VtH
DywzgVd2w0wxQX3zvu4aIF+b5WYIAFSEaVkFiUf910fKUZ7zw+WO4WgHNzfXDdGp
Fl0okwwaiOmpzSP4i2Jiuijjq4+OQ5ipQ7Wzn+FuL+bcO34Ird++a2PfnA/SdRT9
zaGoNyZ++aoYAYfuoModWuFU5MrSlTxixa7pb//pcxSWsy9zqrOzHixg8xjkgra7
kx0JbFsqNF/hB9yXUwmHlAnVQBDBl0+44LXtkOmv1VYaMx6NBucIH8px8CANT7SX
6CGx4z9GD8Cl3jf63MlO18DXR4jQ6dpCXKAvf0f3SXDjTdyRbaOQvgxxiw76mqXx
cUKzXSBPRlIb+S/+2K1CYnPDzPg2X+g0pZJdasRoaf8AlUD3/JlXhaDcrdcNLu9O
RDNyDrD2el09WW3fPUVMWtThcVmDYrH2FaujxQ0N0lbJNQp9hYp/k+X+jgUEA5Kx
i0YYrcDGBcGwdQqP2ZDtU2mwSGFrMCO4VGfEhmX26EkKBwT+XYNAZkf0z3S/GuaD
U0fr4Zp17KHrR5xtFGjbMF7+4Gdzci6eSOxjtupOkD6Kz44bpVf88UbkxtypBWgd
QkiWN2v4Kqrw+79/IYEsdQrbMO1ZBIo31ObDlY0PZbG4mTuChoT2Tv7DxpF3WpNl
BhGXSJl7M+ehdgmTIRlHjxHIOfTZAEupzVJfIQtZdleoX6v2NdlLPfO2D+jwivVN
IXrFGy6ftVp01PXCWzjX2XA5U7JeKdw2ykwZRAhdr4SDZTCYOOClP9DcdiF5gWx3
GR1qhkFw3uKV2HSPY/P6bk5Oox/GofitP/AFQtVWccRKHnuhhrvyNHbFGcgS3ARM
FVjOCR+llv+5sgm/CwW4P64L/Mz0Uml9E3lCIb3Nb+NueawpL3Wx/MD3YjUV5lur
ZSdI3EQbgEOJltS80DsT5108OQOrEEnm32nnc1JIU7sOlagso5Kfz1ALXIAJXCic
sjChruwzhwtPPerVc+PiI8UNPDqkzseMVmqqVFMFxKSz0qa7ooobDX47B44c6zIN
jUcxsXGGtGuacOlnLOa56bRp4jJ+SrxCcsLYFl3QT0+yrwjgfXmZjsiT5NJX+k1M
Q3+i66MV0cAHyyx1Ml3meIi1rddoMm0bGVJLFJMgcoULM1cqtih3qEOFJ5XhkSMJ
1EOwHUxi7QWtpI8uM4UZsI1g8ZSf99+ghBURO+3Gon0rtbjA/CBAbJi9DA7Koft2
T7HiB7tnjbo5vG0GJ6KoPzaTcO1xncomxxLn+h45aU0qLvsR5koEnV45fRsO4uVd
Z7sr+c0o9rBVectXn+aVq1Afh4Tqk+5Q5+QFIflbZWufHh+N9iOiqgI/KgCsu2KU
LxZ8USdvKCQVcnNkpRyo78XiwG/tKT6ZB7vggjtLYSPw7JiCdgMCull6BJZXbfXK
YZMAjhG2+NqEP1z/2mfOBAEv6AxVzihgKcZrTTbq1P4EiNzaPdymv2sD+l+Ml5Y/
yFIsVi1QCGSuygpJ6t1GOhEzgGGmnofJTyk+UaQgOMfNUTNd/7LrczYiVLEj3Ln7
KuUh1HOftgC7NeNdMkyCaJqJWohcTtF3dcgduc+MXtRJRgmcsoV8PvyLqtmaEnkI
L7beOe0YgSepdMIRKkCksd3HQW7FpnSKw8J/9zydRaffO7hzndiTHZDhCfzYPFfA
DnwmKSOo5I7RmHgVb0BsY55K4+Nb2Nx1Kl+c9d61O9LkfUEDq+jwuiYG7hSXFfL6
OoqsrfjjKq6mcaUDAEXofqSDmmcBvHPGDEks3frB9kj6rB4KtGDP938AjgmZITVp
EPkitO3kHfQh8xyh3XTU957O/OvTNmBRSD7XaW01QXpWO7erVLGj9LkbkPSmpXhA
4bxN4OIFmF3Hf2OFo5q8ELKKT/EYkqwzVuGP7ZmVioBl5jr5MEPxPTsDlMwI5syP
N89MZBhjYdkC3K3UfkS0V39geYAaMXwqcG0+UqbtnifiJ5nXeRD6QlFSR9Cfe9pG
fBYV+msHyJ279zRCnuuzCcBPZPojbKb6ktKSRkcOwxABM8qwN4aGedal+4Musbzv
vohy2SRzrZGLFZzVqWOwTgk6kjosd5DKNwZLTydpHJ0ve/Pu9didoBObzr0NDR+9
oCZKOb6SnqWvSTE2wWyOcboWMz3rIO92gSSbs0z+u1EKSH4Ye24hnJUfUlXqruNd
CWx5uKMDxmzv6HIfMTjKpaefMHdbDUC6mqoCTN4cRKrTRf6jnyiAWszS6Bho5xl5
dptb7Rg8wW7Q7pHy6XhEi9L7rf00nIe7iOjgmcNaonmxX4nZHVTFWnjP3xb7WoXq
x2CEP95Lmndo1vRQczaj6+xLak0I/2dgvzeDL0UYmvmqyAd9SMzt5Eued6V19nm4
tLgfgXwI4rxbpWiEzuyJoKQ602d5R6AInkuPXu2r56PI2oVszVeXCNen4P2WKKaV
T/SpSs9xTuBdRaWgL8V1QkS+xNhkQvsEUcT8F0L+GGjitXj6XBE3EQX/ZTggUvH6
m7AcuTAjkgTPovFxnKKy7/7fBSTJvOpjRiMBLs5OaRbVpOggriGcD4LZr+Z1T3EQ
n5eIGjWjTRI3MNtY9BnY4K95XrmhRXstttcuBgC57t63ZGKeNpZ62xW/7izW0Jou
65zwmOaz54f+ibewjDWk6kIFyV9KZl/8w3h9lb4lHl85aG0boy5OHGh3QSTStBg2
veuU7mkiI9f5cSW/tFKrBRVpgeG5C5p8Uxbh4pEkyz8PIXNUzjL2VoC1mWyMhsNx
Sd9I4JUpCbzFUxP8rWm+O4CjU9yNP4QWdBA2HIczm2V5ajCgZBtV3nzlmKfEfs2W
AOOiE3TfnPP9EDt2SsWq1Gn6qYS+sydWq9WVLFPwgewXMRIObxaVy/itLqIzfOuh
mjbT1JOaj8uWxsx83QC9J6EAnuy+JmbuO9xKYz3hsAz65hf//UpzuB/Uo2iYg/7Z
lSfl4ndTRb4ZGjIlDUxK+OUMYSc6f3Cpm8iTV0n/EJf76pbm0dSolX+5cFjXvqzu
RbO4kwh6v64yyPY1XJRplEQl3vEDAVIalfrHXloa4J4lrsufGFwFA+FzVhFIUbXJ
9t7MUKBAELhM5q59A+8g+5T5kZwokRWnzc0ntYVxVuI1/z+JX2Tj3zyZNoTNJhZV
YnKLlKbXN1K3kqIPv2Bvh9JiwubPsz9aw8MrVj9qKKjWE1K620S29Z0qWKEYSVKA
+B8SqGP15c1AijvMPilUJlL/zteJ5b8A8YGkQWA8XGxltTh4Wjh8WOLZ8ant+fTU
YJRcLiN2KnGP0Rx5QL1srHRq4lm5PWGzUkKh8Is06R2BhwuDYTPuOmzIWbh3RFUO
rDYGjWVMOt6DbvyhocPTsdH3WxOtZL3Bhf4HFgv/BFI7ibTQOCfNVYhr/6n/Sizp
JzaFiSKYmeyLM0XqdG4BGeX0janJFL+CopfMeKVK12FeDJUMFL0Rf9sH5c5HS+fu
qH4EVPK6iPpK0GaKjrfTVrxFKoeLJtSZWadG84K1372TV1i8R7/tq5H2MJw0R22D
jBMW8SQ9I/Nv3dj3GCckPNfLvnsgiHmw/eTD+/OdxC7OdeIoWwczHSPjm/ijNVRf
2b10jhNcCfIgDupFoJBbfrTzqZoU0030F6WznYyGzCh8wyaIVzJyxc6zjoZG0Vbs
+YZUu7lP7lKGopLX/h19Z9nTlVq43RaMBuNiQlWAVw1Jag1qRIw2rg5X1h+XpMdP
JNVYlc3afWm9IZBF5xmkUne412m94PT2sYY4oGyXC/5pQgXewpsp3bVeNq+smAzg
vQfryRwjWII/53t098MdsTFTVbqQ20PtQASIAiKmGrJeCnQXPVyze9QOfIrh/KU/
DxG3IsVxJMowlC/PC05bVnqBGjZYypPlPjL6CTbh88AKtRFXXZ5GPu9jo8QgtEGQ
NRGLuRgxR1uQ3V2IXxOfOOmhNzi1v8oBA6eIq5J2HebSmeF42uVWmyeWibT9IYu4
o3Tt2tVuaRMLbh6S2CeKAjduROSUIZMxlgt6KfyEVRl9XKSVnum0bSR58+7R4PJX
pcHgAeG+W2pCMPaESjaHtlW+qjMy5IkGVU3tVPU9AvWJbJUNdtxXqg+K/9Hz+M/C
t1UOKkJHNfOSRXvezF3c0hSRZBOLHdNaVc+adtmLhTZVSn88FiVyhWaWGnDEtuWb
wZpVaRfAwRfqQ1IlaN86RMjAPpsI3X9ez9uMvRlBh7l4FQzhNugKz0YZHWWxbih2
f1vV5zMBf+1OC7HVC0kjXnQbX6diuAeWOQVH3HXsYVFC8Q87l+2xy3RWH9Fvmov1
MrsY3FbyY6Oj5hkbNDE834oLHdjFqO0IlE3ZvOzXvRDwpVw6/9J4L8mwPzOD2vP8
VXYm1LZxaueZV7hjGJqf2PR3MY72TXpIKjUJugswRzJp66RVHiqLDjGE4dM/FPSf
HG7/OqkgIHaNqq+Pi0XFVbP1yea8UPa4+0JPSiNsue5Nq7u7k1pvtRiVOZgqS0Lw
LLBTVDIz2x31owrWEk3VMAS/DnzFBT8JttxKAj+QM7raEti8/meV/du4iwcNQhq+
D7Tbs6R9ey4UmXK00rcpehh0WkIHBtdE0n3PVNGQrdAgGWCzfmda87wMSha/6Gqz
H/X47OV+eb5I2OfVbF56JwbrdEFChdK/57iYYh3boMQ68Ma28IchrlOAcWk3nUrc
dfszyNf5uNBhJx6m5V49EPpXEtfW+ujPY54r6emBMUQKn+6P8CN/WGeHfe9lokGD
nZkrTYYu9nN788fK3HCcB1CyNirUHNm85SFHyU97OL4Qq1UVXPp8dHKoJt/CE7wf
fQgZkoU/Y4rT31FlhCuu+0i1/hHT+Ur79T6AJHrzUbMn7GXhPXn/QGh0FHtjizTQ
SSTpzIn3CZKol5BRfkJGr81qtLE4Ue4zNMuPX/NvLrQ3YZxU95fRNdUFYLLRZv6d
50+2Jq4W6f1MiLxqqRrERFPHgZICWGNlwzm0VmE+DDSaD74pUR5tasq7Sd2AU9cV
IhUgjAar6eU9f9/8+ucLYtuI5BJG8fjVNgU5CMd8h+WU+4QpfztJKZwXGUKaap2+
GYaqjD+Ud3U365DV73GoM0OLGtMBCBvDQfJy68YX0tfBkcHn2GEqOR7/ZjA1JQrd
ojsa4V6D5vfpGEQxavYz5dq0tfOJrLiurZZefZMYvWpN+HuUgYoW2+E03GzIvKz3
IAUPXuOIQb2CDqoooZirAIKNSRFbnFKKXdP5PKaZ30c2QZkYGXcEF0N1yY6kTvZg
xjzCvxoKSQeJ6p3NesD8Y1ONk/rdW25TpO2Xik8c8SadC9oHg40o0gOIog3JRTvh
DHRfHguvBOeTAtHGXf/9Ed9fZr2Qb1JvxQICmNCWNpFTrO/iVwfLFmbZySxYmkDQ
Y6V9L+H2Z8Sq8+SkwBXk26FjINNwOt3X0qNFdPfYtnq8s66APaWCXKnj+MIS8t0k
6xJacJrAeOZGohbevwoDwfIVB1THnFR4mJxmQHEERYFjgonbSXZjVMqTHb7IOQ2h
z1mE2MD/kK0SnWR47LIHJrcCYsO6hy5EpVRESGlx89DOEfkH1U91hBaWKjuS1n1G
tdOmA7fktfmvhyRi/6eWMmYcfpXoYdGZm5QmxfDn9Gh8BS8+vQGn6SVEX7CoJuj3
OamEAbQluwMIR55lUkGbaTA5oqTZXR5mIuFn0He84d3ZZUIOlqaOyppsfg/bhTE1
bz62ZzRUvrS/d2IaSi2T6UEYR73M754/kEJGZZ6VCK+UW9yXE0ORjlAFttEQh5vU
wHH/e5T6OoEgULGXavEEBXGhMfM+JHsufUJpR6DFnk+Js6g4hZ6ac0yc8JRh4R9F
bYWzEjvlt8ObwaC9sIHlAw6G/DzCk7+cRXosDiDt3miPRiAJDfmWmeYpRc56N8GV
atz0ja2FKI3dWrabTaRHGdIUfJxL3yL2sLdPbMR13L+CaJ0MIUUn8QvGBy1MIKEc
9XYKONhA2X2Uq5WEWSjL2R/DjAR8jiVm+wxgXebX11uSavs+yb7Jplgt2Gfuz+Qc
L6odWSKBfXUjnKlriD15OQERtX07Gs77nU3LgZGI0vJEOIbvLZK8a1DLkv79lylv
L3Y47FPwaXnjnB9FRtY/ZLRUc3NorA5sci1+aRtim0DfrAPJdTUOoUkUY/V+L8wr
Y8oHmaLeKXkXsVwEGKjf0iZDoqjRHWjE+Rg/Tf/nKAcPjFxRGzCZ/6fFFDem/bLd
r4IMIngC3tw95tqRGIyQDOY71A0QX8q+pdKDAeolXmNIimM6O68exH625xBO/u+s
+ofwxRt+znocgiorYr5t7XA7zuw3HBw/tD2+Yb4QNgigUDffB+HYYAdhmDUeVvQ8
ZS9qsvMbkhpUgw4IXNzODFgHI0XfquQWw8E2dwqP43G3Ojzy9X9Cn2buHPWm7gz/
Zf1MUMlkWKhCD3JOSLTWTwT6OOck3BkBl70+9x1HKhIpDlPFG02F+Rwr9bCEofJG
bNYdQiQ+oq0GrwVKhxjHsBe2hsRZcUYXPARMmT/3ZWbnArg/vvjBlgJss30cl1+5
JG8pqBXCYBGlKdk/CDZy3eH5/eZXY+fQT6PM/aIxrIEhkN47VurWZgd7/r3l+L6j
4afV6Ko/HmUERXLqDOOVDMfgIhoYzM3Pxk3wS3Fbvx74h+Ah0muQ8yH2TgE0Ri3n
e2zvTueaveG57jqBPP2WY80k74XvvkjiADk0GhM7FmLJufNrEkViYqN01QPTOXpY
dt9e97LnZHl73GPaZLRI4MSLSStMGC9YhWAEDxYi2Ypt4iLAeeM5zWGHvoHRl2Wj
nszb4H1WMboVR0LejQLaASSt5/hlNVw9470tHI6yIcl+m/69u3hlyUtrAKl960Yr
v+ZD5n2o6vUuikbJRHUTBUDodfmZKb55/d/SmUUcwfyZjE2b8E4L1bLdAXR5gjvN
lth2buluk/3abVLl8yANyF30mxjLtatlwJTBu0sQYPzd9wblCF/45bbUMkab1Ogp
hxS9A3hTQmu3Tp0HYBpWs7sho1nhC96ga46MQYMFSt8VRk1eopJaOy2d9mNwhObw
mhbmRh7qmnwgowCyfpzka4HneodXY6wsw7Rwr7BmOBANfhcUbBqZj3z3mSXauO6h
ZdedjLQVhn1L4zO7uisHLs4J9sCp+yY/ZJ/5GEAXgloDJhTw5A1C0hP5cnibDU8l
i6V8pndZBT+XjwZ6NzXzQAwI+KMVdH2Rw6Gy4eEwCoPbh4SWrEvb+vw9RnLoyKH2
K7zA+HZjTFl7uby/OTSQ5Om8W/NtyZtOt+uG44QTl6/bpZiDUqMJLhsyweI4bEa0
bZLWW+Y9KsxX5K/32IrU01r5ScCgGc1hy18DuH4s9qvL3YhDCb5j1ACL0jd0dewk
Da1Rhxc4ch+sxN3tcxXbNlvMnG/qlGIzdwR7AZPFd6Z65MakHwLkEEGINdsLr7hX
93xhyQa3Y5vFyvfEU91bKaRdWB/b9rjR2rP0EA9945txOvboX41xW+SZSGmCyISb
2Imvkupm5WNwEB79s58Fo0nslkZfZQs+2dWfOB9pR6YGozHqi68oLru0imdt9pxX
BkmPNKocqywkhZdXjjlQLzdnJ0dycdcDrAQakhyeI78hlYYIZofyA1//Mp0YhHMS
3J79kH49Erw4e5Gj30arqhrRdCfISrvm1eTjER/SXIpjeUpSTRYXQBUzsjF2eWnG
kzkfstlG5BrJyVjyfXL/z/V0Lw+Lp2dj2XiPePO6YQPsBRiqX8OnjeMh4tQJYmMS
ZFeFol8HtUPTCTFFb/rCbJ64sXZbs1RXp5xVsopxZc8j+wxH+hP0zIlteOBdBY+r
gcMev0BDp5/c8YGYPHxnDZ8EARRXFxVFrYGplAFrbMn7eN/5c0hut6xZDzZAU01W
6/QDhjEuM42nUnAsC6ruwBdvAfnINcag3edeQ8JiXzJ+VcCPjeKQUgnC7bTOlp3L
GrMwSdeALwYN71aWBVkCsk8YAzzid21fPaYQSxfiDRfO8au6Jv8D8RacKc/oNPFb
tWYBLN4x04RSIiZrMyUI2k5OozfBR/jLCosXMlY/zrwbwsb1Epg1ArjcqI5H35aV
7B4gexATihhAlyZrzYgY6Y8Erd5Z1NhpgCKXuYCkMVedvHBatieCj+ig+JDq5Ayy
gl8tyKftOaSvWW5Dma6H9trIQ5brYbTvYfdh67TsOvvWKyQEaI6Q/Gfx6r9AhIVs
jlFuO6ctYabQglTwQYfAKrNHjEIlfLEIFfkD3GdUouOu5HM2L6SvnC5pMvTkh3Yh
302+yXXoKXmY5EnWd4vWC4kJrykLin93DwD1NjTPuwV3Zvj4RgC9D/1gpcbiOvFa
D3mIfj39QomiwZU/XG1Wu5nYp82LtXf4PgoLEj4buJKpiTOWK6fF49ml3ZSHlr+O
piuDBdP0wC1+EIYwIZRqNqwztyi5/anSoZHo5XK3T617KudLJM357jPsBuHLgHEr
WqYRDZ1atEy42TZbIZ0yTzTwJ9zZX2AeCWDOaTArfSc8RYaRhaCoajDbBh/XOS75
0cPETB2TN6qt7joZlg0F+ayq4ufOR5gflAzmOqulREyuX4/s9mZhO8I+q9tMd89S
4K0Eai/7HJpVHpcnJTWqeQfUVup0BQ2Jc9B41s+ynPPkZlG7fCa+RGF3rBMKXp/m
0LCBMrGOXBhM+n8szYHV+ct9maoYmGNptvrGfqts4tTl5zhCiN19wVHfh5NAJYYM
B/7+dxTRRIXKpYIW+hDAA3XcOVAO7aCSB/tenoD38CqUxT4XoaaIIy+U2CezUv9E
rCBL54I5yNd2xba+4XMX5fghJOx88+KLSLrYHcb6YNbRXkvE8cb2BBhib29PBdDQ
JFdiJ8fPQDTUiw6wtGhceaNUWOt0N/YfTyRot6U1TiHlAAlX1O3u5PmEo9hmVnMK
/S7+WMucLH366Gz9WT83IB4ch6oQGGxLw8oqv8d4nIIfs3aettgWyMAa5kAhBQTV
H7fXkmSdUZsYsP/EfoLZZLylKG2s3Hhnj6l1XmC4idGLQctsonQGIj/BkbN9D7CU
KmSOwsmYhz41QfYkh5bfRDqdmnZ68AxQaNOMpl0x7P3gVjsPHR08IF444Q0UKHNB
P6sLU39oijBmtNneDyHlPjWiHw4mw9jdj59ruinOScD1zDf12ZxI4/awJ+VtonDn
QhoydqixMLGHyawh9/JAxwuwMV3jdqhky49cg9u4wp5SuPru0FKNbj7OcUlOy2+y
TL/SDaOBmcwEOsqpM8zh8brTpvW/QrQjEt68BITtoPuGQkaU+fEp4WW/2vl706t/
1IK9iEKMJeOj1jCcPru7FvKIb6c8yczIggqBvymoSA1fuAaXKFw3cZEW9Ncazc5H
NHRD69kdx5rjl95p9kIqfzVMSTSIXJj/s5xnpu+3VpzWN9kEZOu+JqJcgc947wmi
+jzdYaGuWXe4vnjC68cnslNIE04KPI64w4hSkJrEitWW1Dlz2DYgG2Xh7MOS48x/
05INckrvvb1jB96d5fx3Tuj9gGgI2x2Ky4VipNYHgGS2cOOCFZd9Oz7qcOEGXTt+
r8m4Qw/iGSbT67aCi1WbafFWPfJ2v3CUTxfv/GbKd1uS1AfvHJTRIuO2wVrBdBuk
YSeOegC4mZQqbvr1jNz9uFnfL+WM6TgDCf0LzSOPk197JIjw8Waa8DHY4zxRbdBS
GJMgW3T4TuRyFb4oc6woinNTHhGkwT7krgenhxnO2EVS/NJJ5lC7ShnPuc25cENe
2I/2LtCSR1NQWN3k0HlfFcQRFTQNYmSAA/ooiHvFQxUWQEVuLv6qLL63Kn0BKKsk
wru/S9kPw9HyFyTPg85LKTlgTWs22ZhSxBIYPqDum2kVUcfiPjDo+vzyOGexmBSi
qeVvHMWQbfaADLjWhWWGmdiHO3tacXorZ9KCQ/9KGkVipsRyN4wtIczTRGQ1zPmo
kbtJhYZrwZdpdB50dB3aIlfqEBpTrK8rKXVC759LTFIfuqgWlvXU1Atm3Jfwi+jp
e6foYrqYNo64yuIQaWVvirPcNHrjZOocolJ0ACysd8ApMCSpDJu0Rf3BxcmJXeM+
Y/tHtHnTsCBVaSn/Svs3/ADs9V5Ms6JLRlLdwre1Wq7iCnDNiODvY/HZ5u5YQmwH
V5uIr9q77+kDfqoPCKgnjKsNGlK6pH1vRKJ/j6Es22mW4IWUF9qGPqeYCqov7YDW
cXtH9i98bb4WtNOKQblh2u5zTYB1xzTkxK6+ZlHz2FRT4zfDs+l1NV5shd415UlP
k88uqZS7gfP1PmCgimNJ0swfoW/y17xvBYw4oDjh+82oJ9dbgkT3SFcFUpMwPPeN
bgMB2noU7pQDLDN4lucW37bqPiVoxnQds+EyFDM1CzfUCaR7qTWaSF5HAmnusG8Y
VvtqAwXKqASmG95zUbZkHztLt80Snw0cFnLOveoF5d94PCz9ctszoLa10wodLnUA
PmSz4cbANcKn60U7FDi4FJxl4+s2PnWVDOYIFkb3B+sGdjA4GvobG51eFt4Jkuqh
D+341MSmqR8uUBRD8N0yWtn4Zpch9D5TdKWN+ymCgyqtRAYcBXdsGutlWaHT4tvP
QL2iukoalbDzrG/ZTBMS/4cC5GwONq7N4F2e+PqZoZcMuNICDv3YL7m5rbI/90TH
De4fj0Hiw2pFs868mgLZ1G2+wL0X2tX0D0pO6HKT1fBXntAo/YvkLtdAdltefHzm
UKaxkaCRzpL7kKV6gMeDSnvX0IjP1f+gN/IS8SAYlP6wxguMK+xvFmj5h1Eo1t4r
6dx5sH6G+Py/dejBeEiZqvylycn98ac0+4qeNkA20JkVwCKkrKpqUt4ofkvYFORe
8SVLWy8Z17bkapR4JLY3wVl3vsXx7UiRtJZMc81kZnJPElqgU8Ahkn8xHiI+coPq
bBWAWhZlQNFyYrmvhiSqMJDB5n2TTcZ5by7RmRBq6gTOQf6N8Xv1K2JuTLFCm72r
ozE0Oh+4EK+THTlI9Sxb2F/pVHu6r7BPcNm/sxoWzuvstHC1jgkAc8Gy2jT/Qgyh
T1SkueYemG8RvU41HFRj0G4m2yqBTiP9z+V+zl0ZqJFso87anjhlp/DAv2OdchIW
vwH1gu7tQlwTcstdoyxv6CtDBsenRLQil1l+97uTFZ9hCGhTLPnGXX/LX9odgnRC
OlTiS8++EpwteUq48TD9BpklKJrgc+jL8H0N6wSuRLm3gnps/90sWbIugQC44Iku
IyarM69Q3bApAcJx6Pquad76XlWL3WeiKitCCrPtaYNi9kiGPXXVntJUCEND1fj3
QFmAPyCa7gNd2EDcR6BPEG5K1VCXSf+65f48lYXsPCCkxYs9IsJhUJcQZGK1yav3
dS7hkVajrMN+wEAeEl6z4AAv2E0bN9oMBFuhVt811PxPOBdQIIhd4Y9SO5TFVtF5
l5GcYhH6KKC2UNY88UVKBhoAjeVK1ziIGebVSRVZ0aQmD7q480SJxqTP+1CZgjE4
TrBg7PQGBJjMWWD2h5lSJxwvgq/Hcf+qVK9ZHy3bKJ/EqcRvx9YKlbngZBhu8nV0
DwsgkD9B35tXULOdLRfxNxsNomNuzDi4AuOHpb2AMerQNNxmhW4b3vpuFsTxOV9a
wzphiyRRkN6EkR1BQr38r+PHLYZ/uJKrePMBmDNQ4IBz4BA8C1yvibuXjFBhziiO
t+MiZETc+xDBAYu7yaCwXRRraz0s3xoq3xa4gq+EDSJ+8fCtsgtsvvMx1MMRWmm1
Iom885TxSDG2tlS+A1OUovmEzsMXgYtEzvITJ7OKeGhFKT4k76J1a/EDgVMj1xTC
wJKY2U9xS22bXEavEEGpzT2pm6Gvp3HDi4SWQPpg36fENY/6fq7PZn3f9g7HES2U
d0uzAoNM2EO36JQ+hH7FXuWB3vBiY3r4aAtF8r3L9+HMxSdfPnvcrvjGresJV4ib
slsxYJFCDf/8b6hFX71nGGW8p3cZemR+fpm2EJ2nZsfYAgnyWC9LwosI4gMEX2kh
K64OWh0pGMGEHMIDDlIcHj2xgZQIi5a+vWg6Q+VxEnBy8tZYbaV/6ofHd+gAvIFT
MuImpRevt+Jqv7AIhUtTDzV8JWqfwzUsnp15FnwhM2Zqh6OUkuoqEomECyTUoQgv
CzR+lQ5Zj0uDMt1/KoCNwYSgI9dzJ5xlk1CL+XYdArQsQC9n+U5aYBGVRmOH+Zbn
HUmmRIrp4ceoJp00YYqxA8cI7dPcDzWKBGdutIXG+woUuPN1U7AlHR3kwHgUtne/
exakd422Saz3ByFBami17BC+30ssfZaCppjFqXdoBLVYQ5tClLiX/dFmDY7VjbpW
q5YwVrZjdfaW4wPbxa7VPe71z/InGl7Ed16s0OrZFYVX8MfV7exIt3ltPFFFSHQg
i47HCWeVNPfa/VAtRwJLPRwfUcSgQgjW/aEzQqlW/xpVGI8TTygDUm2T2Lu1gIf4
abHHQkE78ZCcP02rPP6HrLPMO8QdGwZSu09VFrkkM/JOkpyKyFelewVOOcEtyZVn
Ce28WsVHiWpLJZjezmV3oIs4VQyQKUy2AyVahoM6ltasVTKf7wxYiwm5u4TMrXQi
tNPTqzv/3mFp6fZBxYseqDsOjeCZfMBfd4yQkt2xgumZ/WALCDeUolXvAOXkZCDd
qa31N9FIWGdBotsZWM0Xe0zCFKWvm/+5RmvMZZuoTWHfYQeDqWwZkvlclF8cDN2s
kSxuaTaCmrutAJuJng4aG9Ltyox+bNj8dt+1Yqpl+MyQKNUwE9lne1HucO94XZP3
RPcTM/fHZMWcmzsRLMwLf63mQHL5qT7jA+rpq/1XxOuc27bdvzm9fz2Eaaw34c1O
ZxiRiekSWUZh/OO3oXBP9S3yxzH9GiKoVQfgZdU6DT3WUFOQ44TRyPUPSnJg72IW
no+Vx9/ds8+QAVQvYtNE/b4875dyrcsdwQmJdI+BIFQAT3IfJiToeP9FqNCnyehZ
iy+tC9IgrYZSyM0+OE2DZOFPGWWsAE3ckv1zAUxZr1ktWc75P+CRfpFKoHgmBXiQ
hZpmYzn3FX5GTyH/4epC6glChhLcFJmelRTzykwFDzYtXWySp8PNkCirY0Y3BBZ9
L3Dd2PPL7lge6pIYiw5g71Ez+J+Cd07LWrN6Ds+lpPJRpHmjODIk9mQJ8OIXhQCM
CHx1jU4LbuKYKZsPxNNyWlWjFfiYpGnJf3nbjAqfLwZ954dyseDDAW85JmHS4qx4
HhypkyEAYlD65FAavJOtPJFjbf2ugtncCQUBEu3UIhWN23p4GbM3CkWMjFd4JhBW
A/AOFkqqWMJzUoV/+UbuqQchmTsdAXf5+HFfBGHwDYdKAusEeWzM/B9NC9Iu/haN
ZphjZ045zHLQrY2jwkYk5sqyyA5OzjBXhITd4NAL6H7GqQ6m3IASMHBjMt2VahKs
c7hXyA03MqoBa7uvnlpqWG9lXvhzj2imOFd7tO0AlgGRFTnoCxA2/YPUw6YEhycM
tQZywn+FiT9GLqxVw4EesSZiWTPGNe890sSKtrFb/+qWEU+OiNKa+1FQ1xraBxt+
U882UGtJuqCAY4iLXaBczRlvpbiYHe7gynAq711aS3rwZ8aLdVBw/LuHK33cer0W
lVDykgs7K1x421dNQizcbYEjjszurmgfEYers0/tVYuCzBAn77+orqkmajGPO6K6
gCZwV3Zq8RGv7+Tkwv+3iSt896ElGZatPyB9yY3e+1PV4o/JwXhAqbSwfgNd38uv
eXJa7k6Ph6qiGiGUPot1Qk40ZcX5EVF+/n4ImH2yzY4n1SRTmyt7IWwTaHMTol//
4FI3nlx1QTyavV4lYLr1PFbJhs6L1O2c8Wp8H4cHkhoM22IKr3/ghQfs0YcV0J+v
owZ5D6s/yxX4qegcmmqFq+bMxKyR/+m2aOsx17GyVy5THKccwuvegVLLavkTNJXq
jJ+WeS2ut63QG3UfBQ2t4GG3NRBa+xl37ll+tU44Qg6VzHON9RQkjO8thg1VjePs
FP5dCPTPVgHtUhsW3wwgGkCmovGpvK0OYnYAFEaQjWWNxGR3a8oLgmiVIzig+emB
FDPQlpBB15WbzGkStkqFUnv8GhWV+28Uyr3unSw1Bo/GhggLvtCE6pLpmbuSf27S
82FKrQvZgtQjNMoaHudOvELPASo5Q5Ig4n7BInDhKy4IyLCo/nqGdA0P0yl4MHV7
CL3PnpQN5r7vpcxAw8uuyS/Mtbg1W0o//OOMmybhi9NvLuA11LQ/o5O9SXhEt4Pz
FdifflyHhsUn9zFxvfnC9Fy/R+uL1FB6dRfz2KnhYSIMkBMxD+79BQ1yptKnqP+X
dwtQUrJOzFu0lVsKhcz/SLDsXNe8BrNrNwSp4F+DZeOCT1GQKzb0WniQq6tFB4U3
MHs0znrncAGUSDAR+rgKSa2WVJbgz5Rhjk1tud2/zzCqlgeMK/hngokOj9hseE6P
RBx6Nn2NBvemR/SBQmZ50MrFuAVyn5F1AS1lXcQDYdJFMERj648jwoQVJb1avErf
7vBROen8XTVlYb2jGJQzNKKo+tZaDbOqOyyYdGwBAhp+WWC4EQ/B40kx4/WTGpyM
Q1UOql8WwL8a3qywNxcA6I2PaLzYJzSttn8nejn6uXzt2jBwJyxfisrg6f0eqeXD
nlXBda1tj8aB4MDwFo7+In4rAPXGM6rUK8BXLB9XnsGUGiNWYgwUDZ5sR20Pq57B
PK2B5L5tJqTSm2u0I41HtUaJeKZgM0hiyHBxHvEB+y4jg1l7dLWp7uNBn3whKjew
ay1V9V7tLn3UeU86jnTz7ogt8t28z7OIOUFl5T7lcOIfrSnBofZwy42c+CPxcOUC
g0KXzkj1ZFEclZ8vZ0pLT2YPSEP+8/OkrmxpyyE5TuUf7llVvN3ZVVdgYPGtugXs
TxcSriWcNp7qMKUcIONQrGypmKgwxePF9UQHRoBw4fL0cgemmecrZPPZjF3/WSpv
9UXKy8vbBliiy8QHD/wMTvZOcpq6N2C0xcnWBUuynx5DF2RlQqn1g/gMrIx/AKFV
RcvVJ2R06xSKv05eAsBP8Qvvg9cKeUn49T99JkktPTLAorFfdf0psCRq1pI8GiVT
gSvShk3tABRDpZpOigV8KjAI7kA1pic4ZN/lu5ANG+i4cQ+0q87jUqcC7IMlIqOo
EhMQGPM4NzWy9N5gZXpLIRnaDL6hUDrFKfa4bfaUO8Cv0lCIWeg1Rinwhx35sCPh
2BK893ilMys+99Hf0oUAm3BN4MOD42sHMSz9GmLl8NxkeOSspYAzrnoUKZZuiKUk
Z6Kf5QqSyK+93yFM/Ak/b+Cfh6g6qdkaSb2LpZ2SHoISR/lUvUDuohSusVAvy6JU
BrmeLktTG6AODDk+XJ7gxEXNeDGNqdQQ0C+DkyT5599xtyJ4P9bypWBh8dj2OC9K
HFeduRqsnbWsY+JZ6VSmUZVhGg+itpJj2Ywbq0Gbw0LrxVRu2BB5FqipjPl03h/Y
lKQK/Yc37oGUxHQMXwYamQqyLs1HAO+zBnI2lXqksC/a40dfcXG3/6YKiaP0clET
J9pB3T61YO85CK2Q6xgDaJ2hyrGwPFPS0SR8kS7f9oSQWzhRPLAIrb7YoE3pmAQ1
XX99td0P8+Sf1ywhlLSw16606unQSpud4epW3lKImMkoTYL+gin0rU2FWdvClizl
LcC51/MtsR8SQFvl2QwbSki5N2PFBG5dwuuOLZWI9YqcelL+xL362S6YEiONuqCa
armCIpftyvNIdV3dDtcJvR+zOqqmLtQiKa00r0qR2NjXVqT46xcJui1/7+CScHZ8
+gGv33A83IvW89Sxd1xsABizhPc9YSsQmzzgj+Ft8Ip6ruIraGhTxDyPzZpDRw1f
dHWApJSDkO9BBR7cQ0QcZwbi17hp5YwBudNocwbCZI5cmAn62JtFZmh9ZFivpiAc
TXLbXMbh5NYn4D0SX3f3JFl+RwzIPQz7ynYlBOICl7cS8E4iUo38STd9on3zAkx9
Y1aV2xp7ibjnKifGWPgzhZ+r9tAAN+NSgZFI5Nv2LNYWT5OV1bgc3Mci0X73vrnA
2dvy32XbwldrYR4f/rthabfiD8cOm0Yzg3ugMrcv63NV3CVJOgfVpALdn3M3dtFd
JGYzzA7M/6anR7KWwF37ofibZs0azN1ZCQyrJjytzFCHGdDdbW0P708yeN341k3I
eowwzAsu35QY7Tacf/kLQ9tALRc8fUbkMKch0CQwkcQ4bttuP7Bp/dKgko2mHTPa
aCzG4m7pu82AZN9VOrNMkAj3EgrXDvCDHDXH8fSdF9u8XEh+6wxB5Ny7pkSPYWxF
TJpY0yMlSEEfnoLyVQSJMUipr5/M8xNsFZnBxPLobj36/U60okYSO7F5U5DhE0Xb
DE7RrET3Yh7ZuKGD/gsHxBcK5VRiZjDwjkFJ1Q41O3lClPZfXy/fDb5uPBL53VIw
SqZxRB14nOA3xCx38onpN9/qoYp2EdUW2wGb3ti/Sm9XCR63qUSLgJFK2HEYiF7O
Zj/Q/8EIfn1OyUaheSMq2fqTTv3VRhAzvmSlDsNoLgoy5ieysxLMHlT8hyu9SirQ
PdJsCt5zm7wYw9DsDfw8aHsDhXrlZ+U19gwFP1ZlzJZ+kMI3/4/yejGxyIeZT/pn
ybPgB9FhLP0+O5ldJQ3MdlrYriXLTsSlY0XYF1VhJZ+447RH+B8kvDQDEFEf/AEo
Ip9iz1c8YKI0e1jOGqNcd1O5iQHSACL5FoGGJ4a+H5wuaHQtv38dqYBXKglDBUyR
VOr+SyRC9nPuZ5t4dI5JlSZqXlWBpsfabRCoz8Wr48Z0bPgFPyDwRBmu3ul52Das
suBM6yQUP6jxx/NV1afOwwjArG7wonc77SJxdClThM8PTnaoTLB+g4I3AAxACZfR
nNtgtaGktUd65mLIdieyM9IrIbHI7GzA/jHx2NVvfZAyNpQhzU7y+lglY5TV2wYs
zHA/PA9heM3gciQfd8Pw8VXycUBp0uXur5eVCRgYXiXTBzMGaEhQ99XHpS3IPSvS
gLexi+E8aYVoExchg9HaK2CtZWs3jF8ldewMouhdMjIuzRWPYz3Zqsb045kmctWs
PWv2xQ+iSs6V49vXRf2Qbskw5NXAaS/1EskTh9uhXs8VJu39pF1fqT6TdnsV/1mk
wPrJiC5KMaZLpQmgwBkFxDY82Zay7Sv94xg+aUF5tsg5gWjFU+wXdLCIKEXXSieu
UjR3vh13bIaA/cYdHFZtHs/Fj5xduXj0wHAfrk7yRqWXaPWYJxG/0pUSsduW9e2e
eE16ubWp8baZcGesUoxtqmAieRLl0mqiN43X9QQkEVOoRLCZa+Q2jKQkCzMJnmwO
Vylj+3/8mnYpwwmGAS4pqw1eQdZjg8xTKeGskXqEB4N3k0cY2P3R27otmfJagLVP
YaQJ9W0OT6qb84nCG/q/dnwm0wk4ybK7itDfKDDd2dqQ/AbVe2wSvQhlZxYYulLj
rz9fxTV0rUpJn0qmSR3dnoyKYU+Sp7ohTmSmLOVl5uu0Ph2C59qlXbKLqX5+TcdK
lhecrD3RsZgos65EAgwMoe+tOLVmS935PHnk9c4ilZcZpfdvQUuIS2oRuRCxlSD6
tFJ4BiLubZFYkHBjbutR6y0xYtzO4HOxXv+ghjlZciuVrKKyvOd4ihM723YJex5C
XqM5cFyoRCw9ql8o3FR3wLLTUMec1PIT76hxrg+fVbAEZLK7AzGPytykIAzP+0jg
LNzvUbweIeR6y9gN+ayLa0zQtjy9YzOxESAkjmj5SMgSBMWc10fvZeLUCLDhljx7
6xRlfvQepxJsprZtthpfODO1xNS/NPU3pBMwc4gV4tws5kffiPdjHz3gxNQDcCOW
zqgCNYWQjYUr5lYjSX6xP00TePEXV6F0uE1J8pPpQ8Va6COG2Z2Tn/UBzHcRL8TL
rJzS0sPgoSjEofjiNKu3L4Ek3DRtCdAdv/CnCiJNtU7xc5rKWNY+5/7XToykhW0B
2tavRx0wizZvq/pFgWltCUoj4NK1hDzd1wbMgCiufeps4dQh/m5f1cCKo2Ou9tFB
ZHCvgdGyDzVx1uqa3ZaizGYY5fxeC8pqrZWpTyX4VqGlKowOeRPGPfD9kLTNHADZ
BHS3wejgQY9QU176DMzFfE2QNa8/gCTw5Nng/tJ1B0FCr8zutUXohWsMHTXGrJmE
0F49DoRGodQ00D4TajBEXMgxVTH3t07Kw8LV3vt9gcrlescmekeIdBF4wAq1b6wJ
bEB4LQS7RkJqXj7Q00Nn/5F2kH4ngU8THq0zzlNv7SRucYkWJ2dMKgnQY7UZ8HS2
eBgnsnt0XbfNqvj5d2PzXTJPiWRRbqpWkt+OM53LqwLilVha7HHoVMaUmCF3MVae
gV0ngC5kbPRTvIsylA5XVsrE/AXthoWFp8U0TMZRMDE0J9hVVcf0kvuQy9evITRP
j/pVM6PejMYCbMLmwdDZrudTZHdi4UtNzDcPHxpRZjjdfz6PI03IE6CeZ/3Rufjl
SJ6iANEM73UIdI1TF9QbG6TJoq/lZiA/2Y5ktbHRC6aG9DUxc/ZdXdTH0jw5l7s0
UQiXvc8RctwoUMCuIFa6wo5Fkbm7cKGSaWvmU2cenUtaPxRoaOVYCCr8XFCidlRS
phlEc9CAJblQpXcx4EmkA7WLVSUHL5a/GNEOZayzdmU3lPmEcWb4meA5ovRvgLka
Wk3MDNq8gQ47ectb+pv95OuM0ZpIUalwcKJdW11e2zCbNHIvpjcY62drP1HcsPr2
yCMF4s1TrYZTdhnLQ4oYwbWueItdXA3ObAKr1T5du2ptV8FEZSOzO3SViM2V/YE5
yMZj/b5mT3KKNtOT/sOWSAIgYua3atceGh8LJ+GhvmPx4056W+5iXgAIVAqtF5bR
fvbhsVvclC2lSQlrODcKYcC8sE1j+/I6TbHlOn47S2NNcB58GRlw/mHs9Rfe9KOy
RooyjkUAeGDNzgdJjPtcrZTkOCdK2K+FsG+OZAdjBePwBU9EFAxCmWcTxGlT89in
xFZcu/c1yN2O4SJSbIm0FZRjcOdlCsNK32A2REA3hA5Dv/MRfjRjZP9Kt0/5EgjB
UW7dJimc6MAS5SsnCFr3DoYDfh4v/VSWWHUk61aYAiN3tuU8zwUkmHBr94wKzwn5
Lp3xBI5O5Kmg0FtkeM2tVJXoiXJQ7UD4a+Hj3pKtsj+aMa2eNyX2Hhuxks4nq7SH
LpRm0OEDvMsrPia8ClF+jQyR8JwFtcMipMREav2A/OEtMCduM+nXMM0FtCWainmf
Di1Czj7r7cM3d/tOvELnvWEecSxyU9pOMPQHWGnbQ9z7Q77pnYXJVJJ+kWafrTUM
mbx49SqZIEoXd6RCoMaIYxCbUU2SmIXKDCTSCEu/ft4qbn/rwF07jkrFzGGAsXvp
oDnb6S/lExYZ7yKAkZqDrSIzMEOM98PE6cmDu5Vxu15QUDB932hkTFJSOeloZt/4
dSEvJLgFAdIRlY85N6QVqvv82pBXW/SsNva4NG7tbFRuR2+NHB2xELiuXWJEN8ky
RxE03PKLPrTYa+JAWbyzQbJ8LGNTJjHhLNMPFzhU2U3bOdf5dGbcfQtkk0ZMd+Q0
KCPLF1BmdSyDZgfjm2KEjawMvej7hBpfM5qLTiaPfw1byJV4RWQafcEYyccBpKXZ
pqA8gBZY7VP+5ueqMotSdMAQCbbs+t2i6cTYBuuUlyN5R9f2SmPTUMr9cg6e7fiX
AyKXAoWP4TyFuaxAhtbXJ9Zk2u940XGYwBGZ7n01hSnSgz6NxRqvqC4fsatFQnJ9
IRMTEtVyLqbVVxGrKN/MYJDJkPWvDEMZG/eS+WvWhkGZVS3qbW4PDlrN/3VKB1Hf
NXQdKIqGy/WaSxobzzfN5DRefLbQhEQpBxLMVz4RaHp5dlfJHvMjDpj7sApUGKap
AzdwLFwXAx4Cfh7Yb5Eu8tCi6cGILM4E411vJEsFNDfhj6EDEWKwzt0smWBbjzSZ
rtVX8EXAtJ2BwVBB4OxCNmzX4OzB8VQdOSBpQqoWJmX/1BFczl+rF2wEEU7+xiTi
Cf65KZPpi7Oml5lh4w7mbP0pS5QICgblZGpKetJUAQJmIFYquusE2wMQOhYK06+3
25jg5C+qPzXqkcYND68c+iTnXYaxXZTb3EB0NU5x71uLRE58jfkpJFZZ4MZ41m4i
o/YBTXpOwDvcU2myg2OSvlnnggDeLu1GWU6v38uw72PWXseQBA2JAfap+41q0M7h
V/pl6YLvlabw+DH/QpQNpP0gTGb9hrgfZTVfOsn6iI+YynRjD2GAGfdf6airqIRF
kDHKou3UvfR562YBgBRVTc1gmS29FsNKHXuu3D3mieI7Bv1Al2yetjc2JpgK9FMK
nfWWr1lSq0NJA+Beq+JUiFDkNR4mXI66UhdGTuGX9OJKrZy6KzNwCEh87T+WCIHH
uygBJXvztVvS9f07QJVkGjK2eUBstsZWWi5/L4N+vy7/jE1/guge0YMZ4SsFrsIU
8jK1l8D+qgGbtGS9dHanJIqi2Qen/Z5IV7TBzZukqX+wORgP8kdNp6sFsYkKcTYc
nXovHkdLMR2GhhuFwyrwKPF97y89ayAu/9st1K2PRThn+lUPVT0ZV5Gkoi5UkxQu
i48bwxznmG3YNEKY+1cGOChLMllTZGxQ/g2mWNn1sPoLdx0oowNz3XvS+VTwm8ok
iJSDsiTdkVrGsX9S0GJNSoOUlCGFb1lHpleIfWjF57sQsBK3l8M93+wXovJETxsQ
UJB3wn/bEht8MbUOIMb9gxms9qdNg/D7TwX5LRpcufeQpEl25n3X+d6Y0Pr7bACZ
PsE09PeHlXFRFAu76kUjm7q7rDFqDReNM0wQT3eWCN1jM4xmS+P4bZvMzQZpBnNz
t4qz22jyaNeJdccSUmU8LdRDqRkHhLESFFKzqNdEEoLsEKOvvsG6PuHu8deGsJZd
cC+NGaJSAti3cp72XHWrJ8sX8Wj0ei96d2yQaVedLS6MDpBhhf+qOr4l3gwkIK71
lfeNZ3kPJAFxEqu8/AkW7QcEcXuxgvuh7KDuH4ejIV+PhlVvaV8ZAd5u5A8GpnQY
D+3Gfna4uwdAVdfe7bB09dzP2/gyd8VzGdJ9RSZ7DC3WgkzCjh15tDljKlM+biBx
bsHnIqTmEYZhdwv/GaZBxXUZS/N3qOkJJOT7/9oYqFiScdsEGK2xxt4D1mEezOY0
YAd594M8a2za6VUJqqZFXsLiDZNKkAtdI3IpxvK+Fvlf9JFW6wBF8zkBN3K7nZzD
71onxywGx0jbrrXzI/Y/bYICux09xaABMmCY+YgqbMzZmHpPM6rdR9KcUVYzFsgm
GdkZKozzbWjfaLvXmQdyhLB6YRWOgUouxKTy/me4u2CmkKIXIz04EuzN2d9N7H2c
XXEVzzBYJcW7ZSgqVLe4MphWPIlENZ1W9HJXWd8U2ZcGxmIcLktQKgNW+4HqTR0q
8Bkp97fk1Z7e1hNGLkYYx0Kg7VF/2/JsaxLFLXhnORt8Vz6hQwFYbvj/Rm13FYyT
5vH4dWpTujyGk5rEpGY7E6ufVhUimOuMbFH3B8UpB3xAFNPNTMDcRWys9alKt2xo
oRWRTCP4Tmv//qmFo2YTNaYc5CSbWg72ri73gZkt/a3ML1EzFUQ+/kEIYAlas0/f
LEx80FJA3SiGIz2XQ9EUYuC+/3NT8SwSMLalNDqPdV+re8A4i6iN8isP5ZSBe+K5
OpIR/oRaijGS07+3f1xwl9XE71fIijNlzjfXYn3e6PitPteEK2u2CDfhFKPNrcz1
2PkmbQJn+46GAiI9i/o8BnykWwxWo0pG1AfybmlSDCgu+YwVRjZmgaWigmyGudh+
qYii+fyDJ/L6KiF3WaPzfMdLznbnTJcu4LCPNzW7Fj/isd9o/m6MovXXagEAV0rO
yWmBwT2+/Zx5iZYtyEaPkTU0yb96ZBYCWmY4OQtVaDhMP8yNIbs62Hb4ug1VBYJN
V521iYgVVzejpkdJfX5HhwtIWI+w2MsH6LmGMn9ulCd3iSv2UZqQD601C3fL+7Qc
T7ne6ha/guzixH5uOkPLnDyYPb0iYgEuQfs4SZCNRAUtXbiUL80YAns7CMFzP3tg
vLc5nUUKGUJ4/vulh6vOs+fdn/pTrSuf7QvwA/w8RAId20Pc96mUicbEKEZoetI0
qNhQW38BboPZa832ydwGZAULH2fsB8pqYlaaYT/fo/KmNPSQ3c+z//eKC5ZVA0jl
W9SxeQjabgNozn+l09LB8Fj0EA8Y6vUi7GCYnIrtU/wquFffHVDyWnCmv6wrlrkm
/Xq+SBNbI/sl8p56T2w1i1Uk89uDkzC0hevyFZwlN9h2IrZMV7YiYgZ/dqKKlJba
AmbvsnirrvFWyE/T5Q1kGOhKabdoKjtolc8/T5DS5HCmbmyAvDJEcw4QwuP/5xlA
00pZiG4NdrnsWw+pmmEAYbA3TJxR4a5wDgoeD4YdUvflMg1XAdS0zTAncau2PhQf
0v1Z8LozkXIr9NT/QB1vsszGRGUatQ56W0iRRA87NFK1qlmnO2MA0M2VZLigQ0/j
HXfROKYAc6+vuaqlqp5HDuwp7+qzOo9PSI6HW+H3HR7KYllsvG9LMdibL/iib82G
o1KuvCOkvG+Ah7zJcTXjj1VhU3YH3VrzxxNex1ITvPmsOSKgcVTvSQRaiB3fScN0
a7UeN+DRfZ+0FZ/5p6RjYLR4K1tTiDBB+pdNrYCQmpg3cpUiFsRZPG0sIdqQHlSf
+sMEkB9AI7uadNDMHvO7R/kFr/XpVRja5QuWkSUXNKkhyNIY3JviK1iLO3ttFd9Z
eyuJMkw7pcc7Ee4jtlBrGN4jjaxht4TQdMTvWksE+aELc3POxSkrBd//LRmV0fWz
B7R4ZR3D1DdmAW1rUv3K00AlNVVRKxobRrTCZiPRnN0pB9R8bM5wOb7otAquJR+y
7CIIg09+0fb6NPJw8BEgnYbJ+hZdyHXenqIjo3q9EFZLkm/umjWIhtH/GQS90eDF
/VuhlxNM/VAGC9DRRGhyZKeTaqHlkXEHe9eYdKSYL7brKWI7cYc+qgts12vLBmMO
YDyoMUMeKkErAHPGI4wXzUuLyp+HMe3tKb/8byF5MY84Y+2MgCuG9f+Gi8H0Z2i2
2yJ5RIst8L+L54WgaObJ/Kzf0L1gxQxK3Zx51PvVPrjatl8McQW9PeXl3bpnUvzG
pgDTzTzv/2Vh3+nxiSCFMeF3Z6XgqnnolkRsAD7KW+GX9SjPSxGB0M0yIAyLjcUf
Fwy7R1/d3TDG08rmjBJcMkPZojmzwh+/f7BoayJBBdMgYrDqGLZGwfGEnrls83D7
S5nMcseqYBw0Epwv2Naw4xNEhEEqt1A3bdOyT0T4IYLMsCZt6jiro+nAdhOHVKIH
ju6mZqbZIKo+Kan/Hll5BJvVjaxI8PLmLys7zoNulEBr+RJM40qZX/VWLrQ8y66U
VnkMHng1/z88FpXla1Y8cSAhSbrVQwC3lqV8iaMAr+nlZL76cXAO+PRHvcVA6TAO
hVakZTtEfReOtjT20Oj3GsFTCkkP95bvmvFFbOZ2BSdhqD+SVxf1ilXD23FCPSJ5
gahy1SzjPTA3cjheh5E4dCMK65k/gAtXwcpbqUsOxVKfnSOb8kUO9r1zfCftN6oW
TrKut4rgvj1t/v8EI1yZRS1Lp/Mfe+xGTxIKrer8t+8AUAQGU96xIQolFPEuGstQ
3S//Lf8AjMjr5DCcAoNiU/JtrPZfOQK8SslCRZ+Mz7qnMala2Dl1FsztyDnZGONw
3gijqGYHUny9pwazEYzvIugLs8WbffEzFdCA8kJXnEIEoICRzE8HaTgelSaS8ors
4LW35Cts91/iA9zHm9v5sNcodEWAXYiNbftu+B/LdFLYgZfYLabzR6l694q4p3Lz
Q6IiqBPKQZ12f/Z3UaesFo1zkmjslhtuk/i1bbCK6KQmENBBTQufWkZlowy/Qj4l
MtLkHZ4V5qo2E+mTy/AEXzFPRsD8zosghYdUVSKx1Us4Y30CWagDiqJRjamdNqHg
OH7IW4k0sj4/gTuxkDNQKEi9WUzjePI3NCqUB5Q8B6JnokgjVPfh096KhlV2aS3M
co3ioyOYfJgw+xjZYdSSBgC2FV44wt5OQSY13I1+tSxKBxgWaT59FNKOzAUA6+iz
4HMm9EROkYui2vMjpRmWuEb538UuKvyt2U2T53mj9XX7IXeCndpl31p05u8SExeR
gso6mFbfJ0l96Qf1ckmdATgSdn9qTefV/vouxLYkYRwEWioZiyraiTsSf8HAS8BG
PX0GBxREQN7lpG9Z13ZS8uGwCY5XtlQ+niIGvUZhTby4m9+s5pxAk9jz/ehkljzO
uYNsZFhaBYWtiiZwcJg0zTb+KeZ2vn9aXFdnyMsyQkzPu3C8FyUtqDCW7SKDcgBL
2CMm8gV3GkkxWeRnVCm+uxxTuplzM+uTAY62YpV+Ick7oE/+GX/Fl6f0EIuKRO/c
kUHdU00d6my68KXIbBy48FJ9CvUBtZ7qBeLXo3MwlOVq/OYmVNBqjpSTRZ8lelgV
mJtCPpn1J0IdNJjTSQ8PBe2Lr6R50FyVRzzMairL7duSCKW3/MGXHXlu76AKQ4/V
GT+hdkFobdk92QzhO4BdDQiGHz/GwHlVS/ElM+ePAAw3AtasWUQvau9BvwvhlZqx
jzDchvHzhG22c0dpP3Af74TRmPHworTYthW91MpKEZC3TDM1EFRuE6CMiWFGWsy6
NIcBbEfk+wi8sUR+jxQbM9WL4+bxYxDEKFmcOI+Jp43nzRmSCRf26p08Bi1hHdKr
ueCURN11iLNBilvZ1h1oMO7eqZcA6jWTTR6w7j2JtX0bWJ5Hir6wCmQdCJE8urrI
Zs75ZenPsxJ8ysQR9cWg8GeG7S6pztgCidzPLEnKvdDAFmfNxOOxg/3KDG2XH+kB
gkcSuXYoO5mIcwK+XqjXxOeGQ3CmPG4HRTCQTfG296XRjVdLFf5IPzxhLH8ZPFIW
5tKBzVCMIpoT4AG0fRtAn3cXI/Pitbm/posMKbgji0EmhgFw7sX0jDlgMznBynCd
iSGhILyL3CtFFwoTDv9kdWWX5cFOjetowH4NatHSVVHLOpSlZhUpScz6Ghn+6ikJ
tW6QoeGyAmEUIJxvAZUM03chZptliUSZkXxzy95J/fc+oAsV2yjctFOG2B9upmlU
QMG2u1sM016V+ttgPXyiJeJNZh3v5FPYpR6EgFe43gdnAYsYwfXKbaY1y2++UdE5
Ot4WnNco+gdU11mx5pWV9gkiCYKEy6e9pe7xupwx6uiZl/PWSJj8BQpGZXDUphBM
2kdusUh+43ZnJcadSrdWQ/8+uFaI+pUe1ZC1us/HFqUu3VI+rP+qlJpLoGbLcgpO
2JGrr9nIprn5EDRrQjvvj5b3Cu25Ngpt5LBTf9svWBadhW13AFipBJFQm8uNOivz
MrkakxsihFu8Ws6nNp3wYci6XbhO2HDW3iplW2Q5vPx28BvfL1u4pinCQ8MM5awJ
QOGQqxagf37Xcrr5Bbo4YsypjRIzd6RW+wvKoSnE2iEUb8vPNUkPKHul5FvFPYcg
ftMZdqmjxN1KTeoy74UvJP1PmSiD+LfG99rHrDCOtHmhOgNZdWlZPdf+uyndXw3b
ONkGgMf6eEHPqwWjuAb4ayofd9SB/+NOtPc0z3zZA+nj3kVuJnyvlIy8L9+FMXUf
cOe6oV4oN8x/SOAFmkt3FQys7BWkMb3PHnCTtC7vK/gv9C7F7cKGdC13YbE/2l4B
FyRkJpIXgzhwDOoGCv+MCUroyB0x7DogRymVl1vvtvsqH+Wmqpi1mSGdv/VOrBuR
qBGI+Y509ubBr7ycHhaG6crZcEmk1Gpm0nvK+XlvrIr+y0ydc30CV0lnHHmus438
o4gZgYJpaCIvgfm6+MSNxAPtbTqT/r8tnHtBy6N8tuNLisrvA4ygSZPetUotgnFH
UuK0mfDGkPlYRa2Ovj5wUM79zokwDphtNAbCVKzeCf7Gs4derCUqguD7urv7Kgez
OF71ZoJHmyZOrE2W+4RYa0g6pxwZ61H9uocmLa38lM5Ga/kO9lB4OIUwtrc2l3ao
GJNCmRGIiVk+ENvalC8KteFBK5EfGM30fqPbI2Cn/pCSIP4CBo9GcBIYzIATwSPY
pWuhI9A/6LR5OqDEaGjhVYhRlqoiZe9oO2yeDCFzxX3huXGxXQd8aMUGZjVAJE0Z
gd1M1rBAwFgtN/2lnaHvmlwRKKQZU0EylpFVrvldJziyD0Qph0hNzVxDFJiPpHxT
7NPl3CbbZ40Ym06NzunQDeOIN4+jikh3UAEGbpZYDN/TZH/L8YBhZdz5JelXZl3D
V4gFhRFo00N3g+BQ1j4UMPeV9NrA1MiXaDxJO0oBfnFXQFtKK1nM9qQaVc7o8SLm
dbRC29UpawVkrYDfZsYlGg6qvqGOy0XZjaKZxPZ76NuIEJacvxCAM4oxY2Dvb50e
rnvZh9O2xzCQwzaM44sJmMXmAjSLnoP1tt4skLEKi3S0OQSZLCb4CqKQTxmf46yc
n0qChdMIUHlgqPurEe3P96NllOXwKJp+vSll1d7pERJg1ikl05YQd1XQoBQX3bhP
hwO1dNR3JRSYQB7sK1R3vM8tRBF86Lwh2ZQ8psj0yldY7Foq6+hehCj/Yjsv/9kC
2RMaK9GCdJ/DFscAqPu/L45McCoTxJVDgHDFssOYex4+yq36chIcQ8ExDjNyG3EE
4Y2Nz0CwDcegzgrEJggpDQd41JgnZnvGDZA3eaEhB6M8UX26VEok7NUQYPJTHvhQ
0fnzYvt03vY7n35PC7occco4roeA1mcqGkNRL6bL9bxdGkyzO8hzmNRnFsES6+0B
KCOUDl3QCadYoqW1NY8K/iWO2voFwJuK4KgcUZyGy1zFVgk6TyMw15sgt3BUy8hw
QHqIjh72e1oHkLpXJqcx6LQniXB2DdR0J3vfhBvP4riANgIBt5CmxQ6aKhJiwLBg
JAnNu0u4/MHOL7LT7tP8OCXA4wq4J9CnlpZOse+sda9dYDH/zSX5j6VbcwoudjgB
PUGikDsdFNGRYZ/wcrZJLePyDiT3vZj3/P5S7gyTtc1SigW4qHzicPSIH9IWlLL8
vyR7zIAcWfrUvHe+XAMBH9UCDiE1XFazPrKHJsv0GXgHmhZDagHk4feqcJ8MFvij
/B+3YVIcTJnUwYAaLe+J+61DDISIeCYMovkJq6rdmeNNQfVpBHg6P4DzKqmcu2RZ
DsSb+8iP1VF3I94wGZ+6l0ocyWggQU7kKnDpWk1Owa/b1US216apLYBbMgs9Aerh
xbF0AsjLVREIdpSFgn3TiX8lnyosET/XKUcvvRtRZRGxW7/x7qiJONopeOzYfb23
eVk4+7zBsUMqTkzaUIUN3lICNeFB2OlOq1yWz1+v56TK+7E+wN9E5krdPLT7/XdH
MAzZurao6FPKhNPLxarjbx42RrDD0Vo7tBGM7hgw0GcbKh/K/sJMFs+a9DTV7eN4
1u6OHjF5xTpFetKtNqhJKl0ycf5Q6B/k4Fu1a0okXMgvyw1hj14WXoLVgPOT8++r
hYcisHYxI56oEw2s1X/e5pXFACt9OowjJpiQQZbs3btFZ7FUB20MkGqg96kIm6Ju
BBbvkVQGSFxFi5uOPl1Di2XXOSkgfDq2dTYBCrVC8cNYpcAb8aii55ixcJGsLZCS
CuEdeiF3PAdci/gnQZpP/SKVJXREuznZCWFoSYmdpZOeaFP0BMZGPKxny9tsmPzH
uK+cq9EuLb8gDmfhsilEBLNIsU93zJBSWUI+6Sin/2nNEWvNrKsxVR52Kbv09gQs
mq+EOena2aa+34RItxG+GZiQKSv82EfFNM7y4eX3GrWrfd489ru4meubeDD6Ras5
3jndH8d6gV8WqJxubh3wKVj+CIutYTM8ZSFmCh5phcqdp4LON7VvANJ7Ut3jH1Rm
ucwgc646+nNZM2I+ZtPtNnlj3ve0r3Oc1t9Oh6Qco6F3KclPmqu84PnM5Qb3TdB9
cl6oRVCNfBX3j4/x/yztvFkgJMPcV0+wBHy5HMayTOt0w2FVArfP4gMc/wJCwHt8
98sXbPSsW9DALt6WVf2G8mGwgLzbAODcZ78z9yG1PYMAR0licYlU6Ub3Qwy9+43i
dHQbqiDwOhvWrrQ65WW69K6zT7Fu4261Q9ufUDGYvrxaXWQ7240O6yWnquRn8RPr
/g2n8XKv/s3kUgJ2auL24L+wOZu9hIUY14gzjFzOVUOjmn8MBrBIlZrS9nBmO/c/
K17lZE7kA+uscx2xl3zm28Xfmo39I3y2BcMCnsONYwNwz4a8TWjFORlfZYsX6qxc
3ZS8u9e12yMqYZ6BnDRxfnM51WC4+DtlZS0WM043i7dIsWrtnutwC27r/CF59SZp
RtNIb/F7nHAG/xAkg75fgdILLoM3gXgFRa3eGEpgMTKinub44Y+n9fiB07pLswPV
K7QXAMSy0D7xNPTHmxcDP8SnX/z8oBm84qZWRI+TMg0xyNnO85Bqe/CMqEy2bx6f
8Otn0yiLgR5kryqxNtkEncmdeSP+QWqbsqGzOvRLYtbRy3Fs6JEzyCcYltHKjLBo
Pas05ETjjwAXEaIZzWxHcWFnr3S3yEPh+L/UE57ECqBebyye8QKlcBbjUc4Mw0EX
WCpFB2eJsdMSUBjnm1SPjppRUPyH0LOX5wYyKDgAB3Ckx8oI/I8dWnc8R7wo/CxA
Zenozie83Dy26hSS62J7xwrJI5MAyFda8P7XzcZ1C6AVysi2XMDR8kENDt/NY5xT
A1+U6CIvYl7nMR2qAMFj9lY4vCkT+9T95Lf4mYG1gj8zBHf1YL6jJwCphCRQvwkD
mU0kRiaelnNU0ndq25wBCcHIPlFSpTQMJbUw0W3aj7Qk37t0Cwpf68tFn3MjZk+U
LnZC25i73CKWPm6Aq4flTWsEWT2p+MTt9jGvqWTmnkTIVz+2uUsRCyK3dSwW+mnH
1OIqgW7I3UqyIPs4fR86pvmefuDgdFIbBsWCnTQ0ZlsYMByDId/PgUeltgrV02Z9
HvMCDrlbxKtRqc3TuLIxdGVlZJA+8kUXz4Lk6p6lzk5IFV5lsdF/I3JjHHl4/Kyo
SKTLYC5djqRKhO8H9gd0xs3LZWMrBZFEh9/vRim5TECY9PvY2M2tzZGNCnzLA3KB
vHJhC/HshhBotUx7fE5WOipQs6caCbtVaLEd4lotwSXAa80vu7DEHVApCW4IB8g4
/+kw/8bTiPJX5klSj52PsOpyrSvuzzN7/m7/k0KWWSGOZHpo/2FO6vnIX4U/RMH5
PMOAdWt9wSwJcB5OzSZSSHN4AJvmtT31gE4GD+nRHukL0EWS7vJCYE0TDKZDRCKZ
qna5i9g/RLkR4sTD3WY6XoJYhT1UZ/iTBmo4Y2PIuUhdfp8DvvpjtYcIyq/M2Fd7
1+hU7AFYDYtq5OpbyTuy1T98P9KPdhG2NhF9/oqu+vM2IiqZsdyE3sZpRdNDmkou
k1LZuH3UU1iGbvossr5r2+myVSqpEh7PkqRebU0zASew7ipEEVKy+0/S6+2d4gTN
DDkMK0on+UfyzrWu+3s9d/JkSwvZofHe+mHjwCIY6gHI77TnH80MqNJla/+Hz005
ipgA8Z50PCAC83iQnuet66F85ZKSlTz8wJXOL5doway23JXkyFtH48OQM5qBzNsl
qx4uYo2I+AvE9P208BH16WNFqozxpGLWGFnXsO1riAL05gqGcCxQKh/te9ax7GS0
1Jm7M45DHf9vqmWP/ksOjIlpHRplFofOQn6NZB2SK/wMvL2P+WbmX539i886H+PD
bUA83kLDPPnaBCsnk2/p5tHqdRqTB8ctITAX7vsL9ctheKm+As3rs51CvekF7b1u
3vtIKHYrKc6oQPDtn380gXieh0/LtV5TcSMooI1MlYzKTde+EzcCXsiRAzrOJjrp
S2HP4V/v5XjDzZz+3nkN2u6yv8gxZk8V3h5xxEnvAEDk7QUfVcUf6XcZovH6zbti
9wDNnGelzPrJbqI7hRwedoBmh4E5sbbJNl8n9bua7/lIajhXjIjHD8t3y5Y54cyk
lUf29RSK0Hwv6fI1xFKuAfpZ+cx6Rap7TlSrYnltTKpsP47/oPnqlj9lF7foCprs
uwaMIU0rsZ++8lyHJdewgZmiwXQ0t3oOOOpxN1eb59pKdf0uLwbJixJBMWDIPJve
644hu9I4A+RzmLJgqwOQnr8eLQ++A9dNyw5wGvMmRj0yYTffnLSAGxwuUIkF677/
m8hASNR1acGz/6XK01VB6wrCPIAfpOAwbi/5AGX43WxacE/S/EZ+8MxH5xQYmaI9
27c6HcrPRZe8/+9PSQ9FuW4gEEFTBFfDQBc2Quwf2Tbx+JCD+dzkboq9oglgIqiZ
+xmYGbGpUPX8gWiCN3YTB4LOv04MAqG6f/K4m7Xgwhd2BpJXqsd0t+Lhpy1NHPas
ey9BsBSGaB9wLDrjb6KXgZKXhm9f72oKNdZgyBXdkgHDgAwuSJTzJ/UajYQ/d76t
fTIr428rRnszgWsqZezbB7ucUGrwOmLpT/sGNL2teSRe9CfrYT0cYl6epi8V3mER
7KSPojZRhWRJvkNT+2CvOf5Do1AiIACfwYLNBLJTEWyuxSgE9jr7bELcqMNnHOWi
AmStjVqeKTIQqtAE/ttijLu/M45ltOm3vL0/7MWz0PHohXYKdmkF77A0D9k3Kzd2
B0CXXLn8sDuw1Aw80AjhgOLF6Ps6ihsX+ZGMLjymPhRfXIAHhI1u5HkJv68SB6ve
3eO+ipqG39xowdHqV3c4zlkXyAZUOp1g4zTCQuv+UJHR6dSmWjL27R3I4tYs65TK
u9qL/+HqjCyHhCKDU3g/oqs9wuogkfTs3z9YdbJBqbm3oLuSy/9H5KTKiQuTHd0h
m9qB9Hiztuy8sSv1Btaq/SEXqG+Zo4BNBmmIA1pEb/NNPjDapAq6N+ZyBf35L5km
B3gVctNZzc7ArP1nSHwngloErWx6XS8UpXSHUcQsbpV9yUZc8mIIuHWNjpZAFGz5
USCEhlTfvh8RsGukVI4wzaILDLLgzFu3IKfCUiXiHI+VZTorZzoGTr4C/SaWCOV2
QCzADR6iFCe3YLtHDUQWucke8UyMRm/0ejVc2hJntXtRRtQJtmv+cjBccszEpGM6
q10cJ3YPBiXT+MvwK/pwHxo204eCG7s1rOY81QuhMQvI6F6WlBISE2TvxV982bNB
R6u5jKTYPxTaueNkYDPA+SuxSZFotKBwCBRuyj05R3NS0zAZZLsgsZhiUiHrN/bF
ED1nJS6mfJ9jTvvGjr21sgyymaKHYPtqHzIFkgQognOlzOjwCsg78bHILWW1KC1m
sWrK2etABO/enSZxjYSimiqzDHPHoKsEuE9T0B9A+okm9123Ic40WOj9LEXtre8P
UgitYFcplIUPufSyWSI6VBFHoU7mrOw6pZhYolnqd14NOwcoVnjNaptoIJNrSo1O
UjT4F4f5qhNxM8OEIUYoONP4ZNEYq2h8XKMz4TYNfljfSM6afHxLO4KEZ0+NY5Kf
FTkOL+SIwh83JToq7dhnObPpi5G0h1+MLDPqGN0/t7xJifLbagfhLRLnzThdQsSY
Ieyi89AVUXDHmQd5lYSw3gtMR9h2LAcVDKz+szikPyKT3rulxJW478nREPyvd8GF
jPm0SaBH/DBOjiApP+B8uz7ucNRYgYqUUvHnUIR/k8/byDPdvlMpBmT1fGd6K3Qc
dIHXrNPpSCqMeobp9XZWoVeZ/xNDWgXR7QdT0UNhtiA2LwAiW/NFvA5Wx9X2lMrz
uz4UWD1rTXYJsYHV781sfREJIjKGa7H00mZyo2jSAK6AnpCPvrMB3W5+HSUZ5VCM
6c8zHbbcYgrkkSC8WHRJV53XtXhVTEP19HQIs6gj9AnSzPHVsRZebV5k4vkSZM7g
NUZwl7wIsbg8GyMPb9XFI2qMEzSCfv0EgHAMYgxHQS70p7U5fo8ZakVD+Jzhq/kX
QLHZX9zqsG6JDN/P6NpiVt8/NwGf7br+TULoTFmpk2EQHsyvPYXXO1nYZ+LrYTuz
MRfYJMVYcE4HGE3BI1LjilInwMebZDTU1ErIR7aYb2Cngw5X9ynzUGJFO6t/KZnQ
7g7V41AWuo/j/Da3HdQ06MLwG2AGMMp8H+f1/dTbwLfEA66wQcqScyDzzjE0QYA1
tkLvL04WB5BDnDmimeCj1YnN9xW+rzg8ZyBbOdbsH/KtHi++e6c024PIjQvekHkL
eyk+MY6JjpHfbliNmHsp1flS36MErFYdEUbp0tivesIoR/+Vbm/sKgqRbW/wwjoQ
4TG2jVRVnrp7hnHTNnCNL9wqgIRMYKL9oo4g19tuDYdpF5EJfxOXLO83TVvyHsnN
3+n9VCUqWLy6IG+Y1GPI2l+7xPIw8UqMTTHY0vLgM2gZk+m8wukpc39LysRZkr/3
/xFe4Mz6QIsPZRRmRFx/GPQ48RVLmrQz2qtBFSiBVqRVT2Ru4j0Qp1BFcay4+dvN
3reEm6IHGfnwW17+BW0URr3ZHjAD6uaF2jIjUn/0H3/fDYdsAKcjkx5XazPSY4TY
0JVWZSwHV9oztVVG3z2WQGrQp/9KAX3njqKzCCaG1dD4ElqSpCPnnXfnSvJ1yR7q
zeahyK2DKciIYi6PtVvApArOGxalCwOP+o8AYOkTsUNZA+zLC53a5GIC9ajktQUN
Uq+q1fvFqQ3EP5Z4QSxZaoEvNih4N8ZVcPSVoJltDRGLnkSxv6CVhp4MZGOM2cSn
dwkzGAgqnxq6xlz03JKd16Z8DDVINGS94J2aZRWzs4nRohkxK3ceotbwIbKd7laO
t21P5IJ+6tszXImYDAKu0WHxSMDhHYVQTUyUA7Z5dlHjyLl0KGQiiWEcTO9wjABU
5jF4IzVW5J1oLtBA3CzlBstFajCD2n35SYEbt+y/dCYxg10fzGnXW3w453WgQLbM
JWj7XQ+rC2118CktI9sgRYGK5Vlpir92zTk2sGF+rUaKY+rc5Y3+aZ/Ubw6vlMiY
WXFf20TktHZShvuDw9/tgpX6BIP7xwAKN32tUBrXX/QJ2YyQTrmiEpWOx3Vk2LqH
fX/X0sAa4eX3uIObzHAr024NJZ+MrZ8Sz25hbd+fb/kSYIgjemuYycAKYrwYr6Ty
yQ0QKSWyETdWMYAMpuT7it+2UccMzHv73IswJMHUGg/Xx9ix2aCbQwG4jhDal2Zi
CdBofSnm/e4Uw1WK0lcUCouR7qfhMH5MaDGsuM8wJWVG7DIP1sN+2MTRjHNRCp98
lHA6M2N/sq9gQjeolG7d+xLFaOJlr+sumq4JwzC1tPR504UsCtp6zlYJjKGX0mOo
9XKWh1MSWIydIa8B2+y1H6nb5o1rNAIDGdZ19ufsE7KfHzlo66YSxr1RM+jWV3V+
NU69hLkR5kllgxx9xvE7FgIeB/BkfZqqJd9/2tvWQX7TOMeRzZvQq+/NiMIi1P5e
l+Wl8QIpgP0F41wp5KZXQA/78VV/ss9YhrYrn94qjPQlWceAQa9tomyPOQH736P4
uXINq5wzmfuONj0LJj/ZX8AYFeEHULaPrFeajg4ky5EvrJ/C8YwTHkzdeWP9YDcn
P6Z0BkaBXzQu4KxSZZERtA0G7Psv0AOyFQKDOP1VJXVIt6mVJB+Plop6IzVDJnzt
NogjZALA6OsR9KM1npWvL3/7AvPrrHk3XA/91/nDTKzMKrLtQmYF/9ziJQRhej5s
e9ogL5eCO+AwZPBQI+5n5BQpICHgF9UqGbC7RBmPVcOs4wKlS0/Wh9ciA3ZgdKNU
dIQGYuOcPDmHoxvTkEO20qtvEL8sIuelGpL/ZR+K8cWtgHafhx5E3WNBATIYUWKC
uFoDlPFEt4Lf77OjpN2Ho/Ej8bRAhH9cRM5pEqFg5DSC3ArxRfkrgVmlbFf/nPST
sdEkns/x0LqzhtvR+Atkre0MXxe5XzPvdjiZyFOVBo86I/dj61wK917u3iRgR0id
TGYzbqoTs9Oh6wxmPEXjOjfOS5bCE959caDHPdNw25tO8qhlo6NJNDRICRtIsBL/
liM09sKDq1N5Owo5WHurEUTfgDalsXFNqRpl6X9vBGEnssmtbSpBwH/hxxArs/j/
IULkC9tlMT5DsAEoIkG1AalyhYyHIqrQvCHycKgAnDKrkEXF89w2ECMBFp5ErXKe
nBH3wk/0Oh9PXbBO4Lo4eTychfxQLky7ptkN60IkLToGMd5OviZlrHL2QTznpx+Q
5Pf3NnlKZfAbQvT+03AP/xVi5INIoyKcpn0tjRo8ORd6JvF/MlUQUk1kuAsKSNHS
AS7kNfWiY/5RBLXZkleR+OEibFnZM48nNQKqKWI+2rorbhMpFy+xrBgUd0Y7aLSy
KxonY6JrpN+CvpqnvNcbFU957PSATeZKGbDPfoPWvMWiiwNNkrexCIPLyfLMK2U4
pYshYkowJn4fNEVEcVTrEcP20uRUQcJa2b1o2bBsil/VWhD4FB+RDgKL5prwM4eU
/JE7GLEPVTFAUsG62Y7nilfItPdix6nPXLmIR12P+L67ME4O6lB4WBxcE3/lTWcA
SuAVpev1ltDs+etSmvX7Pe4o5UYVwlCrN5tGtmUSPf1Lontpj8riNrnQYZ6YAkKE
H3Ku4i7HReLHW+8rncj33k+wCjbGH+q4JV0DaEvxwVXuvW0qPEkrtrAm3h+pTbGU
6w8a8QzxEg/OV0OGl6VUzA7gi+pIlByx9QWDZGC6cYyqdzI20amxOapnwc2N1SwK
gQgMFZFRhnMXd2ukW2XVR8Blt4neQ96mbQxD9oZqc4J30Dk3vMcj+5OVH6U20GQi
7yn5v3cmWOhR7oNKV1cD2+f/pF4Kt4ALjISvjGQ78ZCxCai0nps2F0IHb4xEJ6FV
smM4iqH5AyspaNZDtJ5RTB8b3hsOkjg/bpNuF3YquWB4LBCn9LMw9Y/lXprFsFXn
QqNfcdc+Mhsec1UhhDYWpQo5cf6bvBB3Vn9TgKn5yDj/mpSF6QJOSnP6KZDWhb8z
CxRCg+YPELTBxbxSV+eJoymY0cWHvBQ8kmmKzXKXjRcwd/pUUswRuc/80LHrLDNa
lW905q4mQZ08z/GGblBMiWCL9c/gfN3u8jKyeyMUgDaIn9MOXD9s7wTC5NvFsKP1
dtm4/xAZOll61Ik9LxY1nlDjPnKPb/lVkz16tYIy1H5A+hS83fjN5MeoA73vGzJ3
6ZF7VXGGsG8BEtZaTQTifQVd+BOthjxj15CpV4XMydWWC8anKvlOvlrZTgvEfRNS
JpNV4JxajQiAYPmtCMlBFGqmr0A+1ZdfsQrsiKWj75cPjCWeVI+FhUEqy34IzdFJ
c8xiyCB4D2N71Mnfw8SpczYYvWD0jXkcGkAJZdLqjhj73sLd1iYVyVoTlRYKdf6A
Lj2bZxcyPSZNcltgAbyBntVvLqMo8708CUb7Zmo6A0YtdEoSx0hH52jutETrxP6k
ENTYeTNzyPQpQva3VjKHYkIbC/LKiD5yBvcyPOIxjp+w6tHS3cce9QqwYNN7rUU+
XnpCMD+sq19zbhCsT0JzwomJqEGCPz7XbC32utfhQgczKjuDUbllRTTvMuVntfG/
xnI89n9p/Kywj0Gz9BVzfRkVryBL6LcZpCFGC+AWzODl0/oJalu0CnDI5/5D3BxL
xGcq3ohhqrgE7kYZX5R6l3woJrncyoYSXo0uvTldJpsf2D+grwnitswIVy1Yc08S
OYSghy4mfUjJ0hEQ+ahNaxZuu5OKgo580cAYA42pnM7CK1kJUIFXOgVlVTz4s702
eQfcl92GpTQYnagZloCCpSwZ6x4f/h2R9lh/sn18vkmuUmnVYcFkvFMF5hqfGT+E
iJUu3BnqNLwt8MSQR6cHqLAgmdhahfCr99H3t1Pmo4la+nEEruZct7o2d1YZeuoY
bcghzO1d7BAuwi1HHLZp3lHPiThOxN67jHUPkdjBoKYSyyzgZhUPdSMjQeYOBrHx
BUHbZjMbGN5R/UDFiVeMbfTvNCHewMEHKOT8stgh6704yM0dWE8jbS5bNAlxjSdZ
TJ9HvOUq4hPE25zy8+hFlkej1cGJf6rRrkhPgw0bjmWYJCx/BCpEn+guvksZ6baD
Jn9rgwLuVnJb7T12KlEqgAAGQ/4+cBSqsZwrXnAaLwqz96T4j1zbWk337b0Ougov
VnhTsIiZPFofacULk5TPbd5zAu2Qkcn8rEafgNKxy5P2HiwzZbVxUNHQrXL8mXdF
p4UxsDATrmBXqYwKfyK2XDKanVYm2BTTNTmn2BITdF8FHv3H2Hc7Tu23FQUfmOFI
YU2r7P+uN+ZVuJKGYsoYha9kHBVaLPgIk9rqX54ku0WQW56hHIpQvbwDglG8NHa+
YYGt7C3FhNqjLY3AAmKHw/9hXP9X0cmL4BMlnGJ0dMK2XDgCcfnKkWPohwB2qG5v
rd2oylnbgV5QlEXOWUM8j0R8ByYQgjVaZFJC6oKdgIPeLUROgQcDfZL7mFqHGesT
eOkmx5C+PIEM5l/2WojwXgfF88RhxGAK586m0+cKQ+YWjqw0caFQDaxuC7HTLoT/
uKudNrd8LleoEKkEns5a9vQywcx2JjFKzGUTCMhW9WCCdlYfT67PoKwLUutbRJQi
uymTY8Sy21+3qZoQhWqGA17DmHV/6vCwP5XGMGMstUj0prUBjZ4b0rt7Y4foUDyc
RAHe6WZ82JeR6Pg9VaSV6gRZ1+gDS/Eq6zQNCUlCqJX8uaYOO+tLDkdncaBn63Ld
q4FTSj4KX19uGc3e5QvGAwBplCKjaI9oD5QioK9JOsZyks7l/6mELuBmi7AHsM8G
xNamGGKWpVcxTUTqQ36HNUPNHbzz05HFVm1AxGHzQiW3UMTejpXptxA0U9to9hvK
RknopKlgidLNidrZ6VhnJxqcsGzqgivampamnBqZxLC0bur5LR1HSS51dbMcGmr8
HGQqCuBTsYbaT+bcwo7IVk3pOipZULcmu3ZpgcvYIUOjHnOaG21lSfNf4QLTp0Bw
BrmprpBraN3JElKVAEMRz7wLWQ2E2kXqIoU1TndSwvIW9PrxBbX683OsfADQEq2E
9tGLI/rGis9lm7urMsyozuHFCghTN1m+HM8Dd3h+lTxgs+KO/Y3yD76oc0b3mkIC
Xz01UMVNA98Ht+Yvq/GrM/86esT1+m9o3XkQX1Wta7/ouP2hSsp7gVYfyfV+L6Ap
J/yTyy2A6hAd20zSgi6QYueukM95G1XfNlgCQ2GvQV73UXW7lEe+y+QVbXQzxwaf
gjvxnGf8yKq3LlJbwAzOzalAMknk7c0+IibgAhoRZjBBW3dzZkAxzOBxAEGWr3pY
K8v+9oeGQon0U787qsvHIXmEF5V+oC5wFBNYr3oQZRyhgEh4+eOI2RPNWgEXfuX5
aWYgynvNG2oBvQD/5+1QM4/S6EMghOkpxmjDhdvjcum9MPft3l3raQbqoJ16pWNO
M2X4hX18+i5ODFOPtL0lx7rjm5+yogc4cu6Ah/gjAFpzhWope+AgHWj2BYOzI3cS
h/ry9ypFpjXPelRZRx5vqS2ZKcveXf7C2MYWGKcdp6maxXjqjnGUTxZBN0qMoa+B
7yz0i55nJHWKZQ2Yh5347+lqPlu36L5h4qTYLnRJSqbxSqrMr8+F53Qw9wPb/mqp
ZijPXEnepIek3SC+wCMvB8P4ytxunfmYM/npzsQp/4g2XtBWV+IYRzK9pYSkW4le
iCzS9A7yfBgm45sp0nicAMNQcWDASblLLgXopU9Q8QWHMgKnZF396drn/HhekISQ
uWZLm+DLJUQGyeZJDHzWdSwR2sV9ltfAGb4mLPFPLWRafcEVClrmlsxbXUus8zgd
9WIa3LEEmRFuV3kTM/QP6TbUCL7b5CYeszsceets7II/uXQNBMb3+OD9evm2TGip
xg3Y8DlZJ+DXWDTBYk/ELsSwHUdMbej0N08UyreY0VXA71FidM62Z6xGqYKmzCms
UbJ0xmA5C0q/d0ZBcG/qAsx0DJ50rZRIrwiIhBx3E/yd2b8fCz2u5e7tZdWTtj+l
cC1fkpLw9+GPPcz7YBydBCGZAo+xJlb/LVVNk+y+Tyi5NPaj86fIh9Oxwt4tx9Nj
N5XZq1V1LTzqBQ1GQSmfMryV7yH9Tbgq2wy9K+F0F+zKYCsCCAb9XNjS61SZU7pi
4tzgRhR2BV7QfALtICKqFVvrSvHek4qjgCdHzUTMB3aTT0zUa7bhq6DG1h2B0b5m
1Tni8lVQfnD2YhW8JKcPds2hhFJ0lByq6cnDW4ojKJXw5lcwbORCPUB7zCyPbnsx
YoWw7eyzjdK3PRc6z7YmFNqt05t/MeIZFJj6kBZInpQgIJBi4cZOMe4TbXHtP7CC
E+euq2TdCpTFEVdb0cjdmDd2NQmIvPEqUkdgNGFIWF7icV/+6Ny7zRvnJVCesEC3
quO5uHw3HNEMlk2bTMprKzIFm1Cvv2tIBWK0N04u1KHGJ6ZqPjPuplLTKeTgKejd
F0LWIXfFRr7xd7iB0w/UUKsEyva+kSQEaUIdxwzGWGOIvyepwCJLlLQtftlgIjnX
MeHCY1amXPnCOOMmhwFBxZcqKvbSCMf9AbSWjJUbYbPy1+iuHtzGrlp6r8EvWOEb
AJUOJTI/IkKmggvht6ej164i7GYUCV93ON3RBzy3IpTjhHCfNbY7ILmj5AYPKqQg
IJ+hgFVWcpukoIZMztux43d/duf+4SOvPZBl7fTVbwt6PI/RDNW6aZzUpkMU2a5L
5YxDgmHka5xEen/MYPErq4z05zkss8oFc1192Y1lxE5vhWjIzsSZh1cvP0e25Zzr
n1a+UJ+Juz93U9moX2o/aoy4FmQcG+Bwbl1H1wIulS6+K/auDWkoi7guu7WtjZwn
EKSctOG/iCJbu5gjVcn3JHXr492+fxdMmmsINMjPoK7ZMDa4RGtI1NaS9JhUXRXj
HRyDEfxE8tjQa401wCDme2+lEgFAzaKKCXVQJ7IqS2tzrHD1tIujr7J7H20Ulv0/
fOq87stcgmfJDknFFc9HogqJM9rHElvn7ctp539gemrGTNLtN+UffDHi5jcWIV7c
v4+EJV06rPQbnaBi22+DtG1I02ENv+it+LVYRRIUeTO18TE2lJWJKrEanZjFYEd7
R0x8GT6zAkF8Eirznay8z70lapLkfTi9+6ZopcqOnaLTJETo5HSNs9YeL6Q7mPC3
97lkg3sw18hOVY2gqbgg40hlke9YLOdEKaj+w8SzSB6j1gRffgxPJqOGRyIdlqn6
9SgBhJ24gxu0ay+05sqmj9IfNLjmct8lIrxvOd58A1TKbisIZknOqW4mxIUTwhYR
KRg1FyxH2yOrOMqfjHcY4RIZy9ckCVa7Dj8lz4Ytg/inC3Ax4djuSMqAC4IVUcos
/oXW7lrOY8egfD3kOGCWhSlcJm5kJxO1fxdID1Bj32BCK8cj95YD/S3j62OMDQev
5p76eRvGWo83VNHVwdPk6c/wdXwUCeKQjHaAQIqmDAfzeIAg13RN85eYLieXFOg9
QmN4brYZ5ZslEhoFvHQidhOa29JLhA5ym3ILfJQR8FwTzndLy8b0XzY9BewqXpS4
34TgJ1IATDpx5b1DiXcGXNX+sTKNukG/uEIFar+PoSYNjajxt7J5vOVBbNU8aDj7
UbmV+h+0XNA4henILBoJDU2hJNoVYZkhZ4XqPiiBwCTbF885HbVM3AR0BynqzRPK
p24iSp6W7wL3ukLv2sVU11DlteKL42Amb8l2ExsdbXpeGQyB1aAIBVPnYmar5EJ2
dtqBzSD/BuMf3hF0HEmw+k4wK1Vw2aggg2V7XlihpMfejxB9SD5OhLCbki4Qp+dK
ozABbZdePZ8EM6Y8AqdksoD8MPxu+eTEHwKH6GCblQdXhZpqPiIrZsxwGpB6UCXe
t2yg5sSgRbMtRqD+Oi8zVtWUec6QNIVz3EZ24m1ACPJEbd3ubGJKZXu3S3ysPeuv
Ac2KpNJtY/EwPKuFus8yHHm/n54r0KkGrU3Zs0JrhhFRdTBUEG7DKAHGgZim7Dpf
AvjQSTtBOoKb5pkB7kVDns5KUIewXRFhSn8i5QyqzBwmn2/UyUx9q2KbonthyFuS
poVjClALMy9tXpYnrJcSCKv0Fn+NorGsObNdL1Q5VopOPZiY2y5xLyP6JDpWZbZC
14a/D2sQRL64fjc8yHVcpK6v9d5amtDsm7Dd2FtS35vkicQAsNof0Ge+/YB7CqAg
h8CcsB2p+Efb1BZaH9JedY8wMFkTnyj1lyqzU+D6yunihGveHtzWnrbcto2+Q0qD
zRo1wAe9bwCaKEYmhSjLjJs7bFY+A8iOt6pa8iwj6KpEOFenVWkYAQVt1DR76EOw
6sOq8dCI81RbvNTnI/bhGG4FB7VoprNYT/JleB+vRxA1KrfqA8bpk2G28CoLG9TA
D4KYz7Yy+1m5jWMGoOEPJw65RUxGrK8mDz1fb2NkOGDQxJBaASbfgpVkMIbS+Uif
z9XApIu+mBtIYcU9DU/2bibaotbQPIPwTyJUhPqErDizpgTY0G1+X0owuLuiI5Ty
Hz2qUQ7Jy9wzYVAsKI/1VckdajhHCmsXn3/eJ7lF2/kJHFR7pxtjF/BPfC4OB8Kr
+YDPd87j6JQraLPLzyJ1n/Aj2Z8QOeSP9Ik8IVXmA08RiInF6E7hNcy17Nbqft2w
MSPqKPKTAfem5eyrAZX+ew2X1kD8SBAFH46sfhQjQmn7/SZtrVDE9Ft+rlVwxXpJ
J+aozaS6pfmVcAiRzmE4slXTaHHqLUj9/p/6MUG6Ozs4ub4YfEpz96duBQK/0oLF
eKyjy5Vu0mZa5m58fxxF9V2zUcjja3z1FQ/KysCHuBx3KsTGMG2WopaT6r/fd/wF
PivmkjvNpQbYmU9Uwe5kgoME3GHEzVUSsr6SMxg1xVc+TkA9POn6YdpnrAZCtkGV
ZNkcHLYZLI7Mvk/O2sjCR3QnAEFqkvBUfpJr5idPdHKpJCzMfPdYuHNmFBNRcZXm
cVaxospUybsJRT6+tktont8/xPOsnxYB4rAI8rOa5/m6mLJ7KPoAtJ6qfPCsjloo
D/Sgve9ODyFgTkZaTbfH4Uk79NV1IyWP44LSPgpzoq52HJYCyYAXyugC5U6JN7Xw
LXAbKifZolwI4OY+ykv5uzYFFAi4VK2nLAUuK3ZG3f+Uh73ThraavXLEIV6EccyN
JlEJmR9jAw6dVkRzYQImPneU/Lw4NAXi9woH1A760tD565eTy9cZtDWNf3XvSN8z
ol1sciCccN1OfcMBSqbWNTW/wYTgsbSqjNngtndyX2PrLpvwBfxH5YRlMdv54pHC
VtSmJ1+kMLVx1eOvtcSzkzOacLA9aRvC12JGeraoZwPwp/T9LubU314s5TaNCnUk
Fe2a9rnB8Y1V07HuLRtHEdCueGG+JjTd6yRLWtOxlDssUAObg0tKHDD5Kjuo7yUi
Hn4XE4PU6VrKRBvuT9F6tKXFmwqtAxcuie4csUQyh8U0WsLyApVCZqjQb7OqsrvZ
7GEGvj1EncxZ1fDm3VK9WPEIMCe5AFoQCOcfAJA4w+IAdEvHi/Mzthdx5lF3HZcg
QHEKszNTifZWYddkQNM8RKQ6SjGAl8+upCLbUlOLNzfDvkV0PbggF6eHx6z/vAMj
g9z5pmT27WoTTWV4dLaaJ4KUWc6HQFiEcgjn2CBuytzfSrH4wrdNXFnJeW2h8PAZ
HtCka4J9MpUogsOXYvt4DYT9sFF7l7ihLLvbt6grHT4cPSmjQkowJY4uqmQ7/MHQ
1Lq5m3DEHWkqpocBm2Xbf2Ko52RmIxIgCo/tIF/xM78s2BqN8DuuRr0g0qXitNx5
NN4SpxARIf7xhaMJZw4EibKkFdeSFftGY/3l1NtXtgpk7fJD+zYUkrPrrLx0JVov
LCvLt574F9MBDsyvt9FqCEoKVLYHCYNi6S9sLQilP2Od+/428CrigNt5ViXAJiDh
GMoJDxoFvuey9EP4zQnp9DsG3deZzhExHfpynAUqVkovyazL61R4yuzrqeYXYKrv
m1B3DjpZe1khfT5fk3hWnISQSnNmXykoq2CeiFytNdvNJ2FTvw8XswURkTH+E//K
yZ803hTO6vqjGpgZDDWrwTzE+rb005oqXpPcHGZsR3gBE+a80ciHxOJMkdf1ar1B
0l1botIVicvRPVB9AufRfflq65TsV/uvvDjc9hCg6zLzwCAFA8jTQg85jpuCFA8E
ygiTPNIUWlYF3sP/qS2wd70ohsZm0SZ3Z3WMkBp1c3n8bXfBBhe32+vK/GwnVEXW
E2BoGs8oCaWKnjtebucQ7EwMjAYRMZPZ45CIbdKPU+bOtQf6WhWuPTFF+eYiws1P
LjP89/WXn0oOaddS6Y7Q2ScV3/vCTj+kjwHeINSAAt58G8AbDnOeUoH6nPLxuMw+
nrskdJiq5hD3WWaP4ZmgQo9InEzSzIMgzkznH9QfaZ2QoMstr9irTWfqlfWIp7lz
vfyCsgs5e66fUfpDo72TgawpW7c5N7bLIMaGTzQcQbIpuqjp+/CXucjTrEdOvWOV
HwnxBV/CSWow3Wx0MT+k+836fRvBgCnq/X4mPpyOFiJhiDSaZxFsl01KPddtIl40
L3OYjrufzJo4avccbEjJYAv5JsTgI3vLK7TNKuS1zmGRSJDTw8fTWSpWN3r2p9iy
cwB4kfPc0VbD3gWPH6xHXjZUas96tHQgh9CxTmx1sSl6B0txZ3PaPLi5P3JkTGux
Wj+qjvYefAA6pN1aXDk1okq7zIdOAMi/P4dXli2f0Rut9u/bMoHn38dVKVu+ezIY
jvUsthF8qWJx2DkRoO01eGX/hz6RSDbowzKrJ/xy1KHShdHejygxAXplnOToPvsM
GAPaobMTN5H7yur02yAt9W70ZgrUgAqeNNeRUImPonKYOzJrQC4pulY/a+jSugub
OLdWUO+rt6wp/LOCP9Tt0rTUCAPl9qqh13MCOxXZPfmK9R+2pZAotlGxUw3/DuPG
xiv3dWHI0PzzQmLwA8Ksaj+KwGzBQ6RM2G7RVphINmBjD4aoGP506a/K+j0ji2/e
zsD8eoAfaqokKI/VscXvCRUdlkHiK+ACY4XOaIcuhdmjMP4mRfopFU09DQI5JZpI
DTHaGPoHHCdbA7qYRsmGuE5dO/NDFVtubUyrV9mPu8PSezL3ssESAl9vl0sZdNF3
oOuR1Z0Y7UviSPEaoXJdgJlphIKUhEFMTwz/yEE8GHR1naipkpduOhMob+pxjIaa
OpvyzXScmlJqM/JMA+UXf/ftHeaLmCOAMmlwYNthZacBbN9X/22c9gExZP/jiium
y4E16BrxFyMV/HETKlPka4WhT1oTOZQtzK0f2EVyz2qZLArORJfB0GGZXx0ztark
z77g2gNKarAgpULWjxvodqDzhJC2S7gxRm5APx7INngHQ047D9hsJThJ08fQWgNL
LuMXeYgCH46i0skTexreewKTsYKT2C1x2U+pR5P/X2rCDmagLr+4CvQN2sgXBhox
XrwbdWlyj/sPub1WmAX66ZWxX60eMSeN94maQAU6kcZekxYDPXRaApAktR1blrif
1qJ0zgGg6RVr3Y8YBnDghN0XQGGDDgKoQ3GzrI1CZkWO9FfsejWaDHcsAQTF+crB
65M+mf0tLnJ4D9GM/sjI2kjdRwGE5J37GVwemizcg6NZLVfSDoB4O8asDxA96ma3
fsB9+OUk3XKqKbGnsH/EG1kIQUE0l6v5CAk4EbuwhmhRILOs4mC2SmZ6EMzor6RC
y23bISUSaXXmAl7V9U5r2n5eJuactpnwkVaJtfrFnG/qNrq8X8h8kv2RGYdRJwig
jx0LncJj4IXFWUx3QVKc5xGF/7ezuTzm1jomoUq4lFG/ESfkAOX20h9AxotK7uac
k7A+rHG9Imzx0bE53bjW+UBIz5JDfe6PYOeYq+CtjgIzSyfE8qk+qhib11kNqHo6
5o4adqJ/EaAAuwMkrbgYIyN8WI8SY7AyoK8YhgNL7s5WjSe4R9n4riG4+HTGF+TY
xcA0A3HCmMJNYxhByjq6vX0qg6FaAeRZJuUJNI9yhR7wKgODmSOUrg1xE4EGgpvi
/YxVrBrs1gdrRELUckDYaWjj1QyApe3JV8qVu9YivIjcOyreJOjMpYf8Jd0s7E02
Adstt+Ulr4E5l6oMVv1sU0UYIgPy21aQGAnS8fZaSJ5os4C1HfsOl3OuvGM8wrNv
taaNCiCPqnpdT/sZRw3NCi2ev5mAXIXUNgopeYlG+9PMFd8LXpcWiPZ5Hvj8xsjU
G7V9t0UMc9xzwvd1QSJ4bjyccQP0UoPUbfg75I+G0TMyVIRl/9JSMBQpJr+TJflk
tgHVdWpPA5vVZNDVrcYf+HpqaRuYwvhBnlDFD5wAzaheRddYGKS2NYqQU2cWEtcd
igpXoYKXdrn7uweajnX4nNDcTZGybGInPgNXdd1AQNKaSQJvqiw9Dbt98n2o69K2
T9jeJjhz5x2brT3uYRVlfHcIf7iCtdhJ6VXcQXQ4bM8O4ziFkJ0llZWPCkffcTBm
/O1jRc8qptzkkizheNhtFbuZm9S/cRdrMtooMHg6Loxs4P0BdvEsf2cBdnWxWM2J
DreUu7WVNVqSFcl29V2yHPaKIypmZF5izBtZ9HyollNEwq1XvW0V1Yba27LMoMzu
OSuxzY5agPi30zGYmmcj9Wbdo19HANj0XHUJcIkKhPyQpYhX0QT0rZ1pv0PHHRdn
fjs3vdPPTvoCSVGlcZrHx9WMfgcowpBjWk6q8fIZskOlYDevgFpsv3FzSW/b0SOc
pNq1a8evERn5zqGdkajdwt9sYxUtifYVDdQJeuVzzWCWWr8EnO9KQyHlUXRCtSjC
zSGvEctfO36dt6RfECOJ/wZVZ+ZpEuh9gRo5b4+pQfN4ZJfT2syeC2/Ua8BYTzHs
98k1jyqDfd9lri+AplRuhjfVf7Ue+I/gHOZp4yfCeQ6nROFzmF9lHxMdk6PdgQRG
Io8aqcvCTQnlq+QY8aTmencrkZjIaiJ+QVW1MCQR2sqfqPLb3k++Ff7OvL93ycIW
kI6wh3Ee/3APfIM9uNIThy9PBu5HFFQHAVDSRNQc2UHAntczvO22MvgH2xmIx6IK
LgurH6fuMcdU4VL1feQSXybLKw1JNJ7B5D42Eps2rfsUThlN9dyy0B5+w641RhPI
+PCA0i9Xyf/OG+M56o7FK/ulByBKd7kwOSmcAYo9WICp8e8aXp3t/qL6YtWpgCgH
U+BBNiqV7erGHvPy9ssA+Q2g7IsWUvODXk9vw/hdgmxocHWCE9tad+6AjHAX0iBg
XJhFCsu3FV4vcrplMpOj8TT2dg7f2FdiCncOXIJYCpxTtEVHkh2Ilml9an3UGbk3
Tir22Dpk1NnyP0hJ2BI9zXjnuj2fhlAPCSOHjERKe6SXw5muaJqpR7Lppnj0mcBN
4pYvNUvZWvP/bEZz08SY0V4kHA2CqK0fWnhwqQX62y/XhWZ2syfcBsVEPtHWVo7+
7uoLWhDbxYJSBa7wpLf8bKbJstQTYQ4/wShtFLGcIWvmeeM2KeOGRy8NTIFvP5Mu
mLJua2uQV8KPpxTZlcVpK/nh83Y5C7rBpyrFL81Gjt184SzzsWHUnw0PcuJRz8/h
/+RWDP8RlD97zdfDFezYLLBs+r+xiJgZ3Xc8JuWuoLsOAA4PloAop3irA/g6caFg
YZBlnmeWDQ4qBJklvgH0dgZHF0Bmw/WDe9KkLFObIM0rq9c/a3GAJsubraOSR+Lh
bB2xTikSOJ6q+Sgu3rGqZXBR3k1AXsbF6Xipjqoevn+zJC2C1d+KirlVNCocCY67
ysGg8mU6e9vf4bFTy5EEfuNwaggJFnCh/CMVbtSQKsbFZYurC30Ngs0McSUf2drE
0CuGKmBAgwkHt+skGVYjVPWikZKjyhNQFDPxdLBWLlXwTrNfbrkuBbSAzgVlGkn+
SHyYqDEGja8cWuYgU5DO+d1Yxg3CmC0VKWYxFDGMyBAsYoNP4Vb3IacciB9j7/In
n0GXZYjslAljNP2YE5LWskhxMS6rdV1NH35FQDzHWIyly/Y42Ewzsmh1tmfvvCEF
plZHcaxDSetipQsFX7+g8Lfqs5r+rM79F/E7K0ECK1VPtRBDOKusv13afDXtdvaL
57jv/+ojRNDanlbuTpC0RQ6lq7/PzTjqZ12ZAKSftTsMApITcUl48Bx5+yFSgqL/
5KC23e+GhP4vxJwBark5AJXKIAl6QejI7+87zTrslExFdxostMFdtK0EfjkGCR+y
iB+nf4KhZRM2yvSspPvc12g/KaMAf/OmokidEmPc/RRdZ5ThPnRuSXmEyg/jXmUW
lD/buo5WLS79255llWpkYn0xTbcosTyfPzE3o82BF02fa3ezCc2UgNNAroF6Rv+a
Q0KWnG1+IbBdUVG2FBmUUDdSyZBLSPga08QDPBvbIJy94ItH7w5uM12GmxOwI17v
KsBzTovvNaZqRyy+9uPVojNHtf2zPH7cA28ri5nRisnifBvnaMMTR21sL+Y5hZfa
L/iJ4WjV/qpeZej1YNpr6GtHX6gCpk0IJph/juQ3spq8p99LA1AuWX2oQKOh8o8Z
acY8Qm6qwtzlL40E06lJz4KzfiCTMH2gRGV4atIsac8xGi88wExRr+zn/zyTAuWV
eej8pnRvcr0VYatAoXAi39YdGnC1r6E/fKx/IHLL5b5PNU4zagax8HYE4MZQmZRa
JouJXnK+DAE2ThY1dfyy7ZNMTvGBMkbPOCyWXA5+joo0boiy+1bT7/yT4X/56jxS
WEnNoNci3j1kxWEz8d+Tw0pQ5n5ULmAup+wnq4xoU2g+U9BZYMBz4ut52BKLQsZY
UvNNTFBVf34Jhe4hK5tcEpZ9Coq7jTd1hUlbX+w9Rt/nb+xUCH2B9uektjvogMhL
7GSR/D+rCDn4lSsmL0hmoKb+X+ht6m2yZ3Db3fsqcWQCrbzG3s2Yjz0AB+DHJKZw
tjf17uTeZuvXNky2Ypv3p5u4jBcjE8NK4YbbMOX6Kj6TWtSAdvnnCVu+D9bjM1N1
4fUUaP/BmBzoBxytb2KosdQZVS7zDRcQIyyxPzLiA5eyJc6oCHzCXJGWZazucgMR
jydHO9kCFgbTvUttfbTJeDQGZpspX2ZnrSXSjy2jGp28hADxqKcu9xFgQLwamZGw
c3RNJAlsQ5Rt32acJUfFQCXtMdYAdWjFlAd4nfBhFE0REVdHSSr17i+N7QcdYrKl
wyYY6iT62lmZeRC/AM0Sdmi9wxTLWevUhHURAvtAQX9nuGoN46RxH//Ok9TvT3oW
bQFagfVg94d0Ej9gHXI/H9uKWKC9bFPSGp/gnX8TEKhbchzV5wfiaUvXF1u5kJDR
/nTS0ZU7a2gtqHWFtJskw9EkjOP1HUBmXyvgh4kNhYeWZFC/haphCZa2pHHVYBbJ
H5NBLTjKCqemZcuSttBqY+CmZBv4SYbANWafa1yadJ+kFl4pQ0h0npsZeLm4oANh
16hXqx8BLuElOu/6f51tkJT6/9Dfzys0mPCfegVTRnFINq7lnMnQsnmJ7dhy6Dq9
v0aYztwkxwWdLCqUJjW5a9k41lD032ROM2Vn72fVXStV8SmXwHxqAdbnVHvZ8mHC
eL2LdmRIns938rzgbIaqv15gtNHgbXy2FSsb6wUjEC1sDRvBX2ILKitjVP+gRqBu
p5v4QSo9xdO0tUrBjhV0qQZD9tvRhgvKp/Acu2Rd++H4V9ZTG40UCmilUm4g+Pgo
vRNl6CMQ89XlQOSukj1jbMYrozOGfV4qIKzHFYz/D4ocglk+MAjWRjfXOpKWM2p1
d25qKY44HPfqT/lom7QJ48GRoc9UbYZiQQMNz9IWBVqXN7XW3qVNJrslDU+jgzHi
sRrggZjO3Gk+Y3WcTdI44KZVkltxE3tjKepBA0NTJczBrKQWjkFSSsGOACSN37E+
qyQK0WXK9BwAam5ZcazEyxddtVsYU9bcpuGDH+W7J4OIfO+dvMTdBTTEeTUz7aOA
FBqMZq3b+GtIqrs+1UCUswx0dq0mvutLNvmEnp+MBUWsdcn/ZhFtXJiQKGXud6v7
UCiFZIH14PHOBaKTJ3zVjOnL2fBewHG7k79hGOYQrsJ0nrcCkjZts3ZAHcm40IE6
YQiLB+e+wIR4xwlXFE7fTh8QdGzvM2N9WtxLtfHEcfUkd5hYtic+yJcB7LLk8FcR
7S141H69VN/pBR+BVhsWUwHwQftlWmJfOCn3qBERNy3D8QRau1lsFN2JrgsSC/g7
/wLBNaVdtyE0VQuBJvwHwn/gySshS2IEKKvTZMKlYcynLmsP1aA7Gu3sb4+2W2yZ
fL2+ZURRW/sxa/FbreC0OIpmdaqH6D/umNmHpFEj8jB8DeU6cv7W1cC/MqFYpv0O
Oe3d0lpKEM+y/yUBksYVxsrwBRycCHgG1D/KjcffsUkFxs4Xuel1BkmpyY3mBM1Y
U6mSBbNW0Sj/3KYZMAgpjsdRcTtDfV3rHUdtqBWli625Iq3U5jOgH5HA5tbm9Kx/
1w79P8XpZsAQBmvhi19NMLbuyiGNuyXuRG70uYz1klELliZrjUtc9BqjLbR3cltR
hm+8mU3Pcrrem57AfzyGVC6FkwVGhevX1ZxtfsDvNzBsYfTf7bh0EtuafOUSfr6m
7cAVjA4Qzq8/R9WW0zetraVqaNgKsrxCZH9kk/d3mPIkBvgTKAc8K67VkMhwi3t2
XdCFn1+j78/righnnzQG5jjLZE5eH23wMBVeq/y+VdMlmkgOwLHhfX7HqUbD4H81
u4rIxl8cYirWB2ox28JdG2ScywIHITVKHuxlxqucfdXxAsMKkTEa0UQiKLIjktuT
V13oqD4loYkruoDlk1ugnY6F5hwcap4kGLOxdLprSYViBmWnGnCSOrlf70SMF09C
GoS3sccIrhM4/ETxzFJhPd/5r9AEphS0MeGF17NO0OMN7XJP+9eVJ+byTBBsvDo1
O2NEJZfkJvBAKKZ31P6qAMCrFjtr3oeQ8j94SqfRozO0H8yWoWbXMCZ+YaxqWRHM
QI449dn3FEjXKAko0XNOyM9CqiBxk+vUlFUefeZyYDnnFNEzdEmEeKDVVx3AKlef
SSSdbdtNiVDI3ZHlDhqIU8vJiId0dN2XZDVzHp8j2ZSkxvTIDhcUEZAiYXq35sh4
jIKHJeQRz1+8iCeHbjRzySbaYrKUliL0HnBefXKQ392EupcQwOJIwvTWAP6gmDlV
PKi8m7D3ZD2f4AkwuFlLbbexJTTEK15CeuRWbjn8qgu5xVlE9W3D6Ve0Lk5d0ONH
T9zc/smlyDRhUmX5fapU0rwhDBdxMJxZxl8AzNGQwrWdBEv65MYv8OERZyttI7JS
mc+6qdWWyWi6WwEhgLYlXcDG+6edsUyjHg2H3Qw5t7q5cFrCw1tvAK8QhTmoIFPc
xsX6RphPCJdRrstscx7FXjIA01vlkpoWoLrLdt3g9X82hd3gKqkTc/jEJyACfKbL
n+U7JQoyWZ7c54zzE1njfP8RYKea3va7Iti8usUzAc+6irskKHk55yjgyxy7nhHV
MGptJ7ZDrqdCBWBwmAXXYxIDnsAutzNgbt2dyaTg+CaOd3IYl0EO0BoEdE/yDOwQ
Cht70YV3AsVKrm7ZS+E3FPghcRafZNmcXreQb3KxaRscSIxGTGrseYmoeb/1iryy
6y8QEdjPivZ0uRsxWbccv/OY9ddv73Gvq+b8aE9R7Y8iPd6AKu74R8mGpCdx1e6S
QB9o6k+Oq7aAH87nt8kpVeOh+nMcFhMlFo1BrusynbnDs7LlAfryuBMNU6b7XAnE
RRiFmyMKDLN4iBlUW9FAL5WbnpGcws3E5OLcFo6aNDOOdsIuGoiNULUJSxZjq3Cr
3ctZhxquRVjHWmn9aIsT+VRC6vcwwoGUIYdIAtXSLtpauMaQxr5JwnIFN8uHKJdR
MfO/JibXTamiFDHXMnraSeCyRmwSTM+w3RhTtYKFs795X84FgfTBGf7VgPLLza93
Z3s68uxaGftt8wXIYNaha7BcUTpmHrCjf4DBHMIO6ORYvp0MIcTjtIoMwCVYqWaR
crkfpfyVF/ws3HYz0Q2L0LLb5Rl7rT3o+lwGx1ZCp+z/1NoMlXrDHoNdsykQ8n58
IO7TAYrOUFni5l7F1mPEuEo7tiw2rRZjrgBT1FW1l/K1GX8dppUidrIyS6xYVNOt
8fmqQx9a6rDZtjq4Qa0o0bRLPJSvV3utBg/MQgnsKI0Y7FFjtkqWVg0//gyu76GX
Oy1yM8mywiLrppG3JoZExIbJxnmcHkvp+jzeH9AvcpGbylhE0lgFMksoKDfACOir
ZvloPmcFQVH5d6SoP6FuH3/8cV2eb8z799didgHfLsWQCBsbPzgiNo7oC/+YTP9n
XjoE+x+90kiyZSzRBew+eRzPbczcIjwqEzGU9aJMAFQhO+3DTHpknkzHgvXCp/wJ
/eWCVS7DiGOzkk5wxuxZhEuFYawbEbiJSiyLOUPIcwPBC9k5c4Qhq00CuVVdVU+5
XIWcGsQOzAzT2wQP93Oikt8SoH4n+aboV8/i9BtEj2ZiL1qiSinc7zXjwZGpLZdA
OneXBw5L9t+5Jelbc7la0gXUjMeE3r3O9nRWYrP4zWK9Jcnl9LSipcKUorLb9Whi
0ooPUwyux1NUg03jyKXcgi2SA15KU5IL2jk/vqjoVzJPzDaxvwSyjKjrgrenz2wn
IcfqpUNUi1Lf82/QTh7Pjg8Xb2Xexm7YW6zgdigIOPkhyUEC2QXDrSmaHq9oHhAM
wpNnqACFipVJqdiDviacUE7H7pWNstFRO6YHzfRww4mRLgAW3thmYAJ9RevBd5cB
B4TQrTSxAl0166LWT/iaosmlW7fsyrPq1F+l+8FkSSmugG9Y6FWLKG5b5eavhKVH
pMkicm14JHM9+CbEK6mFjQxFkDbm2HI7l3ExBDhMVcx1ls6Wi+1aznH3qN2JkC81
xH289G0xMAvf7tQzJwIR08SeT54sW95eqoYR+WWLJFDovwJhCNn1aNNIsg3qZlul
Pu9sbZ68pvgSukL7/hyHd9++1fOiS4uoPQqGbi1ONAv2qfMph9zTyLO/VWiFu6pJ
URe2gPk/dHuf07ISPlaKmY+Cyx+B3KLde9BmRe2UCT6vM5luFsWdvyvxNPeyD1CV
kSdAyPEUx4TY4bboeRLhbsF2iGSAkVQttcEG0tCyJVlS14orext/HJDYa/6ms7dl
uwkFjdI7EfkaM9oE8gKmJPfJqglGBrvPpsh7G71cbEo5zgkqs9GbkYH/p6l9Ra0M
xGY2yvble/B2ISgUJczsydokFzPR5SPQR4LoTGiqpvkUZtaH/yv+eY7L0fh4/vKk
lSbxnX+HGzv+rOJGrdK6ukEMSOEx1IzX4mbtL2Sc9yZpdpKD2rJM4dwHbIrmYo6x
6C6tYylNJZVEPHuI35p64aDVRjq9tfprV6xZlfPXNT2fxRByZ9F6cEwjv5FtJp5U
NQCIecsbAB+FPqdWYMb0UqOFGnvbWkEOlUNklnQdDmjr1YhWqpsy1BDZaas9NLF2
a/5i539ON0EKxZela7IuA8yyICbkAUvliLoBF8Na4OduiyR0xgFpB7ZFxdswDmNV
oFBmjMvHoUuMMOA/OSM+Uk7/82OloHtBp7TG70srzPAecu1LRhLIdubqutkWDEDL
uYCrKWCvs9t9XLWrw+KRQClZyUuqQ01VbfvJtRdqcwjJpARI6pNzw+eSiN/J8myV
r05lcEs9idgXUGaBkbYQClh7N4Va9OdT8Z3DloofkOggcUuebswj0W9U3ZOCasuX
Ektiq9NIYdpO37XYy9v165Muw4erw1UuWsFR3xPuEwTGkPjoVaqR1g8iIlr3jhdU
/I/HoIn0llIWy223vV2+3r6Sa5Uhp8GB9wyawXyyHz4752VKn3mjyyXZ+ETjt7dy
nmYgepQra4gcdOsubgofv0FOKSHacn9dLIJbotjwZOkJRCxASgk8hNLhsBTAWNDl
WlLcn8QFCu/6JZXJHG6p/z54RDz9QSBAWTrJOxKYV1Ro/wA/I9amljoeM6+4kjIm
hOvyy6TIrZmfWwhOvtYmTipnEICJZyimNIDOFbYWdNaTkjoUn4zNBh5T+NLWfIA8
CQ7OqkHey+oWaJrqSRM1ScJjCdgWjwyBqPafhR+kY6RW4unx8BMJooSwKXhyV9DK
FGp5jwzz+CIQbrlXfOBisDnTLw8eAPtRB7N3pqzr4cxZ5S9JFN2/2ywsMvrCfBMd
j9YhC8O9xdZvxo2jOsHSS1/5Uct/+vC7y7TzGRJYS95hwbqaebq5ayrlze9bwKjD
29D0+NyCI1YX+Fed+6OKkp7HweLVYPmkM91zeWMkE+tZr/8ZxBvcusdDL0aXCgNr
TRJN5vID3sBGknKxC9ju90BVcppLmKeKuR4vjTGXJokt9TGII/2O/Ck0uScCesK+
K/kzMvXw5FqW1Ot8Lg/ObNMZIotcUmdNVsPvGbghLitzVUAU+wiW05UDXSXB29Ji
OqbRO/gxp7gq1FOhfM4rxUPVRloiMXAmJU6Fot/bEUHi9MPJuwEvffkJ1h+i/yG5
pqkI0TVXwIn0NBgUx0eKSd4YrCJigknJWg6utZ+3ZIrWOe2w2Dhkn9elLxveJEii
UviRE68wIEixl6PjDYOkLXK5tVQ3nYzy39WE4xEKCnMSzVSmSHtgcAb/gI7urw4P
sbiUkoOzBnG8902w4WtqeWCut3YjaGDIFYEmOb7/RUpYsahxS4gIRd2OgehEGUlS
52oK3K8ntP37iZd3/NNqG+Rz1JjRM+IdQ9J9o3711WNGGAhxJLfjZwZQRRj3vwke
IIpGazWBs50uowGLr62KAOMvauqfkWHsU+qrTcztd1/3hIs0fPLE/UpTDW8yFbD6
QCeBVxsq8Gbz1drbZWIViA6eU6DqQ6F6MZhqqhafz66dR5g8N2B9S98mbOshmt2r
bFn6w3/vu+zzH56673D841sWYDTlA7fjLWXJCZ9AhV2/rRWaw+icqtlaUt/EE/XQ
3WlSFmniIin/QFxNdYvWgWvfsFzNH9nap5/hq+bgKMk/O+NLUtMikdev+WkhVYC/
yE3MdJenMIUhrs47qQk6JYA3/BAbCh9Zos0VRJrV8zTvOsXNnmIHRxa+62uWQRnW
vbbRs/sdXwfv+YQwCn5PntL3P3d4Ux/DmFZCKqhMWLyxc5DaYRqR6uLx8mm+w9iF
idDkR8iSjtXt1eP5xIJ8T9P+jkqmT1pDFKV7klUCbNj91YqSdUqK0oRVDHHvb7Bw
vWN0ZI/xbzwhCd5yg6L+gDCd+KnNymAb0qUm0VI68a2pcLw3yYlYQAJqost8zzNN
YZ0o9c7bDgSMu9ydKPfqyfaXS3bUUMjZkKOkDk9rzSz/y+6TIsxo6sYCpNXBjBh9
4DR+zs8gNkGxPtG0DizwAlIQOk8idXHSt0YNYDxdJA5XvVFHO0btHnyWNMl+0rcG
DAmvHOzMTCxfAvt8jHveMpc8EtJm5RxEzmQu2BBj/0HWWDmmAWhu0ykYL4RNHNWu
Sd5tCxOGf+7lCg0TSkRGyEiT5DYYb1VvP+5YetmRnRc4y+YpcKFflqkR7cZ3SPoM
M2lsVWTlmIgLlQSvZfVEXtFd2LvIdQgE87CVkt17Prjty28wtaGygk/eGqx1esIw
TnbacUOGhq3p2Df+m/0/D/I5nS+wXpa9Y7FahkgEfoETWDvHtZzGfDd7Ch6nBjJe
+Hyh52ruBgsfmZ0z7d6p6narxM9Mdk4nuCswi6b+nHsE6eMASm/8lnzrYVlxlAV1
3y2dKTde6QGjXOfZUKQltiw5raHAbyaUKw0XO6b2doH/a/2lWUkOS/GMQFsKHvjG
BpStDbEunUUPRjP9UzTW5n/ZzHHesSoEu3RbZpr74ssL3i+ogkK0uBlddNUJBIJf
eRzuejx+AYsj4wR/C7Jks3TqCBFzB9+8CRYoQ4XDBdVk3Bzyf/I0vhCQyXbsjJwT
Ne3+trzTMb8NjsFqzZYk5jt3ko8/PxXlqY4SAUf+XGwmhV6RxHh4i47FK8ijltcQ
qD1bOgMBQCdDjvF7FrRK1B9XVCtBMFa07NCo+lRQB+jUMjC8TfNCd396drHy8coS
G7yxp72WTwl6R0Xed1o0ylHc9lnZDtUS5DgdBn5UyaMGr3dElxmsfDN0kIa9Grso
SABbKU+2l1aC58IFKVcMdrGihQllE0Ny54ttd5hQtKGVXApdbvt2ejt90cElcjJi
BvoAg4ziUhnEaTSz5IdgN9yYbe+MpUqs9xT15Bt/Wbc6MAZF/U8GOyl1joxqTPwR
ETaei92BeaDSAy8EgAeEAWLu8fA6M1okr35fisXM0AWVRBwvrnJ2/hWocqt2uhB0
aV1YLAzCVweNtmDGL+7JyVgwOipX8FEs4xvLTYIgVAnN2hIIZg508qB1C2CsvWSt
kl8YIqXjslPpo2zQo40x8TlV9LYOT2AtJos3L1PCpFAzCDFbe5UNBMc2upt4q15U
Gk5x1+0no3V3PTwDN2ZQxwlZNlDWWduHhppQKYVs0TsmKVdvPdoOveOHxqeo0nqe
IourNnGzoQgBNl8m8xFJQi572Ryj3juqJy0IkgJCDz0Y1hmyb/JLrKBD9ZC9s17w
kOu9Yb4bpqUX6/aTTNlHZrr0CqTyqLXh3AnYNkW7r/dYGHoC/OZoCa1SqyHZMphq
vhPuX2OmhgWSIYHIDvINz2u+Nf2g+xWqjNXLkaoD568zR9VKTOigRtwU4E2cYSWI
P/W1Jutc8bSCON5MUMTxEnwrzI+qwlF2fA+OdVuzmz2b3sxWqRpswrqfPVYMLV1b
nJS1FcI6MaccMSMXwPL7ScUgfpwzin1QiS3TSWqL7mlyYGisgOOjfoCrb1hUN4kx
D9lJqgR02xjVyRtCo3WQppVMCTV1vPljVstl8s5I8bWr1S+BAehuRiHn7nczRKmR
h4scXQMC85gJyS+1JcyBt4yoe8LB37/yO/7t2d5LyvuRKnE4dRHvgl5OQc/RoStS
GZgGDA+Q82b3ai8HiE6/qI1zpfUCpq1vNxO6dMYlv1sFTv3dp7Zn962byaM1Mcs0
EVkaeV76D6GbtZwq6LGLWMKXL8yUTKYAeWLGobQe6ULdPNCJcBi2M4RcjEBGx9il
7e/43XWuGQD51GXsHD08Hc6Jpk16X0lxGqmBmhSTCTG8YCfTCuIqNkZSyRbeoNhZ
L/AYnDvskL0xUiJtCjYQgdeAs90m400JuwlSQ4IYyYdPbqEkxxe1dc6gPuecv2E1
7hJzP138PSTQrAz/we5Y5s/A/73zzbvv0omwVEYreVcz0v4L4UoF2SjWESz3uSRS
BQxm7e1UZAOV2KN+PZIQs1/lG01N/Jrf2Yp4b4LIQHCnxYhAicYLejrmVf3LAYjg
fTo6L6URF5F/iCsJHZGblRjVFJZqsPwC2vLY4odBncoYsbeL3mAH152duZXWSEU0
XKP9HSDl616PZhKGvdE/qEJ3jfTUkZ6V4XcT58cHKww/kjCbAJwzPiZW8n+GFazS
MDsr3YCRBo5O1Q4K5NBg/2TFBHS/HhH4Wvy03X5XPZtJulN3BBcI3rIRT3c06+bb
A00uPwUBwqxjrg1e7kZx+bKFVwVz3+hPnH244+qRn/QHOEnyCLpW+bnRCHKrXsI/
R//ZPauKJD8kA3P/5i5mZX5s/GaHWSj7kNVXl0HuAcS3od+EXuUj0UIxNKW4TsTk
59KBi5XuX8+2dolQm7REXssd4MHkqGoH4lEKZI9rGDQEuq2iNZkpmf5EdGiRsdJq
0Z8Dq9sc2+01rhTj1HIqMMXadtUYbRBAcpR/ag8EtgAF3sSsCx8qKzvRt+XNimzy
VBBZ/A5CLhkA2rlPjOOoRghVZBk+ugvw/egQLuo4fpt+PT/UC0zJvYUYGgjAFlfv
UxD7UwyRLeu3OhkXQRxHzLnqNNXcziSFhFfE01e/tl9JwPeWd2pZfQlQQ4xwAFr8
evLxyznY2dPFOrcZi91P9cdWfzp/EckC+MNWS8SV4vvBoIUhBEGLS2ZG4e8H3/21
20LBFMbU9E9bd5qEXCd1GZ5ENx1tVmafZlGGMv19jCCB5N5sZ3Hk2IOoyMbIl7uv
KKiz8w17BmE8u3J7KC5lzdAkUHa6p8etAoBPsWZtMMpO4Vugo9DDQJBVQL7g7k38
uTmYVEd0MuRkq1aLWzeVpg5Mv9WFBCBfz1vaX/SnFr8rCILw6GKy+gUz3RihZZ/j
XgsaSc5XxT6JTapTGNTzn8F4euG9+2+B1aijDVHO5Nn4xl0fWe1MVpRrXNJwqhze
rJ5EqxuDEdYWI36sEseJ49ISUQ7f83lwunaqsZVe6uHi66tDv/Tsl6PxenHrWKrD
5r9JZLl9X5M3Ttp1ljTBqJVhZYZ1GsIuzefPy8aAoRkFdn+9Vbgy075qd6rDxD1B
Qm0Hkj4FfVV54xALdwM+b8tI3BmCI5EJ64gXVdikIugK67SsaBPf+9WHrXxiK5Bj
kSLBs5l8gua1AoCu/K9ZCgeuLPDWqk9Lylq4hqsKUHQku/57TbxvUhif3w2rF/bG
eEKP0lX3NKlfuer4MgHGVQPcj6ImVYiYJ8u7u2wtF/F+OpvLhLtizmmThXT4Cj4r
q7W/v5OvRpvdEOupr1/KmbAMtOAN6vil/955zS+Sg4B2Ypo9agPtcHE4noo76uMQ
N9kAC2H7m8+3GesVMPOD/Q4s5HOJleCtMsLe3cElcUFu5BMrbmL5cNT1o0Ifg3f2
O5DV69qPrqfuXIVVzsZHGae+rkL+lr7XSjGSouvInw+y/DY5IuAEWOd1sdUJfdBC
P9MajKD5E2vwzZgTV4FEjIIjHXdu2m2WMQjePfWFyN4JXKhOE+0RH0rGfC7jbtDI
mVjHDw4ZSKk0w3Ee2mWSImJkh7ljyy2NNMY8VMwjEqZL4oDYIqAx5wKax5ttmgDw
OdUEMUJrUFK2fBqYXa9jlaZ6fpMM1yceGsn8qo4V3QWnlm2C7Tb9G6VbIcT95ok7
pqpkDrvA2PlM6fJeg9RJe1mdLx/JqTbfvwKtNS3VyDJq8F90JaJLPQrbEAtbnKFi
oToA5W/wVjLQO//92GcsSt79xPMiu/Q5Aa/4mEUOzfFb4SNK7yrsGXH+5ABqzP76
H6g6hXbAWqVTaZHTCEnuDw6ulJhMBRooT7lmEbYz4ZjXYZbWFToLu6CtCz4PKuWf
i0hZherPY2MHFwdbrCiF2b0fyl/eHfviWKM0pvMl5/hWkUTwLUG5+M0sSjMYJVgZ
vz+YMc0z6lBEfyON6j80Q8OIwsgNj5xWdslvBluGglDARymtOoT2LlQqI17nkl5x
J0QWchGtHf9AT8C1H3tWGXNjmdamUYmQYxtDhAQwEGjy4mybzYm2Ym7Y2i6cPrNX
yBjh5lIODCHkJBQKIkpY6TLxVocFki6k/aPzDOvzlodacEVv5ky5ZTrFBx/MAfbT
NtuKWQZ705E3J1EuHH6TTEyyfzBM0zkXvIb18Vv4OjpSBe4r/cimjUENPuqIK60f
tJYdo7vwBOWx69mlfCdCBT29SYWspsvGXJcpmSuFCxq+Buoy7w7vgoHiEy5Mdq/S
X+6uya/+9sqF28UGYRwYi/btIr1pyfJyEUeROlmQmQCNg/B81vPNk0BVG4Gap6La
u06Fpop4C5rZjCf4/Q4Tgk/Ir1Zc86ov0aOvp2DOIHZeqIWtSUoJsfLhk73SpeWv
WncDzn8OhsrJBUmdru6g2ay6e/bQfS7lAYmWjzkWEWeZJbmjpnRTo/qFsiqF9HBJ
JZOHAWiEXN2cKHH6uDEsWmgbPvwlZj3Qmjic2bTFmRvBeqDKmBYr8zVvacZOl9tk
U/UfvOr8VaMm8Z5ajRgTitO4zg4jcc9/ordJ12ywSodsqdiAUym+uUZzE9V9njhM
0TetqK7L3UTLijtQiPNEvsPrPvNqC3UkPM7Uf/zg5Rdo5y46K49e7VGHwmGqP66G
mRGJEX9Qz5aBEHGjimYsvccw3fwN8J+V0JomYgeGsgpx15ZPsTedI/VLOEf8v2Kp
tH3uwRrKj26DrfZW9Atah8ZUHgyBpG28wPMU5vmqRrRbRY5OnI/giMeLoQR+ywKh
UdHRE90yng72Bp3T1P6MWKsSG/30jsdVRK9fma/2is/BYY+5f5meUxcumI+Nel7X
+kkQbJ0VodRlUpjbb+lM+LOzgrLywlCYYaIpcUhaUa3Xy8OtfGUEqgknIEtrOVcA
XDkLewxbOhyw0fdmzxrG47ea/fmwDhcYBIULaolHlPFi2DouqGBmyVN+TJJa3XI8
C7MK/WaS+T47zlB3ZVcWswox80KTu0cENmdHtcd9EPK2Bwq4PIgD0O2O7t2W3Xhe
Us0SePUiqTaToQhNbm0X4kZIS5QFV7OOHnGxGh32m6d3bmYzMIFoA7fqVQAqwqYu
glPpKylDyDdIhxrlSdISBt2roIjg7ebUvI0cHE4BKKpwUslwZ/hY4JcVKUwcK5IZ
3kKzLoyU3j/QATTPX9hyqMIyjRj0nCdNExa+yWJJgudZqmZ/5PFrzx8RufAK81tU
NTNljsLqS3h6k2bQ7SaCKbUUJ3q2eBhEQacTfLkQM2OKCgQcL8qkaa+rYG2BDmUq
pTfcXYFZDPQd6GC7an0nSj/qBpGhVYlpYEOF4N5og/1oJ19obQ4zg+sVA1Rz+5jm
PByH6UadSpU0teeZSTNxolBd4rzAf16X/rX7FwoZRvpHZhSAyvwmhC4VYyLjHnCm
WKee9HM5aG2uy6G4Yqw8t8w0Y+RoWT+rEiBNSgmafC7E6sW4K+S9T3p+7Qr69USt
4E3eQKEF8/n11HBrm4KYgnoRIYrDQa4RD+O6Y4mSqyOwvJr1p/TPPD/wf1MKR+yX
bWkelY1+Vre2+1Ko1jcYdrQVGOlc6ktzkVtZrIOIABIiHZKH3MciWm7QNluOxk7O
JqxwKgQt1pVAYAGMvFySmx5GtnuPHh2nmifdLDJVTbyEiGhsrtBe6O8iP3zZbvPB
qGcLLHlzds4sKmRNQs0F2W3u1QyNIE7++7ePwdXsxdAsy9PXNdznt4wnJYrsu8mf
p2YZkFyCZWT7mX+lrUhdKy5oy1mAEeJnefvDgSmMmk7trhKk6/CG3Yqa+LjXYtLu
fZRhgLepFnX2tq8QROPaI03+duY0cmpswErlf+5PpCTqTN5GiAOgd+oIiD+wmg78
DeVbPukDJSPSvmbUD00zg8udZHsH3DIzG7H/uCqKRn5s0gberjVBHCDy3dhvWFTf
w2omkyGooVPqGPg7RwouFfE7vdH8M6OztWw/p3J01pXZ0q/MJ6tf1Wt8ctbWQkJU
8m6sbvqslGG0jr0oixvTk7d/fdXBBBXcptyvZl6j1FzqXdBc838NCeqCH7OMIDmi
8UR95TW5TuNEn8uCGsKehVhU7cz9RstmP5gEHgdppiaucpCLPFeB5FCUOOi06qSi
QOaSgjY5yai8DXccJ9Pgq09+E8igCfa28IWCvvN6dlxQqiObNxpyWm/8BIp5P9ba
GpdPJlyR23lzWAw8HeuEHo8cZCghiUNM+mdHgVVW1dyJOpc2EWRfuLnLYP8MLh50
Aj89GzWzPsk3SoWglTQ0MV/kfYgnocxJ48Z2UsJ1Shl5tBSFlPrUpSC+Xy+igRQl
f+9SKt5ADlemUGQSFbpFG7Cd0zrkTcUdb0NksTFeAU69e/+SrhNrm4F2+f4fPBIJ
ZltM+AXcR23eJbqqIlEIXGIyUmxD6VojDmXP0ozt19YgdXCAAea2l38MiJoqYfSK
7ySmg95dTFeFo00acFSA4doh3TC02W2+kNRDhCAkvMFz/KSDh/9dCx1PRhpU+UB9
QC6Fi50I6nu4LYUAry4Y9RqvIjgo6gUZlhAtdt01MObN/E3HCTlSYnm9r+nCwRoO
sjrePQ4bzousgjrh+VOkJD2oGN+EYXsMdqigLriOK1ujvbTwqCOig5Yg4XuJgUEm
/Fto7kljBxO7dt4bPAhTK4l5jgpb/Mlv+nvLCfkF5ET3tbCzZlkjkqrCRvajD5XF
qQ659zPoNAPIZXwBn+19UGUzqMsCTIIDnKjkFUlsDUhXbTD7Oap/VqQ8dI50asII
o0f4OWanb1jCnoM9KObceeFeKE4gQbt4fUGXZt2N6HUEWqxXEO1u/zPXfEmDlmur
Pqtf2WhtNoq+hF/ieDZac+vN/vO6cIj5wBFYJTyvFC449gzs/sp199e02+p1FacO
YG6oR7IXer3iinbbWsTDlunPwOiwiG8O7yP2AD5hJApFB1uP57TsBdJ7OX6p0xVb
CojOyAwqBj1n+5hWWhsa7JEenTaRHBcHeDnnW9ZZ+1ehyWLYlhZpb2lvJP6XyN3y
6Evwap3o9GXdPIm3eNMtdPzHr5nAeqToZSzrbbYI3DjKVOzl9erg8l319Ct1NSTn
TAp8Sxob3XaV5Uk92o++k4w12eTnS8awBR6L1Ote6R42OG3qNI7RutqQNvsf9fxB
ffZrbyKq6gIMMILrKIqEnt0fHM5Dv+JsFN4lsF9r9hi/ekNY+qWNYCFo3zy2yMQ7
QEmNinOr6ce2LqybO5s/nlCx6ZSzkBADHOPQBenWBc+w6GAMDVLutDYHsLn1wN0+
L6qBy6p9kDsWL2J8/EHqe6zqk2Cuu9C1Tjx/E1jUWDZHtrUGcX6GgVaDwx/OFPVT
vZvm/2IKH3O1qL/RElzuBpoVjbZXGDwhs3VuSHp9um0BTU3nuCiGpZs6lfTdVR+4
xPnW9zWOLpfWrNOf7NNS7og/N897Q6PI9oUtA9D6li+aNArsF72mo8QFDtAezoSF
rNTFrx0otxkjqXq0YPSANbZAibdPY5buo0MaYWDLAcn6k70n+532Fi64P0RJmU9b
k5jftOYqcmDSMppY1ulv6bkUKmfqM6i3G1oKhiortsA0gGnGclut2ZS68liFfjW4
sY0o9gxaiclezGeNEZ86N8fkEzvGFAut1ayUDz1UntL5WyI4hdclA8QI6fRvQN+3
Cg6PDj+2Y1Y3mU3FG72JMJDTSSHfaW1HBWFDuyPC4Jv1Scw0B2VgL97uH/BjWisQ
D4MmpdmaHhe8OvvRPvPzhFPr4I3FNCXUk4znxFzK0Fxsh/bMWSaxyz92lywwOUuE
GR52C8wgRlUeMpnaSla1iAnNN4Z9a0bthwjHXpjqpVfknA223nX0gvvnp8/iJ32N
r+6MubnmXv+aWVqshSsd1uFaXLXnIrKBpeTEBK5kSlaR+lPGpEZYQQdLjGC/pT8d
lmFlOWIdjUpd9IsZpkjxPXNcH/4Bn7en+D/PSVfne4K+YXWdILsh9k4LBpu0WcsG
tUi1tNirhuhNhGfW8CxyyvbqkCnw6jCzs30d78ucgfIHmAjDwm3luaxhsVhfIbwX
fw3WcYR8nkcriDb8wSXi17kTzSPNcudd6yvDDLoQ++epiTtmaEk4D/lFo5OtDSzN
IKfMmlDt58sWvvusOBQvMi/xSwm1rZcBIFwi8BU/2nq2dh+N+VJkOtR8fbPdvtgk
0nKOCjAP1omTXSmx3E1c/eFVoKKvZt8ytXYw2TAgF6OliVL3DbGSMoUjx50cePtd
6GqDyOp8/zk0BgMEzHQ8PsIFJq7x+RHS6sCXJsM+rdVTIWnXzy6Ixg2W3TOBRMFD
1saI+IVKHiiYlCBkOV+0Zef2FZbF9K+ZameVE5Cjam/UDuMAg/HZD80N9uB1qy5v
TL5dpSn8xF6XhU1BTabmSSnS0M8j5yDcv6N9QirPVOm7ycF+iHzXPM/JMF21etjx
920IcdqBke7vv37C/WR+G1qlGOYTfTFiDwF3XGzpW3lA95Z269UpYYCuvPLvRo46
sI61ulzUYTFOOGYNsFe7bFnj/NB8Dq62xSbTshvOCm/c296WmMB1r37PLJO2coEn
gku44gi2a1pKzw6Jlj8NdVIgMZURJsbC6TJJGSDJ+NauDPmeZ38BSK/a4mlgBBjW
+IqMxWB0aoNtxQLpc0Xx5BmzjovdaBtEnzLvFJMYQdwAAlVXFdqD+1OnG0O/nX2h
aB17gN5O2MJXQEfLzcFTiOHYEFto3qbReaoxHzlqNKAu0fag+YJZPub4oOIpqHTg
TF+Bi88IWX7wOfcGdb9P02P0F4Lk7UbHQT2jWDWwMkXTdOhd1tVIThwdpD1jyf9O
1CX8RBpxqawg/Zq3KEpHxARdawtbKDf44mdbwPprc9YEKap1O6ciABxhuFqIV0rF
8O9QMVF3+RDQ1Y1q6tAZBUPeGtCJmVn6YLFDuRvhs3EK2/19viancBPTHLhzpQ7S
LAi/OuKZAMCu78VCAMgBGzxLvS7+QWNx+kKGs0fAxeCoGofKoheYfQ54xCLXkzxn
uhHQzATVTFDJ5iFyLfVXBAvMljEymHxBGVAb7lOsVtTyFoO/C9VuV2eIlniO7D/e
myoOTyn2T1H5FRfC5pr7xkAHnsm4Yh1t7oIOj1DJL1MohdPDLNiaknLLg7uuREY3
gc9QwUVuL8Qzhik+qrzo3USuiWbT1EKOpd2lSBdC7U7UxbOdgX5CByyXR/r6bLSp
ybEPbBdk2tnMzIfYySCcfzNK8CKB88CF0m/TLt1vs6XlCUdDmckINdTzCAjmBk++
JrsEtrfbvtZNp9i1ulBpvX+tCbD7HJKKeuLbZIMMEEVhEDFJKgLJSZG7AdZluBO3
ymtrocZq1Q5FFmBbi9OmxviqOhDwKjKdD25so8g6UfleOtSxlrT96Fb/pJE3ca6u
d1rHypQs2fm3W71hRfTTYQJ+XDC049aObSy5UVTxveY+zSSutQc2AQ5+yDb8rVv5
4/F4yRX1u677nI3G8AljTTVr0imf+jm8jzOxXRY+Jblc6CPC9AGDYiRF/25V6VgL
F+xwQaPMrZLw+rPAxP220Vuk/UloHWFToZxfQuqIOHXYxltCCILSaEVpXGYtUi8t
Cmxgiwc92ofAOA6CL4oEU3epK+9sqn+3EwLn8uLVf6uv/tssqB/DEVE/EcgweGCf
VdJZPN+PabVSq8xXZZXO782tKqJqXL4kmZwDLV5zZwaRfhhhnT9Bj2iZarITiP4Y
8gMb03MSIQvisJtSG9on3e7TBBTzw/tcK0m5+L+oRKdQjalxpPjZG/A8MFd6jXzo
YrbnuK3zT9IbB8ZdU6daG7N2Jfb7WMptqF4CZ8zXee1Tf8K2aOsvENPF9FZJ0LH8
/ApqelKrovnT+tF5HncjLta2/bwqdslLGLIwwpq8MKs4suhPxY1nsXXPneh+sRxw
Hod05TU2Cr9236i7OimW8MHN3Or5cc5XGPQtIjqF/+qfgF1ggk8ngKrUBM5TTy/F
5GhB2ohriePaHuNOTwEr/kmA/RxjxzUiFkk11zWsHZcivwffkQhdRycyvSC0Tj8k
kcRHyU2LPZtb6EZyQO/jt35ttH/fi5o6FT/zmag3YRGiWn/DuMogYVY+Wc1chZh7
15valdy8sg0576YBE7H3xiS8rtdvw9XAQB93ITocv3gPZ25d4lM6wxcYONDEqShf
94AdAVDEr/quQgnW4Twfi9LO6xiREQD2l9v/WA5I8cW2kuOFqQL9PF7+zk4hsBho
1mwywT0AI8G32WrqMo26drSNnwvBMKoT8vdsz3RT5wZ+T+BqZ9R2DyVKbyKuqyou
Bm1RHhjKiQDVJEiMqL0cMt8AdqMN5WLvnGRvuia1LMWuVGjjXTLD6JZWZt7Kc9jg
S4amm7qzyyUeo/uV0qcg0hH2nRgn7Dfr/Xm2ckJpoHSX86bIzd2+3ku+ivA0zllL
4Wx3Bpj5OVpx/t/PWv2eA5IGa5iLa5zFrP5CyCngVNEQ9q8xK6kvJibtLnC8Y2y+
9AE998kj5lxrlLJzZK3mQoj5YbYQxNsGRFMmLIx7pIVU978k147ehh1HxHZtmc8J
WRGIvfMBSJyTT97jsJ+PYxlvS/DjG3+7ikWQfTFPzXo04GfL0a/dP/DKYVzUyfRs
V8YRZZdMbfZkphxYgNZ43OAJrKnGgUDhJ51tXtucdcHevtx1ndrMkDuyVYrhFOGN
4Nvg5fQKGTG7wZS4FxtxnDTX8OoECGSm+SkuruzlbCegbZgc9aaLDxAb0lfJEz1G
0CKa8lFwDmJyuZQchGTPiuMewi3C0FR20D3QwhSrC5ELobPVtaouQad5Cei7VruR
kEoLvEz3REE0M+E0+MEgWo3WKomYkTD3+UDtQUyfmRadhNzp5Hf2vXeSlEspR+7K
2IWwd0USVZFfNdmZXQb+76XTGh9n65n/lRyFebg/r0gLXv9VjA0YcwH66ODmCfkG
rXsUqwGZaldBUs84rXVx3rc+gODXJrkCy2xHgH8/PDcWlqVYNW1WKWqvi92ymP35
MJ+3IMikJTd1hVgEtz7DuEOj66/Cbdon1JLt6cpBjToB/bJWbRUdIIrZuRY3QScP
ZR7w3pnAJ3GPj/2K4Rbk4uj3cK7TDBFblah5DLXQHE1JsAHvfviuHWkQ4+u8admQ
Iy+mT5njnAJkJMBTzbgSlKNXDkeD9cY6bLvvrqhlNQo1j7VDP+NWVW4G/P0nQCpp
m+9hY64CAxtpLPi3UQMQJk5UoUIXchNm2UgzeSZCVMexN1KfBsSgEwlNtuBoieBI
dux7RsBAqQZ9Atlmq1pKPll9jDiNOPq+OzRV9IakJ0ISu2sbwNaCQtFd+J5JXc6D
zHzVjFoWvM3gCcxHVu78ag9gS1W3R0T3DQ9Usyu/YCLt2DQBpyIAddCOKoVxcuIK
ifshyHj/xkk44G532JvDeofJcJ+tgNHfcgMJPYllTgQnlAFyRoF7u3hSPZlGelf7
seHdE+cQAD1JqCzplNNNQTn3MpcDCI400hGBPA8L//Cfe88NJPJKPL+xCfP3VR7o
/aWskJjJFTkY5D/7pAYofmdn5ItX/geVGv/RU0V5QkNZxEVtYtzngUIGZMIjT+Z3
ulIPV5FpJX+LxYhYrUn+hrBXY/1PJ7ohELwrqm1p2N/p6L/uFS0qCjr41Tv+oJKA
g4Cyt/XrOWSXmPXpMgbQhUbXIwyU4ySdWBrDnjcmuj2vYEas28nKWgkTXfwf1hN8
2N0bYqgrB9p3bU0nybPhgSA+mMDTRMve+Va8wQcStweR0xmwpdqWqKp16ibidblh
g65DpalUyvmbzKc35T09bA1fZunsHsucDITfF2ypf8wYXo/Yu+AkU3vWstRo0UEf
GIT30eIhK3sPPT+qW3FM7PntPRxW/dbfV4tZerP2GWM4XzXUlmQbrjqs0OfAfbR4
Pi6eFndt6l+zD8Gbam9dnORebIeWHbo/zPkjgVojVfmI8wjMl0nOLYBHumDOCtdV
GCz9Qor7PXIVTqeGPqqBBdLkBolWedIH2y9+VZMB0BCAViCizf8ZSq3NywSyIAbU
rFDa+IHUyJuCvkojlu5Y5MK4lOkLQRqzu0nriKcFyTxUioZs46NVA//IlympvOiH
LzacRM+r0T9sWqiT7OO/cSj7PGf+CM4kj8RtxFhrGnGIF4sMhjwUIwi/4Sz6BPlr
LjyRmfY3avrQLXH/PCe2LVBztP30q4WUWTdpr50L6vAzf+dJGSZ5yCw5ndt06bpP
vJEHcv4dBfPx83TwGLe/63v9B8N04aHEjqWkQck3WrhcG34EduXZmJO528gax+et
NFyqRRdssNAX/kaJsLdxF9ClOSBcmWgd66qffcJk+OjY8NM6q41q+lmppIbEFQwt
ggDH5jRaZsu2UBXRqOj0W1xdoss4DFbf7r8mLO9AI693YQpfceA2NR+CQ38Wg42J
fae0/MgBYQC7kNNyl55GQCJtaNrBYvr4RievzKb1JxP3O4pjF5j31EazSiqf6+C4
xHzIMwOUHRIJ7oXQp9qoLiAXz1IzNIRQ+g5BLONAaB0pO/BZwtw6IUNlUa8vcgpS
kT3jiXBR9dKe0gNzbYD5ut9XB14Ui+CRtn7WAWP/2F8dJ8zdxmjS2Eo5FUp2N105
yfzlhu8CzlzAFiH5DL5KCqwqbjYg/9ddmNJWxX1QsjFAMUpgr9ZAehUmtgyyx1W2
aqQXYOcNOg11/JxT9zNcphg2qOKSRExKaby7aBvnNPyYX/USxy6Pkhz3+8zMu3jF
c5AtBmV+3jJUWIrLXPW0IgzwxRF3bgrH/ti2+zYcmNKQ5da2DoPansHP/JDT+tv6
17/J9FnMa/R7wWWgXa5YZPcDX+y3sM0U/fK1Ky3iCo8mhAg7nm2ctNC7Knd0Kajr
UNmWjSmnknn5QSvwVF0lBNaZlLnKZEXzleQTG6CrkYArK6vt4wTZU/GzEXRn19Ov
pC96GFRSt1SDXPvtHW5xAdFwOHedubSwuM4QDJQ/st/lYaolLtUbDBjyfSkGkUW9
ytcAvjDmrKZBN6xz14sUpIzbQ0VKnjcEURTtII80NxI3uKwQOxDVl4A2xcQu+TYE
j3IzyLIog27kn1B1KNNzlxYgXiAhilHjxoKenNeTCrcp4FvSZ2P92NDUQvZ8beHi
AM+kFEwU0SPRcSE1jKuy2TPY9KpuFv1s3cGKDxE/yLc0v4czIa8KfzOK4MXGVA8a
Qpj2hAf2+PDKWu4ebPpnIC3ADaP+PmfDRvlc0hHEb+jentCeCyGlNNgPP0VtQFrA
i1BmJ6SYpTlOVeNQO6rquaoKbrv77P4XgwSV95TzRbKS0ZSUawfbciDF9HOJmHbP
RecKrfsT7GP/2V3qAvfCgAdeFF9xiwKq7dS/jsspdVNs/mwu8Fl9mTjwSlhnGPyz
YvEPNQxkUoi5P0kPoOdKQe3QzEiAzKt6O9v2xiPnVYQqRxgbaYsYwnuM4FAxrYjT
DAUwwRj2HK59AYqyK3G2Av0ySvyCioFAOHgUz7No2Uc4DqfD1y8JD9zGBKZHO517
gmKF8TTQa+Vlg6KyboIHC3vnuYWucep2OD4YHzUi63RDTFXIquvgHGur4lAMlUsF
zEwRUxO+CcFeL8fB4fCIWVw4IixMnO9L7nFH+5aBOzCEwUAKvR5IlIIzw3XCDI2O
eez0qGOCVB1JGQ7u7cnaBCnnpPPLWB4r/yXOPb/41s351G3Y3cKveg6TxyhkFKx2
7x23XneWgpPtvX0cjWejcKIRDXaFRvuG7tAs1HjwVVY1mZSJB+2BWO+Nd5E/O4ak
1FRJJvZ9U0P7S2zNdmpw6l2DmTpDvlf84IkCwq9IKl+UZAd/uE9SqbVq+OMsS0B3
2RQ6jMCbd8PG/qALJVu2z7JCRgvrZjJO+E/HZ468NNK4SMwPoNYJKEgNcfQSvxdo
h5iohj6NiSMaox8A7aBkt7Vi+kp2OWiQUZP+jRmBT8+CeiBXJdjlmvdTSXk80JzF
umMgMU3G2MVYZ0iJtLoPgpco87dpnsoOrFzDiFG6ZiCGOAxInAPE4UEIsBj5NNdY
pMvxmQ0F5RKdoSqPkUwG103Vhm6isDl/LPGQdUpPl7IDYLAyacwUQ4L1jPs8j+dC
8xy2Qwa7oD7KQDlX4biFFmdsNgnx8OgLXImxaHmIwMCqXFvS/1h/gldd/4sV2IBj
CVmzTw/mHh+X50ha5EMR/XV1O4YfA4ROSrcg1KDNVnFF0LS6KnbKxe0VweMlcgEh
UoFxFKe0eO4GqI2M9txQ+q+hDKTdk67DGQOA1NX6uIWOgt6izQzQfdX7f4CYIZWS
UyP37/HQgI1Jm7jtUBHDqc34xKSH+3pvrgbm0mz94NS9OBgep+XOwJ4Gpx5O8B3T
aSNmKJnkkfNNs7Gc6q3DnPKh+rVD287WXIOGIghhNcTrUGchZcR7UZVkE1z+w9VD
IeunepvAQ8kZkyXMbDYqsDz6k5Ln1j86vcUtVVckpkwOo0folNrqjZCKzph9vQu4
ahziZGxXUDW0pLyIdsIRbOpdcZtCp2XazwqY2hnd0WFR9yClDzbHSYNVpwyT6AXj
NuTeEedVFZvcYE3u9SJ6LZz2H0C8Ol0OEDWK3kdifRspO2sBjWNPNhr7glEZ8mFF
BpFdfsP8sMCuDMxYGLYf/cXuYsAFAUXGAhpghjmyBqeA+3dl2jw6WOR/mOyQkISG
Ac0k8/O0pxS+VOFD9+kUsk3xTrIUKCgY6ofGhZMPWdwcFVTYjDWx9mEZTmZrpRmB
TQvkLIJRFDAWkRT0vIbaIq4Gm13FCc6VpV7IfeWQrk+gFrrqqJgikIqeldi/96Eo
to6dmP9+mF01SQ52LCeyxN6r/SDwAvMoaXaCAY0THn8qX1xQFo1O9T63BHPhcMFo
WG5laYlh6o8kxND1y9X+i43izRPSSGiGJN9143r2uEFO3ijTZ0d9YeeQ5OVKEF3k
iQiy0+eMhAD58QlZC4B027it7lSjkht7DWYypyyDywp4SxCdF1NvtYfWnag9Ev1E
F0chhmsm2HZOH4WoskD2euyWRUms6nNj15TUjAGaaM5MzC1t8IvuajOTh4LAYMDS
pyfZAyHzb05MVfZTjebnju1wTdYoXkvPRS7LdLGSEYKGtxPi3IDraIiGTeVsy03f
+lLPyo4HYe81tD3leqHxyLakgVWRj5KxXuEXQ+GRBq+6A5m71Hnq/PGWm0Vnmsxn
a/N3WG/2tR981I1tdaLCnHRRGmpX3pJfv+zqoIKH01EsViil9GBJEoE3vp1sMpjD
Iz53R1l/egPXxxqpwIxwuMeHkTw1QkUq9XZpBC88I07/+bb+lZ2YKlf60mdZMgMZ
qX6Cm9eB/yZG6ud/cWZbvjxojjFWMtqWgmwQJX37CBEVl6ljUieth/EU9krEyd54
NCo4Yym0g+ETjDoQd+FOBBsYhADSUoqfuPzwQ8A4tgg+ljfg4gzoG2PyS9ZKo5uc
UZZiFDd5c76GGkpZMlvV5p5kRYEGakRmxknf0qSVLrxgQ7HKckG1ps1+WNMD/hbC
8W+C9COJzS7u+6YWqmpavjsbU6tZDbkUyj0yII3If93vkjdZjuANozQDz522BDBW
JqHIcIJe9+196BUv70ofuKIcaRzYJ4ItiA5BGlqdH1ax2aJf+QJ9mCLWT/UEt1XQ
ozkIEPQ7Fhf4K2ky4rpHOGXRds/Sy1HIUArxnmjyKqKq/1Z02oRziy0UJbqSmRDX
70+206OqhgAui9p6UOA2TxQH8S6QN/huOcxJ7QpzuhUH83GR1MGq5psb18hK6Q25
CLgCZt6pvU6OllaUZbMWocrQWCpJLrbTHSAj6E0v0AaMtd4Y3SFek3QscTgJB2yj
UarFPC2OBdNZcWGIQU+zyf+zmmzLphMlfgKF2cZY677S3tTrMDUtbg8PQKNQ34pb
d5pHNijE+MZrx/cb1VXVlWKDzoZ903C0wyvZKvTePUG3jCteU75KKI0ifEbiarP2
/k5f8cicu5TtoqShoMAX2N/Nfck++hDNGkIk1L0ma9HEnsZZ4Souhftq0S/2vFUg
gelp4l2hRqbDAP7RR2Dr/59yy67wgJVFXuhyA69TftXI8xrfeFDE6hFDH7ZKnRsR
9/WIQ7TEo/zhE4g3Xdsf+23Wa7GiTFxeWGyEegZLQjzIXNpXVK6iUJNrhSm/MqV/
etPgZOWb+PsXZLBUF71Gp3Cw5/1kohBkiJx6wuepdVZdN2VmzJrFm3I297PWNcr0
JC10hBFHgXiPBPURqjL5C89VXlODBDzKH6M+HrBEQDDlutfB0UsPh3c3vwZski/G
krp0DrZajuxmbLny+qV3xei9d32cODlSA3NzLV6ZSgTPr/rlK3a8giY9A9rez/vT
chQTJLpChgs3H9jjZ2DHCVLqtRpxPjnkF2jH/SGVISCwWZdoy6M59RE61P2LG2An
7f9HFDpGqmi3/C/Wbjz39QYRMfoCSb3IEXUqor4HcHpAOydQ+twVpNbP4TNYY2x7
s69lPW7IMuVxvOuTPOe6r5Gw8Ea5BG/8ByUg0ANC0EStWC/+fJhUp3AKvZ0imRZT
CYWPpCgdTcNBBgM2d9iig7ydrp8+sXuyzo0XMM8P/G8YlOLflmEdUSASCC81Ok2K
Il7wGdTytR7H0pOs3YEvRIWYhVp2fOenVvzLJ+X+kyZqPzZVjzPkMhjxpACswtzj
UcMBVvQDZC4GOJpSBTPO7xIQYIlv5PS4foeE1ISmVSU97iPJJN/RU6+WD3/brEiv
f2rrLx5QvxqoyxbgMLSh6RMzwgldwm97SeEYVR8ZciRGVSSv7cV9qE7AN01aSJz5
R3H7gFxDHUUoFvVpY9H6Fs7Ut51fM63TsiIAHbN8lgvIO+GapSon0GRNC2nsPRv6
Zr5wSMLMs45/oTZok4rYMgojr+6Am/gs2GunZZvsLH0/gxrjFnng9aB0+3Pj2Rgk
xHv8LMhv+2wFve97Brbc2Z0dZd9UftwrGNXZ1jNAKrXCTxVNNEiZ0XJaYJCFAJ3Q
LD0DBd+gmiq+5dYH3hIgQoAu62XsBmre0Q1Rz4BFCGCqo/8nV5V8IOj2l2hyUCe5
t4zzl9lLjXXUHxbaW7XOW65oG909UynR25pnjU72lfzJGiLr3hj19+gaG/gJ1QCw
LUOQ1zIxuB5/nnkbtwP5o7jgr31GJgcEcZPLKDZ6WzI02Ts22175FCwYyqPldW4G
8n2YrFizYFBcjMh7aR5n5APA2JdOickkcYMKYITf4j8wI8k9lVmmDhi4zOrIHDOs
d5fCK7ltpLAuIW5WQumZtrmKwayHmiAMoN6WPFSuJzdgyOoEE9CVpcL17mmDn6SK
u2He8tUVbw2f88tjFM0TRV5nxm2+VqNRo5fZOZWeKTOxuXg65NIL4IWAea/3b9B7
kgiRqMfHqz2BRsNF7fTW+52ckCz2Azd82g9M2vs7tF9G8FPlFGQeLE6VaSMgvEWy
Z8wwvMbHmrJx0D6ezc9OrTK/0djzU+LXEJ8gOgiqDLWVrYaQD9i0yM7AvgoD66LS
dXnVBE/F12CQZEYEMj5iKZkg0oBS6sPx9f0dIC3XPuY9a1NmP6GMxrOJ0R9kFONO
qjEzJ4pG1nVW7uUQDMz8wH0DBkcwpOMinsxn7I4Ew/qOHgdCVWQ518cITGsv8tsG
YDdKt3W7wt63iDizYjHb+qVoryjIG9RPzYwy0QnnrYdmmRZzpxn4KIoICEdbH3pk
QDnGdhfGpfTv8tXOQ99+Xg3n5rirc7bco1FV/bIwMUj2anf5Zm+k/RlU3rcKSn0y
qe2LYbuXtvCTZBnsF54NGZM/T0WSC+dmnXhqgPx0TuQRMmcWI/q4zwVx6/PTHQAR
AzJzVlT8BRMzG3Rcz7FmZW5HpFDMnVWX8ugK/+gDKvGeerpdYkWwaetHQzgRl6TW
ltFVr7mTbJsnuhJu48yJvbK42CXTciRgCeA4kHy0Rlj/SiMtzo3FalUA+WsuKbMf
CKbPwwE/RPAJ3NHxikSoTNOHCvOo7dbF6fWXXBO/NOZprSXywNz5szAj2J15IgUR
Vynyql6OKOBEETDq7qaIdFcaSZ5nL2rjlL+qNxIq0JnNP2L4/+Z9QPlTOG/eGt8P
0GUz/yeDN87fZoS/ttF28sN/KxQGtBmNrz6g122lxylr9i8oV3nXz0iZv8j9nDGX
RTggcjKuzPaMwrI7Re0PVmTT93wIrKT2ANmVLLCDL02miJ6kYXxTD6ZAxiY+r6Ty
hPkxtuOK+WlcuRlgt5+HI9QzwlN6ZItMDnwuXRDqOH5rQb3db2hIen+lde16R3R+
eAVOf+fBp4s+eMqk5MDnhTLqBFe4LaBVX/SkVo3zDEnGlFPKhhP4uaDELxzhYSFw
HRLHaAcpLL2/9HuT8U+pQzG9WRPtELVusnHOodW8CKF4muX53Q5D9YR+wxoeo/26
eDOtX8H4kRjvf0ksCFP+mwSDtzCx87Qckh41jTEmkp2lW7jfGxGmslg9k+A28wOh
SUfQhNSnu/4MSPxWQWFuM5vHudisisY4ej2HVRuWlmqEa4eNMYw1EQtMSBPYH39l
moOO/VeDVpR+CsVML6V7xY1yfB0fx7VgqshlQ/hrC4r+g66HJIk93wr6VWDAai1X
xdM2wqCPHy4QrVQfUev+OKXgeuei4vA3gxzKxSigU4KqqarZiO9C+lq8P9eDOszu
+n36Hzghtr3gv8Py3UbXqYtqUXwUzTH60B2W+ogReebXWJwmBzaJ05N2WBRa86Pu
Mdq4VeppejljrRD/fiIiE94IvRO7lzRj9fSRWDtAvEj5xEShB1eZrLQfbbxKLJMF
b+VgPnOPGc13NSz49onKrQmP8d9Pl8gEKEcuDKSDS96qZGX4Mv+wxTGafLZ6Vzjm
x+qPUwDH/ktjNruM+CtxPLdz6kmHXzqIGTCuGtQsBN9xdgxlsWs3QRcvemqoS3UH
dRSluPpG3dzn6+KCuzv9WRprb66ulvyy+1xY0vvxgOfq8nZt6/rhBy560ulA5waa
64t13CQQ9cEbHNkA1H8uRbhjncsrex8r62bsDPOxAso/XqJ8v6zagoSAskTy1U3q
qXGWPPejkLipgAkMNy3yX+spTv1mR7Pmbv6PAMUeyevE0p9rz62gjNFHGsMgv3ds
K9g636CzYi27qkVLymd5S126tj53MS0wWYwE7sfYPf1/H16OOTuvytEvUevjh5vC
5Q2N/+nIogdyiQAd/Hm8j3X3Xuva05KhYiFN+a6MTeiWObwrn25+PW/6imaap6c9
+/UOnqyvLV71N9brGaVRyDiAXlrbdcsL+n3iOqgh1IltD42Pt4yRC0NqaiEJNayF
/bd6HzgUDzUqRPHxTxE+evNl6xorRJwtwEJHf0QayrKl2+RuU6+J1VnefhTIGGoL
TUvPsQUPrFFaK3Nsuy9rKY6zVTP4YrkKgw6y7n1WU0bpeHTYSeUb9QuC3TWpGVJW
dwNLUD2EhuKoUsX/2bUsihXFZCpG9wKcbKKlwpjtokT5OHhj58euXk2NX2aL1b1A
bj+Y6QpDuM887jJCMDIpTpAhGPi06u5uu15dcAnvu+Rq96cxm0KtGk90NF1RR3ZD
wUTuyOyizvR+2bGLS/XftjEYLAfwssZygyPofsP0llJOUyoaMbavznskWU9xmJ+X
bMwFtp6QMKYsV8WNvjsinu1iDggxGiz4Inv+5mzcqsQybjkIhU21I7Zq04a1VL+J
EzO7IEInLmbFauut8Rre5bO2PpLDHMADeFZnfCdY8ckpEFNqldTMI41L+gWBBtZN
jdI+yxEQcpoMtNrvn9hJkgGo0GriFaTzHh9J/HITUoea+BsZZQqDxxANmEdQ0OEK
hcLmYDF5TRuQ7lbeNZng5BacQFkmDgPtKpimTwhmfR4Gk1MQa/hmN6bt8Snbxhhz
BV6epUX9wpE1fgCtSKyoUk7k9/UrFs9jUyS5cT4B85E97EZ3e+iiuWvF6mgJr57T
p2WS4K1OZ/ltuC9DpkHdFYtRmK/ERdO3zMuKOfFOFcNt83MKQt1tHKqbQIv8CkAt
G7ezAnw/DgJsKD80Adja93nR/hyFz6afHjbbQJETMNglJQPYxAxvQe8boHkGOTVR
rwXXzOAelbg6Zhm3R6K0UYpAEtZ7lEk0ma+sG6xSQ2i5hp9GO3G0kCP+n+xO/fGD
OAb7E6GF3vkFHmhMTxcqC9d7vHhqdgaCSDPJNvkzAnPYKTjkAMsbomCFnklol/ZT
jpfon7l1v1Daixlo31TPfEu1jmCfGfZP5YCOZbj2zxYC5k9wt3XTdXSJcCwCHQEE
lCezXImr0iTqDLponOyKLHOgrxHP3avqBKAEBlgOXIyuOm4dtsNuAfbUf0qjOMKa
6gCwj2wS3jhrA4EKY0u6QYcwL16/Jj5cNz5sNOlcknO5226g2glyN/iH0oz+fdDi
VTAfKms61vaMKS8nqYna739HZb1JqbdpHUuxDTIENfGbSA96NwmsbFg/yMBwtOxs
NZ0z+S82QlnXvjEBMTPGd6BeFgPfxaOLXlQYN9PdvDwHwHHcLbNBYCL7wtkB/UZU
V7A2PbwznvwvAnZz6EnBol1vwVgouubEMNN7JvZjMkNDdx+fBkPreZcsWgBRCxeU
ErAt48LuJPyp0/E8+h6aibeK0KFoqLiUPbXb0SOArWzSwkp8y9LtXhcvc7B7PCPw
cXUp0H4tk/kJyJh0DD9J6SXPVw9UiZn11U5+YYHGYFqfjHn+mWqvF3lBji/CfGCV
BTbVZYJ9lZsKGL+azLOKLvgMXVpGEDSjPN/69U7r+xwiVcMsRgibOjFNQys8nMPU
r0LOeLX+uErCqMMjvOf7DLA+ShRPLVheAuRe8laxXtJ1NOWeRBqBXN4Y3fk0FqdZ
IUh+dpz/rxZbb/n9fQnsXuik6JbUvSNo8GwrQUtusYebUhEDUTUJ8Y1lN8bdtu/8
v1vszre3QYWz6Pzkubw6neDNkQdbSBGwf55ns5mYbtCdgDYsAgN5LioI8Q3NDK/m
X0fJNALUyAj/yvsJ8pkdrDrGflq7EvjAibArrwCSf/XrdyAyiTC3yvQILKJO12Gc
NpsIPFf8CxfGBhRu63FSF+jbCL5d/V9TsiE31VZOTihAIcuWJqqpDh7fQ9w3fYmt
roIm2T+vEQE83gESPFydT9iBnUKoJ3zKVthZC/AamsLWg8vfRp/K7b/yLR3n6h4Z
0Yk4VxeywLBOWJNyjP9aE+FH2HGZSoV/kUp7cSp8ZGDRte3GNJQ07ErnNCBcvdg7
V75yE8sU6o6nDJCgKuHoRxcRj94nX7bgpw1Z4GvY/8ZOVns6SBU6Vmbsl5rg7ruX
/QhZ81Fh8LbYkCsxrJAtWQNWjbcVfODh1Cl+jwJ481HlzJrDUY0J+gm+vZlTUzTl
lwsw84I2pJAHeyV0kLM6Lofc0fk5ykjodjmWxCGmlWpGIKKIvgjKv/1kkWpIKcPF
Mu2BoYveU1j4N/WkD/+1uHEAKKPp4OMQvvEomNHZSTfcBLMUnwAfEBjq3Rd4HSmt
uzXWqhfUx1r5vgoFdalltcUU9Kl7mgVYqIvGoRxluWmrwdruzKP1NaPohasKpazw
04c42FhdAHWZtunlUxBbXvtvLwbt7AU6lM5yzEQC+AEEMytTIYGihvnnbnGeXBfW
G2QkRdQblT788IDKfNIeSZdh+lt1NmMoRZ68Ln+qw1FQB6SwtmGTOIfN9ALLQKnK
S+eVhCS2tUOUqYhVFDEJ7rQFp1uiJCpYCqNrxLEkkgOzvuGfhojNCLBpyYlMK7e8
Dw2I4CQA5Vp3PFZb6dDGN6BGQhPzYv5i5RQL/mgElfkvuEryZbycHlmz6TQhpns/
QB5Ovu0A/FzJkfENhFWvNfYX0dntlnoj5SouJlOMAOqz6jGuzgZ4yd5+bKQ21gYX
lMP5AE3FonAmGxRN4R/an9I8QAJlYidxe5dno8ue/XNqhoHCX8GM7L2US+Ymw2oB
1Bez5Lx6JDB6jTQzaVXoz8YtUW0KlwLNyJqJjJbrKAvsCoIagKxs1CUjMETIrmAY
AnWKiIW28zN0nsg00IUO8VrATYIRFpKZqp8FacGUosr3RrLAw9Vk7xas5Zovb+Fm
dii5IJG2njz1GeBYYVxihVTgkpL9RIWy9B+OgrIsOsGKkoN35Ehr3kTLa9CsWEd4
iECqx18Dyr2v1EWle1GNYcdX8ZAUjPPK7sWChvJTplEK4nyTOKgW0EzeIC2CmA77
ysJmXKXEy0rXS6r4VnWKR5LMR9iL64XeZCU6JtHav+8Eu2d0R1nJXQRPbDJxC+C2
LKSGnf7cCaLK8dd8/OB26CjY23mCi4B2l+g4WfpI/T4XcX6OUmUBCbfP7U+Uh7qk
KMOFu+7mT+10VEwQgtItFkVZ3SLLP7QVwNNlzsyAOJJhVUtzkbscQxoG2A4ZsZbW
3WkYH3PeJg86OWniTW0lUtib3ZDvTabFgtazr8Z58tvykwebmwjmnZ45iQfHvD38
jX8TJi6+jlW17+5kSOicOxdeU45vOlrQTEu4HeAATuxxf301Jubzdlefa/aJstK3
JRd6o21l3cAO7bhyc0n7sTNLufv6F/qjQJagnkMWZuZz+z1Ce3y9js6EQRa0BDd3
tKjk9yEoP6s/DLwWz01I3NNTuuLZTBKxjSaZ/Rpp7HSCHmLBMaw6no4J3rHGyUWq
7udFBqGwNHhu3xqiN9kE2Ix/L5AID2H1oZtir4sXiZSBojDE4ELEzTOQvRkbh9RN
Z8PQpz97vCHnM8+/KPbzxl71PxJCmS6uC6157T8vaOG79muCvwNAenufm9N7C+Fu
U8MpQcnUleFS2mgb1G5rxmWq4Kg3AbixbWEcJGnm8arT7spC5uUWWoZxbn2on+3S
IxidaHL1B674phZEV4AJYDPBwHpYbR6Ae6yjO4RGuz6+LNnAlQNb4epiRFnXN9Bl
LUcTIZh88kHk3xHUZSgfm2Jj7nudD3QZXFKvZVsuaNpWLPLprdMX8/wvThOzWJCA
PTQSTxA9U2wnnltVYEuF731Kzd6rVLMp8qECI/mpCpZ+OUfHM9re4kYRBOMy0tL7
hEtTSyycuhwxntKuUo4In37eMUDnXebPglL6sw5ISslNeR4gSnVkZdEOPYMj2e8b
R45kq3xKLu0K93XuagEeA6zbVHAKONMYrMa3qdR3Lp6+zEoBNmZv0SL44itag1Iv
tLYviTBgruSwRWiREKIthjeQPqYAdKknvW09qmNuBkfnTrvlg+YZennU9jTPNbDo
YkK4Q9e7cXl8B4cvvJ4l1exZrl7o7snlOwxdMbE3kiCZFpPm9E2rkrqHoAUch+sg
UXWoctw5t1LhU5pqXN84b/TFdkjgxxc+dWMB26BDJQpUkRothLGF9yYgP82+vknB
uXyq1Y/S1oQsvMVXFiorKeSUKWXksoVsRZrhW3bUmCbjX+DawefdkRqZKVUqs3rz
9OqKVoxDAUIIj5WCj1YMrWMkvO4YKOT4BhslZrsBte2jq7EMXQT8uKO73I0Z7AZu
L525DRDRy8tzTdGfPBNsDgITFWEQ/+jpHZ6loLecIRmvWsdQ8q0MC0f0yicFPzai
xrQL5+YhyiD0hG1gPTia/e+LhTfwfdYpfS9R+VPeCER+7n+0fjnHT1CDTUqDl0Wj
SBxxiDg5y23ZQRPM7Xzd1NlGXpEVUKN4/hp6x91PN7S4AX+5my4IP7dstOXm6Ago
AZDkUiGwWp+b8F2TP8rsOJRA8PAIJhYbyYQ9L2cz6nMTSKMpkZTzxqrWMiTM5rpa
zc6uBM4b44ULYQM1/NY9ntBpzwGSeuDB686312VHY4PTCkHFR8N6kLv1g06Ef+ph
W7/uEJx3Y3pCG+jUeYiVxy0dwEdUv1tqiWLfYqjahqXMONpV8ydTBSIeg6T8N3qU
0FNKIkW6eWo1rmpptGXS46wFCHSn39emDRU2PQF5fvk5Xp1FhXIyknNq74NmQM91
7aw+2gi5/TjRGnSjBv1E/oO+BaQ2QPc0FcBo5qpTSmBAEUOu3wjfLpjFidT7m609
A+lUMzuhlQP6B5m1oXhdPF5T2sMlJvmtdGMRiEDVDGbloAB/pZMhjTy3iZT9xYmX
klB4XO2nB/kV6r7fJ+F+GNtBpv+2E/jhJTSn5IHN5DymrJYxsqd/t+QcOvCmF11J
Ezlci1Q8pDHT2eAGfw0lGfgfTwyfrbGE0rFrHz4y++w1NQ7er9sElz2RfXyJqGVE
u8nBxyawgXc0u2Y/KJ7W+u+h3luSm0nV9kSCL/EUv/CRWbXsNNGCgxANu4rVitdS
JEHsmCqiR7n27Rp43AkTUXG2J+aKCbfesvP9OnlIIakXIDwZsG6v9UFP1VX5Atpy
jKPVGO2JFh4oFlWpVu4d6rYtWgunmPFQWPJUWiyDfZDVcdSWajRVJ2wURrGT/oRg
URJ4IO1+TgKQG9n2REtM+MgG+Th3p/u5DKhdcu42XNwNiplBpj97E5DMJrCIIaAY
iKSp16G58HU2xEDbXHYyw8ckgodttQDOA9bIcrahXZQHhtFiF69FnAt8IcHayHWe
lOeIAB0gksQo119wxni3cC5RjpUkIiumCgmhPGzS9cm3xEGI2zxrbBiqwPgNdRvZ
ODMRjIhXNHz+BcGN+j7oZtcx+sS2w7FEy97sRtdaXC6qH3cueVsHCFXBJeIowT2t
WS5d9khZfUhLzUFahcf7gcdTaVWQfoFsrMbXeHMC8lEoiuew8PAMaPwxQGFpnxxy
+U/frx7nfkVgPPTXkNoMhjVpSoL3e340bHhIxWuultM0GQmSMMWFvjTrFzAhGSRb
ICHk+GfOz2w0QXKyTB8JwLFqjP8KmW09rewXPRQYXLSo+P+UkFDtmJyOd4X9m+8R
H6ojhILgLVSX0RF2F/NiExDZD9z8mu6ogjx6S7+Qtu/fbch+h7uLVb1EeijC0mGu
vPfoqupCM2C1Ambk/U5jPCei5bMqep18eCtfXZybshbWGhKDcjqIwCkJlZf/fEKP
/DiIrFPTYnQMOr1xjSE8kKingJEhWJjOXk2YHdwxlPgm2a0SoQbSRfMAbHB+RD6U
P5Z8l9r8CiQHGGy/098wVd35so81imIxep291ppQlN3E5Q46y3cQ5uquzhgY2SSr
mzbnmP/jCoMYN9tQleVST9XJRFaIUQcCTWCig3Hl2HuX+rImkblOzFY+GX1zRJ6o
6TVEouzWytzypgi+WKdMwqNaBVkq4kGSodYdqUCx4o82BVR19dehCBiTOAC89wbl
eHjlFAaAgWiMiDJV3rJOEbjs160YS8N8L8lrzUhr92K+OsdAlt8eFL9dAFWZFBKf
plbh2gvGr4fc1Xo3VUKcEizkPfqca6Kbzq+GuIMSr1qELWntGW7rYv/m+S560qEu
5SjFj+nzjy+/CUOT0WSh9n2uE/7UwSpsnlO8NvD6vEqLGJCeHhchjv3n9R5NrH0C
bn8IGlOgII6dIv0qh6qjPvhusBZq2cQoTOlWncEK6MYG9BosrUZYYdE5LR7iF6RO
flYaKHhnCZ3JTrn6opfsQ7NnaQqPo5XnjOVebMS4H13J/QngolWB8IxVn9zrB4qv
O94jR0xYkhjcmGe0eEzKh9L6eftwaKpanLylKSojYRn+Iox2IYBLBpKQZo/5Nk3u
BqW/t8+Y2Mnsl1SduiXXzoLYh+jRN3cWXvdwSUxCyRNQguFnir+DHop6MMbk1Lwz
fU2HzhgE3nEqLbKMn62JMiXeqEVnOI+IlP28rGzob6TDqdTcIV9gdU6d39MAvPEx
TyzilRKrFtyg140vexNsjZQaftCsCBCXNQShHlxPY9Py5zujuW+0+maQaG5l/0rP
wwsQ/uqUX5Hc3V73Tg+Y5pXJiHylLcOTX2daJDo26dGvtv1qNBY6sbCC5hjjQnAc
IwDEANq7KJ0urLGJLAxPit8DQL639XJuaNeXTkTf2LBCdA2EC+IDym4wxGg2nEyA
vmGWaKusYRveR7xfgaF65XAUocgAQaMINl6ckJ3e6GzQyEnzTZF/cwFesQS6WWgg
y0xDpLeTf7+NHmUeVWbytC4ZEyXQW5/9spQdjGx9L21odysT20fccvGgNDh/3L+t
U2VniZbXgAEIXcdBrTKLPmEIX/9kV2sDLDlc+g/d7TIql6LKNY//8SH/KW72DR4j
mfgyLcIZujtdNXtKGMizLwZMhyUnfKoN00Iylej7smoABn5CmIQSyqax40XuEzAC
aRN69n7MwAtnjkW8vOgELCU78QVQd3m0hCAT+X62oCEjyv3w7CbSKbef7Jzt6gjM
eq7qo4BHw44uUd4fkyJdgPnapafW2f6X72O/hWpS0dIXLO6cMLmnBCa5xIXhQTcz
4fxM7phqaUSjs6NUPmFcxWR6IwZmjTy4/dYisriYm9Mb+9b8VAg5cXM7qchzMrgq
XIgTvXENsaXoB6gOf9B/qLQzb8GicP6CuQz8OMxQzvdlsHm7UU46JuC6VGACZed7
SNYMzfqW3jWJ5ckas8CBdA/SK8nzAnVLJkF4s2eQ6DHjqYqQchQcB42cUUqbGGOu
TR53ZP/aMpScq9JPjZWfbFHqYml81v2vbA0u+bRmCkeFtHjWd7oWBVRbmlNLDtXp
eordc5okdl65O0VtBjHZfzxWQfrkomplmsYD+MHWSlWKNhCJPpUkPh7GMgJMbgJf
77AWbu1ACilWYmUAvmne4+JRhq7tS+3L+rLfB1ubOsV9bNxvsX9O9EkEnWKwkWye
I6Z3bKoroK9H+A6UMhITBvAIQim2BHBwvG0jNgdat4LMmXTuEwwzAFTmP1HagEBt
g6A24eQSkGDjwUYDKZPViGZn0t4nSjqMqDrLNoHUj+XEMnGg/1L8anc/adig6XNs
hf28v5O2czvxact6dkOzbOtcJrvwmqIIWOnmkRDUYmw82P/s2vE7QbychZL0hJUU
F82/aysoqjRoCqAb2HSGJO3OH/ohLkZBmFhDfZHGYyEgYvjA4GNQE7ulrQapy5i8
LKWayki4cBUj/ySuwGYrefXosbmgf1HvoEoZ4vImoCvvdxuilrqByKMz8EsWdOOE
k8gtkIdHv7xiyYBVHlMZulZdYF4pcrX0tORXVQoH6qRIWOQPW/7TL6vx1Ya5EJAn
NyPJm9zMAj76ZQDLmbEOct0db5Obg6kkV8vjDGdF+f5Fd22v45koDSWWwyRfbQuw
EELGNdoaSE+fIrdrZ3Jp8W1qpJHsFzx05Q5fF8d+zawoM5fhVO9nQnGswe4+QPaX
ygHgH8Y7tp95IJpZK8drIV3ZS0+xOVf3/onp8zs5Ar252zulw4F/dEH6v5sPX76x
QarQnbl5rmPhVr9mxdcHiZA2QOB/5hpZirTDfo1p3mdlhhAJHtkZu2WBc2i9CWCY
7/yTezwNM+HOJ5PoXehiF4KII9iIYwPJ1sLGQx1yngO89EG1SyyferNwBEfE6zs5
yVB7T+iHwikHD4oB35X5I267Qh+JYgl9ydm4URpAz4wApSuxmC2xhsWy3o+oeh3d
vMKBvCgWmdq/xsYdzVGQTsAcXj6jWIMHpjbzTQ8PgNmVxEd8ymE5KmbUkoKg6EiB
I7I5cXHSxFYlA76nAVOhypDBx5nsht8aebNLguK9TQ0bH435AdRycaFXIKrKut0D
IPXao+4mgrBlXa+tINHeKMI8oW/MPPuz+UhRCHnBsWEYFRmbAvFRhEDH7gW98Ts+
AV426uhKLgkCt3TD4jvWB0trzoQCJWjbdxxMafuJ/eKpEugad8atv8iyGaRtQBp5
sw7foLPiQdn/3+E5wapyBFXhQX6gicMSQeeIV0MsW/r30TNOlOAOb5tX6pGYDmw/
WZfdOpDkXzvNu25E424edv+1EXOCiW9A5Mo4iv/Ja3e8T5rDR6xtvieyzQfs32sS
26TQYJt/89VXRd30YEa8/yUU5b3zxPw+MHyxrz4Y/DBYaEYtciXNdBevr0xL3GcF
cJmM7P5EkJKHUuEgcaXVvo5HaDHvmQtj7ZjUlZ51YW2dnOQOTfHXMo5yzNIUG5wp
fU5z2ZLchTGWl+0MJXLd/c9NJAKSLopV9+jlfVLIJD5NNq+fzBZP380rdzYfhesU
eUsPdQc0iergkQTwdVTxOurCSgMrzaGNm0d1f/k8tk2vx2SPWwblbmPaIz9qdegO
oBfqYRKXjenDl4ZvPrH/Xzec7bHL+GnhxhHRu59rtHogdLDef6uur4DEj9dPpFqy
nfGpmqc+IkefUhl68WPsQa+4knXiKpf+0Ekbtxfk9ILbNEskLH1b1WahihM/UnFu
wG/3aDdPB/pCXiw0GZvO+U1lWApBSpFv2HMMlsLuBNnt3mPVaID9DSKWU51CIaOz
dM50TgiRa20eUjA7Lu+N2L4DAgF2/vvaVL0S7D9jHKQD59ksGr/0jzmzokhC+qRv
r3k0CLKqtC4J08i1WDm8VULYFPQmzrTJl6rmuilcpCtXnm9zbRIHNSvviVVlE0wm
kLazsIUDc/DcZdzgBfGgmrsYg+TIn97mblSXFZdeaQpwkn1BQTJV4i54rglAKJuW
sYH7plx3GtIEfk8QFHFp29O4c7HC/7eS6k+HwIY9cVhh2jJ8xM6OXMfBsjqLqlQT
T/ltN+3q9xUGkd05SC1MQWQkbMywj/YB1Z8dti6s7X5iiAM3J1HVk3PC/xBC0Stf
5ZKV3lzzegzKYyP4F91ix4Y/tCtmCgGPcUhKkq7qbbgnR1vaLtbet0H/ETrbz+Wm
TTeziFtY8lBdm5qvwEqZ5eC35wD8i8ZvDNsvNjCgefOmoXWVoy0KhOjbHL6RHc1a
sZRyYwUpPVplnTMxyWNBYWduMa3HkUQy1fPnY7MB9IKnu9iWMBgOZDdi/PmmHpXf
rGEnKts85dvqw0r5GpuaRq+PL/nhGDnxJZQP/FMOX0hB/cPAci6ZzOh2z58RK7Vt
vLkXLAOSczmKh5OqlPrDgsMO7fhRFIw2JBGLsP547DrSjqNOjOPXqY8+Y6Q7atuW
6UCrmqOWtKAG5f1j4ItFL1k9r36ZvcNDdCWDWmdwIn8BIhePBCzsPQPKQGchcta/
aq2Bjsw8Tuln2qeZWOYNRXvobYz0HtTwHLYxeNRzYOFyHBHKt4CRQJjYJDfpgpcR
qiN6tI8L2Drr+JRR55fb6a1+edpUCiJk3JZzIIhZjuQnuSnbtz3ddwZqkUc/MbnT
l0JK4KUU2upj++0OECHKJI6DRcXji7Es6gecm4GUsewrhEqOM1oXyIMfhHa115xo
2Pe6+e1klmHTI4d4s3q5cp6B5fro2sQVl1iF3Q7jZMSVP68L2uj6h7xt8MXROYJV
2a1GT469aV1Hes015aw8HRfYd7JqOVCVZZ/TPFslHpETwRRVzb4ioyXhWoL6nrhy
Qf8Jaw82Gq1aJWZ13rXEqSnJjA/QBPfSfJhAAA5uJY1YfXeKPhoNoOJsQTuVFqsl
PyQpcCX2BmoD93dtG+Zl23pJL3r6Si65f2mWGnbRhOlNN87Tmlog/BFL2jcz0f/p
avF4Cwbx7+4HiDfpgFQDh9IE15VoYhkb651I5EWDqQaV3lKZjlh1URr90pGIGiyT
OmlaSBAY04gQRXE/DK2BdxOrgPgxDpt45WE5tB8vTJdWX+4PictqtqgLbKqZgXZ+
dXb3KPdtzlvcHg7OHwhD4jd8FpLsrDev//jHrDCqPUROfiHy7sKw9iaU1E92hV2f
06lIa1AwGxBU7NclKmvMOvHn6AqRF9BG9xjO+PysRCYpd7ott3SVGzSIhVdaSoAY
qBk8IiAAUYD7lQAeA2++EyuHmdvolKLibFyGdc05M3b/j8WhUbU86fWBC2eCUVV5
IuYpGfmRUAP7j8vgmqAjcokY1TudJFhAWAEcykrbde4hTNHnFWicwGFGq8IOLW3h
XhmuCGkhK+DoWDFUBLVwUWFSo17X/UF/ABVr75rrx9l5hLwwUhQPO32WdwB6BYmT
va1ADQ3VEL4SWC2y2N9HgwJ69a5o1vDQrYjbq852O4nT5D1aHiz2Ttz5HeLD+3zs
t1ZasZs39sishYjmgtXWxfUwfLcH6q6RfRBXOkGiUshlA4CVr0SB/T/BTIgX2ZRz
oNOSHzUZ8VtPwe0T3zye9WyTpDy9UqQNQJgmqIm8DuN9qlNZpkk7kE0YNDrFvAi4
Juc3pbCVDU53dN8f4YmcdoxTOlbSfyjPJA4lICDxnkm1fGzdpcU5xYI1ufa14HMv
1CeDfF32wyL/GnViJx5tGcfd1WLydCHcHhvqX9E5O1d+Gtaqsrv5+mTensvEtXaG
9ydtUGPY8dEts+X+fPVk/q0m/BW24UzconyI2M4Ia6q3nbqNNl0GXGg8/2PhQWMg
ZyLgsPLZdvmqLZxXmSZyM0yAf+N7hoLg/ZIDJr8A5lj1KwLy0Jw6XN/QMbXDugcM
HaMCYPu+hT06COxVyjJJ7bUR/4P155qbiBUd0HHamzIoSUG1mDxxf7ZlA8/vgDLi
PrP6VHunXhBCt9OSHUaA/Even1mTOw7yMfGtgASlzgZfIvc0Vxd6y4BiauhZHu6Z
bXg/a1HL2kxb4nFCLR4qeeAhEi9U8EkmLYxIWo4O5W6mPJ7KVF6Iq2sBbxvUtPVh
qKvQfFEeDPa16+QGP4dmYB4ILrFYJQJMG+rW6bFHW3pRkvoYdbnhyEQ2lEa0Zsro
hHdJFfDnHWQKb/kxkvtykDDf/UtHXgkeBPDjP7dH+oQr7BEQtso+1MY67QgSg1Hz
330/QMmNin4GSl/Dvw65F4trIvduIlUQg6um39aESMeKbtxjVqKAUVRH2HcXMA2Y
ArV+cutogfu1n2Gmf7sgSL6tPmxkv6Y96QUDqkZESGA/W5lRVjdbyFUi0wOqthpg
ePJpI4jEzsyZXea6/0m+GFkQvEBiH8vQPIZgMsLGzEsnQequNylVf34WffxdcPJ4
4ArCg6TAnaLJCo8EU/3uHzJHx3m4Ez8yk79aPCdwh0VtHMjOXedidJzdq1SEBVWV
ZtiLolw5la7xuAY87EbPySP9a5KfxLkcIdf/nps5tRM+5lgMVCKiMCfJrvXoxwpk
ZmvxH6FEFrEymGL4TwUoN8FOHc++xmslWW1rMq1jYVDs9ZedCiFiJRzPcyHhTauW
DZ7tK+ZdXEHTV67zpshj6j2nslqRWwRj3+neNAJO5cg12igH9i8GAraj9xsRqiIc
7QBqafh5lNk5QI4KjuyNA4dzegD5LUTpdx2F4aGTZkI5seXEgO6IVY6PLaz/4z1Z
paB4EOXvobEkojM9ROwgcey0/uC+ZBULBjHnc3C97iMIjsKBYKKWT4UqZnLrppbK
c8AZlpQuAFgBEdq9Ei+O+3GXaf9ZpxFxVNzX6M+5/IIger3ly2hZkXAH4JB+y4W1
nucGCErHKRhT2mnC4zR9OntB/XvcxqFj9OIicxH8ZA3Ox6YZ6XMQJMMgnNWzTbIT
bJO65M1PRJ+TyqwhoV4A+D52FYglbckYbeLQZDfa+dxY0JEzRplrlLKfOrqYCki8
o1xA5aHA1iwct9xqWNai3NSg8ViJWo3wLdkH4q2APQQqwknaEEbN2l0vE9m34jep
9brVJy+Fp4VHPWeaGOpiDwIEG2MhoAlVX6uF9WSC8yxjdRoCCqAfzzj5cuPI9wjI
stBUcpdvHxWy1YAp6jRD+Ja7eb1onx+rEgqk1NW2wd68EnXQB7+I6JGC30aO1taX
VAHF23bFcAC79knHSntG8R3Jti20gxcYg+V3HkCM5lbpf6v4EaiVFMvkvjeqi3+i
cHoYkZgJEQgLwAaFqo7GlK8SCukiDR/oGT0hksYy3Rc3pxO6qJgE9kX5yTCHSe0g
/IkAB3IU2T+IgCObJ5//N3qh1pK6a3jAL4clup2Nr4u7VKzqC7zMcgRqqqi+iGdh
/j6/2eRr+FdSySI+vEElCD61RKE3NtKhAzVmEGPSKzV0VrjKbWRNb/PwL6jQXDRU
iEyPbbkxQgJ9LqwZ0Ury7sWH6RIiS9vCiLIpQVlWkHogws4YZUE9K1B3UCNvorXp
OYAvBeXkoOAUv++HBcnAvrTejAF6tAMkYSvRKQV6Y4gDAK/eL8iX2hTWDCH98QlQ
Eg9jeMXqc6AK1TmDeI+PtxZfPi5pHASe5PtPpuuMSWnm9MBvYOFjak1im9xKe5aG
LQ6g+TETNHFNtAA/AEhJMisKdGgzC19JmGo9bvkAoxzrL/9sZvv7m873c/WsNAoB
W5Dd6i//OsLhkGF3UWSGKAmb0QWP2mTetzB4QgA+nHoCBUe61mFJZsJBBju5D5dO
W2FkrEgaFXR7a98jvsYvlXtnmDiixYm9GI7mlARlGx9b3NbYYHVSTUyJoxqbrzQw
55WXrH2VCPQ9ig9ODczNvZvp6hSetF08vaOu1i0YFWXrEy/90zpOf+zq/RL5mR+/
xuWTRVlLVl/I6HTcP37IYKedjhZJ6OAiERFH4WPgd9LXFiA8F0x7CSUxXrxGfivK
Z0aaoMNI3AQieSfLsBeBBWLRQF9GXKQFgNUEh8KO3kTXdyhIeiIQe8Fk5Qb8sO/j
3Lr/GDu5UKIvz+qp3xfXtwak05DtYQ1Xcctc2qRnkwk7TRsCuas5BATfZPcpbkol
ugB58cUJKpUBpE1nO1ZsTMyR920mfW61Yr5uSKOtj0oe+Y5Ujqg1WcyGhoEpm6bY
lL9io6Q2HAVaglEcMr3sjuUKUE5V+yZGMtSR/9jpl8edoij5vlQLp5kFvej35irc
zVWJN3x5i8DWtVge8Uxi5gQU8DEU5fnP+M8udAy96+vyMFWf4MVg47lS41XV9ktu
A7bD8s52ebqrWkKZW675KY0sfQPfw0X8hVi1SxLWbpJZlm//hLK1TFasXZN9+Q0G
yIRqEQDwDmqzCpWHEZjLbHtOAJURHcADMGy8BMucDe3lhHi0D0+i7BiM/KuAWW4v
8T4oxSMIjW/Et+o1Y7WzyIsVNAjVWlI2WXGZTpi72WSwmmu8p4pBt57CX8U466gh
4vZOIggDQvNjeoKgkth1sLl0P1CcGuRr+6WHP9jSgbpDGWSG/zwSeEwODClIgwzD
3mMP7Ei4qRslW7e95utGNayKYIgW2LNHzUe+hO/9CeAB9nme2TKVzrqXX6e9wMWc
v6Kiw9wg8f7xrjdXXyoDFMB4ExEtPoD718dQMlc7muhOyHMS+SdRiR9HaI5yYhgn
/6Z3KK75kzg381IW/cEGvlkY6sH4ATPcikxESkT1Tl0aw97BY6thGY4xzetc8wVm
IjpgvKXRqYXAR+o+n1rNKjKyGXg1UKzdIVV1MW6OCsCT6LtIXmg/5aBvaUy/exSD
mzXqYWRR8Yei12nnzuUjiQhkg74BzyT56F7cCxyCm8zA9sJszwoyooGPm+jwCvw4
6frQ9EJXBcGR/NzepC1mG8EjJDpizPxI39DYqZQX4jLIs1aKBL1BOpBFAelAMZ6Y
9KQlmMw+vqam5A4igSRJFefwwmDyAMUIkKU+O0+X/1UnqXMbcvlpr6oFyLarQ16R
wbO7d+2u+JB4D9WrshR8SXVk+kpp2QgU1cEBXIf9hmPrhyOAxuTV+HQqbyTsHF0t
97kVABc5Rsu9Y9ubzxASlXpxzLCX7CzAu5HCqZvEd+YdGemCdfXxPmuiAGoip0Db
UTJ5s1V39SJ+bMzyCAFPV0Ys9tJL4C2YAv2TPtguEwPjOOkhqbakjYjYcTU1hUgy
52I0YclCslgUBpSNaQgt2hUM7JMW5BbudaeoA42tzRS2LDbpj3Du5dMCMuXcwYyB
/7UaSrn8zxu11rtEaFoO3CNhyQaM9WlT9aWA2ydXA9ygHsttS/2raCrZpr1g+m2b
SFvw6QvR3T4TX/q2wlFzjtoEsV5xcyODzPf/49qBTcy3mEF1HRE0+GTDPHATOmFd
VtEXvwCQeDAVBa/sRb1k/7r+U6nzjSGMGX3RrRvBaAwY6ei4VHEjnH8BxYcJJUaQ
escfL1y8pzsBf2lQc6vr6gHfZKd++YsSDkFMrCkgIagzE+nAEasDvg0Po560bzCZ
djGE0QJGUeDHaQ6EnGNdgkjonZM1p/TTJ78PGuqEGC9mVJal+E4xxtQ3k6zWfS6k
vNhGnqgfI5bk0VvaAsguXWL8/nifv7h7sqj0AGLZTUHH5B1VGWgNX8k3Or91CRM5
OcoO2OC6Kwi8cHc/2Jzval0NIr0+lf4qm0+QTm6UdX0qYYd+FstRatwvAaeKikEr
Y7fpnmJ64fMA5BZYJgtF8y2OJVQHYn+LnfeK9oWtlKY1PZoIk5AIUs1QsGhsKM9q
Q7TXwy6PeHrET2mSi9nE0vGxJ79at5xmQtx9Wd2OAlxNRvIJvrJD2aGhXBJFg5ah
J/RvHaJLaR0L6EJomLPfU5IHOtewQ1f2Z8sZk1z5AZzxB9mSilMpHafB+IT/+7Is
DYfeXPXjOY/vZVagREDh42+pJGBIMkdeVqyLfyObZ1YpTW5XAs+0hceBWg53omY2
yVHewsNB+9ETQhdnveKhdqOvX76w6QuxlgugS5FnUz3FBae/UvXAaEy87wHOpDbh
2rSdIomrSVCDEMPti10GtrtzQarcxMoM3XfKSpWl/FXeJKz60QxkwBF1RIP73buE
Bs+If4CVu39FsW/EbZvD4phxCD+joyBIaoHVm2RI+z4lSCW5bmgcsF3f07b1qHIc
P68f0qgXl83H8Nu0XS5WRQZC67FrG/OGMRGITBgw+ADJv306B9JyQEqlIKCWGFXm
8+493MV0MMUsinFBmY6Hc1lN9lbGbn8jNBjklLYBeuPIfs+n6HAfw3KStrd+yFYW
T1zz1H7b0fiJkuDrOwcgUZNl3XQpSnvuHeL1fDjeCoucKzYJjB+9pgZLinColJf5
XPzLcvyJOwj1h4bV/CG+6GjRztZfCHhUMH5Kj1CRdOWynKQbNRfFtibp/w+MErX/
yGEL+lz0R/IzB2w07KINEQYwh6FQP63HylNCzhGkH2lmn1+N4RbTFUapa4U+ZZ30
htfwwqd+mVkBnydRO9O+MXrddvTmDTKkj7HSARJCTAlFuCxUHEp4uJ+OEHNfJEbQ
ablyI/1IXXuRogLKfSGaQQ7yvDxcaV8P+I+Tp7OQM6LAXyBVMpt+iAi3jFY/2/3v
FqDmqx4GD93cySifUzmkwOXGHbYbjcGzMuUZ9KNadCroFZTPZVO23RAkSiECBPUp
7cZAYgwFRlkTs5jnvEHAHEXqRcYdU/zYQKhe6utdsm1F7b1pERaagdS1ymk4LIY7
0gMp5T6Mv0+nb6QTw14GsmJ6fSk27fg92AgxQIWWQrEtstPpIX3vt0sfHcioLxAp
pFkLTfWurnh8/wuiz9ON6qSqFuAiOqmlfCUrXMLE66MDivaZDrzihbx1pbpBSRQt
OnMfyrJrMj+zJ0Lg1HtnIRO8klyBbSPuWyUGZyX5pHkZlHEUspIKPlNd3UVeVPej
0xmQF54ugXepu1scGWH/TEjcNkDZ1z09G+NGlmgWSbwwcd4+XUqP5B9FI/z7t5xw
kc0BlF+SuGU2yHpg6fBypH2rn62MsP1lgX8vSfrtgRKmiM/0EwE/Kd/xutqW1m7/
2RYZwOD3+L5okG9XD69JpEeK+DOWjsWFc6KdJc4Q9dTkp7iqelkZyhIY18FPAG2b
hfDr6IPOPeTIggcT2azndEqm7vH08X2nz7GccKbx4blOA004AP6Seob91Gu+4G35
UUJp1hoc7R6dO0Dp+2E1uDOLU//1Ya7rPigojp0SRZAoupZE2cQsou8rm6uBv3nB
rI6otHV0W+YId6gllytBZSEa3kZtt3B284h2HAhMLVxFG6xkN+8dN3bcQyNjHRUi
cLVPDHvfDAKaPfeeSZL2xZ/7sKf7zcUs0QD9s/xnX/6vb24g/rX3br2T8VW/xhok
YNz2mZRvw4g0mK8+7UdwUpd1DMN6LuiT5KV87l4iYYx+IxNY6sSXlVo+Oz60Cf8F
RgksYUTEpU8TK52b+MxFfHOlEm+hVos/OC30LiNoNgnk0qKKXP/yqkWC0ixCDEGI
QRuN9VeVDJsCpwY9kmkdFU6m0kroUzEhsKJeTilmXFl3pDjKNcVy7d+nk7Q/0h+n
/sW1+Vz1QBuhSMzLIhhr8BnmEsLHiKRVnti3X+7xzinJQ7NulvJyfKp8V1nJfsIy
vvtAtOL8ExOciojkjDhwC1xvRSyb/d8MX3AcQi/LYcMxYrjK/YGWQOngRW9EAAHZ
zFZxPVQ5lP26p/9oWZ3PuG2aRPVBTpg1pttD5hkqx+4lzY+eqtEamogS4tU7RwqA
eC5Rrs8rbNHyGuDp5nwv7IeEaC9iR0Ya64QYehQk+LCMOKdE4EA6JTL4vo4iksgi
k4d7O1TxbOBw/QL7HCnYo4uGQjzDTVisQ38YcApBh0L9LSEiX7m5vk/ScI9kKBv1
gi+dIPR/7kmDtFMjRN047SKJi+lS5ISlkTwWajLLYX9PALtaed+lXwHSrsdcdXcC
UDbKvCdFQyI4HwQcMtlRqKzgazRyPclWg3EV1wUlPVv3q3eR9cBGbbzkXqPGfKXt
ki2zUiOGINU2VhX9HHLTO7r2PVoh92Lrr0HzR4TO+e0x0JX+ddQU6R77xVpEvHeP
ZlgXRn77WtCsNFN/+lvTAXuuoPkxNl4F78ruHwV1M4xQ73zlT+eLlAhMr0YXp+9c
L99fyODPke5gJvW5lchoKdhD9AYcL9lOqohLxJehH1tNjXliyOtl5z+3VSmVStAS
gDQN/8Zd/DVj6nbG6g8hI1b4WbC9JgQaD5IMkuApqLx45QrOgwARXVEBSVIEn/uc
23+Bi4ptqJRhETsyA5Kdm/URT7MtU6ywIe0i/wVgBfx8YuKOFtJB5dmcZKsx/Nqq
Owknfz88V9iZqOR8NLULp1L5RRQGVfRFy/+wUsGxpvP8hD58viRLvKOCyvXRxj3x
xyqpp/Liq8rFU6RPGuojRQUGx7mp9EIBSkKuq/pdnepMTvAwmHsarJNJUoVihDBS
F7JNxCjJEgq4tq3DsngG6eqc8PvrrEkBJraVuOodJ1wzg3yxBMvKKXmtthlvZYEf
iiQJyoePanz8svujgleZISgyZsUsWKa2PkTCdIS0V9i5fpjZIjeP6Iai6QrFZyAg
xf8a8RRIPPduJFaDW7zZyKKf7D5BNCdoDke8sIBz8SISf2Mpfzn7mZiHtiu3qaHm
ZW311qCpmlK0RAZO73bSTli1u7ej0mnVnkO+7zKFB5RkgDBBofTLl8qq7BB4nC7q
utxv6kisbrAIChsK44U0CNQNOHdlRUT7HCPJfzr/AO9WLydcuDhvh2lXXUovWH1E
xxNU9h6zC+MH96tFmsOMOqJUVZs/e5DRFCbsWXoCkLG0KlqiiN/mcYNUycAx0E4O
aB8DpTgwSQ+KI7N3bxoLPywcCNYbgOB2Ztv8BzpwNRCXecBS5d7715eRa2V6jH/w
4x/Cb2NFuUpxmJMDCEdUVDcaftlDn+dzsyr7SJh5VJN4as5uRKl7dcWpVnHtbcV5
m9K5ngb6WAxit+BSCBVSxUotCKJfavbt3BTAvXhs9Vzfw39NPGbXwjV34DNR8mk3
DW19gSjjPi9aLr+xHFCm5E7jHo99q9O2ljavKGmWVocOy1bbnZjndoPLUrUS8kKS
YtEjeGvy/AakWOkx3LntICw4FkUsf1/kbhgoOpVohZ52vdcMK8dSeJlsid1zAlh8
DVWXJOQMHkU6VhErh6yvEtFtzYa+yhAuCJ7/C3U0YEdSH55xWO3efUczN2iGJCTS
g2GjU30yf9ZE+jarwfhmcwBdVT/rid3WagBfuTROCeQ7cKbe1q47mdUEOthCzuLl
CPlAazuHayailupo1kNL5CN5cIIUNo+JHnr7q4zLBXHp85BLjdbrHQwHUJnbmagh
Y2w7acddn2Q75ThEy93u0kowBqSHGmAD9nqiO/BX8rNNBjO3KYgN4Zrs9WOhV9Yy
8SrpN/VqIxHhqo27/TJ810njiT9ZJVQnN3mSgQt4Sxr/0OiNnN4K2j4bos7TCkO7
35tF70Ndjl9Yqxz4KSkPOqE1bt9QTLE4y+EyxEEq2kRxf6Ye7B4HMu/WKZZrDfoX
+y7PYQ1ZXZmPgZoKL9egJ5/yODpHbiosZo8q8RljpkRxKSjSbN1NW2rbL+DUVLc5
uDOlroTMTXamLRZ7FxS8li9rrMByWQkXmtfRVRJYyC/V6f5m97BPHYkOXWjlaVbC
DY2Wpqon5NVd1I/VWikm8Ijty3WUWJDSRS8yAWbvhOH9yAXatnTLm9zQHWV9ZQMh
GQZsykXNPDRy1GHnBwUfXzQtHwMGMDLwK+PCrhl9i8SRe/6UT2blGAFFcGPYoYe9
6e1pAulnWZMgycE3DSr9QRX5uXNQtwz7znBFh42OfDQwVZFqEPbxkjVp/GFh5PHw
hBs1qYTB+H8qqKt8i+TUh9v4cksaIsyQcL/2SeJ5YiB1mld3TldTF3AmyvzLD2gM
mfJQ9iZsJ8zGU+5rRC2a6VaLEt41hoSxFcc4PjDjMZmVB5e0nRHcuSLWF+7/okDY
gPV0ZKGW7h8x1NZQfICkPDXlT73FY3YObjGoqXZO5+d6yjP6BT2nY/verPcl+QKi
cwqHbDIvhNos5ngdnc9Jy/eLP6fGDB0UypPTHncwga4kRjDzzUfxAaAX7YFNN37X
nMtD8LVQZ4M2cuu+15BKj8Ik5nHHal7zDK3tdF6Aoc51iyBlgQqwOp+oNZNwPbWs
QDFgPn61SGcb1VhZbNuagAZKlR9wo6XiOQrU/AVZuhFF4YNgUWD/9OickuzAh6dn
6nQZFY0EE6JeWyX5Cq7ZOzMCKtuOWFY3ywnHqcQriWpxf/rDmmfYDGPPzmFFEbz2
CmIWn2u+48MAPn4mq+byygmS9hluCpqamLNif7AOiSAy3YwO7DshCr7lbpNT8s94
NARLAvi7UElMpa9uVTz2lRqzkvB4/IVQC8ofdlqrcncgxGzAz7rggEqY6ngrMI1s
kxAS1XtcEucXIsp88robzLesmk5dUTUzf8Z6pqzWjgdwTEd+WVi6ISOOXY+iB3J1
20B7GtH75jE+bYMq9PSaj+jlFIi+hApSGRevCevkm7nacapm+7uHjzMQazAFC3JH
jJitojNDzA8SZMRudBEbPKsZ8XTKSzmbY/+BrCo5R+z5llfImqrXiHvxXUyntXPy
AevjYeXjmgxYLkuQ4chSIE8U5c+sphRzr+TDChssJzQE7V/2YrAjr11RNWrMzDv1
zDUXSzRu96HDH/p6xSTaXb9/skU1caekgI2rwUT/GqNqYDB+lMcCSdK8A+HPSgxE
ZH+wd+1eK4QUDhcS1WBop2FSk05+Oh+CTJ7/7M3K4rUNAf24MrYrLckhLJ22+/XP
ST8YyTsGHlkIaIORUY2+dG1tGW0M0PkOYprhTtpEQwn39vH8hDOZfaziehpghfcD
RVJWJHhGeNdwVAOXJKWQMGOTtznWKfdm0j4QmNMsDQgbi+NTOYOKzrP8aQ0wg3H5
bNiFMRXIOcgRV0SbHx6TG4gX0PLGcQKrwPcw/77jntQFECDKQotiEgSdJNbS2l/B
ER1T6TCM30Mf6ohmSufsCBs5TMWxUNmM7PQbD3fCxzlpPHATdX2MCSVcJ9TGeukt
EZViXEU99jz+vj0Cbg4okRYsYuHU0ksN3wZyImnfsczpYku0Yg1bnhvO6HjDHe8c
2HqtK6sgsJ7oIz2J9CZZI6UJ21jyQF+x602H+fRmmhBdoaxivektpMt4GpYwOBEP
Vs6e/y9kJPVw6CectTrwwBNsBf0tanj5qpdlan47an5ryzwWyAc2AOv+BpF3CnK7
d9KMoYFP39MDaU4WuCGE7SMABOQPp1A9xePkGP5BM6pWOf7nZkWgu53rCwNZiAFV
Q8S5lyFQle/BmZTYmYXsZTDLiisJL1DMKdB2R26GgAP4xky1vj261SqA1iGZGCB/
qLDwAtehRUeowVhUPDfKFpMFG20ikmod4uuksb/P0Rwdr93J+9ftsqUlmVjTHCTt
cWd9N0Qu06Q4FrbDV2kdOPC+LR7w1tWi9o5neg7ox15eJp+1abF76Khvgk8Cr6/x
QzOfE8RubUHIXWN8MSc9ncuxrhXqDZ3fIpHySyUQLxQEmTCL4YrxPV+JQyasxOKV
bLTGIBota+BCGXgMiYvc+PmrQuvIeYHVl/BWxXQ8HcFSUn+x5TrOt1Fsw8vcJ0qK
AhRzfbPrpy0BwrmyMLT0MH8iq8h/FDaupAIp7XCq2obpbz2P4nhmOoDXB8Zm/gvl
63MceVmsfmkjPiDHmiSxa//H1PXR9brbDZjAczrClqqumPeYlAuccS5ls3HvzWH6
1RuwBuyz/peGN/ygWFH7rLkXdOvUl1RKqoel3e481ycTqTsB+tPlRv9vnSfvBzX4
cUpk9mO9Mry1mJJC3g9aiXpuRlikRRW4xV0p8NAHFEmFOEJJ7Hzc+kydpsp/VPfv
oTbdYE7Rm/W/+zu07068H3h2qO2d1auv/aR22X4OvAG+C4VcG1nt5QWgtyKKQDU+
BuPUG7WDXTS53IEOinraSFxJg/9W84tJZx+3L11RHGTV3/0HHqhT2v2b17IWVOJq
SgtPT0yZUe5aTFgQ/Mw5yg8clVwYBnLkSkJzIG/gRC9PynuOYmIyySSA2svapm41
+yftjaJcxNHcaq1O6z3qkxMjHhvunESq5W0uzUNM6vN93E3rw0I0SjYfBx5FChwg
GxxYFU51h8/V4Lbnt8K1bTPSsFjAL1Ie01N9uwsS86KbjewOEfLSN76BnvV74kl6
48OAEsSgtzcHT2uSRz45TNSD3MRBC3HkYlA/rwVJKoiXjcn9w4R8v+aDpFlf8qk7
ZYhPsN+jcuQjruCI8PqK+XM07gnsh32wrpQ8+NUGHhQ0QOpxYbw5A5o47020TK31
ovykW2q1Ep9wBootkrMhlH7GqnKqX5vtjLnyBUBEX1NvaK6yJY/8ah3KGkl/m/wM
cI3vcc1k0yHT7MdA1eLg58kBVTc69ILLzxW5rMONbHhernvUaH3r0PeQKEC0yvK7
7C7qB8o8lMjrTcPy/5+pgidXOfBfBfht2Ax/aFQ0+09YCZTnv6MUj3AEWAKWFT4O
Qd9zn9FLZRQ4l1edXr6mnA1to9Eu9D6zy8dDSl2IDxwScd7qfnjGeHnc7/lX5Fem
prBcU0f+pH4gAEEp4iR3Uff1TNeflplHZb3oJ/vLkBx2wJY3fBAvyZLCXs94jEMt
1ls9DD4ssfX8c42zIzWSkClhtlQa/2ntmiMCd0l4i3Lx8DNqxEiJN9eVklYNNnZS
IFrp3/3q7u/Z5/oZcdLtioxbw+b7euRLRzmUJzyLYcvXBGzLdELbuAryn8RQnFEl
268SmnnZRKWIX9hzdS697Zam38kf2w1dgicBAwcFzpKt7BbibKsSCUoEylmFs2yv
6WHE+RwO4PWA4tUz7yUEi2GGUl6BVkECs/6AnEY8tEvAiLKeRDvknegP7jf+p5RE
ktHvwYo/jEeQxgm8kuXfwqwcVKPTvrlz3ZQovwrwSEOxKRIylRqRpJV8IMt0/9CG
5BeCENVd+QlAAb7ckkxOHzZ48I8v2kpGvf1aUbSzg5of5No5hQBO8c3Aae7jzVUS
HeBchjMStAA3wdyGvOIst8qMdM9SWRd6dREoiP3B3dV0cSdsHLGCGamuuTGQ07yz
FdmNDdUGzyNgr+aao/S3PmiGnqltc9aIKvYslr5RTxjTpl5SGYrHfEBQ4R5JV/vq
JvV3GlvYtLekzwmmx65HNuXDt4qh7HH5lLO7SjstFVskA1LQgpCYs0Xf4av6jN5J
hOuNPyheOAZnSTeDRiqnhG/OQNh9sfFQ2Qm4hwQS17utewkQGdnZBCWdz30SiUXo
21UiPeCM2zsBLIe/jHS2uduIhxK6ALqA06lQZLOz6BdTHqbRYB0QNPcRUV5SDAEi
qb4ZmVGwmszHRHWxtms5aJ3Ixgfywtc07gDcWrcnvHOLKLW8s3joY5iRTHdtUCHz
gIyQwo9QX1n7zMvxVoAFjDdeRmEkriBsiJ0eJmXgDnLwtRIZRL/QQY4eOflN0yI1
7m0XSOJZXzRW1K5OMs1MV1LZszGFRQ6nVWhy8S0i+Tly27Bu5j2wTb+pP3miSkhy
sFtmy546J5i1Z27ziN/uFsU8Qdcu8SLfa/kQ38rWVD/V10GX+32XxTEb6A+d1MSp
dLTgqjq2lHAZCKX5I/UpVSexWESGfV4SILF2Hdm1anhqyB2FkPdPMHoIob4I+YUQ
+QEUsLY5H/L3bo0QScXW39MwNN9n1FJCDuhNZnXcHy1k3SNsc0i/+tcc0tkVPij6
WdwO7DeizuW+U06vwsWyqRtGwqo1dHtcIQ213WXuV0ieXEY291Po4R9kXyhGmZ+Y
PhhGY4Juoojzp6OLMlaKSrndkOQd9RpvhcKcc1b2oA1EtHDV+yqn9UMUfiXY5JkJ
zyciF5ep/3Zg18A0DBnjiw64/0ztjq5BnRvoNIsQgfYpmbuIcM9N5EPBalIHB5Qc
JpFtHIwbVoYA3865VJ5AysGrHu3KLEr8XGN6DXVHNxesWxHDDGPwzUc25PLd2aQL
0RDwrPRDMDAjd+cytmsVFXTw3oID1gBCYvU0usPh4tQ0J8jrcfNYpBNfFt6yjMPY
RxVkGRV97PHw246X/oOkL7LXI4YwL28G+k2eEbJHZRB7unYniwwGeBzHX9CkGj9m
KOmpOqoRKtAIk6VNy3BVWPF0HILeGfwvIM3/cNvURxnMj00RlTlOte1H40kDCTnN
Dsn9GABv9VS90WmLB1VBKv9Ivmp7V38Rl31sos8bNTKzRbAeeAkTED3d2PkTNCJJ
M9/R/jsKKAYBOqGhxPp5ufbzqbxPaYDijG0KZQOjdz/a0nUu48zHSxEAqjPEHens
9X3Z525kh9tyJlR2p2NZNgFJi6ffyrvMPrthyWgtzM3/7MbG3YiV1zINsOKtZub5
1oz/PPV0owKks0Q5/qRczvo0JB9DnZAGAcs4Io6DJ6cbyCwLSXFa7B9SI3dU9WQJ
R73+r95Z/01isTnyEapORmGDF3oz1RvyPu2nvV61+/sKJnIJiyO3vCizTuDHBSe3
xJmpsTqobBIOYQi2ylJfo6t2lvMoqywnlZc/+Wt7coUtGHNeDCwv9GesiDADI+kH
v5vH1stJRzcunMrQsxXW4RKD+PujT5YWJQNCnTRu2ndffySJhmvQ2clTWveW+D9p
G2gREEAPTkPqZ6bIJewLjYSDe4FFvmfU6i42aTVVGV9ZD3ASRUOpvjTztAD4RPTO
Ec9VncSAGnA1/rWE00YV6C6Gcvtg5hhfaq5UOACW+BrKSDt8gIhyeivc4T/sUAqa
mYv0HgrE4GR2l5pXmIkB4an62BWy35FNQJ9Er19UAaA+77TEvw2MIpvzJe+Z1KAl
1kJUM20TQ1w+GHUDA0FFc6wlSq8wmr9v3T8aBhkeN8rKcYzGasJoV9Wcz25rsuR5
QJbMXZ6agYvmnc5j0NuNJeV6Z+Lgb8P+6XLCx6OYVOvq9wbyFYlTBtbZDa9KIXRj
vqkO9PInGpWHWJ2t1Pf/xWvvv4U37ex4rtGN95Es28TyARw0Se6wEMBbC6EhxKwX
/jo3woUusp9q9EB7b8r2pRwgpCRuevGCHGV62vnjvPHw7+26AMBAafSPj/jo5JEs
Mn/RdgRHhMWXxcGKS47wyeqekBb8roYmx2TWLHuvvAm8QWVVKg/GouA3WWvma/2/
A+VvAvZy67NW0XBRcWlGFxMZGjHwQ/JY/yCyzqHmhutDY5gf5Du6s1BAijYNp1b6
btc6pKDAJfgE97YVdYfuaMr7SFvZa4x/dXBTAW1787tKQouToiAGe/3lQu5y4wQ/
Qk6tS+ZbW0rbvRyW5Wee53OAYKV6OAsQRsrj006mDcRHYnUzonk+G4KTkF3lqgf/
tilQIWpQrUMxTTWX6oNScq9hbGV5AA23L/hqm7bRqn03iH8RTtbzYBUYiYdDpGz3
I5VojB8iuYXsc4w4ab0voA8d1WMiXAey2lDVhItstEQ0bFh3h40bCNHOinB2Zi69
rVMh7pqvv7t6TwbuSjI9Fwf2zkA1BoX0Le/paABFFCzSpapTPgn71k/3Cnwzq5d/
c3645aPI+fncJfU33wkXPh+MsYZ232LIyBznHllwMQlXzwQgU7x0E9Jobzhv1F8R
NiwhmHf5mptpYyalxAtz/ER0MNT9nJl/k2vGDsKqv/i6taUWgQnO0xBV0WVQ/X+Q
XTvb+1d80CHSksdHq1xkfCvGc3R6noEg0svad4oMYqMHnXG2T45tY7vs6f7Vkku7
cXjmWE953zQ3lg9XjG0q5CMKWPe/gBDglN7Vum7k4c1ADJokqQa/D7ykokw1Zspe
xdMN4MM/SzNVEg2xVWwuqrBJHfRZ52hW5nA1TKWPNDXrhmITaxShbJ5x6t4huCZ8
gcRxW+Tpy/kS4Rsbfq2O06r48ijF2grKwHxu3K+IkyYlS5THw9ZYhC+d38fh3Wzx
G2OfLErmqEuXQu6W2l4gS/l72INu7G+q4OW3Cfw259m59HhdPnnRmG/QKWfOfvtJ
wtvH9/zeGSBDvg5pLYGTzi3o7q+BgMco8S9gqHUtnC907fZNoTPoT89l0OiFZ1tl
bQKzV/1yNJ9dQl3ysX/U52pC0KXiluyUqPQXrAAJDOtsVSV05pvuoOxau/Xk9Y9M
tdsfxIFvk3PWY0hxDP6fxHpzQbUlNrtp8Ew6HzrgysFESAXrRhuYFB9ts0kVFzEz
/adJOk6ioIAj8LBvRj8uGjzUzs1hvVFJd6T20tWY0qZLKLDOmvJxr9t3GkcgqI5b
N/CUz2FApmhm+B0US9AV1CeYy/X6shuvWoCXVPjZP1STgeAugP4RtggrruCTa9ES
3xhzsoOrnKtqBdjDBqDNEQOsqOb1ZwlNOwXo8pZpAaJ4t+I4UrF784eRNMkw9I49
z0vAZOXM8YiZMJ/W2/10nEOvI1zYBmFixemX2dNOo7uWrXNsjA5R/D2Q+3FmmxNW
+ou5SkTqdfdxcnPAuQJ9FeX2sQ6Z6Iw65hrQgm7ZpRAqKqaP+vF8JZUFMJ8ioR2A
cvH3Z4PrHLOugQc7ZyYvCndSucMZSWWKeYh9wsGDmpFEN7E9zcYglSO+EEHfh0cy
eD9apLoCw+rWwZ+Evc0la9KzZVXYAxyqffd0If9X3JrA9KttfOyeNj6W02wOexB2
bxvkBvT7ggPlgpoiqL4WV5HtK4Oqy35o8JQOXRqNmY3o5oewZvDkFYnGuLL9Clv0
QSCJdFMuw4EqK/+VZdGbBWzkRm1rV2z3R7xXD4rZi02A5bHNL6szaSnDBzROkv7J
L7gxW9FQRxk5aaDaELUcq3xfbw8wYaYJD87lbaIlUdGxxv5nDcv9J60d3jkKi3cx
K4cKQ3ERyqa2vpne4h16EIjof6MA3p+YN1KgJnvSXImV6aJYz7lr7qYz2/LHjVh+
zYT/3ScXeLC0m6eZxr1776Au6ug0NhpATf78MlMFEXV6ZRooW2MrlV5WYTVTulmd
jQGWshMaclvj8R2ncwJfTN3FRcKE5cnx3V3hKnl7DjgUKlvdQWSQrc+ZXLqENit2
G+9o/9uIKPCzb5Ycs/4GsD/b8l/vp8V6kUm31ZQnQXrLWkWsKcK8J3i0tT7ItM/s
KqjLDKFhl7GEQp9wk8ypPTndG83qjFaQMumqtF83nJsy27K3OGZIdeeMdFL9o+Sv
sFRDO6l46VrBmeoUypSXq2uBD/QZpWC7ISy2WYMSeNJplLLkuJ1FA25qwFHOZ/ZG
DTkspVNbpvIgp1SVFIc8xyi3uMxDAssEbQt5tibkx/J1HhVvH0Nd7Gkl5lfq0AwG
Yd8Wb+KkNebpfimKaWU9o6X8t6Se6U6VhVqHE1Sv3aFQ2QNOBueIKzKJGQBMqwSf
bYNd+Gt96z2c+6SsCl4m77lqYiaq3Pn+mm57E5SESuIbOaCgoYwnO8tT8mpEdnwe
KQ6xf+l7Zpex5MavULIwfPgYQd2PuKzKiCX4kUpV7O84oy9hGtecEp5ca3t5gL9M
SWFVeqiFFBz/3qonW+f6A7Y/AQJ/BC5jTNaW+UbFlAGt7zTqCutehNi/tViRchbh
k8lcYeYQh4okIA8Eqz+JugqYXlXonQXTpAaZUCx4OxhseiOlmggUPTCEzulAkFM+
Ic+rD6ecamRC6M/kuzKMHJfFpDp6sozBHHLudHxCibOyAMufqTydd9Vylm7ccMC4
aN1LJqAnIf+gqqy6PtLXjl077Y+5PJKIlw9h/hCzJfl+WIFqQ+IJYAG4CLI32zbh
z7NdPxmAhfjPop+ib1FtOgS1sY8DisaTy2lvMQgA2AO6cj0Yk1iMfs6aCcLSvlc1
fETq9b4mj2mY5W/7BtYeujxMqzzbApBeUuLLjK9H2tw4UZQ+F5RiPs+0QROiFdKG
fEckadowWz5MbDDxg9S//fPSIfb99n/C295y0zT6REaTbdTy3dNOMn8Htx4uk9rg
jT6P8PKc0qdeOIUUlqZyV33zNZpeYr5CgDvfEU2JS2MXX2xx/OWk8iwjBA6c5fIl
tAAv8KzXGHANJJLD6g43ae4WYUqn22ElUPQVMA5DJSz5ayn5UvFoB06Ga1Fk1s8h
SxsK83E5cLWg0DlO5mUNc0CvYq0iCBlJqHRXoRAUPo1uFrJMebICe/BMBDMXOXxg
cjVCU0GDvs+bBBMAoSuODAou+DFUzJG2PxXR+1BobgFNwPebe6Damfgo9UZD4TUw
ZxGYPLmW2ec35yr2IXnLeS+GQTsIQFPNnBeIgdXBmA13sZhok0R8i3vUiAshpkoI
/8SHR4Yr7cuUkr8fDgWv3LFAyboh9ztvYbsHh5hAZEKjnErW33MGJLjmDEMbjEVU
4A2RG/Zoca2LQXe3JNGvcjWNYZ9YOe6IGofYy0uhHWF4LjmTvVh2lo6c5ttL7CgE
/TGUbKBf/JqB1YTS/xrnV2KvetXFObKGTNXTS2OJ9MC1W+r+FHPW5FB/f+Rgbyvo
hczdrfhRGuMNDbEpvWDfyM0xV8OuGtl25jlVAD3Uz6ngPdl9wLPltLGuCN+kxY2I
+wmgRBUPIaBmcBy/Ytri0JjeMmJGrsLGP4eaZbco6EVDzgBDwglUz8oF6ICAYfAk
jbaAT+EWerSoY5EQHh1zwsvVrHjm5JmBoVTPWn1sGscvo2CLntuOQDLibzano8Vi
urh/foC8PNG2SjnL9Sv3IWm3lMxXxM3s2SzvQDvuIcIXdQbSQ5dqJqqO3ZbrYR9S
/TJx/ygM/PdhGJoTXvDJB64k6h8akXxJ+pW2qljxqQFInK56OVrUcXpmDqWubTc+
IyaTGILvFS2NczkJ7K+dhQj2hqo9fodohrRX5blHz71ZRu/4xF2xrzZv9GBigZBS
YslCUl6vmBKe6X58jiUSjrg61zmb+4UvCoLc5xVlpfSp4ryEfZNRiCmuoBZyBBPo
lZolPhBqxX2M05I9D5qjNDxAkX5iTVBwHdWuvonOcYYz6aac5FmBDLm9J9NczvSp
DoW2WwG4yb9iPvla9wJUlsrLtbfdJ794TJYyRo06A7KkYMh1nKwq3J3fgiB5a+hN
Fb/G/Me1nRX4pVw6h7wayXSKImwnyZ7SoDUAab+wza1tg9oPZGwdBt6iuoGEG0nz
WZgAMI4oyC0hG/hPGKJXyYLvWXSQrx9+1ze63H9E/TK2xXdGpSVCa2789gNT6MwR
bCbiWJ2BjJyVtmbfMkTxfilsOIaPDjSbaWl+aXiZKPCDK9AQIfZ4U3XCo/uy0lCw
fvSrg9+oDbfG+TGCS4VrB3eqV1P3SvN0ooe/IOnPDkQN3C1OoqmOmouypVBg8ETV
PS+1HSJqbeA0Pcz91XKHzwfR3A8Qu3PKjGjc8M+14lTHPJTDpjGyCkwHjFCklWpu
hT4zfKbFMncxT+5266KVYCRsdc9U3iq8gG/7R0dgaa+pelcnLZdGPa3U+nbopQqU
bIoPDovCGappAynODTXqfuzPc2cN+uR9o49xZ+mVuzrrkEKkbwLQm3EgcTmmSlWF
dWnm+GsarTRRDI6I59dDj9fOK7/Tzq+UPJmkRFmEdWt49jk1GaLRQDrG2YNJwkU8
5MUjHV7T4uu+zXlnHZS44RQJA+4v39F/MVTpL7ByXkejPNeO1y0NgsZECZyjUOu+
OT6d/q5eCTdJBUwufCcXCKeoCZQY4IbMoZQAcippj4eSXq3ZvtaP119CWBSY4uv6
m70O8BS7sXv6W1uFHSmCGQoRH8pB+lExYbnI489fizrq9IzIa54knPDTB2J2FtVk
ALPIFdhSII9uzRN0bksTqvfQeMvrSxonCAULZhXnh6ugJtMTOOxkudWnsQ/xgtyj
N1Jv14/4LdmXcs6FPB+8ZLu6YXiWoQ0jpJKZTlYej2L4Jc5uKuaV8QWGhbhAymbd
OHhL78OJw8D68XwfUFjmzKEkmksNlcgcgRQ2YuNkG7VKOAw+FjEkQuHGkzWc/Raa
nmL6bDmDgGLnxED6ejsdxgqifkAPKAV/jbO9WrdIrK5ITaikVGCgHceABIb6iciD
TPP9Aoh0JsBQpqh/cADj4StxsBKRQLmZUksihgQcmal4trhjrpc4LRoCW0wLFLmk
MJmqYmFuY/wssiqm3Vqdm05bzuiiCHv15NuV1Ygraxe8TW1voYY68aXZ/+lVZykV
19MiIiqAu4R0K2JWcBQj6J5/cog0gsYWFsWn2Cfm41qKscZxUNl4cOz/5GVlUiNp
jFDzPT4iGBmPLYLv0fsWAfz2ljtvOojwdGNWY99oHldBpaMiuBLEz40d88BZklXS
OyDUKTCD+PzU8To9hemcl77gY1nLwBxceQcXWhSE+FftI28azFOwuozCdEny+uFa
l/F4D+5Nxginogo5MBeH7ONu1lI/kIZjdIJqm7iGnjcMXm1z/bexVEOjT3wRAulK
9qUoCnTPqZIy9gIwqG+GDymJ1qrBssu++P8Jek+qmig3H+KQ/890RgS6TNbm3e2L
H5N9+64s2ZG4LyWYHMORwlC5Z666mXpuc2Lj+Ihv2CzEjvWMLdMtH0MKknQd3Gxu
rVIQJRgSf5oz54JkxZaAaFJvePkx9fI4XKIkP7EUH4RAN/jP5+wyLzFc+K9UXKT2
pMRaVJZ6PefbSj7Q3IJd0NUDgd8BdFEYxQKpjfVwFJdg2IfFV+AFNvBoe0aOMfYt
0zN4571bOShjAXzL6F4jcUu0YxEBloPHaUHfzRAcfSmMXQuNlczB7p3uXRWtzHBz
nLTqNylI9rS8bx2ItMqzhYPt6y6g0/PBKjcYKcFo+vlx7oAB95es1cIFKA5y9lde
jYDZo1sxD/3HE3Hiaft/Zjg3+MRK80If4PMxpY0R4gRRC02goPb+MAqzA+KiZbFS
DqfP92PAVivedNFZOymQr1dt99ST+YOQszIB9TtA6ZuFLdYP2Tybh/2ly6n/9my9
5W+L+GppkVIcJkzMgtKTo7H9KwLj2nOU19SfkFDUCZ/RpoEZ1IV8llQ9K6n7a7Am
I/M9oMtYDUasSCKSnWZB4PKFz0cgtwi8ec1jtD8rdaY72B5ZHe88hTL199DkPpjR
0kLN37NPYhQqZe7WvHVBOKA7QbvLjYXzcA5a6g5Z9mTRCOfkwJqS5oHFtORi+Dbp
Jc8jm1XiC+sLmrYoWpZ3oN5vYosnYJTFmfz8NroUJjpOZIfiargtWD8prpT2phKI
GxUgw98bwKhYkyAtjGMBOc/FRiOblDakdi8o+w1l0m6Ks0jpbbeBxm547naQgiMz
12Ef4FlcMJigJYahPflKI5wLCnCHR/OWrp68FD4FiQq0arLe+iEyxwHIv71fU5qh
np4Uov2ev4I61+AQO/PvYsd3JDFyQcIvHLftuzGTmpv9Hirj+R6r57qfkPyqkrfD
X6g5SyIno/Z5KH+ymmtFJ+Xz040D/SjtTJH/yMDEvljWYArQb+wT5bOi/jwNw3K6
CmfQrnqgiiPht9cbQqb/+kBqX2SF0jE/HuJ+2Rj6DiJa2RlIPgsQDD+7O9wGEXxe
UjkCwAjzkMwZOzefqM+7QvXKnS2tsD4RBzUSLgHfoMSov4dROq004Oq44nqVBnzX
4TvuqFFQuX9VCoDCZ/XnT1AINVc1thYkURb1urZSqQLkyiNw7G7RUxj3U2T0VxXC
GNFnI0aai//0iLsq8C2+qYNUdsv8UU3pSwzcxQZY3XCXvo44V9sbuAvcv2t/TKaM
4sWpY84pMzWI9GmpSr8N2b2eCJBQVHJz17i9/+N0Rt8frujIKEjGuxaEA0yPfaT6
MKUljoMicuOJO1Sgcwo3Nj2MbwIacu1dmCQo24bmquSuy8z3GwX87zxfYJ6KgZh0
Mm3SE8eUduBt7jFCoA1xlh5TKH5Qfq77ZpYhqnu/mSz12j3Mls4MFgcnhAQFgshe
I61xLezx9h95VXFcd6jDZU/RnVsvCNLWssbacSSed2WLFnLVxAm5Bj8WTiGcBzfw
ptdkTtHxt5q60QMXmmsGI1RGvYRnY+Zd4zVZP2jgpPrKL6tcel2SHavdNGqkCqNl
w8tBWnpNlDXPxvdJOwp0oGdXJkmAcF/QpziUnF/wFF9ERJXzYtZDKwaeyCUwoYFo
xCCapLroIp0EB+nb+DxID+iBUZmFDrpBwUooqWKG95nTiL/G12rs0t+OybLQQdjn
bYakIbnd/zN31+XwO5Ppwwg6qa4vI5aRSX4aeMDEgtSGCiAqQCJ0P9MvxhHMY+pZ
fDFEIX8DKJ4Y7g1tM59F3tbm0WiZcnPik/XrZ7oyhpCqFBT3Xj6Pwn8I0HDoj0o3
/MxCbzLEDuRdoLPf3Afw4bPBT4GC4uEDuyt+CZw6flhksFkw0TPkZFbLqIargnh7
0AsCr3gt5Vhn/di/VJGSbyB64VXZDgS6lbgi9eNJgkymQO292koVwfnPUlw52cZk
U+vUpbfuA/CmdTT8wEJLSytRHHEJxdbQHrJ7BzLt0r4hfG4kaoX8prWYimm67gPd
jw499XEsM4mnF/NOCMqhM6PRZCXB0nKlxo+NgpoH9XL363QobsLMHqIv3sBrxLJ9
3osl+R2mTUwsX9rZqyG6cC1a4R0TNfXUovwiZHtn2gPyd7jY58jxEyooHoEPlK+t
SOgNSig0u5LsWEggWw9SI+BflHtt3Pzq0P3xfjoyQdgKQDOjhe+Cz4gM/TtJM7FK
uVlBmuVP/DbL/sp4YTAkkByQYq/SLAVHaYh3hL3Hrh82I3J+BdJy37RdqSwlvTqE
A18bpaa+zGf8mO0KUV5pXLYxdkpT1Sy189ESdhOnM6JInAR2aTG+YmoM0UpQ7RSC
1nzUGESfIb0h8eSKzYagugMLqbVZgVgV5HDU9pqDkwxz7TmgcZ5ui1q3kPrhRlYr
RBZSzCRmmSot4i1FrUXe6n+NyfXf5tvzZo2Hf128ca9ss26BFcf319GUrxeFcrLt
CUrtJpJUgzizRcYBcwTv8sH3V+GIq1RFt56caaPxC1UP3Fi/gKWiNgiOJAbzVPO3
nirloBoCC45kG8RNAFbJP06pxl8HHckRmG9JxcEHVfyOrKcnheCpa4h3xSdYJOl/
jqRa1rrzEFlcgid2voVHxtjJMhgsSPF/5uBg5LwUM5pTtbr8DPMiDgETFjpuX1dV
9yetjW2+OwKWQ2LOBB1Ul+UWrNRR3kS4tFbhbhhzMsnNqIYGCsVIH1sz6cwAQ43y
7Qy8H6W0nFL1TU3iOpBn+pjUQWRg21UelaoAN34E19X4E0Rtt9PE+g0jY9chTmm2
PK1zxmScUN8iz/YSwO7h1ylDZbrxRfLX3SN2lKAtRWiwKX3e6UBEaBVhotnqPzI2
PAtgcPRQLLTN+nUw2Se8KhxxCR0bTo2mUOli1qjjdU3392REHj3I5FnrXEpTLpPl
fg2Aenxe7l7VxFWg5ZK+2K3vMIU+FOKDfD1NrorX2NLYGWo6QJWcWQsT4WYyEAML
czYAz/6inFG9ym4GQn/8h4prilu52P8Ggf+S2B6wK2e/fUFwS41kDqvdt8WJIlY0
kkpN+KCxd/Sq0vR9cbHA7EXpkGTXVTkBbFoqYVy3joSKmgZQR+3/VspyQl0AHisP
o9otmcBpXEEfqZ60tk/IW58m1HZCJcM7lhleANjQGymExmSuC1C8+8TAMEWXYqBP
4I0FOkynkcOWFpGh6OP9jf9o/hz0FedZ5/Wr9x5eNVdi9AhLoD36o7ZeoFoPliIv
6ZnuEl/nkR2GJGGiJ2RhkgHA/FSxP0GJACyLBtxghiY4/nLteO+k2RGiNU3rJHEk
Uu8EfcUNw4WRxn4OIt6oG5TRciqhKYvx8KE5babg2W4+cHZ24Ni1oUr2S6OziVuc
6q+7ob1HPmGP2DpR668RCpNvmlwm99m53txQ6UXdHw+VelSWJMDpalCuow4siXa2
2x9JpyBtxDq0mwwrGa0/01GkLSwazzRgt6kY7lflp3vImWS+LYrKLdl4VYkpY2Bh
nKOqgw05h9CY6Xfkbzs8DUMAioe43qD0YYEn31V68l8zbzpTYevCFcKbcnHt4kLc
Yk3NArBSKmmdBVKbm4ZPqCeDa9iAyWAmB3hlAkf8J5/BlS6+v78tUmRS/lDwwUjr
zkctdN1+rloJaRRhGnRAIXSnBQJJ6k681t1hq6FfNfzdObtsRin7CTXEHbDLgTb5
jmPmSA0Aeh7AxZIe4OxK7XPCg1ppWufc5rrO51xBwd6PnhFF8fSp4LeKEseoT5ea
WpLSGOwGzl+WyLQZ4CsL00oWMyBgFsB4dKjO9YuQ/alXDNVEYV394svoDFQ+1zNC
fHeE7W8haw54jrYi1h/raZc+ANXkfmzWOIO7qqxt2O+M/rnu+GE2QGMUHPkBeRZ0
DxSf689GLxMHORuxt9+mq1QI/PTHiuVa+hMskX/gdTxAvd+Aqw9z+YQLySmUqVNN
CFaEd0Xo/6C3FudpsXHdE0WWFKVCGzkTOOuG/0/PJwjaZK301lOdlNqohsgm1P/j
vc743OVoN1nHlHWNmAjYXDpP9FpKsqogqXjn5RzLlXEdiflQrbEBPl/o0E9J+Sku
pL6aqSIAl4CmyETeYdcFlSox4MXkciYUGzkT2Qs0yAjVlm2Q2EnEQ3Eh54ZRiagn
newVp3iJExeJ5Yo1LOg2HJ2DzhsbugmtAYHCDbUz5TGhMoFoDRyZeS809+BDiFE5
HCXPIze2a24QUGwVOOosjqj2LdSW1O3BEg7/bfO40VekOpm2nAHmffGxcddrP7HF
Y+jH3acsva0nSz2OcL/p/X/T/Wgj4NmyyOWqJbj1W0hpVBwi6ZtpTe1fIQlMK59N
koXOcjDcpBez/Vd74b/VtcqLS7mXTAJAQtpBM1QKxASVmYeFGZ6JTstjP2d++WBF
2XOmpyb1eRhCHWabK0R5lmqZDgQWMfaizGN3AtiM5qvq0lPdgiRERNe1DFyDQm8S
Z0kfkJM2G6MVapAZy0aefgSP6JeQq8MoVgjddGoIPUI/9MjjxPVb2+dm13DYnaYD
9tdF0USQlBNNfiosya/RT5G7qmOKrCv1S4+lm/2/Sk83IEF3Cm6hH0AbDRSbT0cQ
Ffk+p0KhP44rnO8U/cyanQ3bvUDKs7cn52+wz7O5p4Qzw27FwjOFTtVe9ve3Z9wS
c/9MlhEVTm+SlwEsw/gHJqERIB25ZKOBmOULYOVCWpt9iNXPUp0o/C+45icKayVF
pCCwD+qOaSubzSFn08sm6m5WAfsyJBrrbO93e5Heybq/jqE4mNKMYo3wUzQ+VxXe
0fjcpot62mcF7/uEfRoj73R5tQKudWMHC1XHAgMopamjWVGH0e5S/i6UHT40mWQo
jPgRizpAPUZgmZz5EVHKvv6RUalRzpcP325TYwbMAO8fHXSa3fORQy7DkWmFmmxP
aMtXl+D+miOCgVVLpSB9aEIf+Q7goYvoRU8h9QOlpBbSrIKZEqXCT/hs9n0LSSPC
XtcxDWkzscAY7ZWl0zFcwXNotLCC25SMp9N5hSdoDNs59wbkXCA8Oyg6TfBwIpCe
QUsfmWTFT6fcCkw8dVuR8W/94/WcnyeIncp9Lo037BSwDBCcesTlDFL3NXkmVJ3E
o4MoFMHnH+V9wu+eMxySuqO/7IZDth2tkSSARrC43yMdtc79pZDBojw3MGxKCd5P
NorC2UqsQEDChsGh6eaOMueuazynk5MQH3jr5uClidLwxlHn156dK4zv+aSpGGYe
FF5+Z8P2FbqbCnTjLiqc05kBV5wht0umGG+DksE8qMK/2MeU+7USn03cpiglIVdh
tUhLGNmZuhquBiJn5YovBigPWvQUzJe7I3qeloJ9XXmiTn78aEAWxwGZYmvOfIDX
DdxvlT+Twb3cxrQJCwKlWRA5VpdY7a2SWbMbAl7qxRk0d/mIaOU3Ghdxxscl1enW
OA/xmij8qVsH10xNlKphXdw3gMm7zV2VxA28MUFKiGw0Lb6Q2ycV6TBhCVupqulx
zxORrmrAu2KYK4HF3deX2qJ767xmc/YF8HMawNTvKFu2SZvBt11PO14jvy5U/wwS
7ynpRZy0NsVvxweShrNfgk1ylc/8A0UdoN5mJg3BX5+B4ZpOCyHaI9dgVc5ry/fS
icb+/9GfDz7w1ijX0y3vY08TISrZNw4y04OolGoUDMj4zhlC4gigad8TkFSVDlm9
Flflyo4E9wTml5El7hS1uKT5OcRniVcswgC4OoxYHe69WaaFQJshqReqfd8l0gCA
2TZmCJhzGB/JFU/g3kiK6CD6iymMhAS9kgXSTokQZGOmauDffrbaRgY3AzdnFHM0
gg+E/cTbVVf0m9ccU+Iaw2tLjd9ndh1pWjqnvzQZgJFJPmPn8f4BNOAU/ffN68eE
QyR+/rxL70etCcyy1uLOQXWtBO6VDbVVtDoTcAiQAL+XcMiShdJ5AD3DVSosvF9n
Kj6T0xMKsPNbGTKfDFxiA+XjFAQz23xC283vCbVaoqItiJHH4IYiiOjylOjPnzo6
t9BzgNnmZoJvLD1WMcLk9UhqZldwLOQxicbCd4nB/3WHmKANzYLeCnLu9j4DlUZ0
kwPLDMBu8JCF8wA6lk93KMGFRnV6pU7rrIA67jJzPHcHR1eOJjGxo8yTnXagGPpH
HfYiVmAl3NfA+qMcsKWSX13y/EqafNjfVL6OgDxqGLvowsVBCnZdOTKJEDamJwMo
159CTYg8ra1H5D2hbdeVvkOgYIkiC+/7PH2K9PFhh+aw1YH5iUGkf4mDkppuK/nA
FCLdshiNh5U6/wuohsYs5zTJ9GG9cUixKbX3b0RMiBQxlZSmvuV6IeNV4qRllzN8
GicAw6q9EE2yOGEzK3+N2fuAMOswN9TfNulhqAx3qzIqF5pmIrCHO05XYn/5u6Lk
jW84vkQd3b31yetnU5r3C0gVlzEBzo9/0+n6a0BGFZ3adZX4Zxt9VbWsxRJCz/gk
rsnEpNP4w9BtxkKGtB6MaUIupc/8IBNBJnx65ahtyM3/A+Y56iFWHMVJKWQYmrBD
oMxUwt9fem4kNW5lk+9h1si32zsdTmQEFZgHaDGfxI557oadybC6gt+ctGt1doxn
2z5e7j3p/biwhNiErDnYKcsH+sS7MVByDkASVgX3VLedNiFUqmjB61I5OC6GNqEN
z/ljwMhV0jbscqUapq+0nrNHOo443OAVzyI3dR5JOid3akIAH3l+JAEGXkVGl59n
i93cgtZ8nnJ8Cf6qzH4uA4tzZGjtm2SKSDcdLNnCxSWayp5j8zcNfqvF7iY4MkA2
7D5Py0OqAAFYN96nLOj7ejFboOUv4XAEgs5PAEp85mluGptglCPDH2Sde+C7nAlJ
1jG/6WdDF0yXQnfFMI1o8xQT4+huYpFQRzCbx6hMyeR6HLLR2/U1bF9Fzq7xMnWJ
iIHIjaLPG8YPu2OAHR+ei34VaoZrPn39oAoe5ePIaHdzExrX5mrdCtKUSIb//Aiu
XolJdEQcjhyrizSs6JphmZNE/wmPo+wsp1KAtzXt0Lb9QckL8uE8fvc6zCBuflip
ISR7tLeajTULZYhetpGIMcYws5QnL6lSRtEaWbQ8UtP/Wz8LqSivrrYQouyRURMh
lLhhqwDfI/IIJcn2xYv9FzrlGIJhtJLfWFBf8Wo0Q3eMzqQrqvqQeVKsgBHQhhXH
pG7DwEfQy6+2D7m3b3FlnEzVEB9ST+S0ACZHGSFrXpHCEF0659Q03oH/lMtl7Yyy
oXCDx+xzeiY3XsNNPe1jEOONgOHDrnFrjRDiTD00uVL9KQOSkMr9L0zYrEPn9AEW
ljSHHZ1YUwftUj5lSYdUXJBSqM4VPZ1X71xSi7Uxsdy1q8d//iaL1r6bw35JOoK3
tXi9cWTxaLGKGt/2gFEh8ROlLIdSXaDNEmFKQjSWgiB6IrZTJYbfz3h7jrdODmL0
iOtxejq+iXF9EWEfggBoMMUol+RfT1eFxu4evQQ8w3OgudPfB6WGnN7pe1lcKcti
YWaHy2Udo+7V8LA8AQ50V+5P+G90ygbsPUL8JC1HoXsoxTh+w7JMECjA8Qz0nyJp
wxCt3cJQFV1Kx13v34OzGUbSieTMYuQdqkSM0qGFirKbylXl7RzU0xzP9f5GKgvx
X9W5J0aSSlHMt9DgSuqitEbYq35NILSRUIeUYwzZ+FtU/ocO1LCZc/IMY51TK6HN
noxDzxw4Xoqu2ZUJy4XvTTqcqqcqhX9Fkwokb5csKAKIDB8N2A8WygZ46gBZSIFL
Srjfx2ysTByx0XIsJMv3Av20PQHYPbkaM1WqyRDt9BudVI6li+kA3m0K0LAuCtrS
Z3U735iBAmnEy9NWJUpnyZTifF7lf3z85m6RF1rllcxM6StZuo1xIXX7eeYwNe+f
TcH36hdK2YEoyMES92guTpGajozhN6bKScFx+SFCgEmM0GtUIk4w7W1vQoPl0el9
4/wv+u6nd/m7bwD7Cd8mnAjDGiGGkuCZdNq3z3Zv+uD7X2URjjJTxWulXvLOZMLp
gvLeDGTUnUcSc1V0ov/3ApZL3GleKRSSkG4y/+SKLaoKae3gleOPwVJKq+NgwTIz
NSt4GqDvVT5YRl3W0tmVPcyUqQ+PuCj+Q7b7dUliYh/K6e1OEr02l5O/X9emiPgw
iRpAEd3tuS1kpvc69161ybvINaRHfZoegjm4nvHsqUGdCqdZeRs8Un6yp+xX/kGu
CcPs4JCyXCTBKXIucFPR8+5UMG3l7lSzbSGqq3jExej3z1/T+dFtMJWHYUnEldnX
qZZvsIbDRc714yKkEsVzrkUWftjcmuE5ra/BwVIXbz191894G5t+88tSWAshshE9
rajnaUhLjdG2TIXxzAgwKnYlUzOy11Hjz+zH4L9xuR2cIRA+04Flr7snMi4Avg8g
vKWHot6HOXdJVJ3iLM49ObNc9ZGewyrWremmVWetAikCHqhhEQHw8c/fmeUUnPba
+t+pMgrSrh4xTrIseTrH7CyzkFDVcX3un2h7wWsL4KX6pO/+FE9Ao262l30EjJEp
y+IBZEMfB6IuCEZ9XWMuKGPVvKkqXAcOzUpZ1kLBvqmKxo1TaRHawNaP8sn/bXSY
xsnTE0COTpoDGapXKltqQVhMkmmP/twKv0ObkgVoDGzZc6oYSSC48d3oFME2NYy9
wmO23P3qht2C4NWz2SHIi4icznK4r7SoB0w/D+OBREvEX78quctItAenQVHnL2bP
FQ0CbpZEsw463jz11EeYZVituMKtPPkmgNoRzBZlHdvyCngOUNlbPDSxf/r2UKFV
clerwXcbgiLANYfWbvDdemlUF1kF9/iuHwxUmy6EFKKvkGHWnpjUFh0HHAdUmZRb
7hjd3WQEiraZsPMEbqZLpnf4LCy6adOcw0PhKJDAsZXKdehssTrbRTZkEVGDzhn2
amhNzFezT/usbh97+8cpjSeSVGqzQJ5sfx/j4XDXBq50YekwPtXFZDoEZwA/R3ds
mg8b6KogYGrpa/NYmehJ8eu3huqtXAe5Ah64YaOJu77ynhYkWMrTDJ16blxSCXPV
u83Bn+K3hCZ1nAbQ5Qmz5qb2qzq3+iF/1ctLVvV63Zr+MKND6WgduhBfD0Cl5EWB
eI+o3qBH/ql0+jsO7227meJctC9/8vGU3oz7raRaHn8wy9xjWGZfdS2E0VpmJuKt
ldSGUd6Tir5n/062qCXw9eDECB5/+7JxjciZ91td7FDYlSuU41JWxM7Lk/U7FaId
1saUIxQ9lRX9hUlcXfT5eRVp3baDMTEFZVRm92ahf8hUKjZ3JDJIQ3eynaNPQ/HP
l7CVar06wh6dKXjwAR6/JnH0vcc4lzWyYofUJvNUndXbhpQdpsaBd1t0NKEJ9GSj
IQgXIFTwC/T5dJYXVVTR0rVzz3rTWuacc3GjU6dCi4M2smAbdvdQSrB6lr4oi7GM
gXeXXS6gKUBNqgponeEYN7fk4igYFyRhlQoEe3ti5FISbXFmi0qIYEh3fFDc0lq3
4N0mm/n6u5i6xswYITm0ilNj9RV4dMMISd/xsz3yBbMaLq/xVasgAzfR8G1WWzkE
NnMbgIwpAXqA9HNFELloKCFmpfXSwZ8597NWISDiASAzvovzQWWZb0WXQ+BeQksV
GFLCJfrTmxzmfetPxvBq/24aG+vEldUnQDaegMj7uwamrWZBb/LShnDXZ3o5gR8r
T023iNMgY3h89TI02kquNW2MFplGiXjUcWthBvMHvpCsarB5ANAD4lWz/DKCmwPv
6DH4UYH/5v/iSvDW3w3yCc+gXEpLO6zRM8QtoPiGfClkGeC0XIPv3wJWKb89rd0l
e5JZY4TtiDk8xA5RRByvFylaBc5kcgul5lI1j+yCHJ6aTPY/+WWcRri2wLjPQPcA
5Flx2o3LZESMTtiPOF76PZ5su6TB+jzNfiEMTatAplauy3Q20zzuaCmBnJr/mAL4
f2NE3VGD7vv3QWCDBR+7GYgORGOfs1B7lXWjzX5sH+5+LGaCkGMLicXB3Gi81YuK
AkEYOs2yWZXF0sMo/bcV/otDnrpQvJIBULw09yiLbl/eBPeMkYW8ritr7K74lSR+
2E7eMjbCOw23ZPLVExlOV9tEP6ry0KXcmfXQS/RGq2PZjlb++Z+YFYSx+Y1jP9XP
mb2/n74fA1aEiAOzEu/CmSE7xCCq9mqTQ2rSMUa97/doV8DLr36JRlO4O6/3yN50
dJPMCJdSUWxbLuGrHyVvgpaY60vTg6uuHa4rTIm9RXLEJ0HiGgTTazc2x9IDd1XL
nsQ2awQmFTNXmqSKPLm17B5ipxkeWelamrZpcdB9YWNY8uK92eN8kJWkZC9M0CRP
j8XdFGjszuLaZQHt/FqA/K4jF6H5CmeR9QKniCCilyva+zvfV+ZIHFGaS7g4mQPo
ppltfCmdwq5sKsclqsoaQn/WFVTI+pgvzeTsfl+MMnuNNYYw0Nk4sg5cDVSe3nBO
BJE0eYp66zD6PU8gO50s42QYO812iGqtvFlHlcE3XLb84DccU7cUz3hi5x4dXDD2
AGD8NKAhgOWkydmnvMSFuvDBJsMjzt1u2Uq6neBdpfxEQSbfWXs4raNJLP7VZ1Zx
MV1zhKwDiwsoSoyXNZdNdp4jNEoqqp5wchcNk8KsKr2XzJkWkci5/nbVnUubbfvH
RX6vXxWQeKCYBkBiZv0gEjckZyuIulrPnwCNrkGWkpcWo1kG9s9I549CpG/1XY6K
/Gr0A6eCnriDJkT7G66ZFdWme4mPjonsGL8IqWn0jED5a+GlS496lVhzn96ecW2P
XWO84op0PIXxSuDu30M4SUQteDVob/9OsDUYSu3bFbsKuR7smKDsEty5uVtDrqlj
J8iq36LNYB9V81laI5bzCrXbFpPDiAPey8e/yoiPBS8IQDgtGwA3sCCFI4uB5G7v
ZwEX/pQ1AJl/ND1gDBnsYKdhDcH1Oo2pGS25fSVIKd44yXNkMHkZ1Lp5MYXAD6h/
AU4jWCTZ4bQK+gt7NY4YGGPJIScyVAc2fDHAQNP1IqESRd/GcXTUy+V/P1UZ7bsF
HMUHMTP8wqGoFdqKAP/0+XnI6VwEzFb0pR9pPCgcyXN1qXnBCxviq6Z219r8/sb7
xOSPT00xIURIfkQfvZJciZQwIwGLubA1rH84TZzykuSw/zXXNKmTcguB0uKAW7Ec
3Jggi6E6yR4+nUDNqs1KsAMTWY5/Z58ApZAJweFB5emRzG7Rqz0UTpZxU4XB1yiQ
KEiKHMIPkT/fMfMsQkR76l2Q1rLIcRnSNFzSlt0gBdeGvvQajfeXblYxlzobOldk
vomksAsoixNvGhIkaFn6UMPTkeSlg/90gQkqIZWnZrfuHcvKDtz7Rk7R2svzmyYA
jeHEKHNzbVm6T1qvOlH+7O1cer0zvt5DnysOEGiL3jWC5xT9mioeqDYOOOFCsnvE
2r1yKJ6GAMH8dR0zhtzDNdE0jCUPNMxqQ3MHuod3WbzE+ozNuPs+IyKaobJiiGYF
heMpj2MoZ4tuSFFECKF2k9Q4Mg7Vo26YZ354bUhz8fU98MYLnURrvCmz/L8eeZ3+
dahy29ZoaR7eso+JRZqcyOanXmdo1F8LsnotLaa5YAg1+D/gImP80nDvNu+f6OaB
AnuZ7DD1Xm4hLbfFPBM+GX1b1jsRUI9l8JBD3c+DjCqtJU4U9RTkQk1F4JRhg2J/
e39ZNrc6Cq3uHSMvG6odmwJ7w8UutXsUCnK9Ht7rNnWWC7/zL2+RgU1wwEGSqUYf
BzcvgG/kNCo6M0wWPGtkSYPvLoLvUbMCt7c39rfrkGhzFRmSDDvFWKLcfLPTa+qB
b6t59owDcQ805fWeAMw+UVNKViAWjui/Ii1+t4cpCzNGpPbKRw/lhagpZbYw3YAb
SuhM3Q0MvLWl8s/kH+QcBrrBLMoA9+ERn2slJJvg5KXN1QpKaiv8WVwwNL918K+n
Wns17IOLKPWeRw4x4g8R6zHOghCpBCLSftud6ezb7DX/kPCaPzW/wS76EaXMA7NW
ZZZ+1SrlYDph14ZmmrhLlVSV8zIwXIrljL4Xh4RU2IZldK03Ui8eeXKmEXfIa8YZ
C532ZD4rzQyVPAh6TSDuVA6lOaks1FeMnF/qIM4bgcvvMpd/yEXWNdQPKMAXCIAq
ugwcHd8Kx5dIjSEnWrzSuc3y+Kavu8k2sZk5hx4jpCZMzbVT83k2tvmaU3pgcLmI
Bjfca2bTj8PbMIiIF3zEypHcJu1dNOfSQrCXVtv6xtUYZBUDf4F956u2Z0op+Ah0
3AkA9J44h7ig6mRMr/kOauviBmYP25ywWyCBaVaeaJBd38pZC7o+dXbHWM1DI0Ja
3+ptHNFeVX06JmjfUzh/giGo+nENL4JP0OdWfPT9yQALvGIxEGce5tc8ynWHYYEj
T2uH0SCIs1sPuPM3PO94wwuL9H6195TYPhYhYmH8IiDyInhHxNgoZ7w1ov3g8Y+Q
BUIs7DFtidp17J3KflTsHcYO+Tu9l5UthIsI/jBq6u1ANmsAha9KJvdE+HGIgFOg
MwgDJdXDaiJsv2sFX8J2hR5OO6T9iHJYliUZ52OX7sDsQ+QIV+bDSazKJ2JIK2/N
ogZ2fFoeVlAhixBvgAPk+GhnJn+WRoasNiJx9Zd82WUK5ULgsXZTHOJdYc/x6+fv
Jvodkc+2sT0omwW9qgEie4GOtBB8562zQA1UQIGjjAxsxF9j+uSniJPdjr4nL2xk
jH3fALyPetlKdKrmnLctebScEsxq27/APvXdOOvbpVCF8VWzW97iVoDMC3OpwHo3
xYWKnN9oy5uD7KQDjmkuN2PXh4tzj1KZLs4XilcDBcZp7oeYM9q5VRNWjQoCjQqG
WdtkmzaozfQsr2ljA0TsTfKLN780f8PloqKRqWyoKUVrRIOxOAHPxRnwu5Yag6As
KRVzZIuUHCX/8c3mdmx3X54nMmxKzlIzq5WroFIkpIFvfQCys4esZKPX8gOymeWv
3TDVu+TFKKXCwIo2+VuWj9EX8SxAtTHJ0v0rmasN2JfA/2fPCWtDnpHPqsEo940p
ZOU0ie/zZ//SYryuHY9zY2LvIQrnrhyOA3yf9uNB59qJ8Qa1ASHSqiuLFwR4JVy/
KsbeVw6uOe1j+CX1oZu1dwgHhMPcXMmNIegep4zwyO67W2S7qeA6yjC/gqD8tf4T
/iRv7WqOY/J9DmFTQe5Qfsra6u3g8y1yWQIg6DvbK0rJRdEjUN6sX6neB7kwszEf
EV11AZtiOOa8+fqGS2FxhMql1OoAlQm0XOULVHoPEF1iOdJz9JlN9/hT7OsBBjYz
Ykh/xg9v9VSbH6tR8FFbWLmgfqS16gACQhUy/TTNdH6dynUSNh/3m7dGAfVEYJ1l
h5B6vfHowYX2xurqkOrF+aOHKsWek4FJwRqxuyyu+m9ePPM+9iuQTSm2wA43GAnJ
VZntJQcDPCMzhA4iWZGKdbtuKVlS62cGHc2YLXrnEB+kJaWHkZ4lCa5BT9l+7Ogc
9RrP1F0ytqeMicAcclmd1lb3tPy8gLZGfm1QPx6xoGH7GA+B9DwLJBLtgg3+FTIJ
+W2byOw5aBwDR/xrw8GYidbggDwUsELXf857nSW4MRGzhfY6A/+jMZhAFHrn5D30
7pLS1TscY9NMGGLZwIvPRbx9fny/qWkHnW1VqUpmaNjPdCZcuk798lQqsfKyQFiK
UavROm0lox6/VYGjD1swlroT785XmLNFPBDxdh1cXfBZJMFP8kxq/JzrkPjKOFfM
WURQm8GeY6HWS3fs0FtB7k05c3v4xDvCbpfjQQ2v57agYBNaKeSQXYfy+gcl2rwR
AoZ88X7CBcJxNZ7DXfYtz94jdu9ypF+5DNvp3B9emPYQyRYUV1HuPClxZ+19U4ei
eDiuzU9jC+OtsXperAW+fz0txqOFTFvWJUWjWso34pRedW9CAJf0b/sPZuBwReQL
TwNH4tdh3mkB2O8g75qvf5YSQn2pRtzHkUulwZhUZpHkhHhVAFmk8nXJXC+ppwrn
2oiQq3iZRYDLW+oasp6EBfmbldlwfTXiq1iejurY46crU4Xo8Vozs1RKB77a9d7l
BHZX/Ma1cuRsOw+P5Fhg/dP2gKNhIM0xLGTIPSAFJR8AMgvnrw8zi3tY2e20D5eD
ioVbL99vokBO9jyvDwtFR2X9NrylXLdTAobzZ8O9S4wSGXQBAvX5YapruKhgCtfl
eP9BwxvhIjjQ2PMKRIvzwCiC9p8dVP1RCegV5yapKR5+/woAJgQlRxw21wmmHI67
CKc46GoSihmZ0l1zXGCImI9jHlygaJ5fR/UVEBak/UP3PBmoh+SVP+hFHD0gZf8l
sRJ6KHE0QzAZ650+EZCVWoH9FVLHj/XM6GyEBIcn41fcjeV0UXWvrGJZjo7jeRwq
t2kM7GmGPEtKXNUkjU4cpSz+4YbQvrjscBCVBoqJDm1hrCvxQzLy5k16BcVySPZ6
VjrCEZFQkMg92aMZfpMyTgutnET2VA76/jadlgd1AZ3TOylQr3uKh8lUzVO9K9Ge
txZFj7WsJk81Pw1IV5xqe1VPbH+5qXHolLIwqiUhKXV6XK14zKT47t5/AJczzbas
nFShWHoruemecwIbUQmv57W2CiLCTpsuchhEwCptNUubcjCEWY9Hcz7inkJZEpv2
u0KH8HLVXvBhxwXkrHRx/M372tzrLxpFw55Q4NurCxP3xPXTualQoW5Faop4x6X8
8+APBfSb2AN4DpslQa22T0jqzcLxQcEdPVfVAq+DvcnTWL0k7o8s0a8sDOOkMUFh
GS/hYpdw30QEX6e9TuuBypPJ/2sjz83o44jVAXO85li275Elh69t6zznKNWkhSjo
fFRE6KAbhsIGtD0t6wswbYfDFAoi3CfIfnMIgqOMWGuXr6Z+1hQLRSQmv2TUjI0E
zzBvjJckMEqIAV/oSnaJokbhycmprGcaYEib6md57pHJmYx5deAl38YHJnyhVkGq
pAZAyVaj7JPOYa//GypiaOiJA5f5LBCH3NGJ+7/ab5bHuK+q8l+ntEoLQXMv5NIF
JI3ayWitNORlpDSe9zfYU7mZtL2hmmWx+5sFBDq0P/BmRA2M4LTlR1RKAf39mfko
ORNx/oaQdi5m1+9ZfsYCUlXKNGIZKIFZbNanFdMW8E20Ok4UmUcNA43arTVcAaGk
RzlwIHGmNpTPU+MJfAFuJLAj+HxedNCeHtgXWj1IWK/lI3+B+d2pa9T6lLCJfIe0
LeDAV7/ckHSPsSX+xaBc73E00ImIEcrRuIIHjopB+1nYWtZpoNO4azTeh8kMpAqH
sJBKJKTu8+bhUKKJv8hX26S0+vPNcSYH8NJ3p+icHOscsQ9En8k7zkObLSjphi1v
GOYpJgUqQ/qesLVnI9yivsPGp1UewYgzqWz1PjtsSMRdZGSXPbtmpJITM1q6aGf0
0xrwW+zN2TPmPep1qtATFtZyOf6df1dhirIb8UDZxbUFR4GTqoEZ1CANKC4UC+AE
mHjmr7F4xMTtKs1fBHVvQ7LdsYkhjhQcwqOPsgBHaSxKXM2U4DsQ0yIFRYqx5skS
JArUFL04GjM0938ZVtH5emDNCbKhSwjjiOwQGkoRlYi2H6kOKqmkhN4hCavTr+Qi
FxCPPmw5HwYzKf+e0ox0eZP9zoLYLMxVi5xraHuwPdCAzKONuJr9K4sfX7yn1eDe
6u1Zx2Fp61DnXn6SCfJcdXbBEGou/Ln1MevRG+ejETENNPvBoDtd1QzxDiqdjIhG
+FHcTbjdMPBXosugczk4LrGcFpExh97pKFJU+4OJhfzhHmEr3viVlh9I6JfWSfk4
LyePZXYvXO6+6cePZvfcatiWlUwdrWeTxYA1jV4OwdT7D3dZ55PUL5ANvkDtFSuq
U3hWLHd2QaktKzBndpPHdYK4xaPJHaQJHBaj+NVOdfWGMH0HZjWZxz+e0+JBiwBJ
yC2jmznfB5e9EyLYiJCXDMuWLyoWlfzBSzVjXW46LlLLmx5Qq41KJo8CZ0cwQ9Wb
UD9asfzJmddRhuVlkTV4pRjd60QfPvVNNk+v/ptLc9BoJHwacXbLUjZy/b4sCYel
mvTpeqQy5nl3IVhJxsHhCezWpLGhMBgCRx6NWWo/ELYj9Q+LIsDziUAuF276rZ9b
PmYjl2afkdzVJ+PI+C+HnuWs9qiFt7BgSf3JS2p79HKUsqKt3i+3euYF9KywD3qX
Mnl/i5lcil+tVljPqmHtz5FpLHgamJjRGY/EnwRjm60EPPCwFi/q6W3wBe5S6jWx
j5BoYGxdflsX3H/mLgGspWfoNBdicnf0KrR9NGU6DX69V0qUpMRpl6UoYHfojj0c
7ZliOuJmE7HYotEZWKQVZPqEC03Ld38UfGeJkHJ3ENHPj/8WKfdPNh8huhixOi1q
grMetHQ9M4ogzZGqLkIUqbS30HLuwySWxjgnh+Dxa0qmASYF0nyu8ejM7u3R5j+M
xBq7w4DaXt12qYtL+rNmnt3WHC/RNQEcuvNkECN63jVlpb6E3xfQySyTFKff2yPR
90C5x/vcRJMyKV6wvZ3YgNsx3ZPBUM+mrNfpDDCLvnbl1xeQRBG5ENEkihdyIMwH
Eoontc7njx9DLw120VRNQM4cXn8fWyxNPZcuoBlOg+/CcMXV+pc9B+11OIp9PSbu
jY+dxSyih0XaBcmMikc2DAmMXb+jwKZyw6RWTImdsNooEjiDJqJNrMbP5on+4CwW
6TiyG52I777patqfFoyHJQzW8w7kjGjpZt0wrx05N45U6mhMVSilMp0poB2UpOie
vtDUdiybCoIZD03hMdI/86T17zh4flkREYcLJCIR6oQ+SDRiZNX8yDyyozv96jjU
pBiyXKEi8Jw58M8CWRvBqa3GsQr75GfAHceXzcg9jmSJ8kpvmiDZU5+DhyLeHGxG
IYwBQWxL0rcOLNoL4eoudSTwIX/P3CDF3+FZsn1ZEi+09CJWzhhLjd5Cceb/NqE5
Sl+OEEHe6WU4urTUVRSA240WZAnTVS5qKhbZuHzIgPWmP3ap4ln6RyYmbiBLtRf+
BCIaNDdQhhS2fBnWXm8QKoW3za42uycRnoavayDRKRe33PY8eRhnfzi9dzM51zzj
nqifiAc0ae9M7035HItPmVcipLVo1gLNE44lIuCUOpyKp7dsC+duJigqd84RWsbB
iy5kUq+zbyCysORJ9oDSN2mQQiqFBrxl3eMXH/B8KqIXnzMWz7JjXHPznXM/FOxh
W1g0WGKvA7WRi1nrRLuwpqwL6maB5Y7VDDwGQ5WYxpmLfnNVlDiRoyQFiECCmjwF
x96Z6K/sfOQ+txMTjpHXv5pGGMvkAa+xv2O0GQ4H/PfM+wwxHGLV5QsrOdG/OMef
lhMhGPV7Ne7pl9eY+nBc8eNe8Yz9focnczieIqkzxnWusKDd54vJMHGSdLXdwfXZ
TaaTzX7oIBIe0PUu+swryrDX0eXmjX1Ojnuw9ta7y7ZD5noZcS/Sc5jf/4o5wE1T
ncmkXJBlY3fkyduABNs7vNFEkcd18VluqZOfExmya+VerNCefCVjKkHBkQmpzpTe
UZWcJhM80qBiO7lSH7ypJR9VSLVFbiuaWg7FIWxnGwS0ON4dg++FBhHuGfPyPouW
IZM+Qt7rNMjP8BP1EGkPHNGIw60/L06f75Mmaeg6x22rDoEOa+rbN4YP29b8AVIV
0+jb7xwCJBlvXUACMyX0AXlB+sb7fknOUEuCnNBKGC1IWzZWN9xmsoIZRKrKhH2S
siFtHvVzSb9j5bZx7dP5HCqRb2gF7uwLDbKsgQ/xv6IWh5R5t2u0pFyoceWVWltd
aNeK/75M1Qr9MjaiP7S8QDLEeZKB++pUvr63aCYVvoKB5Zk8r31AfqGe7u0TrQ0W
TKTlDjd7UZM7dAbNj7kmgVyAmwa5j86zmzk6EK18UxFPybfOleFEHLPGsFKmlrzT
6+5Vs/AMu+q3vsldmQTFGlcF9WaRA+qlohOWuUuYSdPQRT0/NaA4AivYUVsAIBiA
VM94pBsfv8PkGRxVZS1rqFOS1s7OuXS/n/N+jaUGLV6A9k0vJ6HwHVEzUIRFGBE8
BVN9PXWMQ5j8OaDZJjhi4O1GmHnrBXLdKv0hQ8emyk3tlQILYOP6LaLVacpMMcqw
2cJMxcGo2P2KhCDeQ0UsfH4xgLOrrbUlkfnc0kYJj1TeZ7gD9UaW6TiqXVWgol2u
D8eONVuqQzNJM5XHRLf0w1k8R1s0kDca54jHCsgP94b/zXZJvmaZPbjPPmzIMENc
R9Qv+B7TRH5JpaIxt1TCRQKHP6LN6yyGrtTIk3FiEsdWO277MAVxuEfIv/kG1+6t
qSPwnHezQ1i8HkEsNf6Bh4Ftg3da3dQ8Plz4Gaq6CeRbQwAhi4uao4mIViIDkrMa
8fZPqL5u2AMs+fxgyEDRIgZIZPoucujmkbOET5p5WJeyyjoOkiiNi+QY5/vwA1mf
5yo6lzp5LpA08xV01DULBre9O0HUt+8fKDyvStX83BGF1V3dR4S1XARuMy95VLWk
iyYztxLmWJ3dAAwFekiE/VyIVdvvsI5wdLM0o6ePg52DrGCvnyS52LjByXFlX64v
82ij4rpDs+78RoMnMS7DnsDG7+TGLC2ZAozA9tKR1RMl9CxPZlVdJXOWosGAcsXr
0Frchr8EQLFJrgPRY7Xjdh9ggosLdqaQKVWPY2g9WIWnNBoRjvZMpizvXJm1LDFF
sMoyaVWno8215i9GNA0wfh+bdpN2RIp08VgtSeFsdT6Sr4zD/mpJs8eta0KULGxU
QdhhShklhYJEmxr53VoxFCINF6Kv1yEV6Il0Oc9K5CciyNKTDkLGpkC8krmcEBhq
NZGe6naPjZbcCpagHg4KyZWZKY58e78hnyfCkFiE3wniiy8vubenkkc1JHPp2Dmh
9t2sl2Y7nZY7ekKVi/GndCHoMmN6FSaXeTcNnKvUZliAGkXBeD6CXwsrpXpHduDG
C42G6MzEV1bZ1j27br7RrJZmqQtd46gq6trudTZ0e1joUe3A2k2y/q6Rp/1/UsiH
huGkaAA4pbeGqo/p72uqVS0UuyDKaiGdvjfmvPqG41O1kHJVDNC533z5/ZL/fpwA
TSFaNFzsJt232h5xVeDLEVF0N0Bvd7jhQhUPZof879VBtzsM80buWSqQId1ZvAxG
jTNbQHynydeahS7JDpAj/S1tIPQfJtQuwPZGwiQi7wpRjU5p/1D0lPO2oWxiO6BO
o5bmNZXXUN/1pP5xb3B/MLVM6B3xCJf0Hv0o9V8uXu+PS1V/rbilikENg4AhVlvb
J9Fx58GCcofJyjZrbIz7bQlAPVdmgC1u82cd6brxMSiNWwRLc59AxjQ0igVk+9OX
YhlJW9mOjQ31rk6CxdLRBesPbZqx8kHkgqIVUleibtkBOB5HcoQYBaAt2t5zFi6v
r+khNWmnTJoVdYFHfFGXJ5lUgytyYHXyl6Wx/M3kMrLb+L8PT2V2KHuxlc5PnQCb
AAZRvAtYFVFGLBmKbnGsrboI1u+BFdTRNTP9L1vYFar4FOW/HJNtrtts4uPsQp6q
7UQdoLw61D78/T27nx2Auv1xsQ2TdHXy2WdGKRaftHcbJljd5r/lGDN6wxYIN9OR
V5BkaX96vmheg6uAsaAEtTpjuqfIrYwlTTFKMp2FhfezjBGvv5gbc/CoMf5Kk6cR
Jq4toScsz9vtW5epEpaCPYizmF/33+NNzAmKKvDZwBLxqVBRjjjSekNqYNHn2+T2
uFxVEEy0TA2pgKcb6FfAMD5a2NJLoBSoflTsuUwP+6TXL+VKLkGsseKMYORS5jq9
juM0C5aZE3rle7bAqmkPm5vdUGmuZ6ENDLC8z+ru/o35KxiglhlyHG934cBpuEPR
sDfRnm+nrt1nqG+jLk+QRJeTR8J+HooNJdLAZXByEQx/7Lfvr/j/Pxpc47qxwDz+
/6neQoMQCZbLeZLmwWaD6DAy8VQPx9xPGg8OY8VftCjNymmw/yBkSd++FBwOPecf
dp90IbMirNPG+63xZRSgo96Z33IaxzwE2U3QeXiu2aRl5/ho4YME7CW2+iBGvTB0
I9lNF/On/tgrZdRa6muagdMj5mW56SXGcPmon4LDp0rAbduzi4URfZf1PcU+cexu
iSxvcypubO0qaiZS83Wqz9RashbiSGj3fsh/2Q3Bu09W33HsnBl8Y7HoilizzlWQ
kE3hRwUjU0FCGP/GfuSaqifmd0RhgkooTXYstU31hpyrPWqA7adWpchM0+2IL5l8
J38sIUTGf8XjIlqv0y/f1VvxavhPVs4I4IU3M22ZS/ROMAyZA7bLB2em5gWF8VNP
2izpNqgbWIJ1Gn7k8QKKazQ1RfC0Dz8N854dxlDZ1WSPlvX0Poh7vIS1KI9TQ37e
3dac+YDy+jt4hxYWoBmpaK70wAea6p19FeGhkbbAQTE7q7hghCO75nY+3krXVJ+F
kV22fyuE38v5rgAu7wzGmZLmn1uSGghTiQpZ1ITg9sczNoSgCMB9adimx1TRijzj
mdsCWSMgNLZzVTSnhjtqsEUmflIqO12ecU7yGldwi/RvB+Ey0bMgf5Mnkv+wrs+G
p2dAFEOvaeXMBAbWa7aE4WsPGzgBRIuN/aeGgdyCVK+bAh9HdXdtvBCbXdm0PT6P
S204VqXKqyAeN5oouCoWeXrIxbgFKNOYdFesQiBiWP3xofGrdo+03JTkhoT0uaFB
7Cmrih6IHrV1sc0kePMDJB/BTH+EoqtaOuKCJobEhbiZM2+B8kka/HDYhLRO6zO/
wckcwNjNmO/VN/rUemOCaergsGmK94pbGAcFLEemyTIiGTeLQBbCjqiWmxtJSNxm
Ti7OiqfF0PtNM+wpS/nAwX4qONRege/U6ou8okeDlVMNqHeQqmUB5P0uxzsnazRY
7ihoka9+4QHsLRLbDOlQXVGTd3Nk/eJojqQaUQ/1VN2tjoNuBnxrEY/zGFyG93qp
Pw7KWXXUACz1jbLpYPwTW++kA3UCnfwuI+VduuOIHd9T+KFcZH8vhU7NGQo1HVw6
z12AumKF4RKHUGcqdJroDL2IEy8ESvAbJoEeQneQuTExANgVfSIwD9LRf/9ktxdK
82wfr79weBNHaNzm39hz8tzFsDK4LaQgD2/pZLg/bdGBCeulbssPPmAUvZNGUTQ3
1grEW+saWEWLYjc8A7Mqk7keSN0NCmeKbPvrBInoXmtJ+Q5X+/yRFkRh62Ewk9tY
oDJlJ2wZ8bJJv24cAp0NhbmIlM6ETkN9cS9OaaaMZwmJSM440+f1hMPgj8TcIZCz
n8e3h0Mj6LJoi6eYTClFtby8Eo4uafF+jk+P1kJcTIgsnCq0atjfuxpEgbJYZ6oy
0PV8ju09+WKNhgUCzpvbXBaWiKirweUKqZ/NSnsWDdmuAzqW/kj9mQPjI0vkoDYN
zCxK2N3J8w0MHQg8ET2JoIbmVaGlDU1BPrfNpa6KKLOQMQb4f2Sr/dYnkJgprqhZ
EOVO5Oi54hiLrf2Uhr1SySK7DMyCwkofxRRZXCB3kucqTwz2b57hSuIpqWiKq/PG
UU6Fg0hLnqqAO82J7gUTGOyRSkYyfJjvU45GviM8CB/cTHBZmf9VHoFV6YexKPgp
gXQIM2C+nQ5REF+9gffCzYetdFTpP245SDQY+mO4fExFCGwoeh4a493PlCmERl/1
erVJ0Bg6wFjrVV1g9+S6cJY38K0vY9CgSLEOdheTQ8x9AFt9Rg6QpaRNVTHQ4Agl
cUWqhuBLlr9rZFtQXZJYt8OaATet9/YizVwvVUM0gngVLBR+Aq4dFmVrgcgpq4dz
ta1zVKjhTMRg90KLRZrT80FIl8oDk7Kv6tFjQD0Y7AaI3yxb7JRuBG3r7LyRMAhf
43wjcxZoIH06hyR9imQU9vb+ZHTPmberUOBjtlJ+wti0z2wZibZiEJs473SSMdeC
7U+RyWOmMznkHkUNPi+89o/hIB8/UENsXdSpRjkkiOTyMjwy2f7BAIpU9QdaY2z6
r90mMJop4GE0DPETPxFCVCMGgo+wcT7cpPQ77rpTCpGGbiRe3/iJlnUFypaLhh5J
oGgyUL8oVwCPw8EqgAUJHHxL/eAaByA2FahatcxoNhitBfUtFhL3RyYu9FjKLuCU
TmL5VVANRVyBg9CrcUE7J5JuQqDsJs4jG2YgoChqzZIXK1f/0TMSyHraxsIg01md
YpWXCKYvPkLVWigJqhyhVTejWa6cafshxdAnmJDkTTzIDPub43+48Z4w8XcXkHE7
t5vJo9shHAlENkcwtNGWWEyMwHy0TGsleQPW/jVm9JLfvRHRLPGbxN9VGbleuVm3
rEWlK9RMeCE7Cw9iczcO8T0i1kXfNfvLhTJ9/RpxE4aSxbETbL0GIc3th+TZamWn
Og3lGfqHppyUcEDtIjDv56/aqoV4XqqQj851s9lpB8SL8aaH6y8dhXVM8FG+1n9C
0LpEt1e1CVLS7BbqtFvNeorE3LYtkpv21gdZxD2Yk0ywFlQTWKCHHyLze5EMGWgy
FKKirbPNAs96Ytmm7u93IYWseqsEuYVPlAzvth1f0Sf6aIwNqOerdMPs8mfEWeiv
4z9yo7bI9lPvT989zCvtLfOTGqTj6T/a5yMvSX8UZtV+AO0SrgZlFMSyY+7QhzkL
h90pbmA641ewqPZDPXm6++yznJ3K0BuBbk0ptKfq5QCf6/58hGOmGsoQi48XvvXl
6dnY1NK2IOvUIBD0uWk7XL2M5t/jrR938F4kOkWEXmJ4UeTveeTt5j5gOgN+Vb5W
oz0OJ7R+IKzYMJd+4yZ7U8A3OztxoNiC1sr15a/OfvK4PUBgU2nZXOsUP8QHDItZ
DQP/jvd4leGRTW5XOnBLm1zO6XLWXhWF1MDNqbmCR/kTSsYiTJ+7Dkg58psQIKWt
CISxC6bckQo2v25fbp0ECbWI8TPL640Eli/IpvODpSsHaEJGwiX63XK0FgUlRGCa
zq8epc+3VTmmWglguhJPMgVuNvcjbrQUlDE49ebjMb6A++EfZ4MLbTF5S+R4dapT
sZQEWHSE6TqTo+CZN3Rs78f24vQDULAUHMZUs0EPpXKMf/P0b+H01ivFxzcZ90aP
rAxpwxZKb6uIwywtBPuSvucYqsm3sGcwiAGjuPwaEvRUGBVei6V+p7j+0gT/M01M
we4bKOWH8As1XDQKIZAqOf7Tp5cVzBhbULjinB5UMhceKsu5WV6qVR3ANGLYxQ7e
664f8/dHfoh7fIApsJNCYJNq0phfhDPuaOw86jTGOZZq0t9biTZ80oGP1nAVsBd4
DoR91uZXmuYqXjc8y2tPy+knOrz1QaWW/TRbgSy+aS4aeZcFDt/QnG0oYfBBg81K
RpnhTXkN2QrKnPD/x0dpySQFdCVBJegh4OL3RuyCoWCQUyRJphJrMCAsgKHl7vTG
iWd1D+ryAsmqi1vJLjnMNTFhL6euh+Ghp0z8RDJJnLjLgEkeA28H9Z4aIUuS/Qzw
LMCtNZ8KF2RZRBNW1cylhZ4Lx+UoQ678Z/NQ5TiT5SzpSleGxGYVFU+q3wBdLgiX
F+5yXOR1FE/m4F9+5OXkTOQLEfHdmBbbwcQCnzhSNDinLzcC8zi7WBIArT7ffZSg
rIQvX1LlU8tV3oCHJsCl1MCQhB/x1sD4Y4uqcIrxYA28TZelrIAhuk82GjmXXvQd
fqDn2ZLQRtGI+dgtCauAV2oipXH1hGjo7jPjJuLdftkjFiBHK/g24kO3usJ+LB7A
9Wc/gjiC9TrzBC/Q2rMypMt+ugMdxYzg5y5zj5DujnpGN5w15iyafi4fe0fKz2SL
ROX4sQ2/cUlrvaEzG14gf5aHbes7w14QC98pYNvfBf9Ekpq87R2JilkRXy6w1/ad
eXDe+nlsBjI8WXIDz0FBQIg44s+BHMZJN0mXk/fnlz/8Ecu3jYG+8sRe9HwJDvH5
6pWCeRJFZlKHHb/8Y28keBv08p1eM0FseXO51unb+AiyO2L5O5othuoFZHuhCNK6
B4JDO4+gm8u63qSylkMUFIuE64NK4D6tbJqMAkFFdniI46SPnEeZPJZxXsOsY9hK
ztmDDCzEb/0xeldYepICH5D6xTtEkbZT/6uQpSNSwNnUyuMw1nfvvESiJ09rX5jx
/j5I9CwmXRdjh1Lvev/d8d6OBXSulrecRv7Zus2Nlk4kdbywBeWZt1TKHaH56+Mg
2WtTBDBHBycCmwqUmVvU6dU6Abo9Hd84riYx9JGL9UW+gNO0rwy5DlpdL6KG0Bfl
gZi3o1T353rtH4gVQA3oDBMHO1bprdK1pPSxA1nvBXaHnsJ/J9AdarGrQyYOWxSX
AVJQ1Wm2I8oUHWgPW7VqW65tRGB25xnUUrYxaty+pt91MjLrUgkF7rtv12rETwYu
TSbOH3Tb+h8tXjP4YT/PpyH5biF6F3M3FmeTQHDysV2lTABHDYQkGGr3lrOrVFoA
5M088kN5ZtxIul2wZ8Soz5eEH+suHoy3SwE2eRNVD4HMWidQe+fO6GE2iUgHQR5A
FIR4ghC7i9D9V0xI1YPPhFZGG53wJsOSs/5guq56gWkzM8XbVXV9Je9yILerEc8U
5JeMB3T4fHtyJ4rwPTdsW5+cI16z90z1b3lB3XxLjeHQTr0j/Wx+qaBpIBzX3rc3
nkTWj/xerslKe/SwVgIzUFG2hl2fy3TEvb4BlLu24j26I4bfNSd3pKKIx3cKuyd0
25RQGTg4VQQl5OpJkllZNjdRUUjqFBniSLLSiDqi2wWKEY8vQlaQ/DijOZHxf6Gb
m8HP3bbyeeKD4/KaCKJhWfMVt3LVRm9JxLGLZVnwOTH3YNfdgJfv2vlpqahn2O3k
TUVOi1iL59gMMGex1NDGcNsho40dpU1pC7ErX2bvc87HZIxz2BY0S+y4ioh+/Su4
9x3LFwXzTP1d5KvN8rTAley85v9bCV4zslAFCs+vcYPY6wOWQepYiI7sXJJ3nHs6
Rs4lusSQ3SWVvWS5seXap9Be5T4fNnnTdC0QHgS8lwWaM263gghdQJHIhryB/joe
kxIfPr0hvVNdrFIr/i7EgUebZD4s+6KZhq5Yl9oUIUXQdOQXjOWN3WNpW+HkGgo0
vpJeT4Rz0zYZ6XwC1IZlQqjPB+DLsyjboZNAu+MyGi+nQeSGkfpMbIjMdJT5rgua
b/4ZMQPlAJ5P9QRJZOzp7Pyz4YNUk+TgCeJrUHZNwJ9nVjxrKqJ9Vx+unRuh1E3o
tZfbwB8s2qU+Z5LdxzHiIndWujubSRHtaAE9igdsN+mY/3rLPYB7DMPyt4a5OqEr
nnRHfkyYczJjur5a+fCxQUXgJArwc13+ep0QsA5ZS2n+eqILmRjsNYUVInkji/kA
DnCnI9/w7Fs7xN/NpqJI70F/e/79rjBdb5aTdlmhOGl36PzyzCMEL9zrtbv1ETJM
WowQe//tqEo3zqg7b6qWvHomZ/M94V6/mInD038lvWdFa63RjyVBfqc40ksyS+iT
jFc4khC4Sr4vuG11KHgj3XUYGaToaiZF3qIsZksWNtgOGLKR1YJTGbilkyEeg3RH
b6SVKNimtkLaOFVk7EsEWtNeOlpmGm3fYOgycMvO6cAIoTAH2dwvW2R5F13/kt0+
aL328I/MIkR6bM5TMW0115hLjVlaHlzhLu8ot1HhiHQYQ8003RR80GjSz1W2VphT
noEQ5+IaSmYLGnVFJfivaEt7s0cY4hontqhpMXpXDPGGcLuKew+NFeq2AAczaHPs
MlBt/bVjQAbaemC4UYSgxQKsXhYBBo3+u3S3ZoM5aDW9EGTxF+FOtlmaa/anTc0X
LMQEv+l2iDqzKZz05QjmBmB6CN370Ho4Wc7ULfqxQSZPTG0fOvZKNP1sMjQ9YRGZ
AQdgu50XZbqlWHNPYhbxCyk128HXD7H8/vyMTRJsfMk6JdJEhzfQwVyd/7o7obwN
suEQEQyXFd1wKqoVAbCUok35KYcDUB/9kgaet8jBpHVvlEG2w1TuBM4lGQGIYJT2
EfXuXDFQaCAapAjo5JvO1/urrwOtCWBToj3LHzdytH/ne8L8aDxCMRNeA3X0o670
lDoalTD75e1Y6Tn6HNWvGWAToJVC2xPYWTaUOmoFrDoksnPtcmWy2ild7vn4mx5r
z+U6MOisni2TbOP4qk8x+A9HzQ6/rQsWPUMkU2+2wtfDZ08YrSWuykANf8ryOwMX
+CtpNacTNxhQsxbgQpsFfqEjI2x3FavYGzrosExZQHCTqKypW1RKMdLsFabXuKPI
4r9/nG4FO1FoohAxGqCzFdZRfBhgg7fNjhZG+LijX+u7NDo0nTWa6aFSgzXm/96Y
AqnL0vZMeFDRzaM4mzoxI/DtWlBQA0X5+/RhP55Lr3K9BxF/jDnCbpb3KcEmWgq6
/eQm5k6lhNzKC0Kgy58kFbjmWOBQhH+NjAEpyTg2ZLBKl90Pgz6lN6hiRVR4zxe3
TjVHeuT1+re5Kl0QC6ocSrSyyFHH4C5cZY6YCi36rHdf+Kw9zETlhqGXqG8urCmM
W11LAygZNUC0qiWS4nowWpcBx7oKffGgpifGys9l8yH8coE1wtOtVT5yZeEEoA6J
QFLm/Q6UISEi9KmaqQAOorS/x6JFxZb0fP8SDhmxXq5NZUK6Ci+zXXbyDI8Bd5js
sLPW8VeP4PvfCRSmc2DC4L+Hb8ssM6tsWhqDUygi7VG3cLzQX+rz3u9gMvkuex7h
y7LXMDRXlgE8W8BCPL7RNIhrQHu/BLpJVndioxjQpJYfRuaXBZQuGTmucI0qbUVH
ebm+nkay9GSPKuqEv4u3R2sjjctVq9EtkOYW7GMQ4smxlLgBOp8vbjyspScijYgc
z90A2bqmh3iNo+j82MA6RSJ/kRM4f/PujjM/yK6ps9wc/tQCYU5EQkTr/PGLpNWR
gdAOst5EWpH4dABDbyATGnAOGnjbvUBsGLhnCt2BQGOvC4w7uePe2rt/sZRqMM7I
rKB/OZB6lia/KuZagE71vh7szVFaBxp4XS0dQ+k95JyeJrcmRwydSbcVx39ixiaR
mciaouALmB9ku59DITUcbwW+UiobeMkxv6ROIHELDVmcQ90Z2Zx7GWBWPv9W1Z3W
Zq0DIVm6fev3RCyxFt6O4g0GszZ3zCW5wtpbPRwUEzMpwsHWTz7BWTxrjX/9/huw
s+NBN1sNhjltX5LufDynCGuDE6COcY5lwT/qbodSWeDENUZo9ykja2FghrLv2Lww
FlXI9hODmaT4Xvox62ArL3ccD9x/iTpr39p1WAUxad1ixcgmX2ivDXHrV4kVXJEI
J5rV5224hgsmZL/GADjEk0xpK6GwBWgPIZ7pXXr+8ZrJZj6QcZ6+GO82x9GocY90
pSj/sZgG/H9SF+r6SjTLZlRW1LCaUwvetJrsF6ej+C8A03SH7wE0P2SdWhuhoO3s
0kVqJm2+nq12dgmbRMj9r8r+qYs04TyCfk441MkjbEGXNZeI/4g6Pq8Wx5Izu9f/
4GmG1lVk1An8bmn7F51z4zfQkzKayfEIdzzSK2CbTd//2tTT3JNCywbSh8BwCPay
b9I7YcJKTPZt7J+7XvZq+GMS1yM97unnmmgiUmHMv9tGYaqwjVqvv6CIzQ/zQif9
y4FtgDSjTIIUZ0WR/CzhlaJ1Zcv+vJxDNdXK5a/P6xOwtEpNLjx31WPtxfmQhIXd
24cRBMWS1gYsg/9Hoie2YgabnC6Cuy2ehFbacQt2GShzjP0kKqYzTgMrs2WXSf4s
5CjFZZllrvMrdCwiS5WjsSn0xfJjJuW2WpsnMod/49t3wwPuWUnHXciobbARW8lc
BumsVY+z0ZpYuydqkb5u8s4Bjp6fhBmhAaFFkIYHJqjJhVdt2zHH/t7MZeZnsQYq
LaLX9KYeGX1Og1x7FP7l9M0lXcsvb8bxOcoX64W2btAHoBjaJkxu6yYq313WgnHj
eo0LzgQmZLkpcQVdzts4hzfI9OkE0gsTBCuUypOJXjg6aw8mJz4WiQdNDHCvY72x
a3Aao0KbLSNo4CUKRLKuXVsRjoTZVgRAkSztxfwwM2DqkHNaCEJmnaLHyJMpvhQu
N7C1uxsW7yd3k2ziiNQtp36Dli4KVwaFNfUpeMtsv6L+eslykdQqlUojvfd0QpqM
1Pbt6G9QsI42nKk3mLEWckMa0WqOs2e9dxvAdaQZGgxdakwcZ7ojh4W/+WLd+CHK
qTNFIFizwhsSEw4a6zkzHIm2Cehaiae2uU249kluxLgiVpIYMqEvduLKjh3MDPHz
8z78Nmu1Vo68jX//pJCrYMXPmBabR6D2g+7fiPwRcb7BIFQY6E1A7gBAV+n5NIlG
CEiXeOW1uJfLLeR3xDEu4EfByS/DRw21m/dj1Er5KHivv4LMPnOjnNohpAxcHDzU
H3Jmp3NmcwNZ7PqQ3pVcweKjTHRcrJsEVqjUj4nWVX+NNSQLQ24/FUHgemnkuKK2
9fbmsYGnFlA3da5vfnr4PXAWFtUPWihYU3LayK/I/HfJ0Y4m1kLq7c1VuRBqH957
w4Zq1Xsupwia0XRcRb53NGEB2u7oy1HzzR0WRh7uEH3hH8DJT0JnZRVTiHpO8E0O
+hE7Y7Dbr8Jec6CJHY9DX37jymB6IUfqysQwQvgXgtjlkJptu7yW+SyQE7njt344
CKXQrnECoaiOOBk9Tokn2ScXqoID15u8q0SN1qLBditP+b1FJqVfios4eY0IaDN0
o2QFWVM4XI9gKPSteot1G+7nj9hlFIBNasdzbiIHJQpcUKbLf+ATlrtIRcO79AKy
XBxVGNbxDX9dZAHf0r/OzKT65QpXf8mR8O+YAI/00e7r3ExWYJOEijIIlGjhtg2S
2JxWy6USGNzvteDo11p9RPDUaVspz5NFC8oF4uczxT3Yz9DEs3hVbtrz2HDMOqF7
GwxUYt489EIW9IEj8Ps12RN/qMvtPiaOJj3qoY4KdYK7VPxpFBeoKeiA6YxXVJHU
DbAYK0wG2heNsckOVGJpdehZs2M8X5RmmU2LkONL0VS0DhDgcsFemI7BZ5ei/amH
HEn+bZexHUjZvEuTrMd6juAht7MJrCTyazAPkRZYvbyNt0IaYhiA2LUUIJ9IcYRw
f4o3iQs+Nj8xXip4Gv3o7yo9mqoaHOJnGAxPLyE7B686s9mRy0NSZZkPucY/ITTc
wBYHGckseDLZYCPkmy8SAKME5bc81RzEJCq0Lk2qJC8Z2lHj5VxyLQNpxIEro7bH
bTNNbsrGIuwzPJNWWgG3cdcZSAt3WBxM59wha/S92fC7KEPPB8uL+gmak2QX58m8
gjiSrboqeqbNu9Ew/DhKCXPSo4UX4NYFTaaSqskSFjPUKfLu0wlfxcWuFbCOL0UW
wri4Uw0/OWvB+nh1Ahsgx2FZcKzCh+AUsGvnWxFo8FB31XM2gIFLjGuI8fZWxoH7
H3LyfCETwWXEOvHtR7FH4gyHLCPWIR+LtF2SBpP8TF7n5oAvrCjHBKXaviRvocMb
qwW9FmTq7BmVqtkQvX7PK92Oup149teMCCJVuvjUyBW0AjlKG/cuLiROpxSShlio
lNevFS3IQ0Z++1CNOZsLf7RJYZtJ/k8gMOabdybi5XcMQGqyEIiS9A5kWXKtSx40
n87VKbl7hDaQmAZdiEA/OPOJeuNlI0AbjSsDAkXG0StpPeSSnng4m3d+lJjDSO4A
AqLKBnPTsKgImTV382bHwcJEA7j/hfmAx1U4YX1FZVIyjc5+Pi2VdIv9Xk9hBB6T
KiOWWAUxOyQVIlH2RQy6DNmS2yRaEtaydOLRYyQTevnInIzyjTok+6+kK5QQnKsB
nPL7zs0Bu2N+XOmNgKSLf9gklCC25JTK8kTIOJrd46jf9NRZKNH/+bYBPZjhdLuL
61lL9cSVrJaILapz8gVM2X4IzFnfubNH8d2vrPrKgcXc9B+5J7MgLvOdHq3ZPzx6
0ZS4rt9VDbjCzdKmD0fRHK/Al35PE0UC3oLRBT2/L0mdtmkWGQltAoROBqEBsaiX
mGb1LCz5xt1/Fmhezt8IP+rjD9rk69q/aaxoiueNtJTAptQ7qR7tYZRQFRR9bKSO
QA+Ei/kPTlg/Q/MJ9NjhnF7dDjg0B47ZYO+oVNZes2YNCjjkFmgkEs2rwDrES5ba
iOzQk3rJFC0+A+3pLXMN3w0AgCb1hQY83Oa+fmlzLg7+wCK2jI6/bgjUBH4H6ouF
hVdfHR+HrnySbTlnb8jXSdHPpJQc5/7dXDhOvTvmCCK9uZVbJWKMM5iALucObwCX
s9SvB5HHQ6dgIppunTSyV1YTbTXECdXvA6jBYkrQRW/G3BPqPlCBTPlcin2H1AX/
YKD8I6OaZh4r5F3rSOTBS0dvWqs7ZW9//aoI6TOoSH3yDB6R1SwpDZDWyy+aQuIW
Q1l6hgtV9rBjtm2q6RHrno9DURsKmKAlM7gsaE0Ou7Lu7vCNhJialIJORpqqIgSN
RrKnkCrtQLVfGwHHxmaLi/bd1E/uZtZSHBgKkemkED6Tj5yjILq9BPVxID1sD8mk
TFzT5iGwDhlzKawEhDfFVmuGovrmUINFJczFc5TQ1cn8txo5nBa9c1TovQ54heLx
VexNoW4M+DC+74zKCnbc8KiwgE+nanYhiwjo4s0DhBP4KbV/mxchsqSwZngyCJ4N
Zjcjpdibm16qWjxAKf4EglGVEQB0CvyZy+CFq5MqrutXkuZ9Ajbj2vvqF89ZZayN
mrhnpd4SzNYqhXWhNH1LmFm5OTweZEFcnTgDQlfcEt+iyjlVjvtrTdUEbEfh6Crl
z/GS54su8uEbKAuOT18LsQNWM9iQh0PbffBy1Bf3IRyw2FqggBFDHmBM62E+sDIO
tK0o6BPzIirAnY9M9/jVHUV2yZ7YakRGtHE/5t5vz140mO1Bv0oFM1tOfVZHpmO1
qzmBJUj3p9rFqRX+Jlu5xcUqsMf+lADYPtF2HRQ8Fh8URGYthWpi0m92OWK8Z/ic
NTW5rpPF3oM5PeMRXmps9CToMqGNg7CGvz4UkViXPYhLfeczOoLg6aoKPTJuuyJ7
MSOMKbeYUBhOKEhHuoOb/4iYVjdF0SANZIpFy2GSEjSXwnvlNvZYWb7HeuoZ38Qk
WBr3HI0o6nOhrmauWBpAJc85pEG0JQxVCNSDe4qhusIO/MfQYX2i6xGbNOTbU4P/
RwRX1qvXkjsiyiB5Ndayy3rb7WKQF02I68r1f7mFUd5FThFax/M8TKES12x3jShz
M0lpXGz93j+WEPabHt7haXzydlhtHH42ROx+eGnH76zfKejWF0fs1wSKs8GMCS6o
IcOT2euyzUGjU8ECidIke+aycmz33mN2tlFTJdwtPiipzNlZr/pgtIqZSi1tq9mP
x+298ed/UH8F7ApZYq1ulcPbv3GGkz7mhxxU0t7PmnUY2ZZCCaRN3nzNPitipA7a
49fRne+IqZ8fRvJWMb9Ag5QSSPcHsbpOKCwLspBc9VnGzQkvRisQEW63dWqiSCkR
OTifo/+brarcOaVwha4u4zi58HO4U18vEHYfs+kDvkpiTes8ZJIZqM6EA8Woewl7
d9dZZRaNJDBnLeMutsAxdVHARj7B1L/oscBuR8Nj6Ay83D8z5i13b90gJc/GnUBn
igfK29RQL1t1JGD0pYCWrf6IgmBGIgC2gKP6bYpkFJ5IyZwiQlyRZ2Ny2ryvRR+d
vpxLw4VqTMmbP22bxqY4zjl0ylAY0LkyzlwQwTMA5diPZjdhPkUbAjPeNmhPY1+o
Uc8VByu9klzUL6fwrBDw8M4oakEiARjGqBMEkVG9IhXEfqG8CIqz0+/VA7MoO9Pv
ZdP2vQl5rS5Re3xraMzF2XIYykJEAGjimK16Npbb2NAGz5wKnqmDFegYrMfyAxfJ
mKC7dnSyeTyuExcpjlVPxCXlzZLkopnBV4gGqHz/oauFfg264eXjFB07Rp6LfZjU
H3y+WORLJAulAHSkcrtOg0X+UZGxq0US4WsIIhhyEglv3dUBngwbUUFgjD+xgVwA
fKX2U4ZDbkb91eTX5XNVZPExxh5eGMS1zdCTRbCuLzDUuxuPKfroDKKMHT7yy/Sf
a7LAH8WBuzOH0pkfYt6OAszDe/QLP7thC7axlNAl5SfSlJc0b0/FuvnnRwRet2OO
tMmPQamc6zfPJCz+NioKHfMlbGnHCBlSEHswWdcRA1Px/fd0kKQhkJJmShwECLXM
XyijZH0W6Cdz5VOShMcbjCzfe+26qQ1NdVNx5kNhecSfO8+WWeRanoXDwz2yCQAx
AW/m8ESlWozD9PCMM878UTOpK2Feg5iM3LkfxLBPC/sve6Lt3eL1BURjmCnsWJWZ
iymKLe0NRwiP5vFDy5wZX6juo2xoy4st1YKpJODKmNu12AbipLm6zXEgpld8B+gl
QXf/PlK5bMyrDSj5kFHkrNdqKw2MzSEusgdrrMcdKyuKsATkY5aF+26xC+R9GpqQ
e0ZzhJNW3gwd02FxU0Cbjn6n0wptHPDsOo7q2OG00KXmvRMgDOg/TwPWFINH6btM
3UZdLMTClp5nVcigBBofrunnXoS3hRW4PbVhFLLmGlaPo1S/9WyU89sPGXJHmY9U
A6/KQKxcpAqT16vmkWBUZQJsbKxWftwt7Ylh0kUTcD9aUKGp0oAroXwNTE4RXZwS
9SGmrIwj8hx8IFnZP5VlajcSHBG249tP2OsKb/p8OIs/g1iiIXsH/4sjenhyjWZG
KHcb1f6ei6uUwA/LvEPsWbpu+Fyj8KN0aDBMssl2iGE48QDy+AaaXDosDeBh6lo8
9f8H0z2XHs8rfm2jUU2uEq8S4Y+qsDZI+rXGeEGH6XlA6jfI05YGdYVVJs8LZNIh
BVVJyZ45xbHymVFB5oAnzAx/TkT/DRJgpKHt3mAkya/UrrLfSUDq7XZYmA4TyEmR
CMs1lIMAv7oXSGhmrDcu46N2RJ91tUJettTsMghLKHIr3WsB7KXIcRX6p5DLGUg1
ZTyJtp26h+rnZGQyBGwysMtbWqlTX2FNDjdr6g4clYNDOdph8URKqZFslvnGQDxf
hFy55XpjQPNCX2OZblFXfsjYbFMoxOJhm8WykT0odcwkz9+Mjoh2q1Pgn2OGbUW6
2suIIzI3idDRt2nk3NZomTG38FobDffAo9udMvO+gPrdAF/6UQ/Ct5l2aO6ekWDe
wygrX+BzLb4enYrIxNYqg8qOjKM9yVax+V1I5CGiy8PCkoTWLOA551zim64Nx2oc
QVV4pEY8R/DXv6Rt6NmfLHq1u0RgTJAEBi62lVOJhkvyg6veNRmZtrA2c4JyPrUA
7GJPdtVNqU84SHkPsPH6fSOLIOVmEqkThDu9PM5GiJX8U5KDm7bFh8knwfDBxhOu
LBmfvpkJEbtr7SatG+BW/YSRvuf/fviHtQHbh5WH9pcq7p9ABvF7OFBlOKCCaiCJ
vN3Ry9hVh5abZOJTqQup6PDmTY7VTmhRwZOlRvOa6gl7NuR58UpGNwZjvfFqDRVt
IKUZLk1+dsFr0A5Xo9DqGa9cj6CeYw54MpvC9R5DKsogdC0UfRBfgJj3rAp5jM3M
3OclHu2iw4i0gFlxDk9Kg8uRaRGejk2cFuQGILOHT0jE6KvZ8Oc14MiwTr33DTaM
0UhT6qHX/sGe3JHnb6EwmDD+VfRWy3YmWflDH07K0mp6qGl+KRg+I1rfqpOFva+s
EeRvFn1OwqrFUwA8LlS9t9yI8e9TaCfKonU+O9gYvK/mF8QcN6PTTKy2UqBzPONP
v0Y6g8oKik+vIfWzRWPVLxHdPceA3TE1UylABWbmhwHweqgT9ynHcsf3hFX/hjpe
2cZMdb+SNHrFHxuBWVEbr5TlY4JtjVOwnkUx2TDOdUCH8VMGApKP7/7chII0yB4V
PTyhDu1rAJ7Lm5hAqQ8SmtPrNW4xw3LHQFel9Ow27zSmAc6g3q9jpHoaTCPHC/uL
8N+n2ksFtvWHCH/Jn4uNYuvMoAMpde7tERYS7c/pVHJdNHTErQ5qZV/zE8ar5g3E
58ZUZigGD4KLa4kBQEV5Dhk65K/LmNA5GSdvqrX7d6l4Q2YM8kKDPdiTQ53BSNRS
tc+Xojbj2AQRysLUPUV/63srl1SdTY80haDTVwddNzAdafIqmwD9hTXreZeEn4N3
5922ipZageSZamPcmMitM+AioIqs7/Ui0AJgLLY/LB6+3nXX688UJWh572L8NvY7
hNoLHe8P2PEKTrVwTCDYtWo1BjO6uHx0wl+xbPgYL4zZUC3ZEWSMk6Y2427cRleS
RnOICN8JXpJF8mjKzBQIbnGCj9DGG30hvnOrp7RHYxbu65co0ixVbr4vZKpN90iS
5fCa9hf25KLOPvAvLaR1n5yoVZIrmbT8duZNb/kCgKP7x4WRkmmzLgIp8QfX0KzQ
K6XXyv0nguoHRpAY4u+stM6H0golzUQL/Z+wkZqbeZWAaVIPFL8vzp0o/VEuT4n5
jd5S+qbXR9PFQau+ERUMjIvGovIf6TqznYaxPovdvgNOD63l0Rjq6XG3DQXjIdn2
emP/H6OBk5LRQ3eAhyF40X9vqRti1n8cDTdOeA0MuMsG5thVzmYw8MA7qB1Ycfs4
a80X4j00kE3g1/2bJ14yA/NQxx/sJGE9YbKkh3HobR3C0lJ4ZPft6FkMfknGekYx
qOpB8YAqTlKZTQhNvaCTzNVRLYteadNw62JTDOH4fmND4zK0L/SXMREYSyWSoAK1
a23iTScnguY7ydK/LLtBa5qmQ8fWtomMCnj8CMvEMn+V1Lp3bJs79w7oVi8Ztx4Z
1G6F7gcvZ06MiN3jle0tlvrZ7zJtmY0neKoNRLmk5RyxisVK1zOiMpu4FzPWJm9b
4cF8mvip3BdtycizSR0DK1zHNLeJx/MkXAc7fb6OpIB7wy4qXY4wcMj3DeTxhr9G
q+p1rmHcxWQTmooENQ7uP1D1+wWZcq5cymKknfHOaelsCLWM5LomphNkVo3YVAoO
/6PvooKU/vUwiMdGq1NH3CV0vhw3WDlGID8fZ/mU0Ff/RPmrzOt1y9GQGwt4dQIg
IDxLHrJ9ozLtO5EntkYwQS2hjoXN6WNo/f5Zbic/PAEf270lU2Fs6HYdusuomEa5
AejPM/RytGBqpJS+u+qHIcangk+d6tbuR/vs2jqqhfoVFoJ1OgEJ3hRzn+JlOpik
H5idk71i4JMndBOY+qpdRYX6WiMLJa0A53pHHbSZf/HMGngDoj4HjYxBhIiyaX+b
61OxGftI8EW6+EvMrEjc+4UQcpjNMsf+dKv9TGKd/LCEPg50NA/cz5ISRIuDojC/
YLO1DFxfmlgc1ltnjQKF/kHaDehzkkum8tmpgq342rhuEOJqOobRtXCUf/jGNCc2
6zI2N3qj/x/F6fGNM6ieuvykwp4UqEWoO+J4uyd4SrUJ6jnqz6DieX6keFBuVT41
9tdt+NWM4fJ0kjluJoQVrCI6nEV7qoehzB124hLl6niXtAqD4dDVV7ayp+pXQY79
3qnQydt5QPS1tMOlNk08Kgcb4Jo+aDa3A0BCw6LjC1q26PlJGRCSY+BkhgEtPe2A
S8oYZplAyfTReN53OZDb5zv4faCjQiKNexlqXHaJchjs9lnUpi/wRE9t4+gu6XCP
CPuyPnAKoePXgBQyj1lQuCuNCsROA6kvtD30kehJIK1QShn+k8s+wNv7r+sne3Dw
EuLXaAL7Bz6+quQexwNyBX0hBHB5keb4pE4BpXk/8FEnTgsCg2/PLE2Fr3Vz8c77
jmirC0kMYGOW/vuNTPKnKFB92EGNAts6NDqfee0LZc+obdbAgwP9aJyopPhYtBy9
BSyfejKHs5zuXb1cNcvjyGNtVoYtpgqTarRlDNaG+3gIl6XOfHj+N3upslZDDKB1
sTm2YUXM4cqbXQLgSrTueiOsmYPlL8vA9EQfRU3WcPxDGKkBtL+wphUnjWz2IT3b
xnDZSVkIb39o18IUcLCm9KRUWRnCefMi8HUaxyXL7BwHSaQP/VAVbnwAVlhHRvVF
pPg5JcaB8uwKERswN+Q15QLK/NfO+6JkQ8DWEZWzpScQrxVi6PsfjXn7z4JvsXES
rEtiL0AuZZGirPWznCzywS0H8DKxMFO2vX/9ARKbMmBBLBlQ1cfYYrhgl90n+VRH
MQKD+yd1mcspYT6mturfKRAnkbW7562TyYZvzgsb6MAjVlfjRQPv8qHD5A+cCQyk
Gf4cmRuBmADu9/fKbMdDNQ1pAgp4uEa9Dv75z70vVDepa8wStHfb7RK2UpgDSk7j
W9qEwokdJUOiz9R6yypiz/biv7UjPFAZFsYhrxROJt0AW4Pe4BQBeTNNzrXsCknl
roIwnV7mD05E+2RXXAAjzDt4e1x0Oh8F81zKEGH63XI3pTPx2t69zD2ojvEYt1KU
Sm102TiLoDrOgsWyQgpjEtUMFCBpj12XmKS2gXvGuql4cZe54AHFIoMt0OfV6kzt
cCaUZlJun+MQIYf5D1sYHU1N4QH/WCDQHjTZC5OEixwoaJFY6dej7aNyz4GWuc2A
FS5QvidyXPAXXvbiBMHy9UD7YbvVX9RWwcwo2f5bhakRqH8jTjdpfYnK9cN+8d+W
T1uPtGfG8IAiEjxAaOLgwLyGLmWOzhDyvy8eJntx8pw4L/s8/vb45C3Uez9BhMcp
V2YNQrEgNoKqrF+wu9pjRlWdLpa7vWtF+dLI+xH08cr8envwvz/yIPl0wfVe0g7t
C2NfVvka8uBEFAwqDJuJqH+hUT+DNJTfwyCSwMXd173pktyeduVNOVPjSdRFU/Je
JmAIdzALpNBWILq3roIwRhEWXu/MYYLSqloOkeheTvvTtcIFWGJe1sPix215czij
YZqHXDhIkIRHcD4Q1UHQppRI945X0VUvwdZKCGXSJJJmoqseRCoVPkvRvHimjx1R
HqxEo/UdX17o7M4EgSeKunp/owEU+AiLIl1MPmlnA2yQ+CG8Z6QUSib562Xc32gA
xQTlyrKhxtwvk2lvXOuTxupJr2IepFIlzZlT5S9dpDf48Xu9fG9AMOGn1HUBQxKl
f1Y7FhiMAW3WXm94RDxhaEFiUHqYXCi7qyS1cnLVqaUoOA0NTOr86wPWxDGyIMBZ
Xqn4X2vVaWm96WDbBJT8BM8SQTdURSqvHzOSKKoDknTMFFpce6J/gWjC3+wCBO2i
e8Y1z3E40uEJPjbIMSgAHVr61oEgJ3IFOpklWqcowdzQbgTLb+4sIHl/tySloNhC
lkXrRDtiyttSoOYm29fcPeFgKAqlP59tTLnc+l9KK9ayoSOmg9/AGLg/k41uXZF9
HCQEYYbCnFVmOWORkulpQbmnX6vd9Lmnx5Hj+/beRp8owTnuzmOYfxpCUzaAGPyd
OfjArEgKxgfIPCXd1rS/hKtf99SIR5d1Tgecgb06bZFvwkm0GPZTshRH8Tide6Rc
qPPxJ5//zixgKYWaRWWGZNvT94mPziZSxk4ZovGM9gsRv2R2RfMM5K0r/pWQvzAc
HSyhQJFaBTQO2XfB+cyl/A0OLwgPuBr3FYF0B0JiWr0UyY6ZRex4ncccGEN/dVLX
yTNcORrQ6SBFCh/5x42wdMyUw0Grd2C9IXtAWmUPlkqr+W/5RH+lGQq0Pxm4X9vL
12dcAisXTileGioK524ND4gmSO/36uZeXYHIHdToFJQ5B0Rg4HUN8PiG+RkS+OwS
AUnMZwH4NrQYtsLDc+eZU1KA9EudgC74AmYBedsuWebk2XVZgVVs4/9LZ3/l+Ev9
4BzlPa4ECegdRDZj0L3TsCmYukDJt8gRK6aqywXfgc4K57xsM2/utHvV4a4Mo+ua
yBNSEyt4OeYkakMqbfpUtlG+6NBUJ05T6XPfNjiYHTHWNOEG3JhJi+/VcVxq5FbF
Jb7dCoU9j3GOvtFHhBr6kof4/PvOUmqXYCBPulrCFwHZh814/d3rrlwlBPyOb2H+
0ktosb1CyWqyib4pA+iE09RyknJ5q/WmAbzelR69TYE1DcVl2XvLIIIUwbSEgzRb
oyER2U9tE91OtO2dMj0eh5x4t+x1oI30qtXqrtJHXmyRoB0aRsET7eQm0XqlZOLa
VpF/FmHUlxOcdKuU8dUScsty5zdXXVCqY87WRgwJYluXAdt1dQBPTBND0Ssp6mH0
+ZQA+mNwssWOLC8bEKgV8O6Ei526OTArmyYfcWXEpwRo3gQqxAlDzzNfLygBxEIO
CCkYbduF7ruS8YWQZIqlOmAaDTHB0K0khbYMRIzdzqZOJHoG4Nu/TqP73A5fZdEC
4JR5m2dBM/+kVDERt6g6wyK3NiScitKh1MmssRM7JbOQtwlo2mgG3K9NGZPtfXXM
oxlDdXjyH/JDKW5h0Ra1lmBOf3uYcToK8V0dwxQ/DFPx+UdBy83ovuSvANYahDMn
qgzAR09qrefL58pl1Qmjh68hD8w506/4Zw9ZaUhtpjP6Up1KvQrYKH9p/P4ltVK+
DCgFNT+Pf9B3tjhXwAYR3L2rXWdpB9edCJxd8QTyO/LyYtgvKmyQF+lLV72MPyXi
pxXWxt/xSsjyHIweG//v9vqfhBjUSd7yI6MhUl5dcyg6SVJCUN7VqsPmQna8D9qd
PTul+w4cAblD6/tjeCIwYzZfaColuWWpwciw6txr1ceSJmkVhopJ5UCqZhPJEgHp
o0Yj00W7VA+hqQBrOLo5VdWTpCfieXOaVA4igdaZpx4bflGHoKKDR9g6z/vshUkP
2lLiigrOxNLlRlPSGYcM6N6Zz46PnVSzNBMvpaXLn7PCK+YaKN/TiW93+LXcMXeO
DwCDRaVkyjswgki8t/fsVaOEQl0yJfJ+v52Kk+8feE2WKMWUXRWpLukWpRRfAMIG
MwbnxuG285bmGDX32Z4yytFkD9+B6SxyrKjIXBaD3DLVdPwShT89JoOb8F8lmB4F
2Plfxy2svzYDob6bTqpOWFKSZc0xJJO0bjDIofMQaeDkgtanolDROgKUQyhtLubk
BRflKroTa9SekJHuj6QX5sTfwLibt7drgxXAVxYaqDq2GuE6F8XDIU/B9FT9yVws
v7sdEunHpe/MabxsB50QR8SYtIbz1vIYKdBzANiGUUG5XNZVbiA0TVh59wtbIBVv
RhZX+EHm1Mu4DHTi3VKzshTz5Ry3uZojzGq5q5s8IXBb6Ts/aWpPL6JbozHx9/Bx
2ev3HTId0+Ve+DvdLJ72JNCTSz2M3aW4VLsHsYeD1g5xU0bh1Qwr0NRdL8mez5LT
BdWvoyD3hG4xXjjtSlHrAUAAdyqiK7qlUwf2ubgYxAE8MEUjCI9xtrcOg/yEMns6
2rBAxF1BtFcYEvFg+7E3MVmIsCrN3uBCVXucdsyuA1VZtnIhiWVivMSxIPi12U/m
/29IR92V94xUQCGmc1Iw3TnyDj/rMF3oWbLZZiWueEGVQS3HyKx+OYL/XVMpB2Xz
u7+cQWPGC6bhxJ+TABBtwz3ql2UUvuLDbLNWEamTKEMTrJPr4aKZkuiBub25LpDL
iIb78BTVoLPVASrf+1JhgnssK9KW4k8Z1oTIVE+2w2A13r2sqIz9z4ZyYg/C6p3q
NkHm/sxAoHNerAf0CWfHvIx0RNglcJ0wp7e+eMh1T+QABf5emOay8JqilW+xbRnC
RUEyr+JVZA3z+65ocdTMcTq3jwxqoWkdzmKPZtpiIFXA+AmNgRNG/B7ZwZ17sayY
ihkuoGFOgPHs60Y504X2dd93PCf0dornaNKglkMeiGHjZViA8+woemT9UiNNovyH
iJIIIJn0FDZagCqdUMGoreFkZMlHvtFqAeO/WqHXx8xx+ktBSnBh5vpHLhbTjn6W
v2n4lLRbNWe9QfqkkrSNxD/A8o52/nwOfEbU35rG9wGfst5dhCCyRqzHT3PM/YR4
Tdas7Cr8RSbTX7fbo2HES8Tu+cSwFq88OCGjn7VwZW9blRQoIfoL6OhExp95+tzY
hUYGsaExRG9dVeDFNkRIJ9nmwVj2ErnGQRFLQaeusngclYwbcWA8RArtJ98znfJb
T4ZsDCDR9xzT6Sv7IIpgA01ZEkZwjWkXcqGrpAlsmpzjRDmbSu/Qf9VyGlXdxylp
cykU64vq/7j4Nov6zzz7+N1tcT6Z70AAyLJXJ+EFcTPCCqFoiXm0UTBWze8pW1qw
3PRtR3Qy93oDr++2Fq5GIpCudfvc/5ujJjkG9ayWpSIcfDlocF2LhDMpzsp4M6Z8
dLFqS+awzspAT6hmcEOiY+eS9E9R32UbsaisOk9fxXsRYxtTp1Xq+jdOM0h7HrBw
QC2UME32EbfyGVQYcYiP7m+WRQsx1/ol0SU4eV8aJg9hEnh2z/CHzWLt48DrPUMO
GLj0udfBnn+UhtZdMgJml+28Ia/WomgoGfaAhNzpN9URaNvGvnAM72qs7GLF5gfn
uN8uvBpZBz//hiGSoAAGyXcbXf97sa+Q/1/94BxatA4/59XegGFQtkGCr6WliELQ
kM1kZjE849UypbkrmNKiF1hTPWG/zm0gYiyifRk2dKguWS3S00W4pvMIRsP4n4vx
3HEiPN+EycfuLfeYsOlYWvXHsX1t7rvRvh+yuabdKPbl+Z54/CAeVv/Vrps2aoS+
Ta4SYCLwTTnuDrA4krYurBafX6msUAO+JtMWrlpzlXmXb3q0bQKZftphs5LrGQrH
Dm9GiNDUW3d3A93pSuo17wthMjG3stLrIWh+C6LJg2k8udBwNLJcSFSn0xgWIa5L
voEogcA6kPj5CduCpKUbpWl4Yziich4WNd4uaO9Exq3Cr7afQuA8YhsnB6eP6bb7
ipr26FUGJkLUSbzQ4o5tcnb5xGpGwrHjxZ676tI9x/h2uXXtQbwfTlO/spO7LCU2
4Bag47oBBe8MMdnzcAp2mVyHUhOf5UCGvC4UCW2/wHx3Q2NHTmwnG9YOsjXtUGty
9PWjzIhNuMdlHLn5Hcaf8FFFTevf2jxjpe0oxqVb4SFAD4YOaR1c1jtMJ5zgwWwy
GjrSlriPvZ55ytNU6gdoPrIxbjKBPUeYsUnULlaaCAp8PV0VcA8tTNXNj7gzOJv6
nItBeVL0w3GyvL4M+lXTLJ/hlsTmYqCqj1zlwO1IbIRPnGZac1WtM31MmBE290hn
HmUXM8IT5hjgOtMrMh9i9yqH0sDoefKNww4XvW4b4QXrITuZeurRlqKHZIn5vEZI
ZlaccIGssJ6JVisF5ZJCT2UItnacK3jmx9pX94uMb7CZwKWQwpczHVOITliYq2i9
uTMUqUFYIwEVArI+hPiXK/rxh2S6GFamy9v3zpIcjkRBucXn3heAwsu8RqYxHoyS
5s8KMFzM/nsnpNQJkWlyZ3P2hXJx2VSRxA0M0TtZUOACS2+mVlShlwjT/JXIxhLS
7etjXtPME/aovCOORzJafBtZWVrhJjbwY3pa4B1DTmckl7svhq4YPomC/MtgHKiP
Ko04GBuGvBTHIv5fUm5KMWyGO4OlzPJBZcaZdB0kkIpprGZxgqy8puchuAeyMvC+
fQtlk9ZjUQPaUE8gQyX0+esBho1rqr8oRHZZLMT/V9tJV7syoGzMsv98neaSL+gM
T9dvYmlv/XcZCu71xQ4lyxy3+iA7+GbhEhVknloXFQhYxWZJGtmCJ4bAsDa1UArX
gJBm/k7CbQJlcjfkzeXZ1Eh+JYwkjfFpfDQXNEOZNlzJQrfuoJVNLths6hs8C1Pn
D5gv4EZVYpZJ9CBhZvzt3iwTtY2s6n7m5/d2JMZm5YZE2jLfZUloympm6cUVYry5
vCI9Y7wqk73g6uX7Dvg3CZkQAFhxrweqd2Ar3MqiJ5tIIfmFiuAWBDENOiMsGCLg
11egSL3OoY2OprBy3PLmGWGFSb+Zk7r5nzIBv/6ScEtnI8WiJVqIFCP+OfnVUs6e
f0cJlT4Vkl0zFKN3eE6P+8GwN+EDs/7hcwJTxaNhqbAehxwbz4j965a9WRfXh062
tbE7V3wIi26+/BVE82NjRu5Q+TJ7VWSUOBVS5a8EFcv39JxCN9OUVD5PhS4lWVRW
e1tX3/SNVcWopFqjbFa8G380dexxd8hPNnNxnhIO28r8zXLiBIjJZLRoJOYvOKJI
crz7gej/u0oucGK1sWpCDVoQ9fjIH6XGjXSpkpBrsmNYTsRO6FGx0rtFhQajMA4G
k6BzVTMqVboTDY/cXO+NCI8oByna2Js1lqf9+sA0E3Hw9PXHwMkNTqNCEdtp0e5N
Aoyd/G0SBsRaMB9ipTJ/xI2fbjk1iUFpyqHViTHo/8+PX8Ozb2FAIdnmQmnfFa55
9so3itFJT0Wp7sk7j0FVk7GVnj0bN+M+c6AuOR4SStKkX1FqRd87ItChiQtXj3ug
PQavYfKfGy8UX6ln3m3WyeMF0INiM44Ym+Pa1M70f/w9MDTgog6cu7vEZ5NYEUhM
ZpI3gg1mcrKSx9TlA1V80VFTSX1jGX71f1svQi1Jc0po7NPLo7zH+v97ZfKdjBjx
nPugHDurTRUxAroT+3sJhIbQ/vXRPzzMHzyCwjX4+/XCMej9bOfH/04qjJ/D92to
sFC18tax/xaU+U8WARoTrqndPRG/1PpTOFI1Kuekut5CI31GVEZMen+tiHMVG/RC
dZ7CqB0OE55QJS5SfTjV+WzE+Pc4XbpycVS+H4CPvg13s62QNZQRdjlX0t3I8GJC
Dn6DtMtgux9EbN7+i22YLMaHu3qsei6iqWaN1yWU0wgI23dCSbBP39h+aeEF2LE/
90+jBJOK+L+lzsvlg/MK5dg/01swr8sNHf1xgB1n3nj+gFUlwlBLguh7WTT203no
DdtFTwCxYzyjCQXpwJRRKOZUCFIefYDovdfioT6JMk6Bdd2Ztu8BdrZoK5hPYQoc
J7nBjG91O2V4z2fEEjunTwtUyvFtF6Yhg1sB7+ZtiykmaAaHLyRfUjyTmBmdcmga
c40Vedmw4Xa0xMIeGFGy09v5OYzGZwsLpi/xrvueoI4O1JW1+cg6WUk6NV2dgKVu
eotYo/l1QsWbb02IEqhd+afEJB+RNv933sB9ogNb1eA8rov6nxvvqAahUu/9TeSq
OuZ0uXSE1zw/QGG+IwUeG42D8Gz4B+Mp/aWyoIO7oZYBojqysHQ7Ypr1HCj4hp0f
D20vpo/pUoaVwxKZ4EvBPIV2OU5Rkk8HmYSYMMM+aRPJRFxLOQAmsP8rGYVOqzgx
nQj/pp6stWx8DQgyQdq5VbB5lqaMXXJLyU+NCZiJ+BSbGZPGTeYfgmjIo0i7qazs
XMw+nDmzQjmnPKTJNbDCbT5dOERwGsA/9uNsM0g6AiOGhPk/+PNa8e57cY5eIsf6
EKvcRIZ+yeTuddBFqf2U0rf5ZWmujJ0s6s6QPH4AScmr2YbkGf8UuF1jOcUw6/EW
+lYFaYsLMxqIh4oPY6bvfUII40mNHIPce7apxRl0uoa2+nMygXS7llu0oOSe2xMX
JG9zsU8VCypiCifqvQAgQ/vgCc1YPzJ1Iy39JgtBqse7D9t9AdP1sAZmMm2wbZdX
w0NBKAGxjcitS8yRUH2y7SF7jKrwl+1wMXLnYuap3fDv0flviEXCQSY/g8KZEZO8
T4gF4Ah1FhrLKx0FAOnvQLhUY/7E2LY6Qk/KWQdDQZVgaBEZiiKFbdHHGOX1e514
stwKVXE03hyZ8BvDB3Ccw0a+QRsC+pfZwLe2kWBwYO0S8CLGUPB0GPeGMLQilTDn
ILCeKTUsFJMz5AG/UdeVZY1HOFSbTya3sjRW9nqM+0qX19t5NcOo1lETvgrgGmf/
Zas2bNr1KIfZ39Q0TFF8pSz6uvOvtgo81bRXWfcfVuDIa2qOtOIqBzopxldh1NSH
6qx83vW1WxRxZ2LLYx86RBVGc+skFw37t6f3+n+bCJ76PZk+zWX1Ox4lMkzW13Ii
YfcMaY9pPwPQa3tpjemDFX0ashwIOyDS1Gj4pUKIH13qyWQxE6jDgPoPgRvRTEKC
+dq/p1i6q9+WYLdhNptyPakjM/7aDveF7/fG24ZpVbYJCsd9qH0Bic0y9hJ8Z6Br
A0S+lf/loVrzrQYVYTlCx/fzwICGEil6Sb4FAddWIzT1nL3D/5V4BvYNrsGRdS1o
dORbX9FQZjpLnyNJ4Wlxxxum+8IN4Si3mWsfYfOEhVk1iZUnI6NZrRp5MnHoM3PO
6UrVdtXs0VL6QZZ1KNa29g6IM5LUmqlP+OsirSgnToDW5kiGiCFyKxPLUglwlX72
hYIm02Z5yjMb1Hlqs3eR7amIHlwThHQWN0ECvA3YCQSI5E1WeJwkkxf61uMDAT2F
neqW/7DUWeQkY9YF1qdg7RdLwoUTiwmPSrW2l1Ldd6wEvqq1W292yOW+TJ4S0SnN
1HZN0iovs9bC7NNtvHm22aw315I5QSaZb2CM5STv+Lk6ZXrmXg5+iD3wknAokmyr
NyTtRq+lER8f6/PZdNCC8DobJ+54T1RsJTnzhU1JHmJ6ER2nO8Fz77044a0e9fVk
ScVRK96YjYHsoI489e/jsurLyYRBbhIjr+nXvCWlQ2Vps2tnG5jWEyfqHUmFm+jH
/s3FpRkFcsAkjrciud6cUgLZeVRRspySj3G2TvPJbWQ7YpQVs0+MpRF56/hMhdxU
Z9jneDStKCqIW/EUf4ycrgeqpq7wARcDJPtfHDj5La7T/4qMAc7C50g+TxnnqS8o
cxMy58ifiGzR5rlzvWiyw14+qKthua1/wUEKa4Os8FtMryhBuYYydjbVcgzPcTyQ
rONomjxQUAUn2tmJP6y9bUgpw7zZSJ6rNqYKRrZ3l5yH4DwB3m6IzFtXwz1p9C8P
wLe0t4e8/bJ1pW8m6mR6O2EhHPn47tVVse6nsuSrV21A6s35hztpLv/tFBwg+B3r
XiKJ+GTbOlqwJQg0GlEocSrJB3P97oHiILqZDM9Ry7Hoc/kPbrj+M1bfMmCXDies
BrCX54DFhJANcSKX6A/MXU6FUNz7LOGVp/T7XiOicAJQ/T+OevtAAUHz7AdXp7k9
OdzygOrltppfykqagVG/q28KveipgoAkaw79XeuGXi3EjFxPX6SBZeOOBaBMaUh/
kcM4eiXS4RLpN/IefCQUrBtzUCVUKpTQngp7urRfmmqnhGkRLCp+FUnVeIihhhe3
2/8YzdODgBbmsbh7+CKnwuDLn/BYyBVaBnf96tKGjvz7WvVLNU5jTE7bDuG39n1R
JKdwEOlTGhrDhfEk9gFIHtk0E7f9rMUYudZVsAqoVxSAj5ZqB8Z1kQsVZoTIJyTQ
XvD/LArn+6OaXpQAEpQew47T4wP+KGzgeTrNh/pBr0kxGgyPe4lSgZN79JmqEChN
3ycA/2/Z8hxKbjODi8k4NnMKOlxD2M+Ayq4loVmBJbgQkObbKyb8uVTPEga+VEsK
uIEnKYMnhs5BHbCFLvmwer70znYfc1cJCR2Lzcev0xHEsdrTW6aCkF/ftQLFlRLy
/mN/cE9rJfLz5bfS/rVLpQc7BhGPKu3tYI5Uzaw578eQRg+DkSV9XG/XxrzTjQBb
+LygnpiVsAewLUl4BijpqWWh6j/TLJMLRNiLizTImUIkP5NdcDQPkLjUE3BIPb3r
hf1wvmCLtYXVbQj4VmwznGv8jUJg1wkQmt1CT004lYmE7yP0SDSPHmyFS0fYttCO
uAEREU9tZCYG5uzuYtnA0KA1+GusRkuV7T+JozC1OTURuKYOCRgnolO/pprnATzz
UP1jTczwWFETu0iTp3CiTIlVlhNqIMdWLNNSdz3OHku3FRgK9hGXFeMHCF4coKYT
n+/OVHj6T178Qvn9N7brWVwi8vYPjg+V+QEcysKBhZj4wuy2z1foKYKF2ppKycQq
PGMCOztUtNG+Fxgmz30Rs//A7UPw2uX5OXtn6cIaRfM9BmkUaqTk6JxaVksO4iJg
8M0QPzayiBwbYBp+G7K4/vBbr2OLfXCgDhIcNtorXC3oDA2In2re8urWzHbiA1Ne
hgLYDCjaX7teQ2yJQN4I+WDduuviwKtX+9WfZUiq2s0HR5jI7D5+FYdQFJnQROkD
xdb6GZ3Xl+CAa0ngwcgKDEuQFvC+KYOd0pVvxM3umeixDuz6FgqYEvqhv2pT2IUH
4fPyV+3u8Wof3jMQH6FKPKvZG1pYnyvQ36Xs5Sg0JFO7o0UqBXh5zMgafD8jz9sl
fXE2ZWXL/c0E1GkURP7K268zv99ytB7pvypXkFIqI/Oti0Aj+qqgyPWGgPW3U7dW
R9g7cBxbCm7/zKW4L4E9BnO4oIfKE5e2C5VMrgl4PVrzNSflBkLUr3dENxv85hPw
HG/eVVqtEZVYTU8DDMhrqjmpWHCPlTpPeewn4uzrxRAc6XMJ0Rfx2Co031nAgwcl
Efy3H9jGBbXATeCHZqQnUAOATmHsB9R+kXBbVxduef8zEvPpgjyC7cWlDV875gbp
rXc7LtZt7evNHn7dRMQGxaep5Y4CD+2TXmCNApjNTH/aWJkBGUz07kZQn+821Szf
NbKXtFgdT4YqwmpWppdavWBwn5ZiTf1x4+jmQz5L3nCswVUA+5ze9Dd+l4v0nGf5
lujAlshnA+dXq57k7P1+UDkrmjkNvJ6QeEWofdNiKK44sGQ99E7sCNlsSy4sTiPy
Vtypw6OnwNYmiiMnPK97mnK2vLGgyzFjU4YqNfXjrkQUqIvmofuzdviCd17QD+Cw
hjQ1T/2rV8mLyZbhdSSJA27R5ZiTYqXLDbZX48BF+2wv/XxJOMN9YyOo7m0VOyY8
My/ejpM3Pud4MYLJVOW9gKRcyI5NnizP3480z301JsoClFgmbvu1lrcayKBkJa+C
7U+iwIBTOCVvUQFIg6zyGQtPx58FWvbDhZ2vctrVZCBTi+385znwjUpJTkOIQvzY
ZqKNGovMsVxBqREw78/a+NIq/tNipIrBNv3EnkUA8aJIbHDgKGQsaH/CQs7NXXee
OLH2mYXN3vhWAc86NyMU05mBE3IN9K+KllzCwamRACY21dfNyiRxtD+ihWynYrQA
U9ayK1LFxk09a6nzuwmnDDuAa4jKAqSOaPgVlODFRahO+oCyM6/5+6zRI7B1svgZ
xXFylDhWjaWFDCwADmJDzm3SYJA8YK92puIT4Vywf9BtYT0pXsIwv2L2QW2R9tzH
RVljFGb+uDVNFCA78qk9VNc6taUdcSVK04xFHJs4v98xlKYywtaSVdiOL4oeYgYQ
9UfVSx9LsfU6jemjyv0BRcidFKVFvd+LRoBlBlHLlaKErMUoy4vWqGC0DdlNGXRC
9HC8TM7vQ8tEAh/qnBfrGsp0/ytvYHZveSQHsbysxPRUHyTRwKaLOKKyXG67DY6J
fDSWS6x3/BuAwteKkRuaR1mcW2ziiWPVwLLCSkmUr4VrmNv1ErgZffCwYjoE1dXI
ebuuehh3BJ557FhKkzLRaFPL9zR9kPBqVrtCjrklz8iPb0eEYPTTtJz3QDYTYPwK
uik+rlWcJMYOCjPhVXsjl9keLXHXkLtEn8ctoGeS8UEAPYeC20CmT/lzHsHn2RR4
vi2OnT2ysIKy6ABBuEdpT2Rq6CBHGbRO11k6oQon7/X4Lmtw0To3emn9RZdcbpi1
VcTdw3nvM21hVKYOBxNPHjGz5dmkNSbdaPQKCtIth+4UZqVTfzTA1jg+/n5EeH6b
ss1Ydc5A9S9NXwLy20+DLZhFR3Hmqp/33UUnPR5JWiwQqyASRBZuWYwvj9qkS5oR
TeItJf/FohfFHrJfjle6kHN3yk6AGxBLi2rz4icJUyLOYxAWcArzmWGUclLwdHm2
yYczOMxfYIr2OZu49xcsbvGevrFcOcF3NDkr+/ucf3vw+oqAZAxSq5KzbYJo9Gwm
DBea5LT+pRV5P3RpxDrYumbihwDsUc/sbWXH+nXVKxaCTFjsC/CtE6Uyzwx14p1M
fZ08I13JJL9DrRuSY6fqKcmHoECO9CL9yrCFij3vrjAMzed49ead/NbZoSJCDEbl
KkeL6Rv+t5Gj+sSQKmfGjtA52JAtSnouR3wcQGs5xuT1MBupRVmmdbL406CK9CtU
S0p/NhVq/JsSAJDmtodTGalGDo2NilMHwTXiQqR0yRI9ZYaJTnUFwsSQFCr0NfZ9
bexo+e8QAqF8N0mvR9plyaP7Szd/2N/mmbmyt7LYGSPx0d6HYQYYgtjPt2XqcM3y
+0FfWy0BB8+VuuBfkP19ASGZbvAjX9h4mdF86VTM04SoDW8ovjIhA9FG/91abLw7
4zYlQ9uQz98F+yVNUQ9GrbsSEye60aQZu1SWJ6Fp9aWNcMaH2Ww1gF4KtnvAWQCr
KsQNSb1iDe0V8tGqAMGLhB9OjzJbidPc4JQi9+APMIc7thVd1282iIGuWtNeOXLA
mb2WqfP75mvqXfo/MBjVzi17JPEdOUs4D//5HKnlhJAfjF0Dn6R0s40My1oLP9yy
k5mHrgBhaTEd/xuPaX1JCHEMsdw1zNR1QR4rVkGr/0/N93LzqlCtoVJlcZ/aYETt
s+I53UwhaPdeT2rkucd31K+CEaAEkcDEGYQBSk0MhWSMZVdY8kc8deehW11R/oVU
qpUxi07IS0KgJA6rHwoCsFQImXOcSazz9nJIYLzg6dHlf7+DoPALPvPQs+JI0SGL
2T3kQuH4GGDum6rG4Ys1YIaIDUtOawaMbaRzDXDqWPdEMzPNA3BDNiPrXsnLIKyL
3lfpPmxXssmPD9O6bMqmjgYwV1CdWTNZCUr/v9wTV8A9lpBcIJLVdRa7M/HC2yUS
inQp1Q+sdQUHkEiYeA4QUIjnvgpE25R0+u+UQFujjs33fk9DkQ6DcdWfX1C2p3Eq
WSWBXyv9Zhk+6GZ0y3rSMXyd5JPnS3aFPkg06OXlbUOjKJ1PM7xDrb8q6mwsxsLu
CS1TgOqIoe5PsTOaF8kSGMou/xOywmZiAQtUKIupP+BcjiM82/SRM6mGoejeW92D
3ue7VOP1ZRS7CngxBs1nx4safdr4BJ3zHWQPoYTy1z24n1TolCBosiwxYKLugsEo
ETOc/GZvEsuglCOL0y53wKMGnZUdmQl8vpfCn1Hg/G8FnlZ9a8D03SRopT3KRLmP
MP+HMLGk7r5jgmiUGf04Xv7PuUfh0XrqWlGEZo+oUEw8EmGVGgbpjDUwbrcv03IX
JWae22EeV2LMhvl28PGv/N5ePfwS+M6MdJs6FfWOANiNQI/owFEIqmszQ9AgpxOa
GzXpkBddeocZQDN/l6PSyc7fFT7/dp3EjAIC97Z/KRTPbauZ0WzkKQNtIkH5eWbq
0LAM67DKr/1JXUFzqxRe53iYRhkF0uz4ugbzgCXr6x3uLyp82xr6M6GS4qYzCFFR
b3Gaxght6s6HhoqeRj7mYsWGyPr+Pl46LsSqWTAFkzC82YrU4orgvp7Q4BVmNMdS
HMp4FbEMLezaH8hpLpbXVvMNeva8hOFYV9lU/xQy7mpEiebrr4RfBMWHhSH4CAfl
vwO95jg4+QPiqmwXRJra2c73ohKqmOBFd9Arp4Q+TXnzmTzRsh7Tb9AcKaEuAEco
XBP9HYPGM5qfvaqbflIvrgz2yb1PJujJj85lTHjKL3K24mmD/qJEXiNiUg3Nyo0k
ajhm5d9xscXk0ZGj230n8aguRC/O+F5YmYOeKzqDf9fcI/r3i4q8Jch+2FEPmQGw
uo/xQGgDN9MdwbFT2k4/mAVzwI+hWAbvRnhWAFaggiFE51zFUGMnYcI6va08j1Y9
h2BaQLjGnJeIEqbY61bC7QoNBhCODJhoD+zeivHtDRLbYohuIPKcezxYRlxKEkQn
gotfJmBGqrDQckK0rjOzXEIPv6R0qP7TzCe+vQHho2qedr6IogE0i27nbycZy65k
Ic+NhBows03cAtBDFcDuAL6eeAjjkBy8yz442Z9CKocZoVyLMZ33jI2/VzgjyQST
MATy7sjfrAWTtqKivLdptF/jviYTXP69qfOUM+mfddrRKxmL7ybH8QrraZ/HMIax
cZ+MTe8JXP1yACYCoIoUaALkKccGrcaITF5cAtheCrsycXzbqcpYa4nhWrp23iNv
s2dhPtQMWiyJzUNFwupebewDcWuX9E85Kjb/0HuxzIufRueYVy+mWk2Qt+RK3sZO
FtePBGo+YIBxen2nHIPR8K64G1MkiSm7hhppeHPSKXKWgmLp1yEGDQtR5/3AYiAA
IuPWl43zI2WaQsu86DcRufp+ezvXVpwOYgW43W25bTcUgdLTTqwfYSsWXkWp6P2V
Da+BFwBapafOYHDpL9WOEtSTdPgX1/Bjh4MuiKkozenZ9YWtMel+s5mRZfIrhGxg
rtQS5+9rINmg9VUCl4yZ1ec+yvO6wmtCx/tXSSkWA9QOuLtYJAr9VqyfR8LzXRGy
0fWHyMnBjzY4MMWXsZKNhxS7UIpzjnF+VctiWPki7fa31yi2ZEoVJShoSlHVLNfJ
Mp86jZh6zOxXsjac5siH+gpV9JNoO6InpUDLCXXiP/qG/+WNuQBhh0caqEQ0knY3
Kn84rnTW88uZ0L8ProVCM8ij3m1hgu3KDOEp8Z1HUz9G/JUmW1LdN4jvi9LcjO/5
svIMK1S9QI8e03AkTjMDoFb57VcM6+MAbT22wAIbtfVuot3Te5N8e9ZraLHaz/yU
EPLAQZyagScB2P5H0TfYEPav8zlkSb5zNBqbHjxvUaelYpLcHOVugzZtwBZaBUOT
TsrcDtn6vX7RVCLNrzI9YjJgyBB6Vx5U9TT/WfDv6wvo6c5MBtqjDi70rwPLDqHN
Aq4K6QWd7bbDO9D+C6RP43UfL/lFjNhfu9CEfRtlvrE6bRlnKPEENx0Ug64w4Hbs
Sw15T+xiDm+bvErOEiUG2bjVToktJej1hGzkz1LYNSkir3FakvAXItIewTXvVxG7
tJ/lcx9FIJl+WFrNHQsTNMHsMXwzP4Wf8lRG51HXXECONTGl8veq19ZK+/5hIlY8
B1kDhMpWqrx+kOq0zsEv51VmiTD3BLFQpGmX5YifWhdfRHIkUwcRX8DQPv+AdQc1
ZR7WQt4n2fwdFKWyd0AQXNzGLN2RbSPjT2lfWLDYV9ZCtpYL2k+bgbVP54hAzyaj
55X16Nu5681rPCLnBbhaX9kI/OYsQKNledH1m9sQOCtIT17NnskgKUy7bMpiOpwM
CRhdYtj5xRFgHA3H0wE88JwepvS1QJu9tNAtxjd7HTUXRD6gWXER3reSTLysP3JT
iL+JR6oBj87KGkcdtTXn8IZnQWf2FFBASBWm2Lqqz5B9sX9jaUroEXzqIAJkza72
6hEr0a9MAdG5HiKSeDS+U3zE78FCbc81cNG4Bs/HWXxr8AXffj8CJ+LD234mDTON
JgN0bqB09BFspEufln27BjLmxsb2j5Hj7+JkaK3wVcGMCSZ9hgiC2TIz7Gn1hslf
HFJGDVqTHfllcCIVwz8gWoDkxiNU6+FXw/PtKlQT5hBW1eAKqVnDOLyF52vXOVnN
boB4I1Wb/hIJlBo9wHHB/nm7nMPSpKjWqzOpFLsTTQyr6sogXmI1+9x2WKU0tv8o
IN6ia3I3B1EZ+Cb/ltLHDYgHAd8WSGuNHy7J1QkfK4HqFH+x9K+bdSQ6reSLZ4zy
bVfstm9gb38fqvWGhi00vJyYumjYgXFWlID93thMCD14Edr9HZDYYl5/B5NzjA7+
C+eFCXq8v7iP7CypYMdFI8BA0Ho3w4nyrsRPEsj3lodzr4NfI1k5mC8hbykUMQ95
uBSz3Gw1rTSlYWCVzv7d7URBGpXo/Q8nJuLppcuH9nylS9ejISkpXfZH6ndjwbp+
+qGBKzuLf3hbjNlV68TuiQloI4q6rcRwdVBG0LZomrzZ9V4MX4AuVB+ciD/vu3hX
kIZrtebAzOGvpsbGpDWj7ABP3bKkIe+IVxQEdS5r4jogsbhbQW2LojYdsilFlVFg
ZOPhhYpa2cMKUnuYsKdIretdBB4ETOtLmdilqPryK0vnhj+FHn1sOjcqWnEpL8Ie
BQ5LszprdFPvZnSt1RFBYxbxjLedWYsYWpNOONuJbnli5GxaHtZhYAVB0Lw35iy/
hdzpi86MP9rnaKihCRrYx2otzbNc/GjkvhGcfDRrK9IfMC8+HB/Dz9CJ9UrZ3HLs
ie3Pt1LMvrmqLErY/j9AfWR9cTF4oU3oGG1dExfj8KoFxeA8+AqyZvDS1+yYClEG
PPrdDKtl/ZdaPagowPYk/18VzDwJmnnQOPy2s7OsW2ErUNk6XA41lMKLsJkaWj49
1OViOY8P0a4P7DcCxryCzpld2b5UlFdu9o1nm1qrkm1IrjN7Kd3iGcWdspxgqiWc
sjr9PPhQRb2EprYV/uMZYRdVglFDK2CVJEuUO/q343caroaNGAui7rIkjCXDX6sZ
LnAVgns+cfxpyBaC74+4c8LA32eAbUvrzfooqcrRhO+EcXV8ucofrYE39bjJmMPq
A2KhGen2mtTV/jjkzDr4rxM4l2Su0Z9JalgglAlL6RJfRX188efM9wnJfFzR1w/Q
IO6Ar6Si7l+Dq1JCBdmcoCg8cyZzByCyuIClAZ7kKR7N/jJJvYI3h0J3dFXQ0acJ
KkSl3TUAzncNRGVCG2QGkrrAqYsvYp2EBFI/WZGCCzDNUCeQF0l0ElRwKzCE/SOp
sPRUj4SvuB6RpKk+eFLmKq+KycqMEg9SbppIMTuZgojn7KrRPh497HtLSoNXY6g+
RVaE3jUOzUCRuV/9Snf+qH0hV053+i3vloHlTXtsC/gl/ZfWnmk2Su1HF7FpqlOp
sSAqAOLH33eHdpZtrnsaxobeHBdSyt0ZL/wtXUSbNZlKmdIxg9qe+wmYINCu6zuz
gWQboNWzpoJA1VMrhqUI4GcyLr5Z9qc0TtRNUOZRQ9RFqmxIhexWWpzNHwXxmReT
6DV5Qq43hhdWabF63vKUKPPlDUJEhVrIZkp3dadk5+68Fiy91vqCxkdMMg8Q/d1n
V5yms7sts1p7Ccf4HhGXfM7vFobFrCspNxWYK50CDMwc34n4JHag5WL3Fe55QPpQ
K1pEMiR0yM7w315El8Xd6hRIZ+wsyTGvmFkI4/SIDqtfY/EDgUOe3byvYfVTmybz
1tvMsQ5v9HgDzhk4D7Iu3wPfWDsX/mIwclrXAlHwSf5w+pu4cyXj1wtgbEzkYSxS
eD9mkdT1losEewWf+7JFDmWJm5X0JomHS0l4YUPwou5ReV4DHnlm9rb5br1jpMBD
JH2ZIOG1JeMwFbH60AD9Wy8PB/3s4rQrtcdkpA+H3tR33C/yu6Of8LWEkSyOqCwQ
qinENvTONc/DecVzcl3PBU5zU1yLG7j8lVuSjNBL4J5f2AOhB6ciA6p/gSSmeV5x
BXowm60yTHufXcZBkXb0DapU3V85/HjYVnjy8RzZXVymr3E2ZqOdCdUODmP8s51j
U4LUsck9N8/tCdcw8mvBHexbvb5fh4XL09U4nMcAeiDtzzOieeT5k8lZWqjFI0vp
o6l+hJ9F2fl1jmfBLq8NzYBEWnERntxV2PoOu7Jj3xPwlFZwtBjmLcMLcy/xZwTx
FTOxZ773woZ+ilOKG95yIpwpAix624naOs8lfmBh87fvE7Ut2hA1pADN1+PrLAnW
XQdgxeAQ7t15GFaZPrp3uVENys0biPQXTB5OproqtE2ecvaYjM3xH3mPSUG6k5kz
6DWeL/mD3XmHqj2xvmX1CYJ+Cgs9J8AOkoROzKJLYxYLMk2v4Rx4RupHodc0+x5X
RMwqgZkd+l0hcJyemHkj7aDI0lHlVCZ3t7TXFVD8Nx1W8MISPyvWZ/Tx3mpYwvoF
ZXpgaNYm0w51RQzoDJ6S414VDJu/KEjs9EXZssp3iWEkTveC321A9IG5V0gOywnD
z1kMLmjKW9XssGF3FjzAT7KC97ZzNaaGqeRnCJSQGnFh9Ed+s3KnA/nT/RhoZSnC
gtXjuif7CftEU10f8UCSgOgXwWlQmNrciS4cJFbZdGLFhmyZJnVA3wdXB0r4KHOr
FjzObxJ5oOkgcc5pTAHjYO4Kx14ABX+perqW56w8UfWroFfPfWsdXgqUMk27xEPi
fB1nATDoyE/nS5iQQNgY2wStyBroylrgyMp7GgA/CMKy9iLy5ETTnqjn8ez6sdAb
OKzZxE+6dgsZDgmSXcrnaf0Z8UAbup/SIqRxHuNhLcLOwbkN71Efyz8sNJhIXGR0
74Br+3vJ1yLv5w1UoDWgBeoc3B26aLrhJqzl4ZITVliUGcVf8u2XTrsW3JIwbV6n
NOg5iRa37YYkt1fjyZqrbrrtSMbk9KieycEfLQ54+UPGVc9ZAg4EBXqZFdm5Vjzc
Cj8Eg5jaLE8uuheGEoDVLaV8fsnx+UgOclcgMmQZ0Hz21T7A4wTqhuvdXG5ekkpX
JoW6sPV3eWNpzKSZhFASaNGUR9tfpSY7t5xXcK5D7Tmtg5p8BxVsdso0lHOor2pP
kEc+O2eCJYxSTHtBliyaMr8bebwzlgcoqISQyjBo/7UtbeagjqXLu3t9FY+hykq3
0wsipg+NZy1TZ1trnnznE1I6ycHddf6rMDK1ZrcOxgiRBAnE8AVRdFog9L462WAS
7k14yagG3FDjiKYnPKF4maAZeyAHpFqE3ZTxEhW/IsaKuJRC/nXfKwekrRG9rYRV
+fR3IQDTZF9bsEpxZFbwKOrYePCm7fcMXnzzOOj5CcP5fmPt7Q7U1/DiC17mxcyo
8U+PoXtW7EzksYDUC36Y+4aqymvC9SIsPWMX87KLhfoPMrSIKirl1tRFpRUtvn0b
dS7TFYSkDcooinxCAK6+/ujMHytLiJtXp97556PzzWiyQeuYNstpT9L57RWt83o3
laMlxIiOJjAoEUNaOxFtpyazPU6BznDOwSO8WMtEQcQux43ISG8y3IYQkmEzV2wM
qZaYCdi58VpJtmdu5CkzYF20fWk5fgsdT3iNXUcSYHhfPRrOHHO5FMgf/SfAU/OZ
md1RHDRjY7lYuSAPQigF86CTXx2CmLsM97sxraoPQO5hpIFtL2WDvkdus5YrmqP/
evnnecWCH2/cNNjJZEh+cIX7cRetPwM5kcK+sTURCpA+ty+0Hy/16YKsvuqWVJ3N
pmAViasQgebNqPADiiYJkryUSNV5PDzAsJqj2yGu4zybvv1A2xh6wusa0lPlc6KV
Hbrhz4Exs8LvHglBa2U5GCqOIOOjz9K+9jf1Xe6BrFcaXvPHectLMGVstZ0o4Pka
o7UPsYbcUW2UgpFpHWkSfgEGJ3lxnuzYy+aLiqdU6isx6FS/HCNar1id95suvFxr
AS1+O2QpdISZbcuPSEZjKIf7FPJQ7bg4VGp6hOTSjcGrnvBRd+qj1GUTE3OWgk+u
AEFaUv5eZQCFfipW26G9HnsW+oPjSuV2RRqXfP8mTw/wSlO5CyB9YvFBhCkugc+W
JZIgaSY9wnlDBt2x22C88z6EvtwxqxJP0tQO9eebnaN4aOeOgHpqvuMsrWuXmV//
VXWfC6i9hpBANv9pH1lxexPK9TXQrZgg5hm2HxSJLZTjW4jaWKreVXP09eWfFizm
Zunw4uxreQbwY7eChTmhQ+Xyx6NsfnjoVRSPnr75+TKwaXcTDUGPBxxzqUEaYdoG
UDSDiB/5uoIdEjDKanuGFhK4oJVyByAZfl+O5Q4573SLvcghJYYl+QpoEvhSz9MD
s8St3cVLpAamNOIADNA8nIH3lyb/8SfjBS/JFWRaZiFLE8k/uMIAKi9ryNgID07E
gPuY/FjsIWxCv5gh+88rA26zhT6t0j+Hiyqn/D7Xu+9egui+ZgkAVzNUjW6N3cx4
K/3KAJkJpnDUuU7PSZVH9fhPPQfToGpYKU6PWQhBLoAPLk5LZHpiEBeRDqZAQiNM
fvVgJFk07T0YYwru6p+q68T72AeZk3Awn5zpAeaY7NPFXUX2+az7Md17jnpqiKiv
J0KoSQki1FCrWdpM6r8RCZ/YbeQFQwfIuYY4miQsIMACynOAyEj7COqWzLhz84K4
O4RCFvKmNO5/fKr8DUbPZZicmiNmmh7XYED7u62ziWpIm7LFg3OLQU5dFrTy0ehk
i70DKwhstEYE8EymExYqt2g+L0U3UaRD57Yelr6MlUbk5oiSJr43NB3i9/M0xEdQ
z6os8AtwHJ/tMuiHpdUOegfdgSyN3twaA1ELxTs+392wO+4tVaWYGnuttmELIMZu
YIR4eCFblgLEWhAoRgsISu5CwSIZaoUHZPKXtMZ1b7JDw8XhQ9iz1Hje4+N4AuEj
VPIi0Fe+rC4DOtCADKgCoKx9utqObFGoU/gBLNgPS6mFY779pnKI6GceY8mUWqqr
CArf4hNBXmTQNDYDGvgxBkNWpPNYiQsKw9s9G016CzrajEYybtTMQTaJEXl6B5tz
LjcnXT2S9NlLfbSrfnjVgg9cGRrq4v6PPN0DSHanWCa8ZktKVM/FMOLIwIwUAxpH
6PnWGY/FLGhWlwXx8yZNZMXfhKfIgPcWuF0EI+10svM/kxGYndoqgOJRU+jK+AX3
KK+AdEqqnoFzeLfVASjfaGmGCuQ576vqPIWm+5bArGz9CDVv2EZz37LdrX2qJevH
pq+rkb+B3qoxscdTswpoSUpVrTBaVUQ7UQPYNv/Y7i2tCAJlD3zYOqJxTohfBOtC
cQTKnpbyEJ1aMz0ruJHy8E4iO+mlIc3dVr7va4p8+qYE90dXnT+J7yQgXhbrHewA
sVe+cl/bfmJoT2EUB7rco/d17JOp1i7qCMd97unLnm9ZfsMkpD6qMwqgZGSiSSDs
Dr4fmgP9wGgfJbp97KxmKN/7yXpciiZMHC9YYpL/NnMdDqI5mDxnnWDYuK57Grhf
u8cthJyWRvuFCe6/wefAw9QS4rKtu/nlaJo1wSSC+bVoJWqQfrB7WNlX9yCyeY3X
jsKhwqX9dl4oXbi10FfubB/n5mrK6T/Ocv/VlgXQvObN02SqrYuEIXhjn8qGoizC
pFmBEzDpFk4wt55eCk4rha1D5Dipt/2Xjg6F/cTEDgWGuepDhK/tY5+OASOTjzKo
EAqP3w735qC+wg+IZTn/vwbY7jl2W9bGQWM4Bbr5hpc+TLBAHAavuTcPQysxPN40
eN6iAcjuafIoHFoJ6Y24b3B2dPFklvut84awWjybe4eeP+87UTjO2rEWZpvPjUmk
Rc01Wl/kdby19I0msn/uH9vG4T1LGPAUtsEoxPF7CFENfdOBFZ7DYoWI96tgude/
hGQvg7XUX50P46XnQRB0vtra0db6v85YdicDXFsBwnQR2WJdfIQk9P6L/aj1xQ/7
izJPmWAIjzNC//UTrHCrrdWAczjB8GnAyGom7Di4NmF2LG0Eq9ovvr95S4NeWyCE
zMTq8UzkN1iuo88l2ye6PvC+1dDAtsachbX7+dezy+yriFybXdYMwMrtS1/VdQ7E
U6+WKxGruhgW9cqQGbKuJalHCPGcqgaWsgL80QZE2rgh/W4ksS+kVSgs9oEfTBeD
fNzKQAx/N4Q404aamGeyuLgrGWIxyOk4xzNPyT79vAeyFwlBrR5Vf3zhGoE39z6Y
nQM7J298JzRbYoym6do3zr56y6p4ErZr2T9B2ABY2uPx3pnXOkmNRBrIPuSNB5C2
EHvNGOhQElLv+OV9HYE9NGgR3Tct5QtVFPRxV67/xhBVrLRrpL5hjdR6t1iRXZ/T
keTWaZL6XbGprynbBI6w8eQST+Aw1fviNthIMWdTDIaI8tKkfyRa4B5eipvycO6a
dPqJEZAB24OScDm5O/+Tl0fqCuZH+6m9NgDj3vp/otge7TfoRckyq5hs/xKlsXKR
YEDdsXTp5NFdiB5UCXYU7P4Dd8tAk1zmz9yiRlE7w2VdZz0g5rT9COCWFUVD+biX
XcWfujcV47aEXWU6m9wEusLFNVcY0UYp4ZFWJAuPHvog+Md8hvn6oLR91C1aPgV5
1Iz8ipF88OLGEv19JkOl5KRuyVL17whN1fEfivRSY9YFjw3GqzNu4PU/2Fewp6fX
wKHB8AZ5krhfFj8kSGvuIhwVbYKW9eeIJlrysSIYs+fjgNXAbTYEFkURwQEIgjHY
D5qyCWn/6SpEYVAVHEavgv0gcNbuup+d7jLJPFqtEqPiUHaDtNAvrb1dHvTJLAcL
lYEmZKUJ7E8uDqCOjKfvmbyBcu7rmpYWsuaIobjBsvuSKDfp3ep5KBkkZ2zn9gMe
QeG56QUXcbTJxHbAZdYwKldMOsjIAihzN7RH7qKtKa8dwN1jnp7dz0FZgGR6xN1Y
43sLGY4u7SzfGxiG+1WwoGWkFghztxVDDRCrPCD57lNq/Ew6UlT0DI65qm0CiRzk
oPTstOSm2htNEr0q5DKenD5jhKteuCt7UETMzs3ZqUrA/7R8vPeEaFoHsFlDLHgm
cUcjEBWf3K4c7uuV5lJKtBl0Ul8asFIThK7G0T6RU04jJ2DeRD7c4IVGhsCG9vNz
V5h+VPljtt0Bbu0yLuzHDCYhP/nf2GfQR/tjX/6kDHzZBl+TBET3ToUlvbxZhAOw
dsM9xqrS9sZ6IZYAPPpQIwJ5QI/9SFEaObtd/FPAVIUNgqHRpEpKXSGmL/bwCf4v
ds1wa30rcghuaEn9vhXQ/Lhdn9ThMIXqQqmZBqTELTv1h8egfwX/D/8akgE4xH+N
7euQjZiWcJ3y9FF3Ofgk40KNrLcKYxNraSa+F6Ek9iQ7gpn4aJy3fex4pVWgxF9X
Ja8A4UFlyp8fUE+a5l2OTsWolblnpgbqnOXEoYFhDciiXEITU4r8ESoSo9FJvpsk
i3+YORHH63E+fPX5Ic/rwFJyn+9l2XFBUo52D8u9QQzm9NGCY+8t0hj0/5fl/+bu
2/kVhErViP0sp7iITkNX/QWxFPcTaLm2jcgXh0dEXvqTNeTgdxTRV9S7cVRDgmST
HMdi7fEaSbfz3HpUzacc2gR562IZ+Wc3oeymQ2XTfqjh/6WxQ1qg2xERpZSZhQV1
FMAyhNSrzdX7Y//Gqr0O0qS2f3hYcOww4NAk2SKr6NdQ/2P/9MFtYu4oi/rMFv+L
f+LOvV7TtpJY07vZAhI72hd6mkHZmFrmB2g0Qr7U2igSFldcHBY0iS9QLwYTecYk
OvL6ZqqaWYMebEeeTJD617QgA5Ex+D/7rVrEx9VzHKt0ldVXj/iklmUktltP0sCG
/mzaTVVwN9LtZwnDVQKCo/DF2p8lhXsfNp56JcxQoTpyEg4ipJI7Y9AGCjEL91nJ
kdzVbpf/D//ENNEV7JRLsDyRg2C6j3yRDDccqHTxTnN1+HmseciNvsVUl0SpnuST
XxMhjE19J4GT9Vw9NloHIeg5AS87VZ94LIZA080NWmGMZ1UKxk0RH2CjvSbuoosY
Ng6WLr+E4eVAKKPIQwzxwJFJWOvqvLlbdYlNjGwd7hn7NasJ6z+JA3zQx4KtpCoL
nH5NcBZwauzBK/gatoufpnAqZlK2bfE5cNmy/6h87vRG899EsgC6SVEqTSCOFOSZ
sXfFsqqNvl1UT7NWqwfClX+CO3XS9PxxcATEuv0bsZ5dyEhRYiQFfRdKqEBIIFDt
D0dKP+xmAkHDdLcq5QmzCkQRWHT8YTw/Z6ktBhSHBTMAphmM/2HypEkPy+wrfHQz
QMiv6m6r40nsY8aEQPuTGHn/+e9Mb+zbIQYbLqYhpCeND8E+Vqvc+xp6qhC7HOby
atvxbuLDar7lIgmSHN1s/JcklTfMgZCPTMk3zepocfUv/6zPNpzdFdNk6iy4kitc
Umc2FEY7VMeUOVnmQQUaplZ7Vhfnuqq56ejsS2aI5n090BSodJ5OFYr9VqsEECdH
dxvFS6M4rWRs+kGlOyq+8UMvjLP11EmZf35Z4eeAiopOKSa7Uwb7Ru53WDwwgKbB
/JQ+vZ5K/BcpKfpfqqkaXC0jwHPsiQ10UfiX434FBoz4g/GN8nToOWAju09f8SJ5
fVXtWiZqkxd3fRbIO/w5rhSq/S758XyzOP4Wfc08siQyu0cHLpjEXd2fRhRWb8qa
b3l8o3fv7zmRx+rx8vFQweiszfRqNsusEgPHXhlcesT4FgpW2GhLmmetOv0WvDLy
Cn/Hw2V0zZqBoLWQH3nA//jkLLLMNJbVVeFqjTsbDhxJW1kYZibs07Z8Ay+mp9ZR
OunKIllryB7pisrl2L8AmIauTaVmmVbAxgAcq90vlQuwB4wmPNvINJLoFYc253+L
IcPhcqkBOHAZDh9xfWzOdgHMcvSkS2B0U1f/lr68bnwviWgqvU3W+8+tt6xZALB2
SIXVtvPn6kJemWS0LVeq6I9//xwQ+H+KL+Nh+gxIhASxrwJXDHKhSyGFRUXSN3HT
p3Yjtc/ILBCrJPJpZGED8fS8jG1tQ2gRB43JAltXVVIuPSlm4W0gAt02RJp2blJs
nnJqD69/S8Y6P9FobADACZ6fx3r2kJqMv2HOLmJWf0hGfuIj5lxqrrd5MZR+hOzw
TGfNqUi8gI+vDE+i2TJEcQjFBPkmkXTTH3XJ7/n0Y6EY+NmFvKJs5piDGi/rdryC
muAThqsDUrOCdkg8ut7fsbrAHMhy316SYbojUDstBkrLifmo3Sq3GbdxPQqAm8NT
ZemFCaM2nilkDvTUDXTgki5kt/vAhOXT6nmVmicoJO2cr5PJ4GKDVY5Uzjg3IW7P
3Eh3uPtAb6YUuBN2MFVjKDjn+0ISc1d23QnUIUBAIIdPXBIYpL6wvhgArgi6swEE
6hk2hk0hZS4aRltKWu5ISGQHKZX1C4TAN2dUTGfkUnrQknWXl5neM803IFAbxciP
mLUxRfjCx8KBf7x3hn0HXCIRyz6Xr8bPmpbpPrZh7WwIJP4PZoCihAZcRVMFlIs/
/15wvyhOTByxGbaC/0S3PV3Q85q49P8jisCuQ8W+GQdQvZnpfR1zsJXgXZJLQFwH
kOWwSC/1YYAVIkEbhSQj081nmbYitkbB/kEtZTd+nVhjCYCT59mwlL4LU6UT1nTm
3Yt9knZGMNny7//GLxigmd7HdDPf457tXbItIuFpuX/t1zHDCLt/HeFDArfWed2K
FvfLbzRYduWAPEn9L0Y2OCFxSr0ei/zWZcEs8nQmoB8hlGyb4jATd7Qw5wBD9Su6
4Hs4KiILLqna+x0a6i1LiGUHTh4l86yeX0CqazLdDHoFwt6VJsextXVuGXnxjELn
18UQJbhAJ++z6m7KB07CQbux5g/k4yyc9ZrBLTl1Vfl3vRQORINhkZT5TsahS6RM
lmXyxwVkRlYzXVKA81ljydrOGc4KM72Fax5rdZetYsnyzZtOUQiI80GzlGlf07z0
5rVOk6Z2LRTMZhVYW1WlFckJ2JYrQ4AON6HeavVYQHWHmwoPXT4hSH8zhTbrwecz
arnP8dY6isVTpI7YzoZbNheEHQ4AnFENCkbXkOg22jQmS02DX964mypRkVl6JvBz
eRObWDlBu/48ytIVNUM/qlztJxmGfA8+g2/Vv79FHkyTuyhyJiVINtJ3EWQUWZcM
uFpN0SDAtK5NzVAM3HK1/wl7hAkEmFRQujiu41N5NmXpeL07DCCsgA3yP1+eUZsw
cKR201ETIhodhFTy9sbqr/N5XLGDMNam4/fnVpxYUQ10FC+MvoedPN0HJioXRxne
SHSz4ydp1/HScfL+3QmW4ObUCkko5WqKqgvu/TgRWpVcDXffoCpr/aF6NFNAIRNV
RQ6/zZGXE+0WfvEwoS8e/oz5D7NmF9OTxHl+MF+1SHpr4+LTh2OTxCEyg8lTWkci
OyEu5yL1PrXWbPASQ7rZrdsv6PCtDzUK/9JiyUl3nr3rg/lQCKqM3JH8xJxA6r1M
Au4jGKvhdI1zdDVDrBMdJz4v49zfsikX9IplJDTasLq4lHWzkDnu4OluB5qBQeep
aA6Qxms5aoh8wykV6Y47SU7PeH8m0RiQfX7eo7hzNX+zXRV3XD7jlRqY+42Jyeb0
qmHCMgji4xApU3Sjf7o6rQ7uEtZQBW52CpNzcG/+OFooYpRcJFYwudzCOMZHF+tb
E3qsypIW4rOyTLHmdwE/l7VYnr322DT6BoM/v5vrJnn0fkZxRrBtZeJfvm8A6hoz
mSA/OmCsrnYs98IKuBZtVx6DZB6iJcj9GfI6bUBkO9msN6k9rVyfEkYxMVmzsnYX
MOJPRVd/lk1Y+08cur1GcCLYXe+EYnPOcBYKkqGLYWzAWwng2yt9hoBakXyAH1sS
IC5io38tWh+Xdi1RaQQTYtzwxrOaEUdRqx1fP0g9r2vcN84lx+jbGWSzOHWp174h
uBQXrU+YGO0FfufxyfboHhPKywlYuqviSAkLZ5RNweUeNv0LENmXsbdcO1M2A2YX
OCT72SXgV40WME/8CqEEPBwFNSPGd9kwrprhgjbE8eavN/zDnDnKaL4NAzDzQVer
wrfR14AjR5n9SvPklZrNv5S7DpgE1eK3/Z20nPfLCJjQnGlOFmZPF3NnsKvSzoGA
79F9Nq8gopKnGod9p7d1i1I8LFc9qRHTiAd1AHMiCqbrmhoa9/3gA5VyrsrWyfkt
kVhZVFMuvxy1IyyT+hWBgfdzB/wn69r4GGS1pyCifRpnsGja2J9bCwhGRSirza8t
NSRSA7is2CnEdHB3HZA356YFhrkU34xYW4miAtbwuMRunkJkRFqKyfqlGHVho0W0
lPPOzPo90m9V9kJCb+ndm3vnalSjoBu8ODrBXwARvTzB7qeqef8/Vn8ZbY9GVhJA
L5/xob0W1+B2v6f4VAlw7SiJfDvIkUocLNBgtyXu9b0vAfUYX26Uv8U2zb3fFBPx
ffhmJik/RCRIsldc1He68liiPg0uHCdqApMKOSBf7JizBPlrvB+MDPsS6NQFzib7
n+g/RnIvAiiw7rCdcjIpRTHIUFcc1zt/+qu2+rw6KTuOSYuFAllz/UNn25mRwdEs
zzUfffwPmBcVLYTGThXVFkdjBrMLfgWOAk0OGRWErNYLiOz8/VeiAdPGtIADoUuK
RhNJl9USKTqMXvYc7xz15VRK/jNHhLAnXq9nMlTbuW05t/XPpbCikFLPPdnrGcrk
LuY0AUd/r3wd9sQEZJCNcJS5dUaTxAvFQOQFXWxMWJtomOTtWINHaS3XCBBAuYyS
FWb4er6GXKJvnMZglqsrd4cnTzRdyQ+JiJbkCBOm26FA2fkncMjcb8vpUXMIH2l5
kzPKhGlT2sRwelKtLIN+dTZjg/NESDmpoL4zLq+bnFYBY3oSYkGv9E5r+iXJhaEB
d9/QcB15QIB+bHPKsS9lQtUQnjpXaEn70vw8A+Q1MirsRc3J1yUiQ14jvDJKt3wi
LdcmKfJbctMjPRiP83Th1TBfuExbL2+apHUQKYvgfb5n2Gcvv+dB6uyjaDpPw62Y
PIMhZ+BjvvrZyKOmVhsE7NSa6/lmY/JsIXMLmqoyufuUJkFnMUSqQa0W7pgdKAdr
tRF8v6niAKvEjx8UeJY8aQduVPPwwbAM/6OeQ4oJGMtfVXXGXenTaXm6hTAzFcGa
8Eeemy1R2PXEBMn0947eZX/MdZ34U1YplAkyYjrtFtECyJ96QhIZ5DJfqxa0RzcV
zK3ZRSoF5UmWmvgVILEKiG255NGwg8mwWvYzNJapvCSfx2wdPmgUiqLcD1xI/Hs2
YUoAu/ZfdHO+/PC/Tyk9SzF1WwUfg0XitmIVA/YaU2XxTBcBWjfCn9Q3IMcb1rrh
V/hF0mqwR3A3/rRsFMhjCfg+eVl4plwufBw1Gpb8Ehfl9DyKqfwjl8B10r9OcfTa
CDLTkCPFFDnsAVjvHUcjU+BENz3VP4Lmh+xOWtq/M+PtI+D10P+1GaU2HkcNhHKe
0ZEc8LE4yzNdBHD+Mem9ukNXRX8qaO8KH1sm4wUNCvUSMVEAEz4fGayU0uUhZ79S
mgqc+SQP6i7HI+J72PVeWj5EKl+pz7gvg25GqnIqcc1by9e3PUxYIt6BSvr0HNMD
73zJqFdDiUGnQhLD71tBnTX2lpyycDxD6OosaHTbTJLSWlWOAxoobDqS6UoltfJt
325GNqTx4Oo/NFT53O5ga5sGpmdaZBN/gLtdTW7pOzlgw2aipNbA1S+kmTwPSG04
RHozARdedry8YnaFojcjWX13x4wmVpauOAyk2OhoH473MeNyv3Dz7FOtO/fiKCZa
Z24TUv+KSSvCOmxfbyI6tC7d1vK/2cd7zZOHZd/Qtv4e8rCFObX5s0rUUB23LYyp
YfFUMtHks2wNRbWoYECH32cnxleRgWk0eBe0bbGcN52WID7nVJ4HqZElJDIAH/Yq
tQn9RXE7hDLohiU5fRYYKcSpAaSHtsKA8oMqoGTuvGstMeYaebv+NvlM2LikDoqA
+xpmsx6EBebageuDtvrIrrbvb5QTcSjoq057jdmiAMSPcIOscYJszngINv2xJV3X
ATFyGHcq5Oe5C5kN+egmNPBVE934jE88cDoRlfcWJiumdBIa1v1TKXk1qdyp6zeE
OH7brEeOQUDVjUv4ZF/2UwHAPd6V3YAajjiYx3KRy7BZE0M9P6bcimAWOnHzMa5A
LqY+mOhdz5TUvDvCamyLN5EUG7yUGVTduN4RDBrQZ0PRWYFhY0UqhI3LPniKzkqe
RzR91dmePwI9q285nOS4XlTmx9XK7vqwS4zuNsxZgDixf0ryEizi0GfKuN3t0gQA
yNn6RFkUKksJYjCnKuVDcIpQoG3g9mjz5g7iO9GO7fEyrN8RP0Us/XvolillYY5Z
xdWxUHcRXbmqYqQYvV4ob3Cr5XhBRCNLbnQgt5UYbuDXVV8Hf5K8s/Qm4jGlNZnX
giHz7BRa4YrZ7QAQwIo9FpmYo3YHV9uEY8HKwHCFtQQHTh/L6gtDDkbU7qgFQqru
xwwZZrxrpUjKsFc25K6y0Af6eaqkencx5fBo4gLyuO6kJwOdZMh3M1sbOljtm4xH
CXtOezC+sRLUEVkFMO0NTrxyHhtHp+lOos3DUpKljhic4I57s7bsQd8l6nUSVwQb
RKikrGttOQK1H9LINyyAbY8oIVBjKXIdUTGorHd35Ux9Un9AlCn710mKTe3ceki1
zF/7joZi9HDDEG54qgn9tO1AynQA0jr0Z2tbikwm6pxZi3JfKG4D+1DenWRxwWYE
ZelUK8CmHhGjAJqL+4cT/BfbNQpjA/Lp6ffqPf3lCHv6tTj540Hv6vSVNgWYZ0ir
zBbfNv13RONBOXk+lbVsXRoeItthj7K6n6P4HdP18ttom9qM7HFoGqKceWn4Okbr
uXZ9RhLGDIFiQViHzHL6UzN7OV+1D/s2vyfOKxHh8SVXm/Wr09pshH10UAZWGSu/
TYrw4/cxP1yy4NSD1Ikg09iFopqbzpUR1R4PK9jQ9ZDZ3Yk54J1Fbv4pDCm/QSBO
CjX1Ni7Bl5CVscCGkdHXftfKXVQlWLcpwEuP92Ts8iLsjYCTT1t53M6ZeMUuZUCr
QlM9v2+jNHrpfPCcaw5lTZzn4JWJKEztNm6X5EheJJCJj4BrC6u5qmUHaaRjEJec
QZRNCKvR/LgVSQZQ6vmw1g6JmohQ8PIz2xOMX6RuoayCrkOYvJ2m+6zz/LET7pCs
CLunGGisSTvX4xboKECKEs9cdyyEvSaF1oF6d0C2MYgfw69nunpHlkJ8OUY0DiQi
ljORL71J4bVflZkPLOX4lsC3jj5UXML146DBsTPDgvitgyFsMAZHkIkedS30fvYz
vGcYkf+CrFQt8MjM2esbq8q/zRxjo4p37g7Git0nQ9D3hxLI4gU1cjzbCVpcDmnD
SwPAu6S2jUZdKdbHDtM9ExIiqwFh7i6+yf/oLHViFwOnKT+tdK2V4qjS/C5Zf3Zo
zhnaQbSRT5sIhgXejIVX++PmVOs2H6KQaUCyDmK/eJ2nvcg/S5X39a0wQezscXD7
RsN+XwrO1Jwf2QzvZhXiXr8m8c019VSPEOCsqbT54JttXoUTRshnn9NnYUG1bTyM
D7xyERYsYg6HwYq7yMkYbRK+cfPZY7jQq1usLOtsgEOKLM+24X8/bb/lKCvcNRdA
wTkX5Ipb0Qdg5Z2V/DcuTP9bQjLOKWHRsQm88uUxXl9bTGlQ0gKrP6KJc2impt+4
YkMT4sOiETOcyeuzTxuHiKglibEqq+ESWQZ+68Z18/W4HpNo72Zpz1i96jgqd0cl
Cc4k5h2Hxrn7aeG6gYaWWRixi6/ogX1uPUo2pEOseQFLHvPLDVtVYmwZ6/2a01Mk
ZvR8rqLzWx5bJRJOQzK27IsdmTlFBJMAX7i6wEsXM/5vJ+XirxBIX27is0LZ4bIo
nXeFvKBMOppdk7VqLofJrx/h7XlVsBxYIVKc1BoRiMpb8b7SHn3I472DrKVVT8Lx
P/NggP9v8MiwWJbmPkURuRr8h2eWsfwR7eg0RFTAnFan12oHkyQ59xe2tmovrcbz
Lo730V2uxVp7gfQuXIB4uWL6ZjF1lqNuHypne/dSe9gflx3vLfN9dxgHHQVf+LNE
dwrjfYxlzX/7/9b2DMw7W4A6XEqmnfkVHUcjVWt3yzhemYT7Smyovd+CLudSNYcF
gVjlzUALqS9cCzUE1Tt8Ku3mSMOZnZXdtpzljwIrKNSBNwLBEzTBsdkF3zhkerXy
9t9Pc+iRiqk+EvpIwarSpKATrFgXl2Jva35/fxotarUr8IjFgo9eXX39rs+fDri5
M8iTgeluhd6Fo8SofCwaw/1OdC9G1xcBEdE/LKCrqQWoJB6F8AwsLorTi8dNUU9q
cwGtvNvyDaMCGSzL3AtpFA/LqVddF348scM6oqr0a19lDPQ1861lZw1HMfynmpjE
Q73ShQ6vPVs6kvHnyzl8oIsG0a/jKmPsVRapLD/73nCz6/9gWYXhwP3nMJeHAC7i
tm4v1G1nr7avZi4NRjuoSJ9Rnuq5d81Zu8JoTGj5NaCQiKzlM1D/Yi8jIjpIlRwJ
0HWm5hoSxBWSMcNNZF+H9GzN3XyT5h9zCU+5MDlnRZdbIMRJJOlqayx7zudhmpQP
lxlQaIFmR5lrlfnIxs6fAeLG/NSXDmDe1vjJdIBPzaihI/JJm/uR5ifvo5XeFHi/
adjwGGDGF1yfkq6O97ytZ+LsOnQn3kc9SzbydOMbH6amp0GXOFfetuh2/BsK5oRQ
MA0uH2SwpiMrBJOfvBcPTrSPp9PRER/q81CRmGL9EN1jHmJa26IxuYXBwtL0BTQV
3FRvH7vezOQdT6C+zEssyDQzTwiL5YoBUzFJZ0QSblwOya4teQHuhZEUb8LZiwfk
FsG/YYrFDmzsBJT17kgGVgvhtD9ZKWybGAzPE3fDLDp7uN0mFiN6R436tMGUu1hd
2ruyw4TCkd9TYhAbsgGFZp/nP5eLjc50OdHpfOfIVlKx9IDN3WZxY6offPUwkRPX
e+YYvtYVDjALmnvGAOByDkYZxlaUOqshLDLKwtFX+YIejNf4VQQb7GIvhFTRc3Kv
4xPmjJ+F5ytycueS2sNqzYmmhJ+RNc/XENRq6onNoC1s6AWR6o58wobHytpHMjh+
JGMOuydGDpFYodlw7Ygx5ThL1BLCyKz7W/XZBrlBBf0Yj9EJ0n/xNvIo3RZOXDX5
pH6Fgqze0iZ5tCD/Z8Os7BRu2yUnKI+0qfDOYxhbBOXRBgvljnYl+HZj6aLQHZBy
cltZk9jnyPCOKYW+0CFe0xHvG+TRZN7Rzqdd0/QpG5Gfdma66v4JgdtvEHned9aS
xrZl3tXz4uSx6MDD9q+4Nz/KhJLSl7n949qHDTQfO2MCSKTyK2/VxNOcKJRl158L
dI2zox+svLuCS3p0CsK6SxAf2XKMJDZYc2/dedn/c2B5jdpc3dSn1FmEkzpdVX8f
HYA5pJsmOcbWqtbK50yqgHsF7bPBrRLfRWp0yN7Qj6ok6rbEzcdHHvB8augOaFPE
JTH3AFC7SjV3Sa2EdTjS1z6DhPlYFQ61u8h1kZvj2qlRfkGLmYUWP78Wxg+2iD6e
YGRC8EYQQmkFE3rIeah6etv7/XTHVYlA/NCXQAipc5/TTDdzWmzgcrUFwpeA6AiJ
cjrM2dG9GfG8lKKqs/+Pyl+cvgSvrH/SpqhNw1CHUJv4f6R4RlGGi9Mj/J4qxSJB
YLfpvRW/Stg4VMwM1sMGzNZIuc1cthSUKLRJjW87ypoAk3zJ5BpMF+/PUTdULpNz
phyF3FtrXhYclq5M9mexmqUJ/kySG/waX1edVF9JR92dFLeDtWJPTTesTKzWIB1X
6vxWqfvDLcRKY9A3yRf2X3vrooSUfmk+8EBwMbVEK4osOb5gj0l3uWWcxbSu9myj
npAhsmPXB6eBgJYY+UP7CPeWvhAD0q3osTTfTun9cbSvZzwm+LDaMFwVdpcDAXQq
KfXZDu5xwdYEYCzGVO5VtDi9aswOMX/lE1OaLd9/iOUflS1z0kbf/K+BlD+ypo1+
MwStHp96b6CNq1Q+AK7t404x/lG7vpTKJxyrBv3rc+HdYzLVurE46ehFqwnom9TV
j9l5luUrLxsrzium0NDNHuw4DD3uDRRxM96mm2aGsl2aW+kma/aBK0yLBLSUXm5N
YtPH5WJpoXgn1G5zSV1Eb5h+gDDAKpxZcAy1sA3JMVKQTuBGRI/QQh2l6BXNFtWs
5gdewLpUOb24JRdPmbK0T4+gYufPO0kALunZpYFJ8M2jnJYWdkH6vju9q2KDbT9N
EAHAjfgwoIJw0BvvY4LyaEDePWaq6k4J4iUJOA7D4GRDD4BlqYGOQRXhH3D22e/y
7LcppGxiCDkmVCguzaMmHDzlytNKIp6kNiXJCedfZoXZM1/3boJRgLXx5a6FHh23
YKiuWAoP/LvYMFF9CE/AJNV/N5whjVHeNzmU2aEaW26tXuBnccT9XxVTwlkLpGn9
ZQBNCryhI45iyRrYlJ6xyGiExM+lKKOx2Xu0+NmqlGrkVP2BZ9V93CoIilBG6TT4
SOrrfoF7VZmhLUaiQsCWRK138sIZwtq5U/kyPgfvOAbLGLPTxno6HAnbwIUIf3hT
wHc54GIkAHFFZ7Xm8S2xPEzrzs5NPqwJT/cW1CxCyi007asoOAYnonfKZx8Bjhcv
yYKmx68eCR34QuaA3tTy42/VE5QZJfWls3B0bmOeDUsCIcQgV4ccecH2Wf35/gA0
SYPFqNy4ecE+AnPQWa3Uigx9DyJ2LBtq8tk+lyxfZcoCqY/Yky0r9PSAoajwcXRz
ESeZEz3viX1nxSrrjf3BoVQmZxr142+b9mkB1UBfVKgJAkOVebLva4MF4lcXe2uU
Xq/KTY+OlO/J4cbYk37Dkhh6tItUzKUc7dA153Hf7xS12NgL8PNHOJeBleGWCBZy
7PYHUz8kQRIEfq5XCDpckulebXqCjaM6Ms0OqbK6VU5VSPy1J2reBECzwlFinb5Y
wJYq8uqluxo+yapvoxyI2Zg1QQ/OqFmf48FzionZfeGCHIodYIv/xV9xjxQCIZS4
sfHZ0m28VNk/pFs8d1GQPAZdGQYGxW8QTYkiUyZR43npbtZJ7xwMoCpK4GztrMPV
3vwwTRvpi8VLNOK8OqZM7V3Shp7K46YNG7nqaFUXWlCU2NdxAloEu5r23itrsQ5p
SPU8YagER8RD54QHq8XDeziEdRLz8TmuiFPF/HOYqE3hQuK0sbvOZ9IVu1QxYoE+
vz5JHKb3GdR6Iw7f4QO1Vxjwlg8KWTvyr4qXorMoDNCb7qntDr3eBsz8MH/kiQGv
9cL98q2WabHunP3zR7n7djyX8ycFy4AD8KP9GQLVx3tgjSQg+lU1RTjStXOZ2up4
cEpzJMXySz9kL17kE0uJD1I1PUFDBxCAfptWB6lmC9WXyu+kpy7Xz41gbiUTt5Gf
UeQOZmsORtUIAIdJ86RO6HwHGWHwAGM8r/Hv+167KNt7wsxSidaKrDU3FviTmwYC
pkHlrjKxVnSC9z20A0bJWhhkaJE0fxEkAz9SAOEsDna0edc8VwyyH+qoZXNf6ndn
XnZwz39iUWDECTsm9txaTWIyOamXxndL7lFHFh0pZJ+KSA6XJcP0GF3rbAScPSf/
nQxT2uk1D1SBLGSvKGCfgRCrVPEuk0Y7PuLnsTrhF+jKpZtq75QN0Ur6gHUKa+aM
8wzjeXlyAZ5mnrQFDkh8+IIOJyXoIgnpxppQqXHvq7Z1ChXTUqRnmOF9el+bSoKA
QNK+JxObki92QZ7DU7FD3HjfwE4v2DsrpKzHPkWEYgIaTQLa4+iHSZLFrlgSFfNA
Tb2eXppMh0LTwmYlTRs9BJTpTeOMv9z/Cx9IiBxxYC5KBDXYQGsNtbplc8xY+tJs
wc9ZLags8jhCumrNb8YMZP1648e6No3Yev9WjAA08HXge1HPenLry8l3f7X3Fb/8
INH+hMRrczlooYSnpTSwLWc2ZmHNf2QJD3az6NXdbafG4u2NmXb6MLc9r1CYa8Jo
Rq+6FXHurhDuc6yJWsXXEv1g4JhTAMLNFC3pMM03vaqI7p539SPn6xjyhsC85HXc
La4EFUhemnQTSydfzgbmXz1HonzxU4QivunTS4+A9jVyli1CzMMuuzVWgo5DP/I2
oE2xmWLkY9N1PoDtmozFAWnXt+qUOQLEkHnv87hPmUOrG5eenz/Or00fkZEWhQSJ
Df/zi+9bAeciQhYMrULwrrC0WY6phg4Ai0pQJZnomhcdfVxRlT+j1sgIXDdPblL7
P8zZzxVwl/kj8Y1hAbb+yvktOM211FM1jm2ogFxP6nw16burAwQgcVyBOBJhrHaA
dRdMV18Qs2ZALLyxiMz+/s7SWgK/vxGvplayW4AgUppVOUhzXCpPjAVan6e0QBfR
bvKCYSJQTLJcLyNSCSvcdJwnGcCdU458fY+412xAgZMll28zl2rLzbXNOJXe09J6
4b90CeCEypcH6CsjfxCSRxfif/aB5UKcaer0l0BFxz392S3MXloUCNk6IGCGwKiw
2EbbdbUX28bIsK2GrPZVVyTrgwgpgwE1I40jhUccIJpF07SxZ+8DDvwYMT+THLJ2
vWZ8B17bURumLL4te088q/KPgARWk2MkkNX8Evhiw58tc6uloNTmk76s9ude6otq
ifrP6ydxR7ntIcb6pdDaeSa98WrX/a1Dzmlco0dm3i0gniTpn9JxfWko9z+/LWJl
6cA4HtLxW27V4pIjKJXHS65hjvT/TPHaKqNenyNuBlD3xBW2bvnOIlh/pa2MQ3a/
Jg/MMBuE/FGihrW5oUTVflxXjh/Pir7czm7bvgeBAn2TTxfZjBoWnj2nFKE8fzYt
6oUyzuOLWjbOSGBZUK9Bl2h7nwp5ffFFp6x1JjxpVXlSU7EK3ZaOxv9M/LMPZ7oK
6vwjGJuVMGGqMhJtIKcmO03/yYZD72oldSPvhXHYc1CL1GiJU8daMxrszOv/F/+B
sCjYMS57u2D7y7/B6cXZ4NeFhyEu38+s+rJtvotM+Z7dy3SVw1pc6/uwc4a/Sx8R
xVx/q0epCDfJSTXZyY685bDuZEfB1IsK78RXHypWw2bql2zbVLCSStywkoF4mx54
dSuAHa2SsJpeUF9Zuu707ZpE+wsX+2dNzN9V+4SWFqz5XVwIQo2y4KdC2p63MUsy
qYVnjWwNU1kcVeI5C4EpienG0B6xfLMw/SMm2DyQ2CMJ+dfipkMwuBpb78o9IBAp
LaMTpyPWe7hekBsSwcD6DzFlcGLzpiqvYl6b1X23sQX/wMYeMpFad+G3zHl9VXR+
D4+j7ZrKWv0W4fEsPim8cJflHVyZxSuJA0fyV4ap0ZlxrZQb3wqvJj8CWmIIRObl
P17EhsSEZw48pBOIFogSA8fO5jwXeH2nr8tg3U1aLolqq51kEraCRgw11LEQtYnz
Op/NdTCah6yeo1N6MSWit4eJ4bpOYQFn9maikR6jVapan4v7o2rcbZeOs+miM8aX
B1CD3VfgBEOv1vSYnUDVKVg7oE9fkjuMQJK4ENb+gJ4LE9PqBpCtzhiaXV/LvG0q
kFNlGxicT1hcdr9xsjIZyveGqNXC2RXkqPp2Ydv5vL3pr71pwCaP2aRikdK6f6Og
5ZGJYCAqGJeY1m6ffLpm9R5vGq82NDJ2jLBE4qbz6k4428ggAmf0D2E9VNhQmXE6
hKaRVz9PpH5LljDrPRr5r0OHx+HSPVPBF226WBGU119DrtCqQjz115LJbTJWkFM4
LzHMJHVTF8HIyIu33fITtD+NjucFB+Cwm9D9TwpU3VVD3oKBkzu3oJjNG74IdhCM
mrowRbu6+DAryZIGmDv4Ps3m1EqACZhpjrgg0BmqLbeImKgCuP7MdDHHh0XUSeMh
o8m57eQUs588kdUQdEWjh3p3nnlH+ryqFq/6GkGV5HpUfieWbFVdO8kqA4B2NES/
2i24ya2xz6uAjAVGaDoYdk06LJjPn7vVCKxxnoPVlaJTFXepDdTFYpR7nYpwiTBy
jcYedMhR55jzZVzilC3s2+9uS1WCbl+4wDZaCFYsZQxW87oOmsydYUR9VrLK+xc3
rVRRE9fP/es2cuom1GOmylf611Kxwss26h31Hu2ELn0QIKcg32TU0msz+L9nfAMO
GD8AAVEqwetOzKg8d0khZtSDRuA7fPS4mFB37PXtydsnB0yOl+kJSr74HhjjcTll
+P8hDqEtPXgI5hdMUtYcN9zfkTK48+6bw8De+Jlrnx0/hdLP6l5c9xDLvHbTvkv2
gyL10SJdvcu47pZPxYibrMb0XiCaTuAchmKSGjkkUT0dJBErjYX/ZIZu1a5v3MF4
9/5Vn+Zx4qGuRirdBYMaDrPX654U3ZI41sk3NRJn9V7/d8AufIs3xgC+cdnEsy6j
ObhCTp7AV+TFPlRQDsT2XJkxjqQX0sHx9Y+A8IGxMbuyBSVYuowC4wPhK9H8HkLE
Zvn6qcFMMQcPW67fvVGGYjzeq0IBtKi1jCML+iOyF/YkkIUqJUbYOgc2wvgT3PtT
odvUiOfvQqztMjJX/HHi6BSzG5WBzUaqkCH4CaBH9Tq3r+L/BOgmzz6zTqLURsDE
zPXC6n/tPPwFptx1JUWMv4ncJsVCkwRMiFI6eziGXL1IeYjUO5On9hr4a3opsSpq
i4IagJNdyil3GH7+7/rQ5IDIZkyJRgMDMkfaaohBCgeq5KwmqmsAmJn07wsFeXaC
q4y9JHt18TLywgi+/jSifLCbpwRADdqlN/I1WJRTN6Tkjr1FznKfBovvE3EOofFU
EbUZPIt1LT50+AZyUDR7lr5FdRgZ8KsWae6eve56Bb0sXdUVGriQ3NQ71tjqYqbV
nmO4HvkXBrXl0c/C4A2FCSj3mmYSS7+vGzYWRwsdG4NyVupYBiidtTBovvmHP0dK
ywuq51FPCsRjam5PFzHqAIcmQisW0t7FwZ7By8qmwCXGOl8yJ+0ArnO5NmL6HpaP
sK53I+4njPJkiqbfR6LxTBTJCBx9X75chea7ep6wu7mKY8hXb5SCuF2mdzrt649N
ADzCw2atcFQfBvvk2GUjHyy7CZ0m8um8tlBwcaBA/8Imrf4FQw8r07Zy7k8UfESF
/7gYZl5qDAFQ35mJPleeL5UiErzzM3sGDNRRDBjeHy8ljRxi3fZTFUrdeyWOjFFJ
CfwYzq40ZGHmrmoNoVDQDVvxrg41TM1yWZ90ahvigWS7ebfqewlniqoKqD+G3L7P
i1pu87gS/z03hYispKDMdb7cF2fC/HGeok9SBsY1ah3ybu1sPYmKsI9nkvm7ugFl
wX59xD4wxTShQS4RPurBHqOg1oWomtJfGv3TzbdPawoWE24hyjR95aKx23J9nwqd
Lf6TMDaXk5vt8F1Fx9jWtE9OG7Q0CCJPUn6T/63+FbIBySdgk9vVYXJoi+WrmmZf
U3MAdIw6h/y+ZHfV+4mJHiewSBUMiW0qZlU3krM/ArQ34IyNw2ruGzG5Y+LFVkIv
A3s+PlSbKao2lsC/349ToA9ZcgVowI4f0PnhplJOsih2gfaCIsRzb0O+f/T9taDx
PjLOOtdQem2AS+0xHGSuPcjg/TTzeNOGln2Ey0Z3R2tun3HvncEET6GLBTJaukvu
q2u/+RerqVAPw0tAdrwGKLJC0pLK5AmDUwI/CrAQdao3ANfYcI5pIjU9KvlwttND
zZ5Xvaav9sqzw4khXrhR42gk0NI/oA2LlJHDWqHonhKTzmFRVJY1hnDDPH7x9XwG
n3pkU+i1rpXb95V7dv2uEVsnroERdrjsA/tbb+ZpD0n8OWPsxtdpeSvd4N1JfUPN
bFhKtYNkd7xZ+nfA2l/MsDZnfJuc1td4todzXUcdrh/IqDKXbei2s8/5yzkp5dQI
g+Vn7lu1zp/SESCWk4Qr63DaFrBmQ8XROq5XEJBHA5EA/c2BJAYrgQ93GfBoyXDn
YJuFZS0dg3xp34j3QAKEkjJKlS3xYrP1t0pYlltOSez/5W2w8sNBVXLL++taS0yi
cfPQybOypYNVAzmWUDQ+2zECIDzCWw2Od9GhCEu8tkKnEyY22hbL2wRO4KIq7XVC
Ft/MgGXKqJykCpq1FzcD6Kyzh8Vkg/8COYKySmvKGitrvRsGwVSIEozxap/xvAdQ
RqlxRpd4/NYplY/VeVDCk02+G5bRLgLMDEXSzZ4jEDOpT/oLwwkJZNNaJsRMlJmr
9ehcH7hovbHSIWq/MB9q5bAhNAQgDDKYqbho5dLchMRwECIQyKEbQBAvoxK1wJo9
Kr6X2HUEzJuIT7OzK0Dt7LKmjhfmtij8ELCzKCkRQIxHq7f69txo9Nws94KpVruO
fAhCUHqet2JayDlYqSyxwlr8BL0ILiwjRMig681kjT6Wmo5T0G7KrBbwa9ng+SVo
yg5BXmgE2D9nkAJ/ji/2BIL/jiMjtfLbNBmGx5vUHTB2ohiqhXTXMnyEjvCZQmA4
wbRjF2aJh0hiDc3T1F7QZMnnFUuo6Rr7NMB2X12h9jYT54ca4e6Q73ByOELD1u9a
4ylJHp/RBVIeh+cMQBbKTCMCMm1t7bG+WkzSuv4CjvwjZQJKnUq70ObrFo0VqiXB
KA9mQIrZvWIqX56SAbX/XwA1xmqIYB+7KmuHZrrdt3OzMnIZkqkmyGdSHTyGIo61
kBWL3Ko43erTMuanU+AT9MLWi9fiNDexqv2/gOFXH39lxZpiuq4pSLEu6ZJYwq89
OSIHw844whA+WKpn0kVUUbXw6LewfmHBE3Ysor132emwxhNZNdi5lw/9rUOcTwCs
enjBQhtJwLECLE9qf/lVQPa2PWrB1Fzaq65okbYjHYsG3lyuof+cqMpBz2I7kzOz
YYTypwZcKkrgyFsz308cu00+kUCTmUaQiYwyrDjtUeqyzgxy3qHR1SuwgAUWcscW
RUjy4iN4THrYTe8McBPetDYiFzmWMuSyGE//sGawJqoPOas4SINKvw2d8wpvF4VJ
XwGzfsiGC1mC2v7n8LWBB2HRKieO/qCQXuGDviix2yXetiF+m0+3tWZfrLssvjHx
A6+j88X6wWlTb+841tP5XkVUbA/kfaa/+om95k5nv/DwnPu227nsg1oK4KHgRCg0
BvX2uAo4eHPAvUew0KDhoaUQ8OMgu81I4m/LR6VY1Y9OS6OPmmrKo6ydHGKxng4r
jX34fZpf1Rj/YYeow+Rf2Crh/hSFidURi5pemFut6jGJ3Nf9oo+/69rr/ghCMrUH
eFn4l9mPUdCbYHLd8+c2He1gmm3OjUtVR6dvNAbGenFPsh7jIW651L0YYuLOHDTq
eKsUTjVRURRZkJsaFWYwZ95j3RQRWE/pX2DNRBYalCaKX3FssjpHQFNjss7gOaYa
MsgfSHf+78aWBY7GC4foZjkJlnbsUH0jaKd8H/0I1Giu3dHSSVq9U/E+Ct6nbBMY
AZz8ii6Z4BXEULGEpajJe2m0bpB3kYTW5JiV934Bvpypjw72J9WsVNm3R9dv/4aM
T9EjcAnxs52KkEwLEJ8Zos5uVR2gusex4cK9pi+Y6ekBcfISo/0YtcTUsLjqd8Vh
dAGSOG3FaaJUKHVf1dtM5aXnCvesPYDgleXGp1G5zuN9OTcYPn4gD5HivNcNRuVg
hgb3PEl2GhHW/JCJsKKhS8VIDGIIdJPXwBxPYvxvCAuQLglKEIG1cNuXB0SOanwm
e5Alf778LLIky/79N0lAGWP1L3K7QtD5dSSY4s9ivGmAAUO9QkaiLC1OEJ5EusjO
Vpvk+cErbpj3tESe+ocZuDx6dUs/GmQzm088wM0qs6/k8RMIvrQRUUVXobj/CW7v
Kixt59Ox/2zEZ0BELWFSRGTB4BWBxCljNskGNE4gczEjEDK8z/UEkcIHbEEKjEQB
Gz4/iHDDjkj2RSQt5CycXlhaNjkny+2Gn456nERhq+zAyuBAt489In3T3ifx0qYO
KGdrPl3lJ0FhEjpx5q57Dop/GxjXF1SlbXEQE2vvpfqdLGGcN9Cr1Zm1VutQYRc7
COCvmpcwKpM1psvtLJtEe8wePTfWruIQh/tnM1RHq9Su30LSTo8MMkNS+EYb3iaQ
CY6+QofU00mMARdXDvmhXsn+qpBwZfK+k5QJab4VPJ2VuvRKz9a/Sn83oKc9NLSs
/SXSbsrooe4gv5KSckKF0bLfWIQNCOpk9LBGfdYATCzlSePzPeI+oHQ6VUfITml/
oICQWzp5ych9rDz7bTvnnkZhhEFdJY6WO2nqfZpCX8RKd12p8P2vwxV6TK6IvkeK
4BbFtzv0KUCpk4cf0D6SHZZP6b0kSfqp+JjSKGt/h+WmIQe1pL5Kxq82mhi5V0PL
HtFQ8LcaSS3Yj1u7nr0tt9roksAFifAHZ587p6IiRWsQSmre0Mhhurj0aD5A2XDr
2j4L/jWfGFwHqncvEHJt60c6LdFI6Mwxa8A5R2nDdGOOYp6+xWSO94WhjS9U2eZ5
18xrAkzHbDih3mggnQwdW6VEFt1hhYMHVAOhWFVkvTpafMnRAlRDGgqQQly6gXbc
6O3RkUCJSX9HV/xkdSWTkZia3WgXY0BkGFT52P7ilfB15W7cfQV6On4baG6Gquuv
itdRmaaT5mHFYzwIthhsvvpc5I0UXgoa9xmp81KHI+5pKG7ZsjDA+wQg1jgQjR85
erjf0gvfw1nPxTn3NN8/+lvedaJCrQ9970bki4wx6lVfQ8QhBRgMOxN1HSZVhDbz
nEwMxI1gjXkQyEleQfgMtSrkfh3hhN8oj0H2KRhOZRW+70PFUTUUIxpEVYc46eTm
GWZTk9fBpQ+4vho4pE8azzs852BTczujNcqFkw8XscjoO7DA3w5vX0e1M1Ef9nY6
ydYOD0OHumWMomjrmYEc/Lz88qqFfuIKfd8VoPSQomAyFk8HOmxWIqN7RQFk5n9f
IZ45cFN8gZiEn6y0JGefn7IgHExqZTn/5WylVHLv05kHqKvHJUjWpjRvSoB8dJv5
c1e5Y6W+VxLCrn8uL4wtK0n9FpO+rI7ySnZwpydOu1RTC3m5C/0bN66C0wDgjiFk
bWc61nGmUfg8wrS5/F6e0fGGCG0d1fMg0FJwdVWyiD4Zv7b8uiWiM0QbjpyE6PTY
xWF5S+UKg5Fg8I7P9RDchpIZrkA9kI6A9MPITy6tUvRnjV+UNR+2EEa5+flCdpbP
BKjdel5Dg44onyYvFpTteCVbRxW0Daxzb+L4iXqlx8c1S3fSU1U2AI5DPnxfRiNY
VrZhRPKGzeQ7X1FWXFVGtmw0t68S+QEBf0RT0gZJaOgfrOMH+byShzgRImvfBwK7
CZswfYGgyqsUyxd2L3uUSs282KMb9HVmBA31o3Oz0omG9sVNgpzxwRiS9Wr5kC63
QdN4fbyXSm5aM68IKi34MdeSKj8w3klX6ES6KMiQo4/XoXTbnPahHxHBmlOrjfpC
n4kgExVw16GLG7spZwYAptGpv/cOkmdHIYcl/+MSDN6JQ1jdTwuyOBB967bN73aL
datgivpnHqUdDBiJWAw88vGJUIf12p+eCp1z5es17qdCVGfVGBOojl0iIJCE0LA1
YAjZXWv3rF70GpOxk6QRHbw/Ybi1/NyCo0zs49CZCS3RLEHujzZ2+NBNOLIBHP2D
Z3vwp4o8Om0fg2/FVzOF8f7zQqTx6EbK+QDVZ/H+Q+sqxeUt3GoyQu7XA/xwP711
8yfVdRsonF7xZjPZ+9BBeYr+jJTdL8KX5Y2am1ZEfCg0jLCEwZhBq5HtQf3K5L+t
aMdzjxctHNqYPIjEW+ekYqlGqPflcZpazw215JmN8N8r1vxcDu5JwPLX7pIaP82o
SbPxNyCsbeua9qxAyyk2lZQ73srySOxV+dfC7O0VxGIK+06afAb7FtmAa+iGP3vG
qYd5UUsw5MApdp4HW35VJzX/fM6X1nBXhb5M7V1cqVvOjnoM8bl8lyDwaFBEU4Qq
WzB59UZH++Z2H72/7kASgZcAzj3UbREx7P203b5PYvMGuaMi+9ZPCDjKkZ58OkNu
wfmjj/mSMYGMsS9xWGhfDIVuHMCA9z0r1ORsbcSGljmVHcFr1k+bR5s32V6FqfDr
UZGId9ssM9GDv60FXLLkuppW15BBN9rz4ttCnnk7nP0gvvMD2mQ2+cUT70yPzH0T
kn19siXP0vzWAGwzNlrSuKSOkyANLkAwdrt2PUvyR5KE8kJJs8cU5LBcFteFjNxa
+/biuQsXBqaGom7JWfoVeW7R5eqK7U/w1U8IzZuTP03irgzDTE7fSYLC7EnuWinw
P8noKxj79RSMCeVPJoLkRfR0T0TdmVwXDCdiMsHUC8nQuAp27km8baA+BV3cinXW
98c/3fzN8HAmENJoi7Els+/Lav9qV0CCtl+HGqm06mTaB0SvdaUOnJco2ow9KXae
s9BKk52om6enBkkE47GUeebEJfCredtGVDuRColWGKSp9mrfX6RksvahLRdzsP+/
y5LHDpvt6kdI6+SdyMf98iiLR9ya7YL5bZ7e+Dx3Rmj5N3AGuWrPEwRFpSg0dNPw
OLPQFiAV18ieofs8eWWW0q5OHwkPCAIFJW6U/CwRoJFcU+pafyTQobk8hz+VQp5o
mmXzNaoLROdg9vu5pMo3H8bY3RgaoYtLFcet3NGQ/IK8dyC1LEPT2LwG9CBIQcLA
BFy8iTcbRCl4nHFd1e27gZfVd1FKmn9GZfNTDGJl2RtpyiCi5ZsdIwMZggazYjjj
vMmXQ5LZAFauj928V4peJ1GW9ZV5qF+1DVHASGqKrKU1MkjvC84uVAoDz8pVstnJ
Ln3cex/gSmS/0Zw/HNdfFH0lwTAQH+G/hGCFpVQ6TuBM5E+j5OielR0SPzHjAi9p
gmo/RNHACpMSghEkNamE/+R2qziY+DYRxMj61j6E/W8QMZSQ8WEXNuqJ8f/8UJZ1
iFvibcZmbbh79/91Y0K32TqShVOkj+NVTKIGFJ8xjnUVQfY8UJKOlXs+toLvBWxh
CXcy6eOVrtxr5GWjvL1ZkQLQDJEbCtiJ9MMaq9/L1InJZrMd4ekmFJiVRTGsMhMm
oQydUqiA2YKRoBc5LZxpevhxrabgYS8xboENSegiqktJcqziIMlcaqyOme5BY0EI
SN94M+D9ip8vRzfs9D1ANl7A/O8iuj8PT1l7badxNVOcU3esCftlcZFnqNDCWK1N
jbtR91xy17LR5TJd4qDCP+xsBd+QG8Md6PmDbjDURkCsIWBR7q8CJq9hV6bie76s
QRRgRnD+VN91yfW7ODUV/C/eOyoAQo8PbUGnj2vEeFIwgo4GQUn8RrEHsadkdioA
03Kxaz8n7vt8E5wZ9Kjxnd6D+WmWay6+UthjsqjCacpnpd+lMmHDgUMWnnAZ/h8G
S2+KJ6KJLRc/0tmKQDCefXLkUK3/NoUnPDWUmCkWI4lv2lunElSwbx8r8NYdLDy5
9gBWAvPBKeriDTRHNTEHdvYiSJ5ZL0db2jlZ1+VUx4Hk4igcIqs7kUvoWz7hsnb1
aQTxngBDIVyQRdUOMg3bcoNEbEbXxuDX2zj40VUeNea5i3iBivT1AQGcfL2qHVO7
vVdslGPnpMyE94eyNvL3YJP3BDovSZRThmDDI0lJ67ILRx2IKAVL9YuhtSF7lFNo
6xhj0we+SCm/iGMWv/UR64v30ByuLn+jVQElalhDroTe2kcq7MufJ9drdF4+tfxl
DQJ/u5yGfJY+sDJ+YyI4apXPl+0Qz4jfDYXv/Wo2H1dCIPSvGdvpuEOOZykbqYi0
eY1kjlOUoIPPyxPhe+lNhc1oMURZNCoJBA+SGUlYiJcGUX4b00i5E81HIXx1DNGY
igXt0Zgarm2JBDXqOSUuXEkjZYpXKg24iSgb7FXkubee0bAR6Rdu6CdjX/9d+R8W
9JOfcLiNKhPPZnaOqNM31V9sbo7PERD2ZHCEtwYminBR+KkF3SMCot1GMVkB1BzM
+sV2kLxHk7ddr/4uz4NA8Jup0AAi1aP2z/luc4uuLQ+HKhLSxU6vBXbPYfUpGO+L
CIH+CGZxP6XOtgmPxZZoP8GLnOCQtHAgBd372zDm/Pdt8QLVDgEQbYqk+/1I/QJs
TOxdRNbl/DFaEnU0AL/nnAkMGEIwF5PM0h7MkLPZ4WLNUxNUapyc8drz80BVM9w5
SVu8+n7CwjkRSiesftAxg0DYJ7GpXERoqzOQ1SJUYiZ7ayemKD6ZTc5qEUydk3F7
WbgzES4CiBiAhi8L2N06Gs6wV2XQ+f8mufPf4isV+btjyPlIjGT0xUTZ0KbVTyWS
JmNpAgRPji2vn5iUqchVyCzgZr7sZ0LH3W4R/1ZQQh4F5tfVVy7OKL+qNlsgKTgR
7S+MuvFMYaGXIE/T0aSEQ0KWNcO4BCbkK5mmfd018+15H1zFnrvVI6550EgEkjlt
OmXDjhX9WXSsVa8+r8YMW8katxdp+ikfgVfxFo8id5yMyPOMUCDcmKmOabrOuD2G
rVSMGa0jHW5V101IRfrb/BeirkgT1n4Xn3ZmPJLps2sVEN1zYetMMCXisWbMMTgM
ZF/VYCAEnotDQ8dN+vwZwKXHXSRsg20A7PIBwQgASesrHud/97x94och4UuwEXEH
58yPcn/yc5XrDVmzAdC9rXdVk8h3L6NA7D6/cYTNJipDwvole4Bup7GBE7w6VGRj
HY1QM8pyF51DKA0pWXszley9KgF4NSRm6Kl4YrjaZbDggyy6UHAPNNNIt0zeoFGp
sX++DLq+P2T1L2MdRjEbTa3u1Bk+4REGR7G8EgwibnJ1z9yr2wb0asuG/qe0Ku2j
SGWkmFE80o9P0+lRlP2wSncW0WN4BaZB+EVafI5wb9uRfmElrc5q5TevLgmJU/Mj
Z9XmJWZy5nrkQgT8XJ329h/8lZXnHO7VxReNrswzZXXblJg65RqRzZUcAQFgVE3z
yb2arsFwpQGe+ycTYyTPe1igmLEFs8vCUM8vpjhQ1+yIZGEucuDk6oMzqr/1acpM
FdMfxvgbdkykxmNncE+TYXpa2fYwswCXgBVS5x++lScX9zpDxnwAvNtaxlieBxAr
HE6Wh/YUYS+NTulf9KnJQ5c8MW6BM74/GROLSNzQLrbI1h35PUlP9Ixv8mKuCyzh
iRneia3qxn0Vnf0QULzI5tHkQrpzwO0jsHIjombkUE8Sba0FqoRRfwKSm6z/eVXE
k7AnRyUAU0Ke/mHcX9dbzNsDUf8qEfs9TFgOsABO4zBD0DL63rX0aQptuBGuzP4R
dQbGhMxu3VZn+iOkI69mbDsSBwY55KGMcKw0C45GWXocO5MeRB+CDsKYWDhmCVTS
xyaVFA5EFa72Wb9vZ8a9gsYZGXEBRpTlYJQd1RAARl5tCoSSVDjQHXKdmczKFHtG
p/b58YLN3fXQWgZd21NfMAz9+bHPZNDIrKuleR2QONVQ1XrsnlYm6j7IHG+o9Dn6
e1AnTcO0DobZeIWr8XzZlGtFr4JA16GqgXimXairppgtOtkn6+UyPagpQwWwdoM7
Po/0gR99J+8CcTvFPUmQwBrwXDXe+oBA3fVyWY8O+Yd7WOloTJ0hnkhyLq11B7zx
bP/zvHblIT582HwLZgyT73awfT70XMeC29IJSkk+JECtV1IucA4MDxpQbq3sm/UM
UWm4QtgkkeKS6Yjg/JefWvZh8T3sIFCgaGP0zs65uRBwX+kW4/B3/hEDBWsDXsiR
0CpiWVtZiwFNSvk+DkkgOqoCeeKcSfGs1QXoy+64IAMp22SF6lAK9bsUflh7n0mX
dgqTkuTF8QbQDKQ2TQusywCd1AqWvVaEfKNZ2efP6GZZbvJFB3pleq/A1RoysZY6
4kY79ciKi5HodS4yrzrJf82Jky2uyc3Usl0TNoDZuIbutQt1RMNnm7v3Ns3jpR7R
94G85QKJQn3F8susEx7SN3EPRa6qSi+vqKAGQMipHNqMOpzjf789nRAs89fdwdeF
Oip4rnE5NDdS29xOf+51YUxJ8wqGcBHSHJEkd1NpNyru+AaP3Yao8ARTZi9sSmcE
C9N45zr9L4hRytKkhI3/WWAXekSxR3Wm5FC6nalFNCjoNE1QRPOIcy1RcCRz38qt
CidCloe2lwZeM1foiLswSWh8ZHStRxazSBcZIYxm89L0c7vOA8AMdni8asx6lgxs
h+CRcqhA0sSCL7LRC28u9c2ukthtGqVXh0opuDHA0HZxwp2MSJSytGELiUPTHiBh
oMtWXEdIZWNV6RZ4dN0itqPdifOdNKxck+OdEYIWVgh6RQHSeSkh3PrFemMp11vr
WivmE19CyRozHXj5EriDO3FF92BpbdMtcaNguoLK3PnJ4SqI1fQ5CpK1hS0OEXLi
dH+kHlCVw7vvARKjwIdkm91LiTrW5YfRF5x78nVY1a2nJSDKM5U+Fkw6eDvx8cwU
a9FBWFyKV4F/hEh9WwhnT75qglF6k8zJDRWTHzhaq+RkAit+6A6n7cYN85wMkXvM
96vTnNriyGQ/tv6MDO5Zd1UEt10z/o9UQyXB5GlDmnV0qiaD8rmX/yeF7qa2W1me
npMCR6MNr6b1tHGkZSJYr9vhmCF1D11y5+SJycexRvR1wCcslWd4d8WI5W6jDys0
XJJTp5SQHjsJ5e60CIm3ln/M8q6sYuBXpt4+kNH6hL4jHBIrfG0+8BenMkJb3mQT
dzPQP0Ucab6+aRP9443MtFkJ3UHb4YEjub8Iln4PvrVNpSNw9BqfAVH7eAgA6uZw
y5teLfW7ZYdu2Ro4TdlVdn/U+7Uibbt+3dw2P6CDCap79nNOOMm/Zw7TPeXaU+iA
OCkqEd4Bw5tFFuUEIH065vjlB1U0e0Mynsvv9qoP9PZ88bTz8Bvzn++/Q8AJwI2j
rmxjd15D2PLy9N4qmWQXhRX12Bq/9dxgqKSCWSdaRwuT35Qjpg7S6bxTfY8T16Un
pXAENxz1eqzCO6xOHFB10r3vLFAwkUYN4exR0fx65Tw9QDwgNrsw8b9RYF4ucnz7
NONybqqGDu+N31za1aPAoxsjvecF8BtYjfzNfX6RI494jfchgGDE35ae9mBtVw1t
Hb6YlpSmfauNSxFSjEptKPIHNBQyMwHo/zVy87sFtJQqOc6E7ovJ+5/URM6TENL0
lCKSHstLbLUbVyzPywcpy7oCehSVJxI+FUKSDmzEWeRHU3fHZxQ06dTVGOYaTzhT
aiplbpi/40ClyDzEceUktWMB79WNijyB435jKAb5FLK2rWHU77EJ/gTXTYHVSkqi
q+tywk/F6EWpFvIg0SXLwN5B5TQeKT8eeoZGlyL3/yHvnSvdl2CxGBzbHWvjjIGg
1kSl7wAMH9RePYuP+JmovsAa2ojnZFzKyCMJCD/GOLW4M+EnZeDuDPjbDndfjTO9
XAszx4a4qnJlMyXfgAhO0ukBq3z92IEhRqzIB7V9ImoKJtQFIMPzMsGIGOFYLo72
/xhB+GJK0rAcYLMPpfrgNvS4Lq9iIu3b2gB6otgGoOBqHcGQ/F2+oS/Zc+hHK65E
FgZQKVctXW5taB+Xbeezt7bicx0UAgrsCwJq0eFFmclkvZ9Sp91of3dcBXtXyKs2
KTeQ+ilxFadgq67TLu1ujCmEfRJ7MvAsdKbr0/tWccXe09XbuHMYw7o9eX7oKJXU
fk8OQX2msiDjFES4fQTd4pq19SZzxcrQ3LnY5IpOBzi4i6lduHYQWwSYD3A7S9Nh
Y7p9DOvMKoEjGyXV1d0hwgQfv+oO4Rgh+hBKoe/k0D8pQ4NL3ZU16ja/So+qw8eT
EugK6/c9H93I6mz/q/A86znHUiwW6/zdC07KzvNFRu66WOBed9KUNmqFtrnsj7IF
Y1jdVYdrmBPibAhY7DF+bUfm8ZzSIYzMUBrDzEeLGnOq6Cil7x7mhWz2Gj+Hx6+A
4+BFKGAmPfcvAar9UmdPBgSUAkubdWvN50VvOCLmSQm5ntKDXp9t3oLjnb8FjT0R
3wjcw4PQ1Qqj/Msb8McREAKW2vjo59ccEG/PQgVwvHuolrBGxA36PQVv71YZyfMl
5lgeFLtu3jdA5P70fh8ULMr6q8JQRoKLxi+s8v0Gs5Nq44NPeiyrnq2Nn2Z9beIt
Xejmafn3Zxmm6IA6jXWmxL57Mn312nqGzsgSy51lfYJuRAIeF2KJwZ+q8kynpNQe
EJqz99Wygfn11TMnzpPOHdzuk9/+KvAseKtjjzD3RKxPCAhJVjfQhzwbwgw2b7yM
R6r0s86pYMZPjqai4zQxITjRaw7ayPQzuhGsYGBUW/0tthN4MmuX//wNx5LS1Ca6
LMt5HhFIfF1wJicWh1pdGdkZ+fW9Rti8q7A22uMFW9brNx5OwKHBNyZNvMNvxmn/
VkbWhpSctBGcoNsSGP6BPqLqOIhSTmEF9JM+FhahlgJ8h5YqBTIjS4fwUx+trNjC
uTc+CgMuCVhkEc8ubFwuBMEE7LeBHXxJGaiAO7/X4KtdXGb8O3asWorPoxWHnrxt
lNc0XncYBPXUtDWdgINaL2tfOW/UgttKbKl5SFX+nDL7NmtSRx83jJ4WPSV/4Nk7
toR1nXZRVs4Ub7pZGepk8luhDiBkhTsa8LBliOrXOJ5BgdAwv0bi8r/9FMqhOvya
6P2xgoBTOjBIsTPlSI30Dzzwj2JtVWjugnigAI4pX6do4lKbEZN/JZgR1xX5/dQ2
fbKsYMiXUUJ0B+FDfMNrKrfzGOID/lL/yhzBs5eURXD7mhRWw5YZzSUUI0hp72ap
RlyDAHNzG7XU0+IE1bzgZoUvAVjmOqgLnzmzlT37HPtC7D5L1ndWbxzq9+y8SKdy
xz27lFFPRWYt0sfWhj4TgIHpHln5nRkyW/NW1YwIqnG/gC4iPVmoBckRm4jLOL9p
rnPtBIUZvp9/SmmcYyasDUQdmf2Rd6XPbjUnuP6MwseMoCpfAJ9ql2ZPSqyHZoRn
wm7UUxHuJXOpsT8GMt5aXPVh9TCF6tQLABH6IG9JhySWX+zSbG4LR/AZLxQCnrTL
LYuYiFTBayW/QM4Zzm2aVs1hxZ/WwTwnMysls0/lwilcQUaB6nvIsIOUKNBpFTGa
wj4YgBaa9B8lRwabeG62sCEpdGRG/dGm5H2KEqpY2Nsk2F56w6PufzV7ymXzpPap
PlJQcJ2w1oWoyAaNP24LqMYjqh5jqQpQHLXIW4J6Kao4W36ee08rUTLTpgrUMaXm
mkbi3UTG7tuze4G/Jp5OOcY7cpD6UyXe2IDqP881nRRiJ4jcSy5eT2K1bqS9OPrZ
ZF3mpSsGXXWeBbWg9HkiTgPMittskiahyRAfsw7AGCNSZ604FklQrq7dDjvpBber
WuIEVKGNAUdzrfgjkrRSqn0Y/jDOvW11xMidmcnerlru4UdvhvI+IeOrQibxCQkk
hPl336wUV/6F/aIsgkOzuJpvtBUl6CT0yDLwHY77crTPsYVMsKEBKCevgGhpMKL3
L2kaaybVw/6UbAh+pN9qb+IQizHRZYMlqLXJcgl2Evl+hv9tyx6ZqQ4WNfjkZ9Ya
OAVWrdccLGg20ul4nbgc6rCcrS2WEEDMCrZqe0wbju0vebs6Ni4i1UIgGnzNtG4g
wthSP79K08Q9Z5VxLuZsDroA2/ZWTcI9NQCHQYd3Cl49aPi+iZalbI5wFyfSxJOf
MnpIFWK6hM5mLTli2IVQeAwKp+hAXtfvkaZJaHnWhseEYC3VqKMRAs8doOC5Coox
JhfhgHByThcr07dWYExpq1DLGf+e/C1Vvez6TtZGKDNIk0tx7y72+3oGggamXg9N
zKCuOK3/iWgXZp6Vr7WxOYNwMOQi07IOWgo4bQaMpp+AgxHONa18oHTTTdNR8BFQ
GkjncLu3G1picAoYPlJeV2OVNI5yyWTjVCAGUZLB4vl2bxmwCyZndT0/fptylfGI
AkTGydgNL+gG8kw0tpVswjjQcIhtxIEnKAqZWdNSNcwfHXfTyGp5b2t7rQN0AGmb
liy997qx7Vd9LlJ5XxS8TXAFileZuYm+e4EEGkrqaWZpnvRFVajCkTCqS7iAO+qY
Fwc0lrfR9YqiZPfpte7l9daIEAKquglpjI0frC1Q9GsGq8E6T0l5exhxKXMN7rNP
FCrLPKxNLOoQLWTdNQqoczI1TgNXZPgTgNpFLNwaBTYvsriwXNp7kIqfR5l+7ZsU
Do+Kq7RG8Bv7WQFHlTGPyv02OTMhGl57B6HvGf8ZkaAKLTqeY2NdpVVs8XeM0+Iu
hkRLUJ8C/Nu3HKT1vU8Z7aRVPHAvm0JBci1Vacw9+v///M8NvIM9oc0Sm8CNi0od
2thiq8Yh9Bri3WPgfhr6gIoHXtGNmBaTX+thLG70jeZ0C2GDhcj/SL7koVf5YMtd
UWARSZGewswQK80Oi9MOBjqCKpids9az8f7QIUIh2Uu80KkMBTb5zQN6YFIYVjss
oLJMM5sZarNCsnM8MuTx7mhk1T6Ale4lO/2Gqd3PXY1TwmmZBSEZLMKXKExi6/JT
ZV68A+346HTwIlSDnlhASkszqbluijyvt9QO/tBplphIRehyugpr8OKutWpookeS
T6cq369ES0MmcrdS/KNNx7625USiAmeVzKSVsA9BCO6+euiOYYHqGdcazQJrfotS
T5DFtX3e+ds2nbfKGqXmrQ8RRGsvUADL+rtJuhrjxbwRkPDDwXM7w90CrUuXrqm9
Ai2HQVL84kdR4QwmYa0DXtn7nVVH2deKdHQ4v644oz2XqPmLZupcOi0Wt6ZdiGB0
GdCs+SO5L9sBCSoX98c52uPtG0cbqnPUwJLQMeG/QpCSdpsCKTdT9kXdiSSquEg8
sbdkhOpPTcKkHopU6dd9klE21b0qqlR8U8kEzt2odiKmzwo968OLu/2NJq6yZ7md
C7FaU8FZdnfLWB/9ibJR6wMk/MSG+cdSKm7WSk/MDHcz9AdB/EC7u2QDwzvrIfXi
XvytfeJdrGUChRyLouVicJvU2xTw+whMJ6UxYPoUy1dquZecbNgzjUnfB5KLpqtC
4hoeX5Pc53O1KhFequQu0lmVPxGGJdgzGyhpu3kyZV6/Jv+9zXlT116nbu72kwPb
LEpoKcm6J2I9rTk1QX7ICa4tm0ixfogsOPFuezfucvQZUZuIO8jZwJHYZrVtDfRF
uy7nqaFvNOWHQ9mgUo2nHrK61I360a+cxrggp9rQnCRKZ8zMDkOgxQ8FN3movPbb
sKCCWHjm229wXVr9FL5iBB2+GxC9Q01MpYVr7fnYlnLL4YAAcoYAyFVSZVwU8M8Q
KT2QThSL75wKywKhgXnIkDdp8vzGWkq/jDQKRc9Y+5S0VktK0dL+Nhi3reTdDfDA
qs5WGzVsZwDnz3ohsipIQ9mKATRKdQ3WhQEI2wUeLs7PqKKHnJ4LNpeSar0gSRgr
bH05GF2AKw8DgdSlKU/60W8qd7XaF8/Te/R0trpRdQxl2CpIua7NGz+RAX04huBc
MYB+CRiCpRoCisGNXqcRZFqpAzX93BQ4HRHtBqIsRLb1KZgHjqahgyv0xAg05ZNR
xzWdnvj9PFm8/TS0a9ndxhLCAuGCYmrjQBU/bg4A+PiH0ltH+SBFHbXMxWQNi4qP
bjOYCpawFAcOq6KhaeYgwG+5mcrvvA0zKSiAo0y564LcI/g9hyIpYY5NK1j7iL+b
0XFWTxhCXGasPW9iCq+c81eF2v0skVGyh/a4cJNsK/5+F7fgtu8pXAaCnzDb8v1x
7Bkff+O2ncMmMaAPiMPde+KD+G8Uu7Bw/ozkqmI8GHFhPWZD9TZDoKlwKJ8Z5gck
xVJPdo+z1qTouIawjdld4R0UgAiM4/9KwVHgljunPvV7mR/V0gRLpW/r0eUX9pb7
1ok6bqyFohpr2w/u0e0E8Rx+8NA/OdSc9PjSRKM0j/jp9b3ePn/sc5/Dy3B3dgm6
3GiUoVSrepavXmNBFAp247qtkl7KBRwDXgydNlNGCV5PpqD36XUT+sYibURelno5
5z2ZCidsb/gPklDSX8PAaX0Xi+TiVpBzYl3kzv7OBYIkJGDEfmVZgosxcFWG9ElC
+XLjw86R8CzyztTtqbF2xKSn/yO4l0RybM8FXXFHRaZzHUtvZ6scojh8d1+PQKMy
Pv72VL/O87LzFXRcxQtHryL9Pfp9tTQE+uRLVOAJ2ufK7rUlc2519YdO74qv7q/2
pQWF7jtb/1pg0HSRYwPf47okWI7mlWBXAEkZuwlHc9l2npCo4om4Y1zKcBKAI0IW
IB4qT6mBIpLVADtgirR5ubjhrCfJa+/Yle5tWc1VLBjR3y86PmdO1Oc3QH0wocAM
q2mas6ln9DlLkedDTSHeOU0I7Au+jLcmTK/rkZxKmF/QdTgy/0dtvC0V5XFCGF0b
OHBpqjeZZNhpnazX9Ddd3V3hq1A5p3UdPO7RYWM9I1eAn9UOL3lgj+FW35F+9f1n
+HtaND5DmhfNBnC4xJOKU0aiBooNSVN0sJuRD460fXmWjS5BuURig6Ya0yssn4ne
zquPZI4VWbXAVFCM23OzfkX3f9393+pPtyeL7tJ1I1rRxixgLii2rMo2+H/YDb0v
rJjtcfhzD7GPmLgias/bfVhU1gHg7OvjXlBjim1SBXeLIRnjmUQTQqolDKi4Y8MJ
YJfOl1ufpsXc3F8+x1UbiBliOUP3snWXrb1n3iUCFXCsTf8tRawSfRq4O/QEhiFa
oH6GbeHqGFrlw8BmEmaBDlgFFes7ffeRt6Ytg8FXjwEx/M090XP2vaFrGXTYSf+q
eLgVpB35o7/1LEvYCpvqhGkYeUuWyWewT5jE+DJQgT2fZpd4k2b2A/NocUzUZxkc
e7Fr+8G2d0BEiy3E8RQWfDAVu/8ya82AhtjZ+aw6MzXWIxgNznYM2eDPi3OUSZ4n
cPkuCjWYvuEyLbbA1PN3vAAUEH4z3EFdBdV2qM8uhaRjfDiBaNbrcZ+35VnbxRIT
wZ5sq7sTz2FT4X4vTRLv24XQvZLARVobqYvUq+xTe3XQ3IXk6AShB40v/L8+5d7r
9GSKUndgeBHvEbkL5Bu9zcjCgn52LiqRd00k3OtZLNhfmJXlRMCiG4FKF+ahmnDS
qj1S3+02wGo4dSV1OEbVGeWW0CFw+fjkVogOh2vmtY1VEILGEChZEbeNle4gQNdt
zxd7bR/PXAGvJze+YA6/OUguXGzxBjZG/6wj4A03xzxi1btzkhiGxyjR/S3klJCo
Ind5rZYpOmhIDYYhohjRR1y7nOGli575NgDz7/wa9wArNgQn+nbKeIw+uyOkPKj4
2Pa+ZasAtZC/qr6nAErlTCn+GcyV4zjdDNOgn57bvlDUaOGwY8Pl0FNylVAyLOPL
k7zOV/CqDmAdXPP5QqjL/npFnXFH0vfr4Pq0IQkL/2fM+YQLmUDcc6RV+Q6Puhyb
z2Cgb13sbX4N5uyddPztsQh3T1h2xMfbuKQDT5wfT5JbZxzcnCciImByGhauI/zR
izD4qu5jRYFgSDWWkBceNSrYvGBuZw48Wch/uyMAzggyGSQoAMqCb6jOa4Q9izTl
QgddifN9jwuU+E4K8T/4NYDc0MJsmdVOXZNHIjTPYXwxGU4QEn3CuTMFXvBdYUo1
iIpQWiSEqYqFI68TazZRlPz98aurAFRLQKZrsm+4SQrZLVDo8cFVOYxHJUiKsxeO
p64cWU7Qa2tYW0eGCz7EHoGimgclJTF7qjgSdQdD4d3q1XU6N9D9Nrq/EoA6xQFu
U1rBJyH5pxyrxDldmgQ6fImt3q1Jh1WV1DOtKbaU9nQSOONsdODB2npH+ucEFjOm
JjoqUIiD0N2L6lXvBHJ/323lSxECD5JjVdk6AbrpyYxaaNC7h1Hk3/gHFI2JnGGD
sLbpHf4nYVCs2hu0N5EJA+NxsUZMo2li/H7RYCdz71tD2DkmZTgQcGYSXX2hBMqj
8rCUnJz32d9D/pftzaAoCa7XFF0AolLxA7j7BMwvfvVrJYPWLAU0WZD+kE65eyEd
PW+nrOLuB4T2cERkDUq5hXaDM3QEHJyYTfDSyTdLF1JG2FUOQH5scmE6F2/dRE00
qetzuK4Wzfzzim4VbKosG7rCfaPMBPoR5JOyLP9fBucd8e3JAfcffMiN4p5gtnOQ
3sZHDcQDCEJhUUr/QPWNIO//d1Q8D+rsYV0NUysUIkLBxUrvxQPQx2T59sZSf18Z
K2X1kN8t7EoE58+YZXUBpcAVeXz6YOrhZI244XRCrs7MUH2mJgcOynpSubpqZEwR
/QsvKNra50g551KqZJLVhK+3Iws1sExFrPEBnZshFs1lF3/RPSZy2ZLPz7DJJTVR
5wvAmdRO8IhENqquD6D1lnv37ZQsixuVRI2p+x6AjMvVyyHHuHLaYG6yrTMW1s+O
fgitYn79tkiWJSfJJiChxf8pNjxGuWiWtSnrc9BKnF3vj/KpvcX1TSeLcMQ+hJo/
T+gwSZB0+EcIAOsuxY5LZAFClUZmHwbDWaz/Orkz4xfnuLWyBwB7zlMblrQZDc0o
zdIbtn1WhTzIy7oAN6t5zOTsvEVf3XqsU79J/vj0oMRVk4pBWgMYmA0vRQWmdRiE
R3zE0qKDKYfLCaccG8Dbkf4/j4jnk1nk2gNNtr+1zgPArkxVq0cy2flApmW7UWb6
Aa6vPMEK3zgnJteDRwUcWAFWDu3DtUg4W/PzfoKleSC3oE9ixRa/dEGHVzPyVch9
y7Aa66J/NhtVN8oqaDr/lqavSbsWp5fvlWrBRtK3UtPi9IQnQC+5PQE+s71zqvK0
CXEnZ3vor3YmF6p+DwE542va7tOv3Ovp1cPR0RrFTQMxlXOUhRdnpMhe8sA2J7dC
Is0uijQHlrTZPkeiGrmzhlIzz4jy9F28MIJlAbqaibHe4NB5iUyJkSSzH5VkNEwa
YInq8dYKfyjiQ/pkA82FTc8D9PTedUfgYM7kBw3cB8VzSTEcA29aA8oc01Da5ztP
hb+xHTpQIiTu0uj9fchXF0EnWIqyfSSmLbnre4t3pZguvH2fFJCPGLtmKYdr5qt9
SLQ67BKG+NLAe8Y3cqjuI9/vXWi3oDxmlme/7Lq06jH/tkXZZSFvK+PvL6rcfmz2
A+t2ra62rX2Suas3k0dC+EbxInYZavIJ9AQDygBUhDW+Q90T94wAynXbf4H1FVzi
5GWnLF2dJf+CPzImj8JaztdCBoNi3q0VOkc7A5tlacc4Y1EjYWmgo9AmKNfgVMFa
DxTuvffl3Xm4hiMrAZ/gzVeTN3GIt0d8Hwfvlh5HuaCfLvaXRWsTx9gtKUerlrlh
WQjTaPs3+Zj/Rr2QdfjR0kcxqUenLHF9DsyP8lcfB1IjuR2aGrrgKwt1H+qA4Vux
BSS3YK59EijLpkDCw9utKtdDom+rScpH6TqAnQQgV2JCFP5ZeuGhiuMEebqD7zgP
8XkM4h8FN2f/XKYXjWZ4X8ayo8iSFBsLefBwi5FRoz6JGVVGSjnLQ4nJW0/cQI7w
jGnF0zVUZpPioKIXXgiiyBFWDBYPutHYXEGtzBTxjeAmIvg4KXKf6s4wKBQPop0o
qYQ0o5zWl5MgopGfFZwrQyfgp0Y0D2QbUaD5IPxSBMNUaD/A3j5itqu1eEU9bUxY
vUcqyhT7jFbWaBPgXkAuDH8F1Wk7ei0TidkdL0x0sRW/aBFA4rQOAtOVUhqjK21I
gRB+yEZjBKD+gkne+1m1y9SK1VyIyv3aWEcJ9e5SkXOHoB14kI/EJzs1PQBSHEGZ
mQ9doXHDSxuNdlkTYeqS63pYHw2TThlWNZxbBiDhmO6Welf+lSzPCyVijM5CEF3i
6uyon5UhengNNhMVlsGw8Y4J/t0LpiglCij0HqsF7Fq1fzRTgpggZF+slQXO4jVm
6tcOOlDBV3DRl+5d6SqaWdfLjMiux2cJviYZR/fH9J30v20UZN2G9GTTPZjd/S6j
3+6qWFmJ3z6pz/n+mgq5wiFzqp7dSRJXS8SwP3h6HmboFqiPU9Peh4MtBDy+hpfd
sbbx5aB02/dajM5TET2pgLdUNLYZx5BSXC3kqdfUl28pCRn/b3hemgPJwDDdppCE
47UcvgbO4jCSh1ThR4hvBI7ZnLsoplRerYbdHV8vW/8XEekEweU3aJSMcvV1/YdF
4eoMv/0JxrWkQlE1ufIfV9Hfucx0iwk1JqprceYLxSCDmF/MaXguaL3OciFi9cAD
k1AuZW+iR2nzrEu0sJN8Q1dcFbpAPIp4YNZ4FNkSNwYN/pyrWIDEN5ePSP6uZkv/
03K7oA4nv86z+oz40IvI7bcVsqpLKlRIXV5BqUYfwjvEfWtOHKNYPXbohpnCmedy
RmOsYEXmLD8Q5YlxiWqsVwnXbU3QiobAuywoWu39FuqJ0hk014cRvBPsf4eTHtVn
37lrrjIw7diMSRECpbJ3rGTAXTdoCZ49UWvhMBxR4V3FfI8Bz0s9tITZ1l6KGLh6
j0WmyzpqyNKRMKqrVup/W94RQgZsLsBrLXybbN3D8bW0sjJgZP7oKAiunCM2nvXo
JX9vkzpWwz8H/2ilwZDzmfwDMbgVwx/ZA7xJLneZJ0LzRQRBDikjjxlEh+TfSF3K
u3JwigPFqCQ9Yf2Rh+RjFBgGygc1/vIFXCjV1ogM/8+El5yIStyzpSOn4SWg4/H9
UCoZonZYFPcuhCxArRIc68WNPqs8/iPmVNGVbUF+AkDfd0fHZgM3wPN9de95ktfA
BbIh1mxPnzfrxcfOpZRTawnxX07Z1idG6WstPXB9tEWDld6GLoFcNl8Z4WLdSukc
B2vVWkfoBRV7+xkDZ1aJriDZpbwEurkj8nyDzZZ3L/WBhNhJzb1a2zBPGIfXy2mp
chtWXx23fFSXGKs4UBEX9WyJfE488hnpTcw8ycRAEqHzR9OKJDfEUwndTUX2647/
9y95bAemzNDeFQjNp9achjFmrb7lxlAa2ZYPzsClGqT15P4gUVAhfg4Squ5/xjTg
0g5KK9fQomQNWkUkJjA+Zs5xjru4ewq3wHZ255ahX7aEMdO1Hu8f9pWcP77VCzm3
Aa+l/K66o7zG7nORWMocni8mHaizZJRpyoIJF/IoL4+l4upFz736PTPzrbNk+QIL
hKN2B6+hSIlDaVZqFQrpY9EYiafzZmDRslOH6aUQ+sxI/lx2Yxh2h00AE4mzRxdJ
l+O1GHjsJs+LugOC1nhREgmFn3s3ElVtu5ioBsoHCDXXLpHZCtIG7XhVzPbfQULJ
Q2MpyzR1oh9hc/RJgZd7GLyg0JLHbQTnKZZzK72nioe9y7rPiUwdREtoVEsWVgR1
LuTpBWtiAZl5BSdOs/JNJTniAdr24Lq4jbz7/ldT75U2HtzBVZteam5f7ZZ2GpZM
0yMIpwGvWclZS54DxRVLtuSFwKKqgnIaAQtYRONToRmRVLus3JzN9pAMNFR6zCKl
dohezT5KFtc3ytK7At0Ozba+Z98ER+nRqyxCl8qf6a2fymuALpYW5Oy8tbAEPxQp
hFVygv/Flhcxdr7NNwSMp5s+v+rKW4rIBIkDCADqARzmMuQF3np0rNoFYE8Ks8ZW
+cQ+jNhPIvGvu6GZVLenNYc92caff1ZBsnwiYHV4Wcy4WTypAO69qCr8fci2uZQT
z/AaKOGtPmPwwzPtMWGYX5dwtMj2u23lg89iQwqEvU8xJfqB7MBpRIU3nAgwmxpR
ezXD4k07cKykXO2FK8lNBV5AicjomtQZpnQaeS/idCe7OWo3eyp9WHjCZeXHKNkn
fTljh4rqsqnA7Yk6EGXe1jqpeVFs9huj5Z5h563sv+Sni6nAC8vnKgCzap6Lp8lX
HaYyCtx3w7cCbso+YcMCWuK8WvwUsepmn5L5OwN6MgzGdYYijd2TOGqN0Y02i15v
u1huG4fHYU/8MIEEEwicjE8uZQe9k15fcHftuaj8CwoeljptVxOjMbswNd5tB9JX
RrH/GLqxWf6lfH1FYO2AXCQsUKgtG07Rv6puv/wcrhZQj8GsAV7UlPbq2Nfvr2hl
tLNX3Hudeql9L7dMsIxBJIX4GS3mGGC05pjZj0rl8GPmO2S7Whn/JdBY4fEgiyno
53HeimrJCyv7rO0A+wr1wegJgsUNQKVnypPttyOTT5ys+YyXnZaP3Btd3fwPTGH7
K79qUL5jCzrO5H/2t6PjZD1zxwmTGEO1qUmmHmEGttULtISuKcWhrzkzGOz45NmP
4j5H+uE1wKZTwyccRk7d2J4Am9D9S1wz02ovXv1lARcAc4gTEs4axbEyd+aAf0na
Y0CCKYCEejW5d0SlhyZ7V8VEq7hEnJYs0Dh/jAK54z6TP/Tw2ILNf1SABlXuQxBf
WsrxZWZsXX5v0JeoXv7ccmN9CHH5FRP8tIwDoT9LcN79B33dUye322oLhpV/J9Iu
qVTf7H6Z2pQm21bUanmECV7V0lry2vrFQD7sBbSi/v+iWdEcw16kvnc8WbANA6+N
ftMUyITeGa7iM7WtKLvGcCphPpfBa8qA7Eddsn30+hJ6y5MIML94N8PlZypf4AWJ
8Tqzb8RhMufWpfodlquSbGppqmDUzqUYQflXWdA05BXMvqo71dllJiuE4wILu3hw
ezffk5wXmRY3oAj3O9CvfSx32pebPncTy5mc45Iofy6vKoTJCaE+R4N6OtijXN56
I1hhjZA27XypB71A60rTCBg2Nnr3xVlngfNkBRIxh8OspgMfutuJ+2KfbsIR2t/Z
x4w1/wKi0ZMg6Q8IInc7+myuNSG7X8KSKmIQOcqAHuVcwVRTdq0jJiHYVwW/AgQn
y3NcYYMSCEmarceeV7wTxoIHC0PGcyDtibdUv65R0LCNer3CJCfHkp6hCXf5OL8C
1vnyGeh0l+HwbT1h4usG/HIW9NiFxi9SkqTL6mTTy14uIOHvg/vcpstRsvkiWP35
jnfnCeM+rJ3+Xp/pmfsbFA25RnESTBBVhNWOqIstNViDvI07Fyc8v5pNGYzXNxYD
R/gsoqTWx1k7V0QkldCobafUkcsto75a/E6pKhcOCKBgoYbH4Evvnad160EUtCxE
B9ASOs4xcc7J1HgGLZPTHhzj3gKgi9u3UnSovOdQMof7JiHhFHKVDlCcAz+E8RmT
L8SjsHqeLQa04bhTMmSgpBoq11ss63zgzf83PmL1ncxeBkecBAMUruj2F5c7AN17
lnRjN0TFYtKTogVoy2c4Qeg+ev0RRnNfzy376KTpeZQJULfMPT9WRshoMuTail+H
tXGWOd7HSRt2hxNz2zyeV5Mm/dKJSollNEhWf1zTYD4xpI+6nLjMHIThLsNaTEbB
FH3bXAoV73xm/G2rlBEjpktuCm+VY/EWPunxIChCmfe6dhciThfLN2tB/5bEeUnG
sR5P/EoYFYjncerg3anMlBQM0c56jbnNcHs/EmDswbNT1hfW2hUZ6gP3DjICtDcS
8mLmZ+UwvCwgwl2Psu0o3NDgbZxBfCTwaKwak89jYhUVnhvhMj9kKhAnUgpFPGUb
nf3/29c2YixuTzVPLbDIcVkOvpZlo++zZMhfikKi7THQefTU3HIkTIYTw0QP6ogy
VFa+NZo6z7ZU+4tzWoc75DIajn9tH20ekp3oHJqaoStA7FHKw4cqRZSvguO6x0GV
oFbSDQlh10VkMZrJc7QOumjLeI6cxOfIpJUwyVV6RB0uPVqPTe/g4F7ltIqITqwL
AR1TdS4lRATEG2ZSOWF8sNOJXqdxwV01zHi9hwNHEXLMvPoUhvq1gLj63oUgZcEu
z2ivZdvu8IqHazQADTV8Xrlo1qxXUN8HQ6frh/g5hVWu9qO1baC8S7NKtQwJKXbg
T6+R4U1OQI9/8Y9J7C7w6PeMvLOP2lQp29eV3fs8rV+3KFtUD/SIJ/ShWIblQDdW
2qpOivSPC51SYFJJUA6IvKWQXfzOPjNYWDDKioKg7ekJg1TlJB6mtCAAgDnMP7UI
/OIZF8juniGTNFtV0t5rPt6CNdCY+YtoN6WH1wsMaOUQwCYzBW4Sz3fSucWZpY/7
mcGDwLJl5SmsPDpnOzKIniaZrWPY/pNY7sD+RSG5uDffzwMbySvY0XFzO+7LFdRq
9Lduu0mL5m6vWQTvuOHkvhj2aDmDcnHDDXxC7GULjFu36v+yWpy2KxsJvbw+a4zS
IOccbg/G0bZWLOaDvZrEfCnA7Tp1TgePlj+/nHYtLqMJGpHHlxdDqlDCoy1wF9Lu
R1tsBMcf8E575AIWpF+n/039BYx3nUZLWkRYQWgB6XFS7H7WOFTCX82BFbnRR5mv
aZryjxEOJgF94HyHVEUYSx7y+6HRSd88B9+s0kNVBnqcKdLgVnWAt8VRXPzBZfHS
x4znEzsn+KI0bnKag4fNTYopyV/homIhZxIFYCUs1kLG8j04lYLbMN3hnakwvt6f
6rOb7Rce5nDKmA43lLi2ViQJLDl11IMn9JYqCYE4fVcyDhHarvmuTqarET3xlrYY
RWhD5LGvVFMpOVy7tMyNCdAwBI2vi/I3/IDRzMKO5FYi5YHlcXkUZeAfysOwLufs
gcSMxAURtee9nZGlXW32DCt2AZNyt9LIiCgXvoi+n3xR7gZ9j+V4rIblE1usavSg
p3EwHrQhkcsrPwFIG4wphJe02uYBqOeTHvYXR4MghFDbJz2LgKZVofwaVcScAePU
UXs0RtCcjUeE9dInX0NYcWb9Bc+4vw73TKeRvVaTi/alz2wHvrIEIo3PcRXQp8or
FHcJMBuPrJkSvNdnl7QNqJCpElczV3OfYM3ADV2j5KkWmW7VitPeilTam5N6rA6a
0j+UY00tNLJC3r28VgJW7kgF3PCdTDCuVXcWOS+pHQRQWbezmSaXog2ZEGhvYkGb
JiV1mKAh9hbib3CCUOlR/diL/FdN0y/4PGx2lIESpgkMrKKOZ5gdyp9moknzgOUy
ocMfzv8jHSmNSsKhV1huHnjsA3v3TGUiu689NfTR4k6hB32vLfcGX+WKPHqF/1ie
z3XeUV9w2rnrHbqZ/VbOfwI3JThWb8CR7ccOMayxPMF9Nj10La49MC883YvAyTgM
c2QmTpBWCODZlxI0+5Yi2cNS/bQ/M2C0lemhVyEsNQ4qV8BdwfJ3w4uNjauD2Onn
HuNVtwjt1wJ5c/iwMaIm2iz0u9rjfiMHCDZN4S3SWFzEUBww4oojqiB3dd5Ku/u0
tKBkS3CEH+IHsgtESLetbdFDCIboaXARHTFzDC16K6SeiVaKxhy+dv3xOXvVImVI
EcMZMWX7r074YUnQymvp4pRFwn2Bx/ZHUv2oDe3F0fmZebgP4SltuQ7yFgwQyYd3
extZCK1NQCP7Jyac07dqE/JOqkvgBq9UuoeMSWHswJDMJF93CHE7vHP6CBwQTJhT
jOpEw9CMUIiXKMlnVBH8yKUMPPdOfnsVpOK3oO4Cs/qfyjD1/3LmG0q9t5V6BXMv
/1JhOQ+NOXZDMK4CNmncOgUIMpXh9vG4asuyLIpj/4jXurdHzjHs1fS7j5oZb50P
+xPFfVpiKnXug+9M8tb4mLTieVyFZY7R5aV0ahE9BrQ9WYyChObvhxgzbCcVsato
ZBMX3vRqPJm0j596tS3Yj9C99nS6xa3lsj/j0/Iwz+5vnBS/0nSD5rsTxouTFh94
HuqYtxPfHRsZzhXM4NvEIdue24l/LjfzEJfbLGslHEH+g0TawvOdVlTaMpWu90+b
ls+HrXv9GL5p8mNgs6gsMAZauxSdpyhS93QZEQtIkjNqSbPSMLVLN6Jci8CkE8Vw
uh2ge4JlEWUpaxu7KU2tSE7Mp0kAIGWac2mwFD5RBvLXgTxUzsnApUlKaj6jMhYg
oSazPVcziQTbkRjysSJ/yK4i56YRlbYRgaAp0Ium9cBGR0iAgcr9L8pkkzW2IYlz
IrUeTv9KHAOQpygGlpuT+hBDtEMc0a8tppZzrGho+H2Cwm9mVxdl7Mzr0Sg2eeXX
hqBtm8zv2gWzXDRXLFkrBJ0XUCCmVn9872+AWokjgaursYu4kjFJfY+4H+1ssy1d
n3kdXk9tXxt6NOY03GOvX8bMaG4ZK12qMfaN0IiPwTWv0U8k+meKR/aiLsyy/hBL
fqfC9Yx16OOhLcWaBx2zKtzIxBN7s1+RzWtqj4je/k3wI/s3dqOMBL7wGU+9C+zE
sF3sYjuNpl7kQwfUVyGRH/Dqcbi81Eaqv2pnk6vzuc+/70yHIz5ZtI6uIjbpEGX6
Do0KwRynUGySBNtnNZoHmkHe+fGKambGJiS5Gb8DX2o4H1NrmDd6ipuk9Wp4U1vm
RRB05gbFXGt0aVjwiHiCeslcA7V4IZO7bZuoNT+O0wyl4+U3GRnVbSwXIjIo7/nx
7n3ffPp5z2p3BSmYzJ+UbOC/r/Z03Jm0lTTDezOI0Qa4JaoAjBEg8sHLHVKcTWkk
BaGHXWbq0VZ2/7wRL5DUqgCjzH5rHG++JKIfY9evhSVw915f6Lpt75ud3xji1IRa
4TUBhjmvitgYQufMm2OAdPKCFjcP+9TOETjBWHL1a3qdkgWc6+LMl+olnSoCut0r
HUWakaxrYB/OujAGnsYHhxv37WQFeVcnXuUtNqpoiAIQ4m2W29Stk5xm+LftFWHf
ReEIKXJpFjTyPkieW+gLCMIrau3NZoVSRSkGz5VLZrG3cp4NbR5ILg5hsU0piSKY
WPpJC/LvAXF+Q98QzeEcYHS92C2tf146wOntrUURb73NIdSVMyCPuZA0ffhh7zj0
jlfT9MgSpA8OjP0kKEQpY4CU6glTjKu9n+kbHiyEmp9tmohfjk7BwbKoGohjdyhF
JmjBCN3YYylToVvVN7QnvGqc6pn+oDDqZh3CvWxDi/AeUOWZ65Hl1VdT5N7zlIM3
RQMFDhccQ9wAQh3N7XP7HMq9klejnKP/4BPMf4L5JWNltCkwytJBI8ZHXc/GdXkH
gQ3H9al/B62SpR4p0wTrPiwGXSVQJDAiB2DA194no0f9LrT1yvD7+LXWVPx9LgDv
EaC0muhEwQi/cRb5/CXDwCFShHoJs9wK6hMAN/dALMawARiczwOSYrbNAh2kqkp5
kYSxJ+AjIEIo9s+LW0tHVoQzu5sBcWO2E1MW8Q2HBJU4NR5KS4nOAtPxe/CdkpMf
gpWYPhn9pee8ZmcICXvLkx6cItG11kcDW3PT5yvJfzWr7FFHV4hQw4M/YKgvqk/P
cv6FSAg9Tj/FI7bT89r9WJg4FFEj2pF+rH66DTlQN6Egm5QErDwtFngCg5QIcc1Y
5sTcs+WHkd+uClL0lnSDJKQ6ZK9eSTlVY0HBED4josVNBS2ZIQHjF1cJva2MNMsq
mxijHMII3Rr7CTvZpUEbUSMW4HIP9NVt0GXsDpYuE9Mzmsf1Zf+cimoBmqI7DOV+
S+81oB/tsnDsB8jyQthHQm/S6okiPqcaVNfJbFu6hvfYfJ9VzYhJeWbAXNVuiyYe
5iXhBoghjRJG7b4DwSTduAwj7XH/ZsxU80sfLMELIuyON8yBjOgIWWHXDvRMW1uM
gAsXIIMnewwYHtR6miwcq6Em50R81WPeqqxmsRk3ax5zekvOdoSAin2CYqRasRYp
gVpKOfVpX9w7e7yxu/agio+eXuuYAi/MVipxsn+RckZ4pMhRPjvi4ic1hbeehvlT
5/hYUPRWkuQu2ROYxqSJ0pvWQXiOPiyzvgOmP20gw7Pcq5WYfJekKDg5rEV2tFGA
RdS6QD8+wiMIyGZCYE7VS9HM9+0Hw/xHfKtKcdo+itmV7yxncRGdiuN1YjcaBJHr
Rm5YAIUVt+gAov3YOmXhLL98GRQDal9qEMBE5rtUqKedCEcfL4Ax5ihB9mr8veTf
N7lV0Tp+hWnRbLxsyDJo/GNCI2CTyEHhG4vhAh6XIk4I9I35OxKSOTT9GU0JANKz
eqPjJbqvxJtb9rBKdFGvCERBuXgGta/ebCcSipIpvMEuoXz3sVKBaSIT4zH5fNIu
V6gPVQSdiQptLw+1+ffLv5EqH2kdUo56tVpjlR9AclfSStvY/TdKUgCDppjkhf3R
NABJ1WuLJF7A/fF+U30cAI+kAvmYvJFv4MsdSJPtdoTCA04Rru6Rlw4/TbieEknS
kQsIculyvx/XYFoSXbjP0OueqB4NJl/BkMReiI53YgPkB7PtHIME3pb7rCI+lu1J
n7hT28aqzozYfSuF6cA0UCKj4idt3v3F3xf09fhbojpnZID9OnUAteSr4yfMYkBE
uCfMbvSMQexbVcbvTjzxGOOGqvNs7JFz79wfkCMbzOghrATJHgO0EA3QblzP8fkL
HEQRBlOJofwFKKR7p5e0Y6y6Ivej7WkQkJw3hjy0HMeyxkK/v1v35t2CnMO3BPf+
QqoADmD965w8fW8y9kZP5xNjQGKvVVrfvciEm7XUtBNB4yafd5T/nh6yOIcAMWYn
IjIgNZDqwodbgVlaeadmeGBeK1tC98LXHWeLWz8cXKIHTm2s+6pG/7PJlZ0VWOFT
byOsVUzzm8ySCrDllxLaDXX4GSuqD6XuvjjIbteBbPpkAh6ROIm1YHRCEtImUOZC
8DOamnMQpb74Or7GMCQ7nCVZ2AhDCc0In3kFiO2r073EGXcDsRr3fQqng5cTk4hk
etnuPkjFdJKzuK73KdAEOlN4IjnBT2KvabZBUkO8o1uptXwkv35fpzmvZcAA7ctX
DCaQ/8vDBVtJDYX7W1GlJpMuZlsjpBY6QInCld7MN1rwUmm2kQBmgE1SLW5Jz2D6
SAK0pp39QUD3lepxRC1jErBpOD6Pt64a2iixch/kPkECIqFRIneWFeJsEY970D3L
vKnFISzh13O2xO6pUrc0XQqSFHlETbzHGqcpMHppkwYJk5ux7U2Ne2a5RZwq9OHc
JQz3rmX+S6pTeVJ6x6oXjwjHIsx+lUl1utRv6WVZASqMctR3UroQY++kPy7XEBUC
tLHKIunJpyv+0GBUZtFGyIUPL4ywZVGoX8ydlUprzfqXzLOx1ZqtDwj5IyxKCXrE
TENeBtK46lhyn7e0vBbs41uJb6aOpZJ/w8CA0GHeRxFo/cLmb/3QMhRUXHLEzkKm
66J0DXCogsmQjiFNgCYVpUn/+i9a+gbwsf5Dd5DOIXtklNFcDjs4eWarzkkBs6n8
iRA0XF24KhciiFv/2zVEOX4O4k6lJwbozAu3SgyYYL/BCBFa+4p7AtDnXniJmTJh
C/jxDHgwDpNMAxS6d4c0jyrXNiQ8lXzLkFLpCHd5JSp7UvQc0xWS2WJAwwfD1DWm
Bjw4fd0u87G2q4JyA9UYB8dGb5MZ5sGUf98zbfHp5HZoE/wTTJ0DIenIIWc4laPK
c1tbKY1j9Vh9TJvGunhU1nRThrCAhALUdv1q5nllaGU7OBT+MJzwqVF0hyduGGU1
dA4mGaVw9C9qsSgw5PTaOTxMQJq0qRfYD28XbR3ZhYEJYeqFFeLzn3jpjHcUgv0T
QRoa5WBlbJzpFMx/CtsbNEUtzB1MTwXr/yu2g/AgnXNaGNiEIz87XQqaj/p3TlW5
VBzGbJko1yg0bz5imu/1WTx71qcdj/RE0NNXn3lNaABcCec85JDf2qX7KEDLX1Dt
rFqE3GCcjUDg0ah1FSCr1OPOAAhxsjVUJ2E/k5HoeInI6XUwC0yRoaVBtH1estmU
a/Q6rgyUeWqsSmoAN4M1h3Qmvt3IFJ629/IveaZIOkaF8rbc7dxwwC0Dv2PaNZ+r
G3eXXD7Y3OKQ9JnNT4jiuuMNkeogvbqh0udNYTei0iyMmOGu+tQ4FKuClzf8qfNp
Aeu4HLyVf1VJMoK7HvkdcrnCxVIlcXoyDBm5JPqmS+cZkxnpMGmr8ss8kbgxO2UC
vQ6Dgw7SITuazVY/1C/tHialihgM1Lz4fq3fODKwAmsA3Fk0v9OOddM69TT9kaVP
SVPgkX/uMECF3pRJyL6ASJ5A04/EmI3MmxnR1nlj1uN4yPLxlaJ00Xj4Lfu4WWpy
dVdG2ykra1x15PfaWfrpkGaf+pNzNE1UxbEswbHZnwxLMZiORAAaujt3moby79/I
cfiGroQ7Wyxq3bB48J79vH/Rie0B/r84GZ3TrqQI/fhdY5vYMXMP+BuX6BZ6bUki
8Iqd/SPL4J1OO8Gs1LdezMjTITjCLG+5ka1bYitHzh81xSpkI8vzm5tHZlvlu6te
qdPeAHrbZSZOT+B2g3rbGNQo5eQAE3xbmbxLce+739rfyzCZ3SKOhgJ8f/JZu7GX
oceIu0UPrK6QbNhUmrcMSMg54lyzTGHZw5PcX31o1aCwwfClpx3L3b6nLgJH0Mpa
FCGR3EPgW4OWtqGSD5pxqmN2xHVzWNizM8Y/+U10Uv9/ZpBE3kAljCgXWkN2bk6+
icullwnF9VoAbxnUHY7fdiDxJqRUZWDwbiRiguDrwToS0nRfSShL70XWFCjifBi/
jsK542mpHMuycWlb6jsZzoRBwkiujRJ5ovkhRFFV1w7TRy7Y+1SwgdBsILoEe/kf
1EP8WzYEQ//d8/R4nzqDPfDlOOW2GAn+IvJnvzptDbsFl3iNuJidxNBVrldhtI+E
NvlSAj1WaPFy+MsSsW8VUdjdTRynODWxqCidZSt9TeiZ7hjzO0c0Y+X0UHPxYp7S
w9GAuUQsR/H3q0MJYI4wzqB5GLpr4rzyDpf4nN85Hr4KEs928G/hP79UhwyiTLDE
95Gfcv8BtCT30sAo0omGRA3kRu3MMp8+WZy+X2jpaD21Xh1At7vMBry136udelGl
3epD2S1Qvs2rCK/tRsVQ0iKDTEakB2NtnYfhcHwlgB1+/ShhRLXoHED4P+2qQq9+
0TDETktxskbwj5mdOoLHxcxNXMQeS2q7ZuMZMKuD4gcuAZDSiOMAWCN1wEdYns43
sunY4fo/putQnhnk5m1Ajhe6okcAXtiE8bgrrGUNgRh0JIkCv0OXM02ySTRYtWZq
+xedLKgqGBPI7FScIUmVZW3cz1JARtFLFVBZTCwxuDtYyoHMpEaicOe3NFFNg7oj
e2G75T+WLYSAhS+RTdw5t/zCB2RCHI/O+2buVdFygpn0eP71bmydda3cIK+quX8u
T2/+roYxh5YGUxeWa/9J+Fccg0AoxcJxLDewQG3VIszg/YmrAziGPor4QxNkgBgC
0CswrfYHZ0PqT49gGiKgp/nbzObJRYlhVfg3Yr2EsJlQqoiSHJtv8uRNLpqZkxFe
UC0cgDUL+UBI6rmemsFyKo/cyyodnqtn3t5BuRA00cDvKuZhdTvhR2yDPXWDASL4
37LxjmWR71XetiWrnenxvvL3RiigOetbsdeGHLVQHgGoazhS4tPOt8Gw+Jilk5lo
gIg147Jg98hRAClTMCTBvqB2A+ZCv3aLRB/ZNTgRyJjRXC+0IJkQg0w3RNcTp14M
mIR+Dok2p9qv6SnzqPA9S1/zh8yN2Q+iMiML2tqWUkvdVjsQjUaevVkqF9bLVAAx
9Yi7brKvSrmcN0WyUbh0tQ596jRSmrsG3HMsU2if3cZrU6wjdu+ThaT0mr552dOw
N7J5nE0SoU/L86S/4VzccQMVGY+GWs86I3clTAYfSyIdjhu5YDK8PSdBG1PBxsXQ
n6r83+KpAqnwwnkWo9ybmQe/nxwDy1TY+9n5YeY/07VAj7tbfGnCmxEIxBk7fLZQ
XrpxJC7+OaoDI7GI61PuL3wwYBaO9anLJK8gN1KO1sVm5UukY7rjHg2GpvolIapn
3X6ernm+Y+YPWp8fY2/9kuK5WcatLlmR571QUW79Uk2lh6VejgTWe58Hx7tsU13k
Hkrhut0vdKOu93XmtfQ9vnFG1Iu7L6NYGwH3k6C04OfOrizg2ciK0iCXzMAabGA9
dGIlwEpNxAEZM+e7aKsF3ZibZvUPrg6KlfZZTiFxUpCrX69DLqJqcFDQ1pFuloXH
3ADQyeWhFVT6/jOgm6moZanGLiZZPUnrtxg/VGcc76Oag4Cnd09zdmOtBHHJf55F
BByegzSLESYfy8mTl9lYlrsb3RFay03prEdvfUahZ5O84g5Z4WCeXXqjnOBpHIxK
06AfE3gZw8hfwJFop7cSdGnMve2GKQFsLf8wcAzwJnuZJmY8x16/YD7tw62QztGw
agC+tnFnvLczLeSKYQLiveOlQuuQlPqMoGLLAYfB3EvsDC5fcMZ+yDcikIZhR+UG
0y7B0Gqf0GjxATaUUfztS/9yVVbkKGxYUNl3FmK1DYrnMDzf/cdQoHurKGsWI9Ut
9MZDHHmzWcJDhYeZ8rY/zDjWtV9oeS3tS9dMjmGBDD9KwwhYOsvK92p7hlxV5nfZ
JaZtrE16M3Bj81/ko+FV0tLdv0HMXKBOXN0kpCfmSp7XeG+/QFt+uNosp6fZ+FR1
AFx9BFK8NF5pZvEAul9apZBPd+3haxBd4/DNuUFfYrQdB7j7rQXprxlcjhjJC/Fz
NS349uihr2CxqbYev3eS2wI+I7hDVfbYfV6OlHhXV7MejCAjgCstlX56hlVM6P9Z
wSdowkRHxouSwgst4sg6gdSWqPgVjUXBgU2qwIdogBf3QwweEYLLrn6lbi5BBjLJ
cWDuO0PocyFJEWXdNnubFi8AQB8SxTGnCNfFrI3aPEBHR5sWMCox+V/d8dn3woEf
ZhrZjtQpKWX5xpKaAz2RVijzQVeo5BEIaXhi6+PlcMxxUFYu9PMUEhhDSQLC9vXd
DRKZlbakJWXd0cZ9gTnTiS5SwW7x9uXiySxNLpbu0GyATQ9LIGHrisgRMrRZo+ya
DBp7mr/L+YeEcJD8oDbPXkSPrvFEt+SdZtz+R64Xfzd5j0EubC+m9EgerZevHHA1
qEry5GjkOSirKMgMjCgKL8k6uQ5ABi9whFXl6K/lXiQY44OtWYsDE8a/J8pLFCwj
kPdOv4t+HBYjhL/rWr3moKsCWvtHB8g1WSJEB86mI1gDo90ZDwg1FowzPxV0qYlL
5pUXbsvebJP3qAupzAaqYsXhJiwwsxYdP3u4Yrcf17GX+E2DBZ701jbFG2K8TmTm
W9acKXZYJYQ/vRKmvhz42AOC9iE6vmWljoPnS1vu738PrBKZkV6aV2FwmKhqEzqa
mTaekxxElqrEmRtJy7sPc8elc6EfYwmO7PqJcNhNHmcN6hVouphKlzOaXJ5yKkv2
LEc3YHXOkL/nnx4U6bs6GmT+YUZBZuk/zEimX/kf+o/xVbUYcNdiM+dpCUPAZgqZ
rZ6NLFR9gs+risogg40iJb/ak8J2Epi1iIzun9Y+cO1kUJa7iKYcWQxE668cxOLG
vWpGTaQNM/g3lCJsVjTXisCu1ehZKtu5QBPnJ4Ui2OQGR8iOCVdt3dBxnMgiempW
bMRXG9Z3JFxOr65Dio3nc/80RXrrAWxE9fy0Aw7tGYnI0aXAAIV2AgkXbTeFNf7f
EnJ1DkTwMrwzoadog4SFSOi1IK9jQEzd8h+3BpaJnj4H0if9LQrSz2xCv38/FVyG
8jKOxcXlVh9P7Ve28a9jGrj6tUpdwCK8B17jfE0tWFdKB1lscDFtk/Qt2i+BC3+m
cI8VumfoOBcVWRis8EhcZvlsQq7et06TvmUvuuBJc8hQh2VF/eqZb8gKxzMEvM6+
h5KutADAn3TDA9VaOjHuOrJiRrSsdzQ7G2V2rwLc/rrVS/4a+kuSQtBimxv5uhxA
yK4PfTeC7r7Pf9rU/OGRJOPru9JQHbKRQyTNX6/JF5XEplti8Nho0dM+cV84/Ghf
nPS7J/QHs3BEbL77ahRacDJzCmoVmv6vPbIJ8zuehVAqqCFVD4CLy6utLo6TCL0m
41DeJ4Tjz/LyOXCCFvxtINMHA+DA83ooJntduCF/YsZtxeNEAp9cjG6umsXO+oRh
K2B4GHc2j/Sz6sK57E7naCyq+PqS7XMU+tNv/WSQW2i/WJQnd1UbEawu03vvHYHC
HzN0YTYeXdn6BXM/Ds+7Wl+DPjrKHUxYaZpqtY2x2UjvvJ81An2SG0RyUrr8eHiA
Ly0lr+nPD+chJqPjzRSo5gnX4+9C9Ps0YwP9zKE00os7W0n33eNv9xZ99GPhtGv+
CjHYJo7jEVamtsKZAB8Hs+ci2IdlgOhKk49MJqzEixgM2dpBX46UqCrjHy5Xq7lh
4ujFfFK5rI1aif6lZyK+nMSFBJnx/hiwylXdD1JaaerJQWY6DdmJHHOESeleo7vX
LKoDmeRrv+rxJhK9ygDjYd5Va9184YFlKXxXQ8+jHjNV87N+nyD+/gkgLHwIs/Lz
azYuEI1HEkhz1OE+AApaoDI5oODvqx8NuUysyt2TTv20Jk11co5pIzT/AQ7yMcL9
AZ7ZUVlq+1p2bE5p9DC6O35phXpk3omh12Epa/5KY3flRXYEeQTXdcC+fS8ykfU6
2RABZipkLj5Q4M+LWR37AWivo+hIShvrktYnKGKGsyFdRmYdCRwo8uGOcae1iENj
Tk4oojrB/H6Gb/CjXFf3Ll8tsdE89mB9ZDw5VNe6FL6JIqULMo7VMj1HmQuqzYwa
U2b4c12NVBrMoJRF1mTU7IvXjPe4hOv7mAjxFqLzNvC65fOb1xZY110AfNs1efss
puvhwVww52TjM1Nes3EEqH1XCyv63UFFEgFIrFCviTKtp7U+vwgN1hBSLsBk39Kp
HnERRGS0bIc/WYSJdRt3A2zI/E6klQjDrk+RW5VvguDdWw2cYjq+5/UA3sE5JYua
F4m+x7jFr0VPQMjb1Td5uvLDuATVVUhDtTi8TxBsNKckyl2yrP0DSlbao3YWNB+R
KQc+Jr9qy7TKrEi2QkkuRw0A2wHDX3Z/IM0e0QdbFUwKm9iQ1s9wd61C7spD0C5F
9rmLo15kEQQNz8UNYK1Ye9qVH+Y/KF2BK5iXOmA4wO6oceBBVp8YNHnftouVuL0D
1pG245LeNm7zclKwzKJJtZWFTZDNErdKEvVXCNYR2MBcCin138PNrtW0vmmH1/6M
v+KjXNfNajbk3IC3ZYmZaNQDSr3Tx2HrsglnwZ+f9Vuzio1tlpwHmcefC5/leHKq
hHhY9WZMMpUX4X0cCPGZGu5iG9weWPQuHQTtpFGBPid70n5ALD9Dd7sMD+Bc43kC
01cSVeU3k3f4O9+wh+yuKXki4C/hz9Roh2eAwhq8W3M/0s9m6pqwD+EZp+3JR9vs
YrXKLg0dL522MKic50mJ7S3kx61eUF80fOqsAJImc8+8p5MXwwhWlUoehMbHGdI2
wvCKk/NiaVwaplZDeUJh28x14CvVNyB3I2H/a6ChdHRN1d5ZQtk4G3Oma86OFvpk
JVmG5mCzVuUFO+iiW/x8AHX1XSbKnrGSU1MA3hKMGcyx6Mbf90FovKFJ+/iqJ1K5
XD4WBfrfyCw9/FqQViNcR95uMMMuToGz3hZM82DyS2UkmEgBfpFBM+/E2WDAPykS
ifv6rfCLtbweXjicoSWr99Sk8V+/IjmZAQ8vi2iYWdgkwvtmVRv+IOr0CUlc967h
qar68jxg2CeEeEF+YxeKSgH8RSPzhtFTspO6nfxFn9PRTCq3tkDhHIMKsLlsXMSD
pof7+ZhIRfbA7qocq+ukb8rO0qLmdH/HVfHkO+OvulAowl+22zOaoiZBJBHfKt5I
10FtEUPziIQYMMaNrhJrYb9cYaOLQtKMqzrWPPXVMVS/gzxdqVKK8JL79oj5vnM2
6PNOGE0gyFZ4MrrD/Fs2CdIlDohZSm3/SMIP0TFZVsn/UQsdm1b8THqwrc68IKwf
EvvdDhqzV1fc3dD/xIgpQ1M87YchwcGnCdmlLH645z8+716DPN7tzZMOnxd0U578
9/jQTZw34RnVwjXZgDdSiBy/rvyAg17eb06uWzzvXHJnyV8CINi3BBzOMH00wQfo
OoSyE5MVefMYPahfthRsXFxSooOg0xJ8ASdUdFSpUIrlMocCAe9US4sFbL3kPye5
Oeeed0qC4Hejrk97lNJaHmxjAAu+a5H6RLBB37FPnOXxZiBItm6rL6SEhjU+am3m
QRKKiQGhum4k+5YLUWo3sr0bQcdHiOwPyXiO2H3/8uwlevY4CeUq7T0u3vwXIl+f
ut4DQThNQsiFcDJ5mC+Erd9jGOQk79Isxf1oRLDJVwWzl26/OlTpUZ4016MtTL0L
IgktQJa2zBc7ag87CjVFD0B0D7vsp2eFZvpAnyH+sACquq5zOa75ooHrbcZKcqcJ
4/zwxdqkb2wbNJp/gB9/NgipBQnrpAtu0DjHUZJQWowfMmpg5d2y5YaIkf69s5O/
NnexnhOdDGkyHQfVPJe6fhvlI7jMXI7Xi5afVkcpUt0cBFlbt9jdu0OTO8jmk93x
LDlkOti373x8pUD4XOhWkj+hLh2ctRoV3KqOzBLTpDJE1ndcB+wEobmyoVCHmpbl
gTcmE/GjGu6imZh7Cy5WRdNa5gmVBIrqapbzSMFcB3DROWXbwkpdVB2Ks4eSVi7N
M5L2lpoWdwsWZjRVr98cbMPQzs6MrzobFm6a/QwWRitjl0p4+McL5pUzeBJxpT9x
8okQT0KoXVawjjVa/jLrXopBz9APxF6iR8Rhj+szT+FrxPmIaNpvBEqAPIb29Npd
uyI74M5Hl7kqZbBPk68BHKIZhhyGRigoETSfIIKqdNELbMaVey0w8OMQ+zfAUCg6
4MxEpuk34xKwvrsivKma27jtUrXMc+5g/0xKGhp1BJis5KCbhe70HvAhevBDDGdG
90sMqnf5TnM12afrsNHZqL87OeTomT2ecX+fZy47a14OK2HXvWSmLamDS3B5hHa6
FqJMKeqd0YbPhpHr7eJqEhaeQlrY9mw0ZoCVGRdnzQ8rEs3meORRpQ1rSlzpv33D
fYvPleV+2mj/aFiYEGSxbDiGCsuLSqwUt2h6E6ikLCG4D9ew6u3H937dNzbQrS7h
/d6kiRUuzKEKIPbfJrcXggE8ge/zW3AOY4uYdfLl2PQ/AHXPQ9pCmBckpV8pW2nn
5umxzLQl+YbwGRQk17G5gbl6bct4Us33U30GwYoMk9eduIAUrToPf37+HYjEIgL2
GChTrVvMoYpFUsWKE+0DZYsqguc2/TBEHLGu74fLOs5ll1U7KbMSYRYmnJAT5W5Q
2DSe/8lZhqLRT6aqMfdtOovsgyVb3CnPuYO0SLfI9klzr7vUTShIVqD0MvLWS210
8ZFlZtJS8b9LpNFO2rmrMrL9mpeu/jS5xGeGwh0Lnk1WNtRn4Lb8ZEqSCpZaCAUy
bXlF/yq5fd9u4+7VzULic2lDbV1FDBSaFID009gnQ4FsiLBiHCUaw9Q1+Rb82gX/
Q8mL81o0RpaT7xC/wwGCc8yjS0ixJO2qT+FN0I3yPJuq9IJQCeblapNxP2pL6jhN
KyVVxg39M0A38C3YknTnajsq55XESE3eMT9MjP1XZzpAAHGhNRT/JXd++lXwsRfu
yaMf1X+FRrkFotSYZb8T3bbEWyWMT9zVb4r1pNyCn2zoj8/KO4PgYFci4n7AJlmn
RAB2CzyF6PkgTXFK3BKGDV3+wXoNvIXIrnT/HNUZ2SUCwvTMRaF5xGqyyFCGma34
CmPmcaR+RpvaNeJ2MYaKThHgovjw68bE5YphZAqwpIbk0o5haQCUl9twbgbPb9nC
AQgl7m0XEkXeJhWOi9wG6CcI4ZSCqdCdBtY6q6E70hD4y26qmuqutMIZI2fhGlod
uvhEIIgB33HOZB/wykwIPDdJnw055eoLVvjQ1R+TUdhJFSPGoFIkvh6TIPlZKc8D
b9OOiKpl6EV6lAjTadkd7yL66kR2vmZ4DW1hsy3YnweMyeSqvLorWQTWF+af7TNU
KKVKqxy6Tq5r75XastrmI9+k8fubSGXNhySk2hsafyUntYmi2MMN7lM3Xscqk2m/
j8XlReC+rfohjM8szJcTfzoemMJCZuiLb0ZW4K6LwAi7ObdwuBfIwW8W4lRGNF7z
jGZas1EzuqeAT3YtMhwThgsk3Z0sSM5p6UHw+ghT1Hd4X4s2UQV1+KgmdDNwMDu4
sTQSZtHDjPYCEOZXN2OAfPDlXeZKhY0qH3VKpjTqVpvnevs/IDL4+Z67vWkJyMIW
jgudo6eibsB99ZRAc+ReqUsozzp0uu+YFeEODBUYTLGOYuUFjRgtXbvVJ/cLhXF9
UkeefNfHj8vRu/njg5o7jOYRJhAID3Hcn+yFgn7hSM36M5OVRc8r9RAhm5DHUUDM
dxdIJHih4Tqx53dQXSYiymaT4Ft2rqCgRS9Ikp2vddsdzaM8Abvm6LaYstOdq1Kk
Gny+XGNetPlXccr0pCd5XVi1PFqK7BPnF7rUQEoGv5yj3M9zkjhUYL1+EB2QvFkJ
jJiy95+dmt1EdE4T2rHU/T3i5SGR2xKUaqjNOtcqDHvAUkZmnT2FItlWf1iOCF3U
y9IzrC9tQ8EvrfsFVVVFxVh2FAntDNdFEn9ZGwKM2p1iW4sJAwJTZF39a+zjDoQV
aMzCo5DQ1h0Hmv1eFyzY7Fd4n+v4NVwJzdCXvAErCJkaIcyKvCehBcPz+Zpm35VM
huUEBFggHkQAMXxtbVGFj7+xxL4hxgmqHDwLkqRg/6K6SHBc4s0sayYeKvzCt4w5
ODHAtz3hyYaqCb/8F6LK+VAy5m29u9qRs0bxRRvoxhgG3WjzdOKqHLIdbdP5jZXj
HkLXwDGlS0KPFhUcMaOUqYru78QezaazPhYICcah+Kv0VZbExAuGOY3N5g7NSSd9
Q++2fQgBZ7Z2QSxhaGMemRTxWf+fJI0UJ7+Jtp+70iDkd33bv0NaMbFOnZterWcC
Z0y7h0jWQy+M24TlSI0iHUeCxIGyTju0hdFmjTLmy4VkkybYDIgKiyi4pFC2hAkT
32gJFKMbmcqwiIL93uJR2d87CDFyfhOJMQRQLFG7OryY5phMuloxxzTHqRoSoxGH
NW6IeeLr4mRlATakyS7g50q7TP9RWUkxY4CGGJdSLCRgVQOduVI8g7saiM8S1vtV
81pXoHt8HQrYEnKrbVMZcvsC5P2wNYtgJeaTDTsQTAn6xJ4sXS9hEp4cs0/ibMQ4
CXvhxhh9Tk/A+5yiGzWa7Y1T1qnVntLS+wW6HlZ+bH8wwKPYRkjQ1KbU/gxu+0M1
i2Wn6AXbms09UECaHU4uGGOVyTX8FSizL0Ekz7v+l4Wp4CUl043WW2DjoDHGMJgU
sm3wVqJAubVwIZnc3Dkru71Cl8P6Xivdvr3tqaohWHrJT+zc2HGG7rrfbjNs6qPK
ACyeUc0kDiOLSVO0dl3TNWUBg0B0UyJbHjLXow5ZlaYKjdW0acIj1/eqIRCxUuHT
+rGNMbss6VUwN6Jym9UmPBTJmX4u2EOjdwpT/syk9bkeg+BXOhInRWRBg0tSARRd
kKN6cLIxsj/GERc1ftfqMwG5QUxZfxnyKpYQry+LCGJbJY9TF/UWe8Wc6Z9P3uPD
Bc2UhOFeDzA46pqwr7DLt/b2hhK1HWvvlvC966TkLoc8oQpulbptx4anYJ7PrsAL
jkvzIq2Q5XLsAM5Kdqg6W3qDPD/LnUphoXrwy9dy5EUvTsdGQ2AFn3NP5WgukYYO
BpQUV67lWrrqGU2VYOPj9uwf4SbDUkX9VsQ2DsByonovQB2DQakobfHf4M3NFIrq
udO6DfIykPW5DBeAbz3AxOAwtFyw6z1QuoIwc2/FEAqZvN2lk2BcRmaTC4USBsAa
BQceBmJK+my2/Fm+rHNY8s6gigKcKMukbJ5egeAftchBiw1+JABZHaHZ57lHQR8S
f33M2DjpWaugh2d3XcBiufZ7A4K/6CLv4A78VAVud2xMt+yuhBQEde1VLMP3KcEE
zfXxIAkdWubsQUUCFh/09DtEaekJoctRQYFLQYDpZvwlJF64mHYOTI6d8ffIIVKI
OFU/L2ekRgcJy4fk1r3k3BfVzmySCHTHcpOUBjXRBYbvR+6m4lXEcxHLIiJeFQm7
ta0WAWIIg/E9kaarGBLxl3781fWN6/oF1sWYr5AmU1lzC+ZTWHuRyoHw7DHMugL0
SmV79/YiovOOnDYDUbvWrUvTB+GZog0BrIDeL90QJ/x+CatcHbEQMDx5BqtnLEsA
FZWS2bj01Mx8TDk7A8fjwyKnRoTJVvPfK7G+KLZAaC4RQglOyWSP4jj55N38HBEP
SSD0NicJr0hNYAFuGSpptmbYehjwkloZQ9qF1IC6wezLj9j6r/I5LodGpQdzdd+p
AXUJkSatKIf46/0PR+TKR0DFfoc0v7hcaD6DIdgxyP//I1fKheefh/SNvqxTdxx0
qpW52CTS1O8YEURpMfzqzerxg8RfBp4UVoddDOgH3bfC31f46clemMB/SOCIqN0E
YWuGjFVvqHGCxlxGaf14i/GU1SNF0fimmoZuYhC0cNNKoZfRZB9rbcmMiGDxleIx
DwBQtoMvXI/hyTWjTHGdfmqA2qxLVgN7G+CMUN3CdnDl2X3PKgB1+HKQ7bWXYex0
FYDiT+dLm/rcN0t1/99WYIRDeIdP1C2Jq9lDcHJ6OslDxRZjezzi9NKg1vOSJekA
/cOghpBqIXcZEB/x1Jp26OJ+kQ9t2uMGQxltYj/3Iw9KX/A+hjKzWkNuGg5yRrQh
4z9bYViieH+pdaPlgk9bcfBuVtO4PQ3CS+eW1I6w46CHcnWxBKVdjbf2GH5BAmSp
gOEObJzZOxkImdL/IXuggI96wGQv9PrqhsEOG9+q4f3FBHA0eUN1eB3RZ1OIETKV
KZhadFviqOIGslFQFFGPyir2j46WngBpz5mGJSFOMCjnMF8ajD2+/6ZofunYpluu
gr3lo8/+xZS5O6qhsxpGRqtEpKHZi6JE9l2mMH+Wi0ljWzdhXKj0yt/wEDVwRaoO
J24E9L6e0Nv+3C50cwWIQdxy5p9fTlVtGgIyO5ui3w4eKFNl4ouv9KMYFDwmH6Fg
yKQZHiQCw08z+s9ciAfEV7Y8GkzmkCb951UHNyGj65bshMWjUFOwqu/+iUV5jIxk
6iDdLhiTTmWr9u4lnB5zkqzZ7HxexQUVZ91BUKkmXt77LwDu2asuRwzXOwL9ewuF
POhZZe7CK2uVfvq7EnvIxniGsTiyaETwzNUsG52oNWWmbUOYrdjpDvRL/zNgYlbM
SDLG7K7j2NSm9gZuHPoUwbmO41NznaPkepNzitVHYAuNJXF2PctNOiIqp/+o+i6o
oVcmupWY0S/edgO2ijFS/s6sol8KMobuK/4MA5stCAuZgBsz2DKrGA49uk/12hyj
v0y23Df9cDd1cejHXvdWCA1529HAnBHsEFKgevPRLhb2BjT81a3Il9FKpWW3bpc7
QkpxVseZRhPvYwDzP1G6S3AUBozwqOXjpoOiYZFlLrAlgRCMZPrsrP6HDy+uitpa
xbY7BfFhSBoQen2/C4CgoFibDTdSUijW3E1EfZx0VfhEpTve3IfNoURWpiqrErGc
9LTDUzOzQKJ+HEndIQTCKr7Tk1YbylA1Y58Fosz7Vh14RIy1CP6I45XXztCMkd6h
2dHsGVbWEf/a2F5isjHH+rSojDMytcWKKTDbmznL6ko95P4LQzgn0fbo74VSKIO2
3qH2u0gaoeIv60TgjaNVTKlsZbAwazFn/9TR7WlqD9Z6z/gI2i9CIB2DfEgb9Fuf
n12yiBPPu+eU8EVQ7GAGWJj00+1abXNpaAoXahMEf7C+MIRj84eC4a32hL957zw/
GdXEfhesCNoqDR/nt7R+lHyxsdUJePbAAzy8Lt9xkCKo7rk1HpXXVMzulZnIcZMC
l4717Y5UR0o2LANjmWW/bxxJd3Ah28i1RRgv4+c6H3ZYVQ6wPWOdWyKUaQz1qNyI
EknGcROpX72p/MZUl/OgYY6rS6GA/zlX24JuYtazWT9mHbqDTrec26fmP7EvinUL
La1WEmrOPuCBx5f4zm4KxgamSNrJRw27G8TEAf6oc7bUb/h6KDs2H6Lt1qF6lAl2
ZyYGbBTyX35n7b3M4TplYWCIlhVAWODgEFV7ynNwzATx24zlbZMxfQ8yECu7Da2B
9VY3ze2A5pisUVlednYwuiLBLSCm9Ev0zZ788NsXB6tO8nh8U6EaMR0PRpsbRgsz
d7KA5I5KLJ5PXRjFTl36/CYYEfU9FCuxwanFf7LPWUSg8TntVcgD+cIR9HSqHekE
/jXO5f3f0BoABviNxfM7wq64SkAVwGeVPHIiswsJL3GbNlNXgkh0b/jW/iRbBpFk
aehKDN/26ipiPJMXgsZFXO6ZwfwgrukmHIjHF9hlE12coeWI8/mE7uhie7oKOqVj
MSgjbI2bpb7HyExJ1CIeVH4eDrQ68mPo7Ga1zYgvM5Q/l6N7tDLo4W2MniYqoVdA
DKjfURGNAti1uWvqNMdCRZ9rnPo6MKrQNALC3lyno00yxVrXtiwsd7VqmANULvmL
Tcn4pFPL3Ls0EPaPoSPMebrTniWEBLXxKAyHeAzGcAUAnAj1rf+cSPljZ4u2VweX
5gwrxJvZZCFc7CKob8+CkyOqJStTpb1+qiB5LYRcWOu8Gd/oy6LDxAsEz3+m2rhO
FV5igETfJg5kb/4TaI0lqd+8lddLc4ju8XX6mMHwsbDwnr6o0k7/M8dQx6lWm6bF
FhjiBdqXEG5tvleMgoVBmIXHxVuzRVcuDxNmIsrR5HVufYY3mwubPMu9ALpndKsm
yo7FAfi3tAa7if6a4JTNWtqouNkOMdVbH5IFrRPt5Lclr0GiCU47KelVfXoIlzNJ
ZvbzafxppyOw0nMQCJsrXJ/zu+9k17gIdh+oKyU4wAFjBr3b1gE+RnSCxXxDPKYh
GpeBQIYGUp71ZpOpsaGjSBg01Xn8apwPOPScFBctKCusn50eOBfHRyPlmZ35CxUh
RYDPfH/RKhn9bPrg5g+W45enUr5nvGtNleGXlxeFh0NlT7kCY620ICfosF3YaqEC
4fbwtJ7efZ4+IRI7tYtRJ5R0SqZilCuyqhmDQ/v35SbhWdwapsvyKPFpgNgTn59S
uklzf2v1XH0QdUMV8lTKCxsWV6h/tgyqRJugqj5dp2xi4rr8TzmnT+eG+JTEKZBg
cMB/YTDKNkzJF2QElUDKaEqkXIGDZMS1GeD1m8I72L6xfJTPvwEIzYXcJ4LVz890
ANJbEb9DLtc5wKWiP4gEkj+oHYLBMdh8AclBinEqZRyzxKjhKuhj5RRCctucLzID
3IybLMZ85aCK4/ezKupYFfo5dnwI/RLi+t2M3gFsjtK7B7r16NygwcF/Nh3IMox1
ZXpYoEPbNPtqdXQNsjJiHRXScSloWOznQAIlQpbSn/WiFXoigdHrgMwiIOX9HsWt
Si/TOqXVHuF5Zl0vlmPFYqpXP3UfszBsxvRaEZ2lrkiTROEFvnlr6QlwDOCBkFNs
c37L5EQNsrFlXoqpaJpUbB2KpPInFHPxf/dlTZFH9f4/8Qcj5xL53FCfINtDVISo
xHfHX8yLLCnJOXcBhKChnC97FYWNP1Xww2tuD/X/KWdFKTlt4kCg+uI5xeKJajNC
rYpQUI8cqeQg/W0882dNYKxEf5QwgVWidO1EkZn8RfC4V7VCfyU7//GNertq96NF
6vbTiIDUVJ4EBQpFdawAXYiCMcbqchb1jSbHuRn52kX1g4Y2MpU+7XspM8IxdlYo
7YX+l14DkbT8mSmLKvm3Ona003YcWq8PX/C9ua1hx+ZIpyYgEhmfhvY+CPpPECpG
yjGG1PPnW4XT+7lPr6lP9fELqo0bwMWjRPMIaVxtpGvtO8VBy4RCAlkINCuDAPFp
5dPNAYJMH6k760iqgjPWLB7vhBbb0PTx2N7cCudm9LfROD82CWgvIByvnrxCdbeK
lyGKa/8fkcPobxgJQBb6n6h0ytIyjm1L9nuf9SaCmQWvubL5zzUSR79UnLiKbupZ
wFX9UhWIlNclDA2fYXDqhgkAZu7URqBC50lQLyoaNK3O94qIYWGrTl3UoO7GWTYQ
DiTZwIQwecanOZ/HAfpg4SUqocZtd7uLu49pyyBCPYVUyvZTUCIHfQd89pNSbvLf
/0e7ZXkZ8iRCVwIHEmx0XWe1a8FTiV75Ri286v9DVZtGXZ7jKsbKjCbz+AyOWeC4
4NMHWoZ2FjNbSlJPIHcvtRkBT2zSg6CTxb3PeUJ9evnttbRInAmmLZP2ktRdU9Og
3/SD7ol7BgBMO7YZ8VeM669IHJQ8uS77dUT+8o+0lpZHYCT3ARWmxZbNKMO5rWrQ
4eGFteCg8FBPISlpJ7Pga9PiEdG2ApEUHP+/84b/wWnZcIdOI6YkJy6UKZ4jB62x
YTS2/XP41MqfWzUP5sLReYh43UhgbqIZQeLQfyqrfE9RpoGHnmqU0NV75YqDa+hZ
AVxhKJUdiEyG6PFzNSzLzRNmwaDOwftSNVCGZYqtU3uKn/PdEn6OD22Z7E5ocpmy
t2aW3xv4KpHN809PCY1h/eUrJKsdO0t2LMBE7mol3x0hOQLaT6zcS9Xv7tRKWc4n
8+VkVApYKvQ2xtdfrTdXrlnDz4Zpyv8ynsxyjjozm6satLrFZajholZ7sYCynySZ
CpewdPMfd3oXW/6G9SNhVP0igsfXMFSYxJyX/Cn5t7wfPUTkxIZ2EEaLveJCErwv
ETOClH/0OiecL4Lbu0lqV4WOCCIa/oWTed5v8bjKezPT0xPtGrQENSqCE6IcP4rN
eLmwHDIsMc1+h4ATs1yjXxc/8JB3EmAa2CKiLoiyaU4SzdRP1KH32PMaz69KjgCl
9i7HIUexfU4//4u3V+e0V7Wqct+WCdFng7l2xdGOUZe5xw54Hxs6gN3c53GhgkHD
GPBf9+kWuz9JGh8ahhWhwX0DC71hSsbiY2I2WLPUyUdtxMEPQcVeABiRNpedWlJf
CNhM7RjqtIt+uOQ19Vn8n6GaaLLg6f+xr/0qbUmDZsnxnA01FqDrm6/4kP/K+CN/
s2m7j5xbxdCH4gXwQPvPFJqZXKKnZhrL1nKfDg0qLobUc0gxUFz7cEXFzWQgZsVO
WfoXZh6c7tnrw/y1Ke1TNJjgwkufP7zGKEFV/vUaz2s+wXs7ta8c1sznPEp8VIqx
7OobyrtUSW9ofA47Su8JZN9dms7g5e90ofX+i+hPK6k7FKcoZ5qih3AnO7AOvChe
k+kEr61vgqQxSMkVC+EB9ViZEFAcnO5l8XUn2gC3F8qP2Fmbhh7g64peELmFU2NM
OgYn5iQQw/huaeNCJqgd+zwDSkZRMxyHEB5kb39cqCijTRXNG5fgHqoGp6eJrJZT
nC4vAvT/4G8e8k6PmbSqlKfaNmlwlTIjhy5Phy1XozWWGrJe0blIk5d0QnM7TJj+
Stg6aDlCB49OR3CRTuhVhfqOQDYY/PXAHuYzGDKKy/RUYR0Ad7y8gCGvu1u3YTxD
bmAK2lDri6FPlM8YYs4MkZbyGHoDH490DuIjjuXZ9nCYeryed+OKNxwY9q0doU0k
+orktSo/0T8BDKqiIoMhxak1W6LEZobsI4vT4459TEJ9FAL/oJ4wwvqlfMWoq+7i
VpOhIe58GKvNsu+I3X5/4eBUALCIXCgDINaqokn3OGOMclQaOHV3ruW9KEqR93hw
dKPDpIoydzvWeM/CYx7NYCmENNe5ttyNzhbQx7U0twn6Z0qGAe+Bb9RtRFGXXwsF
DyWmtR88uoOsyzy+HAu9bsWzGt9d7Hl2d0+NJvDyPA+ZMnp1F6Y7dOYtZiod9KjY
v8fixqFcv4Ehmr+EK5Mmj14Vz8aZPe3vsVx8H8mYyqHUFJFVr2DBt0koLw8Nyz4T
orQgz9Imc5do+Qzd/XLwA5yb9jXXC0NaThh9gPNXSrsxbWAPovw9ZoW9ZOD+fw+l
6Jql8sPh1cBhXJGI0Jl8NXsPjWlKbK3M+IKY7rLfrunyegezK0umJbZEBFvzPYUo
t9mPEYr8vT7V4I0nwJbj1bQCB14mIcdQ6so14/DR/MZlWFrX7zsPDTV09KLIObod
Epz4n93yf2bJ89bvgCd1WssnZqKqDVThI1wWHocZKbd5AdXBOvNWa354I3y81lUB
Uq1hmjWqsS7b9eT/HZA5Zn2EWcONSQFq6L8j5Aj0c2zAlFIldKxzQcQw/+eRe+6z
tDZexwYKWpjARhW3NvQGWf9/GkrtYKpzNycdj0Zvf37gbK3nhtUXDVgHb6xzySvN
X8wrLOyzPA/nGwfPh9ayUeqcB6ltp6IPG48rKapxXMJgVbJSPXywNIexsZLfz+7x
Ee9M7ahhW4tj9dKS2dTLm23N4aHGuC4YjGsqMJ6dPA3gHOOHlHicW2BZE6YP1rlF
WZYmLBzSeikHk+Qvce1r+0RxhkzfkZMJKadC/GJPL+osbbuPY449TO8eePs+8xNb
Dcxq+RuFozoLeOYzrXOp/7836DkI3Dj+c89jTdixDsQCXEM8JsbwQih6qF6bu9nb
MYeILQDxxAEGMarq/9YOV4NHCekgLmkScwNliq85ERMQ8N9W5GipVQNi/9im44Gv
+shP9DW7AcBb/9tk1M3dR9gZINb81TWRqmcjdgvqbV4MaBFVbrzDRy/Ie3lxE6mg
LyI9OFvJIPQYlr5AOsr1QToHV3qmWQJM0czuPLHXKdkcqpRo4mhdN9MF88FM5UYg
RuX0zNA4iIe2q7hOWGcZ3QpDlWASNiLI6lj4uy9A4MkOCpOekGrr4WLShIHLzzHy
8hqyh2B3Slp9xtxm4ZLP0NIeMAiT171zMxIjBw/lvZj/gQ3UlMEZLyNtPATmgvn3
ygj95I642AabbecLXw+ewwt7X3ioVGlycyytxdN2ThMMJzfGpvRnPY3blNWrje0s
MHcrvm7CKUss8AMdwXtsIHGAhGJC47yGh9fZpe6E+AfbXXBPANjSSluf99s1sfwX
BqrrP3CfTDq857G6zL+gD4efc2Z+1fwFytXh8sR+39ketW49v6vmOY0rV0COqtNm
jOGyNWPrIMY+bHmCKDDKzgPJMQ6USLJ6D9FruAfzW6YBRFkhHs9+Hy2d6sg0Jg4x
+eR0yuRTwNbfP5W/C1bOucKGjmSC1l951BnAwq2MROpo3hXXq4ph9oRcF8xAWacW
b50QnUMrPemKOUdrKk6kOhnj786FIXrabUGvIKDBQEo3hewzdvHgy9HZXzmWgNNk
2rMZ7GIMPyv3C5UL+Xw4UfAefbmtMZ66SX8uwzNTSkEUNtxsVhJtOAvJoBXahRfO
8g7jLinhALsd4+CwiieEnsNnHb8hz3oQ3+97ppvc3MGf18gefxBpRKwfj90QaX9T
4oStFSseI2oUsX3lYNXr+huhVlNJegAB2X2+1oG7B6RWJ6zY0P97Fth1LTxD1vY+
kA0G68zav0Wlvl5td2TquDOx+Rp9kyLRzfFdz/lYmW+ipBGw+kRgZul+ElERCfgr
bGEXVOAHeFpYRJqO2W+9XmFU38Ho3DmqZ4jJK7ETYrO49CngbcPHgxUUEMoIr+5Z
iov6BNnXPZVy+TwVFhKIFzYNCetmX8UefMNNAunZmWmq6Ww8y+F70l/fPgLRJqJH
FAocstRz7oW0G7tTAifXVwUH0RkP+uXYMgEuYIn/3eLFLy5Siq59eJnRmOfY+VPl
YcZQM9JVPM0FOGjiOQVedWDK1taIO98DLvr2fhrMR2T44F+Wp8OLar0KHc0AcnEv
nkUhWCVyTKZoI3IkKrvJ5uOpi93q/mdNJUUZKSa0wdqXg/l+xIECDr0w0AFgRB9L
nGS8NyPkjwnHJwpNeJGpnamtV1pq3YaWTgo0w2DWVtdE5nWEpHIN+hUAksqyezRn
LYv7g1Q1jSLzLh9V6a0dL5nVtnZNbhZcEEqiMUEDCQplCPB3gCG/D1Fb1F3RTYQ/
xR7kvVHWW4JshSNrvPIj3y7zLvGbsg6JLZkoZeAB6lfEnjcnj2JcGRp1fmJZ47H9
PkXvStUKIasPDsseuF8Y96CAkHCyr0GRSJPUF1nKD9M9g0cOhsuoawsuJZDM3FV2
OUps9W5owFtbxOME/Scqdpxp7nSoUOSGCUE6EkeanJhWaybux0ga32M/t6f0M4GN
YsoCSWO9Hy8dloUBGBkjkFyryhos5MAZ9zs3v/1Zxez3JEV1Ovw7s/grJRITFGcw
GW/JXfjLfbLdIQDuvBcRycfkTw+a5QC3HzPXIEmKNT3lWW7Dc2TjoRuai5o457/C
H6DfST5yih7WVGsZqMTnNN5uWTEds1vUAdsLrW2N6Dmt6PyUrXtDFFwz3Hx3FoOZ
aQ6GfvQQ2jgBlDqq856jmW1x2xpaRuJjEsXHXN0sWqj//7KMZeck8Sl7K8DRkDKk
6DwHjODy2BN1ZW2g1e29A8qyARlgohg8pD0uA1IDujGlOJoHySzWD+J8Opu3otCi
40K61tauBmdrMKwWlpsuFgYMran6cYCkeLNwtCFaBnGwYRod2m+4ReVH1AyJciM+
P/0qt7PHZwPCoVtByiX3QEgIoAPAeuaBqdvHhHx+qlwDiqf1ldmbS0L4QGKfIdpG
DoUHtLO840LK5PGyKsdB/SJV53KQtKlTtGBrKzkd/lDtiC5f+LhqPxpiC4it7s7o
/rLKoeT82sFHAORjTX/n3QwVaBgW5tVpUk+b2wk1w8lIO2OcKpGJix1QqTmVE0uO
KYL4pLLA0g/Q5Z9nzz8OvdE6IXQdsZC1gM5y/rTGq7sbPWtDJXvc/fc1tX6HUjXM
UDGTV0gHQ/s+95HU45L/BLuG/yqR21bP9k6CUNh7kr5OLIRlQBctXN0uRrHwGCv3
v1xfOrrIqnRbGDyUqyY005MUcHsy69O0eJgIAxwqdkEKHlJv2t9tbaeWX/WUjn3R
6Kyg92+f9H/hOLcfi+A0BxUP2Xf4c1oxJPP81cbpCkFxIv4qAtsq+1LQ7cZoHyFM
mfaacBTuZhMCdsjsesjPfhNiI3AQ9ou3rVQUqlYWy2tT06o0Bbn0VVFlCxvdII0T
csRECDw7pEI3TdfUlybh+MNRctpFaocxWnea/31GIIKL13YWqCAMzpA5dEuh0zag
AojocHc1nbVPAGoS6QStk1mj8wKZ5gNbnxmz9vQ+ZSSyKINlc1NxEYjnM5cgD4sQ
7xx4Y+L+i5bxsdxMTnQaw0mYFC+q9pkwI6pIkQDJrFUfTkVgLTaqX+wnVFKpZoRp
YW085wYcftkR8r4PcM0QROUVCu4dTkUIomBw2a2ZDRKvx35BXv0QTZzErASc4hii
/w0OUZe/uwtvoRrBtTQtGr2NwaYqIoF8bUqwz36NT0yzpD5zES1v2ygL6sBI0LMA
4Ms88ZsqRb48xf64eia9gjR7DxVvnA3oXaWPQ1ukFq0GD4cqHQFo/QJL8YEKWaz0
pnNBbFSM+JpmOdYp1nM26tBuDf/KSI83CbwbSfLNOIpaDNdWLjKUhhvJOBSi+U/i
9b+vGb0yASNh+9KFXJama0EjjfqXi3XvynjxX1ZOxSNWPwgL2FDEaA8QKxnc1wOf
FKR3Xg1hdVkwCyhREV/+MSc3RLxqvsS2QlPltUDr/joPu/SFr1WylhLYXQeDdLDs
7vPjwA5YmJWYhoaSKrocJGKNHQNHsUjkuR6JxVf3wVVAWJJ1Gi7R3s4I9tQN1z8v
y9d+swnAHtOEKH9B+7wAAFomiGtND4hbEgPr8EEsv2xdRyqRoQNGZUWjiPgTC21F
aEZHVnkxsKd3q9ZyDXqd12HiqEKMznyrtBjj7TWgz4pYFoVGTm1CA0q31fB8QMX0
oODMxRoZLsP9zXnMGSdFqYGn4qoX5XqqdAEB8f2CT9JA30BeKuiwqMhPreHHzlCA
OLd2kebDDagivAj8JNj7mgzfWr8cmRO69UU/Oi68qcqZ0msT/dYX1szHwEKZxCEd
YGTk1/E9RuPsEV9d03qvnbBqkNT+Ld65JNPfAXk/s8El7SEfAmuDWhPYueJVyoMN
7lO6SMBtFpcxOdJInUdu96Kyf1DXOpPzeXLvq1KJDFo+mEL1L1N7Yj3nV7lrSCdk
CN/omJ3Q4jNLlMm9EdyR3KAql1NZLqw9O6+00eJGG/g+yORZtrgLBGJ7obWqkAdb
3eRrT+MtFDIVy2SfH35yCRAVd5Vj3cZIJ/eaIO7MFKjWYdnEAjmusEsCKFbI6rFz
BKlKvj0djTB8LM4XiV/jdHLgqbgFoVV6kMpsX3a8i4uRMvIXPzx7MeK1ZA7rQn3L
OpjFotIYHHL2wBeCAgMZsQICMiukVW3d59yUy0Q/ycNeeCYhoe/Qv13xRSg9U/E2
8wGaUlQ4I1P/WLaMDeUNwjPkKSeTQhUBDg+/N/2zCdUC8AeC3mUbvmExhreMUwb7
9zB/smIec+MRpvv2Qbd/7H8CG8qv1NBUE7EHCzXiwsQFoQP0xSLzfe3IfcNjbibM
I2vGjzFLrJpFnXdn5kFh4hvh3Am5R6iMDfC9KPsHfSEg0rtxIr880uhZ2etys97l
+vkPiOaikkoQ4luZ+QqV0952H6hJzm9JtMoV+u5COX5c/DrqAJsXVePmXUKOSeuB
Lo8VvGWgrkhsl/yPagJK+KOTxBjjE4XgcrU/cbMcGBkqA5NgnspGQrhILMF7SCZV
cGnpdt+AOmgxOoZlie67giIVKjnth/deLE7oSq6Q0+e/pj5LWT+1us+nl/FgpLxZ
Vq3uK+Z+bWFItYDKNlI4plDV7YzPLe3SMP5OaGrfQCbmevKs87JkDvaTuKO4Ul4Z
iJs9ujjyVfPx4YmVXQlnnlofjJDjzIKhYiCd+BjH+QRb3BSlY3Z77D3x7mLI6FZF
SyBP7hJuAs9oVh8Jobyok9SOrRkOJe7qnLH5ytNRZpQd/Q2wvT3qIWnLlk//iw7J
+qk/Vl7Y/PDOXZKYEJEKOdhJBozzYGAuFWtQUISkGXAMcsLAyPL5jN5BAlDhaelL
zMCReWpWhr3GUKwn2Ax4g2AbAFtsUI5+0dXOzwvVd+3j3eFPXJO9H8A4/Fqojqaq
x82x0kBhLiBbTwGYSFdoTJprP0eqn7I5l6/VH+5CGT9vUdIxehxV8Z55RS+AG+nP
HE1HU7ZIIJM8wGdobq/5cTQ3XBqx4YKlxemTchNmDmqkBwtk14JWo0v7aGfHOH0N
S/5uToHSJ+LicJSdIPJklblbXXJBoXyMwEQi2+5HtWY3zPQNyQ2+Hlk4X8+o+w3Y
K+BtZP6OpjsdfCJ/ecIJ+KdmViZgZi3Wnr6bBzkiqzA3X+VNM98lr4+0MFmQOPW8
Ou1N2BXaJnUpA/nPqwNFhMPLb3oj0AJhucP+2UEkKhVsgrklsu5+68culD0GBFGH
Fs1Zu5LwWGDYSNxQ0uAwzfdF/aPitasmVcLxPq1B0PLamMLq8X3b1OJsGF4CUqPE
bUJxim3yX+5zXikYaEjhWVaY+CgGqaZSndCpgYy4HTUBiaWZfECGYZQa9hgogoiR
sdq0nKg1pA2KsQMkTJKQZRSmmHMBO8Ys5vHedzYj51F9tl/j/dtJ17yjXgtjQVdq
Jd+slzBuHoLoBqZc5LEia98H7b7fUdjMo2kx+6sRQ3kqlyEWCZIPaQXMncPdIY9M
SwTJ9MjsZwYWGJNYjb1imZqnrVVKEASelQb/50/PF3FSgWtcFAHsODBogZA7Fpnl
tp6TaxqKxK0xbbnC/OyUIoYcEBTqSgXV0TAlYEVGQ8zqmDdPfk9HYM/6ClgTPu97
uDHdBgc2FR56O6N3QfOE9h9bqcxEkN675eX3oDpQYT8iAWiEeIH3uGgFZ1OfPq4j
8I5x86/v8PT2M061gaDjY8mK0X+kgRp6Nl2yL14p7s35fa/jeNCryCYk1Kjv9uPm
wThsJ4p4T7c9j4nYOBSS74PFxtSrDpaMVIXcn9LQeMyL82H04PCiQuqYoNPIcnBc
znyDcha/sVy4LFEiSYgqzyMMdOJIRFS+F0Y/NnJAvttJjNV0X2cwqYPzC9UDJBPl
LNnwTpL7THh892rlpAivydGHbeOhTMFAJ+br8JhSYoGqFExzKO5ZXSxBWoxgKAML
BsWHD61R9nfBBxA6v9y/ZWnaDbhXjnO1pI9wvS3WPKciWFR8iljvR1ZQWXgt7vRD
SFCP7sdtGQyirtXncG+GI7D6ePDqFN7RLGNIYmxwvAAgzEQVh25YJZQ4qV4L5Ql6
VzisN2ussFMM4eU/er9FOB587SK/n3mUgpNCI6pzhcTqrCoCl8iduU+8ANUIgR9s
SPHQupa5rVWNcez5QJvt0YItMmo9iCVAHtk8tunVG5LZ8ZN/HeJXFqClC7KN5uW4
XLfZT3/QnDmmAg0h0eKaWuoCgyCf4EagGdNu6Rnr5qh3ruUvxSrm+OqG01+7uhEz
KpJy3xYmryZxE9T/r/nTe4kmYYonuz9SILegfTRqdgAV9W01uOppzXRylN+dQjMv
yq866/uTEjDORYQpsHhcQKKWvtHkzPqtqt66kB66wKHiLgpN1elnu53Y6Qo8LC0Y
/nptdz0En9MqUTiZoos8AENvtPBsRIHhUFOk+7DHX9XrqpiM5eDM540pYhKw+Jar
xt9KU02Pdq19aL+U4t3AwNHevkbVXGAPzODMB69ITgNGX66rsOdNk8+t+vSLlGb7
LKwvHQ+jwYPe59wRfoepUSOfngILBnyYt+EFLY21ULydHI0IbNOA16YM5/xk+DFl
e1uxk3Li6Jccx2pLXhSozVxPDCdOaNB4CF1df9f/BVL1+Oj8lRWrCnz8SHPrHm0I
qHT5cxRp7StkPONzi83whZ9qbqr6bi1LYSzkdjq2rvnd0mBdB/qJA2Au0FNbf+ug
kIMeSoa/e/d4vP4EfykPDxqcsZ6MdJI4JIHDOQhfkTfblkoCeBJQJrG5Csqm0Y2B
k6RK9g5So3VBPGpmPffXG6fr6FoaqOBhRhTBOWXLaBbDIOUr3y9InuZOTT7wfs9K
kWq3GTxBM2oK98/biNlPPItoeVTMOMraSKmwjG/ciAlJVBKFE4w+R26yRaP3iWUv
0w9TuCDtvphZy1J+MCj3EranakV3cKgE7+SNHu+RaX2NZRCvD8jtMIDPv7jt6p/c
N2oa1dbQIUHfZPTHmCs3qAbqZ+Uts2X2ZoPDtCItsgyH42ZPi0FKSGErG9rkL+MZ
WMb5zepNrqd7+vptabeTndQLpf4A+Qsgty58C4Zzbfj9hKO05E0dV+zB/m1/xJ+P
RTstIBeygpCEiclT65PjYOH9dCWQnh1mLRvZhOu18mpBoyHr693jzYZlUWB8Q95H
GzP6PhzrrajjhN+0WOxJSgMTANIfsQ42LG1caCX62dH2K0bH64n1Y2/nPeg6V0dW
C7tNeheimJeK/bWM3yV1E2CDhaCF2+/VJkvRpn9Nth7aVVdXPhd7XquE7v2rwAhA
YNGwaNVqTy5rKvt7uZONMKzoU4ZvusFuGsMrXcRBjMjA5iy3cX2R0X+FTMpeDplS
bEilmaAReNhOt0BBOno2VGrW0Y/dyfwzrdyqqrTva+3g+xKN3RJBJiyf3iRK31FA
u77hfa9BvkVsKrnpkSGc5gohplqMZEqvH1ai27NyH47i2K+ifVsjWCqy7eRN/0p/
jbvcrQGVdlzODa8PKBTHHegn+RbZ2fkgDYanXmuCihMq3FyLr4r/VWIWM0frsUC+
P1yCz2UmSElrQ9ayyJmicOXUvCJ2cKeTsFBx0EHRuCrNFw1wutVKv+ab8AwpeWFe
vCTvnFz2dj5MFilmzaa8usmwiztje4SLtoD+YwzgE9KFum1Cg6KhkCCzp3j4dx5v
RtG5AYleFkE0b717i3GaamMPcdVrRMFDzUvp87Ts5jYQhfd0pa1yOplj6EAeenrb
pr2tTCibyLohAX9CO1LcyUW31o+ptlhHGN8gr+mJQsYeew2kJpMccAIpnf35oEb1
nk4PN7vLnQCTfS9sYj6B8kl4MO72awLJhTqLQOqA9QrUvzL5B04ngo5Qz0lsF+7z
Y2NtR6kXXRxayTSKZc9wkiGyfPUQ3h02b2oQlCMlHV+IDGwF3rnfp+3ntk3f7d66
7tmDz6r7WwJKA7/9aNw4DMENbeN4Q8lSTb8avae6HRbzBfCchGC5HqcFEN023KFf
vxpQ6UjCMi/TL9gzAKvRMwPTkKek/ohCeJ2UewBjzex8TAAEV0hkcBqCL4Chj4G8
ErfNnymTwrxdbrfo4qCDd/IMzz8W6T4Nb10nnofJrLdhltH2ytyYUTNkOyFcDa2x
cgyOgE0HXnkfqHzWyqERVgIGnvDyuvv7Eh3D9tUu/ST3B+UUH84hc9XQrIsKzIAR
qOoVcKTLTD3NakYRMo7507QkmeYoCybAqHk7Ajy4X52I8+iojC85d4gsw2V+NDQw
EKgbNHtJUpubRxCd3GZA+uzFBLYlmfrZ3gYKEiZYs7B3jscRJJARrEKGezMYzgbY
X8f+3t7h4+SbuMPnnMaa9IA2VmsRvr1Deo3mRcfCmqTUWXFWH6rsHQfhYqHHTKhB
8lH5WM84n4s8Dyc1GujWzbix5/z14Sy/r+GBb2/E7fI9J1QGW4fAR3sLu6UYdn0U
HtnYncHd+9zPm6IdFwuz6HlUMEpy4RYOZyfRIET2iVrgeh4HckqXDAuidsWTkcI2
xeiLfQDEFUlKjOyZfuvZCaex5EQ0/0Tl/OEx4nftehB4ZtpKFk/MEH9bAf2ESV1q
cxvDoddSRctROz78VxxrLlcVRTejvdw0wAUz7/oNrGxNc2W1smZd2YqQvF2ghJsr
scIGYZp26Bv8eMGRlBT65n9U1PBkr1jq5VTZg74Ho77z5F5GPwFLmasEkvfb4Ei6
Js956WJlailEnXEzQKGMB4W5wNmM0QLRSelWBPXQynr+saMxXoJaJMQ0Y8SWWIN8
vAlXWwysNT2b1c+biu7isMDL/HohmDMolTvM3ruRkWIggS7buromzn/sJGkJYj9i
CqtjUhtevWXWYz6qaNUVwiCozceNQEBnhENeyL3Wpt0TgSVQA8JNU0C598gKcQZj
rmC4/u4Wx+q/DF3wAR/6BAHVcb7lEu2OoAJB5Xpxd77D74UPD/SbvbxlcF5FiWzy
aAeHaTWpZ8SZ/kz5qTSPgIIisd8o3US2g1uxc6c3PhSBS+oiDapiC1NvifJl0j44
hFyC47ScTrlG5oMfhTifJ+pyo71hMcV4A4ly40jJq1YQWXY58QQfE4T2LA1l2gvN
ESQ5rWJwF20MMLawWFUPWaPgTTCYT+bhvfgk/Vt0m2hArrwCrcn+FHZ5RfOodIwS
XoXJknZTL4oIGjgu0qxrV8+vwDdiCRg5rjXnS4+Zd60KkN6v3MYt5nyqHK3lrFsl
Ctw/VbEtNI6EeUVH6EohKLudZZyLobx1uxmPepY4e7pis6fU7KhIiPzKm9MXM8bk
XEkNp7WrIRJe7pgdJozq4jKAozk9qkqGBWxNhlmjQ7SJ4iySa6FoyMedDPIUMZ2Q
p5vhLiTz7TmBS1J5j+/EPSMKcjivIvPxT2XodoFB2HShY7okZaZpdYitI1DunYYM
gtC3vQiHHrzr5qjnLdVcaVPrB16CWoA94Z3CITDUbLi9Rb5bELMDnYEoXpbL1n2K
MZcTYT9h47e8YlrNNInSDaKJd7xeEA06M7atZJiPEGlDwEAmrHUmaeQ6ysLab4hP
wMfxTvPTrz52mDrcxA6ylif66G1LQ1ssoBH2Xb/PZYp2o5kkj9mVB7RRVvlAZ3cW
FypKsgkW6dAuO4VBz8WZvyxJm9Gqs4cPX0MQ1qn7EUtFToFAitr3ygvnK7qvQEdC
ZSXADZYEV6HDaNrfzBZT++sM6fdOz99Ujca4guuwXBo5rxbjsD+Uv0MKPKmnpA5q
q5uYwTgeFw0cV6I4m6afvKHFa2MmufZBCC1jMSq3Btnlj2DsKTDzeUzs5IpkUW47
Rp9o9uW5Tct7QRU69lQmyHpZJFdyYcuANnh761aRk79z7AnBQeFRzulu1gVwuybi
VQyLnJn2s13FVhGxbGEZPczFMcpWHlCloMq2INqLOoZ+b2VtFdWM5Xd0I1IPXDPH
UM+nUXQ96/MUNdfiKS2/aKm2+yaFGhWy8junf75uMPbKGQ4ANGew4YrLul+8HWiO
OnImGm16KeX4Hb8N9LilyxDoomkif5fgh/RVD44X08XVTOVgH8r03JPumiF7C5DE
rAz4kN/HqepT2rXn03kXW9GekJ0YDUea/1Zh7F5cSZM6Gxu0iljAcHPu+BIqVpX8
blKg2spmmgkg3zr6buKtxoJw0OwKwNpJoRWGS8GTzQRPk6qvaFqt2wmd03SNYVFm
zOhvpxb2Isb1VC5WzOEJ1lz3htPEhKgSyHf9xQQk1OJ817VgCbd8heoNoCmEbu46
XV+zGi3EM/SZqgDpbWZjgYakv/NW91OuZJu7mc4yFML01v/CknuQ6gJCm4seUJDx
iLGhhLdyRIszNTz77qhQMXh4LcGdnAlalhEBr9POVbJ0Q3LvlWxatn0/2iDaom9C
ZlwV+KglAymKV/vObGkuHWb3/SjeboOUWYUNZM+yDAeitvJQxv+GiuJzAK6S9fxg
UyBApTThX+ObW794NKRoe44ZAaWSDNNjVSki3G1rlWJnnPp8vV4IcTKFd07lVId8
NxpOk1Hb8d/QEHUeqBBA4WuRRqnt8yRDoQrON2LhTWuybdOlfoRAW0KmMeQJhOe5
OxHjz27RWD+a9tvyvc1KqUXXBwBfZX2gE9sk9RoHNwO0oi5B9FP4b0vrWPbcwAFx
UTEkeitHlaDwnbP15cK9gPnvDRAJCSOWtTVhRn7Npy8P7d/V1xgyMv8sbBl/t2WW
QH5KwW65m0SzJMJhEDpJ7x5vlH19Ar+ECxtNxPxjuvgwwRs/L99cA4S2AaxtmY5z
9OsPHiarkLdJZnFh2NqRLRBTgut/h1iJB5jExqHT3bNmR/lZllM0LvTi2rHTPhmL
h2ifLPkI5n7y/cf/F4kFZJ78ARe3L943khVZusJqYuoQMpi08Km3O3upHevUgTbO
zc3OAgZpTB9MWcoFjc2Loxb14jKyQQu5Av8xH4eTqtzEX0F3m+4lGl4A1s1kWper
aP3lj4yO4QchY7dTfB79UWt0UfIQGQ8d52xyLDJiyP+6dNgj4+kfsbXEwaiESHKg
9GYoaQqzS285s0Ar81NfWtoZj6TlwKEHD5grcWEtRM8otDnQ5FA4NS7FbM8pIWUW
keeuVXIY8HwDovug2FM1MNdjFDq721Aou5FsA6uYmnUMCH/utF7s/fmRYskXz6DD
/DTTYBgZwnXjb9+WEVUHPA1Pyi2sSv03FyrlJ5J/nG/5sKZlg1nRjU6z9rNn27tn
5Ra3y/fEOdK1b78alqe+/ak+Nq4x/COKY2C8BJbQ76FDH+u3yGEM+VM4Nb1SahNh
0MD753Z+DXfzphYQHqx4H5jmiPUG2ozl28nnnJngJgqfThcbMedVfXdj4f55PYTy
+m1wgek0qDG+/26Kzm02s1MlcGmN/9PIyRMuMaNZJT5KWlgIjFfOeheQfI5ZNw0S
C07lu8METqGNijjwoFXfXi8g76muToXDFbSSiszXGpbmhzLaQOBTHhqSxUiQ4lMw
85/21+tna3kmEkdZXah/Vrm8GdS0OGsbYqmGU0CdvIBncs2v1mUe6wWNOVysjt9H
lBnYVvfeq6pCPMz0PJQ956bBPfV8ZJy/40e/C0ObWmoE9YqHgA2u2qO3ElzDMBY8
LDY/xJxiXWkIdIg3I2iC/w5Ftm2GVmWIDAvymqxYU35RvOXZVuFaTusoxatvAW+n
bhIE87fcHh8P/rXxCNKyKXyDn1WmQ8iuo1hAr752cRI+In1iK3SExJyOOjvO2F9+
v2ubSf9j4jB/PASRllMl9vc8lN/dJx+uvLim5eKqzM8Sc2p6L6P76RZYTg6pBJ/K
/9TWTIwHZeOTrsScAoG9/kZxbGrNbBIzMa2xi1oRGkAhWyrUEPqFBD2eZ0QPTQ3l
I+oPkoT6uWeQtXkAoBTp8EE2moNFhIobGDcqYhnSRCNAmulbnoMguckUgyjgvOaS
mbvaAmAnNIi0Bu1OEPYsqLu1VYFX6rEKjjO4gu0QbFVDtRUMLhyNaGx5DjnsXBIE
MM/8350NAf6RgOo8Bs0WB0K4/purn71GA8B8WbtIIPyfw8P5n3Lnt9p4lqaJjsWu
jds81JnT9T5y44HR425IHQNh3u2RQaCqSIRbiksFm8Kg+NABCXzc31YVmJ39o2Ic
jJ7N7aUB6KNfD5AW0FFqiCIBzI1dZJB50JKZq+lyYh1sDcnv1mVMsqp7qaqnSkuK
wnqy7QsgSC7lU1oHQpnvhwdmBEJcW4XpdfHVMtgUwQjAPMyEanOXw+ku04wTFTvd
W29oDxyxEtNkqXpN74/rF7f6kUQns9AVJF51yocAeUONJfoz+c9hxVtDp1IrPm45
RIyrjvJZu352379aYqulKltIyxEh703GXO9M9idVDfA/O8zqIHyssokWy5AttisX
0ZbGGDJCe3NOvc9P3N4qLGj04hljg4Yy3bibODpXmHKcpa9pZf3HXA2mgi/RgKDG
kV2VkGJDAFlA8kzP9jXA/fnm5ykbQjBXgBy8cCZWh7jv6BaZKujmoQNn1E8jBQoa
R4gyHt+NfMIC2MPa4p2gDsZwJc5kMEKtm88QBo/CmDC55V7D4UEakkBWSwWENAae
3qm6QUTMu31yrKgD0TQwV2f2jdEOZBaPWbGfnUeoUlV9kaz0bj4psiCvf/cBb5ul
Z/Agqs8TbR6B7h4yToMQPaa2gVEVUbh0SoBjR1LvUGDseNYhp3ZcZ6kfDQQtxvhv
T7EyooH6/fq0llnn0DwO4O7PuI836MNOL0/X0Z4l1R6Ug30tme3s8WYB6pz8wsVO
7KmUXHOddeqfVh26TLOeVV/HVrg3WcTZuiksBeHGbjp6T5XnHx6sNmY+K738d0X7
g5+4m16V8ReffOBNWIrMtogTT5Jc+CPay7NZnDnTn7TaXoPuOPZGhPqA9W6LAP7r
3kxX/Aj6I2Pg7/2SZ3fsRcBoBrNxNO+4yliu6mQpq3SiQLflCxEGH0EpkFvMkpm5
sfcW6v+M8U0s2PfT0tTj+qxTfWo5syzZjgUktDPEmnlOJdVzuXixwEEUZ+FvqLZ6
MZd+uyd0QDmKkFABMBDgsaQyhMnzec5i597gkmA5lFJUyT7zzCw16BJcrMCC22RH
wi3IGJuhORsAwpSiblMRxG/hxMGucjOgQ9ket9Obs+EIUK4NP5zLX8F4sFyzr1Yh
s8CW9Ovr+MiRD3JeQljtmp13FIa/po+idOGMU2mgB2frpudgaygln3GOdbkKUlSC
vkqUK+LGRzSEtxd+MxJglJ7ZCURbnfaNsZXf2YB6CMOu7naa/JBt0QyUOxWIvwmv
7sGQ42gAidpcRMxo+x2/JhjIWj/iTilh5+450vI3R59W4tYFsuFuHSpJuqMgtbdY
48IlWAeXKJwgH1HU7cSB9fy5gVmsJis7C15x3hb0mrOXQ0SxFW6hpsI0xS5qRGiN
sGGGmNCyFiUswNOzyB4Bt5aarATJvvDEaGpbTjCw9emAPq6SK2L2BOQwA6y0EVs3
BA1C42QOcgCBhUQxevP47Rm66oxBvtTrBty4RE6rJ19V6VpCH7txlP7l1U9nz8nt
XV0MIfg4RpJ1aUYU1bqZMSwHSmExyII3s7UWu4sRia8c0dMKtMbgw1GyY0yO5otW
HZVlHiRuRsdvyFp25ByYE0jf3qVFP1ez+ApkDuru94+/H6mpaUWQtDSAnJ3VbNTv
OAKpVq+zYe+ocCIetGVJy+KsxMjtDAsmdakcM0tyhijP3TjXNEovLUKMGzakSpUb
8nvrJuiOOzqnzJoufTEqcSlUCsl+Lg/NH9WyhE2X5joKdygRo1XgV/YoH2JyMpu1
WOoQRSCGRADf4Srpc/6Jin35g+NBPoazQrBr2J9aROfEoSPrNmgeESiW44Ek+iLv
6yhmpPGyp2Iy94IAPMgN1cgxVLkXIM1GNn4IDbJkwrXeHtf14jt+0rVJTu9OJP9G
t8jd6v0Pm0S5MCGOKy8Oh47MGsLOT5PI0k9cDtVAJNHHRrmGy0i91t7ojXWf+Wld
4dgSaSBF+GdWQX4k4EFNRWUDn33GW0E/XjCnDI0DPw4/0nhXVrDiVmV8sIHtS2l/
+Ujg7J/YoK9UdmLDvqMrap8/ZdVxBSTQSLkVP6O7eANfAbVUey/HJk91SwNCeqIa
u29WcaTPiRMVad1AEVTUz08CVDwYJcJYAFY3HKh5xkXW4gtRUsEtujuBjJ7sKA8+
1/suzfTDWFdpkLv03z/OKuFE0ZGF/vMEGH9E1+8EWdsi71+0pVCKCqb14bz3Rdjm
6o+jis98n47Cw7lFiB+wVXDXLl7qHN1U1OWRqIur8nEp2puHDAYV/D0C7680kjsQ
n83S8fmfzrH8HOg3sT3v5VtcAp6usQuCo6xspwnKOGkq/zBG3qZjhPt9DeVpPyme
YS0HkDu589vNI4JrKkqFhEozIfdzNwOxc4BbnkGNS4oXmy8FfiMCRCvDeFX7jPC+
6Vuq3SqsKgjt4LAruFxpxD9Jg7XJUVhYfNqmQazf26TPyI6EiIa95umHusp5sdlN
dQmEIyrE0a8VbJ25w+bgWqFjmY6FuC2jJ+ns8YCcyyR9duaTtfXpqpNWNBA30VHo
jQGOlLDnLiXwGdWI91QbPz0naEkdB9zmtPM4VZMy0Ra1xeOUL/tQQzRCzz4By7IQ
a0HH8zZ8yLGuEOZC8qII63zJP5tpxGJgUXHd4bnJVh8UfbU7b18XGZJqnsnV/CGM
sSCdR9+vTgz+PwMN11AhoPgr9HL3Ll2vnHKXg1apnIPd6uNQKMXNrLlXD9RuEqkW
hGqgzJTBhSErAe0dii5BIe8rc8gnMy+HCrenOf3pjJIjLRz6BKCowz4I8iSAQpdL
MUafJbNgKu7+u+P8yrw2O7+iGUQmyr+LsjWAHnt+VwkDnui4iR0Z7pcu2kWTWjuu
TfdExLNihZQxQ/dYUwAN0kay6+Q9fAr8kCYGg0OzxRdgma/cbgrlYn/I5lBy65Gz
NRlYnjsz4pFvAHv6zY4HpxoP0LVxSNzJBFAdPgvu3CJ7w1ahbZ/ztAFmLmwHHEVz
JRLJly06tepP+evvkhXf6n6qLSZl1uhNteAe4oMH4JnGosoa1LEywywTIAgtZlma
Dtwp5sYSfxuubT4WcuVJ7jqpC9KVuqfPqJc8OtYIv6i2/DWNcjsFKoxH8u3VaeBo
sgK0Ui1lCiDy2dv2QYDuyrvwMZREcGnwaHDyfbSnl5zMUeGupZv0j9yLMcTiMRc1
dBmbztNVE3ezWOsKWClRYY+zO0JWA/rUysJKIpe+QHKaIuGWvGOiFYFBHGumx8rt
hHM5eHVXmdIOB5QPc4YxszmKiPg/d5/bYS1VFgV+dY+fwE4DkJuFwfXLamiPNPr6
llB0HHs7jUCDuJhGWllKSBpUuzd4TYxYltvvFi/5Ccq795usWsCFMCKL/G2ibmQC
hgJBTN4gKXhOJKRe8CfrB2hIeZhjHvd1dR6eVWHdNUJBuEzXUy3Ct2VuP62wlRkB
uOE3SC8ERvhQ37+W3kG88jNYktFyGYLbHogrlSWezUM1DvI2gqRLMdJHwTwvqyZD
6VQEf1vVdZ+UuaV4yVns1Qz8sl4gi6JfIoWnHjzL41melD1uL9e3IJMcmOZmAO3q
oAnt5yBC1MlPJGeAGv/xir6GINDSy8/uxqvtw21gYe6ShcjhyYtRSToK2Yg8ih1U
FW/1XEe6sIafy2MsYsZ5vsYssHjXzzor8W6be8ZUo3oyrmJ8YezuJCWjVlv2QqZX
7110164WJFwz9hhJWNPKeSJm6d2qAipshZE3FEa7tStB1vi9CqOheB/XFyuOI9gB
8+coqlRm1mOfQZk6WvycKUJyYKC26+dnvfuP/5kAteytLjCmlo9X5SvagCOPgliK
CQjqGzltGnmirk9LVGfjLdNxCXZIzovMw34pOsv2nSW78v0WvpBAODHdtzLoflej
BtygXlSOv13HGfEIrKjs3rx4Mlyx52PrFRNbgRFwiBaRQwqbxZO77bgsqlkvT/Z7
DtqjtZgV+pMqqgsK8qLNF9L8CM6ATCWWwCSrILxJ93y784B1c2iv3hLC8aNw2rP8
pmJU7jJl59UAia4bNt/X8XpUky8mAR/vaKR4jxA+XSAn/thqBfA9lCGYNnMNdhpP
7UsyX/t6LbYhhj8qYjLreh6X7Jfw3jnElcSeX1a37Rk2toRQRRc60/qSHkMyz2T0
Hp0t+rm2ZaFZy2yRonLpmYsHwfNaGNxeNAueqYKysWc4DbNusi3h0JgzSXoKs1fu
ORR+m6G0cYoKeBBtG9uW/uYvtA8ZOOfDAt3k64KK1cM2uj9X0RgulpVdN8JojDwT
Tv6QYYmUQ+rUbagpymOG8tnKmKHJkXKqG0chdAdGzWWynE1ypvomHM2cxEL/Z1zm
2UpurIVMaOG9+JghWf90B10A+OZZNmqY5kLh5jMtI3ziae4re1v3UQxPSSWFYUz0
xLc8EVexe1CxYAlBkC/PwNwr4JcnCG3v97LMi2a4KQ8n5u12ek5bjMvNwqeJ24M0
wr5EWgs6TYd9p2jNY74cmIbCm/XiBIV7pquBzJ2STUhnERDGE8pnzu2z/2aF9GPt
8B/ESBPknrfwG8HKtKatfhtIL3yQrT6Jpn/9r4ufXQEIMLU6LV2Cm7lm5pNt4UWI
f0Jqrt9Dc9GF45fDZUXn+jfYwCphEfW2KHHwMxUvMBuQvk9kGe50FW1tmUAf2lSi
5ZtExEfdnVLscVPrvwjw9rqQYO1Uj2cqYzeV1R62PNWLZve43OaFM+Z8adCl5taj
F6VPKWeUXeHeZEH/79166HozQsxd7BDylZWDum8V2ewjNY8SZyc+TWtXDecb0Ek9
3liRlIncqnM0ySA6cdGQcoLAyjCeqTy/eKgUMuqf39e0oSXe7UH1Ba8hT0CdZctS
jvTXgsE35I4kIaxTqgl5qp42qL9pRmUCwVejqTtQRpP7lxjZgCSjeIKaMlrPwuhc
fsfpbLY06x5wyxlILRWGwb/0SQ0b9wXcOOOTRAXA69nYpaEni21AMQvffUCqU3a3
5A3+l8x7vX27RMcnbfwzYF7jzaNpBuUgAYw13maGFypF2eWG774458+BE4Ae/xmF
WLmaywTc0LYCZlhv4u516SpssflQ/3wD6VhTxXqm4Ro+R7UGR1YYi3levco+/EQv
Z5+BQ2laP/HhLMQu+0TTttGt+yXdHUQgB1CJ6BBbIBJtNxgxWWpSfHIbHh52h46V
2tmqHCnojQm8PdSo/ewqxiQ3YQtJBdqavpwf8o/MOgi8Pt1jLxMv/nlLtsiwNyP+
h2pVKIyExmj+xEWYcmT3tiO8YXIUDmclJe8PDhQ/cmVY93cQUQ9c1qXNXoyO1DhG
PwuotBZ574Bqen6y4H3v1lobry/eKVGG/IkCgoH5qd4XIdJ2+Wot8Wn/+cDpWpw/
2LYtYB8dABM9vLxa+uTlooE5rVv7GOdmly8YE/KJpGB4DxawhPsKiJ6/wOY6zm1T
ZIqcAWe+V+pEqFrgfNToPD8sj7NA8P8VxohAnVJMdcaAbe/O4ZY6noCidnk5XDRq
9BOzniJBC08WrP3eeSoCxy4m7wf/RrV4z38mK5ufyoQAMf+xcqdTTmpzGYN250tl
dDiNlBGZvY2SNV9WWFchLoXqt2pvcM3Fs3ghKYMR7apraEdgG518GzlYJqVuittN
ra9DI+2LNONsA+h1kZnllq/6kkxV+iz987fkdndB3Li3/m/VIRWzbOHADYNJ9TS2
m48XtmSWtn06Mg+Ef156AuBLbSKC7i/UQbmMg6WT05KssOZrR2HsJ+SGcG/kj2CS
SeNGhX2xWw/q2GuPX0KiKEp9yZn/Zzq4MR2MLjv03RWbx2SaCLGLmp50J76FNs2Q
9VBnbxpjv1H6YVYq8TZAIxfj6cqRROvqdrtODqyEnuxVkaY//cuIW5sJY0g5rUjJ
huTtqv+npqinvQLx+kaCLb2AdbEfJbgOaudnoBS8sBLvVB5HxuLYLn7u2Loab1h2
Rsac0ShXUqdjanMb90PnN3PsXMsO+fdFS8sodrODq+dMufEbgfHE6t45un4MwR7g
2rKINjdmTeusEy+HSXfZZ4jrQ8851JddXRb5obfC4t28jYGiB2NfWOPMhEWNMqsy
kg9466XaA0fmV+8UGQw5MbWSlyUD+Y43K2Rpk/e6BgVaf9xtKjG+8PIONGWRjCg8
4eXx0YWE+3F6OZ7BVZLVRyeYnsJF+Ny/Yi1jaPGXVCrGquNdTpDE0TCfb8NSZA9o
pGTnutoKyMgoX8GWa3YnVqgTlsa2M0vCXQJnQUu5aT/z4IN6TC4fcTu2GgztIRfj
K4X5moRW+s5hZyvyC7c7x8uaHO3j8jyXkuTuaEN6Vjk6Pr2Owk9XEGbFUvwkz3UU
jcOmQo5yjNFtHbpWEwfTX9RImumfZcQQ9MUZ5+0qf/on/K2Ncoa3BR+1GcEYIk+1
pIblkPvRbgcWXHP/2qZRfKUPE8wQ9axq804ACeapHvYNPY32vSP4Pb+WgReKFUTc
MMlLpz4ntyeVcmJXiJS8f9rNBko2lvRRP/W1lyczK5UFyj5E8Oe5pdYxU7yoxnei
yG+WIplKayWhDheBG0MMvlTf5+ZHnRRhvv9iw6ax7oZi5szaXSKzSW2veeOgLfT2
pbTt0tsbLZ3hRLLnqmePVjoWeGZYj7/v9bgF7f1yIO7FJP8iaFyHbB9IM4gsXsU/
mXcT+S+vI2tBExTpa24VLI9yWyQEpt4+pkYxCSC3VNeDt26TUgXgSlBI8t3+vzgm
WKUUyIgox6DhPALxBgsuMFLWtw2NN9BvU4ZT9iZ9Bu5ziqSRJJL4wWlUDc2GjtCi
Ako/GL6FwckiuB7i6yAQMKWInr09bYvwZ4t8HSq0k936fLw9pPXlI6s9IQs/nzYz
x+4nKE/82BB5GWo4nymbhMB3abP5U51VpB4oZBPy/kxsmgjD/BLL6zTcY4CiOGoH
LRSZvOrYBRyYTMEfu8pU8s3/rSyrxZVoopu/knUxTqESTObVb40i53AKeVuY3BDD
cRH6zrfFUvfn6pSY/r+o+3mJG/4/LnIGyYJP3gedrTDkhjS55tiPabEzNcyxR6v5
Pby12voarBx/vlFysgkDwXaJjga5Bd68mh9L9hDIRtpks17K0iYrZyoKAp6Dol+c
SDvn+3BZooT61lNLRDTP8spavJUg4iwydc6wN6YdMK0NhLQfndaVeQrO1p353ian
jpW0moWb78QlBIOf8btyccmfK5+85/md3zuxfTxtktpSpVwdC/0x14dAzJK+/eir
mSfDv5pQhyNCaB01xFSw8EnajEPTz5BDXKAZOYcL18GeXYcLAs9C9Ai8McORFpiQ
8QvSRX8ROWkBRTYDREQ13UE50BoI4SY98/pGC07igqkA/imsrQbyjWasWgD9lRzA
cuKzVqiKmOyQQVV7nIV+iVsOFpT14/jSQpFmScLOaww/Ngp4T6u0bYXKD3cJE3al
a1/R5tXzIuMSBpqwqyD/q+y37TwwpKYDZ+BXGxFAmCFVYhtDWnx0asUSkQtqsNmI
KwEVLkSUdPlMt948MWpNvMxgNAFVc0IeFEraCDAgAznMDRyPqR/FCV2VymfumBuz
DsHvDbjdt5mOTExWgRDkpttm5Pmx7TEyEB9XtSCJCh6msyzTx68SNxn7H6IbDNBA
rx2Q8IjJNkt/nwsA6SvE3GWLe7E/h/F+suegXav/l6jjdSuYO6PdOzwY6DZhvaF7
loBRGjQE1LpNb6izLYFx2ROvLHRaNBwnrgjDX3VbvIJKUzT9lq0e3T7/vG+yqW5i
RJnhhtovPTUM2xYTjSXCbFb/gTPbHtAHqRNiQv619lkMbxfaGDGEru/22JronC5S
Ee1QeooOTJr567Ly8QP1CKwIEVG1uh3yM4MfQlbDtNR2NskjaWq7a/lmvzyaAeru
bpKf7N5OiKXl0RzQAvrYGEPRL8F2xXV04JeGX/2ndIuYF3m7dATANsfcL52uKS7R
1/Gd+CHNHx4DBRh/Qa83NAuJ5JZmstDQ5JzE9SjjOKzCfLQEY8lcvs/CfgFO515e
8mBou5fN9uz9EI108ZgmtcVdW0s+7RcaEuxAfiOoALXI02Cuc272MJD+h7IBrUgX
qtHKoSYaTwE9viMP8HNJKPZvVVQmSzynJ5DwXolULOUxfu/9BfnaAZ3AEyq5Pd/R
W0l5fxDRIw2s9ei42z956c+eJjOo3+IfIJtbW93OhDFWp01kxodblAAWIboYzof1
RFS+uohpEKU8Llyue21BYLj/EWHf8hy/sn290w6gyGyY/cRlCgGtt7e6hEXRNNOX
09EzTvl5dDkkRhXQEC/gMEd4iCqZNEK/hrTsKe53wDen12PJdHON8cR1ANtEw+L+
JMfCuc227ToOsXW8YqNTS1zhEvwVjHf1uPuqACuT/1gI+UZAZrYS9z0om+aAZOfu
+tB5ikKkWctRbK96PoJ+Y0SMoOAwGkbk+7qqgdfN0jWvzG0++BYNnQjcg9iTu/7O
VqXAfzUsz+ru7Vq6pSwRvZdUnPV+M/eikvFmjQ0d4tzgtRJ9n7uyEskTG7euIaKs
DaVPFdy0Qc9bmTkZO9wOQHpHpB8GtSO1OSL6HFHZpxf/XcdrkMYgyHKw54sg7kqt
CHBfyjcQykquZw11fxYSLlY7sMFveKRbfTtt5okgtFX75p6Gt8s335cji5tTvQS+
R3P0ufamhlpHqKqq1LBnIZ8MvFbFtUEFDduCbqXZ468LLgLsH/bcMC0KihnS+MGO
l/gYoTu6Ti2mY3wQMd0dCET6yCLaLluo8Q6byRVzvVug7EslXB4DX+FBcsyg9bZi
DJZZfFcswr+t33SQB3YdJudaxHsyZorq9QsCXM3U5Mhfhdbpt71YerPEqDz3sKdA
Ii4DuqAIhWL7FkLx0OJ5PdeVa97WT8oh5R9PDFNOacAvgeAfCKQ9b0Ufw8Lu9/VC
DnLVYbKPbVOmssdwRpqhPENsES/cZfH44HpaF92VOv+f5RjXBK8oINswkeOqniFD
QrW1Wz07GuOoI7YDFlCD1qPteBA+NwRkDhZtZ3HLaVE0zT4FU8kkTc7zXyHtYtrh
Kt0Hz6aAFTkruFLr3kC5iX5ys5hhgqxpQXn8Q56kKlEulWld2fzEUhHXIK2tOgjB
7231ogkzNzOdD0/WgsBfh9CxWyr59l8NHkd1G5T0OAgB4r+gi59jh/WHlhgpx39M
8TiuQswcTLImSYnomGRv81gfofeGJ3/JXqgHjzHs+8EsVEYlT9MRO6OFjv4xMvUN
9Qu2P2HPsCK2iVbiGsp+7mnMvfvj34bsJ9c7T1XWBFKZabPumHxhnoGKhOoRlho4
+xcAd1MwXSaXnJU8beforUBLBSxTmlCuVo1N9aaRcpgriEbUQc6iRTELaS32FfCj
x++A8EtXik0ZeslcCyD+Bp9a8j8SsiHbS95itbiX2mGMq0R8EF/TuL2u9fHGs5KU
mKC8lRwTPLewQZYss1+sWLx1v66KGZG41daHFGaAD0a/b/7AqHvuzvFJtWPaSet+
A3WaP9tlEt3b9FxmtoM+ubmLyHWePn4bXNSqR+wDLQ8ISJRurSAHtzkF4J0O+cdi
DHs/626PwuXe2tsprpMoHsfJaJXkuoLK1a7OhNzxLDBjUgINYhsmMNeosFaqTsU4
f0U4GPcaBmW+rhqSchSa2nwQ2CJyuu4ejjBySqs7q3XM/XZhM0PRQT/ep0TmwvEF
7JWJc9UnqUw/J8CeXza3EOFIazU2ndsa9oRrWovlr9tdHoYKLMhujJevUPQV8Jsb
ZjBJ0FgUOMCi43pEP0UgC+qO8eSf4ZWqwGYIwd8Zkv6Lc/qxHYl45t7WNo/PCuRy
WowowpLl1/wRF53OALYbZALOAI/VXTTql5jfZ19qs0gX1+QAoqggoaoor4k2nhzI
gZoeiNT6lfNIYl5Fs51vebeMHAZQS0i9kWNTvlT787OC5/4hjJOpFO8w8BfXE7Wz
6YCLOQskfqcdBKCyC4dbzrOOuEUFAn8fxtezfobTaxYwRPZXOnmJrjM64IqDAo1J
1+p3q5ue/akts7bS0ch8CU4kdmqsvHa8yD/sCrXqRbGMxtX74pKf26kk7Rowqy68
57rwJGFvPIZtrneaWCAPu/I12/4RteGNSVSPteEOf8N6HB3R49rIDX7mTKncWaeX
JjErcgDmiBN1tSINqzhAefijDtU1HxD9FMCDlr2+uCzlZtjMsBXnReDMjJ9w4Hnq
OANfYoj7yf3fMVlkYTaUtK6GVj2LLTva9LaTEauOKiOK7IfIrgF/JynW5xRspEZV
2C4svYykpg7rYOpKaFC8Qf1IXnPLnwoVZ0pUDmUqvr4BJ4epWFAUjXPoxlfAw7Od
kjWb8YSiOhYjI+GUngYljw8YKEiZL3nDsEbqB9OwZ4OkhmKvzD/ldmPPevsvO6sJ
gbhJuDBn+fGqbPk65xplNLhpMXM+zSsfg3uP/7jIEfhrz1py+PQ78qjoT6hnYkBx
BuUZngWW0AeD5WKCXPelwdgkJJFa4QUEiui/XR0XDKqJeNzyd5778tnLTM1rRfFN
IYU4vb2TV8wZcDXtvHmhmIC6a/+H7J94AKGGjUfG30X4FM3PcMRnj2OlnqiXgNz7
2p7w/BZ13zHotxIx8G9LnDr04IpPY7qHKDOMrev3c0/+wfX7yK+mynmgTfWshNUt
W2R8ToANhAA8dj6xaV6UygzJ5s2OjUDIq94MAHK6suBSBH1CBc3pXXA7YLFJe2nK
5YskMfwKUPCQpFt2ygpTMkhzw/PjEO49134qH06UpdSP6zAL9PvCCiwWhIMiBu+x
b5x2RghOnc0UTztQ27DWE2WVCVB1jZHJ7VJ0u5mw1JdU2RSPpACYYkGcXYXq4pbc
ok0xBgSDnpFOvHB9vTJtJSrPw8YIgUtHHeXQuESm0DppP0GjLbgrWZAgaUZOAv6N
vS5uquEjuBEATe+Ye/fyB/4VmcOTIDaeZDSG5R9NQM3IukzsFKDx8S8sqQ7/BCOw
kOkS73UPKL9ozc8CMNbK13HCF86DPWuu11/wp9S90SCXPjwwZ7Vx02+QpAr5zIv2
eXcAnCkqE8KBz/ms5MBwnEy1pUxarJjQEuwlzJtA1Y0Fe+DQUgWVlJwh3IfEhXLw
HRzyJ4rGsbuaSfub3UhGiI5fDa+nC+xFcEs5UqdOtMRhpjP+JgmbPtfgPkADoeds
uZKaPxpmTj2MRH5t7OXwK+pjN+dvwnx0V+l6VJbMmqTWS2ZEYc5BYUBFRpUYnih9
qy4vPcgKT/1TjYgofsJ+LszV+f6mGKANxWoI02UKkuVPFjTwTUnT0W5KEHnbwKk2
zl/RZ203zb3pwr8Vf3WNALsOsVf3LwlO5wc8H2w2ZsSXW6qMyYINoLH6IvWsA9OT
VYD4yG3o7pxlHiqaLs0s3hZCIeR9V3fhNLUfeUdhCTLLQWlHlevxQ/EpuSNvJW+I
iI32V8Cr8VzNWMqwF6gsN2IT6gH1MeT/rsE4WI4g3thqPwuy0HaXwPKf2qvjhFV+
Yb2CsLaWR7U6G0NdC9qrBt2BoW8C+mhAwa+wpgN/nxnT4JLRkYgLjERdeOg6WXvr
aSxtIc5r1eDSr0KnpHTldQiLolcs2ERa/ID455CB+BUOWLAXMnWepl0DnphKj0YS
8izC3t04OXIuFoKQp+ddn2Lg4ZKnRKPC6g1Wp3EL0QocChVK+TyokponACYTgctU
b1yXD15TTBxkXKLV6cVnln7Q78id69LVTZtRrnqLx8VWh+1EA8Os2pr2q1LBMArR
vB5mXTGnYkA9T1gfKD1LWrxE8kYeIgDHCXXqnd0il1nB4CfHUtnjBA5HqN+JGSqE
9tD1u7VOGImM+XWfXqwxRCx1065Y3H/g03RtRbACBQOmswcQgdtyyuIMKz9ZQg5y
FdQr1o9/dRHvXOxmVfptJQmKGsL+YwY10TrUj4Oc6C1y7YgzuIYEPlL8RIFDTNfv
FVOKSuRRsAWHNFe1xnf+6uNOpo0u5DKe5Jnd/UUHnK5up3C8koMtVikjN+0cLlq+
nAVh+KbQqG83aA2cltOqUs7UTLrvtFsC5I1YvMLjSe34c7qVxRSVp6ciMnHSBy9w
w9WHxC3aUYiDSvAKYaT/eefHbn16nCu5MQ7q+J0bHstFbf7JI7VSkU0FSIKyzdCn
uZ6eK3zvtukoTCzdjdrt1ovHgvUDsV1d3Vr6qmwxLLgHRSoVkA3lHJ2tpHsV4LT7
8AVoNY+Zu/agB7+a+oZbYRXb79dXZ+VTTB451VIrDTHWVMKbXY1b+gEsKFj4ZZCh
vvJC2jHh8sUvDswonGzgCjD7N97UpSL1ShNyiPI1N0WX4V6Cnmrf9l66RxkIPk/g
V22YorsFdE1eV7H3r+SBpQATqcbdtdSlMRoY+9E7SinR84a9+0KtcDqMLTaK7l6k
RABEAK292qj88Q0boPR6tdNiGBJqE7Yo7kjQPmBBbJryIDcN3xBsyVKjuvZD5oN3
ixeAUo2AjqEFyWCVqMhK0nPCqkrfaeO8GugRnbMwC2BfolK+KigLt0FDTCKGOsfe
YtMe9gNtcXy+wPNFjr9EfewUcP0Fu1ra7lCg8MLid4WjO1ySmzjL+I+wk1+YS5XW
IBfczSpcDA2kTOSx0A6P30Uq+gJM0DiDBRvUH3V7TALKnw1Sdcme38iNz7LzYTIV
qiU7/nIDJ99pOyIuTzm0HTr1zyZsxmXQNHUfIoU2MKil3hhpJdDECPDGyLxM3DHh
L3h7ZAFHrHqSNjbTuGbsMZAOhy3CxW+Z6IZYvSCAO6BjBu4UwTXfiyaAFZ57KP/z
fzO2wDw/BHTXoCVpQhbUBfnsPGF42LsYk2sfUK0DnZHIAk0nagzdTPCjlyZpUiQV
3a022DxqODrRZiBT08g7cMNXZ5Hgm62iHYGruyTXi6zkqnHtdc/rEj1eDlve4FsK
XcXESaU+2JYy6CyArzVMJrBN13HsezxnB1+b/ceJO/P8L/3yOGcUYRPylqCuXyfw
uUfErSsoZq4Q3D1/z5uPhW61PiTFxMZqOvaJrO+tRb/svZUyNjaAA8FZubV3oW2g
rh1fx8028+vHFKz9l9xb8sVevQ5tM3HpyF3rm2GsXT1l1N/BJx1PXTItYSqMBvnw
HtXOvi/UYCmNV+LSL02m5cXfpxk1Kj4xefJMTE6bbES2ThFrO4SmVgzeaT23DaFQ
nzLEiHNOR7h7RBNq1MkIYuuf+W9zAMDUXTGbQL4EV80jOuq4NwSs2cHzPUiF6+wy
z5VW8UcUlr8TbWWSTm8g6mbN/5WYMC+D1fOnqNc/HhB4vTpgp0KBZ6Y3KwWsfiNU
a4h1RV/jo8UbAm7VA6PrNItXf4ikNldqU875Hv+CgbHnem9Q7225zeu1fyoL5A77
wRgyhCl8EkOKt2iAs56RwVdq9GeyqpM3DluxyKgSoOJbKhXOvTmMjDgnSu+iKVFi
AbKnSeTTSxTgSJEW8HQOLogE3rKg5A6h2wIg1SX/EQQrV5johCpq/f/EsiSTjfKE
QgjYLyJZDzcaxuH+4HwUrM3/aBednKzxx7859yQRlXqqkIrB41Qf42zxkwWh79Rl
hstMN1Qmm9NDGI5g2tlBJu7rBoWGMY6aOjcvTaBAjnPyMbyLrAcEYacHnP8UBppg
kz0nyZwVaAfuZU2+Lvz2ahJEPBo3xgD6jnynmIt0v0qV6Qd9lVgw/nrAb+OPYrsf
ZqZIFweD5AV2ef6QdaS4Y9Atz82jmCbLNTm2zJAaGEB00DOoGNSZz/E5dS4UTCGE
pTpCWHY904mjY/nbOZ8csczGzsMri9PuCSXcflziChb98uV36hGHrjIVlUH01E7V
1kZYT8tQzMP+bZ3iZFeOKp1dlWEzYcT2ex93P9rLxHa3diyQo37XakaQshjqsdaX
KHRCbRndPpav4tHUe2FG9cGW1T8HLLtJq5C6HOm8A0JdUMJkrTfyK6oUoHyqo4n+
z6wguQEVedbVNGVoFuDShNoGv5zBD8Y06tjuVDqf5nGbmiqKJrwRdHg9jvXcL61B
ui+2Uju37LBBpoYm1mpsWm5kRrl0g29vLl7MLnZTEfcTUD462lzA2tUgXcXwAjdE
npTtmSTlLzwq1kJgesadic15dHXA7y/ldE2HbWdhdBtvIVkAnhNfCMN/0a0nxm2+
lhgE4DOBHeWviYWKODJG9AXk+WrwHZOw3/PvL2x1UTSvgRpFBq/PCzS4/ApVkswc
RYBC5TAzJTdJ7LGwmHXthe+EQRInwZhDN1H9BUIjiQ9SvIiRjh9Cz7VgM9Tzy7Jb
cTspqTYnnTXr7FOqHBSXsxXtoSNcrFcr6KTFK1VQpxiOeOwEbYKjS6luic3rE2Ig
F8zKBguwjriFpk0mcHV5uhmm9gJClPEMOX/5l/kgpmgtzgQ4CscXa/3ys/5tjy56
X6YR5OU6ZRozuWJsjDIrl+WS85CTF/vFAUX0ScoSRqOPWqQnHBoFcOAHuSq9sGwm
DiDCeKuq3te0BYrD/5/b5w8mXsk5GxiAor+TMqmrPpi2357gKkzN5S8cDJ/3/sn/
J6x8TfLNfeLXkHPjPGuJ6tr8uulpOtybLv+sME6km8vSBOmC8wK4lljZYQLhGZ2Q
8mNLcPPG8bvAFm56jAN+N7UfcBLA78DvsDmUAR/rIMflHcZRdOwIA+J6vpCX2/jM
5fupNgfQ99+VaVUyDvAGNGJfsptP3uRyQsdlmBuVjXEhKF+7WKkwiz6Gf3F82KUA
kJdw67RoAjofYEADNlOMv3Axb+j3fEQ1/79iWYMmM/67AdHeVr8aROxcVs3Wzly8
mAmg0qctq0FQ2KXjGsjq5LGIV4gVIJFw95TYxBq2S+ox/Q8FwWPnpay4xDwP3kKC
YkWY3O/oSm8CjRuZ8LNDeXiImbC28Lj7LWNlpEeUSz8BJAj7BfrecZEBjK4WFqFM
/rj+s8OpyJjGC6DgQzj25GO5NJXc9OOdE9LorTZuNRed+2i3GLiFH2vgCR4u87nr
2uV+84cOtYJhUzZJI1DjsIiCuu05pnylqdz6l8257Lu2HhtvZ0OHpWUGrN9CRqvi
BfgJq6Vl9qMgfdOoqtWQ2bjT3cIFFrv0gupZWQ+jokyticH3FYweWNHNVUF6EfrY
v4ZtRgWc0LQ03UYfVN39Obzx1yOodDQtOqqO8vKtmQ1AL0mGSzZ9KyRF/QadWkkt
i85d/nJBXJ6/t8O9BAtxVAEZAoo3cbXe7qP9fUNYJ3iNxQnDd6mSyW/0sfCbE8jv
ge0L++xrYhw1uMUdGzYkuK/MubyXgOMmPm91UcBrpzH8WQqRAlMsODezZ5oRjCZp
tFsNhy067v0qReD7Ehiqx4HJnRL/xkbupunBJI5E2ylb2apFkTfYXbNEvvyqsmBz
IDeMYrJQ5NmQV7worMNcSq/RTdsKx0J+cCui0scmluIcdFRcNMQ2yjD0KrEUp0Ij
VX6960d335h98wqlyYAtdnfT55IareBwgwi37VhbGKkv68YMdynkvP3JCZQ2U53r
4iw9k0SySeUrvvHijFs5Z0l7VPbB6MXn0D9k9Gra+uz5S0/z+85GASstPgcflIZ4
T0kRbQKQinT7V4EBFDqrFysSxecjwNaSmzFZ0awqfGwuk2h31t0uTGNoq+B0XUbV
rpYvsDmOvztr88XQZKevTYpGGjIwaz9vpR1nQG7vY8/LPeu6yx6oAE925h2omt9r
0k5GZOm+xacnOQoKDNShKl5U5uwhRnvq2uyUkap3pprTPPMhx1Y+YsdjdaXMCZfW
BNK1SWMEf81Wzx71ha68P1KNzEiRf0staX/nnbOLtB2bBZm6Iwvz47CWfFCkntEi
hQ919VTxX0yLIj4yjENwk3E1BuMbR6C4rID2H53ccFDRNwl53qGR09d0JbKbOq8W
RTJauzTFiNWCAdwh2HIgpxAWLPiCdP3RL35KDJ8IylbSccNVD+S1wobRsHENP6Je
9d5bfxK7fScDRInn9B0v8G9SaEOKNtHbDuncpypdbt2b6sJiMKkDGZBFB9FFcRNr
ZkO3Wjh3ULixURR51essUxIFaOUKvWKAD89xRRFt5v6N1ycywFdrfi/yESJc7uYU
Y8M9vSN0D2mkC3HkLroVy63Xhsn/axqYgmpaKAdqjNJcDuyKsRpPUukV3bFQ+BNA
+qyB1GL4zWsXkexljzxL0UMNbkUzIO6s6OUgfXNhwLT2d3YjAi97eL+fIY93TPHk
n3LCGNL2KibEO3CfIXmG/kwICtUzGC3Pa0sS2m1cokhAUVeAiZmvWAjmTN2LmXnp
hcE5xiKHUSDst+rnYrC0BuM1bi2OrXUTEIwKFx0xf7wz00GGzrCpVZZSxMKEevLg
0TKsNV7NFhzDZ1gmiE05uSp9GEB/apoQYyPMo4YcRxwt9STIR7jzDmWDUNWNDPpC
irX1jd7Zc0dX+PK/XrM7QGsMnFqX78KTrhz5Td8xL+FGomIzry8ODkbMCbIShVdL
OyFquhM1cynbwjIjWTrnmr8eI271Inc1t+NOzFJT+X42AGuv+7Sqjf+j5ojsevuu
m+ok0Za339nLWKbVmHWOkVCZNezhBGxJ0xOb1T6X9wuHY0OgAQwGl2kK0ElvG2sW
pSVVFx0RgT+0/TBpq1YhTmQLZwVGPnn0UXVF+AWc8g/+8pL8KFbnm8PVkVcZaKQq
G44m8G0w599CwfxCv+g++thaB3qRPk8BNdDQ5kNln1dOlI4fNRXL6MucmY78ZcAK
BoaJtMwqJZzpPRqcw1hM9TIL3vCza6SDivLU0Es0VOj/AlSgp4fT8FxWvj4U7lwc
sVvWW56sleqqVdy4Sw8JiRUAvawfZbXaVHjtt8qNRg5J8nQ1JzkBUU2FCD5HUw+J
aHIqIL/POZ/uI9QNHqres8lhahNPOAx/t9+Bb4G1Oea6AzRPXLcHOG60NJ/isBdf
vpmTIRX2BYSarGgRVEFlrJplbw5N2KQveY3gZiXN05Bm+aLj2jrAy2yQpzB9SatR
4L3uwn38Z4PdU1bAh0SrDLrJb2xBnJiokPum0zW35pQl73CLGDO/FPGsfyObH6sO
y3E8X7da2x1bVY87gWfv7tMytVkDmdenzS0Acm9ddwYmKDTtswA5LYn2o7crkP1c
IWwOv2WA+7ceQuZwBiiecr1PBCH/Zzn4RhTTuseFy12unrbY2r+yXw2EmLYR0qXG
Hqt+TFg2sNeu84XZmZH7va+jkPzAw8LTjjU5uGYO3ON2U6cSXPyLeYq/nVhLDRPQ
BiwExIDRAoyN/jeMsRgqY3wOkAuj39Acxn8pQakl6oJOFdIkVs16He46+llnFnRU
McwWpm+vkQECpXHuLRRlixrnrHV+kqJ9dkbJExh1FImCNuTuPkBJHIPMpmp1Uax3
pQ9m8+Y++WG4XXnycUhQEYLBnr9b5/ZKLewEF6kflo+3puEvqjjjrBDbUXqo7EqY
sZ7moLf/kj50F52dK8r9CRfrSuVBJvJuZ8XV+1LWVri+NgXuPWtZvROvXK4THleK
eBk1vn59lF8utxnMBgr0dN6ADyNgDyviWTVWLq8URXAqzIChCSwE2iUGeccUVAwW
9CXCfkHkbme05kFWjU1uDLG3exvBpePDN7Fsk2+QABYBNPl/yc6j1RCpt46EgvPx
HO2La04UhdRAPZhc0wKAWj83Z+frph8hhQtzOVXS5DopRQuqQaPh9sP+KdYo7kuI
iV2G9NNTjINCBTGjSXwQ3JJIQsYf/RBJuwhsg/a06pazt53IDkAtgjDNCF/gLF5O
V1MvD84tCwGLwTP1AzSZTC/THqxMQnEPQLdXcOUzYPnIGf1Cf96MS8yOAk2s3BFX
OHixXXXSOj5ZaulqgQiF3b7USvrpSzCrPFtvQx6BaIGNEOZJOz7jmoeCgscFFRZ5
40hGW0ABcgF1ywK0RMU8x73myuCufj1skL2AHFM3qwB3+lfW4+NsvSzvLZs2L7H/
rDMHLPX63uw5Nt6XqPKrGPPbq8gcDqUwvdimWgJX0D+XduZRk+bB3nobLaCASgxu
6cLmPYUYHKPMPfwMZbBTL3odV4Ot1uOefZulJvEEVAW/vUxzY5HGOH1CYOG09y4h
Iu8tYJNbIOnLJVo7TnU1ROiqpgfMTjzNkq0dxxDsmnxigHecopQUC5HrVkgW2A0g
yhG9O1YuHKCythE4MHg8YOZXmfKA66Jsrjv+3ShkO9/XuLm4FLCiRhhiXQsFXkiT
2b5ypyKaEWAB4IHeWyGfs7JLDdzlMFHnKMfm/aZpKbhltaodoa+gCDAC5zXLpzFi
MU39QxVSxOcZ81gSCE/UWMmfJNDJgzAiFtP4fnekGZISfTIYpuJ5P37VtP10lbKL
jGpJyS8iBlWiZrb+ItUwMvqs3nn0WVrSsLbQenvtpMSx2fp8pTat206co+lbSuav
JHvkbTYQ8qvqoK6MjQ0VC7mZmR+1D778fUoQPbZaOGPuymUnRkEtmgDdXpT+MsDA
5diSyA2YJKXAIx5+qHiJ9jxS3Japjoangk0/LmjX6U8jbx9aDZ5wySSDsHjmP8gb
B6JYX1ghOFxc/xsOSZeF7uz7P5iO9UJ2XKb8w8bhYOzgR43JtrND3Fb2GMDvBgLb
PzI2HGuxh7XluGuJsytJD6j7CZAyMG7U5dbHSPdcFxl8NxK8BecywSmkSDFn7K6Z
rebqJKKvuSygafazYqiJAd0X4Y/NPFynkMzX6VNwfxeyQ2MJQS6mExd/ZkW7CEkX
j1UCf0PVWO/XVl83RJrj8CV51Wk9MUmDxbUkaefQDCx8wkH0yOiCVGGsvdP6gBA3
A9Ugq9zqAscBowZuZsMEjNRQ1WgwtGUuHzldOEU1/VX4Xbl7nsfoDPqFUnY3iPFJ
NQUEToRwxgIQpOMtUkE4M3E7WpLgkY/41NnMUk+S2QYB33yFBPyPgIfrTOd5ORZs
tjCdcdW8NpqCH3SugCYxVIjkkytqkoarjMp8bh84f8LkyvySb7dct/RiFNAeyH5I
aYmz7dBcoua1cH1a/FaY9hr6ww6f47q5Az4/3tXR2abK002Zh6I4/yS9P5y+p3pg
bXPFvwKHJww+OVqEjci6LdprUji6Eu8lUbmgpk3NGJ2pNAHmCU+sXXgNzixjFA3U
XoM6qBqJ1rtXl8SigoILX+7uL8c8SmVvlCm3YkTh+K7GRavDoWQ176cVCts+Ywds
V/pjZSxHTqAezsjIF3xtzX9x37JvsZSHnbhI1Q5WZ6yE/hrRcd1dGwCOyxKiXJra
9GVNRbbbfDTWCD+D0NpwUgItNFnubN7C17wqt020zlpWU8o/Ghfm5F6wKgq5yfi3
wD3EyTSn4pwqCCW+9z58TSAUjYZZyxGSng/AuHuI2nVJDW8BTvQ4wRfN2pJIBoFm
eOq7d6HwaPVzkgUp0lNpL010Lr4R77vfHUUC6kHXsa5A5oTnsRMGIB4yiygMrzPt
M1G0EYmr9irTVqFbrgwb/1eSkIwpHouLEQKOex8orUAIgR6Xmi/6wZeJP3kBGpi3
qd8wuBy7QVBwphGHqh4KToCVnGYwFqxN+8FsW9cwXlsi/2tSEKr/sJSu1mPYAIiY
uuX9WLgiFp+l6iVXxh0HLa4PeeCFflcBRU5/KCX58E9HjiI5xpyyogp95edHXxJH
0Bd56mDo4IpXXI0uxKgzlCUvyeogc/7iiyu7laix/y6tjAKZ9PMQQQPzGgcINY/3
qTLPy+6of5BDaWqLsTxNrb6v6lY0lraua2hWgydAmP2hNIxcLFHGqJYwGHRRArAx
pk6qI+T819zytmkraV5QS893JHc2tEH+sHKIoD1oZ5xFurdL7XkhHQLpYnVPQaH6
Fufv3V4PdzE3H6IaY/gM2uH6wJyLMfniP9frDQYKuX0XKvT7cFvDaXDCBcTgKYfQ
BkXvUfbIqj2JFnVMtjSs4sxTpMdaHBGx7ryhIRCpnPuN3l+m3J/pQbfzPWbEBaQ+
L9gNZGV3N1NdVr5KJ33leeVUrvMw9avcyxP9/x+dU3BSuIBuTMogv6QTuM7DpOl3
rj3zJTgflUQ1LkgmeNZa2UTk6eZYunBDh/bPESeKSe+wWJgei9L+m3MTVyOGmtUO
V+JRpsE1n7mLu00gnCpZwnPBv7IsjrYHNwFn8hXWJ8UPcjerO/XTdhFhy9XTuoJl
nZEpucxUZdA4x0LAEJvfLZpT9XjCBm1VMfRcXQi0PQuACSDOuzDDpR//z7HWiO6t
JQkE3CE4Qcx6woeBaRTWCFuwCy5tn/crKiE0zUoqj8GHdp7WMkUm46pRNwcxSil2
NTaEPKKoqsmqmnbCumJxkIJWxNFWNHO3RibZvHt0nPg587AkZyjP6+k2ogFJ9QEh
F4lA4eRYKXq+xEGljRcLvQ0gwMFk5MuStcpKN1Qkoccj4Co9zUAhvgjRPyIhri1M
iDM4bTBzCLLM8w/IT6SaSTnY7+CUmFZ6fXnW/YOFWEYbNkLv6bAs2LF/jIebfaIf
yzme/oopMduP6MXzfzcE6TNnCZALLufBu1jC9vFbbLZXBxPato+tJHxBcsk45Vrj
Y4147MIaWmyy3nhAO+4u4dClK9y3XpAGb4AMDC6AvpQcmtna41qxNkKM5Q5GuHgs
nBA5DTj6jrOUWGVQmh0HwbruygZM9tPtYLa4goAboZM5oSSxxTSywmTmBDpmECwe
G0dQWxzbyXrhzw8PrUgJ1ihXpmferXKYGI6hn8fuq0cv/PqvXaj5ccPv2pHD1fJK
0cOqj2FAkYvP35nijsBWbOPXIcIXJ8NzQdCLfEMaLXyHioD5z8ylx9IX6fFGWkDO
n7aEIEKoomwddin60BHTwYAKXhF88EqHv9zgV6UJfeUuZ6S9uHkFfU9S+DQsu1TS
+BJ4lVXo4Iz0HONZbJyMqznU8+f+HfbkAbr1OF+neNVuZPboD7HG2x+nYLccV406
hZfAAQeLMLGF2qnfJIthSBqpzz0tdmuI+7AJdacF9K3wBRJqYp7go/2qYMtvoiAM
HRKwbhC+RgFUT227pQtGMXM8tsbgfzu5uD7/FvN31zFkS1d5cAErI17E3UwQ5Eiu
fKN4Fb3sRHRyH0rMaHXH+ntkP4/92ieffP7qLZxPW6eJ6eTcCnZcFaZXvskGWtht
PqBfaZjFhUJv/2lqOBNk5kD/ZuZprYuY1k7sz7ZvfDD+H2SUt1wdYI+uFc8OgEpU
3Qaxo8Rik1Dd+4zhPiPBy+UHh+vbTxi+eCeyzmlvaiE0lM9BFnSdQtOXSaRWnoKn
rSHgekihvgbB7Bm75qRWpLHB1XVH7GXQscbhkW+X//FNWAaIBh2NL2UBt1sMD3RT
MzXVCf+0ooQrpBR7K0ro2EiTiiNwlBtjQUsuOKcdgAqfbbT+a1D0u8ajltysHAVX
FnNGtJGMB0t6qSwBeTOcwzs71RwNHB1hHfP0auQZpvQ+Xvcc/blLfODU4J4fxUuw
+IU8tCut/N6qwcHWcEX7Pvo/usNv3+C48xZav1oq02Rj5avWUrRDtN4yBrX0tD3Y
mm0Z4qQ69olXT4S9IQyiqCyIYmHAXYhMg9wY3CoFKH05ZclkW1+cahMojDivyIBB
4crP/AnObhvHsJruv9qaVMKoE9eRAxrUhUzWSDgXcVm5T6FX4gORUcMh/KELwTMJ
hAeHRwzPwyDvpbQ+FcQSsTcM5Ge0KHAQSrMxtBRBVjDR6CFMHb9vdUc6a0jDbMAt
BTdiO2eqL5c/NHJmKdbv8QdFqOW3yYwbSgHJ2g5eJEqsbVRb+JYDGcQ1pSKjYMcF
hp2lkIOyWIh+P1eUmM8If0VxieaRVADw8ZhkrTu4Qn9JJWoTTQI4DIfkJ7R5gZg3
9fW0i6UNWJm/kDYJ9dcXr02KgDnMo99547lw0VZbMM5ck02qK28ZzoO1UIfNMLUo
m2NTsoa7wfeTCLy5PQdjIdtyvLt0FG/HaHh1rAq5WgRHJAefRlSFuRbKlMt/FXHb
bZs8fkJc/fCewAmzJHMMDrtcBO7a1rM7YZKV3SCXKr5jNQAd76P2auPuphKIJ9l8
Z2yt6J8woLARnTz5X1HexHBnoaZFmii92QE78g2beP0ceBNVnXIh2FhVW3beepbn
FuvlCmP1J3IFX27oNdUfi9ndxwwsn6BXI2cirKFVqHq+2zL5PU4eb9A6/tgY/naV
S3nSR6GiLatdo1d9+IdYRVqOH28Q6YexjiMIqlm9agHxBfxUV2/wmsvjzylJQw8B
vB0xlJ5D5Wv6NTmuAEi1+/h+0qo4l8xMkRUea1IQ5zsgumBk9xOx0K/xC7T/+dGr
Sf224q/Nv1qNhItWW6yhwLVDbl8gNP45RexUklMfDCFKryIEqYE3M03EM8sINh84
BJkkTXRbRkbGa7ZwSq0Az7zzvVwCqF+GTPTRIC6F5fOn/np9rg2G+DPiWa5LqJwx
3W4U5B2N3OsFe4qFq8ckWtZMeP8zotMy7RExvpp5s2WXEDlpAdVwKGO6b5PJsrHk
Ne1xK2/zDZe/lUQvM3xuoXwNA7vZU4/E74n5CFeRaDF6b4zlhdB/iNU7+8xAhbOe
Veg81srPOlusb1jkQMb7lzs3lgYebk+RET6GAsIcvL48HQGwa7jmuoR80MXwNoxI
tDhI0lPY9ZjJOwLfrhgXm3IwhpNN3C1j5u3aHwOr4uDen30iF2nF/9quqpNzwRJA
F4e1HnTxUrlxHuWcek7ig50UfedZ7okjJvCEiF39yHZPvpLzJAa4sEqpz/hBUSA8
SRcWYeN+KDutOY6cZnCBEtLewyBfMEbvwWJWj4fNeyLbeNYlKBFaHKjs24rgN6ID
bhdCmOXC0HvCsfJrhG2Cuf/wXN+gDdY/rsO4vBky7gQgrvLTO+C4TF/Um2k0Bl70
N21Hr/rsbusFBu7nXtiWNFrc9sa7FtTu/00Np8sf2XFeJMmfhwGgKKo787D3UX5s
+7xJxTipDTBFB86rKXt2H/R/0+hv0MM61iA1PRrygnUndLGn72Ke/6rTsAeWZDjI
c+R/Vd4ZUnDtcsqldexxnSin3Dx1hoJI2VN3iWS60OQZAJJ8Y0qb/2IeCSIlW4JA
RzzrYVoUC9pZ9h/OOvAsv/hwyguG3mf9+OuPfywXZAThlhCer7nV27UlwiGBIWoY
t9PEqbb8cdjkxTYB2bJKQPuJDdJpGkW6ecNQwWx9XgCbTaa0r2QpeP5chPRESwTJ
1eNWSmC5LeqlLCtc0qdcJCPezum9fCX0TDRsmX1d6BkeSgfyUfhcUmmcJQjGT7hR
Q7tGmabhMRxKXVD4oHnup0nnxm0aOUI/2E3nHbXXT0PGGKLoBNVWkhr7Zr4AEO8d
YOmShYGSQq+yPElg/Vu9oCLbLGD+S7zeZTG8/XO3Jx1cWgmptNGdd6QdfbnHf07W
JnZImAJE/sDJqOxkToAZ3i2kTs5IGgx3YvJdT1IBuJS5MZ1Eo0f/PClYCZP22+Qc
mxIqEqYTsfdDa25+L5e6fhlINEvO0jxYICLB5kdMkbz6iZ5UOr2QVPffWRqmiCZS
jDl1Rcz9+Hr5zOcsmrOk9vIfaJR6XTrmALvmrkqySyJGs/kmuA3US0rj7qpkFIAu
o6QKmILZ4zuHxNyT6sLzAamzDQLMTcnp+sBP8jLo7XWRsxW7+U757Zs+7lEbZrpK
HmQD1NWtDfgOfKAN45sBxSVGqgQf6R2Qz5nKmNId4+acVZa3qhKM8wdjI90ev5W6
vEow9O2fXNmIAQcyXWhsgHibaalTulmPCQ4/JkcfULr7BML7G8hL/i9sbcYU/ijR
a8sM442eBsP+ICXrqtzKoCmc0putXkn+hh5XkxHgs44BGCxKMTvXh5ic74P85gXq
83/Rr+v4a+cBsRg6FPz1qlHrIegsMgRe/vSRSVhWZ9hvxg1Ev01686sD/ihJTswt
UCo8bMy5Fauplh1ASJZrgeoSILIoPo1Xl/6NKCnPi+KnSWhOrtau51udSpnkBQw4
/RXArT7KE3PfyCtqRrgDHB0jZd9hG0Vr/1j8990/nwpyQUxwlzq3/aQ5kyFLqqRx
/vNyUmkQ254fFeKHZtadHCHm57o8lXuOzWwEOuyiC5Z0L2UCgs7MCDc8hK66v5ua
7YulaxcazSXOdJCkFuB19N+GecCOXQTdCWdGHk+1CM+1xPCEkaKJrKAiJqZlrWCo
D1khFvpKso4RzZqCqIR5/kINXicAjXyPQb9xALVg96U5q+94n7Hv37E29FCw/uYG
9OfxZ+oOEzzxLK4LnkbR0sN9pCJG+CfUuvj+t7EM9gyu+CV5dZO0/0xykuJI3bSO
UJx4mY7uqOjamQ+jqx12MFdactWwUiPfhmJnVTpA5WZLNz94cqFTVhSpvdxBxbs3
JFEzKr2yYj5JdY3ABTn7k/1OTSUBWmXN385j1IDKnH95ooai8VmbDWSqlQk2AZoT
jVwWOoUKi4yPyLmVMO8YjJ2/OJyoeOPOCYzM1L2lPYMARz6x1uwDZ4M/tMKXqD+k
oYrTWYAKEwSsvj5kGgWH1zMOYCnvV/yqR7DiNYvWPNZbMXXxXZQ6mfTPg9x1aM3f
FqYqoP64HiD7VoVzNuvEIS4cEMKfnXIKlrWzskUn7L6oQeCRGbYZC4VO5N4pg7cY
7NMByQaSIobumxY5t6s0FGFL25iGS5fz+CvMsSN1+Fx2RdsmC0VEBWEra1+W3bg9
qAXhq0k7zq+4XgTZ3hgzKpImxuSpPDCGWHCl5ThCTWjKL2WrtpPc4ogsazZtamIt
oftE6/T51fdPc269Qst2+SUV6BQMSlwqDTwvql8FqIsC168Ftl5Ss+yIfKGHEoVj
B7MmT1gxJsuGDHxC8HfjCY3PmLFUoIgP28nc7K/gbA7jXRvoiJnv1KmHMCqEC3RH
XVK2TuMZgfIigGmo0+74xE1D9vKJxR4Hzw+wuCBYbrKQComX8txblEshic5wxwM1
QVpt9iNT4jkzB5IRfK80BtewcuKc87e2dq+spKNxpszSYrXZZXmCpKe2uHK3aTJd
lwtfgiD3KgPzB9naYvqi7JAmVRUNBlWjvzrr80W6/xusI0ML5yAyUwohKGEkPQV8
9pJOKdPy6j5+BOLBv9vCHMyGRZauzS2GOQfB152I8aaTK4a93WtysikUlpAa1lhm
lHLwlJ5FX72ExHacbejyIS0sIEXvXEqn0/SFe614tJeBeKHnQWRYT7IcMvlEXFf3
fVnuv9zY+r+0gteMWqNRXdTP/p0dU0jO1wD4jaVSDPC+fqZysl2FtmSQcwi15+/5
4/TwQSGHbAZn+n/VZa+53i/tleAIRNEAnnjQX1LxcdIQEL+NvdY432nExTZMFg0L
8IZs/D3k2GrfclA/NIi9xBotgarE4bEOpoWzWXBv+svqeolOium4txNYzAH5irbx
uKgfSAwrmyku8pwZHp17fsNJG8iFuu5bI3/C6ZRajqDL+vEopXASX2HxjP0eIYIl
8Mk/4YvK+eRdgwaHJ8hGhjw/2wOuev4bYMZJcWnl3uPBV1j5HjXM5L/1UUX5Jh72
3RWTavFA7lA73eQEdZGMig4yE2Dp688s8rqZGVGeGNdz9k4vB1OBa1eqFiIvVTR2
9mP+9mKVqUdutKKDuKe3S6C00PThACCzuSP37booDU/jil3gf7McL1XQif56gcCN
dk1W8tWrHD/x4yF85PvPkPZqma/A9L6EKZ4tqG7jv1C7+fc+DqamfNWL9K/5c3lN
d1Om6QL2e73rgRfC4RMqTQQFmZ7vk5okk68J/qCoz2bupupmQCaUVo+9HGQMx0ZI
N+ZK0VibsFoaKlt8hWQVGYd3ZwHRrvzLrVWwS/LQGiOtVxIZ2kAXW130JRBwRA3C
xI2qAWzSI0zJb5dE6RLiVwXrglUJKE7ZYb1VXkJUH7Ipxatk6GqNLZpmjJyT7IWt
nBdegdBC0OKbWS4nuibvpJI1HFYOx5MrZg5lFEmMyutsdwMSKOAdGmWxCJmaMVow
Nmf4HbWFCLsFWLlclxTQMYKviGPCy0Nb6agZ9rGFsxbiHWKSn/M6Z6xjU+3WdZK8
yGZJIN7dCkN3512MKOgrLEqdZZYUPf6Lti41o9tCOqzj3/pLvh8oYhl7cfG0vq29
nD+5sSLVmfRzEmJbUB9hQtdrm+xwVtWz7Gk7X45ib63Ujce7dUVDgWDT6+VFp1WX
2hkEevCv+aLbZB31Kj9ZtkoF4vRtOm60zCEh3cPRj/mVBYwNT1mPw6EeLs3prgl8
/Bw5BmlPJcBwFiPeESIGWBw14a+GS+JwUBtPNLVpP14uoi7U+eQEnGeur3vbcglz
4HcNJLc4nr/8QsIICWERu8Nvek6g5BHQG3F5xiPx4FzbEtEXNfJ4PVTSw1/1im7R
379pa5Dob5zVhPi8EibkvqT+36OizDrcAnqxpeTViL5ziqqu1Jpja4r3G7w8/LpA
4kV1g/noZtbDj4zxZ3KUaPqOreLWu4L/bTV74QgLaRrcH86/fQnz97yCA0giRj5N
TJ7J7M75TMJJSEWA/p02maz/DlDF43RjpnSVWujMaQqIocpxh9IBD2HEmrlS78xX
ddesVqmsnuEvrG+iXK6cTQGPCuQYuU+peRbv1hZrdG5V/XLauviz2sPUmWbE+6hf
0XQYCV5zZhBlGMGLpTyws9pF8SjW5fp7i3ZGlqehVv4ir3d0AcPkJ3EJHht07Hdk
VNb1OCVu50hYK3fpU74vUJrwOzD31DVZ5RKRwXA0fzDvWWB2rlSMIHlORI/yUOpo
UrENuroyQKox8br26qgmb2/ER7gKbWPiz3D569O3+pBGQeDds4ycGvRiaEDi5GhM
8fNE2UYCAUaHP5zbiegKHt/0eejQ/zx/CkbyMritjQtVLAR1NJ/XpnOSh9L+MLgk
SsbxkFRfnSFUcJ8qCc7G1y+5ROBTYvzwtXHkfywEJr2goFIA1jEpupuFoXfsejZ0
UmE6ZJVJiPnrmPPqGccOubjDWisofsn+QRmaaprWfM/4FdfQb/7rxAGqL/iQunFw
/FU98+pt/jctK9p5p27VgjE1XX2NhgLkvoNQE8rAyW/JtOFDO8HMUK5EX5BE+4cc
GbPBhA9StUOkRIy4J+KS+3MfcoxJuu/AXgd9ZGVR3fN7jwHvYK85c2N1qI5aNqJ9
Hc65d+jOIqCg3W+TvieFvBaXo7yMcRKLSNfELrQqSkraZ+/bBcSiaH5SUUHm8h55
e1ayCp9HTqPRiwsuRJD0GR0RVrZmskRmKdjz22NFZDsMGU53t/E4Vh90FF0tOZjD
b5kbcH6hMMZtdaf4LJ/Pc6+G+ISY3z1nok3RIerPqclGU3Tzc4D4hMzDNbTBFflH
dU1Z+ROy0eISqgLfsDYi3aCxBwn6a/LFNbyMPaBqBuLwoQ9reRa9+XXr0bvZepea
7fCgbaNC4TAAnkOy+VvQ58BF3cf1+lseTd4e6BpBKcfKSwP3DFDALF5f2v2JwQ0S
LpyDPll1TvEK4L4bE2cRTvVzvA7xpoNi8Lxb06hRDXYIEg2o6K86Des6aZm26zP6
EmDLOUbpbqDsJpHvDXrf7UN3NQ9qC3xQpMtGgsja4q3xYaxZ8Mc266jX6cg2rpxa
C0DfJrITtwcEloGLGsPKPYrG+5oVnatWY1+38P9audvDV2V0eeramDuWUFOPF7wB
ubGXQ9tLW/KtrNsExwPCe5yESxNnckIHnHMJ4PWXAN2IcwxpmHKGrH3b+OUpMNGX
wNFrAu1YMMn8lxsZ303ZI27Cdo/FIIn8+Urb9bxBBYRebAKe/9w8Hpq3FliGhFno
CZrMMKrQ2CN+co+rEQ6aeeayAWlhwNKDsHoZZdE/GvS/IvTaloGnbnqCYACrbm/6
wFD/8/MTY8dgmp47TdFSTDSiB4sEhaUsNuy31tYWmPfffByS2OK1MaxYwI/VSu1k
LvvpDzScz3p/slFtq/vlt7WcRlX6VMbLJcjPZ+4WlCNd4adYZokWZh4PqsLS6XKj
bRVqNISng0oT+Ks849NLI9KiIDwT8VrHWqcHolfHJLvDrt3uSVhRQcj7gMsDtW/6
qBtQ0WBqP/HK5Ry12dkgpAVq+nVkk91Xm4XSyWICF/cA3PgVU+UITrdBaJNeoZeT
qmSSU5w34Ygcw62tJb4w2pU7M0hkHkLLc1nbTUuG8hPXdukGDdRglHhMaN0vUX2x
muCiRWXuMmskN9XBOJve8e0E0zXujxODnyUna3ZRLKNB1Y/BU6NH8w3tfFcQHIRU
cAQTOA0MvxDWz1zAA6VqWb0KgRudkY6PtcLj52SD7jfj+H0l2uHPnrDH1xavKCxd
PDi+OUt1QuN3cC5+iRzWXXv8u1WDPEUdmJFKqcK5plZ+nbbN0W4cMsN4kwLdHIIm
zZLouQk2E8FQzcC6gLZsvLX6hp0ULeWEmDs3tia8f6C1HLxBLR3MtbI4B/YJmyxO
d9akmd31mAG77Qv0VkzGH4Jsp/hkfc8Lt012YLaITqjy0Qn0VMuajcO9ss4DNybe
LY9siZFQvosI0kUgtD4hP9ZA9M6mZFd2z0zONhrSP4p++WV3vMXfz2GVNU2E7OcA
ooK97N7xF2meprPjI+djERyaBHEiculTtfnvtlJZvqBhwhHQxUk7brzHizfprs7C
/Nt24PhiTEpc9Lk8/H9lMojZfgeGn4Vo0uIgkTla/6cRKr37S01CsXNoHUYq4HLX
SWaxd+Wiuj/u/xH9eml2yfw3aTRPsiOuy2zJ8992dwtrGASwPdIBB7TKwYX8UXZA
/rBQqwDMDght8x9IlxPEXGlcNiLwwCUAb0fYsjWwkY0ZqM5xyl9G24KLGh+wOls0
VuF3o4lhc2WiLj9q1p9cbYlcByEI75+W76V1HgxOSXjjOR1zJ9kwFIjM3TL30vNo
hF4AtZbg4SvI9OYnrZmKKvTFsHkvAfExsGn4A5Agm254NVeICotAQtWJZFtDlpmV
xqYreBSg1NdTbIsYvdLuMIyjGnAXqjuZOvyAKBmMCfRoxgFT74/ANyHeQj44AWMZ
oHgwPK53QlE0cFns8nePyxyCnmZKmtR9YNvO9QlO3FME0HBpY63raeylVwe5MC17
riGPNBbeqOLO6e1ADbzx1YxVreWMJyvAqXk0/JxjzcJmTlY5IHq000P8oCFYaVY6
r/FDRFKXMw2fB7b8Ajz8M4Fa4Z3BdJSEwSavvKz3MBXltMaU0J/tM1+OiMa1xLIg
tJAMrjtTFgKlw2YPc7U/mP8k3CFSbY9Tyz58iLRbFxeZCbX9XRhYIOR9lif5x07+
ZMrtmLtvZXOWrvd9qEKggK2AxqhSTgcpr9grFUnwgzbSMfQl7WBXs0PHxxPkne4V
33DeXrI8Z62VPkNg/4L27EwgfYMJRikXOMz/YJoxGRLehTF9koyqcEp4ONbVd3n+
iK9r8g8qGsvy5vhZKoKC8Xlr11QWUK8+P9fiVkL9/Ld1jGvbmtN8u+E5UyKqnFD+
ssYjLGZihKxrsb7+odjEeJWsmLS+H4bSWl9I2bmRXXFuTN6264OEhXivxGbpbKVL
CydXIe3GqcwuyJo6cyTs32G8tD7yysx3cRmDtaSKb9TXr+4Vfawdt7L/w8UyUlGl
Bt5xxYYxejxmsh49cF7wyto8vAewE6V4l5BRRcB0VJAXKcbhsrVURInm/7yub0Sn
Ho/H1B0aV8H3knyTHQ0hIJhT2r2agYO6W99p5f/5tQsQ5yA9o/N6ex8+ppaoPe8D
FUt8N6AwdY1DdPdx4MY+A35UPanDtvQfiAXwIahnbsPNowOIcmq7aAlrDOtqtUxD
JZ2vkREgJEr2/Fpr1k1LdPDlI3s5mWmC2HpB5M/GqxqSq0hosokkeKJRlqQCK/2H
tcNXu0ecAT64xVYyXm6N7bR3dw0B8I4Mk/dFMUg2UviBpU6NerjQAZyYKYmWKl21
8NisQvQM6DOphiYcaRXnC9dFVwxGvFSaFFFPgrJAqRjUDA67Zh1YiGPUKf0eKd6k
50uQ3p2jg75fBbTFjhXCPh1iU2E2KOJM9NIxjHsJYkZTdl+kTWPMJyUseH34Ca9U
MJc3TUHm+hRN1VWWV/O7ZzGenwGqvNK6ghL2E/qqIupZvxW2yXMXE/wZyKPJMwfW
PFy62nWOPhRv4IKy9U3uISQ6A9wnUD2QFfu1q51UYWwifoeRtw1RLKPxUfR9m9jC
l9mRAvBQ1PIG80r/phxdpqCvHx1y8ah74HoHYby7S+FK8JmSYLd36c6oQJ7MnHph
IoKVlbAiNilXJxb0XhI3ki94AYTSs5jQo7k/7U4aiKitH/oyC2Ds+MCZHxIIIsY0
MnZyRDH8trQiI1sjb84QqxUE3Nd9l8vNUnApci8F/7VgzcxSk5Ms7G51W9S2UgdQ
e9LEiVh+LH0k9H+xbkRmTTtuGBeDzgQ8Yd03ChCRepFRCTGgMT/RQkl0VXA9KhNp
Pz6nOpJ1G8fLTB/NTua+ls4dAW7SKSZVmtsivDa3gQjviapg/+SHHu/JPFUNVsuC
gqWtlshoEEH1zv4yIaj02fl01uwUDnW9K0ZuXzM/kuzSabIO0FjtJ43aUK0k6qlB
srhSYfQGjShwDD75xnfNRfj2vH/0es/9kjLSSW+BO1GKRf0duN0xqugQphaPlmSK
tv3frxXJ3PdRJ/UfBCR8XMfvi1ZnRlix64CHfvIMOP8WeLsMPgVDtousjgA4XRUn
MkDQE5cB/iHQCu9uQGC7hFX0BGRxzoBmfAsPWrKFrL2WkGdZZHGNXK2oW0Vxleb7
3e1dEXombwvYX9DSMmkTXr+VzbzCshlQKIRYylCH/Y4Hsqo47KFyF7JRCzO+1+LK
2aO8OS/jgbtO1KgvM05Z0i7gRTP/HD8zxC4jK3G7NQQRXioWOJ29ov4flV7ht9s/
wCoV298+zhyZnVirZv+9w4clZabfzaZhrrMjiOivNMnCvIhdPXjnrzw3J+PD1blE
Bc0o6KZ4uvzL7UqBF/XYPFPkAHg0rngBh8xs9o/nwQmvtycdmgFG/R1r2rxYkLPB
OwJapAfEHm0Y8UBgPAvcgiS9xWNi+ZjozlLkDQt3dVb8cppLMbrxLVhNncz93lE1
WjsUA9mm1ujXcBBIh7AhYe6JcoIqZdLmV//6xUesQ6w/0BPNNlHEsG0X1rIhyuRf
OVrYFKPyfyHKwaqkRlFoUM5jEcJo8/FjKFNa5Qo+1D1ekprgqm26obVPUiEZS4Kc
YFjoqxIp2jYf+Z2Wn9DU/V4c3NWmHEBGzW/3/QpZDUvzuIPANX9gDOiH0SWmYz72
nepZ1IKjFeO7OJAFy36Y8tc1NJPlw46S8y+uGIR/N2upQgkuuXhBY2S7gV3rLlFg
P0DeJ9ZGg++WJXVRxyg/NotuJvp2Dy2B5G05B2R81Fg5sYJqjLgZNeVfPjj7QP6y
6liFUlA/yaLGg4U9ithjQ3NYchXDuRge/o24cMR+3WMkYi2gwq3haeTZdHXpTk1x
kQ6UH/aUJ0Hs8GbJT4bVNxDD2nBn7yZkLBzKHCcPFg96XEdt7qclaTENmoScrOJF
EvUU5zLcdpM3j8xoFdLwMAfVuhVIEDKUEF2QNELOoTInvHUZ9ZCirReSd//A1x0D
3MH2xTbl6+QsFYUkKM0GFJGXHrT3P9FuFYs/xFcgkxZHWA/aBY9DAavivhVdPNmE
SkSMsgx4SdF+mGRmf0mfwXNeRnrKCU91Ttg1yewrX/5rPSZxuDgfHW5FhJBfHcSR
B3nu6dz2gHqXZ0h4KDggue2g0aBEXs3YlywGFDaRj1nztmWhzA88FFOwRcLFVfo7
qUTpp8hDDDCGAXfXL3kQHOoSVQZPoUgTx+b+O171tLEs/dYT1VEX32iUhAbwu2dl
nXFczxtHXUYR1zwBFTmLtCEKx3k/2Nhzrw+ZnGUJMtKhTl13Vb9trWW6u+wrvKlO
vMZbrwhVfaUcCKxwXWHd/QIYmo2gk+Qx7gU0PUmWxjnebTlXsLewk8/qH9eoSDCV
SCKcLr1tmrk1h3f/7/TJdSKP5jtctxgWoeNVx09l+skk+/mkf93GeogFRsIcDRrn
5iXrAhs1Pz7WoSQF/mC0ddPSupZvycPuPsFb4zXM+0US+rWoslpGsQ03Q3OdHwpX
bjpL7GMcrqs310YVwSeaj+bUlNZN4eEXGXtX/Ev6GcZI8n1sCZP0noB0adSoy+cr
hWBjN1jGVjCkfNFwMRrFChJ+abCuDICGCdPKoVCtwCiHMZg+B/BVPkwkatcSZpHF
OrYIfcsinMUEUNzNviwoZ21U4W//Yid25Qw7gAC4h+6XFlU5gohY18Ikqtf54qJL
Ux5QrWtxjttm4eSfHowoGeFw9lzRU1FzfWoKhFYsDhqhzfqVT1CMZNAursk05LwJ
RumGWNJNIXPtKRqlsQKnVlL8Sk8qWXU1m2If/cJ+IA6SI9YoE2FkPMYffqexARIY
PfyqCDHkXq7dsCq/l3qotWwLVsbWO1FRigFHetdAji/+k3j6mMVIftrxDGzDC8F0
pYsnw7l012JQXPNXAS6ThFNMyrIAalgeJmOQ9+XVBwiiADoOh/kA+HkDAKutKX5j
bWAzc+0ozsS4ipN+2xbnKgMP4kR5a9ViWBgdnpYpxtiIlM+Ki6p4Sf34pSnRp0yl
5htNMbHJ6g64FZILeUh4Y+OW/++4xFehy/2W/FkURCxN8BD4nJff+xU5pqLN4sv7
wLYALDYNU83lgL45Y3CPplcuIS42clZr/cvtpm6V2Qnjl3FOSj/lPEkUSCV93wfi
OhAZ/HWgmzS+CqOIOtltonvYwH9GEBMYqvkll+z1pFwQDS1LUTUUNAPNBYEH7WCZ
DRmufVnagxL4awpbBo6a00bY73ZTSLZGUFJ3H99Ogu8BW20u5XuoByETp4gasq5x
rsIjCJzRuZPCTByKXgIKyIeXLxmWHXgKFC7on+XAdztiS7AVEYK0bF+m/cznthQx
RlemRwnG0JhPepmgKfe4Y1Xk8aEySN3mcwjNFFxR9U7hh4uOsN+sJdcz0EVhDpMw
2fZWjZqLaXhPx+OJYAf3BbXakjyvX+XPGGI45k5p/oI5fPo8y4WwWFHo97cTvetx
yx7wjZ1xkPEMbyAW38+kWdc/H/LauhpEP3rfx+7OmcW/k0HJLDbEb+RfKQQzbMdW
BX3TaMq2x1aMMiivGrpWnu5WzllvnlHWC7EwnKRqC6ED9iom0opUdrRqklO4lAwd
m5uoqkc7Xd83rqBNtoDkMqkG6/po/sfZKcCVWruJInFOphuJyS4RF6L8YM+pVXHL
6yCw83HhT3Phjn7XroWZAZzLoaKHLymvbHQV/GnQlERccqIdSXMVn+4NJ4qA+wfc
q/Hru2pwCvtaTnM2s4prmbkn05rwY+6EqmCHLlYn0WXpCLgTmSDpJG+H315o59qy
Habb3cy7pChZENmjGq3/GxRHJfc7mnrOWny59mbKsyb/Nc0es1gDLy5x4Y4/eKDV
Rq9/KTOOZGs7uSZOaW/psF/KK9a3OVC4vSooxgIkNvf/u8+0vJ6SZwWK9Ime70ks
DWq45BS7kEgIcLeJ19ds7uybiossqGmfwmVZCRxvmR+wol7Y18g5sU4+gJbuJe05
eWoCBaQKCdwEfFL/6vThj8SxSFvS/pNaDR11aqCfuSk3Z2RewGZCWtp1i5qG8fja
TFGB9O8p2svFT96BFKeymVERRdRJU9ZWJjaFlEaJJ9tRL8dIQStz1NpYp0pEk/ia
2GwIhbLOLeC9aqwJM/Yjt3DRphKs+4lLP3T2Abmg9Z2bJMiLixHy9n3v8zzIgW7G
Alp/B11JFns9YeGKnoEt0HY9SWrFOH7QPKMhkshexb60jwsuPt/CoJkWKt7Vudin
q3Cl5i6j4FTBGCZuUnQ852NN8BZ9W242CMOdINiiPfOlT99/x1HzoHoc/ahdg9Uh
SjSjq2zL2i3KnrTc6Ask4bpiLkVoyIsmC1YQ/FYYGdd7o8nqyjR3DTAQRjjH9xlz
xQB3k1BCcWCd5arKQhhxLBO/ogv+QNza3veTagJymHnWZYAvX7yJi2R70atam0UD
orUmSMEx72oiB0j9Vuhnlx1CPozd0ecpC0Bp34IOu/NAKM1hJAthjy2CzaAXaRFT
C4HW29flyAaVIt826dRFJRPkpswQJT+FeCQUbaiwhjMWNdOYghh8HeRGwe3iv1WK
MRapjnpD/YM2XeYw7F3ofHKBXTkazVupsgE5oN/ascr6kuIPkwMdTHcoWX32scci
CpCh++sjToafiXfIuc8GojYWX4yCS6VNtaFjSqku25dJ7Y+hwx/rHZmk4irkSb0o
VIg8PenfqUHZrwlu+jIBMARBhwGgkK7rwuAKdIBOC0g1Zmpp5OW9SHnzkNCF5PJj
U4vheSKu7q2OmnSULqHNlgy4EDxMUz+cfXZCqAjNVEJFxM0XdukEY0BQhaskrlQN
IJyes5VxHEFUpZduHSeyQf3OSu98zA9Kh3IVTQX7aIo+BPwAdcnSptmv07fTbzWd
HTdruJP9Tgoirpl9Mx2JoKRpiQoTbEzDDPGTEgj+JlZFw2IBjLMiKxcR1a5kUn+s
ZPFDGGpww6heRlLztfsNLUXnsSH1aXrtAQhsa6UyWISGgEdm3XSag+ckOmZkljH5
wRRCE9PGmnAjOHW9tRweFI1RAhJfcOTegLKjYLqakijqdceUcjeOM91gJ3LzDg6R
fXNJydsp/BuPuixxOy7y0PSaD6ajEkqUjCmWwlb3Fr7j8XR2q5CFqaWx2mMEUzis
1M41FOYoLPYJ/kwnc/wyHEvpvUsZKwP/mTClT5ThSegOdkni6jNUDGBjvdmVNmOw
jQ2IdVoIUPDAKjmyDC6MsUYlOTaJRWig5sqYaYTrqbrTYzf9jwAIVoXkITZda+0T
idWF+SCmzv6fiF34qU4x1HDXYJRDhJ4e14RJbuoXu787CHMaYMiClAgns/BRSAKx
mQICrzSk6Uzpd2GaIqrzb/mKpzP3qdqo+67AnyatMUXF9Jou8QmXETJyZrQFKaeA
dbno2hdLtbLWzNfPlkA7moz6Q6B+PeSbdWO4+h690E4rB27Iu+xXHL46K5mzlXCu
+CRNRL0qrIZrZXw3C+a/yJKMSrTM1VSx80JuGXUweKQFmCHMZTr0Frs60smLDtKF
QPIhp3U1bmZj2ut5YFk+exa3umhK8HZAYCM0Suopb9On0rZynOUyjPKmWi/SQPE7
dkJKnolYEIm9CkH19zBBVcJfXNb40jo1bU4toZJrAztkonVN6SnGkw2HQv3NgU4U
BQej47v1Kq13EZ5qnyMQnbgCm29vvohoGSeInFx9KlMSvjkxL6AeMTx4ux31LWgF
U7r11J25+TE1HOQgeTsTv/G95uwFtBx9hb0qXSt7b5QJ5z45hHwcUmIRdbGsQeZr
iiDqUPoAqN/zs1Jh1mNxsNt4/L7cRy15SahwLOC7kWMm3ayoCeqUR1zue5HUnfvL
DqIKG3Ny152KkX0abaoT2btY1xCbJZNDzfTt89ikhDm5bhJZX++XX6eUwhYS2P/A
DcTnw4QvpgrTe+VlAKL6sUooszX8akAJcUW8qT53Jj+nuJGDZuAm+M9wIHVXB7Qs
ZIvF1zNLPpjkuzLHgG9RvwsIlpB7tUkU/JxcZ7o2oCR4mwg0yapznCrpK/vSKFG3
YihlEkjqisQSitXRifE+vq+LxXtULWlDxqivAiIKKlDwOQ8XaO3EHLksS+GbecLM
sq7CWRacjNgg28EIw8N5gEdIPziZKQ0i6k7aL9Wgv+kUhchygKB2m0bOGc0HyQi4
vYsod/YOQxBP+z8aGXUKm98es1p6Z8oRp0s6mwviLAKzlEzhpcEGYsA56RVc6+4V
xrv44bgah6MeMpmzOEPITeZFRvdjZQECpOY2Y0s20NM7rIujjuPyc0pJywU4jaTQ
bNVU7/Hl1EEY2OcO+tD2ha2kSWTnLjzcp6l+P3nj3IoFP2IFIMDndSGjc8H+7l7x
5na2u4ronhXt5nehTDQuseU2QyMkdI7F8Io39aJsLVQ1PPrSrtxgpcJKeSkplMKj
3T4z6EGB+wKSsWh8gc7u2X2Boa83f4wfpi4mEuzHgSIUj1wUGVneQWDVJj4xciiT
f5gLqM3jyLk9w0+4i7FEivXDuWKIoGqpWrx+rdTz6iJb/NPvdCVAGMroCAXQUQ3M
mrZu1o52cbILSRkBYYNyqVHQ/Y732rJMksT65fu74DbJICKooxn+953lsEKP3TcT
CZf4v2yIk/KXpZzC+WWsL3Bxn/cKw4xIrABq3Sb0+lQaFMtVbyR53y1bFkKVzaeY
FbhiNUGAMmVAMzVIdmsnA+8n/3NG1npYqZWmcw0J8ZUATsHNPnWIs5iEUaagPyhG
0eWhJv6WkhVtBqNW/UFh1/wtFIilpjOdgSaKLFfnESRspy1E+V83d06O1squEjOS
8JBmpbXhW34tajj2eRzj201TbxyQ1H6thEwvq4AbZMtepc13H+lYqEmdrNONV3RA
e4E0Hbp9rvCG9ScD4deeOMS7JkY9LduL0PSvhdr1he3rwP0+mt978azSYOjw/nwT
NpVBRpaAPZ8ct9LQc140kIpDaockhvPAR6ydFhsv8f10elRTODNYy8FNHFnxRnky
7pTpcxKXPbYKi1Vxrrd2pvYOT0kQpifuoOaG19wL/3Aq91yVnlxIa+j3mCJdTe3F
3YTcd5uw5GxSn0NIrQzCUSkJ39qjc0qQxEiZwODHnEJWHN0Cny1iRlex/qqgXKuk
gNSiW6PJFoVsTDPedCiLKlSpfJ2SHKkzpjy0MssIHFfw3KFeWSL9pSkupqfOQG77
PKUufZPNuYsjaK1rapPH1DgzyY6JBQSgDV3TubxMI407l2DbF5a97aF4ykvJyGdV
wMi1BoWsMdu1p53kEFwRpgwfjBhh3jwJzYV14rm3Cgr0lKer63yREDJdhD3Lp/sh
GuMNJgIBrULNCG8TVsl51NQzzT0LpUgMCUF7wfl2CYIQ6VUJtjhi2X3HgshgraAc
MCzP3Ky5DnDzL4L+vQD4Q8om6w3dLOlcnvn253BUE285veHs0m47shaSzWaJobox
QajbiaOZzee9QytEJfCikN1Pzc6rZqMlno8VAoPSXWfFPvTUVHfpUrTiSfxAuyii
rGfF26ylV/Htm18w/ePZmlHZoLbdEsfKlLrDC8v7D4AxOYRuJov77mMGmnlxX+6M
MDb6yBTMEhc3uMpSklFRYMiOuZlXbzXnZnY+F2QgRsrcZo/CMh1JXXF827e1Tj3m
tmJSOKzDptZUQABCCy4Yi61iBk4RsrAU8LllGXGyig5VKfEDHfMZBtpA0YOzig9F
otv4e2LVlKJDsHo9+YWvmD/5rB5VCB6tnrggs1WU3sYh+KjxlCTihp7N+HBgjG6/
9oVZ4hmf4teLxCJhtXPGA5gIHXHzKV69dU91PlSZJqFEWhpJdGFOJRNIhcbO47t5
IF1L0tfNB0ApMkyhWFWmZ4E14e3pSN3sdl2jxCayM3jxRAuWZx8VFKAyacGDqLRD
+s6VVqlrJM8kxc2fg/ZlKYdJe6cu0a4Rjl6HwcCvSw1xjHYTcXQ8nJy0lGv6AIB1
kozpOhG+OTO/hGQcdoy4rgow1AhCdxqfnKWduDukwKQGq6x9bFnpMBQpeQKIUy/A
aqzHy+wEgIArcE/+zPB4IBn98buMPsmRQEBFxfRK1PMiY/P05d5RGio1XDfXiYu2
QnFs/QUkAECAWqFhFCofHZagbT5N9KOX0eEva4QCCo/QWNeEnM/8aSn5EPGjEqM4
s+YzYwUjZfFjakbimjbXwYHlnJcvlHQSYOwhG8PcWL5Bfcwdn2v5dHO9dDMf7M+F
7atdxnFOUz5e3hQiArL5RwWrqLyJtbejgUMMDQqB8h8oY/5Ht5Sr3VTzy3ir74we
BXlJtyBUbULAdKmOQf1IG7aW0n+L4TVRKN7H2PJiHoBo9g7XF2WTtrbXPZamONws
8L3Eo/bAg+RappKQ8FBCrv6hGWapwgiA1UzJWK9eZS//8is2+p6DR40qyS6jXN3i
MeDG5nvz+v1xYIr5vYdFMAXryHsDLFiPZaOFBAHTwyeuSQWK8yTnP8n99o2oA+r5
yxenoDjyhbHjHhhbYTM8dxNF/E+R631stqlMOINQHuWuoWS3Yu5yGNKN9RpzjZEQ
CEYGLUsLYDWg7qVJtNw9wMtqczgnswOZ60rwnEUE0IOHs2EUErl5BPtF1btUl/nm
/VhR1KtQw6tW8Hf4ohU3eu6S1yS1+A03lGsit/8HmvTRy8LrHy99Hhd+so4ok3t9
qg+BpNxAgW4r2HkWemMEmJz4PDp2rbNHab6YRPIvArRIKSUwoQ/uI79kgphzlYG8
GcctNzZzSNucXYFCKrNPxIopv34pm0giOOo9okIP7s6EV/4AoCoCwyE9jNjAlQEf
4P0Dvgq4KCL06EJc28Nf5wND+zjB0y012VEEFO4xRJs3IwCJHjx8xYQD2+ZBaOkR
plm/goPxnQIvpdv6UmiVGXBkNsI83lS2L4rdV9cTxWqNYuFVLYteIMB5zbiz8tPo
akAtEsYoMyqlEQYyduNDlA3aThfOyQkKTJOu+6gP/REx1qaILvCCwyVNE9mBtUHo
tSUsRDVPDxnAugD/xHSsFlwKGze/T375qhLeBx85lEjncEmPcaRQxFauEm103UHK
jTs7HIkjxW35spkiVCvaQ7hQc+h432mgw/Cwbbqi613jPjwT2NYHfoUKUSZfcVYD
6LxM6B7MzNq3BTKWfO2h6XXy11RCoORriIN41tWPff9vdA6OCiGKsks3NpXurBEr
x7FX1+uN2p5RREZk8us9Okv9S666e5bOqBpbyC50O2ADA67DnCoXij13TLMr84pP
Q+PzlIeCUJtAcPVh575FCFo4y1ltv1Omb/LhJIIFpvhR1FWHNGHzPzKSUq0MVgs/
jX++oooDVdzSB25mE0lx1skcENOhqT0LnuBGp1reN5I9ZUaHSQrm/qT9VSrKTbiM
Ce3bjrW/qXj1KJBrjca8wXm9PR0cACisYbJ1CQEgcLV95qPI+dA+yW7kWCF10Ovi
9RECK6VNzZf0KpLdKCFt+9F3ZkA7dd50V1gFewJz6nHAMfLZCkoVHZmbKE7w+inW
URlZBgQ6ZpVf4xZFzoxqjiAYH3DiS0+FPzk0WT4nPHw9KmYyfH1AfgXULYgUrjTg
4kFcbPHmtkmWWG4gF/NtcRnSqyET2Syss20btBhcoltTxLDR4k+5hcheRPrtof6s
r7xwY1bKK1deY4j9mfxVf5kTfAQfIHm/XwyqPiRAQSMppWihxjgk7CAKiQHQ+GOy
rH0aYJGbnq7AEdRMXQjr8IqlDwInWCKg8aYGpBeY4YNe2UzDfd6flliiBhZgLe4g
f19gnBemsNT7B0i9EoZoGsKfx3t+Qf4s0zZCH5qPhHidMm4PvHfu1QAGa+4U7MqF
X2RmA5x7LoE2BzsIVMEUTGaUVSXSA6hRNL+gfszdsTJ4QCkHXH42Pk9k6pnL746r
W9Ds4LcyRB1nUl5vH46Yf+K8xeaS4+Mr1RZDJeXzq3TCI9xSU/5lKHooynqFkCdo
bjzGYWI64R/BGnS8GBo3Lhd5lwnVYYc0nKqk2ETkzHum1tEvzPykLNHuTMeIFhcD
wympq0CAiJbFzv1sblRqLMyw45vkPTYtSS5Pnyluv5YjWRd8vOZ4wtN6Ajxn63IM
4wYCRLUxg026ISCmm4P+vq+ZM43d9ZSkyAmiqJ4LYK4/gBtx9fjDXof8Vc8Qgh40
tuNOmk0UfDJC29f+hgKyg0K+FmBLiozrEi5av9xYYIQEp6UttspxJvIdunTamudS
THVBHVYRcgbWExvYLQYCW8VBWQLzojw7PHWLdMHcFpml5xmr702xMoAqElS0HOi7
TWnfm6ZP13nRj6VgdJX2d1q+9H2fKCqn3sRYlqleaoPClPSt105gBSKbOnAmUDYc
YyAl72Wgp/2WQ/Qm0KV3bUgc3YKK52XVYHvgEX972HgqHnXpXWHct64LmZUhYPB3
mytZZ+0vUEiNPp3QgII5A2Zu/i/qz4n3vWydHXCm9VDKDl9WcHvnuXRZ7lj7y5Uv
+fgjg+hF7rJfbl0sMiBblMOwJ+k7FnInOHYlyRie0ceVmMuhq+1ImzYlQH/3nnXG
jcNSQYfjIH3dBcdtup/AaddQwUFVS+jgwPAMwkA+d30RrllBL1fslVAsCQ2mjjBt
zPYRk7EOF0RCRkurXewJeOLHbuWUitn9kVE3EXs9Q+NE8WHdnB1MQ3ZquTTYAR7l
YkWazXRgOJnmunpELjOyWnj2rtr2Sd9qemctxZ/wm/U/KZVX5OBNmHmrsq7K2ni3
/0H+yzjtumkcax5KJO2MUu0sfFx6FSuSj0SMI4l6emY/X2SsNTq+ygVq9sFhJoeo
kcnNtS/eDDSOm+9l8cijwFKVGnfAmkrmCL3Ob6cnslvseyoo9knQBYBgPiKYnkPY
lKHmKy2s+z/6FDSm1fhfoO6qXpfMitjFCRN0v5HzBehZs0D30UjS4leDOvF7fB8A
mFdb0d+aNREn/q2FINxWIsbL/sFqasXHvPbEZxBs/aw1raJOQUUa1HebLtbnJfam
1nweQ5RoVaiQUI+1T1sEEbbOvNBmIAmAvg5SG7FdneAxE7lYJEQkpfrgAZxS9tTX
KUq3Ol8roCsAkFsest+wLMtCV5DD7LdF5jmqtzH0fSZNs0X8gNNY3HN2Fph/4gtC
7L/WDtJIzWbM3zmzkDEw1LXYINvupBmOqiwy4h1e5n/Zggk7wuhRUhdrUxuzo95E
cNt8euDqon3XLnF3yDrvVUvl2iy7ed1G5YVvsw/nAmu1FkYXcJp5NgPC7ESS5Cen
FnTiAgKbacJO1XzJRNKzOwrMps/1DCp45kYpw4505XJsrJWtgRSiuqD88+akBo+P
fbqHhXlywW44338kY+SYzKbmU2F2qKsm64M/Dn5xfiV+3OQC7fCdZHFDguQJm7DM
GcqrnaoEWOplmTz5t41In0kBIBahugSu9V0JSDmEdlEAWZRTOYIGGMzvf5XBXwlP
BDXU8ghtZ1QeT0MyUaRLDpSyaYA5TGzIVBI6zG8BcEsA4IsqvtAq78vyO8vbg/PA
7o1fW/HqiA57A4lBRQotpXwGSielvgzvabTpnor7UZE5ukCuU2T878kX/Pp4ULO+
6l+eFJBGcUZlTwBmnCo8dGZ4K5dOLiTSnzmpfVZ487FyW/phwEt33z9R7UXzLiCv
rsLpSdhmADFvJ+bth+YLfXckLJQPtJp7f5SNzFNNVjOvo5r49J9llXXgdm5bjcsY
xuQT2yH7loY8VaF1PUwZubsLPfrM0OErjw5THWrNX4lJVXCSJMFg1gEpyEsGMNBn
50khILP7jcEtRh6fhrIypwVMz1WSLFsr1AVoW2NmppPBDhOngtJiU452BpRSrJht
2vgXpLsv6fvwURR0K5/G1h6Jk/TpGa2Zz6oyRqZXASo8vL5RAKLHNG6a+oe/vj3W
AQl4Fkww6AAR2oO4yX74UGSigWQRQeroIl4r2C9HSYrmAAInLYVsQA6oofBUUuL5
yHVeD8phu0FWFNaEc5Eg6LQT+kxwlmo0nonoBLbqokDwiGc6uor7B0RXqNLFiy72
FBOQqJonY5FUpcOWSr3d3dFdTa+5xiBzFxh0lbi+uAvx5bYZMS95vhqNTfIqFi+4
PLyh/tHvQITrZP3x728Pj85DsGdQjCb/OTdpR2KqGNOlpmJ4oaVjixDcjEMcU0Uq
5qrIxoKOzSxhJ6q+6fw4FBNrQD+Qe0qZHeVKvVdNum3IMXaQMUz/ncuQjictCui3
T/awv0wZAZmhzTjUtSgJ70/YSCVcLoa2HJnC9WCEDOVS1iCapaZtyqPsAmmWy01O
hQ1v0bH4qtphH5RtCbaJ6As/+Qkjfcrx5mpjQzM3heydKiKcwuUK99625NFNfK7F
x9845kWwi3k+yYnGB5gXIHYtx+6EV1T70vqqFQ5sYr3IRJDdzPCGPg1vv5zVnful
zuFQoPJxkGVHz9Q3YCQ4+qBOkWlnp+ONDB6wgQhQ6bAhkd6oCZCXFsfP+Aea4fLr
dIY0KkV6f+T0Jd27nw5Aol6bfRzdJUnhIO/iG/Bwl0p4tJyHWa9RLPSD9Vbrauln
TLtwBJeOA0J7nVVDbwZmaxKTi5XxazydXdB7095UEMYEBLhGoY66dn8z7Mu2KQXL
4nRqGsgCfCrNfbFPd1f03rHlk+PpprDRXXAviF6RK+ULrLuoVr9CMiV292QdtwlA
75JfAhTe/XhvXEYT2TEj/Q23iJ7kEBZsmgPnKmjhhxLsbB6ocTo2Z8ayoEVRSvxK
8+pqOAJqCYxEsx/tjFr5pL6oN6Ui/LdL6npR1NSKeERJSTcUgvKDgPDUslrsbalU
IYOVDIGEOgGSiJdmnWcVdDX56/Z3LbN8t7Nmxw1KyOCPzZ+MM+RKlG43khh6xwa4
k6nub7gZ/1HNM8WO2jEhSE/HXX6rRR8/MCOjYsyD5X6aoBy8Se7UeOP8GjpZaNHI
vW92broO9af/DU+1t8oVBgDRsgDwgYMrIV5HAqEIgY/iFwThSZS1csYdDB5MXot9
8qWBly4bG6mYshT5KGSCb7RWY39aWpLtGLVEs6lJYGb4kN7/4EZjjbJ2e5xXMhzE
XQdapLuz9AjeOQVNzvuQzrnrn/H43UGujShX9pus+ftnVKxfAMFZnY23T6+laa1H
/mzzp9QAVdGwIfahF2lfjy29S5Zy1VnSV2i4RMih9RhthLJo1G5cDgLop/V208jd
Q3v/Ff86MeD/jKQIyT08idNgxrXI2wcmaVBvDDXBN8xN77E1sNc7M3PggIy8cVyv
DrbR8hlFSziCG3gAtiyLxDUyQLGtgEjTWwSO1RlesGk7c2rj32h6NgEhdXI91Ve8
uvweGXFMq0I4/2rtyq679LldCJJBwC9Coc0QSGPBBWek3P/CuY7qPcWFMoGY+7bD
5kcU7fXfKGzvkn/8LP6dZqDZQauyT1eVKol69Us3TmfIlf+s24Y16e5PhtnX3mOP
fiFO58xasywolNF6xAiM+XHzhmEcVIQLNIpSlePqPvT0gHobISQbfynEtZ1q1Wzj
KJg8m4ZuaVThYIe3jzW5i70J4e9Blc/gdMT6Wjjo11NDJei463WjzZbfwuorqhqD
MqR88PrOWmVJZOuhx6REMunkHdxCPBw9CrqSmSxmKqPguGBiH0TixIk5hQXBifbc
dZ9ph4/8tBGryba3O2s10BjFSXnC6c4SZUUctPnR1s7m7xCBbqG5MZ0i8KB97hR4
C0/AZIC/vc+HrByjfyOpEjr8e3Zo3aQnfwkLOgt69uBaoAKFNgu3WgH4e8lCw9G8
4gVJmeFDChEKxOAXWPXULtk8G1wFQ9Cf1QomVXwQs7ZVCEoeV872Req3mE+lkRBv
WG3WSS3lAqg+VfYVl1ZbC0by6syMWwC1pdwjNLoNj0t1y4D0ACZdsbsIJ+cahmEI
JCLa5wwZGOJmCcb2V6DXPkIK91HXi3srCCijX8k9lWThJM2/03TGBRZXJJlI5POl
Dbb8mcM0yq3bakcm04uqaNn5nTzReQKS2zW6D6k8D8fxBh835FPUVmgJAlBKnIHv
Ri1ksGOeTZDnYh9BlXuQOqUffomHFJRGel7KdqlhcyPX5YSqULIDGlIshsB/tmhE
hkmCdTfw5YHZgqDsyUcLy++SxUJCjg+ae+us4i10QEooj2xleIeGRwX8T3sd2rpw
zvzYHDWJMrQEf0zT9SjELu5EAv0UjAPpu63kKK5abqpYfj1uXKHjwZe6WfR2Ab7L
9dNeZRT0ZQLZjmOGCWTEgcxGFUAAurcJZfz9dngIrJ1CYHaREQaF5zKzuFH/ySf+
RJS1S7J+KM/yHIXSBGBJhbymg9hgKYktJ5men1oAI61llEojfNcSQTZUiTZnQrM9
6zcjVmbONFvRRS7p5zFl46HOK+2a1D7H3RixbGZwsUn8KncXBNdpKrxkcp+PIC0x
pJojvjcnDz84bWe6deUSD1ej3QVyL0+uIl+m5jsk7D1cYH7aw0nGfqBBNRUZUcS1
Xb+t+kNj3o/kDCu6FzYJXGvXIcNubChbaJl9eEHOBZW8+jg0BHI8OG+AFnH5oXLR
09uZ2f0ZCW459drFRnR6r6pLDqu2m9tXXuFkHxTqmYD+5Xu4TKC6UVr4zVb6n0dw
HKLj2xRlQBr75zUnx70J5+L/2CTlVOSyvPHv7p5NyEyd7FawEQI2Uz4UszHx2RWt
/0NTLRRLtL+BFszfYUx5h6eMLDbhL/+oYZ9HqCj5+nUtD8aqfl88F9wXYBig95xb
RbdCdEsWnXl3BH19t6YgSUVJCeZ/gM4yXhEU2k95T1+jK8xqZPzDhGf9Y5MIz4f3
zA8degsnJC35kzshyL4vGUl8lsVc3fsjbrnrHIrc1GN2lwWbf5gqfMLfaAi/0Ka8
b1WUh5mMDhKa3xUqDWMcSm9sjlR/tiPAcnE4R3d9vxC2Qf9gfQZWVYcpI1LEleOB
Xt9wlIIaPnr4NoQcPYBCH1QjXoL6IND/UicKo0SGyPdJntV7rmjC2qAWjeZxQhC0
lQw1tSwvSyrdqqvcroX2dD6OOSi8uIhLZgEX3y17imnY5IbVy2UWSHgkiCKSor+x
IdyRRy3JszpImnP6LxtenAQpNfKQpOJhFSn0R7RYgkGENEcQOpUyQZ3UenYT23QS
/GS4fcswFjp83SIQ0ppdZHWxdb0RX6Q3Vnge7aAPRkmICxaSUbV6BiSfw2C7iItr
W8hJyy3Sak/8Gx0J6Y1F95eqvWf50EXQ08g+AfSqzumoNrsV9LvlyXAeb0UtVqaQ
vVkP/z5Heu0nRxUbx7PwkFvekB9wWEabtGmtJlmotYDk8IHttaKJVYxlmad9t+PP
QzQCFX793zJ0uGyKTVTf3vROrXyqR3JEb81pg9wNkuYFJ720C0FLIiA1P5VRTYOL
Oh6d8aXxH0QCmRhKE6lvU69vLbTGK3u04TjCewOr6tM6FOkmAbWp83DBoV9p3KFm
lZH+gKfC90yt4nX1mBtNP4gyl/58y2yTyFAAuxcn23u6l9dx75B7Qyg6MG5sM+TR
Uo+dsYLc2X03OzmrfAsbrzfRvfKPlTaFxJiQwolaBwdjD4NzNS++TqWAl7mV2wFH
6hh1VV6ayeA/fPFrXvLsFdL9H05znhfjcZ08YXbRW6z0knd8rgNew8A+GQtUx6hJ
WTKeGhrhsKApxLpJG7V1zXOD3zri3oQz4OQ8hln3PmLMbTWRnvbbrNKwBAkATffh
Zj4I5cMpDYmIh6uxIWA1dqvh1jfREyXLLwfBXvaMDNFBvmlOwTU0JrMSVg+Orcyn
HXuVHnI29kIkCYe/z2RRE6uGGEfqgAxpP0eT/fxkpnUe5HgmTBxWNwGsmttpLKjq
7XA/bmHkbpmbIR9MYQnJsgif0orz2+OZqDbSn45FuGWPo7KB3EsD2VqRL/H3YE2Y
1DO1+KgnR2VE+ac5pE+Syf3KDa0WHuAIuPm6VWFktklH/4KwTPlPbtymloFj3e0Y
kjY1q+lZpfOp5j0kfbBxRfaRibJ6GZBvIm4ej88wn3kOn3lpotBDzJCL/dvNC9X6
4HjKs228mVFy3I/QQtthfAgLPvjrRatGusAq5AolDtgqrA9udQacfpteg0gOVk1I
vrmcJi293hX1CrPO997JvE52Iu8JSxxm8WDxJ0w/XjFYFNwGwExRcgKhhRfdi5Vi
JWlnOAts7BBDqfkngAANNB/X1jNumB3Mb6CaK/1d0Ii1tRfWs3yg+jAlzObKqV8j
dfwxZJSdSniHIrVB3ALmiXZDg6TZIhfTtwwvxBZMdwsVLFAlZM0KRbfDbHTqMHcL
gNgNRVbFWGWMuR43YslRqnDBOOWnOPXVikeZaRJJIC0YaO0yHvmNYKXytupQoccY
I+AKgiSZOQzjzloqsfnTL/IcBTXOgrGfWA6fdDBQoFuSEu29BEUHeFMPkhiL8wpP
VpoBrZw1qq1YRLP6dsnThDjzIiYiXN2pW2lWkEXySQ85EA6GOgVKLErG+t8tLxq0
p/yY+LYnNjTAEDLgltkUX7ODW98P++oKcZjm2cq6xG6Zv54C143ZCvvalXZ3By3I
syMln9VyWAhyoReI7H7tU9KKa0QtKN9hDcGtwiVd4e/3adJ/Va+chJmtYtn+BgGf
E1Nsqxqf81VuBCTGk1EcyQ3BleFoDLE6hpc0b1PEhWYGhNNBMDO1ItMkXw4sIXHj
UMUGJ3bJO7Iq3Dx8Cg6QntmZXzreNkl+UItwix6xv7rcDxPFIOJTCvlrTjkmiFN3
hg9wU9FwIcKhDGjWBEi6VgY/7912sH5pIOiprWHIqpMJI+s8uHsENAeOW+K1WG+D
ybG8sGBDkMQQDoycUpVfym7I7AfJcFBkTfaMrEo2v/ZPZV1Sp7GqeeTKQnuUMYCg
PVsrz/xpA3tNy99d3Fx9t6RDgvp57IpwYVKwb/nUs11Ii7urryxPQzqDh4lXntRi
eaiqJQeMS1HZdX/fkIEbfKTDW2G7FoOjN+OjfoNuioqhWwYQgi/aoUKy2Nyk+MIw
mKErfWKNQ5AASLfX5F7i5t6IFK1/VWrjZuDkEvMEfvwhwuh7exzHaeK0CFhGs88H
cnhgRmleWMr+jzbc88zHYkfWcnLY12t6+/naAgIJKWTIYrZIfrgUTI04m1MOY06i
hmEzQxWntFLAm9+b+VdGXDZ6rYiBNdKOM40+wh6MariFgVae/eAEcWEiavwfAAkt
0kCoYcOyjM2+eZ8uIy4h8sh8asN6wAivu0nFbWCJTCBkPaUGuymw5LmSZYGRgvJy
6YGx0JeNqh9if5h05w/1HRmc36DaWFOoudOQzjKmBFBKJgAvU7ighnR7ff2ty+9R
Eqvp49WMAb8ViRGFZ1tBY6zF00PeWwyPpQ+WT1/q4f5XvUiGzeJOgmthUCbL6AOj
hKU8PT0KPSZzQh7zklvUi7bUIVcI/RG5n/QoF/Dhug32iqDwgYcceQPXSQMOSMHI
xu0S8hl9Cv84t25f4WvjnIewfWvK8ZubdiHk39JcSIC3xdtcQloghBbnpgxcC97c
kydJ6VONZ+RRD74qlfmVDtO2dB9nEL5ixvBs1hKjbtH93WTZmePogyygmUKbcXGk
lxwSbC8FjHBj9Iqgs4YyT0pSobuATqYWJL3YsxY6PqGF01cH5K2IIZzSBKTizmlz
nBBiCj4p8qmMM4rslagzjchtfh+g5h9aZPxAjm/QD6sGLUTVcPXY3BpcB9bHtdcF
Wg5v987yt9yrKYUn5Xk76Vk4T5g+qGfQlFyn8fHynfVA+Zg4C7f9OSwJbm3anwmH
6Lj024kj7H/j90BYBbrr6Ri1vBweynKbGbh0JfVDNFcKfN5wBs6HmFTpfRHpEwlb
FBVGwYiOgwAqfShUk3BhUog3c2VZ8mP5opG3TaCJ4rZafx7zINNuto+YRabU7LWk
P1yx8bTGRoc1Y+5uNsLT9NQnoaZ8Lnpr4efHf3fOzhQSOc8Cg+UpRnqnrA3xOCSI
Rd5QTdE/L3d9nf1jelslqeY/xPqhs8LJ2sG5MdLYH8jvwi9T+1Rb8Tv3NQyHvomL
1MEF1NbSGmwvBioLPc4OyiGU4Ei/NI0vhLopRxFWCbFQxlp/BzbpeRXCeXS54i08
CrQQMbn9wJ+hbipONRIIkyeXxjNDma60lrbn2ZWYOA/Ou694uYlkMD/kXcEQIAXI
YY9mEYOUvxyjxSpRq+9rM3cLfXbJlMoEp7L//7ZW+yTvop40JAjfj93YhPgjXXVN
SJIOAEe/2vzVmxo0THzndwd5oqbLUmE4xarzlsoUa+Ik4mIMk6T8HXfvXpO5Haxn
HCfH3PUWVPLeaQBFoDJ/e9DWPiAC+xGY4kagjzIGtN8bgibG4xC6Xuw2x7rqvozt
aZqgArXFUDxJjcEBijmCwiysMX1sINMdqHbeV/Hib+M/FMXLivvKmAipuR/LoFqJ
cOFEhST9FO4napsJmYu5IrfSMOG1CyaWNStUtBRfFSxWOUDQrbF/AXE8xPpcwz84
Qh69zwSpLGiKKupB3os6+qSZEO9BHyUukMq9h44b1JBL4SA02z4bc5zf7+RIxxTI
nH4NEi5F8DUqZSbFri8cOVhC7Q+ydTdfp1eaqzg+rRQiZqoCMFPS+lalKRtSwsvs
4w2mUw5sO6+/6D64lk+Eq2esQd2zRJ6sEKkAbpMNZpxpTAnJnABl3Q6cyJbBS5O7
8pRbNiGJaZBTjvvbmt+4LBBi3qXO+69KHd9oOtf3imHI3psV2gYSESOrOT1KEQgX
pr7ZH5mXSlrkVTyZQp+1X5kHKok3+MLKKEzKPudyfMq+fCRGToRo4r68Umgmccfr
6rM5WsRNGYWoAizuDHi7c6hfcMePtfAu7Na8C3rTafOYFGQAhp926hSqRFirSZx8
mk29NINWBdVyDJVFu8h7Le2CQfg+DmCOkuhP+G47b9+zcI9orxLtXUd8BVWM2XIf
TtcCmHWOgAekPLgQCqF3Evky82C2R/I4e5QJpZEEGi0BZ7HrIUCyCzAgOSMss7xD
g4OaggBlW+y0bzdeiR6pV2Nm7GvzRcon0dpwjtbg5PQxvk8GZUGg8Yj0Xk12lEWz
wbwR8sYjJx6wkn0ehPfkHqeXqWAJ8FfoUEZmbhuCWlTQLmIbQwB6Fjfaf3GQl9tX
KLJzLM3jnGlF0JzqHy53FwgxTDsvfA1wVN3aMfbBXa1WEGplFHNAHlT1Zw3YZMFm
Y1V2lSBo6Qo/EQwidnUA3k7UPJeFKJ1vtJaDOHcP4PxaMuPaxogVB+F6rJ8FjCWL
KYmFMTyTV+royUq1fHhmniDd9tKEvCLQGHKR6+DZFXAaq8siys6Dj90k6p5byH1W
5V4Vcqbn46btHTJKGn9cycHgyBjcNRmoWKJvj/oqnjEavPSvvn9iG0816/Gk07IF
qwJ5dZcz3byaWW4mlskChvi3E8RsaKFpAKKoXVRLk5wbOCFW0hdBwMW7oY/m4lFO
7IPzxq8ygU6ILMB7rRipnO2/PWA/w4Px7ljTY5Fde2bO5HwVb42PwkN8tBr592Wg
JAr4g5TK99Ib9j60dVvwP6zecXH4MudAkHjvRWclWO7aCHSvjAOhquB3Crf39D5w
RdAMCNiHxkcfWo1b3nq5JCReCC2X+78Dvw3Rq533l0OehqhFxAX4deF8yF3UIzxh
fjzTVcBZMO0lf0Dhxn/zA35fhX5WcrY70b5iYuntB7zsjpQu71O1S/LTqMJFr5Nt
aKwYwLBD3HXd1wvdRBO2wryNh2L+Y04TLSaMgmVNKj13gHr+lZALNedeRlDTcR7Q
KKmVA+4UsnSG6hZlZ4WhpQBOCG6GQHs0fgY8xmn+y6aOQ4hXW0qlpsFvKHMsIfqs
D0Q1OxW5MKmKNbhMPvGcJyF6OHa9DsddcUT4L0E16g4YV9X0JjB/lqfgzc9JOH8o
XcfYC1gwT/9lXxnRM0NcJyGnC9dO+X848r+uYaO76rZ3Mw3zp3qWCEtiqP36+abC
57XbAPqTh483YrO2zHXsdV9xEZdl0aYQqjuEAzRwKyElohwJdDWFeASZzq5dOr07
ih0QJzc6eOhu7LPZw80JaIddIj5tt+iIaf55LQ9us33AwsBw4ZufJ7kA8MiTIITr
PntafFsZRuULZeNxBbkxOZAiCSFnlxVpcw8O4ptzu/1HUKlKrXjZ2YEvT410SWdh
/GjHnYHdWUl0+gANYDQrov7qAUrcVQAX8Jki0Bd57X+V9sKtt/LNVb6uP+mBOTIh
bulk8SBOfMVoiB215q3MIXN9wAzRfL0GeTgmP0YMtmdayjpsJ4Ik/yML9YXF12Ra
NwPVjc1O+7VSIonyThO8Z4szI0FGklj5s33P+dgwfXSGLmeO/HTdkCLS9zOQrNBC
4bT4kRnisIGpuAAusyUuwNvYiRZaLEmw0Z5/fxjVYviqbduTcXzIOkLi7tXKm+g9
j0YX6Q3XeBcExGfueK9eHlSOu4zV6mF+MV9cRvPa1iw5iU864CmtJ7utijtdBVIl
CPYJw7V4bnP0McMHxaaX/5TDr2+5+Ken7xfmgdvgsr/3T0MkXcIpEnfDk2k7r4yt
3U+IjQ80slMLk2Ie+iQ1pqP3vT9L+eEcprz6kou7hz4QRsOfKpKik2yMMPCeNfPB
seS8TPw8i3TxKVdjEq0XFDoV+2z+MQWogHyGzNQIeJSngIqpafSPZpZlVhCJjr4n
KUm4BYpkHnNYgf0YbPz60n3S7q0wEMB0ylmKQM74i0z/8wX1g3mf7Cz5ogFLhLc0
HpHDMc4ADZKaKdb7Okh/t8D/rlj7BYFmUYn3gTDwF/72MmY8tnbk9AX+OUUWf7jb
q4Ro0l2Le8CTbgeg+fd7KSVHqjTDauOA568Ye11enI6M9x23Slkc0dBECPEQq6G4
TL5E/epkfhHhIngR+1BoeC61wykSeZ4VbWVrJP3wZvNiNJEnEe8Y92uKYlTDJNzt
VnmFkQ3lpyicI5FUkO5oEIRo7VZKfuiMQgZd6pIa05QnGKicTC9ur2Wigm6vD9/k
ZVB2LkcFvjGxPPyCDLB4LYTXdGlTt6BS9pyOQSv8A53sVPtLBp5KM8tR951te2aO
sA3rhArKlSwUrirKpLY0sYLCDSparznr05fOmMTWxsInjZT1y5YMGE10bhAEJvlJ
e3zK7BwS4M+OHFnnYRXEnDk2yJy6afR3iBNnY92LC0rd0xJEtqIY+ooda8nogl0v
+lzatU6XZBvUr/2F5/oRgokVgbwV2digL6PH/D3CEEsiR1mtB9KftnGy1zk+Wumw
n+hMG3E3sr4xXeyojrp9R6s4gQldH9hJKmqyKZ7oqWO7ZKSlOg7HgPmkI1X4b/Pm
+Yb4eiwAt2gbXftBt/vAoG17n4plUxq5kd1hMB0HumOQjFCZCE+l9xgR551vWzro
R8VbDGjn5Eo+/hgcHUijS4T5d8OubQHW8NVkXk68NXlkauT9IVsNjxkjHUrcBZ9/
dGRwwjqggHVSc8S7e9Uqf+6uvfVH+cBAR+WyXdpsZfDCxe+TVQKS5BE7vp+uxfR8
ZZ/K3xtuIiJPhNAKf1uyJPjt/3aX27d8aOYrD5nIZJiC+QVI5vHT5JMFNdllqAyc
K4FjWfAqFhoPMv7posgVzWaPq+Ax9r0KsMN7WF6sr4urEOEuW990mgaId178/jEw
IEp0pqhVFhZNvTbxDYG6f6E1Nu+qOLPEwhMDjBGCDc/diwvyBY2Zlnny17DvW/hH
KpUx/2t+0HfILH6iJFgsLbWJ0nFS4C3Dfnwxsq/MSMOB8kPt2xwhWlRJz4YE+oAQ
yNdX5ugok4Bglusp5YXoeO3AvEGM4h8xidunGD7etgygj90dN/kzxIOn99IDFlPW
c/OD9H4wUEhuJG3gRzrSj2K9zfAHtGnC95+2yCbA/bocO+BZttJkkIuCX5zofYJe
upl7cC5NRaM0duv7xiHG1L6d7tsD1C0xdMBLKdQkTuGl28ZADKwVMrsPCgbJrfl8
KKvxCKJfamkD2elrjnByuj+sVgHnoA6QTjkaTm60GnZ3YpeKQkm3vo1IioBHxfle
T0U8mX6twD6tg8+iyDJJhRC2Zh3PZDWUAvZgrFEbfrPvbuG2ijJVa97sbKePQ+WM
NQUhzNVI00bWdk2LbCuuRH7axgtpyT5/JPVh/qJB959H6/EB3FENWG13xKiJ3OO8
B7qF0YLPac9lA3GUhMsX9yfFiKMP9SJQFiQZ5ZCZE9VhymBr0V2HNnK8wBFYKLE8
SkXTax/kbAeGCm699EN/55+F8OgWbjvKg/20lTX//sKn36vkVSFkl5ZEzM1/8f+Q
+EXngQpTjjzG1t+U1pqcWBC5JZPNEYpxeaBlllFQYPmna1UDkRFZlOPKZX50PdHy
ZtzytfavIQPHIqdJjrHhVQXTSzvm7YRv6jIh27PkUrYz1DdVm3bqVhtyupZkOfDu
QdsqOjh2B3k+Kbn3vqtgDL6qvWIiAH0lYZ7Ql23A2k/XNBTQJzTL3ZT+BJ+otRnY
PM7Fh1RdpFHyuQ+jpc4tZsDZHH3HM1AqfJMTvhYjlcfRa/9H4Cga9BRLjKK4L2rj
aS2m82FVs8o7uEFr6fgO+V1UULZ07l7CH7VefJBgkpozBIQhme0jutTAT7hMIOsx
fQFd6hqxoYWkOw0U1NVWepB3DR3NySD1Fqfu53KgTpF/Xa3uwG5UHSxzUihw7lTz
zba+kmT+bzkenour6+dGgeW5uzOsYYMODrh7Qrbf8ZCdNdrcHMN9mJgR1wTRHQbb
4aw0AaZM50SranNViC4kdQEQL/9N2R+Ge7CgeisKrf3Qms2MEXmdUqT0kRqdYvor
B+965MR8TxWhm8vhrQD1tasQ/13H5ykoaydom/zhm6ykkDAv3S0VX1Zy+cpRQyFu
H/GhU1nWtjU4SCMypwz2ckMCSe+sszvdt6mkK+OegkO4BXVhY3gF2LUkUsLzEhDp
OS6lvvj8Gcw4TFv15AklAivXrBUhr9P9v/p+M+0z7vHHuzCnKMB/ZXbZc/RNXK09
aDtu7NZzKlRGrouACebaXmFKBEYkB3nzMo04be6ZiAsl22UkLqXgO7L2DCC6OSC4
2Hu9BNSnrceWlH7tMm+iPPp46ohbL24wWZtKx1vDLvylOy1z7EZorfhy9s8Q1LOS
W0O9BJslSDOZtjSRHqxsn6WH8mcFFHda2uVJjPXxKCc5yeTmqMVezhn3ynATpWiV
ldNMVRHX8zM5eCGJh92SndgEvR+ReV4jmCwr5p8SvB1OOmdaZIbBP6P+f/Y9Z5iZ
J4fP6TSyMsIs+ONRVvYOHRv8QFaTH9KGpvD0GZome5p0A1QOiISlJWDO4hYo+Evw
RPLzvYQaLXOOfkcZOk8bgXJWYF6W6V14vQZgrISz9q1iJSGPGjrEhRMDsSpmU7TH
xpZ8Dz2Zfrpnn8mm/ZkEO4MK2xSdZk7iLXYZwDkoMZO6R9y9B6DrGGA7OjzExRSe
Ul0zKLdkIlX6DbueHQHtIOp+Y/udm8oJhUybQhtZTFmT13D62b0QIDeFxq9DgJGP
TUWTQcPHbmzgodGJ7a0clAvKpDURZRWl2MusY9jIaNnHra/xEEnfE7lfuMNhiFTK
dlQEgSWdBLc46bZ8LCr4O+aGkmxRkv0jmN86LiZmSiluRNXLxjtTZvRgp0gxrmXC
n4Kd6Fygft1MLjKrs/Jp1Y8ApgqiHEkqN8jsZAOrY27xWU7JNydA/MM8wu/tMOan
cR3abva/qpi713b3LmDlGMIAflukacWOYZIc7+Da/zeMvrdwKiA6SA2PM/NCov7M
hzoaIjxIVAm4nIQ3FekWbtFxHxxjsuWU8gl/F9WRjQO1ALIsVB0vM49350uwYnSE
yUQbS9jfDGzpRjnhATDj9oyJ2wgnBS/hMXlAzQW72KSdf4tVJsz9jZFuvavp6T5u
SgmMycjdOTImuLMrbcUhPqbxEEcB6i+UHwCLlKqyvey5ETTtYeRZabdVpuHJR699
cG59RXkkVNtoN0ZUcSGmy6P96z2FUPOgKiZLBPF9mfo3AXACg7dt6i2/zkw5AA9k
4vIcUFmw15Jn1iomap4p7HzT2mt5AXLMELa13SLbWIYxEUoZo8VLWocuwwMJ/mYp
CI+Z9D9VBg4cwc7rd8u8hFHyaPVg55XbMH3uzUI/6debpGV/4WjrqCjrpAw4ypCF
l9x6ZZtd17/mgAzk/VjhvzUSBjkosDscY2qh7Db7icRhwPQRzdF4XSkjuOq1DBcm
2kU5Gvug6ddt6sibUmaVG0JmMlU/Hy2xx7BiYZ/eFLBjDg12/bA/t1mimTQmYyKg
+pM79ZUuz5L0pTdNtq4da/n4b+z5dsyKRyXIUpiLX2NCY1CVZY3Y+BzHnlC/LJr7
DQEu07nvEXKPgcBlW2vBLHcSj9Vh7f3TqPceF8xjstnwOUbtrM715RV1qJanFfMN
LVSRcPtfvgfCf9rsmbRl8FibeNVLf0nqcOGxC4QqgLYem8tQ1Z5GeCWjH53YshXn
r+bhQB4lpJpCXDnhtOp1R+1p6xjkBO2t8LJya9SCI5x6QuzqQIrNfT90y9EegKpK
7RCQTZAJ6NY9Y/pWqFgSVJl9Gk3jtQNhoWuaihI2nDDjTRdZ/ZWMoQ8m7vWM4LyO
8vUg7k15EUKdO9O+0w/cgBBYEkjQOnEzp6KuU+azp8gonsx0qX+VI6j3h8n2+RD+
Yxi79oaHMRJNvtFvVWVt7+HzkOH18CZD7pH9QvTFwE0Prf7u4g8zWNy6MtHkH+Eu
BkIc6+gC2zVs7nrk2NoUtpFenPpy4nTTRb+9veu6i7OHkn2kRxoWIvr/YIu6TrT9
I/HYGhlgKpRhQ1JbExc1UqOcMAkvWdicMBfwZU+guN9en/xdzymvvjZyiSRzrfmu
2W+2fCVmwTZh7KXGU0SxlicAQij0oAq2IwPSqtTSLeYMxFaF+QdFLT5YVZRijSbY
S6IcxDX9SKjW5YXVdHWc171wzhdI65uYzAnEB4PG8BKASVpOXb1CEavPibmWanfT
9co5LbBPnJK8QfmxIE97X/2u0Z25XQdUXjr5KKrypmh/qlfraa7UnckhuAGhYStc
C9ecZgoaOCv5ZJWeTFYm7ETKJ2ch5FgZebIChe6swrhoVmuulrSvhfc+X+HgCgs0
9qh2uIQrv5pr7GKP4SaEVSHn9NABvqPY8AtPtWIOJ5+Bnwu1BFMYwcXJ8wH6ggsm
/pdlFz89mIe536Gjml7PFE6QI3p0TEpNdAM0QfPjvgd9oaYi3ktJTTsI3m3yzGWj
/NWGglnOP9V/P0I6SppZEqODzzit6SgzlDOhWCx3LwHwsUrRlpLoFzH8awEu9Dzb
u/hibv+dJUTsipUvuTWC7LLTgErzM0zUf/fx4oproaFFnxrpfPRxlHCV99WfzXDB
bUh3bhU3H+lgXcfDyGKOEg0S1wZwbHW5HM/JSPIgA6cILjoa98qhZ601N28SbwOZ
fnC3xtOqN4pBDFCYD48AFNuUN/CLySAiE+tiTyZXvExyEVRyuQsyFmV/fmEJD9aM
yjCEM6EJnofUIIbXyBHoGJG3JC6j4i/56bEKnu/7u0ybLoCmlVSBEHOxS9SOXu3b
OtiSSdCJBYLCgCeTYcqR/kTCYkbKskRjBPb1FLdpgT/b5Zj+Z8/dg8glow4ceQID
O8ElAMAp7b+f25lDsLOGvIkwSi0KhfvuBUFrkwHoViuyIbErEmX5ObUkuzFRxIew
xVrxVF1XikJpgCJkozwwLSAia3YSQ5cicYbqF/+pKqLBB/ShCWewHXHaLhgYyaB2
ALj4c7aYrngWaBCXCWR3B3gRMBJhm3pnCvQvShdon2Zfw+e6PjgOFtki5wpkPucb
1ifDy6ReDlMgqKhv6omI/xOdUH0Ul5uIP/ZrfK+Q7c5erZ+dYQY+YqTC5E3cD3cl
hmsQNcDtnbFTL7XqDTbzVWanUHyAroirLE82HKb0+HPlI9wir2U5PCBeMCqlJmYp
3mjg96HJeJRP5Q4n1/vdXU6/I/y24tJ6Vy55HOzrXay8WLx93e5V5E+R/Hh1kZMW
r0QZY6Pp3EBqePSstouKh5xGaF8LKzW6EFz19p+6OI8n3d9b7/3lM39szGmaeVJH
sHm9PdgWxPOf05OaVAOUd3qZnURCR9eVUTNGZMDCyOy3NU0DDkBsdeArxEBa4nCs
L6i56V3KIFcUyQBVWueHqS1iqJSXYPfncsvbUbHg9GFMW2Fg609kjesSOBO8PhWJ
Lv48WHPa84iK1FxGOa+idyQN5qvyQfG2yB49LxSbqam8Bgywo0uSYas7WoXOOAXY
BfgXSM/fI18FDbmcey5gWwL6+bntM0mgkSEWUspr8SHLqhk0p5aDf88NGEQB88P/
dTKcnvV0oOM8y5zJwzB1nct8CIfnPpSCBtFUwya4nWDB+1qn9uzj/ZrmXOvkKaOJ
6AfwsotTA4eC22FZVKUkYjOGpJZuPDed8wTkWyj42tHt8lMFAB3SOntk6cWTusK8
9RTNOK0hd9B0Q3AaFjxqOzicP5PBqsQ5Cc7Im+X6T4Ei5DDpH/qj2HXs13Vfb3X+
chnEtVtJ/Z9lJjoaTbQIiaaT4vFCt108igHnW/qLmyjZCndg/q4FrMCv0rx7lfrg
9K44BCj4UY6kD0ydf/NlRgPPPhyb/lyhm/ObIKyeBzzohGL7nLb5yTx/fi1vUrtA
LfCIJ9yoNNAjPPp2O3EQKAJbXrJiza0GsJwPW7PgSRKYnh2lDKDz0U7V3fBOtrLM
bz8ZDkCxCXuHZuSJjgkxcJBYVM9xN0ZgfTjEiep1A427LW2ghJtLs28LqHgyFLB6
/aZhaJJvGiRcjw3TK3a+gzIUhboeVL828hrG+IISk78bLiy16PmfjfIMYYf4v7Vl
F1Kf+37fvZRwh+BPY3a6K2HheagpREJaLtkhImSlUXzPd+YpEzW+/cJagouKZ4Oa
Oi+JqVc9FcbplhxjxnKmlZS/q+uJziHkxxOWxIREKTC+6uhz2CI0rYHNhy5MoAIn
jcp6rsWimv9V2T6e9yoc8La2cosqTBpfzaWzz8AVlLlKVXD1rFAa1TrrvVHu1swO
s8zKGy22l6nIJcl2gqwoMMNQMEaeyiKnzGZIYAhRpvuxakZjLT0LnYONcFgpCPQs
WGFZl1dnVrGPyAvvKE3qM3EF1G7JyT1xUsNTbmIC+31q7ptOrN770WT5ndr1mhhQ
2JymaFf/Ds+7ynSWOKgK6g5SXb8POmunI/cAX4IhwJEt7kh4j4QmOOAxJYbJXkhI
mbq131m/HYZVhB59Gql7irXao4HRHdOPfRGZDcKuEdXzuizscAdGVaLJUeruMiFt
L6EnakbocYAC/YsJ5w1tpg1yArOTmL+vtg1hdT5f/XOmXc7m+LcbVYIsRnAzCYam
TmBr0gfB3nQvQhIEZ6OV39IRZfoYYQYrDLTPpVex053XgwNornUAbuDut0MmCWn7
/MPdxoAwD+Ei2zH4sIcD8Dtt5DRksUs78HHgQwOnexQZ5YDkujfPP4U67LVUtB0n
mxZzPvf6t4U++3EI/588RCm1ADS3QeDSnCBkM61fuIOlZU1yEjSYhduCa1ACN4P6
aF5I5FoLyXqI+zqliVpiGp2R+9Tv4nZZDFdJfX9TjutVcRymZNnVE13HU0EZ4C2C
YZG4s9Z2Rp8ryW8Be8s4H2sk7j//HV/fkN+TzTbg50LvU+LonsNGU1YsFp3Gn9PU
PXFKmpYSLO0DyB5vWrhPiMf5DVUyfQGB4g97AbphU3jaSlY6k1Rg6SQh3fhzE466
JoTpKZ7/dWokri+SLiWmyM32Fb0bntdivBLuHqvlP0bZvpT66lZ//6PRXYX8pZAR
TGKK4d9cLpgedchDtEAPY4j7iRd/s1iiJ2HZdvJ6pRSVLvvJ731PNPELAXOpmuce
4sysrlqus9+KWjcyyU5UiUDBrCvY9VNkygmcLA/gw/e1QbbeRZ6oBEG4tHSlIqUp
TE7aEDhsEIwSrrcSWIsbUjci5/8L27TJ7MPL4/tMntDd9NTgodE9EnKlM9A7icpI
VMyP25wCfw8tr/Dt578XOVlDuL2jcdWJgpLNxGj+Nas0TFpw01KdLoYu+lp4BNNG
C8MWpQbTQEENfKyxQBtKVoUV33O3dzGSIfDmfz0pfzlAyHSHoJJxQX9ZrzVRc44w
j3szKKBhyUqDDVrAWPlTMSMayy5sVt7WBrgZLp/4xa7XBOYudJwbEOjOAYgZhMNH
s8JNu1zPPE8Vl2hKtakWJZ5CVIONwHqb8yuFkOXPmbn/1kUbqttqnF0PBVQLpEkj
SK0C8/HodUhULGM2qaDr+2U6xZ+p3tbd8usLIwYBPunUVHFMK8jibGC/R/stjGvS
CPD3mvkZ8FcjTBVR3PSE6GcyawvV3uOXMIiGHvpi7XUoTbgTnPdOowk37K+ALvA2
JV1d+cJ26D0WTi9sCtVoqlS2z4W0wT67jjYaee731xjpAtPGaVi7w0VMDlJVSjWs
SoZZpzSBSB/5VdZCbAS+RpZolveepvJfFo2vd7poF7j8wuXtsywPH14kA+Z8+T2M
ZbaAwn9RrzTLfqVhQlNbVN64GJz7I2IEe8MPKhTC8pm1QF08ACNshp8+GCLr8feY
0Og99KK6zLI7ij1TTokGtCuQWml4RFxzdONAqLjoqK96gR3wfFkcin3TVCEq4yhr
jp4KFWAJYQwUWpMuBwgdggWxv/K5m20lkG0LgULgoHNgPCLwf5EJuQZJ3ZfcjQxa
SWO/63SqGkNeXjgD8unHsqrtGHz1Tp+zBMjp1Dn41MBsWdBetmYom4DnORGNWDnj
Z99DvPSbJioDzuJcWEmO/Alb9kQpJBcc70a++hcaLVJdO+d/jpjNfYXB7KVc+Gvb
FbGB2RV437FyOFNqEbdnO5tihi/iUjVXPoJfO3Fm5KtE3sCD00x1Cc/70IHBfTvu
lGxC/fdJePeZWAzyQPxE3yc4ubQlq2zaHfwUe+Q0eenYPHplQJwqXUGqSVAVCjoq
/n/Jit69wm3h+K/dK5GrPMxSDbx925EnL4LiYDlSLudaCEsDZlAEBeqz+Uu1UwgO
nXFCrldylCpXBivNgZVBUbd5BPjZdRrfvEEIHtah0kB6OtChnexxGQezQXqvS2sE
OATSZeSxIZvmwX/F7ZlfqKWu3qoaSYHyk15VIq5/B6DidOB/mBkN7/ihBE0lcNA5
QvOecMSVkiGfzoH2u1AB+Y6al16e92oErUOEHRh2kBWnsp4QF9D0lr2GQQreJ53K
aVmeoWeWBSPbzvAde8NTPZXMBt2oolX6LhoK0LJO62YW23GCh7+n7yZ7zEB8aNom
EjrtUgZ6OMquC7nnpyEj4B2Fe44eClUClD5laUXhKtE6ALtAM4+ptEGQ3wxxhGmM
bOOB2BY/eA5fjxVdR4ai7l7xPAR3am3+oQmdsVISymSLDDZin3PSTk586M/aQvHm
xx9AteoYS6GGSXGfXMpJHihR14YqGj5qt5fa36hP/VARHQ8YZ/jMOCpD1x6DNRTO
lyFqdNtx8dPlpBpcaDgncCJTuiCuFzBn4sClPF01xo2bjyi29BM/EGM1Zk+lzi+o
u95+Z7wU9KBZuzjIALbCKK1zAK0upYLYB+lBB7wq9qUqxeZHh+UbC1QbWAwakkKw
zI9CsSbcTCTg+o7lo8/T7UGAmmievt78rQ+3vc6Aj6S7x4lWCwaBuA/XtWMZ402l
haIwz2t5ooiRuo2qd/KBlw0YSHHAnvsrpyZbN2jrSgYKQKyPsYOLLTTh4ucP/zvK
aAmKe6Png1iraddrJc2z06mo5hqZ2v2OqJ7kjDIBXrQgWTZWY0yF9zTBxdSWNrbd
Bn6KYH4hhwFywARVOzfF2DqcN/P/f+mNi0tSMphZjaKxDKt7b5FHnn/93BxDHHOz
fO6RsiyvQJo7TyZBbZnBDxJPXFev8d5seNoW5D+zvwozpJqHBcjbRy+QF22xnvry
NKyhgOmfjncRKo4mlgDY6Ftyg5/fhSsrY1NRbbuOKkNW+ykSAVpnXSxub0gVtKeT
Y+bGePIQVaGJXlAiFOU6HO8BT5QYtNPjUc9SKL1JcTspdyFu6V9enFkwwMEkpJrI
br92N75bW4XfoANgq5+wb5Ec6i+NvWrqeNtV9H0NTr2WD9pXUkdZsJqOLM9IRbkN
NOu3qEBN20RStG1dFoeQwWbejSFA/FWtLD7qfgrIuvnKcl7WB4kW+9dLSHUEtfMo
KLvKsMAVftMP/00eJ4a9UhpPPHOLJURH1byVVDosgYxY6fVMCpyquGeYdU+iaI+W
qMXkDF8jw1IyUOPUYNfRWKEJkkzmiLWnDWC/RACFPxRKWaxnBNTF3/7+67Hf6UWs
rLncMeqiELCP952M1peyxQdcSHolAEQh2qZIK5O7Wx8rA04fBkyowpKnacSx4Rj1
WVLRoGjWSOcSG3wDgh6IezFa6KnwgW8wYgCsfrdGizo6CnQyayxIWN07XGdgMD0J
Rmhmf136oDHFqW4C/CRjzLHu9Sl+P55mDgoSTi47fa39OSQBFataTpqPpDooy5Su
YUuSDN+WrFuYc0S5JZcJ5NnAZx71zsWj0w5GUTNLXhxKhEXC/QIQGZmOPUs3R4vv
M2mVZ6fj5bBpGRNGxyj0fYjllChl4iNhkuwrdgDhvxbywhwuRtqWChVPdXy5Ik9l
TfdYJEGDAieTr0ipy07+rYF1s8rl4PHIqv3jKiApboUDGdSa4hZ5lQgV1kbPhuuT
7JYh3cE70VvlQlPpH3kc0L9afqpVwdmMZpX+2BsLtkDQqftL05ap5/eodOc/chhN
laaGtvCFcoMtgCOmuXG+gKyl1D6dW0ehhDydTC5+uS6/b3IK3lXcuTnJZjc92EPy
jHbJw/iwOq2HVtDrYp01/8XbHYzRUgQvLqmiETUxUmsbv+Y3YghRHgEhRkSC1H5W
v5BL/vbMhAxG+Ja3VKFCTs0DKFp5tQ2EHGRezV51XoHZW3pMizmR7tt7kJ5bRHoq
SPld4zyqMmFrD/sg4eptgZ4+hTKMjmD8dL6K5ppFtNfxwLUT6PR4ypiKrRY83vLp
Ogt39oyXk6pJl4QsAhGzpNz0wZUs1XMYw2hZkPfy8xaQo10majFjnqLxOpt87Rd8
PVDEBsbzYFun1Wlfl7q7GtqyQVtzYgUBGfMzqwxk15uxH6C09c+dTpk15ZeARCLl
lVpfN0PxPXBPzxnDhxfyMUK7HEXwCq4eLHmndvDoSRInpUwWMyt1kc59NICgLC1I
fkuvcEUrIa+U0adzstfcw3AMhL+CPDX8wXRR+cCIbMKYETL/E//94Z0QgO9CeydV
OvZ7BX8nAM/Io7iQf8jzWdie8z1y8gOCzZrAZR7tzKCFvJGht+y/K4B6kpS3GPG1
Kopk6jsC0bOUOq2h5q1hVvPRyBVjgZJ54bpFXvJR3IbLWzsywZjr4Wt0PFcy8IjB
fjinnJU9Zp3k+tG6V7niLfbOKS9qPEiqaOQRNB4Zg8+c+zOgTG2bJKClswmX37+N
1swbxTH1kEgCR97fAvbHaVfMg8/mbjR5jLB1Gzphi0yjPeqTuyqijIja2ReJyHXg
I2ilgDBg6Em7eh5OmRpyqKYHzz9ba2OqDm5lX4mrQARmsxxWA8tsAe0le6MKIDv6
YGjbsIxHJaZnMYIAMJLjMXvKZsMtHruG0rqfOGNoRfRoYq4XQaNX2599lesut8F6
5H9SEp8qKOhnSDVB049SvJYtXHlwKv3fANCIEooP1mbTf4Q6veKmLloeIOz8PbRs
moIwFD+3UCWSr0WM0M0I5LhcdzpTo/3nu3tt8G6um/C4olG04bU2q159rzdrxleE
g4e5Rty1MzeZY/pP+pdB3nJBxITFRcGjGIrDpFyYl6wh8E/UrJS6BaMvY2+BKI53
gO5IJF18s95coDPkJwLR8Jdt0AQ/nKi2ZtFi8JAhaLzs/1KmYdYi42/ToTrCQw1V
zpqzpRXaVHgwp8P8VAC8EasmDAhN6as8ZmO7h2/oaZ5+ARROh+CmI045BBS1oMos
Zjw+eNbG+JFxH6dc0WlkjRZqASDzKCi+3I6zOj2tgX9r8DViLe7n1rPoHf1efZdV
Z8SM43a/8I1ka61GV4wSkGbq2cx1kX+Sqaf21dUCdKdtX35GwCwPa3HdTKA0bSRs
ytQ61aLPX30JkEE3hpHLFXvnVgdGdKjOMDgWGNDafmh2c+W4MHIFFk1pdibrZjF7
CCgX5FqqcNOrgtfMglHKRe/2vSSPWoEM7CBc1VFt1bCaJOvGEBuLqdFWh099K2g3
qWoSvu4kkWBDoErkTigU8fR/5uLBY8d8JKMVCtWfkXa6Z4wmz5j33yrcCQCinC1S
mIDb7sTHtQS+6+2Oki85xwDVIoXLxzgkAhVbrkBg8Un6tep0dCT58xuDJuMKU1Lj
Of597C8Wjv4b1Gmn5iePwev6W05Ctjbe/dyi5tpdJEb53hztcAkAS93xaAcWwiHT
7jAghqC8zEchG/PPabRoDoGlBZmiSdnamPBUHkrwkJpujU0gu41rfl5WUyRDls+R
y3c7it5dvJCsblDn9/wu2FRBhpEcqXLjoiIpKltYbnu4GR1i7P8y7s5PigiSrRJS
YGdiHF528WWs8g1uo0NbrjCPmxTIpv2TdsTErfgZyEpcsa16EONwmuoGar73t4xY
vNX4r1P+e33fYOB+RqBgV5HOWq45VvgM+zCGPzp+KRt+QP2WD/bLxbgGZaHV46N7
w2hSfTi0p6hbwe+xJU+vAUVrie6/v78QjKdrZ+AlhOeXLcR3mhqOhmc8yxoLT44E
UXOOIpFSRWBErEMlFjL8OLzrEjxkRnnEkOUOwrzFcttUxnu5/si4ribQrlzgEuvD
hVYaLeECuP4Ned/3cURjDkhLRBaWRgE9sGUecqmzC+lj1zmCjosZj7gi2shGC2Av
mi4ag/tGjMkfd7r/HMts9QituAt3rictgRw3E6M+D1ZR/XsdKrZRd0P6ZrSxqUqB
Z77i6ansqDhhOF/Ru4ejctZ/lDoj7IY3VEsgmT+s6tUOi2+JSjkordHQZSiGJhy6
WwG3Eebb7Lh/jrP54FWUrQdvKN8yVc1+6UnYsWU5y2/ubuF2LpJZKyD55abB1XlX
2X15gY1rv0zLSTUfODTGHzbjnEkvEQazNuO0Mtbsz0RbmE8RiD//MumAuwLVonK+
JMUSjlcvyqjr9NIyP4Ljdyi1VjmqoZHfKfgy+BtTYrrSzrLBbIZ08S7n7630q2MO
zotSgs/jVN/KVL0/EZj9x1K/AIvXoUbLJiMzBe1V6Z3cuqxUKtgeUD/LBOjoKGgN
XVIGAxEI40/hfHlUYbV/XTgGJbAl0eSbFLanUTyRDtSNiCzuSW1QqyuuWXvUAR3k
HOm2KkZ1fp0I6soVidcdcub5m+XEUtMmq4ApYW0qeUgAempfp+8xEBNvuSDXOgdW
PfqZkZA0rkR/UVGM4jqifqSoGYIsaKeIJG8hPdm5UsEbBinWG7gqfHhaVWtRiQRp
pvmNAO0E9kBA4U2URX+LcOEVT0QUsae5FkA083V+yMxXMktdRQn+j3KVYHnm+iQe
yRoOKRj5IuaFGO4sPKHaI9z7HJuaWGDRFnfTpLS1X8+iq+pjvvsxTiOntE3OxaZK
qQU54utjuPdMMHZjnJMCmDGPyo30AfGm8oCAUGwkmX/kthJ/hIW+ErpUQ6oZN+o1
PsjPDdh2J0sZFmFZLxqy+rNMPcHBVh3gLI+Z2BZj+kCG4BtS2/D24ALSzCKP4/Q2
a0glfvpEf+C/SFj502B+TN38qbWTvM/1PWKyvpj7GN8NxxSfUK0gsYMDDeXaygI/
t6vcasy1sdp2o96KFb9MOQ9TFVm1m3eueRbng0zQQHGw+5l+pD5/ploT1abrqBZm
Fxu8F4IA2UujsLfcN1ZeUUAOGKtTb9T6H3mZKX7m7NO32FKdnOBoNOCAcIiTjLCD
7jlgbz2s5KPVqLJ+DC5rXrl/Fhk4SDpLkVhPdjlW0kdkbziLMtNXXMIAXfyH7rzj
sK3yKFLheJSiN4pwTU9F5lKaK3p+53H1sjss8hqV2rB9mvC8HKzR5GJNA676Nz6u
c/dZNoKbH9FYG8E7hSPKFYQn1YY1iJlavMZVKWVqEKera4hgG0/98c2EL0+hlzKA
rV0j5SAnnJBvw2RmpXsOkZEGmjLC4iY7Cj5uzvtlkKslZ020sEZKYAbGEHufum9x
HZrTPxTYh1W50b1taPS03Z0X0dio45Rv+IZH/Eq+5mQhywf+OZCJXdBzg4qo/38W
aDzXFslizPHOi5nH4D2erGqfk7ZgFT+ImBI9YY/z75+ve88jRpNxCd/MN211TYT0
vOl0+WJIGlqBLqU+ef307jwpRBGeB4t51jPEzr5LCfNXkNioe5GJ0TU6ZvJSfiO0
s4vZ7GIPnVRJXryArA6I+iXC6nwbA9Aed6/eERRwSonY71qcaULupyqaWkNYGsLh
0DgAvpsb72DDb4E4QfSW7Kh2aqtMkDTF+nf+LGfp7LoClRdoMaAOGgD7BSK8BGMK
d20t8+IPBDAcvKYyzaz8qgxX4a/HdyCDP0c7v+GGyanPbpECYdVDIL7spAgmke6q
FbPcnI24VdB3wENHNKkNrOB2/hr2cXEztTZg4mOdahEyavbzBDHfuT0RtVum7LxN
UaCwEMeTIG4ic6vd6CyXMVef+bdxtZRBwytmlEWBRCCm/RiGJiuUjV/2xOHA64C1
17rgXqalAQOf/ItxHho4u69iwbV5ND5PBgcEG+Jt1PPtkMpcIErz/MXesFrSXpF5
63zcRbhsTy0Ugn26TuP6uk3gPoptq+Cc16gtZjDFvVC6cT1tAcEafuub68EWSsQW
jYlE6VYnfGGDa5Kxpgn80rBWimNcREOGduUptEy4qbE+QmJ744W5H6lUaUWRa7kW
BbOvRGx8FINiZP1nINifrIstAznE6D9i03BnRAsJInC5J8uHCD8sDdsnjB7an6Vu
iNN1KPdXTdODxO1Ci7UhUou7qmNa1EcceNWlgpP5KNaGZNhJijnTnBho88bmSNp+
KnhMvx2HkBWbkaIZtKM98gDdUFGtfbAV9cycjYbyIA7QYf6HvSfiARnRUINduI6+
4OZq+JfXbTzHhAceuix5ijYGrPV+K5HMFa87t1/T3e80Ax/cMqn8w2eJVaqw6PsX
/4ZvppNaOertKN09uwLrY11p5lsFu9elNcVm72D+oMGvKySfuc473olKx0g6MXOY
aYqNc5V4nmBORGCkqNySw5D1U+zdFSCZv0goDaJ/FeryIYwCwqsFWq5yd9B7GkP7
/fbtgCAMV+z7s0cl+kUknkqrGxkqGyHK8WxxLk/QaPwVct+D7PZnXorLqP0PoaFy
3cLl396S0mZfIZKXk/4w1PoGmzaPkq9Fv6XbJBGBg1kCeP7VY48QwgJPTlzn3DxH
K53jFHdKZLYlZqUaAdhNp8TdUP0LKtYpXyL74dvZcSAu+bJHyDfJmbgOnA32LP/X
Ob0qywZZSHA77uickbsUuZfnE8vSmptRopdxJsq2ECD6DfWVsHWATpg6q/Ex2JQT
AP85DoSQZWCF2IwkKa1ElXM+Pw1JbOtc58Vame5XUU6C5mq8UhS0nLy472nYxQiC
ka/Z1stLHFOl9/fnw1pN5Lnln9F44ZDuuNHPmVMtNyEXvtpPMC0d2OhpXWGR67rp
ekqxuevq5VyfzJFO5RtoPSuzlf53MwzM7uQECgM/gMuu6G5dCVwU5ifk0+Rf24i9
WEQ0eNUu1xwwpu+J/iJa7T1zCfP2Prs6sd9E+Y5yRMUCTUWL3EPlUdHX4HanZIqY
swwbsGnjjJMZm0+PK0CgFKgI7gsyZI4ydBKXJZ8ZKxae7ZsPF3A58difX/Gz2Uh0
AfXl5WkbrQJfXA4iLwwlnDlQsKKGGI6kgjSI9T3c1oFREGQRvI+62W7BmrW1rzD9
6pXSIV2mkd4pZmo587wsE5e5GZrrhvtRUWibTHZdIyQ28rg+0iRzePRIQJRs2z3i
k3mCEZ/Viw0BqTf1g1QUqz6k7s9KGS1LxpgC/eVc+yBSR6neK1kvilo8Te9bALyn
0ZFCiunr1heWMH0NeAT3WQNymjQQF8LqlXbjot3GfPmoOQJ79YvnuGZq7kxDjSeA
IFz25nQDV4TCI4+Ly8Z517Wgwt3U2nQk8QQMIV1fqQfQivVuMeorfPQTiRjszRXR
pgxyJMPhFl27iZpsKpf5NF+8cbRUhgiRQoCZEzRlL3K7aJ7XNBTpa/0zYkimXvlb
yfyf6kOwkMsnTC9PFbhnr8w3B72715WkalNtCT31cQO7cEdEVZvFg9PXRAmc2yta
slIogftc194DYAj6oHRYwOjCtQ78xZXxY+DRZ2h9MQpLYEK92668FRP74m/ZN4oo
cOEtkby6Dbjq2ggigQmZcJFdIZVgmGwVZ7ysNTfKZ9mFcHElHKQIQyMYbYaJ2dAA
XtY4CJ2jRAZAE0ccyEl5vDVq33IRkjKqtHiplS5B3pcdCMGeV6+QOrA5LYhSFT0a
f9AkAVaggCNEV8Ta92+stgUaz1ZVe0wbg2X8a09uxyCDzKbqnh+l5EXZ1l1QHAXJ
dXPlweI3pWUWYXqkGG7tjsR4kJNix1DKqeU9WafM7wgA7NkMeACyavJmBF1DOMMh
HO3fX021PWs0ymWT/tF2KHs7OjyFbhsgJIz/63ZVusmWFE5Ga4vTmT1DpBxlIP4/
X9/1OOERBfZJ0hZZ3ya4FmgNm0jPj/qu5h2tZ8z+vTk7NgX/yEqzkzF04DWNOaOH
NnvS4XVlXOhxPkZQoi53JY+Ebf5iqxB88ynMGfsRuKTYXBq5DW3PArQXXU9JPlKV
eeHWy5StEVdEcN98ataw5pm3iFzNBmOlyEpb19Myg1LOkIFMOca+N5woBW3OVzYX
PaKsvyhC1eFzAx5qyottYDNspDh+LMONdFcpzwkbmurVtysgKqApqt7lnSMsqI4+
7r1u4LIqH3ctUyfCJLSp3RHif4moL8QLXAWuM8mg7CCarfceuVyjVe36bYcriTNG
lQ4l9uvtccfpZrF+O4vNfTKkU1B3ChqaBegGhOJJRueeIyAmmqwodSuoQeCLz1CA
e0HHAZc4zZQKh1vCPyJo/OoXd5uR6zrejdGtQM69kpSEaff1VOFNDnNk/AsSal1F
v6mbdWMaiZVO163J9i//t7yNOYW2UlnRrxDECeV9rtKzi7DePl0RHf/NMPQAsBxA
dA+6fhq0Yo7lVSgRJ0GapV61n3qf6Ao7IqVg9IjbpHsDSuVFsJYbWWwYx1tiUZFW
YBBFXcracJKxvIT0DfUh5YRAH/zyDvcxAn/tWe6L+sTPr1KJku9v1i9Z0RpAbG4z
RUjSpRmzeyTVB/Ss7QjkOhrnI/Ege55h1oAwpzvebRXfYFNipo8BR/kcLTWXf+MY
AXwGEov+7z8O0habfXP6EvapmcyaF4DJM0YduyA//G1rHrYpyyAIIWH2CmSa2hSe
EzFJ0DZIZtwGARmmMs7OCQxyZZPltUQNeMCytaDTnmSeJmEnnkg4vTClAfqosOHC
9aoJliWoGAAt+hsyOdKxRqtdHF4Bv3nKcYYOvqOGE++lDyj8o1K8Vp/o0efvBwkt
Pc5caCgT1Ll1XwZ4ZBz2xNNV6fAu4WPHbXOJoBhDaFLJODvMrIbc0EDIPpZMPr/L
HURhpC5qDoJpu4CSDJj2Hi7EQkE9GKcujNv2YEeyDw1RZXY5Tp0CoupOBqnCgp+p
ZAlu0ReViPoYL6YYh/d+3tGjXUKrKNvlNXy0vGDgrNqLsvpVJiBvgk1CL57PdQRW
9BavyymacLGkFp1AUG6jdgYkKEAVTpeQq017ONBgFcTSN7Tv9nVylZMtk8TAs36u
uRCwlVSFPKx384bThUX8lWMNE4TcOLYF4ib5lccSXdE12o7QabkMtLtBUuohM8aB
Hc9FNJMGgCS0YpGy8mngjgV3lUlbMflooR6kvBeJ6n0E8vFN7qTMGAjXvpUT9RhM
1ahyqeBGRLyX5gU106zxR+HGfdB/gqoyciXGolXfcFunnefWBDaPMd1EURPtKe5P
TfWxily8Xznb6BG8SOtGvpG5eypRHyCXcodtEJumPqJIacbjdD2jzZdUPavtWam9
zjsPGws1NWe9mT5fKYoIc4iTXtrr6oSyMZvhwbd1KikLi63rCJUf+CzxNy8aib6j
eB43E90SmcbWMKdSh/uCADOH503skPvArzcjKMEYtTJ+NfP9VL4Qg0cc0DOfHKXy
pjTe1MC+BvqP9XmVihCaURibly/I2zB0UwC7Cfw68Fk2XOKHFyIwj0iVCqPXTUhX
W5tT66hWuD24HHHU40yFGOps7YgRaM9cRpClGIQ9A/p/ZMnsvZO/CzT6eY+IrDd7
nqvfyfiCaokYxgL1DE3n6E3fPiuEhJOcCOmQQrnalWqsw/MH5lVELDHfYWLlR2ON
EUtCXqycxz0SbIXsCniGn6BrolO4svoEqio95N5mb85BXULv+Jn47V/MGYPHBgrr
HKwM4G8RwhnvV8FmytUOrehRQb4ZtJoB63ICyxULFuL02+f5CUh6PXNwqq8oBc2R
Jpye7eRvE9dO+VNdJQotCXWVAYL0IRqZRRIxzbYe1mzuFNYyu+CKqUka1ADGVoXR
31EVt3e/jCuL3s2plzQAYaezqPCweudapBMniXCmVPggIa6gF3ytvMH/ZZCuEkgn
JcPsq8PZ38iIKdIy2NbORjHjlagLP6SSQ0M3mtaoXwtwOsDXAdmfy9m5kXOexAvx
rqbjt8Ss4wqXHvvxIc6YeSVeYRQt736WOGYgbtTGUpLZhqQwAETJoRUZwOXnYyfJ
nrdWsNmImPQKCEK2GwWjIatCvLcuMWxWyurWBKuW5bOgSP0e8D9U7QljdBBzoMHQ
TC08H7M+o4e4iML7NvKjYv0Rb2RafqrFHXdUndaKwcCe5YuCaY+ARrzZnPCrS3/P
9nZkffMLLNxc5rY5JQc9FktH2roJ97Z21mYrpn9NEaRY6n2qI7rtms23RQASlIkh
fm1asMb44x9SbAQMrEZU+6mLaaWP2HNlJeLxn+wIeiEumtgYAPNZVXu4e9Z2KGCo
ioNBxafaWZGGRKd6+tc/OLPUXPbvd7ngOll0vuZxS2v39ddwA0lLcRy2YdHz7uk6
FYVf/hCmYVZDpyTABg5rANRxqaSzI2RiaxgucULWnyogq2S8e43VCCUF8BIDXdAf
oMr/GvsVmAT9rlBu6oZPlkZWBwyOP01OZg5d9zmAlgdhkGPDqc85ny7nUMYRGgsR
Q/gGW/b/5/e8XkLqw0KjSYhFWC8/NgIl8bC+3Nb0pAxxdZ/zM/g1sJ8e0o2EORWM
dqbz9ZptGDH2zkoDLWGqL58wo+hT4KKh8lk0mEhkdfa5bGnxGDW/yQpl+S4l/ljC
YYrQXWu+8iZ010EVXYV2PXeOMDVEmLudQlok0lBhgbqV+M25iVkrwrUV1ilpCIdx
nOvxVyy2lFdPD3aWsn75znjPw1cSrk0gvbpjAUPld7M0fvcFmzRy7CXl2WS+8Rym
Z28FhqQANpFXk0qqQfdNDQJ9KXgEZBmYK1aa6CVua8Entr1rQiJa9Nbg7byOkH7Y
lepPgriE25I6mXOGgJ0VWsA0CnWBpK0KxSNa4hkpEI/yZcvGuVSYuCHTh3CpCAni
m/gT8NcOSk3jm8AD854HxXRCwj8rXXPt9WA9+12WqdqmfxdW/Jc2i04ufjV6hoKE
ppuBNhUMmTAPwNMQ6zgsbIlQuS6WrjFyvOGR1p9UcOGRB2BEfRnZMzd26m64wpCK
hhhGcD+HIkU3KRJL1I6cg1p5mYLcTxz8OUd970VrSHrmXLvRmjN4SeFBS22Jff8q
+bxlMVi2oNMrcfsRS34CFLzsRPPeJyIqIwnN6sf+pqbyPKBZLytaaSIsmBRBAWTW
oYgytCgyfhonw2ROJgW521KBPc7E0qFaZ+vGiGXXP4xtEu0zaojx1A8bdIsXsCzX
Peosf6kUoFjAi1u4gdCHZq9IKpvXSgjFyWykQsSIRIq5mQEUziWblfSDJrTRxycq
IFkDjB8Lvc2HacsjEtx2ik4lSDMb6yv82DdPxYjlMujUgyr+tswv+R9B3TBOXrOw
pFr3HwmyeCdcY2DgtAgkRWFlhG9Y7SaeqsacEnDMnEBPB9iPLUdcN3AqYWPRkgFj
4TAp96X0FhH35o0x1ekBmgbmViswodlDiew7e7ZKBd5pEmAMDQqaprzh6CNUUax6
V5XFSBWvNfQK9HwP9sBbSYyJy5obVXO/aAF+fQebvLgTdauAE+VjjEWfRR9F4kky
yEfTprbn+c1g5XfHgH0yo68p+kiFk6lzTXpOh8wjJKqJyRvwedEDByEO6h6ywOIn
lSgXQUKJP26MEK/bI19h/DEPDR9iJznp/Fns2IChofJRsFvCzteiLU6OqdkX6uU9
Su0tFF/j5rbb3Eogzz4HgtcWJ6900Ig1+JlkMCpjfYyJnwx7pxH9ZQTiQnmaztyO
ivuZQ7/JN3mfqVdHAFl4PiSeYB7qJc+0wMLElL8s+xgEhvnAn5pVLZz5uSUDRCwZ
v5eT9LRqvSZtb8di+QLUNN2+ANCOrYiiAANdFt04gRlqynTIDNnArkNlEGMWbYlp
9j6+zNvz+SEh+JFxRMcU6jF+yxvU2bRji40myFbgtYQ/InU8J/pYrw0Ay2Yn/Zu5
ZcgyVDUgz0Wp1GenPT0qdD7JsGdm01IXdbHcruKZMWM7EcfUgh8NozWhE1D91R0Q
h+n9qwh6TjGIjhcxHvToh6ioilC8udl0Gr7WImiMcTAnk7UjNNszBgB49I/ejG0z
GKfNZOfZblmQPgCIF+aq4/ZTx0tKbu1tRJsyDN4IagEKR54YivFSJojpAlr8VT1e
YCvGn2cfxOCAoaIRgpEX9nS8elhHIc67CVUefxtrmDelF7n6qNU9bmPMIMt4AzHc
p6ox6YsIV+zbKoVRRmnFezw2bx1OO2d2g0UF/wH/UocQ9WBDSer9GwTQggtJK8Nf
sMaXIUorgNkYwqaaU2ocy9fb5knj3Yjq9M/GxHYHD298/Vc6ixw/8Qcx3sZvOnMl
ufhP2s/qDARhIfS6aZiPQnMGLHH5mw/uAFQdi9fekS2QsbhUVYWBTZ3u/PhV5bXz
XMqWoc+33o6IAoLtB+7YAaQtIDpPm5TviKn/85LIrq8vJk8rNBJssGHvsOmfILPc
X+lO6uoO7cq6e64Oohi2a5bzXs59HuUS0pK2AaGBXdZpvgBTMJexXBcAVnk5hQwm
PbuRpetAe8lljoEo1NilW2STdCXL2AWUGNwl6ge39QWdSaXlwrYJWhJYmT+nxAWX
v6GxhDPjSJnU1w34dmsfko9V8I3Ydh7BwUx0GyFGdxE/uqH0yZqDbkMZciPOCCJG
whoE5Wa33yQwLBj+sQ4y3Ddglg5NOTvv5qtEThBsViQeIhCZX6lVJVxvmu5fALSw
Rb7r/asWyKfjyeR5B17gYZg+VJoos76tzpQiibeW6kCqHvBjpa7dwc2ZaL4imp/S
V7hdJuJTJrK8r8k1sgJyXfFpUFzusboIQm+i2MYcQ2DTFIeQ7JODw/uln9zhtr3r
QqNm8/e/PrAJVBQs1TZCTsjETjeiraCF7Vi2YU1anVBLqh3eH44qH/eTrifGQWRm
3/9rOpKjWB2fGRhM8Hw8c29Va3tDCAu60ye2c5ufLKEvMFPWrRwYQtJJqJ4/TqPa
E8WVAB5EWUG4HsZogmrHGE710jL3fDZw+tInbHpt05RXE70ScPqAZEdH7b1H9iEA
tdAcN080A//0tVORLe+8gK+oiad5uVh2co2Z5Jk/6dySXNo2UFqnTxrSH5ejXwJv
NbY03SZXTIX6PpzvVptn0N6akFATfM5TtO1hVDp8OWqXa9PuJGg4bP74mMnt4hB/
RcAi6GQYsvoyHEnk4LXnKZ2iMWc16fHg6rHpFqCnaHjQJXeeHfE1PeosPHtBPFZN
j46LZ6OgQbw5D5IYwS2AnG9StjNfwC1RDNAoqVotPBviZu0DjAuBmTOEYCWIxOqz
ZLLEtOfYOkvPTlXqiv8PPfJ8S67C3qcscULaN8HyVU5F7Vew1ZZAk7fJHL3BFoFD
SAwTm2b/fRgfKuZYy8vpTZPYXnEzK4UZMN3FnZZjgITT4zncYHOQEBLlmMkSFf8x
ZUmcU1IAyejSxstt9GxbSrG1qpMMFeQM7NcnvBKPLVuPuqKFgJ3I91zkRKv0D8HX
OCGui446WrcgbC6FwoTx+gFWDpqdehqU4CXPH/76xvh0OXZ1HVEaSIDpKuUmAfez
0oDgshrJqv8CgVmyffZY2WtJgzkGtRjf9bpGwFWv/HLmvS1SWg+nT3x9KNwjhxCV
Bw7hLuXKh98IUzbqzsvs+0Yn+wAR4Bqsj28yAQzlEiHBjeOFBXuT1peZ7jfJ037Y
z1OvP9msZZr6w/tCQQKaFZBhHjMctCeYbl9/vTfO6svktAZJRAvkPT/Iu8kQ2s1V
UCnGptsIiqEFKr8cSkehXI8cSRudrg42IWvW+GyqqPvlG7/SXYQi2BuHARtfuycW
kQm/7EromYF3TRk13Fc3axXlxrpSrqF9Cup61n4zofaoYCcZ/IRnf/f2DZCh/Yso
H0awOtkHHDWIY5ppyoO735QmNaq55wmQI95RjFcMY4taK3HASMaf/6q/eHA0swsD
WeQ/wPPddo16wGQ9UphRV2314OoKhQs4QZ/e0zwiOBWupnhgzVmueAt/ZULwdQR/
2ZrfVy8xbYftqESksIn7LKYAMd+77dJ7rol+c5JqiqZQ5TqPPPY53DrMnGpR9oUI
CTU/TotJOS8SJN0O+46IEWiTN7xx0eudeL+jo3EQdNS1rcLbscJ6/GxyrvhZAZhK
YMP1HvIEfUnf2MAcoe6PBU88wXPtwV2oZo2SoKSpagyYMV72HuUJ02fH83VCNvwK
vWC2SxrDTkn6dVhaUG//MO66UyS6lmT5vJ/5lYMeMSaxy3RW67TASBlzOCq/KAG3
1WEuF9XxNGKbp757sYYQq6XMpkI8Sartt7hHOgNaqnLBCIbeP2szZFg/lU9l71SZ
49c/crIiFmI2iuAXfssVHWEvgRWtAviza+l4BC0oVGMQvZe7VkiQ4TkHOJkTcHt4
UQXVsLOTTqxJLndmkXKyjj50+oX62IuFR4TzQ8Q/pmoK8MZjhUpVA3Ap5DcmZymu
f3tDQgvu1DugSd1OEpDq6GDAKYhcGdGWE6Nbo2yqT0z3p65BvyM08HC4KOJkXSZb
ATgZmT8oAdrOLXntDSoUAKtwkhJ5R30qm71W44LvqRjWW3Q77ALCMI/v6TrOw/UH
fQkKI7eikBHXo05VERplx433aourQyeWmJfv88D6DpUf8RnfjiKzhFs7JsoVRe0M
tPj1LtGjT+Vsmadtmfcq900d5CLZMA6qMCqKT6oeFX3BeJ3tJOCKEl+I9O6CX9pp
bNeQDz7wB5gwrq5K6hgr1Nmg8UaY2Ahy+g8cd5VP1pPEnh2px4qgLm+ZG0nbS/HK
SxiUrlcw0w7GtSE0uuC2XDEZUdrVaDjry0E7BvlbWdo7yh3/qYO1rkyun5sT/8p6
fuV97uQB958e256UY/jODo4xkgPWyCWe+xIrxsJYNBA0b1zeqQEDQQYNk/jesjIm
NgY/S314sSRuQnUTwcfkhtfSKPW8riWxDR4/e5wEcjue4+P0mi4lOMDt7uDR9h4f
RDEXAORhZS2NW3p53AaF/1eReF127Lil1RFnH6XX4eSTQ9Xs1byUbV4oyOMzmnj0
GmyLTnFR5rh6e7ArT+Er+tPEnYdgMd0t3lxVbH7MMkpyFXygtjJ/XebOUiJphl7X
gXfdlfGvTe6xVxWxrT73r9B1FK1Gz8PY5uGYMCZ70OLXk65SbSsx/xs2fYa1BAWt
anSU8rV1/90E8kr7PXzH7qcTp633VrahjNXSyybwl3JGjruXVEQKVffCOya/sAvM
xcPHNnFEZfR3OTkz50OibNIjWt16+qLjF75IktS8yKzEl4c5/Jhe1R0lQMCZVF80
RY7n1ucOFrtD3IsvXeTlThXQsyrzMazg2odakORhekzVwC0EweOwodTSZ/S5m44Z
zDF1gZVM4e7w0NElc3i7AAQLZY8oKoEJHEUqL9/5XECMsk8RMgTV4P89OdgdkP4P
WFTt+sCvW2+U4Ghqpk1py0Hmn0ppvcNaObQ4CuPTmg4xunGzZKlqCfHwE4m5bAqB
BKIj5edDZYiMQkwvViL/tzoJ7ixdlg6rPn8muOmoZgy6oEnbHSYP3D1cG9VRNsSf
nJyAmC09/G4EhYNSols3tjHMaXyaY0eycUELKAVoiuI/NQ18bd8d04w3XocQhkNG
OKGnZr98RPHeQDBo9AGAdFHg13zNgCrwrWGp/eQMNRQWtBvFoUHPdduFa+uLY1yl
H1xTkZU3C8N8792APP+rk375msTbSdAL5ZoUz+3Kcvr+KtTGWSS6KmpB3ncLODmM
NdDYz9tub8Ji1dU7Ptcb2XR7wYLA86gkpS+dSJnHhlaC0CNl334USIQzByuZivoV
CDltnPE+KF3QT2Ct9d62cZqbfaXkVEZ0dPDGqM+XuOmIiXI9IBxypWe7m5Qem69T
oq9rlD+uy5oDn9OS31n2qaqr9m7sDGQ/izSHtVedSlcwKBPdZhBPpa7RTA2VTHXS
MzPenmWEnHI9Nv6fuySDSDI9ME5jnvq4URI42LJvZQpw1st3lh8qq0IVJHbzHTog
rkApuc1hSKbdSX1/UqYOZYnGid9i2svSZ+pASRp6rVXkBGrfHTs597J7eZqVoE+M
sTaMA4QbGf4wNhoio24MiUNVqRGVn1Wxiw2IPwXeuPn8LeY2hbzDy3nWx3rPDCn5
xRwEAA0Vx35weHUosb//B5K+1cdAwtNEtiI28WTmt5M0XEL896kjeArWADj+2S02
KdZXZi3NlVvIlWu/+5NxCROvCkzhwVQ7f4FMrFLIV1QJ16f+GuFpRYKRdWlvNoVM
l6uXnvJExn5SA60W9CSiwRdL79U/NqmB+oxSQXxpQvTg1F/e4IQmEijM47sdZJA9
YPzxULGCzOK+Uz6VxC88Iz8NMsIF5LdBXxc56Kld7HyNmUcL8y1aQSJx+7VwCf3W
1C3S4yy2ISXArPw5sDKRPUxrdDSE5QeatnZXfe4xma8/XtIkuB3DPAKn5j7x/i7q
YZwkc8fUAuoKEg+FkNVs5qs+0+jzInqw8WbK8cCgpXIpdMBWlEE72QxCPKdi5wds
Zv49QvMAOSHojUc9wOgIXWFFcT/7U/JPrLFLC7E90n8gVjb+5vUPaw73tAc4QrCc
JrODtl0k6hZFYMurG2BBt0WYavRJtC7WmkMpSPFpJmvI7U3Ly9tKDGSp8nbX3y8N
a0ekuGx88H5mLr/PaGU/iPh2pV/JJT/PvwvWQxR7ftL5qMvZZsv+WI3RAfBqdBOf
6MAOEDm6KggrSXhLFgIkUhd7cZeFQ4N9itxlIGP2qm1syehrBZVR65nVC0F1ijMs
HnaXzsUxEa11fEwffDDrrDnAajyzSV859UE4gW1u/sxgqfijpkCxpimZ6uBen23+
eNl+59uE2iAKV7sD+60R9sxguDH8cEPwnJ6r9yNoNYoQhgNx9Hc+Sqq3IXWE16eQ
S08zGu5vhi1LZO5JH/iXBmlfTKKObIDYtOkaoH55VGjb6d+ys9RORTRtk8BCb0/j
6m3RYfR9qa/KUOV0B17fTHI08NpRGQyRtl5V0N45RCOwz04w+TSAJa6K84nNBS/7
wnxa6eVtpLcD80RaCW6I746aetENwfrb2NtNT+xsqWsDgEZ9UvJ3JKsNr/LDcWYF
wb+Puf54H4FUexmMTtH49KaQCPbOZ8tzTMASHI7+cFS/jEkaFNCCCm47CV8KsA6D
YEFSGyt4QugehZplieWUmDTRm6rI3Mye7qN+uiVBQIlZP5Ckxf4YRmMxlc1Nhvth
qJhfP0q+Zy5VgH+DAX/dTqnY58xJnMiQhW6Lyd3hxyltNr3olC6rcoM/OnD8zTpA
zo0X7FssX9zM0cO+sow1vl52gSWBttRBfapO2SxoxiiVubJo+pfwzpyzC+uwcrwV
Mc0mVQGNooe5k0+0tPCgKBRaZqoI7M1ok/vS0P/QYBfZL9X00KU/7bQBV7UBRcUs
rTcMehteWmJ+W5cvqbIgA5A8g21DOM1K4OmLXRaf0hdv1q9BKZhqeWD0xYYScMrb
haNFuLFG9Uq3KLUJi9AecNF/a47P6lHCeiEXsbOLMa0PLKgj+RqkUw2W8zO2qcK3
H6Doo26nsGRzcRtKorYu796zeDa8BXf6hNUqcV58vd6zUqp/zJ8DEZoySW+dmt54
lk5/q6bP9kkcgZl8vOY0NE69jAh2Ct7RdKQMKcO5YdfgsXGaSu6iVq4UL5O2LkX2
hrldlK7IJPT6csTq9B/z780PPCdlXxrO+MyR9iMMdu5F5lFq+D35GIbMWCaj7I3U
Q3LS+1hbHW5Yri43JknLWRqo9Dhnmcjx6aS7cbIdU5N/HG1VNJq125nGylkqoVIK
ywO+qDE4k+VRJFzghUST06aZw3l6bU18/1KmJwAbxzWneOUnfiIr6kpUczMBCV3k
/F+eMzsb1V6v85V2/JXz0+NN9KzKCToAYsfQby6c+eG3Pof5nVKfa+6Jp2bvM8oU
NEaHcMrpr7xohLd85t1bH6c+VA/Gtc3WcWGHWBHYm8n/U9/pkvE61rXKtBReM5mW
A6UFjIyGefWSQZb313+CKVWAwclRaW2INr7Cvog8FFH0sqVJpP+U2/U8TLJjAPdw
X/ofDBxEfuhucvXmb+jTj63iCTUk4zap8W36upbqQO2wo/2vf3I5FkB0u70uW3gQ
Z/2+KLMyhDeFI/eFbk228qpqLykyAO3E0Fv5F83fj20xn3sFmo3rnT5uf7EXdMOu
dStddZILa6hLZ/uAQSaUueF+0Ji3KuBtnLUZtTqG3/y4K49QcUsKCgYft8s93o0u
5Wh8dqcEBEmmxSBDRJBePiXkx7JyrNdsbWmWu2qwsCjVrUH5/ZCTGoigLxP5h41D
0oV9YbtQHmKC2Ls0zYIUMX0odFta3dFhYTKB9hQLk3MF2d2yKrb5Eu4caDwVk6Wu
q8AX7R9r49/DiE3ftLtOR9uayC426ML6PohSViHu1NeSiTsAN6acRlzxg1yf3DRs
SYZb15ijGvgEPCJioLwnyZmmtGDED/tIS3/WF7VjE57XT3JUYHcX8Yu7k0oCoIib
9S+K/YPoEMPxKYWN3H/tEiHliEmaNzt6dc/DdfIzkW8NRQlCpZB/IrTUaNjp0ylD
kqZXxri/O3vNx34FlZICKGnIVLYMaxdV2uxj20rns90eQ93OFOxvNdyY+7wFz3YF
tbGIxgGaACuYK/5za22JoitqsMgssrVgJcG2nF3xFOkeV+lIdAtxXoKNU2WlJzsk
xj/ra0ZAb7M1uLRrTDtNKwCYuzILP9LXnx4oKHF4TQe1PnsEhpjOUPM9BdeRmArM
IJ+tFg3AAjDoNIBuJp1oxtpdoyXRd/etHrLD94C3kBcMkUEdaX/T8AWTXHRYcUBN
cQS5iXkDI/w023aAyfObZ9HYg3l1On7u0csVcXVNtfDh2ypwJLaovmsh3O27nGH3
dA2ciJopcSvxnjI/J1dtZLjXh6yZ2ysCMYWVQjD3C8FYg3JZDAUCVp0T7GCkSnQ4
qkiF2QwwPZzaZuY2A05Rn2ocwQIcSXGSbYLGWjq30TUjZRQ8NRzh4XDeAQHM4Wva
z72yrJOHTa12w3YlYH+LKzakaOCVxc+VEdp0F16E5z7w2O/gV5/LQNhNoxvuQ+CP
hfRN5xPVPuFoWRXf4HcwfpiIAHfARrnl+sCz/U2WCMbWl3wdlz8YINLikVgEaXkQ
NJQBeyUoVYk+fvn7lPwkJs8sFfPsEuvme5fpsAZLZL5SpSlxADzUqxqEQYCeIZ7T
yrrKycDRbU23KkXP6l0YBr4PsUcL8fqBeHDToXOaNDVY4eiZ7AwTv1PgG+o1/rta
nspbf2zvDMlke0zEZO+gRoX2PWNr27YMkiqrNcG98NQsXPo9u4Hi7ZQpY5p50rwM
H/oiGlG/QKsCxJ0+R/EJB9kGmf7Kw0OwpwJqyncFL8KFUAgiuaXNBn4XvHM3rrVT
BmsZuu4qW8fYtIg2v2Y/tvzi1RTsFwRNzmDm+JTE3BiI8g+LphEUX5ERfSnB5y1X
juUOOUL7HW6v9e5dtPSeNtgh5zx1vSvlPXxaf08rQ+vTnkMEtjJGNjeP3P7gTvoz
dHaFN4AT2j46A3O8PhtIPNAdOX9lPDmWqPdAWuiyEHssQnGKr+AI6xE4gviYJub0
S3QT6s9rHOCnS71N1hqBscpnwEmhQ52dTxxBuEKGLOy4SHOqcFSQbwLUTtptIdDb
ZNPQ4c3UJEnaLRzf7MxCwvHPmvMT8mDhx38uZ3lkAN5qYYVpFFoxKe/bwP55x367
/gDC0d8lQ6wBdFNsOFWPM1AKVrEqvh2wP9s7heDwi97UuYd9r0Ute8aaLDOWOGrR
Lcc/R9yfBd0c33Uva+8/ZiKnI2nOaTK8Cg5nfQ1EgCHlixBs+pe8v7p8K+w8wfTK
iUlWkEVNMA2gjDXnxwmBtZ14YnLhyMPM1zk2V2I3+RqDs5rAFttDt5y/2vozUEp6
rgtvbCm/R/vtFaODoJrssH40zhywTqOB8kTAmbgaavEJLbAfHtibi1cr9emjJsJE
P82SbOEIhAEr9lBhMN1diNRBAXdbRftBB4r7CTyX9nO0W/ASA6N49TH+20gS8SsW
O9BNsqmIZFd3IDXgQQ/lOuv6wJeoj8fZhRr0BcbmCwU5W+baBBeraKjQq5Go8/aG
uqhOOuzeZnLFEBpFbQ1u20ls1lvyaJwNRZU2mQyDnLENdDkXs5U6O0tHu23UmNm7
rHe3MJ0gbPTGH03NBZl08Bd05MKEX5SQ/IR/PXPpmNunBaTelyWEpF2EqcA5dlwe
fbHY9QGVTX8zz2JrlO4noZvQgXwfu6P+FLxiaTv40FlEu5fzCecd13Wgb/XMADDV
VGni8krC6kYj7jEJoHO0WiQs5y+eaG48QMbtqbQfBUCRQOjRp/9ErzWUPTy0XS43
/+QOPd/29xP58dxXD5Af3MaVIwnr5Yf+w0atT06ly5dj9njLQ1eMnihBKcywtK3f
Cn+LDKSACGWXtjcclKPy1eugFeoFU9iwLxfxs7Tn5gC/zwwD/uJNI9QrEg+jhJeQ
09n3F40zrL7fLnUObVgJQOdz810i4beT+WyUBl4lerNfkvCGYZy9MixmhsQS5zNA
FDhsSzDyceb69/1RNNNIYp9bNasahYpUAfZMdfaanKLGARbaKKfcBbgl9D2hQBak
ITKUjfy4McEghEDBOpgZVSF6P9eXzhXRT6axcZCspGOmReJBioiCZveikUS8xoVT
dMszfE9lcFKmHMCtrlbn4iJR6sM/RldqxrF+yJ1xP97stzzOcoDzDDt6vxj4a5kD
d+Jkhk8nfSCG1vKBca5V+rcO2/uN2tII1LPecouc3WaTQgkLgFWOXsWqM5DHAZsX
KsGiyccuYS24L0eZYxIm63vuGid/PSbncxJ+kalEhGKOAdDwSscHZq69CCz2SKUc
Rm3BIwLEbDjtYryKU1dQLNrMLRzWNlf5iDlr3XbzifUi1w/WzzNlvdEIxjEL4Kom
Dm8HCYYqvIh3KAjo2qr0ifDfsLw/r9YjfUCFzFoJfJLGMMK5+ZpQVF7DFEyJq8hK
eDaYNQGS/Gvq3gkPprD/0vok8Q/YlaJhSjZ2nEN1C1sIylrqBCKFLRVFMkvYjGsO
TKKIPvyDehQGwu2iKlFRaictCpamVps1yOtR7NEgPb7My7+YWEyYOuhXDkdj47vK
ABlCfCsifObebgs1lRMhmkDf9fa6yNZoM/YGb6siiB43XykumgbyJyoOw7qliHNW
/s+qMmGbBw39GxBmBSwyCnZA23/3gt482kPzPs6zfXvZSCAKrxYLkQAhfDxfUb/6
LQuhnp6cEsD8kIu3MFeYCaLOtPgxrN6qd6StZ0M1Gb/EKjKcl6nuUaTnLSN9tKNe
YiQkdk30S80Iyvs9BuEkUXKnEcSs4a1FSmFuMjDvV7CiROs+FvLwYCmCpPvV1Xk4
VRhaTwx3bj7OkpSZq7jMGdBl/Rtp/QV40fcrM1BJF68fZ4PF8rnCkdTlQuQAqlvA
KXX1GeX8QkCTJR+AhDAJQQFtLPzia5V2qK+XeMfdbB2Mrlq4h68v9SQUq3P80PfP
gbYpga0KXcSmWHc47lCNOJT6JTHVqv5JPXz5G+ALIp0+PCiLNIs3pL0fSW0yiiJ+
Fj1iqPtyqwe+s9UQ6/7jEJS5Dh2xQ1zpb+M6LrvyvCd9LvbT4/PPGexJrz3LAQu8
IKYR8sbBuw+0oqhp/JH4Tupm30baaJ4Lq/p+Qwrfc7pOqkRmmeLvOw1AFanN2RjJ
OSj419ZUU1H/d9MSa+oW+Hm7OgR0BUKYTyCjG2uLxAz9LR//oJDFzZTYtAY0X0RG
WfoNA5Y8L19hGGRftZVbIdZqrMUS0w1vHIV6BUXW5TpHHV0AfCrI+L7J1ithKw6r
49oCqP5PVwS92mrGO5suIdlip6KIIKpTotwsKos/spQG5NYeWQoiRcE0hNh3+Mze
nHXGyEtacQAVKRibNfHiswsmC8qV8q03/vbNqbnjeVyQbnwEFnqzFie751G9Aid3
i3FdQ7n6e35n8fRaAD3CNtVq+okYnd84pIYoORAkmdVALSI2Lv2jkGgS84f9kbv6
Fwvq4WIC6Ky/Gmf0YrbKxjzRsKNYgVAVnLBAvit+hsYypG/2bW3p4y8ahUsmpIZ9
WHx+Q232+CXbp59ESHFzo4VYP7G2ihG78EftYuW728s2qe2yk5mpZQafcSjK/fFp
bF0AFPUTrKMJIFOC/zlItKNcWSXNNeGytGO8WpcS+AWjiavSjmEb+hQoECdCB8bj
2qhFaYHQlTAB8W9HDuH1AKnBQRcpLY1mIYgLReP6TLN3OgAP04TIuEZqLifBO48P
ZAwep7Dpzwr7nNxMJmwIVlynxv+jQV1TXbCA5hlKaaxhBbbdlD7yOLcqXHBcIccT
zFzfSJg2HkGB1dzx0dUZwyqPo5K7lgUQeWAK1XOma1m9OwpmHjgxxQ9dSze++ftU
w23T4KiPTPlPc5i9KSdwce8ucundqU0xei32nt+ov1DgjYRtduJTv8d0dyY7GXqS
6t8v1ADorNJf3xKb8f6J8GqJWSyjomPeZbheYsKNC3XEXW39ZtOnLCXqJxF0TL3b
G95PEdjlaSznGcUSltJWwyFmScX13M4w4YaE+beGrjfH5f+5Te75RbGCmHVk/cWf
mMtNAfadoguzq+ulZM16hKOqZFnb691UB0UzUYLelfj1G7vJuMvqRX6vSXsyJRaX
esIb1u4IV7yyRxkfh0889iLHmTWvhOMj/3GXRCA4GLHaGm3vH8sJOlONRFQFtPQM
y0PNWHqvHtYXxbU3IX/IvI1UQFTPgVF4j7kg2rHLf6ULKlR5jrGrkQqB8rBQwTjh
wlbFsYmfI06ZU0yuZO5ow6Qop4Ig4tJDIzjKG6UKKOtpqK7iCkof7CzgjaWaNpTC
xoIOtWxkspWLs+jnXktKei2+27SnIHJxPDxyuVPvpU0QUXRcRzlSBf7B3UDBMQ43
HQUfy9+JONApMJF0HNS8ZV/yDRey9FAnHefXfPCCUSz53yRM2Xm+c0WdKn3Mby98
5H9PRrGXu8kVDpwKfrv94rTpao0zhUpnuTAewNQst2YA53EUjEWcxUuFY3XRRJue
9/ThF+46XvTVRqXZxlU7nAQa5+fPXQWKe8Bg9sxrOetsLdGfX6NnS9cE4PYnvECs
uvcSurz+7LrYrzW0ofYfgHn16zAwrY53Ne+CIz1BZ2qcwIJ5b40TgVDEjE+7BpvI
fpvYXmbEMfjhknalKy/3EPBlJoQG5OGNbeMbvfRph4duIjto0xpsp8Rn90HFYuDD
wnOCRI+Br/UUjVle5UmIWKnU7KAN7lopcf/q5j8oO83shCFCze2i7UIqlw+eeIX2
WHk2JwHu5XxV9Kry7rkpy4Vk7+MCCRlMZ61NsxfQrlsdq7n+FnOf4zyJTPmUOmOt
BpaPvPmDpFMQ6Ie4XvOGsZedrMgWuVWcVPAGku4NupFV1FNODfu06xQ1pWxgS+r7
xHTMuR+pssPJRj/RRarsFXiXRL6flPMmIM3rVGBrcd+nMOyTtoPbhU8jAi9mW3lG
wCZhzCgWEZhN8iujVfWJytX0kZ5g4ZuTeHdvF2SUFewWu7KC1sfK4zGR3Q0T4hhw
2PRwXzi5oHMbKTg8ITRcGqc/roUG6EX5XpR7x0nDKgD0VObv/m45+YV3yvMxUixA
6THCTC2+nl7O2ZnFlgCgveM483xuHtf7hqYFtECxhoFht27m6dlw0OLZoCLSBDe0
ci+tCZrwwRChcD791zZbqoQE7jAjSEmMKv0zvhDmeyobD/JJiJBN2Gxphcc0YaJm
I20TFTvLYlvoSYvDMGNorEPNkNBXZfg1/+kffk64Lg/HgGFG/JEZjcpjj42sdCjG
R8+5Ay+WIeYQj2+dqlWgta3IgCRHIxrt/rREH+WUlnU34QjooTXhmf3PHQG6KoLm
yXoLI9QYSrHK9gYIpoKyPVGHHgnTMRz7b+k60appBWcn53VY2uUqrEsrismiJU7K
DPnR0mlhFAuIQPTs2XJ2hyXeEKR5ZPWTfUFzf4Tn1vY/Zar7Ut5AMC20GqAsZwVK
PuYNqZNG0sXw99gMiI2mROg8wmJGcsNNacfrICipnDI8h17TpThZIF+4YDQvlkvj
+DpAgjH7YjkvbTAKHPbWWyTS7spSlrX+dawrallh2ogB/lQtdgqv1Z1Ftla9gNMq
yJlhnLAbYJy6lSv4zuqxV4ACGRhBOcS4rk6smUA0weXU9EpXosRUv+brySXTvZD5
NOymFepqdva9OAk1FCxy3Pi15aDoLDnAVTxly85iWq41oMH/c975QexhzjHuMR7M
zXgFLVmLrK4PuQadeFz2LipgSI2cyIT4a+yFTR3u9g56k8JBSVC/YLcwqBqDpb30
q52380t3rcxWzxGwLQVdBaz5ALB/oM1Gbz5yUbbIwwIV6oFOkBlTvEq2uZIBVXE1
ZdvCyjkuARAFPJiE5Rs4dletbPJ1+nlhtzE39fkUYqw7lidQhcBAXH0yj3nIXfQP
w5YW1md/3BSVM0q2iTCFEOMd0fGQMnFj0l8Nxy+pUd8OsOM24MXAfo1SbzhjI26i
H5QccOfuxutlmLSzLU0rWH851s4xjDVfuL5dbC7mXWkg3yD3/DxTtv3oWjvcXSMc
5EkHngeNVbJMBFQX5xFOMjIevlaCaFtsUz2V9I/CBdjqcRa8kii2nrWFMRfurv+B
QvYjGflecoVHr4iOpIybADjtA23aG1vEzFsrDCX8Qdw7KUdgwY+6dQtBLODNcl0h
xcZXyDu3gBLbygs9FYJwONn+CnoRbRTBY6Sr+KQ5yrdx3AsMQm27DZCjVGsKiVSc
H9smNbjyDChDOPDI8zLjbFB5Uq5Cu8W0Q4NT81+rlbpLJKwbQGGjCVo/fCsYCdIo
JUvfio4DjMZgdTsS8KUP5DbEwcmG0phgcnw0sD542uy9c/PkWe3JipKZ4kBs9Ktp
wo2Q+BVlbkwhHszfiDqNwoCcCXYRNPFypiYGexRtsgWol4D+RjUKTYi0YKzjkK7+
AfrYwniKWqHf0e71yv55CW0q8nVhL8Qz5bZJOE6zsYqFjT5LmmBYSIMn7Bkd9fjL
/5eFKS1r64KMU7b9XtFpfaF5eyY1S+L2IA4g2o1LzwE74AQOG0WGt6o3tJW7d0DE
GAKOFVcfFq/d4rRUDyBcjKI18973YwRDjDyI/6Q0I4ObKoDtKcrTREtLpI6qklSE
BCBKiJbISTxbBNoFb6GcS2Rc1QRVQdMej64rdNLk8kCYroFwLpsrAfvSc9ZVDcXA
+l1mMHXRD/ifiDnDN+mDWzFkd7qDOzFUnrQeXlqrtzu5zV/94LKIBKrVLXHJEIuU
HhPdFNCPEiuaMOMPMQOU4r9wopfGca1RtPLvxiWM7dUYi5lqFuY2Wu0ybKS+yVsK
2PEiFRhETvJAsPf2Z6+2nIJSNOeYNDmlFQnuyUN9ECCGQWUWoiFSSOv6HnaQmtEv
cx0KcXWbIvvL9b2hFi5LOVUPaTsCpyQ+xjOWhoRkZKs5i4CJGO78DkwBC9+z+rlR
soNzf3kbsO4plordN3wt8bC35ZEyirbR7bzinwLk8wxVcmbSyDnBLPVEG1CPO7R4
WCowgsIst31+mw4nZoZoDXqKovu/ZxQ1pn6AmAPKC3yQmQdy5WKKCj7SCB7f+qRu
6fqdHpUKzrtqrwaa4Y8LbAfip7G9yW6AzIrYa6rHh+nT+2pDgf+voiRNeGm3GmIO
LFPtK9g0sUVQZ6zFFQQrARuMUw4OKEYmF7zFf6GUCvHGsUvVf6pD3tOpqA2H6qxQ
WwrXO3yCjFkLRMWLe+0nDuPJ1z29NQm2Zy0RJaFMdjvt69xFN0BXCpa7+CyqMxHi
aKAl6Zd03VEY+nBi6QIJ0cQ2i8w+MPzgs+5eLU9mO2BpkS7I5jY7TFSQn40IyqUY
IZflSZX8lSGrWtg3S52TM2Uym4M3uwwJlVKfX37bRgR1E++UGoM/VL2Jk9sqf2+X
ecQsZaqv+F91lLDFm3j++1ZEhmECLzuxaQia7YyVoibVr1+i9mdcdu4G9i+G9F++
dXB9/0sipX8DcNCbtZm/opW/zMrNnye7Y5vli1CjEM+YK2RStj53feLSYgP/BrUW
R8HylYW4Xih6aU8LtkrL4BjROPvLkc/pEMh2TwZq7jGJnyXw6bAup8AZS/JQfGiT
RKeynSsf4lrJhO72RrOC7O4q7eAh1VON5+MWPZqQ24BPW20qbTOdtdoolioGAgD1
+eQihD3KXrDjNmj39HBnHpRPWu/esVGTzRH5Bg9DbDzfda1uex0WGLXLJjyhVp56
+I06YTsjh9hNYCbn7SVMwojCjm442zaoZyat9A9k8hXSwNrWjMbG2Nmcj6hpeKJx
yjHMVcXYCC4GlaoqSfSAUT+0QChoKMEu5Wzm4blgx1jp/riiKBPfw9SwYpBdpv+9
H8JlSaCMUBFFHeNIopjE3+wQyG79UVHplBfPs22T7N3iwLE25QvPwF9/Ksova1Sl
GSLfM9ohGg3DKx5C/nbbPrUbP9OCAcSCvX/cqXNMIt3XTZom8gxwGcF2Z92a0Auk
+4OO+N+gSy02hndBu+A+PzTJKbAad+xcpoibEQXUgd2RMK9pNBQfKTDGU8OYYWjt
yNUniBtPrxQeB6YR3otxKp73YP2DrF9Y/XRHRij/ZyBm4S5KikvfBM+ROoIvSYm1
NGMhX1wCaQH8gCJxBhnMalOGmlK34czK2wr6pUgqU4Aur11DxbZ9kgAoNnDz7xrR
dgyHnnEsF6Ri0XV9wp01vXYwglxDmXPLfO6eif8y9ri9ztiw6GhRBD2zig0V5ljU
/6/s3SO8WnNZp9b7DRn/bKGLrm/NM/9dqDCDqsQwG0TIAzdDIGJTzy6Q5nsiGsVy
T/usn/nzLzx9yvAU4BrZUJhc2pVckXMgX6DMuCU01T0ItQEtdNyQFKCzUDtHRSCt
KCFBncFqyY0yufBicCiApM6xvJPkvBmgQysO5qFp9tDzW7Ro+0YP8QopVi/7ND8/
HfSWTq1Zh5n7wXnpZN4qs7bPm135hjbLDOz4282v0pspsZeEHY9eQOwWc4vNdj6F
PECNhvn/pjQnOhcscIcTwsUnIhYeiB86NBWhT4YvvbEer8pdV4NhAuhvmsUzcoDN
QNz+FOwOOt/UIABwkUdyoZr+CY9Ph49Ywbn0Tw3BvrbbY5EpORbapOIMTmhZx2Wm
gUPqoJPBjwScxn23GwMCbDdWmv3am1aBUDSK5jilE8vxUs46BedalSsT717ak+UL
mWmj1oki+3MvJJWeQwNhi7GqNouSpqhbcQJFJ5rlMN0py34OH2gx1sHqvZvgH1ds
UbFXe8KwPFhi56ryOpGvENsejR4owNec+OBsdwZ3Ow/i91P7iL4bYkcV/tdphpN4
4pZ1Pu9qNzGxi83b2rV5jOnU4QwjLfqn42+8CNu/Kel0ZPAo8tGbCksvMhMEjIU5
4u/jbJT4hTrfEnctDM9kRpU81XLJ9ZRR4TPzndj/9716Rdn/tz2J0J3z8rN+mKaC
t87WICT5P539V+78lITe3m7ZhMzLuKsBkIO64Z/IG6jyOJbiLaKdp/qotS2+hyAP
aN5DbLKf61O3bJS0cm7z93sCrGR4qG4a5H68yZr9jGTQMwDnLjF0LBz4ewf6vNAn
4ERVU8uZDHZYXwynWJ3Q0O6LJDyS5w7UylpXJgIVgeYTcF6T+jJsgAK1m/oJeT9I
ToQ928KHTkk37zeRVYZD+g7kCroXxIdNScHpJeyalJveUv2bXbLVk7Zeom/Fbhp4
W+AgGGCw4QOLoO0qtdFvNfgvClg8LudqZdbvfQj2KlSMtYwcGp5SPQZhcbjWMySt
jdztXvFIaKnOmYrARpdyTzdee0d8E93uPD3rJR0i/clEIuE2ArBLaJb6lYFmXu3W
PnqTfsukyM1w6cvSro6d7zc5tVZiErCZOe9bMpEOC16zrTxveS11ss3krifJNmv+
pG9yKWMMga3yLjiwnQk8IVCvnj81ogii5TMaPheKMwzUPxg37lz0Piy0i7p2wjFO
2m9Nw84RCovAE3PdEJv0s67cvAC+v5UuaoUXtohBjAxL5HKg6GLj5g9mW95toqG9
sxctuPCYj7BYWK9ehJlh0osNGbYY/dk0muwMd6Ptk2Lp1ilmWzrKr4Yl+Fjw39cb
g7UA7hV6lriUez3qwUfDo41dO0ZkdP7HYyxWRNet3p+1X1QzrvX2ji/+zeepuCrv
hKhKxS/B/TcLC+WLoK3scyZdi/tnIeWVca7Asf68G3UjoL48TMr9fCINP0A/lkYq
8LIJs5LA3el69hzLi2Zu43BqUDcWtWhLOIhjEEuFhSWwoOhHRD0MyoDjp+mK4sX1
eD0DXUjTXOA3MUMED0pfwYBGsQ2b7hCphvn3HOOXMFry0zlrqD41HxU2+iqcH4D9
QenipT67zXqcgT/clSHZMOkLqVPIyF+4ON/E8XiRXqjNgILJeUXiMoGq2IusvM/i
IHmyCida3LSjW4WPATwljNS1hYz5FGFsDnJUZiZlJQNa48JAT0JqRRmUOu5w+Shm
/7JkDfwzXzFVcWfG3b/ZCvpj1H7BnS1ZS1GUN0XzeHzrfTEYngtwU35BCD+hsmQN
IJKCG2J09HsjUYWjRaJYsoGEYMDLRBCE2RtMO7M3HLMNeTOwL/nnW9z0zMWt/OLf
Xj2VemgeB85ExSzOdMGy8tvgvrnWg3T3/lfKbII4bmuGtd7UyBKZd354M/6oQwuo
kJJGpPFa9h4zJc4jnkXF6Y0gixILm0W6sLmRT/D5PXlrC5Sl8Mus1hsh9T7JJcF4
BbZfUH4upVxKsyshR9eILNykJhRlN7NGHQFNBi5zyIogKxS9Qn/zXEfYKzcdzF0H
NBuk2wcPPXjPHgo7z4l2D/z8TVWroXUbQbFB5dWTdle38xO6q4KdkRuFEM00wy7k
nu03XkNBkaYHeeU7Cw7e5dVEhl6JAEi8endoepk0RGmypCPrEgBkaqtP1+K2BCRu
AwE3HSYbU0u2Qp0UQrph6EjZ/gYuALRPuo0LmkX8jcMBjF4ynE1wZZM7WOohuQu9
w2ZhGVQw9qvNpPwEtGoSsNb3esRVBoC8POk3WD+2N9c/urlIeGnwi2JBheLJgWoW
LjurWbbX3YFAAXvVSlOVs2yfuI2EEP16p3dAHOOAVj6ZV57eXN1iziTJ3LHJMOKc
w3DsIaic+lpQuIyNNAZTTvkXZPoItqvV8MxzfF9lXr+xTFlg0iW07E92oAgPjmw9
cdIIFPeMqF7rMdT9QMcZeRieL2M9gtueCEFaovi+iXyImroq5lak+5FQnw2dzkNV
7BR/UOOihGvwpT1oE/1bsCoYDjF2iA5w42GVGqGe0lNjl9aAK33dwKAwljo+OaMm
+cCRbVSoScawql1zjZK2tdMBqDokgz2tLjmS7BXkM8JuU4hOEUCCw/GHUowShjDD
P1HQDi1kCh6jn8Pqsi2wBiOpVsoEJa4a9b9g47kE75DPQDXViCp+3aAMWSO+bS9S
zUUXaYGRcEdkofOjuceeSkrmXxfBH8NF7CGwSAJOxA9VzroW350hyaP8fWcCNixi
cN1Foej5xKF25xt/XWr3szl54Ak4akgzApdd7KvmFvJpEzpWYAMJVPGmlxJwZbL+
uKnxkgPr23Ii714oNBKxZaJetFrPjaol4YaSY24iw3C6X1X7L60cpu0E9Yb46Vs7
Qqit3yoOnyq/fgJxGrnP+SpQXKKnVW0c+WZ4R7b91jwxesSL/juZR/5SAVH0dZUO
Je5UlQKlE0TEF8Rgq2v6+aqgShg0SBkqLQWtrrCX6kfOA4b9qtE/ASotLuuiDb13
zFysbIH4ngvKkfaLSahUtZhVKuaftghY+BZJiy/h9FM1K85scMWkodjeR3jCJHac
tPLj0rm7sSWpat6QHej0tYkZv3K613aLcvpC951Fw6JVGnxXsRAJB3bUtolTUxDr
A8BxpNXbRG12YLBGKHiFE5Xu1oxEEUssBwF18rDRxBCiX15eIUY22VUwLS+9WfdH
/3456nXJ6//UAuXlpGhGLH60WlSUjNXJFVFWi3MuG7SzdRs1t2SSMdXoyM4DjDvA
DwRZYAXW8iIvZgLhNYlbQDW3qUhy1LeWnQy+fH0QzjPtXYw66JlD9Ao4vr3HvO92
ox+1ocqghAVcdL0XyoydvruU6gJKQ8Vvn0F08VCEIrpU5//qQVowD7+S4jc9wZ/C
MrSUvIk/e7dLOpOW57QBXJSDvqIY7hCWdvQpu4LEEYPVdcTn9w1C1iLR0M5Me/Dl
RIajfF4sre+ARuG4QEBDGH5dsoelO3kkU+1kPbztcUIE/8TLHkXdI5G7XtifqIaW
URIdtJL1lX5+IW8fn6P5LRjcmUBFTRf0o8Fbq8Sg4P29H3rl2VrDBx0dw3ya6czK
ocVBeFvcVMxqFtzWZmIHV85UytSnz5fe2cYmlKeQQEA5tIZCH3WfdPgOxELLyBfP
ShR8+iWDR8PYpHrIiczDr2//IN1Y0eYXZgjXWUjelmuWZT+JfIVTqkfSf+heJ80b
B4+YApybmSoJmqWr5yGgSYpSfdPfZc6BoYEwOr8Bl4z0wEmrbQUkJyHIpsnm7zTy
VUdInJ04I7smk5TVqwddbgp0D12S/YDegXo+OP4VwWM8RAhUJQ2AY0iNsxKLBT8f
EMd1DZ3B3m3vC9oZr+V1+RALM+EWd2q4GaxScfTBObF5w39Y6hndZqgTZlU2plwN
TI/8dDayUa91rEw1BmU5v6ceD+UR20C++BirsA9gKHpbP/eZtUXqB/B7Dds6C/Dx
Nh8GP1TqkxVedNajwB3dhmLx3IKL1EzQEYlKBC/PEu667T9iPEVrssvFVaFl53vw
jaq7jKnehCo3BLxhPf/KhKQUM3SAULViTVhr0kqB9q3BAnCfneOnfrGQWkWUZt3W
ybVxeEXwAhnmEdrVx/JckHJkCQGLEDyR/XXJr64gVw38ycptT4qHhJz55zgg+eH7
xm5IDaDIXTyjXHO7DtrcqPg7ocVUbRosCI/YMmCJ8kMpmLgmDErwKx0YdpNVjD1B
UVbgRrz/QH+/qhSzd/zwduuFfjbbg+l6dYkGSJg3WMG/eQQf7+gSWA05UAaMGpR2
cdUPS89cJpaAVHf90QFpz+Uwd4gfxVStocpmgRF/3tRxVy3Kzv+O0mkmy78o/xwh
oA/A5WcyeC4joGLzf9cAEi7o9JBwQmllNdchwpWBDIfYT7DqXj1LR+bUJtY5EIwg
yntj1WiIDoeqNH5YOdmW4kjO5gKlGxBj2O7u1ddPUAav4O8Rqi9JS2xXeI6Qz3W4
nbuszmYRgM0jN0ChBR5ArWJHnGbUofrys06HwkPNBhCY6a0RBTZoP5PyoPruccVZ
NQH0/XIljslaNFnNw/jIP3NGnBJXjiTZEfUpakQRQvTUpF4GM9HnstSTxkdNdOiJ
dJAPXZ/ZtHVnXxNNBhu1EaPtmwj0UIvDk7TdXePMFMoVbCvwBYMzO1UdB4PLhgrn
aS7jjI4KZHiPvSeyaB6LQ27dpP/Ts/XHu2U+g4xvy90KeKE8U5PiyjVTeqnlvwcu
KciFPK4nnx/9nYfClfjMcB1imfJEOW+HAPjg2D2GTQK6sTSwEdPE9Xb5cIGjCY2M
gLPg1kbU8iqt+gXZF6MMrs6DSefR+E6dNE4sOC/pU0cJCshpyTVnEgDJAW4OKfXr
t4j1uNgRg3jcEat8MWQFbo99TNeU5XNq2cT55Ruf2SI6tqmRLthcEWLiMqNLn61Y
PE1hUWTPT8eNbiljEIMhtETG6kH2/0lBWEvOKu1rru+48TO7T1o0y5vEKJmkRyfL
RcliIus5lmfFpniw7pOLX1fKdjYWaHco6EYzodBU19Acc+MaZVVv2l1Toc7YMcgv
m4LX2WUiBnuTaosHZsyKai4KYCJdcdNwQ0QYEwa/tdtKoH3G8KolGFHgqYYX+/M+
ZHrK80/UDLtm5eNNB1t4iF3V6jGWDrmLyZ3MVtcKtlDoBZ7Rc6UyjcCT8RnPUKqn
PNHSENYaGisVVdJujjP81g7WiRJMO0i3EzaKEDwZ5zB80gWFiemJBQfoEjmB510V
acuqJKkxaiot61WO0upRDp/Y/QUnyKxed3AO2QosLZfrxMVWpvN5qGM0cBoyIWA1
dv/No05TrWdOIcL8zybzu8x/28lcTusiQnhbgoUm6DEqopbEWH9gZy0zA87AtgEl
+6iFuX0hscRV3DyCp45KjeKxLGzeyQpsuHDKncRrG5mVt+s9hCo53r7uiWsHPdx+
sceNHKxLs4699DnOGll4eWo63w44E2IWdK7r5TivcDwgvDQE0fX3ZLUNNqapK/An
0fJ4/dLrQZCd/pJIiHmpFiqLm/OQwmcGMeI/+ptfhmDKHfYFT71PsSEDTkJB3k3+
616Dv97SNZ07J1TeAZvZzEkAKtbvjcNkROMbEWxSqRT12SbnWFhuwnvcdHOIhsrA
G+/8SCBDayVCEhfdcBaKk+Nm/U70En9lF10MVtFH5n2JA3ZZlOnVyyoaha/zWXP+
lJduVdUVnnuuQILH0hYG8F5CKT8qGG/8paRG03ktV3jmtl6p0pmz4x0lrRoDDDxY
GCpdTDO3ISNyYrhnp4UGuU/VocmImCvL+ehEQB1Arf6Gaw3uj8cVGYXazsG9LQr2
GFofwyeJ3icrYyDL+4xYF52onT4JI+86ZtQJIF8r/DlAdLN6R9nT2fh2WFUXKt1f
1wwj8C7Z+8+XFJjjhYYJuqlVTTwZk8u4R3/bjO4WGiiqFwq18TE8+FzdXvUExbGn
YriMdlNpwmrJ4NUvV4FkjioQ+JKf2+yvQIqIE2UBBMsk+B1HmgsJJXiiEnDSf+uJ
A6FY12phbPCS2y7TVTosWFEll2hlRr88zhEWLGQLqSBGXph+EDMImDK/nb14QL/s
69oc/RjIYo5cVFsQmN5O3lO8LOMxNpEM69tDLwQF0UAS7XyVMwP7lt9ivf0KNYo6
lNgj7683SN7bCsvIEmpx4uh9xlFr02F/MHqUzo4t5xXPLkbYKQ3S/DBFfdelvc/J
zTe753WaxXDym34oiUlf6riBo9LYxszlJR+dmHw6ft5HhrrxfbdcUitfVo0sIE32
tlYcPWENt/nJ2+I1rineJDlRISM0Htr+qid38Ludk3v35tuSP2563qqCFUwRAPPa
LjYouBozI+p4ZjeInsb7Z2s/7z47mZM0baospZbYcMeQxDfAGzm9KrD59ikssUcr
QYT/fUJY+4EWaY1cHdJNtp6MMgJcW83xjzJw8GwSf6wm3E4HAZN6e2zVBsQmkEVK
JIiZiycx6VqurEdD7N+TrwcrFGA8vgTO1g3VAtWKVKz+1MNJ8S+xHOot35OzEI1D
uaFJrKNE9PFeRLcQ6CvIU3BxmvUWuiRdAfAkSguD3bjrW2/qH6816PzNFUcVJE9A
NBqgXLrOBV3YNnmxwkRBgpCLa5X2tydImC3n99BH0h9zTPePslktWPkA1TsRiWvE
KDCYUj1r5ET6jUUUustNKO7EnX75BeYdZiuuijUsAAkEwiBvehRvJIK9+T/Fcnx6
foSJfhAshYhSpQhMtXDzcll8eLyHWG9ivv29NfkYA55RGSdUPsyfr+zNwmUJYPWt
4IY+M19W9EY1v/eDwsbjbq4gTgpE3JdrhVGqjC8WWCGEcVp8dnaeR+XVL3HLK6FB
1gqRrp+/NR1yBpr5Qup+Txhh5Su63yVV4g4NoDSqdk66AAm/AL2zn/WqH7NJMQVc
TWnUovz8hgtNRzc/JVJViEMG8ZsiJGmc1QfB1kSSJjZPAzzxroWSeaeg53Ps5CM2
1/sRVJb6PXfATJY0FLX6mY0Gh6wTCtL0PDsn04vaNVOkZJmJsmBrhrhLW/hq2Tx1
5COqmyS2wp+8MMoQ0OpVD/2S2fbqr47OMSRhW9mDjB/eGnRqm8vKoY+HrJn274o3
LsKL9c50O0hELdJvtm4Fqn/AjELJRqQErzDxAYvi1GrMrGoZtHet2w2YwcIcvkCW
RsRAouRXiKROhZeRsoV9amyLzMUrgH7SzCAosZVGXwcsyKnwfW25YCeKROxPedkP
GdBFCM4xEbW+3JA+kfypAOSY5OHEn8nhWlFyS9NBQhlNpV9vpXA2lwQo4f2tRRLR
JlBeqD00BjccJ2fjRI2yAr03MlcPkCzIrjV0IfDTLKttn9MbC5cJTDsnJBbIDDCj
8g/jR1fURkMfoSczqnn8rBMij3zFMbSMn1FfqipMcDqULZL/s1z+QSpN/ZGMXfWq
u9C/v2IeAT5tnsfGywVkyRZmA1Fmqj6HX67QDBDmu4kLsgrcHjtYrAG9iOrUXatL
gosjJAjUUB2KE2P5kPj/egK4G96ij2dzBZLkZaGpQDj0rVs+Ue1RGKGkJw3SH8oA
JZk4gOeveQAvtxS4nuPpPkx5VdOEPNSMhFdaesmBKw9jNbjxuR+Xg6PNyTjcgn34
86dvThutGsdvqFhPDCaP//NKTzdFOVfO+wK416rdzUdAnXifmV3WhXMig0ZCgmLK
v119Oi2B0WD6+73Vwm6IofAUWCbvVSLrVEDWconIZcqlu8SlmErMIsbEcaAvgA68
q3136E4pliRoROYlds09R6CDCUZxoFFGG3NQra+s5J15Cf6Wxi8KoxWvfoVqPvyp
0E5LBEBdn3u9vtC6RDIvyBICTs/g8cgoUhSBJiqGVmDCod7Y4SLZN1l7m4Q5FCHg
UembhQysYD/v2/AuJG56+zW/uyfQdylgXtKn5NZpNJr1voYIgcejyqr4qDYx/BvR
O94dUij4zYUylqpl9YkVGFuS/4RQ9aSCow9KHymMwj23gzzWsMqjmv3PX1YNq46c
1mMDVev1mJlj6j2xqB25o//SpVRqVdUqL04l8UcYXDtmneQeYsv9noycG5/wQ8BR
yhue4StGZPoZuXSlCRZrDad/tr7Jj+CYtacktxtlmGBhgiwUFcVIDKGidkKSKeLk
N5pImv3qMaA3UtlSg11GOUnBzwQ94tT60QkYTU4xGQZbK8cZQemmd/Io1uSbQGdT
OnTWZELT928Ty5+qd2WCkJDIf+1jpScAV732vQ0OM+htGdP+Qx5NXsV9pWCshnMs
rFs8ihYW398dbEwDfx8TWc0tTWumr6bOtIyfHjNidl+kG9lnGJZt2mcvei1nKmRq
kEjDuR2BD5YNrLDzJslsNNtSgfenBmLboHgtPo8MMxEgKprj0GxzKYVJfeEFM2z3
cOhxxlyfC+OIdRqX+zrZzPCrnIGickrdUs3A+hgza/v2YGHCIzMY3N30kE93/iQD
c9uIdvwMtxHFKIpvs3yAD+LkyikkKHKrdOf4N4e/AcruAQksF3I+xx7euLQDXl8g
nAKm+PZIE45nhkqCQjFcCE5olq+ZSTrFrk3Q5BIkXPWbeMeb6SvffUSHeoGNV3Br
O8LprvlV/lHIfu4MZHbqXBSKVmP3ndFHe/pc0Pdtl0ha/eJx6qWXk6EhY61LT+G/
Jbqs1DUwYom07t8Zb33JWTHxRLpWZqSRdxQU0tJJxzn8bqpkyvLhbxpF6JZDjiS3
s828L8lHfQISn2JRjPxkH4IWCuLDc5rCfCwyYdJji8X7CvY/Yz2EzPybe5s03FLH
yIDJexEpe0g43Ef/m8tZCqIFFAEAd6GR7GzhYnW5OsTaFod4EJi+FbZoiD2iN3CI
0bSc7RX7/jxq4bp12ORFFhKU2sCZWQmSokQlZuYJt+wf4+oM/PYfbctqTvH21YbD
byo30uBaDX4jzMD42qq1D0Ru4ikz6GA0i3T5p7KHZIlclSr0kwgqCALI88r+DxCj
B27HWfVBXwrTzC6sz12jEChHF36ZxgxA26wSzfhyXcTio4c6//F0szpXCjrTb9tY
8al+GY3BQQSBOQ7d5DaNBVW1Ee7Ujs+kyAddA+osmM2xkyAH7JAcZJOfy/xuDVeZ
oN8tp0yb/r9A5pqSQsdsPvqzED+ex1FMC56J24hKmSzYEnVMyvgzfujmxrY9Nf2f
ErqYvcBDJ/3vdwMq4OB9can4jLbuSRpfFGuuvgR7d1WZcQYFd7xZAE6GjvYJX2Kr
hYZrA7lKcUb5VMKciCtnsGmlltFQ/J72fQDGp3x2Bc8hg3rmVI+uQvFSlBaPHSP+
EyyAgRA9Hsx5TFCCXzwMOAJWoCcIX6l82QRQmEM3kOXDHASnTyeJfdOkw+oke3gF
IrkUOvcz5Uxi0Jjv56gzeiVx/sc5MGluOss8N9VZ5gwaQ7sD1xIhT5dOmJ5xgC3A
cnAzMRuiGnY+lNRj7fe4W6JqXJo2OLQglkNTzh+hQS93O23ivVBeZhW1JD9kvbHN
tWx1ZJPWLn8U8BCMunqxaYEkXdXSv3Jx80kbQMOTy4YB17nUWgy9kMcD93/t+6Cf
iCbPxJjKDkX9kvQ9sdRlX/JJYel68b3DGmgZ7CG+1hOcSNOcjM6zb+w396VwEjeU
8JfR0q7zSSCxqn5Mlg4WT0kCGBHYp5LQafWmGYHfDLznt+70u1ra0WyECjmsSM6F
GQVXbt7Z/xrRzog0cn7EviL8pHL+W9mwuelKJ8JtG5uwleD3/OaMh6EySOSAAPtc
Gc/UDheelzullSa6lQudOtU3ezaJ60+nRJovFrVLjmmEZQLx2at2h4c8iHhhXjUA
bsX44oGqHVYw5iiiPyxQA7tozpbqfritymZrnlxsJltETNcTXfjq8mhkrPiHihcP
JnqVRpx+5KJ4naDWgLxZtB4vD0XkpOwfmBwOh9pcSL23jnKcKT8reYppw59s69ig
9lX+ro5a5lE6ZOyARhZxwovbTtczyXEvUwh5TBTE0CIE5AAfW9SfgOSsF64N/l03
YQjLms3OR8miRX8PeNTYzi5DPOOeZUu4rKJLSwbjVAEUz4DtsxQhCDJvKk93/rmb
ZLQazRQfvOAp0Enjw46TVUgnL77r8M/mSa/6iOHA8g8aHeM+RMMsFh0RXRmcijvu
prtHVf1+SFKOWzna8S1rOwmrar6p/Ad5mx7yJvtZltBbctwCY8QN/a1iNPM9PWRa
0KWUViPhNnaxmGGTExEjt0Sn7OuiE4YffRH8JSyrDEBlr1go3umtEqX1XttAudhE
dSyHHIyKB4E4YSv4ug18HNdil3hEivTN7s5dayUrz0czAe7el8BhVYKquHX6zY7C
Ub/XVnwD7t0ywz6SNKhYxXpsorYkvy8H9G4qUGtVWRt9miEaTCXK96vgjIGr0eG5
w1ecRdUEDzqiYlL9f+PQo/LHj5MS9q1i6aLPPXyxfluP8U2RBlkJ553LDZsnFyNc
WDcxVvudNKLj6eBRNWJbwG7KMZ722cXW9vH3rV48XWdzUiVnz7LZkio5U85qPW/I
xshg097vhhkx82B0v+hHBVWGYIhfQBPOKjfwRlWuuNUG59b9Muvw8v5m6Gg0WdtD
xjHxqJlH6fQ0qSuuiDbraX4+TWsEeeuEqNTenjVALwnNWsskPNDHfltKg6ruTCP4
pBMOQl7yvviM102BCPoWHp4ZuUWTQK9deCVEv5b0GS3t+0g6RNMwwxfWx3XNHpj0
mu5wxkCiL6Ntu3iU8vY9xOVuWBH53UhNc3Cre9Y0qLlM886s5lg5uYt9GpB9X2JU
2+NABYCrTcMoPZc8FC4Tpnz495IePUus5QvZeewZZK//iA8t/82iDizau+EbAiLY
wqKVZ+TdOzWVV1rUpjuAt2fZicH40/i4hw1IsUut8KGmSB2OyvT/3xcyxrpNxzuL
d88UKsKpdtZswD/jI8O+iA8EESRxc1XTFkOPdZQMBPrdcaUS+AXgdLX2y9iuiATP
eErvN/ysL41YXYFeqeli1/LPMpOKFHR8vE8HFect17/R140piyxqRrxdNE721Y9+
iZSNh8+GLtjPma2KMPDigMLi8XzG8Kqh5gog+KH3nszozeVuapT4cb80XeK1EZV8
ZmHruhzEzgEkwpxMknpMnN9wmnDRuX/6KTo69FJUmbbiZ1UndjpIhCQgNxdoKg+x
A3EmkyC0CxgmGKk75RMdukrhCnvzDhVfOEjLkhdN8TKFSXIs8+LRcD+rBM3fl0v1
ELWNm3ydpWt38ur4IEsadP8Ngcgoq6NDR1IBQsFhFkIcrcB8DoHjgmKMafZgGqqK
6zsF5HFyen9m3UcSjDFbQ/Dy9tJ75xYRzhwgyVNMgM5YRyJ+VMw9CrS32QN42BFc
KnRW3SBKX4oaBFhwtAw5Zi35U2Iz31O5CV8hvBb7meR66MvlX6bPBisUbqxdtQK4
MMwUIOM1lQIogvU0sptKtzh2CPUJ45CiVAYDg1YDhdqgNPx+Tgr+T08xgazG4noQ
rv69DB2VxXS1OJ2UjFcOXN9OCCZNdy3XI0D2W+dsmtgYXAU/5RJ0KXOp1zbwgsa7
QdF2o7iZ8ejxCa5u1etmYnGkpgn7H8cFEOiZ7J0QaBT4NvWI2u6fkSVQn5Hi10lm
YGlb+FKarNCKjD4JjvW8GH4C6rnhG7B0otpOpWnMKrX+n3xapoa/EBk2ggH8nQTQ
s1/VKvc5UU76eXStODgXegrTaN0GI1mylU5/QIEOebzsZkWMDly5bGUAIReew+LW
6Pw5rPT6cq0ahcaFjLHkYOoV5iZsMu/H+IJh1BtQD/A0uvSSbt5EhOYmQp20qiCv
AxhBDkGSxCS/7s/G4tg1vdCd4/j28iX0DjsuzAwafxMWazUFEF0C6ytAnPVBytUe
GU94lZ/ouIFQ3bTnA7E6QKiv4mqR/Q8NgVqJ4sedZhn4Fss5oTYDWO7IHQSANbYE
kaGxgWwnfD1TRhy1E25ahgdLc4LhKUaqDrni/H2V4aRaKr7L0bVvfC79tEc8s3Vj
u0pSgDTJnUw9eXIMJlmUNzt6MJ4/L5c/yxuEFCdOdWpjf6p7EJ9hBOG/xr7h5F/g
KrHE2TIQyvMomC76WE1HwG+t1gQsS/VhBe42V1S/Q3cmHSlawDThz0XKj4rEUQp4
KC+/THALmQEN/pZk/OsabVNQoreeLuOZFNkkVUuc1MFMWZELCq0FEWrV/KQ6AvDO
/kqMDcAACmMe3+l0+VmNlGqZUPRRL+kbprUuITn9e01eOOua+Rf32IRVo4QuebjK
5ZCV1w2gSLKo4j4x8wDRu+ksotGHREHC4R4Rk8pk0FoSusA/cdtQ+giKTDEaizlm
/lxTk2o5st432xipCj7DmcBkqvxFXrLJDrbwmTfxhbQSzE+g+KlRC2/8wpX0xt8l
yl/pjsMVLukR6lEWK/ZRDDHpuSxWUEaEHzRbVmn3UiehhgaiLvL/2qkoTXygqft0
N1G9xBMyX3Dxm5JsSaEqhtFBwAcb7EhHmFgRyDzbIP1i5ZHqUaM4ZSR+pJTasMr6
qr/T2Jfx7DfZBb0Trggn3HLLRIz7l8SqcObbQznxzK72PIIw8edVGMsxDQyc+vaS
9pKnFvgsGTlKSxD5XL+fd+8GvGdAwSoVcPB7zhNq0bvxH5lsonI9xV+bTtNpCZ/S
hjjK7wszljigxUc9ICR+Y2vb0GDLR+hImXx9lA4jcp9VkozsKyIBXuUeBw7XD+Hq
dQq0GBFH5vl/JONHCS6CeaCnK3oniMi/SW+/omKNQA0LQcgqntvI03nfXb9kkawX
nm3xynylc3thUP1CfxjoXbE0svJzjnuHQehXKswVuJAcm92lr6qiWkmqH+30kivZ
5n3xy/2Zew8qxFA6LimjRbieMjEIwbdVt73kr08k7W/ZjEM531nKboTqtTdjlmAT
ndOVckswU89JKNz9/vQJdWs5TBJfKwcKcXuw8kcn25ghs+9R6G0CklmN9SSDeMT/
H6iIxvnWcDe1IfLWIYr/FQ+F0ULRYzWtdLFhmWfAhUwdQEvPZXl7lmE+4yYLdiQE
nYKDPVWUYgEtonaJ2kd8i389jHUBeI5V256SdyinVXnsbSRSLlN/UEpIzQhtcLYd
rUO1efZ1Zq6oMm3NR3iwJIe3nW50FVolzDP1unN7IDpQBgJzjM358+f4HR5peWWH
2Kfs4LX+uuKlwJFK24u7ZTw4LNX3RIyoQTsYEfbsQep4Gcl8w2WwE0boQHMMxSll
j4tO56zXxkhAotpQAJbBnlT+PcZUowUlg8Zm+7CoIKCNS7Vl34Th4mJeQrYfkH/h
WQc2/jl2ehhTmvpozdSsT0+jVV5IfWAX9vjeuiAICzY+9clFNgUHDiBBgrE5J9yM
JSCzPJHKzwXUtDONrLxeZ/a6FCWCaGKeAItYR6hlYgYJLZfD67IqdH4c5xtH7ig8
N5TSNmD0w1i3dqhf/pO8vWYj0mZGJLC9wf9nfo3sy4GAew+NP3Za4s3dE8FStZaT
JGLo1HCCjJc+pxqWAA9GuAJbWPFCmma04MJnl0xdIZfdIltyYeSxWUgUHat6szub
IgVdk2tdZwKoTVQTCH8NUtis0m/lriz2gOCoIpKy5tm+k6WNP1fEncL1vw1x5FZN
EcE+HqjR/fB8bI7kN3UB7DWZvariaDdh/h6KlBaxzX4VVjRi769TY7zna0HeTTCo
NBUPi4MLACzyOH9xKVW+gLFonPJnZl4L3I5Zpwo9gynsl1RI9NBUbGaIAZ4OpHBe
abFQtzEO/Bb+2gCb4VDLy+9ta6Ln54E1tpizu5hDXZe4FcqsVcIvesQPukThZR1W
SulynUnpC4kiVe5hysOsgrV1TLPBCU635BOS4RKlQn5BhknXl93TSt316rLgqUBF
7Hc/cUW9g8pJKd/MYMXgkuxXVlpVJJqIRlDO9pC4k2muiiWz/w4WKhy0tDnEtCnD
22asQBMYkoijYa7NMzMV/uoYNf1NwWokURk9GMQw3i3fYyIVGIQubS1ru7P2CqhX
1CsY99H+XPaejXRCtm80RnVsdTNv6eU5CvI4j/5vsLK+/P7haLrByE/eeZuIm3Qd
Fpke2rvNUbLpsqeVGhum1uX/5Wbp34kAZbK09oD5bTuzcHmTNbz3ZYUx9ieGgQ2S
qhWdG8CtEtbhsDwIyA1mCz/xDk6cRh9DWWvKtWJN5nCXymq+QtSgNxpmHqom4QOG
ufezyEeZo4ph6njXJz3g5lvkflGtV1Sf5Gvw9hG5oWt/2JT5nPSt6GoAUApUJ9FM
6v5e2tiRpAmDV9DV2d1Ivhm5Y95fWKroGk1ml7LPusCp7gfIgVw9ISFXe/sqGCqQ
9SJxhzyKM4LrnsBTHM9+qt7GHPHRohqcH90L050QVwi4u7oIEYiPUwV0yqEAeqDn
phJATms/4Cp6UWrmuUqdGi5HbYz1sekLvkykDpOTP2df/t/A03BxtwO6rmzXF1tD
m62u33fcAmUK9eqsC3W2eypu8xr4Z9GWoHmaatzMHNseAaLz1bme2NTGcq+rBJp3
tg8pt0sB3n/avR4c4hkHhIzuBNCmcHdA6wMoZj5i4TGHGPrSzcPtmUW7vRplUfC2
IuRwuj0neIIr+moQuqbRzzFkaLUad/06Oy8Xorh6WDwrT+M2dBidFWdwnNMi2Btn
dR4OycceacwVAmHeBl6P5A7U5a4nZNI+0l7kaM5Rhfmf16xiPbyfAM4eaH339eCe
V/BiS55OOzfOPsIZxYUZx8Qm1HPrlU2o7eCewxkUWM2Wj/GkOTaSS0v63xzQXKnU
utOOCIqeTvKWpxBSmPPWjJyuy+SjjDjpge6Z6dUYxHNqSvUfyW50SowTxT+wdlSG
QbIPq2OhPuHQzJ489x9evxiDryH/3RyTgzTLlxAdZocrbDfbbkNVlH9i9H+RlDBi
RY2xCiIrZLzNMglhDKC4NrPA0QWMrEsDPciqoVG7oQec4xkWVQwTqyU+QvHkZQcL
93F2PdxEqE+4DGGCfOREMrIuk7hHLupb41Q0NVujy7L1675V1d9Ji8e+HKkKSNsS
VZeWgZyBtxbev6z07bBAcVGp1rFO67Nxb4+ewhJbOnWz8Sf9U8EZ5oD0rdP1btnL
xe5bJzMpLvJuPd2BYHPYCHqZwghYgPuUwKoYDSvLufctAkm6FMtnGTUhNBjF48Q5
5h5od71okh6ETe78srYl6jWe6Zcz2N8gWfQe2S5B7AfAd4Oricv6rILseA5PA5Zn
iuu6CvD3T5wPE8rYCh3ZrWxbnb7Yhf0aFMM3GFldLsl4eoQBRc7FW67RAAoiRyPq
z/VH8THdXtN4khKITP49kJJwFCGoP6qSa+mcasXzN0rMhBQJMblZ7x5l0gklNbjc
0EUuCg3XFPKUfCmygPBZqcsUK1AifYzIm07FGmKE2a+pE7PDvSWNXJ9Qgma0WtG6
4/YfS4N2lvNQzxw7PH30WBgYwYUKXtLBG53pZ67gopvlq55UB5+xUgSq/s5+dxKr
J4nLYkOk7k3KeJocUlp92XE5t3Nupm8JrSp42jS9ho0EHrSuqoEg0fHOF8AKGMT0
VZjGsMdiiWRTj88STxzPHiHP+lp/kba8LqlZhl+WZbgOrbksTEedwfWcFF84BF23
+NskMQ/N5eerwB+wsBKGKSF58OWbloXc24bh7zU6F8xr56ktAFHEvLIS/BJNS3xx
Zo1/7bHaGCdhATG51aIaZeIawX7iXMZHyEUqcYKS4t4bYQtX9SWJoRcuOfGoafe0
oNt18NsKGBnaMkMygE37H5+6A0AXbcHgLUJiqaWwmzye/UnKQwhzAT+8h1AJKutD
wKQQ5aIiP3tiJ/H9lIrNL/+qeNA7Ctu2M2neXgecv/mE7FxtHLnXJFVxUdvC12l+
c6Sn+FqYVgiE4EbaUfI+P1Zo+/yoFZQ/fdgCu4EE5Qr4CDeIl3aJjYr4NxnpSwNG
11c0a/tj6BJAGzvpnenviTXaegBTXAZIwcSCt/8gSa78pigXXVh3L2q/e+v6wPB9
Xn2aoBcWj6NhLAqU39VUT8hTgsEEUF4ucGM7KkAVEvczyeNN+hp0KAYMGL7xwZh2
U01VvJ1JiKwEIPSqr6mZ1EivWcLBatisyxWGG02lTgHkr7+vlwj4Y0+iymEaNqxg
dMy71O2Noxoei8g3JPQs2WdUNMosh7xruH5q8BW/j4k5k21sszVmR9sxr3W6VcCO
F34erIvUKpipGPrx+GJBxyrBKuJ+vwfKzGNjDrwlTAqtjZhyx2Pps/GfYvZcPiD6
m8hIEMpC3aIY9r0VqBIwjBVtCrG6wgEdsZuHkhJxiReSMwS3g43qiJJyOUs4Ioep
KPCw3Ci6R8LO4/JE1uGqJ3TLAbetSKiM1IC8fkn4ojhvcYHhaWn47x1C7Zw2SI9W
S2T5/82HBFLWGSV4dKMVT5v0gQnKxFUAySuU7tPWznhU0y6LTk/ynjyp78Yt/LTZ
36h2SvJQeWGT8DKxNBswgGof9UhMbIG4S8Mg3gBn5a0Xxq5tG0qNbUASru71OCqg
nCFaRbPIXFonck4LIExeaGR3zvOI7ODHEAFpe2VOn341bztXj+U9pxYtJZUXK+Bs
d0wK/xSJ/s9pCuNUXEFigIGl7wAm9gzPj7n9EtxH4vTzOYhkSQc1AJLet07Aq1oM
fy/cLgLOQezavSBf5xnoK0HCehkT2GcxJxD6vLvhhTARoHMvuau2I6bO1zWy6wKD
hjuvcVpRzKq2z5DZo6YfJDIPTDDbh9N7QuDZZHkAWkyID7O8XwJ3YrzvXOwDO7Nu
+D0EQFiNcfWmBuInL9ib+m+gkZaN6fy2qcrTH6xt1sX+CG7vsgUomvQDw4MIv44b
vnRCcNPKznUcqQMm+OYGq9BP7eTLYG9rkhCg2TXD8vMx1Qoh74XMNVTjdUYLZfbh
dRGFk0QlY2nVP8jj0Nq+fTQihEVwxWraDwJHhoqzhgjhGgkzSGnQeOKO6xH+C0bk
IJF8UmvpGTZQsjGaz+wdGCzKiqwBMAtrA2cE1/iOZryZxWT+A75fDH+BxZ5Yf04g
gz15X8owXjYBsL71k++GxXcp4kmmBLXIQuLZcmz3BlT76IpJhK8KOlt+NA2B4Isn
WMXBnGH+xOFbN++jwxL1eEc/Nqal2tu1QIjtJ4a0RUd5Ddl670d6gclaumPSUXLC
4L9z9X2A5e4nRZPd0bGGMAblLRKmFr4ZKlCpBKdN0FdOy9mPwgJyDFYjlRv0DX5s
0pnO3A1PHpWP5ziOuKaeLrMuHAOkAHKEdalsMAloUAxKYTAXcxPgvYAsMgFk3DCo
0PfEUOQsUy6zD9jv1LvwHpPlDTXPiUfCuu8IO+jumYp5SklN8QAFvkH3iqkiH2Zv
mcYJY4OQe8uuBDs2Gvm3qRMqo46S19Gci26abopqTtDmOb/M2yJhRPdx4cAs5bMf
mkJULTz08u/PXj8711hfvKdau8WUnJ4mQEteG7LCL++zw2TyxgkLfFdV2uO+wVFx
CnV+O1GF0naZec4YJ+SWQYlShGMZer6w0M6EoQDt9o2NAXPwOCZ3L1Jp+GaZyn2x
etg2BxyuaRNU0TFQbarVzwqsircc4oXBUOpkATTF0af1kJxTCI/m2oheoW0tT3gu
KsK+vgNmc4HaPLAc/rRV/1THHYUdEn/6velRJHoKWyuFumOJy0RQUdWNQ42FWjkA
ifD2DbSiuG87Ub4E2mvVVC4Y0++lH+ernSWtCsCNYigGub0NA09Q0/OlVGP9thDc
21Z5mt2AP0kXc+qbt9dFFtoxNB8ecWKffOxNzS//DpU5rbM8d1An3rNdx5tXGwMN
RWcVirG89qIdND4s9Gr6/sdAM8ijcwSpg+j7PxiwOTSZ2LOXoPknnqw9zkPP05pD
ntV8LE5GX2DSi3luAgnflFeDs4OjMwWH6CdJnHFleVuOWcxcomGzIsNvZ3M+X+rt
qFfivSSvLR+Ec5rlO58pQdI16kUv5azDJkXp5J31PyIy5uadeBSAFK7n7XSN7M75
DMXc81COwpslJxrBEVt03fvzrshOByOMyyO8iTa/ijlv74lQRpc/bgSIv6JmDUy2
VELDHlODGr7RQ2xPK3UPEpAJcVyg7SK8MlQMTdhQY44CKWzkVdkiqQk6SqSFqWJr
zdzqew0JpBmGXduWfCWLWVh8iyrpyercWB4lr64/YKHvuUqXUUBBGB0xufWnAOrU
WdkLm04Vu9HjJmUTrTC+CtftzGIl0727XMEjP2+UQgwLmYb2VVmE9Kwx37YTzz3Y
yuHJOKfVyp1vQMOHTG5W/bkfgUpA1/vEnP4cz4+MYM0+dRF2kj3FMR2C7APg8XHY
evR89HuL2WAtE0zqSSR1TkJv17skQjj5jk/u5OWOWt3VPqVRecTJUXkCV2ey58BQ
948akpyJpvy+HpZOeyFLSM9XD+jheKYUFRosw5VyUoNn+I2aZAETlA1mp0UEMNZW
DuJi6dXVCvRvlf0F7L/iNehYBUflpb07es8KEEXkVoEP2Dr8qmJMvZnP92o4mBUc
aoBqkRX2ymu9CJEQfePyDp1RoVq111YtzF845MfxY8IESbw6/a5minI1GJgzQYwt
g3peSNNTebcKXmvFX7N08taYP55e2dsVTU9Xo1BCCEWSGd1J7pJVXuDxCVYMNqwC
MFzBxNsyF/NYiy8UA0vh29NJLXV/w85k5qltYZnQpwqdcrqVs7PBDLaVqTZ9cCJl
3+oGf/Z6W3ZYLcgRtTSO13VAixB26t5PBYxvM8SA/gi6xvr5KtbV1DcmaAPN6Hny
H5IsKshhAvH7+3nWKskqqxBg5/4zvfrGJAWUgQAGI+q06aQZmEQyeBzvukwUCvij
PLIP/y3O9PK/IfowpYuU6anSasLg5WRzH/6DL/HzS63svMGlcR58eHEDp/BC1Igw
gW18bybQVR6fRLnUc3ZxDQ7mutx18lguOJ8JHUwWtOXp5AqCEPHAd+cBPns3Q5VE
A7lFHNszqymuQieMUQlphCkUlv6r9Lq7Z/Lf10Js+l61YhH87rbyE/KpwZRPYeEN
gGRxyLf/9MSWuxPvJcobboHyVAxta/DUA+HHFYAAmVBkuPnQ2/RprtsEDpTwy9vs
gaOxpWPMScGvG5gUM4yMSUF6zTUN3ZzbcumclOptDcFzI6CuyvcVKd+sof7x41/3
IeFjjSUi/8QQP7bEcIs2czSgcy9x4jL8HMyjo1ndGD9uUrpBrOXeP4ASuMYHT1X6
mjhKPSjr6M5l2+ro6jmHTmH+EuHx9o827H7cm+H1gVtmX9k/wNM+iG3TTE/q4Glb
rK00i2hI346tT2KSMoSf+KkI3pcjzR46qlmT+gdTXI9r2NiVGygQOM2b4aiPBfxf
hvS+RQr14wd6/OKBpRKwxvZvVX1jGAWUDlsNgpEgl1snRvFtS/KkjDah518hp6Ap
clxyRg305QP7HqGoL/OiLF0KacLk0l7cCnsRUrN9szV2zJluULn4utEOTZH/p45m
qeJp1w9LjPQftgG2kgDDA3/B3OEuBgxdKgKL1ZDUrXKt0mfjUhH9rMp1OqJHYQcj
eoez99G+VBWrd2g1n7CkYXh/+lqaYYUpHuzjiFLM69FauJcsR1zNt290OxTwQFbY
FdOEAwt7mCo3VJh8fg6MRQ6QVzKDaiB/iypgDyH6TqwQldtki2trMiPIWgMOQntl
a4bZWVvnLFhRXWBiv5wo7gfhBWOlWbaUl+j3Gxy1rCT8DQFXFZ4LgdWMCU0EGOLo
4YnhqZVzmaP04k2E2J/hHzWPZMhgKh3bwsDuAnWs1aFxyM627DliXPsg/J3XRCrn
jDNyUoLnyS30M6RNb33urifEMpQTDgUuZhOTg+muvZSBg225Zev9kA51dypN45FX
yqA80AXWHIGJZKMeCn2FgZpJSI6Yq4FuebMeHAX/IV25yq8GcT+dmXt1MtV78u3h
NRJYSzdqTL5i5FPVb9YnlGkSd1JtUGF23vJMJDO4UWH7EwcWBcxJ9UVNze+kzTEh
bu4qan3vhkUVQyCh0lzE3pvciTdshg7Pv5DiFRkeiX4MmBGZ8CncO7fQEdqd0DD5
xGgVEc1H3PLSvyVzbY1as82/LZmwb0BW04V8CxFAigzSeXgP9DPTjev9RA7IjJyR
lj1SgKUoRUx/IKLYlfD238aFHUHW7ti5kb5Bnhu6M2zYbzIPXznG45xE+31qlJm9
Az3NcnKBOERrGwwQX6e9uysaJ0M7ULHvHTqsjcANkU9egTRckT+jsxFJ3gXvAmJn
jWaI4eW1v5hX3NA0PEyg0p1kXSQWcI606a+zRJu9lI9YP36j/hRrkGqsOv3sHdzX
46AyZaENHwvTSEzn4XKogoaLTtMZdDq91RRr1WDtYZjf7x8hw0ZmnQ0zoJueFW09
QVDuBm8XG1RHSCLCyn1e2RTSdoyz6hXzPWEurERD7uFCZypFJkw51DLB1dyAfXxY
K/IwFAqaKjWgMeBPB8JM5xKTvAZK1alFyCq2CSyjWUBytqjYZcKur+iaRGIhdT6x
rsfrZ3G3Rbr+UFhRve9BKmoWpFtjKWQs/5vCX+XS3wZ5xudzDLP+x1rJBd7nVKp6
agw8ijyMVTrUibYqijcb0Fxyy/+SAvRFko07Yu+7GjwR1AqDfiu9Fc/byYfPIVAk
tsQD+m2xHkXWxfdkySaJu0qwMUObbYMFDz9anQqTczge+bek5FKp59FgNmzgTo7D
tUKGRYIUNS0DjQDlAJ7bwxPjd3olrBIYweMYlUhQcQA5bp+DLEoZR3tB0u6Fsv6d
4dDl6oHwUUmRG2fJS34sxAE6ZS17CO0/oD9bIxT6m4KQ1/CZi+c1+an6AzjbR0Ss
Wnmz1WE8ofrKlYXwaHwn+g7PEv89uSKjvhZ/YtBtZzOsHtXt48JMb6gBrSUOsfu+
JSMAIXSnliwOlnFWR8Urjks/27R0pXvrzXXTaGXIOsmYzryqL9z9OFUDLyrUrSmv
Y0lB6hDO93x+JiFj89u/G7nCp7meUAwU6hCLjAr8iejkCW0xrCPIQlFfx1uq/+D+
95SH71oP+Muya9Gzka30LjDShLiGHosrWzgGwhvMfylf3S9hPTK4E+RmlE89lfX6
bR4EbqP7FIWSA9bHdlpKgr+dw65iIVk6zKLniWM8lGJ74JsedDSm6j9MOrOBkBGw
bCuYSetcd5+hOYnbSw7IjJvsnlbXWnvjaMx/nbiG9fBnSrh8hcIHd8KQ3GtSkgzs
6VkxlzKUSs4KC6TtqC5WBXsgWxPey6enceEuAO8IMXRNh+NmaXoXGHdpCbjaiazp
Ean65TRCXJEKgT6qJmQBw0AgcsSwnAS/yt0V1VPd+1MASpQp6SllBO1GkPI4Z6XY
ehXF0brigL10a1K6Jm08Mn2g3csCZrq0MAK8mfqN/fTzg0Fr9AXedo/++ThguVsb
Mf7+xaLYSq7pG9HAXJGLUlmEDtrI/G4H1MBS/hljQvrNFIvlT6gWeL5CKcV0CtfV
zHqxISnV889lOvqMsTFn218wVHpUGmpK/Zhv6LH9PLaLuN6pHJ4gHw/wQXpPogAf
Mad4ypdpo4lLCJnBgRxNf0LIHhynXXw5++Lz5WM5GRk8LGP//w035QoKzqst0Nyu
BrbRnKTbJnOcikoc1Uiof9A2OI5EWJP/WH24q9ge6qxDfuBt3cxa8HDEGwEuaX+D
mGRDwKM6zSWWvqQ2ELTzMU36d03cfjJFlFMVuj+SQVLuL2gD500cUpaYbe7f9qj5
r8Ho9GU4VhNd1GUN2S+5kV+yIhjwQ8Apx33i5Fr4qrGia4jxhsHpmQWl61QIc2OU
pzL68S5SJ/e98/Pe8QDuwADmeZiu4sYHtiPZew0awOT1YfKYEdtsUF6usFO3N+h2
sQXfpQndvP9ks7UCAoByDvy1COe0302VvNTNQtdgsokxf5Zt3o5r3tkyBf8mDNUY
X2y8Veo2uVi4s+VOWiGoYnhZ2/k/q0Hs9X3FmyydB0uH43abA7GocEuw99gzqyFp
McQ0tmXutdhvHsk3rXpM8o5X6GLuOskBS5T54tAhThgUHOr54yMWEglXmSiAoVeE
+Avtq1jBRTThIFEtQ8BBAq6qZuE5jbtutbFE84nz0j0vTRz8dWPzs1/ydtbjPJ9w
zd6zTASQPIQQp+u+0xUerDZe5Y/4lEQYMyCYFPzsbkXLj59FIyp3o3d4b0drNTXD
tiG8hwQqZwkYHwK0BmNgjIRPjVA0hLzeDo4LDART/fxKHIEQRFB/HC4GdgWjD1Tn
bRRMKloevIgwOQKwFI7YFdr04/5k17CwwfLcD9kxeMjO8t2KqSbMUpmqpH3EH5Em
o0bEWLPO0EoBRQAFeft5gmM7HOtYepb3JYU7pjOVFBFuILGpBe+L6Nf7hncVljpE
QmjcvQZbandxsFEPAWhp44hJRMUrO8D8W9yfWUHYjJuqPGCTKc0EpgnT38mFS6Cr
mAwMAO5xXk9BZm2VoSO9FfkE23NjgHmVRTIBQ1dao6ilZ7yK35chAswEfdeFRSxz
nD+uwSC8W+DQb2zkdBVxh2gWeemXGi5Dno+v7uXxq87HHCrBSfXakS8qkgKtKQfB
gTnWcpDHa4cHV36FwFkv3lShQQuZSQeKNnEGV+mu7rfR5TYwRwser0ZyG308dE8i
v8vD9ROQPlYXsl2wiPYFGN3NQSN+IQVMmWUgrYuPkTKOCi6qYN8XxFAMM9L4mI0u
CsSlbSw1ZMS6bupGmEZ+r1N5B8wQP/MtPCLgRlUIJti1P3NGcoAAknbHOIMovjqE
66xlLlkJYCc4pfm6J5zyvQTv/6DMqvWuljl0Yxy/1tfg768XOGTPWi9vlDNMehnb
Fs/tCDt1qtwmIwSs8k1p5c72nxkGnL+aeOJ5Ix5AveZfUgDUoAEYjlQbkZj9Ws31
KieXnovy2v+hNg5wm3jogzBNldxDNe3rVMMdjLNHeLMixeEBoK1CrMH7YW3GORxR
bLd0rPWIfav2QlF/pakG262iesU/tIjZuOQbqounIn7iRYt7fg1XEDn7H4kKRuxa
7cV6pZoKXqoQBJ28Gxrwsf1ttCWofFqSRony7IhIsikwkGndU0RJrIbwsNXi/uny
plHMvnmSS9QvL9fHbKMXihj3IuXwqYwySuqok58thdzDBorNMWZQY+kXutKs3Q3n
O/SbxODUPbW+MAhC0xR4eDuiOUkdJW9RLBlUSuirkPBMS0VbJABBSbcgxpXW9DNu
TJL6vI9x0Bw9jcwsrPnWH4hV73BCP4zfW/wdbZY/zlrUALqB9QQPzornfLr5TyjZ
8OIn3NR7CVsukXWem+lA4FPyndn55F2n9tU3/xm4RQn6pKJzXmWHa0zDk43higLD
EJYHPg5ohttbHThiPIXZFrKH/Bssq6lJ+CyBdByVZxFuOy95fr3Uh81KNTQmu827
R01yTybsqWG0CemzkTfCAnVlbxCn4O+mdJXzEIyYw6cfVyCAws1Aa2mS/jDoExYO
6quU80yYuK94QGQzx4bkJn93nsIDW+fRlmcdOL5DOGc7cXqrpZbVbH7gGuowuDn4
fwXaYj9NleWnTnSY4oIMmxxeH8FfatVmIPMwZSWFK3xeKgHvLzJmfnsab3ZCihLP
GsXmm3sr5MdRRpl0z78ajIX4ZTAP0ZFapuI6o1Cpzx8DMgSH7l6wmfCXtr5UHebb
zTP5u18ddLOAol3wrob4eHg4HmNmGpxmnkF7Uyy1ukgu6cKwNoEf8lhvYZ7xI0rE
hQ2HDwnDdD2rHZJ0GrzKidd4/uS7fqdC0elSZjTKgbn52XJvCEzxlLi0+0v6B1oH
WszGtSig3eK7pFeCYi6ABdKfWcewwktUtBjw4S6DxiIMBL9qp6Ppci0VxR7liTbd
MHS0fNCH6Ksla5WuwfMndv8arDpkC/x/rvEbaq5zWKsbUJ0m7DNKhOYE2sKUNwPl
qNeqZZE7K9Q1MLJZMF6WFy6qgiCr9Gmh+nxKf5kqwdgR7+/aDo//6QG9J05osg3S
lLoEInv3Y53KrlUGaBhDdjU3dZJoECcJcEQiczYN8hm9qenLjTBUSbTx9Nmwj/tY
sAUDgrQ0dTRaWPc83dTnJj7RXjWz4u7KVIVcCzjFR7dh3gN85y/4e967BbL/wR/2
kJHu3BcSI9TdkYhQ5/rnDWJY2W7gZ2MHJL4hGUuESGpnpU9CLt4gq7T0J9qXam54
TPMPCVoLpOk0JPNp9oXfoLiKFJIXd292KLKKvxL8b9ylrJJAeHtLkHAL8S7Xzbfz
ygWQZUW7jRqAOhVtglnChYe+p2a3pZwbMwIfdOBc5tDTv44IrTcGuqDj2feTvHB6
FXAS0W2i4qCXJF4vGl+NcbWQLsvTMZXLbnvhSl6YXYHu+Hdchz2EZt7uX62hn1Ui
JPDZtmHz3nnKuEv0cJCII51iNjP5BVa4pvCU4BZPlBp4H48x2bJ2EOboy50EUtja
FTvcr66kDgAee7PilDog9V5YoPiX2x7SNqyVCQ0ncT31N9GVCjAl8wU/6XZ/2Q1P
zz6PwYODl3ISqd5UTn19ePGT0jtlfV2d0tel0ug33hvjHP6mIfrpQDgWhSQW9V4d
zx45M7Rhrv1AJIdHBbRqSB2F0wPMW69V05zWusC4yFNeLYHNfeKITB9f85sLp/3X
rRkrRM28mFUSW5f4eIqdBb8V1qxl1sCGTh1IM8NYAyr6TIII49Q0RCb2u4p3Sfmn
zA1eQzvUMRZu6CoaleYeqKFt2mh1uVbebOGgKBawhmoUgbt3DvM/aJ14EeSYQvTR
U/FBHrGVvPTDxl/yKHn7IX8dJGB4D2/8fjV49TyoYpnB5NBixrFzdQLs/WKhLTDM
EEijb4KKRghrQ61fGX9X5ZFaO9MD9mzd+IdJEgSsa9t96R4X1abFsTRnVdA9NVpe
RpU41b1VNEc6EZh22nfq+yeZIyQtO6LsdJAjOq1E8nE1uQp9lf2qIjMNSQyxx1Tj
LCiMGMiHwQhFNC4LlQxWaX8WaMsazvyExz3EtUXAfGv76vwwoF5xgX8LozrHQWXr
YmrKkTpxvpblro8UbTEW6Mnnf2yRD3Zd23zz4BhRWisR5g5yryJ6HHBlsVdvNks/
Syxy+oyhV9pUa2Yxm2g4fdnmkiAlu4+VszBuPems3nVhf7IvRuBiUyg4tplI/NaF
QFknZg0BeWH32pFqN9tnEUWeEVXqGGz1Utb2SdxU0y0RPDjs8bjPVKvqZlHZBd3f
IN5P+beIHbR+Iuy/hpqLDNNAO5n5N6vpmxIwSrUPnBi4jUEvKeCfoH+dTH6Apwj7
yV8v2bg1fKSkFBU9V9kgxH2L8AAhAurq6gSuC1RfTU7qVAi8xXArUlL2o1xn0IE4
WpE+FR9BzvSy63vqxUTaP/LeBv9jbeBfPB9X9ROwHUIDtjvkGC/0KlYEnbrxqxjL
JU8KmCfP+AENLoZaDDvmVtEOGTS1WfIPhfOks3rar4TzpO76vZcIB3yLgwlkcdJ6
UA1TSVvpn8MypzndFI1qOpBGMg9yfwj078vst/iCH0mLmrewt4GogbEeHbtIC/mK
Tk+Wkn6pV375Fv0eCwRuU2jeuvwOELu1/FFp2nI4VSGKUQzFGqZvfEet3RjR3RKB
yr6Xo1KMDQexJcDORI8wdQxVQnwSC9Cev2MA3sNkmZJsSjhB8rFSvYbJmUv+jN/2
mfkWNi0jzgG8wogJSRP+rCjZLo0yKv2WufqfmVQ+aV8bmURxfGrZZN8XkgvBmAsl
ThdwEwkOQBzJ5cAGQuSGSmIPEmpDalvWdJxK+fglc2wOUiXx4EWQf0X7OPwItIHZ
zh8RtFlwcxmyHYRkQRzKpEOlD8zPnRfQkpUlEm8LgPqtHuBUrqrGcpgyBm3z9QhC
anaduIdS++GanFvwd1mm6vguggdcdVPcGrEWta6HP+VAecDTK4O1AvrreCwobw8Z
egI8dF17vrHB0Yh4bLBAF/8e8IU5WzCTFQt8M4wMi05uCdNBkRI2TM7CHlyoiD0D
9Ubqa527uN59M+5jHuuIciTd1TsAdIthp5ibmyHIK1dWQ2af0pQuwofr9Kcg9k+W
FTEKuhGmQ5rD4/pC//qaGVaXgBxKwuPGsPkpXq4LlK0QkLd1LdMXv2Bz5dWfPjxF
WYtpniOTmzfNu5VijRwindYGf3hiIeDEJ+gFfJxdCPas8r6KuIBZLU+oADdGBOCj
dH53TGmtV4RwTdLryVGuKOx1oRake+iAFUrrED7lsbRX4QYmo52ch+zqXWzMsHJh
1roV2uZIJiJ1Pu89RtHER44mGlXcam4y0+flAhh2nvuvK4xoYFWiuZBAD50w00Y5
XtrnsbtFQhfyP4hX8rdU54GwdXbmpfrdFQ9nydjAQJ8cv8yCWjaf1UlhWppXjtrj
xzVZT8VeRii2gJ1VzU4re/TkDJBQK4vRWzHVZxn/mw2AU9PG6ibZHe4GdDBgjhph
L0Q1IKibhBjgcbzxIDezajt7IvjSezV+w6jjW7Vg6hX2J5d9C8PQM7QDxr63BMpO
J+s9v7+04+U7zCR1BOjfssG3WNPqu2YZ8Mxu33e6lZCwiCrih3+cUV5vhosS/T3T
53OMqEQ0SrtFPybQDG2p809XW+Xnq5v6tjvfzgZSQXdCT0Pii0+DlNmTIRZ6FhmF
CGAJFBKvjWDzzeYVyIM1X02PnEE2+CLT8SHV8i5weUhn/SmogtdEHOp0HxnJ+kgy
4oJeLJn/n+YfXDoZjiinnyREFaTiN5zHV/VsJLFSzGPH0YKBU1vqnZcMo/QKaIfS
i62cA8nY4W90qgSY11dbTNWnBlAZL/rBzACyb14L25IuuFD2N6KXU+0t1NNPejVO
erLh2NujIAe8syo/zo1FuE7bqaJgS9A7vJ/K2vHMdqeGNxyDV6F9BDFWnpylFiSB
VJCJ48ZNhArOYpDyiR9pm+MPBDIVDwoLVac0zFeyz0KXAs0fDsMmSYgm8D39u8+O
6G4I0A2T4b8kv/geC8O5LZirgo54rSdkV0JF3TwLt6C0w3nxxWHiFtyRn62P1G0F
LHdtOLJ381O7LdtwoCYYOBqNZNPRA1GzGvsNPZmw0kT9CGDsrgNQBmAYHSX3ozh3
lT69rc+4KmoR+sW9iHtdOynbB8/F81Zp7vQjlUBeNV42DKQ96Y0PE6cwCV+3m/zQ
dSbdtD4FhyybQ6KTxc7yZj+tsjtZ5FD4yZoKvZCsQ3WgmnFcnVcFCGiR9mY8l/AQ
ACXmrujB3brs4DR2FY44O0TSPJkJa836ulcip8kDgocbhLsO3ijaLjXld90CrRW3
c2Gn+KUHbVoLRKiETh7Qs+SmdlsUb5wnvsDgmY95SD+QwypcahIGnM7oqqiFaH8g
CMkx3qjKSroFosFRv4usGd1xzFNzdBFycC6+b2jGuDEBpSITKWM9asb4AnuUwwo1
fzyPkTaXFUU1xoD/0RSzjdYv5y/UmyfNsybvvZVvThhK5eIBXO9cF6yo+mnQYn1/
yrQLwpmfAqVHh9tjRV0jbxW3IoK7DBgi/0nqmoOH9M10j5T3A/IW1SY8rLVdLc8G
bqJEMJIbCy3Y07Za0hGIGFtmsKKdRM+CktJbE3j1SRJqQ5mErffEdZTs6t8JWCNG
bGqYHAwhMpBU3HeZrKwtOV0Rpqer865X3ErSxUY5NGlQCFgEjHgfcd2KYcLKayGi
m2X+uUWxx1zXWIpJJdEWD7yG8Fb7nIth5hfN5Sy28ql0SBZ968KwsnLWI03JCfVg
Wbfmuort7tF8YY8Ev+shkKU6sDLTxwyLbUU+a5DtMbpptDTA0CAp+zcCaz9gctJU
vdLvv++Rr2rhqFAHwuGwl5UGBts+jvo5jiscUxqrdzYqeXjZhbhTqXoGloHVKJQx
nDTlIiugiryVmoMWSskUODWkmaG9QgVE/6zmM3zulqoUPA95Kw4sdPygRzABILAQ
pXMgVKSX5hOmgWvBPfHrTJOSeMnHQoWGmv5MPawSPBWuU5oW/pPmhr9mpS+wLeGh
4/qtSMPgmImaOKFUdTJzEWHhcUmxBZykVTMKiQvfN7UmQgjGuUUmyjbfvoOdSPji
OdbjAGd7fI7vnJMOnDM+Z16qaqzrKO77E3QH06xduzToHKOIkYkoYlAQZSxP262o
jM++GSgoGbA57rQm6bEnDmnkir9+HPd7z2Gfr5pXCmHzOHn7n0Vur62upMw35d7f
HFUu3WRfSTLAIlvsacAttQ5EqHW0mGXenRohmlBxpXLLQu/Lv6HdHYvhABID1ce5
MRd044+4TEAWulKuYljFDD69fG/UyhvmmCgA49FZHAjQ9yEIqbixBY2/LD+XfNo9
mRUpZsTk2oa02JmivJTXEngTN297IRx68KN5NfB9e/LvoJZAfsi1AgSOWaUrhPvF
oG+wFVyuZg+MIJY9Sq4S1eDsQNqUprVtGBLDY9IDap1EdtElfJJnzNeAJKpeHL1k
k8sSid4ZqJp0vPAtGZAL+D6YMfJj2cYRDW2QCHfZcsckKw8IwAAFzVrr0oZ3h2+q
v7bhYIs+FQ8Tb0md4G3Gz0+Y3B1rPqthb6T0veHD2LrTppyDGSbgJ5j/neuFBXM/
m3n8XL1lG4PH7Gd1sMgCYoIhZZDeVDdxLznewKsXONzZRkCxYthW7880uKmrdpfl
Mgb7TLXWbe7WXpUKSsf0nONz7hV2h86bHxysDzCdzy1DEcLVSQ4xtUYERHhyEttp
LBgwfLY9n46qixjpBqnHDrID7cwp2OTQrPGiWfIyd5idi/yvugNI2fsjAsemZ8JU
EjTzdJsEVusdyiApjRCVNt0ls5SEjBz3gcMXRzA7Y0HGPi0AL3p7/P5PtMn5utuZ
KzQXxJXaKXKFRezNxI+mg4B9KfMv4wKE+nqJ91dso63qoVg5N79zfXu6B11hanUA
ElmQMQBfN2/q7PvIfLFsXzZ9eJwRW0+H9fm0wzUWqu8xOXsLJGmJDDl8t5P2Tyyf
w+9GXnqOi6XVUticY4M51kB/I8Q0W39FXZtH0npXtURe5Spx35F70DNh3bqsrnhf
uhCAKY9Y4lHvf71X++usZdgS8ikGmXII3vgcLEgWOjgBqszKrj0jUnSwFzmnS9nO
H6SWiQ11khGv+7yAaqz+9ePWudelEvrpHUKEY9ojtbvz2mI83Gdscp+skKGuyE3T
s4nf/Llkr/7wYmicDPymgdu7n/OWzgwwtVcCRlPS1KO8DaMOFCMiqWrYOrLEjKI/
txIN/rnz/V1rhe5x3TuicLVPi8zamckKvxMfHfwV5Ram/jTz+DJY1HopyPIgojX4
WJpzGQXLH6UQ22/Z7BtTMPva+R6FGPdNqTe4kLv9IG2H3jYw6H/hmXHH30qf/qy1
JInZb6eebPvH72d6FzI3c+dBfkOFDt3Gc4ogQjvQMf2qhVS4oDGdvdsv3rFWax4M
oM4sVifyf/IU5JO1HBD+WSyaw8tVtBgoU0cD/Os+Ezi+BFD80OmSCBWMQWE8DfDh
e5eDMExD6g1ZGXI8OJQazTlXDAqrIprJ6qOOVp6u+q5SeU0kkIMC0070NT34LTd8
D6AGp7FAU/PlETDvJOFW29e0sJ70OGUY87VFN2fnEQONnc18qf8rLINfrjjVsHm3
+VtUG9W3cFIEHk5TvSh/ykrVY8ILrELSMJ/R70ZLCQI9Ltf32tBZqNdqBnVn/VrU
1fo0lUhfy9TXHBoaefGYw3zoCmSRa0nAgB0xmEJZSaF3TZdJ9vJJSXNlq4Ep9+6X
qYpgiBIED1fVMcIOu0kJzRAg10a1Ni7QZrMXq6JMOx+bpNNSMNMYKmj/S1KwDa4S
7JLIczwJovMOAHXUrap7PUKcXb/6x46KLGZYPiDcbMDpR/4wWTi84on8qR2kRQcp
x4nY7yjTy8QTp23y/jGWTI5MmNqqZu4IHuqpX2erOc1B4WxOEq/uIvf3zNwyixrv
Qmc01+MFyvNqh5nG1M4DJN86RhFkQBe3B4dND/ra/zalVGC1Maw3fpeC/ISwK493
VXIEsFKq2KaSr2NqDI3vHa+/Fz225UkfBfE0aw4yODsCIbRfwYyna5O56cQk1r9W
QrnpfQQsmWFl19fQcx08Zxoa+sKscFtXt4LYk2aBhG8nXqPryfvXuZC3Dk34dauN
wWr0ZKBHq5hRcZalVuRq/hJ1vhfKm8vY8D2UYw4Y10ysg6PpSactlf7KHg6w3NcY
4FbazOYQNWWM1uh7npzKnzHzE+U3q06seicem7tb7FgHwNHyNwohKMzZPadT8fzx
VG5pqDpYsQ0oHeW2jEe32qCV45rPl1pQmmXNot1pzApyp2jh8OP3D6rScUVrbDLh
XtKy8iHsy+2nrZQ8yYbuJNDh4ZN1AmRxIsLUDgJQijZR71Zmy9lfpiPz3kGJ3vrP
QC+PcGrYcEr0kLlXzg4HzxIP1fwIQD8vX388+YG5lpxTxC0VlzViZnB7/qxE2YTG
HcG9wYjs7sq6AbCMbHy8OFz8k5h7xpvLfziJNE6hsc8XhJEnPiHBQUd6EG7ZJ2vQ
Ma5Ci61OSTnsC2y+WFOtvslA34HgihNVO6lGGjKOTMHyTcRzZQ1KCK3bpoDyqMsf
O0UDqQoifz2Hre7FR9RBl07ht+ce9Yjx8lKnRiJl0L5gjjXNJaZjWZ36O4+N21En
6ncdPA0TOxsHWuHxtHxqPzv2SmhyXj2Amyog55PlWmC8Iyr3N2UCkjPumkwmwde5
NmaeXT4B5y9qECvzpF4sQr+qo4ptLWkvcWQfMrxVKCn4DEJ7f4MyxFNah6s4u0H8
MvdTAPMl9fz0xVtiFCw1hhnf8ouB0NJSChfD04IBz7nyRUzTXfd5EaJaCGsIjobQ
wCE9Lla7G8/s1TbKVV0tGbY7+oOBekGMgIN/6r/CmkpB8NaLiZDLw3u4u8xRDm5E
Lt4Mz1MzpY7w61wjfoni17qk1P7o/DWwr0QFl3MIsUDhT7uwIcL6JNRjm85VH3yu
oWvT7v90QydR84ma492rgn4IeRRtF5ohssN0NHWaL4WRsVIO9EJpELMY4T74ZAn4
qT2ZLR4kHTLkcWGxh0LNyLgfFAvJnfA7xdyQgncUjGSuHZOy9OwmxmNZV6G4Lpj0
x6mwHi3zW+gvsVyiinhLZHi5nBLEaVWijyc08Gp1Br9xEUI8YFjVOmkr5O8Sk/3U
u9vpTH084bK6Kg8zfsE/UqAJbAUfhR2e03xzWeWGMFKQGMgzkSKFM+qGSsw0k8KG
qo2hShVtKzLkjynz//C+BcfhvQ3flk5Tbc6dpI8WwL8kCqfx13e6V5glVF8/8hUk
KGbRb4KjdzFT88WS4eeDPfRrGAy9vF5Sc7o5xmoPSGfLBxY8QpeiygbQqZDg1VCf
4vC5tyjFrbHaVhZXQTRXDD+e1LRWXde/VtgrrhTcIKQCbN1A6JLYO642EytbdCiJ
UcpaVyXrqjPQAd17ZvH2zPEromx9AIwIQkuFsFlJ5NmT+ctTu5j3S3aZwqfExrcg
icfb8FO1rUfE4qQ4KdZ8xsTCN7cYWBnZKamRYdEfCIiLmHTRbrcjUHFRVIiwDeoF
UqEuo3NThTJSfqd+PyueC0wSKfgS+rsursBNWg31RVxHnxVFmpv90k6gGkae+3Gl
E/+VyFGr5C6UcuVK0hu1srKCQrAGu1n5/GZFMwlBFGa2Q9+ZJKmowf/Mfr8r3GS8
KcCxVT0rCzQq1Bgr3z31DD6FXyRsPf7PHziQsVbiuL+6AI0aUej3iNGdukOHcCqH
y+8pKLY7DsYZQ6RI7DRRS5tgtsPv6U0hOp52sgpnv7q9W/sROnJBKM0PrKpqTx79
VvNs5hHddNO/SvBoVhcYfGd2z0OpQ30tZz0HLa8Z0YiUOUlBPVsWm+v0uPIwnSi1
lSEIb7EyegMiAPDP4S48jzzjDPhX3vrMlfnH7y/wITQwRK1psICzqP6E8n1GmmXk
iPnaY36pp55LfIuTeZsGbXQ4m2d3+SRkdwedsx4BTFPKKdQN2lQNEN5RChmmkd0j
aLEszLj7ZCA4kQVkTV9yXOGWXHXrz1HsrEBd4f+iHxWIWHwq7l58smsy2Csw+sQR
SezvWAVaUIYuUW/poJgvHxYgJCVvr6oNhuBvry5j7DINM7tZOdQ/8OHncx+5R7yI
qzMH0tKpmSr6/7T5obN5A5MbO65OXf99Xp72Ontjs00aXaOnPYa/v/POHQzHN4dz
eY0shrMeYSsj4wYU7QJlLxzLvfUuRco0rpVjcxmEqUSADjkWOTnVvijnXhgczYF5
dlVbPd8BT5vmjOJn6hBc7Fe3W5Uu/nVTLBBr7B5UsmmyTHkpxGB2w+k7J/dGMEV0
Sex9QSyRqL1IqEOEMqoRoWRMZqTXJY4qXhnSbM2uuSwVtbG7pm6TpMwR0nFCWbYA
Th7thmxz9Ez5jNXe27nTRqmkEFQszoh0Qp21nniU4fzzICDznuk+caPiddiTLY0r
Ekxdsbbh2VJdIfNjfx8tHwigZBYh4xP7k5XuTvzfBASUmo4Mz64R8UMmysuWNrpK
4usKpbgzCUH3P7ehiNjbSrAyD+WokBqG9YSiuLo6MmMJrVJL9veW8ftH97RPntff
uc0a862qc1Qrqke/MoHocOHDDy/3j16W0psw9as7YtD/0Hwqx3F/H/HV8odh80IZ
CyQe/hCft/+Ua+ttrKrkgen37AOGLofiFbfITpco150frUciNgwHL9ulqkvbTsPQ
JlpS7vK9IXC9fgchSprz8XocrbnfELmPX8OeaSwr2kManzZjr5G5PQnfgLsaCB/x
a8GeDmPWatxfHXUJwXX8eURXw/Zz/JxASFG7cJWvW4KBobPlEmcPWn7JlmuBrs8S
1e7E0h3EKmaV9PUW3a9mrudGF/N0dLAnPPxHKYXyipkl9REuFYXvZVH43QTfIvzR
5Lr4cwRcH69a55H/zabpkzzEKxq7PWYSBfkL+Hl9jaSsDaj9FymjiqvObW794GBG
OaljSuZE7czxkG6jnLjufGTybrETmIMrdBxBnz0cX5lNrmOm71WBv6TygFai8AUf
6b+sGDj4OBdq6/7eFNbY+75y6a+DPjTG5xsGHuJmK+OngrXFMhaZoLgU+fl9qZG3
uoVisp+djIOXWKbJEVJ4DtCQKiFpjnsI2+oQlC3dCyrSr194KGs45Y/9FhhZaoSq
5h4Saeyc3agfRI41bgUjCzy2ei0Qw8ppCKdw5et3SlVeXY6stDBSkndfUB2feNki
Lw7xZmAVM9+1S6aU02oqSVU6MECokpUs7AeMCKTmMdQdOu8CzOmYrzN7IQEEyAe3
xrMUt8zr6yAirv3HdzTyjfPre85FcFIGrZJ+6NNFNuRHJ9m5j8FmAJBDqTM9W55y
MU9XUncRw5m4bejWloQn9kwnT0tN65FPs/6ZDGmwxNluFk6jx78OiLWSSD31WwTT
VGK02RvqCOjDiytpU5lCv8vIKDdKX2yJF4id0UWHZChx9s4ZGQKbo15zgTxzUnKq
6HZGDH4kkxxevWwPT3uPco+sMZq1uEH6316eQx74XxpWupAqXimeCtatLdEugzeQ
aFu9BryC5uQa/rfdu9tGoLpL1z6BDSJsmoqfEc8pbg5cD1Qx14wBc8A5P4IcF5BF
rJjVE+//s7M7Z0AX5HF67jkIxCwZGHQ9xVff+skvS+2moqbyNNIy30Th8XzNNmHW
aWKH02bsztVpe/38g9OEtLuQhgvjigbjwNBrP25tgYGnF3pmrHvV0hIFPltsYfhI
SApiPSCwk7UsCZPXhz2nY2MXlxncf9At4/D3crFyeg9k421fTzSqldOPXVtXwbBk
brfp4uXD4F0AJmKOOmdqCdy1nTCfrG9XF5z+qwTJlOGcZM9WcPqfzKCTuvQjan9j
3b0u4RELyr1h23l253Em9j4YWyS9sivYTFxIv8npkeEX1spRVD0RGG85Lw99cMMn
aNNMiW1f/Xgy0pt+5BbI80HgBdBAnX+vr1n0seboCSRUcPpvsoazeWRvuopZzrHU
DoeRDk5yswQqhrTOM2OakwDA9M8wrJPwMyg1q/MHQA6UQuBW0+SXsmJhdK0HTeq3
av5QgW5yPkExxBKg4uuoc9redS/jezs9EBjvw7mcuB3WXSb7EoYLOkX59Th8vHRh
0ui4r2hA+oabXu52mFowdst/IJC54WqLK+xSDMplZ1MY+hWx6Gu0kxHQk2D4mQO1
KTEZ5Umlbfc4yVhC2h4WOkSAMCjhWG2cweqWNwifri6L7BSc5JvGP1ruVwfjkig3
9/eisRLnUIES7Kc+O72onMwZEPt4EWKwG6UFbpx6FmY0rS53HKDJgHUXfiYxD/KS
xaHkUTOj43anYN2wZRTs6lrs3NlE/hsZLCUnFfAUvWsmtr6uXGZvOzMjYnZZAhmj
ikgX79xjW1wcJsiZy5/lUrlb2py6JxsfGESpmOojSWcB3tg8FRTvCdCkj6bUeCt6
cMIQiuHDJLFk5GEdtxmXZx2HGJfDp/74mivaZi5wyEmGB5FOsuZUGGdtdBmHzF6q
Pl92CJYbSS9fJmns2e5HRV6tBSrmPS2mUX+/BA92qqWvIb5cbBFduHKEOF2hjEbO
lxZ3+S+p/M8nm4y36rnfytlsrbXzYnw85Z2Idj4fqlPc+t3qVyozDotziRWe8V+d
qB3RohlvEvdByyJmqnZ4jFd/TKUySoq9fg8IfQHMY16p7WQRIBlqi7gXlhYvRU8K
mcpPhgeD44uVAIHBmrTKXHOI3TbZBzFdOmKQQ/4BigJYK4/yibigWlyh1XrrZGHx
x/eNkYaqyFiAMcsyTKkMd5+uVPftZo4i82tFAnVL6aJzGbaUjux1B6vSSnlJUz0K
CU4yNTNpxzkNZydY07Z3rMaq7Rpq0ggPGKDwNw7V6QpUr6fNJ7Bame/16YnI5UVN
9ds0Oa0OIgKDpu05vlFhb0Y9nxOInJpordEjyNfJ6zFfeKA39fGEXgKbZP3B/JPg
Edm+7jIqv/KKLFQ37Ia2Rdl6JKNLrtcEOcmwMnKbwX+u5oIafAdyfraovrbJmzzq
0xqI6gf2j2hV9DHI6VRuCoCrJQpY0gVuSrCNgXL69/gavZF53w8MB3C0dXsh7Fop
7nJZk93QSYCTSQSDkqN63mG1ckKLCFd2MQLGFqa/GX+xMDA6yvcESTO5k2icJFpQ
/FIa7k1orDt61jxPDkPCShscwitVTcprunUYegv0VopHgLTi0P5yPv5S0KzneEj8
O4M9i8Bhutv1IJp3QhkJTB7xjxjoZxaqIUD50Al5RHLWUhmJ3MvJDdn6vKEQlghf
6StomKMMUU0+nnPm0bQed9hWURxZRrLVMNIu2w+v3SHLC+gg6gzTJsQfTRlmqY64
W2wTaJ7ijFyCL7Yui4QzujpV+eVE3Xj8qBsD57AejD9zSC6uP3RuWxLCHLyx9+d/
GmJBtX3J17xXTHEQGcSxD9LZQSe6DUNcq+9Ks4KHB/8FCsDI3Jiiu75NTfNVNu70
Qb1Ce2rq9eywQq9MMBBK1EjATorUoP8usIaM+v4yademkbqOYrFZGD2E0D8peLIG
SdlDDHygrtHXG04wBs8w0mZIQYHdNRGbt/y3oS2uWG3jtxMasXl5jjeNb20aD+nN
KKIWsHw5qtbOr3vKbd5yhSAhkZZ5G3MUCIZOR45OKOBPwttJddA9JvR82A1J+9kw
HndWxYqi94HULP/Xt6WlU4WXeyMjhwVtE99icgRtp9Pc1Xtxch005MKghiZWgHZG
nvuYJ4GHTnAbl5ZsOVO4bT0YArrEEx1/PqrOWdLA9/z8B2xcK6yhvcV/ZkDbWHa6
QdkEFeoVqfvFd2wXI4qdu0yhl9ukqYU1YP6g+RgFsFBJhPyFWOP769jBiGgaLZ50
ARgoTCjbXQM7L5PfiDIBsfayiBV/+RPnCr+aANjnvFy5J6aQQk3wh7sG6hm0MDXg
FD3L76/lJHZxeK6jKdIPajblO1+uTlH/XGpi6/Z90kdmjYV1V9EcyskYdmBfk3/s
u5Ie9x4krPgcLAi4VVXfxZwUpKPGR4k3Uo7VgAyLAShMap0dPQiZ4edYJDSv20su
pOpzxK1w4CUVV35dx8sgdPJSLXeHWpYY/0jun6JZIZKlgudMHBZuLAF8fSpvryyf
qvUVMgF0zjGevcAn3u+njkh+qCO/CGSXenJh6Tg1/aI1r1NtcSSH3skurhhl53S2
ah4Gbfv034qBogny1bTF+j0R5m+eP00gXtI4CdVYVXwAaow7wpv1HXFK6264sh7P
lbAo0MaLPjsji73zgCGUVVNpRZLJX0BP3rcK9Uis6G6yZjbSVPA9mspYNBZae9Xv
cxo3sMkYViF3e8hFzD7vwNErEq4TjRgG+SFeVzjk5n89nXxM98FN1aF6Se1mFvNV
yKwxE/T+dlJ9WSjb3jptugp8LWZ6y8Bl7zcXXUi1I/TNzYFU635DjxtafhlpJsl4
b3ckHFKzjc87ta5S8SlTPpZC9QCIyPpJP6wWZZxU08lgNoLklpUcJ/VzNlxdFkL4
g5nZ0PVcRp+LUQBV0P6bryXoIpcEyoVIRQmHEetHn5vRQBH5ShldIZTr/JGQnaJg
/cpxWFSX9O+rpudnLqp40Txd7Jc6kWXdiwAFYz/PtxQVAPJn7W+j5xv6eX9pZfPa
ETjqUppO3YDuLzf2wS099qI9jBA5hNG2CAUD6cRnzB2mV+Fbo2FZH4tkek5CUEKk
WBVASUvLXwzSZXqtlAYdvHrrjDEk5aDJ0E78b2/ZLUEVPS7QZUzmz4WX1tqK5Fxa
74/SKnHYOQ7DpoV7ZfPvuqwS3ECF6iwMPgnYyRIw39Z8TfXA5j2+F36X5lPBu7CQ
MTjBV+vDiSh6H1v0XbB7YYdPGjT4Cj9MO4d9uMaUGpMWkG3KvJFAsDNZ32Ps70/s
hRriISt0o70suuKHE1oCfrojT6hkFqwzxGabEIwAr5cMkYTGehEhA632CbROyCYo
+00U6czp90XhecvMLvdgahOOxlGUdEbW1Ltcmjq5zKU27tVoZZaDY5h8ExdTyqtL
DS5ByEP1NSHAE6jZqa4CmYb1KK9LTrVvkESVciW9Xk7nCD86H5Bd6ICJIGgrYpfi
AiXWHeGxb62IvTVKoVUT2KjeXTeXSbtwpdpG2VdqSFIZcfGrwz0GCxeHSLclGVtb
u6xE29XghOxFeRdJaEtw5cvE4VH4NSPbm5n1rBi6+0p6M8sxSjgjVJlsSD1GGudW
l+dli8hBYHzbqjaElGGnOJ+unJZToxtMKZtfA8DxJ1pPXRn7ht95oAz83JqOT2Vf
ugDa8b497lDCmy+YVll3tpjiN1YUD9SAKzwmDYtAM8ZF4M0HxF886T4X6xFnLMF0
2zg92sXo0h3j+CqvJLjoucAHnlkWiRB5+6wM4lkQIndf1KcOpXMoIyuwn00SnxSG
AP/vs+/EGqILAMCbIoMaCCOOj6bBnp9NZm1ZsZvCIZs5eWG7GR1NCRAxTzCO+NWq
DDjw61LiwSlOP/Y6mAvNFbshdYs88+6pqPyAAp0LYJ3rNATwSOaQTZd86VctWg/B
zYoCfMfHffkKgUZ3pSaE+Z2GzVPe3CgTzUuhvWE5W6RmB/cKMGF3SNjoPGANiW5G
W2Qj26fMzYHd7cUfGAIgc7gjSlNQ/ytnZaQlGvkTo9F9dBltWBjUnSgpMFHnH5sk
/+3jf3NXaAz22N4vtf6LhE6ODG3vN6F2/nnYdlrx7mD7+S5Wmv4ifJjgR0xvNOqZ
gQ+BrEsA20W76p/5Zqp8OShdsVJ8WHvg+ZkaTo8cRup2sPDCV7K7xPetMphdwho+
ls0IRim1SnqICB+7sqilT0pqNpvHjoNgDjP5rUkoITXs5+lUVG4ZDN8xadnPBer8
gG2PCo3MjHCcKPNdoUwOIBs0s5PkHr7rYYWduI3Li3hvYNsJkZAMaBooJIx4bS2r
friUlnnHow+aIsWsTEgPk93zf76KVZ6zjx4cprVCV+QnhFc01Bp6moXZuhiihXy9
Edin0kq9MhsI+Nbk97/0QePK+/XdrbIrdjVS05ItQfGhkhxtOXHiSrtGn+FQLZ+3
VA+TzBnqlOJzagWrivx9zJOMDRMhP87Qv8wauroilHMkBT6vf5+TC+nrN+NE+Rj3
JU3fZ2YU9Z35U+/2DQfJ7e5+NciSTYvALFtwfROpWBqYvGykX3ZKDcbMB1tdzRPx
1YFgGFI4NJ9cg/jQakdnm7tlfsOEffRfwbgkA9o+XBnpDy8dZ4+DvUzOA2pF/g8w
ol9PZGbA83UStwvskY/ce25G+2Rw+Da9F0Bm5zXzNbunhzRePI9nmOM+bLFBB9/2
6XxUe4HO8NRYflpP62Dnh5BXWPr4s9oGKom8bG/150Tpy4BGGAjjYVrfLSKb42/X
hQU/Ss/vzQaePOViqBK847XrHinBH3GMvtEAsdwL5U5S9oKbguZoG61ZCcJkdbvI
xf6Vjoh6PRvdRaUeApkYWbV0/wKmqHK1wzScY01gHcubMIhdScH5hktKftb6mDI5
i0+U/nvyOjWUIiPOoc+InFEHiWKiydqB/JLSYL/osAj7xWnpiuKvl7+UqQxK1NME
Fmvb+gIoZDsLS+qrQQ3qOgxajy7LNgwAub0XFEbxmDo37AHBgmYJfXPQrIlxiDuZ
439qreD6LsioAZNKeaRvrkzsDQ2urnDiZGEGK4qslz7mKeKK4dqzQgTaDRKmmuuj
7IXgNv70/d3uHdl7lPbFgJNDSSdOm0NK+m03KKTuzTOxdqucB3t0gkqRblZFM//H
0aEN/4EBTkPvmFSFkglWeKF6Mzphmo996WRZjkKCGXvTh7NiDwpn/43HzA8vumir
a93aDHqgJhq8L9bOeuAVP3dHMx0Gn2awfx8OlgHNxwnwzWtvdixeTfXkNzMT7PA8
+3ogq/aTA5hZE5XVvUZB15vhAl7YpYhh3vlLnnqnrcyKiRL4e9eyxgDf+gFBhvkG
p2O+VzkYZLucB7tr6zXx3PYyNUVd+6t6L8OfBoCMeqgRFNNnb7NZ6qmJn65SUwU7
pw3LqE8q8NT++gvyPFjl7CZpABmvqLucG645zAaDYDRlfGnyxEdoJZpdybd0VSc8
FBmpo6zvtsbfa+kPRz8GT1Cs7qsJHmNC19WEAwgUXD45ps1u0P8iS8z40ElgWmH7
F1L0ETQT1AzcdnH1IZcxDbXI09eDUryDATPEZNv0KC9hjrjb/MZaVm7YMar/SShi
FOFEoaUZ/xCJC/m7RJlMrJleXLAuZRifstdQ8osFkpnpkfcCipPHf6+j+R9KjYhm
oJgo9NQ4tkSBzA3Dr5zqfRXrs+NLwr8iTkXXl/w2aB85zS2I8UtfDSdRN9nYlBba
7urqkjb43sJS2zQXayE50SY28FjsBAtcGYIqbWMOLdQBAsmIHsvI8p1BV8GchhVO
EPFxTvKrJdx7/vxbY4+umUcWYK5Qe9BtheM7EdPy4jX4hnmxXzUv7wKynXdcWWI6
hpf9C+XRMH3T+K/JVFoqzxTwePfuj1Kz44rEv2HU2C/PcJLDuzFPSZxwJGLT7r5Y
/FN81erGLnb/Rc0KWGUFC3sF/TFm/KZXh4dF8evNYE6ydNLl0Rxs+thfrYu4NZ7d
nW6a4LhBO66bqOWp/XiAwIWCAqTo42ksyz13u9SPattPzZ05ogk9JW7vxgId2FcC
M+efSqnIzkYchtVL7mz2J+O1MMJMjkz5vRwIK6/mqdiqFdjx2lyMUJZ28U4oDtBD
X4rfeZgmyuFCKYRQRsJuwHwx4kn4O/puTXQdmYV7IDOLdjaMNj4HCrQTDYVMT9kf
CBlepRULJNG7dsQySmCiUBeBtkBg9WrMDXKBEdef0frmZlvg9VCwM/5m1hv4wkCe
CLqgnCGkpuN71OFa4kQeWvQy5LTYZItHEwgJc2dI7DGijnKFy8lhvkdKY1Lwxnge
BK94TANfBwXMSs2360CLup8pXX/BOhhETrWHB9XWogMlVYkGtAdko/LHxoiQSxPu
GoJBIGUQdvPbQJKrnBoqUl5nUmu5S8H94jQMni9smaSu0aQQr4ioVOk9ZBYOhJo7
d7r7230Dep70w9MfJwMNeSqfjHb0njS/SVFMJch6EbK9IOut+f2wtAtuUY3EBS6y
tvnUh9p9nzHiXug+aRPKvdrDvmdbWJQtg+j/1NhojMZaT4Wp6n+9DgA9xj6AAT2q
k0naXtfgSC8fJdBe78UFVgZJXDACpFeH5HT7EwiUDOpXS98yEaD92qYJvNoyeU+N
In0h74rWYFdtgiMR9i1gbozbgxmcP8nZIJAdnBPfxAbY30xAOo1/GGnhdHpkU21M
8x7FkhUncfU0GrHzG+eN8/+CWGEo3uEJ/nKQIvwTJcG8A9bbuRXFuHTVHdSHMQvh
gC9gbr0izcLY8pXmH9dgW+1x0XOEfj5Vvs1tY8jfMoYFeCKjcpWhzw9Rhw8l2Nh3
AWhP4S6lnNTTYzVpuLg+1SFSl/qnSA+AzDlJPDIjyBmCt4Fi28hMkq21CrE2ojsm
NLpoY9jxSRjZDQGKegUTyLPqhOG0CLLmhnqplZNhRdMS2UPbvquK/3hJGZn6d8mD
gWm8MmKTR4H7HVeEUAohIQoqIol3nRUiRnmywYtAcpv9cR1rYjPq3RRkKQGvpz1w
6LnCPqTWTgV1VD4YaHi1stUW0h5DCktyOw0i4bNxWQo7W8Sm3APdsIb+cuoQiqPd
DEGNi/+0FU6t3RFbpZ9SSNbPJiUqtY90iPBr91K0N9r6wyN12yzXsulzbk/ihgDM
U1t++Kw2jonCVVOdf22dIYVeZVZ9RHxN83foOCTt2Cq6EciEpobd3l6BfKouxFdb
vOqs+AFbJxCrnE6hl2/RYDB22xoMrJypY7eo5t/C5GzJRX1fpoZ0UbHcMUZ1FZIq
w6/JhS8LvIL2D77BQf2oErnyTB9a4+v5gFYAeYaAlYj42qx8NQ9vfxkfCZ6QiLD3
+mg/wLSFkpJGbA9DfGyfgxD6XxIyfsmSpFy93ZI4Nfj2NWoaZhfWBqbeMLk6mRss
mRWwvjbIgxaPwJkaZ0IhCtLsGuoEXgAhZ9qCHNl/aQngzD6kL0HTAJGo+lEXya2P
EGpdJdtlcXXcONzzxNogMEXiFM4W24YAbGXWv1VdcM5Au4abm+2J7DnrXoSTqC7P
xmZa+7mRCmoIkb4G/AUPXLyq+WLttTZ2qTi7pCic1bM0L4hvvbSD5ZY8nes0Taiu
ag000WApVOCSVTecTNg3ONKTd03LsCXxABH6+K0U98rmFAyXmJu8wwC4ru0PaJAe
XMUimKwZlym71jsX4liP6YJFCsN8Cwm4tmMOk1d+q31nZWmpuatJ7D6NS5dfVyS2
/y9wsqOYbvY/lH20uasCxYgPd1A7xBs5cnrGuZlmvubBpg7XHpCMSS+Vqr15LEEX
bwnRQaKr9xEZGs7nX5Wd7hOlax58oRxNad0oCRc81aNOQ2zED2+6vKYCkG/FqERq
6vH0w449dKTEyw14cyov1XYl7U4f9R6pAMJ+hWzTu8mvzvt5Ge7QW/MYgZPKm5me
E63AyXBrzkYNVeDcqlixdzJGypPA3msami99hpAJQhlI648t9PzLh2MoPQ6Pcqne
1ZvNPMD/p6ZHHuOeGa3EPHzBTXgHhlSLL+qHmqgtjlBkUFYejiqYgpZKNLHTB3qs
t9bT4ocEp/fGg0ll6feSW/oOHjPwpG1rahe/W5UkqM3/AdXyr7Se48AzadCjpF53
8CzqOYaTpnCXPFSQuBEwiUsjr+RQDQb9wQVkbvwWuOog+caHZc8kZpNTLm1UlnTy
59bU0ESXmriGNu/pgNKW89JdSCn7xfQk/VHQWV4SZvOiv6nLUDtiwX5PVTamFawu
g95VQwZkvX0rOB1DpVVz3Mup69JpBmtB1EnSAI4iRGwxm/PwYD33d3U5HEkzeQWT
ixIgwirqRaBZ+9e2BBnPgIiMMbJVvmzMWjHxMqcCI86i53M1iehsgTb5mHfWpS6N
Sn4PpJQb67GT/jZfXiCeXmW2+04AsHmgDuxynZe4ilRsCO8z083BYEsobv/W9asz
fiS+QhmcO2uCw/rZqE8/PI9z218yZO0VZekLP6gF9Nb3wuVvu51bdo89pGWLTVK+
hTo5vVXAskN4aom3rB+gnvhtaIRRZA5cp73l5XKAN7L6JTcjd4N9g4cqmabKwev+
6XmDvVJyNwe0Vg+W5I7RGfZRypY1ryRQdDuUX22Nn8udbcrHMzAEv7PvBCysAJdp
sbmVZfR41VbeJTshgNYM6yQbyHoRd9tOMOFfzufGbWXsLQOvAYEk5yy/OxtSSVXp
tek6cRRL1jHVh43QUaiVpuNiqBlWTu85P/UnN4txRg4EwEUPIuPgUjjzFIQtNjOa
c2ttvLOG9eYytRxupPrpwfesX8GpY04OCwXR0+fNpUogf1B819rkCyjNth4HyPnh
CPqjwlz31nd13ozFqIGGUcYWjd0JSJTzL9JJdQpKtj81iHs0d7JvgNrUWbailSGP
wu6SVwBqT9iiE73qaHlLdNkH8F3mzJKYzqKOdrXwhn4GV3ajKkbOU/AYMHHJIOXG
c7PpcFl+8IpPgiPg3ew0bRI5ttYUVr4/E3uXW8I3PaMO7LKxeyZM1bp+K/b+y8sA
0dL1GHgupSWBIKLjqnZc1VSI50ie7GEYou6cHUtAYLvwAEUSC2D8Cq8x7nHD7Z+T
AVHprdFliOFz56rZnR1vVoz6fSXPypJA2bxn2xNhCbhmiJGOPVVsiJwnVHX4H4LN
SW3O60hU4zJTBUEI/ieoNFpiARiq39udHx1odIl6KFX8wg3jubj1TJYvbou8Zwr9
oI2VWFR7KzmXeJ/7an0L2zGYLLmpxuw4SYneBUSTTUlJEAStq9iR6akm+1IUB69/
4rEHva9U84YF7/JphWiMN+jjrRkX7+u3PAMzqWjJhBfkhBZ7xhPxqX6QWfmn/5iT
tgUp8z9AomD0f6rkBCxAqWHXaDdzdxUmlEJkipSXHwscR2qKmlH07kc4fZ/uf8jt
FVKf65h5tF4jnMY0owLcx7PMptJdt//+Tdd4oaT19etpOHt8nMHps+SdI03TfR6a
/H8kcLtcO7g8VeJFXs8ml+Sjzev9o/gf8I3jLMwuKS9048SlPoFq0Bm0AFIgzRVX
xPdZ3FnZYTxv/4K1b5//iaeHReNP16Qh4Uz8uzvhgNAcZD4Yg7vUxRWNaPCu4uHH
24ORdgQFlHiLFCfJImJNwU3tAzqhvxCmTr4bElRgSKP3yVGfuwnXt9t8+bxMInmA
cmiqnWgU5Crkyie6rptBWh4g/gnl82Zh/IBq37CF2xABr6yr8k7Y5dHg5a33O7Rq
pCyQXKcK92GAFe2eofo/qKW23vnXNeLKwZf7Gvy9CIx5qW6aZcJ6IzFI/WhbDMi7
UO9ypTWxDDX93ixJRa0n9avyoiyCx1YYtxEb3Tg8INHGwpm4iARJAR3Pnv/P2Hgx
UaxT9kD/tXAuQAUimwdfqoxUNFqHCQ4szq00uYl+F3Tux1nH3x2VIv4OE3aDPH7N
UKtAKDUIIPbJTk5//TJVoL14bdxqo0OVm/aCFJdgfbgwiztbwnz7HRmDai8wnntk
0jwDbjRuhek5NKBc/SOuKI1RIj1T7g2SgBIbAIgwe+UZ8yf9jpbx/vwuhyf/X+UK
6yh0iwVPZnukpFwWjbJtkjd1Gk+xp5M+kb9q7BOe0h1tnKSpbhyrME04AESIcthO
BHw4oPAPrtJxkqHGFkMoWVII1euKdlP+Qj2Ce/p5YD15OBY6W65geQO57FPwglRZ
0QCIaBXvAqZasMqvE+jLbpAbHXx32x5rzHOWw/qjuDrtt/HWqXlFF9BChMdeH3pT
lGWZ2aN5xXKqDmgX/29Rg4KwMEwOcHgaA5GSkAXcHIyviR8SaJh3PpJ/7EUgzT4b
WZG76xAdHuX+Rt26Taf3qhjXCEKAw9+PR57PtWKdcYFw2JygXmTZLnaEvjF0bjQL
IUkpMCh6Gz89ILeeKQT+ftyK/RgWFx7zMLCYQrBLc+kvGsAXIpjGwcmmgIRZSK42
WSfBleIvlGJGoZn9UVKabr6/GGvKFSh7Lh6mLtYHhifde+Ymxq9kFCT9El0jtqz8
zvDmyOiV4sNMlOdSieYGYjmsCs9d79maPiyRIHTIILOpS1B+7ut/ENCIbodOBGPN
e1Q47NgM2newmnm1SUGgIISHRfI9qWPausNqyjvIHSaUyTLJap2xQlFbugyj5QM2
p9oVLmaNfeTKGd2LMngVcxa+rgRPwDZMLDiQj1XRVaDWy3scFLVqhjOZ3zIxa3pA
NDODj4gYe4VIHiXwQ/rQmOPkAKFMQA51X4GjpAP0hWDhDkDOF5BQS1zRxn6Ph7cX
VNaF4WnB6kntujTLONs12a7+qcn2JVhKxCVagbU/lc2KDO+d6SpHWpTx1kgtp1bl
rsujkBHj6PQlHGfoaEs2+09LJCK5gdPFGZIdN+B4aArQlULFAtHSyyKwOw3rcTpk
5hJTlOto5fAempVQ0KLYZ86pQKmR7Fl56MYyhLPCHjVEOBYjakc5abaOBqHl9Ey6
qD8tnVndYWTFV1Kf6TxSpJGNXYBbdyIuCDVj0TbEL7y2nEEZIGqJRMTa5HZDzMGC
ucKissaV9H/Y7UETWW2Kul/ZxVLwVlC9ErNfWT3dhhxlIyDvhVn/tMLX0hIJv5+0
jyAyF4BBvcBr7pKsN65bckYCjy3cYLBvbMcNmpschNTyWC1J6KYMRWHbYk1vt1ZB
mr18JFjJgHoNNJ5EadrCOh+Ph6aqhmmRRAJqdDxDWQZTebw6/4e80GdU7AN3UJNX
PVShJnsYb8/nvWYZIiURcvLN1+NRusfYde4t0A7DtZ5MzEdc6e5NoXt8r0H0KWHk
j69uWCnMXojYZWb2w6+EMyradZtmk0l8/N+FaClnnGexi0twuZw+zLDDg1cujKPf
lpRhG4TwH/XAb1FwOnR9slpdtGLlDSwJD+FAlKDpgZEzud6NWTHEmzNyr+sx3obs
PhdX2ZVGkFlyq4yWqHSqp4FkplZQKb276DrylTF0i8v71xAcugD1c5vEchGaIjVZ
6+kupV3kMMaXPjFKfZikHQJFSAxvAyZJlIi47ZuE0ilIFRTDn4cULKwDwHtsTxwj
Z1Ul3OkSh7byd4Vi4EQBeCI5mxZVzfpn8cdAx6wCFDn4KWxWLQhDd1wnN6VraPPT
FdKByMwtZZ0F9vjDae1wBOlJUlxTz81lhq022gKe+B0Yi/d/MTaLAFNcqHekg+iw
h4H6E7To8DezK097VSQkO8M4LxxKnGksewc2h5X/BHigLYtUi/30ldK1wK70p0nK
zNL1IAfaYVGzh4PMYV0JLHQFMTGfEYKXvrIfhUVWPyhb5uiqOkU7KWpLojGIcEd2
jPMTz1HcxwXASMhX+Mjey61USt2+54T8YeDDzEbQhFtAGLO0AEvHLXs1qFwMLD3m
4rP5OkeUBxPf81TdOhiiDyB4rpai8exOdmrDlErIYZSawJkflWQr4pPT/fGQoZ3G
QuJKiUiqTWGCKS4oIMRoVFTSpfwQjWxgfblc1tIN6lqFxJcdVangFj5WdQ+IhiST
lF8+UELXQ9iXNJ9M0gnwH5w2SJSFBANWQpk1xbcnybVDBm3LeKQJWIcNmBUG1A6j
V46wSRVHBFHKDQl2oqIGolLSfFE591JE0yduvtN/OhJ8eNfWg2DkbhlvoCClJ8r2
s0IKSoxC9PDvcSsDJ9aaWOBM8ST8ZnsBQsckv5jKsnHYTpl0a9nJbMuErvTkE5d9
bBaCA76ighOdgRxkF1xKpN2ZtYAyPBeX2V7FkLDK66E7C2H/L7Vy+El+NWDa2g+p
8hgU8aHXnjcmp5pw97PED/nb2Xq5VYajZtqwa871oOHArLiZ+MPCgWKsORwweZnj
LXUQ4C1dtuq4mgIJYX9V5kC0Hf8frssCGI9E5O/Mzz5Us6EDqNW5lKfrXUDDiy8E
/jT+M4p5aonA2AtaH3ZN9u7thohrFvx+4gPt04JR8C/O5Zt4HlW6AonfUgWYcB7r
/olHYVeQrsmbAqhwJn3sNAru8osK/GqDQqc7hJh8lbkU9pto0C/VGUUwXPDwtf2H
IJlx4f5kFPfBbm+3bbcxY34RIcV9hxoB3cjHF0fzDePJH/5ApP2h8DWFMgAV0asx
AYgv1iAHGt8sc/CXlUev03LjS2SYDHUJExqsos3pNspcoMumlESwrHVzwOvj42up
/AaLvv/cXTvYyTOIHqUJHqbei37KJ0QazJbaZYrBybwS5sLiSRnmWFk/GdY8i3Eb
O7LCBN43IGgfBZSb5+oXJnhx52kRC8kj6Q/RHus51O0xUexarswblukt0nwB81Q6
t6Sg2KPqa3QviXITc96KHwO0AZt8DX8NteLU1czPi06OVg5We3IOMd+hP5oYJyVS
XAZaseqJWiZp9KQWgWQw4Q78dnxmctF8yFvD7czada2TAN2F0E9FX7WUs9CdqBqh
2StBjBNbpdsmIbDHpUMVunwcsps0dPY0yve4wFrALv+fTQaGHbrzSxcYIh0/lUv7
zCFo8bJ3ON7XUQlWpYuDuC2YkjDAHZq0jIPC4iPb7wudbx72jyqXALCqH6ut0cuv
I9t3fu3grm6Q2ldeajRGfI12ktYzKey0ANZcdw3e8NNTV5eWn0Ya3JlhS8UyAlIg
mfl47+lRVVW96iEfYA9wthDvtN1lVVeMFHIzBuvTIjyRtZuyO4U4xogcp2DD5wv9
KI+PcqX5QSabcmeB/6sFRE62/qUQVvpgTVTxu/u36S8XGCGdKGejKmSxIm5rpydC
NXlCRg4bkgCpYmdsBSFK0rGLi2XEwXAfPZGlVQz6sRjsE52Iy0+cz6wb7JI8bpXW
LpDwJJVNcrKSpLQAsOoQfT9WF/EafyXBVeplNEYoVyRKU//YOOOljb9nF5UXxzLg
P/XGxSiAWTHqIVZ4ftLACgWPHNMj+oFJpmSPvV8u2xKoWVPJZJaTAtP9kqt98ayK
FHiZR4H1C4V4/57bz5lDKboLCkrgHCW9vYYFqt3StlWsB00vMKp4Nez2njpE7DHn
mq+sLxhAkr6PA9HIIqjnem7z8EsHxdhb2W7LC1SM2uHZWHhOzK5JcliaKtVuPqjY
T1eioeAusCSw3UNC0pEC+rUbBSD6wxRwaD5Cs2Zj+Jd/U3UGQ1Gss+BbIjHQwWBJ
ozqw6DRzEhCitSuGtPPqI1qVtBlGq4aLpPKk+0LhTfWIXJLgLIcZ/6lRvzIxp73P
79KwDiPZfC2vhhw/DLlBOIf2CshmY9gUfBJLnrdftlXU16QKf67E1BV4fDRsuFdE
U6e5isWT3LE53OSgARAroKFB+kyaB9RDMBegtjdRo0jIRc1dmWsnMr49WZ7bIDDc
O2j65+BymvDvc0fXmlFAab/x3KA0nLxxNbZ8x+jNL1XPfNqvzysgV27xGJHgDByy
kkbAeoC5Kgq3RvFlR3jPgKChko5CIZ+erstP+D/Q4t76Mmr4xOwadspGzxj/Bx5c
JzNEbzdJahS0jZDJSqF0az1Sx7qvsNTglHVkwOo/DLcD0HnK99fvaGSh79N+3rh9
P9iVZJx8/fJxws8VHy+0ya3/cJpR2PyuwIuyGVmsBc5gKZyoyAuzsKIKP3PF2yWe
vDvyzx5vmsLEAH4+0EY3ZPwd0D2Rxs1iEx9TqEv+/fYMXj+4Cc1V97iVnA7fuw5F
6nTcc23Z2lW6Qt5wgGW4ialB96PIAGbOnPmVFHrDnrxglnN72LRlbt6dny8CWxyw
KNJ6PtE1I+nK86Q0uQp6gBpnapqlKJULo2oZSSqy6QkhOQZYhmZ7muIJV3eDP5Wt
6K3y1g/506P0ZhviK4YEuX28fvC3lD3VqFTzN9lggEFyEoq5kxzdVNBWR6ms5pnR
GMKSVycudj46zXBQ5HcfeWWbtS3G2wO9Pc6i2EialQ831Xj2+8QrDBjPssIamE98
95YWCZ2YoGs2a823p14NdOODV+OgVpvJLHVRhTlFwBgKHEVPdWE5sYZ1nsbntTTe
lvBF2gQwDZ8xjEfaAohNiI/wg9aDLaCnF9nEKXMcHdwEYvd64cvvy9hgH+h71eBb
zU2Exx1l/8qCTpp+ZAHBI3LszXzuY7qsTxxgGFq4eLOQdmlwxG2QEdQvUT04CJfu
fo6uKQmX4VxWOR4i+tdjKDSNENxMwY4P3jubdqaiB1Uo6JufUXyTxHJpk3T6RyD4
7wRBoC/Sf5MWbQJ+0B8d9kaX2axsgT6Zur97ADDbo6XItvSUE3G0dhBXdUKmN8Oh
IjMewnsV1ncb2Xup7FfZqc7xsZVTywQhaW6sBL4Ec2d3wW5WHSOdx97x3NHyNeWu
jDRm9e/6Wj2hMXRtXy/wc2L2zYSLQnWC/FImhKB3+kFV5/SdzrqpEg3e/9raDpRi
RZ3BMdbk23VylFLpM2l5+qebHYCfTzdmoHRkKtL9R+s3lnyCWixqhCtavFMqH6ct
jYSVECC8cawuINc0ZuRPjtztuWKwBXZxdYaL8AEWPy/YlOcB0HLjx9eFMJIrtrZq
WBslKLdvP4tfeLnN1cweQj+16ABrjJmWGLPtTsTU5pKiXy8GJj0Ubc5zAQHJ55vX
O3gBADgbAtX/tPzuY/plpMRCvTmg4fh+LEI1pSw5M1fqJzcrxN9P/rVBNBokG+AV
iXM39sMx1eayHQs/DecWKF53AnMdqn400u4n/5OMeK2f/cpAFpqwxnJxsGAXVSfX
bcun4RLLt77QB4dgKtXakf4eiXbuCTmVTgLn1RzWw+jPyYiNtJ3SYOYzNPdiYILs
/dC3G3dEo+YFE7BfDhehYnSBRAuLgUxq4KwA1Lv7VFzffISN388mMczzsH0uSTPD
WLFK79jRfl7ddjRIkftD9r2bYHRWI7FjLkj3LK/xC9CqNTV7MgIwwiLl8GkFR6RV
0e0A1K/0s+C5Gdh4rhyTwMj7QCaOHLqZjy0LrRxGt1XEWsDLjGabxMQZkqyoSjO3
nGQXaPNK3+F5Ezf1NQk5vXn6d+v9gOpcd5/Uu2HZ8ndRnlEUnOn81Ox4UJ9IvlEg
JNHQOgKSHVuw5PT6YJvK4VILB2cC3oMejPxrE9Q9pzsK4oVy/ZtY2jr1Zqy0QOn+
hg7b27rzS3eAZoshNF1/lJe3z9rETJF1aAmV5APChGfFJJhv1WOgl2uDdjnMEjzU
5oJ+2KjNPMOC4+rm2SXfZgGgran9SBFu8Hlr9Hrl/GCCmApL9o7SR0J/nfXNUM9k
79L28zp711d4gCn9H602A8PBOx/yhsqVTrh4uLzgY/vHINFCpEyChRPd8T9kjANs
CQ0KTk5YBjEUqN+p2fBZHQNZevPXLWBd9oqmYXNQnuRKigguFVG2I8YhCqxcsUYj
BCZXaIMTpD6Z5Ecl1hyZwC8VuyuUsWE/OEH9RmxhPeVKYa6dXVVCvcHn9HFFoF0D
e1Hr28bc9aihhSW9Fk4+qxz6zcjtDTTUrQaDUjEWLP99Eq+3y93dtoduNwvDn2mH
aObmRW0wnF2+V8UZ8IEctcXVpZpJmM74Ib71obt7LeEaO1XXCGVsF/4rqZq0miZI
fluVT4CvsbbML4pd+2J81wLDnBXvXdFm8L9ZoSqQ+7vNfgITKy/suCgTWKtgJGAQ
i+TNyozohc5uu64NO1hWapkkVEraA1WBLqsx+8twEM1zgBpuM5VU7ggl6oDle+9q
J+gjJ2oNbsqKBXi6WX5HNGsX4iM3bcgXBa6TZIVSwhcTC3BWleQjdnqESeuMzY5i
pld2rf8+wUfHvM9u8sKMWu6jB7p5oaTTBDR4XrfmhoHfskOCQppEA/Snkev1LCcq
Ir+rrE03jE2B443zQLGJBttaZcK/BV22M+CACaAU1V1YfKZIfpbh4K083wX2zcSc
4PU2FgMLZRiHuACoUviSH7jXVZEYqRiE2UZyU7LfXlEGYrJRNmrgH+dAhGPNqDH0
iK2Cyhvrxx7vmxwYn1I7G86KAZ7Qa/B/4K3IEAxQ4me/NUQTwy0J/e5Ua7mn7pu7
5OlstLXvkqIioGgg+b5+caGc61dCHFkqgK4jJiDleVc0PQTOzvi6bctR751jP+z3
/Wu0MyRgxizLtDCGTw5MHVjJ2FHTpo6sxJjeXIfSDsFFbq9Le4DKp2BTsA8vNgBz
p5bjzrbv78idaBPyuDYPIvzOmHnalPJ5PdonlHJsxUu8js3Y3BPziXYZJPe87jHY
V/mRYB0/p2Fy1p7mEtAW5guwgHjH/5/bUKwrW5+vdwpjBAyOR1pMZsXtmA5MkMU3
ASyuwzgrdYdNWl4TFbqGfSSfQCj4Ztlu/BTIPtLR2HKCLb7JHyBVNIlPVu6RAlwi
hBG1clt0YrS3Ao9FhJv5aCKEmQFD06IX7IVP4hKZCMH+u2juDO+3VUkWQpzt+3xD
v3X3F+TZcenpdHd8yXtUxrbPapOgll2sVCei0g7PSQp/TRCMaMmH1NzhSIFhJpEs
hizH8r9aEZzp25S1pER5AnOxnh6Wc4t8JV1YXMYYgSPzpFlXtlH+ZvYyicZyfied
XZNfqQchR0IVva2xExXG/K5qSZVlqp356C9+VIpZU7Y4vXzfIKe9T/MrswORdfg4
mbjbHI5LnmJ4lQ6KGuI2pmPggNayKKDSqvxbWcaG0U0cBS6HxT6PKe9CFg9jGPgY
U4cn8WXrVkqjFCM+1St84X5CNWzCx5TYg0fzjcIfKUrdwymoeD92D1vBQkgiqlqC
QrBJhQrh37doMSICv+SDYvp/uTUgT/Ukpa1WOLPqqbAdptuTMpd/dycioeyiS/l8
DUT5nk0QG4gjfZP63YjqI6eTiyPrX7oCcwJp73z0++VvkrTvQ2lmSd33gqqKBxsd
Lhm56Nwt/Zz65Nwbf6jyFLGdxaHMpyasOw6ERw/TYmguRD1YIdgwqkr4QVdVvsxy
qvww/tto/l0vjQrVRc3Om+6FfW/k/jLIaB3AnszyB7OeNmIEYDGSPyp9lJq3b2e5
nq7VJBgxo1fsWS5RfMuTp32Z1KqOzsKoq+mSEAvExfn83kTuwhwW6Htpf2ZY8mRd
oyP2b3rhrDD87JHr17ErdvV2NU4qciNkDmkXnE7RUP5OtN4BgpTeDE28k0YfuCpO
kAeRvPlCdtcndxwfuFCN7gC2PTfYAIfm3vWIguejgkjXl5z/NESKP0Ii+JaH4Q0d
PCP6GMXKV5khI5lQhyr0dYOIqBCcLup1bByX8y0Ih4RG2ELplqRSwugHekPWPrR2
V2Tcf1iJeMbyd8lcxEHZM25vSnVZMwG7BnZaTDVsw/9Z4m5qjuy0tXuifP2hdsqN
OtiOfH7KKk88daMrUL6O5IKnD/CMYuvKoRKUWZQYqhiaKBKIvJGOllEX6w3bHgMr
UNGlbKpIzKSbZxv3Lmlj51x/VjdWoE8ZAZNZrg3eolzztpm0Uo2IVO6WV7MMZQFx
upJYKPRku+FwjO/w86zEBlneHvBVFS/06c7m4zNBdUDBuA8VjO6SsQa4eM2pWJgx
W/pz3xIRO2g5/meC6/crb9NeWhPd4VcgCMG0DB6Ai5dl0jSE4xjsMso9MvnK8AEa
DkmVLmaqkbl/Ds9u6nxXVICRejyCiHg7U7zxFo+v5D9EOHwuUD7RZC6VvnUUxa96
YFdglsRQbC8RD/LlB7tnr047st0MYFgVKnC7XajUrHeurkg/+z846juGuQfLQfaa
QlI1lXd+24+sZQdn8ZDvwx2So6cWPsdZYleJtiu1Vnr/TONFTpyVqpCCgXr50XUJ
7tNTNdR8kjJCqmt62xiRXB7vGPXw11zMoOEgRI0ILHQvrANPeaEl7xRYHqTDu3ro
zSSLo0L1ZapP3PGIPFqS7QAZUkaVVPKIS6ZrYaOKkCuEjxeGJYWu2HKTYunbJxs5
Og3EwHxAf5CY5h2sKZ5do70VMwvCy83wQ5oI41DqR4wg2LE2xavhX+ZJ+QkpQeTW
2W2nImaDpQQP84Un8aRDICU+evbCY2igDIqyFOGhFYWqS9H9oU3lcUnNRihyBprI
JuEMH3qrrBeEPyyhZIoK+LanQeIVEQmpb85wTLCs//j+W6y3rI5ZSN3uz+XAM2/6
DHpEy/Fb8dMe93LXiNpQ1RkpSgAbKx0qDIAHzQex1LPQ56tYK2RvTi8WB4q6dgR5
PrGpdq6jpiSbHl3GwWQ4ZVYUnEntzAjN3D28fuks4O+Z9fQLuE+AhSZ0dvDarSI6
r3qq34gpEZ8unmJ5t5kbASY/26oE2wrsq6xRAqbaqS8kFHnVJa09514uo3KINSmo
0mxwz9mj8C8n5w6EHDTFrRkcFDoUD0toPRyfMVgFmaaKD/cs5L9xMONWVMVdAZYV
J9lrU5mfEhaCSJosvNnnjp44m0ctZ7829BQDdcUT4v5hYle2617T7TB6QQ4OpnPF
RsLnGJ7lynVAmGsd407yOB9wMjglhZrgWpRwsKA7HSGnNg1etAZEeftAzkqTBfV5
m/pVbKgksVQ5TBtUVWM1hDKxdnWZHAwlfM1eX7XpzF7y5kI5bAAHENYVAOOCwx8z
Orv7IC7b87vETj1QUSXH0YLdu2qpEjioUnLozxxfXI81bKfr/HXzcS9sRE+d9MwA
wVmBMlswo0ukkze7JlF8wPX+T/Nmd+JMVusXrU6Ytqr3i5I17UnQ1taZDhVoUxtI
AmvexdyWuzCfIvuHq3CJYpw9QZzqwDKzlUDWVnhXMzHMRk0eyprBmAm6dYFhNpsA
nW0F2SMPwslpgkB/NcJFwc5Kzb+t6TUiS0XKtGllvwsw8deeTy0DfWGVo/+2/xvS
7sPvKIrcNIXU/RIvDxhLAqw+l3NNYiBno2GgiPZHAD3rY7ccyVzeU7wEJPMTXnM1
vd1wouDC6rC9FqvlYhfF2EIJEnjdkcEiHMEVvZ/VNv9y0FJIalfPo7mMYkMNSl+A
aBBhFO/3Pd55DXoMdRvM012+IDx+C8opAGrWQWcM/K2aUWyMGS634Zj11xni1OuG
dmx1kBqiIVd1PIiYvhn7mqWd688m4zll5ynwUm9FADqipt8mJp1H55vypjF5oWC4
comUKVqYGUd4HZjFsCuynOPXaY6fB+Bgtubl9RWaBT3mnyVb4kOT/e4WDsRWSw55
+ex4acLWSvkAdbQtadOWzOmwpODqzkFpoXuU3RZOo7ZkqpwMXZL7LOj+llQPhBy8
zlWqXX45ro4ND8rrKXvry2LAMyS2E6ak6fv0EZkGGfWtU9HkwCX2bGW1DBBQkpyE
zmDLkxG5Jur1SGDE6Ve9o8HLxWkiDAQS9OWpHyHccTEWdLAaEFeLSOidWWjpqepp
AJvOm1TNJG87/cdhi9aUwhSF6h78UhRxONP3W0zrmiy9urVFcMQ9Xtho7ysbAP9h
PE3gtzSLHpknS4p5TFi3nOg/1ortprodcDTmfCBDvGulftHojZ1GyqU6MUQgw7Po
mW592tBhjyuHbfMvWByAeLGCrd5DVu0JE62UIi5IawhW2GqZwyRnbJlXGRCwe4Bv
/ezKZ4NYvoofC1S7WVe5RsCVKlkPxPP17VK8mNW3IxKpfgqB0ta2PX85ipmwRK9b
q6dkIYkVtIqhfI+CfUyySgUoHznPB/LAk4KTZHrDWejqGXqrtL5xUMpGpbPNIOR+
8jGi5CWPUrWodaUbFOFxBL38zpR/0BdpHWfphrCWPXtOx9nw7GpauzN/1QVDx9iA
8OA545xept9xdf1CBD9xn4dAEr75O6NydHK5n0EvEGmadsIX+KFq7NXd0iml7WYL
wplC7jh81sC8B4UISPOO//j1YpeUbi7H2QHA8QL0ekNt9gFtUrDIF1+92Xt033Q5
/5YbNJzBTZ+poWk9GiPBZ0alA0VG0gqPDuZnhZoFQhModf4xCAL6fzgxfdE9jTwy
W1/sZzJawljL3J0bjvisC6E2diPaNvvja9SWq6oGPjTD8DUDErckVWfg9wp0zwEo
6KTqmNKf6iPlUHc8AEYGF6qCS6iIszxRp5OEeFiaapxOipMS47v6ecgManEW70Zd
cl/Qzn9Ddg5TFtsNl1YrcNhOiDhsNxo7cX1RMhQJ4ZDHJId9LnJMOq7fywvvmIlP
j7p90F2ThyGY+/TDlG4J6Ws0rEQimQhIkQg/comPH4jSyGoCR8ikom4REXZ1kzv6
uxbTPIIAeYG9ybr/dNhz8UWc3+0O+hmZvBhdUmtjfv0lPMVWhIG+PKABliNHDlCt
x5xHhc0VnmhvpPCRRUWUxCb3IA2bCDFjxDZ/wTHnJ0KAe1NpBALbOcapNU+ZlHOM
bsMqZMGJc5IP8nhbL9KoageO6/LdTmeWwPWpV4wIJl9ndjF/g/SKV2jkvgOY3C+Q
ZiYplrCJwFM5Mj4TQ6Hd8FK1ecC++n4K1juoDukCyKTgDguGNca3u7Xl/0M6I07M
6Vi+8rFlwi/YzfZe8vMmZUhU5ss45wdrptD6o4E539FHIKj2jW3olKnHGtZp87q9
jVNc8FR6f1pLbtYRzwPyGV0G7hZHmn/ckXDqhkH/Ds1ixuRl+70WYTDr1b0aBp+7
F6FRv/gHZSScLVpvXeiVuV72nwWuZq/wLZJ1zZe5YCEOKMgu8cmjFynbNMgSDnS5
QlJWosl5A+a7AzyYyAZA1y3RWrCFDB6pNqnsDbkPfWM1cx/PgRBiTsMYe7HTL6C4
ePLUBcbKkELzK/GVcviOaHAE4glO/qT43Syq1dfRuLgxEAqKgivmJoc3hKeJrLmB
klapxjvV9s66SAwNXGkIbKTyY6cRexQGPkbR2mYoVyaWv6QpNyjXMt7MFT3veNst
ap/DSSKpxaK1//fdQp3jcHW7KuaSVy8B8sceOwjS1BQDom3SDv2CGJqx0UuyEOxY
FOS4Ecad3T4gp8Fk1RCuamHHIKfUcQiAzlaINwm5A1bueBXqbvwcNz1anSBF1SuV
3Vfol2IIEL/NwBkMAlwDGT2MKfr56n/uqSNztjk2lEUil49qB9YbWOta8QMYJSxc
hgx+cu/IhQ43+Rm5M7VlqLWy+UKeom0KtD5HLAyYMKFUw5C7mV4HRBU8UlNB+sgU
x/825ZDon6HEROZsjr36ekIvWKUcpmpO3hEztCPNjO5mHSIsncHdkhpMJny3eg3J
eWxtgppGMZ5EVypSX+9LTIbxVRdK0ESuhbSBHsRZpfujPLAbXJitF6X2BF8bg3LS
Jls1gxVudRsgxvOBHwiG3Or/tYHr7UysoAsVp4LK+P8idhbtfSui2ccR2OvHpR9m
e6U9C8mDxJbdi9GxW5E0ESMNTYOBY+aA7aqZICWZc/nJmGb24tKSGZFaVGWODL43
Z64lhhCs2SPKLcIlFpEdT2LcFoYmI4/TPhcIM+PB5OaHLb87cSQBDbzmODytW8/z
sWYA/AWHD1Ou7CWW0XLcOSe+aP36uWkhXiebCJ79geE60xdWcl1u/f1jiKk3DPyx
xpbOkJHELGHdFvy3g5zv5EaW9Rr+UxMpjgp7KhmUJ1idAz7rmbe3r2O0X6pOwpwG
prOWJ3vNr2qvnWukLTzrqefrtOt/DelbwIQivrukmT1CVyDj1xekiIwaySbp1+0D
+Ws/Q91xl8IZNpMym0sMI6eBiAfzDEN7nN25NXlgGMuyQ6o8lBKF+RgNrAy/QAgA
20rI54CE2oKhYOcZRgMe5NHwIpGRJdHHGiwLfh4EWBkfkjm1rnXKQpIfYBAziqQH
sAXmA51Xhy0oPrVGirve/jc1FQwsG35mdljcKZlurkBpnzlRowo4MsJ2CLGipkfB
xfspn+rAozPPlvNmlGJh3Z+4IAgO7C4zn6idPtBGzVOJLtEhH8/kZgpyh/muHhDG
5QwErydtFmSQLfKXDYCEMxjQHFLJpAfPbpqtfS0i8qcsFUqVUIrruE7fLM9dEpCb
tI03Qzk7z3u8wS/PTec68Rx1nIM6gXNRhOsDOEkEIyUiSmVSg4dEhzvfDjq/z1I7
U6oOEWqJcl5VTWBOEUitU6XPoYeAcohnIzR9qyEoFP4wrwKmxxIBgebn3be4bUDm
DFIpP+bp+VDdjzWgqwIbxikeonYvpGRFEnfa3erE+ZP8IZaooY0CKZyDhn5uzn+/
5yli8s1sYBJVL/9yuTw0rrb/nlJQK4X2k00wAa7dxDzzenDe6jdk1JFUYT/TWkw3
SPAtPFBrmY/VuixbvIXSE922KlGz+ghBl1h9nmHLjonvV70u/S7lLtyEJOgxcYGv
o4BzuMjdvjOxmKhkZ6aIKHHfn65kQbNGitf8kCLMGenQFHWHaMclVhWng0Yip+rq
XLkxY5QCaozuL/tACRR33GXpHbDFAZs2Ns9dc34c2kbTjw/qmWuaJqMwArJR6nhc
kJkdylyC+PQ1zCUIaVW50valb3xxRmYmiIYiJKtMFzKZ27k6gQl1tklocNdtvAAR
LK+6NVdSd9+P8lS4pUUcqCWGD/92zVGRb0qTHISQp3fuGSoV03V0dMxmF35MAFV3
J3HiHYIrYY90+sJFtD6NbPEi0RnEG6Lggzcum3fMnbHtG4+RocoqNRV+hEc8fKGC
9327RO3amsxi5gluZZvClvCs+uesA/UDnVYEB0nBQoN08mkCMiW6qEC9nr5Ffwzz
6GcbhgeV0xOoA/K/3FwCdyWahZ9hmce7VqYMk1lzQ92so3LomNK8/Xrxewd43won
409IwNW0nvcqzLgdP//i+t6LUm8o7sHeoT/lcxaW/kNixe2eoOjrEAz5pM+35F+x
Ae+/AMzjc3GmzW3NosbSVtL5pww8vBYmu8QYzOUMjGm+Kb3HeoshjhnDiEWOiO29
jduCJOerz3BlFV3Cpl6y47NM49D/osQln9/R2lM8YCSbocJe8btjxZSoZUMmvGpR
rS2SWIPqQUyI17xgPKa3TM0wxJvdeSj4vHgfgSaOB/aJQ0OoA/m5Fd4NYXKGw0g/
L4VQ5szqk0BgNWgFDZnmz44kgPO36Wr66aun071cWsl2JW9GznuWCO0fHfV9oZ7V
4TBRmEEuAIsIzVV7h+p6bkcfrdVY+xmJNvH9Ys5PgJwsdZ+tPZtJaojVkRDr8qr2
uZmpMSYAbnpRLxqnTxHBDO6k8j0XbyuC5+pHrTQVTszhJvLLjUTUy9EKm8vgVNga
UCrWbXDgFkj5ZNJ3gbr8+/70SFMZi5PAnFKb6FF5voVHgWZA+63HGJ9LMCLhYq2F
emlFnr4AHCAh7DxpqypAi5rPV60ycoQvisnCNZUjnLasyOVDi0o90CwMkllihnwm
B+MlKEWYw7A5LgWIEBDujYXT8JbTzbpExHn0OAyzpJVfRlq3h5VUL6bLbY2Fx+nX
/NcrLRVjJ5Dgm+9idFdc4DVF4Wj6yBihO6kGnD9jmTw5NVCgErKpRYkrVHsEPEwK
XWJ+OrT3vke8QBId3uHbOS0erSrhjs0/ylUjY+5txuEAcFT89vXPSa4+svtrZLWX
vNrfV9cR7vAtTEXGVSvU+XUkMgAyReW/8im2aoYXyvBDbKCGqBjMLVyJjFk+k+O0
OALqXcl61JNMCO0SE+m8wniW6pVjuICTl/85e8hgMIjrtyrJJomotOw9JM0wG+x8
Rjxm1HGm00bKzJQlKPxZLyV4kpNQfdG18PocvUbAEcAJkO5vdvgR8PlWQ7EhWd/m
EgPBJxP40+NIec6RAoMlg45me49D1OaV/T930KVe3LT3Y4X11fqer+G9k4bbI3xx
ywGoFTSrgzz+oQHqWANyT6lklC1bVionUD5nPYq1PAoIWHHd6ouQaO4KR8mxMnGb
a6+ZRduuQUrIgBZlM+VVVg1whLHIcHz/DoF3CQVVXUgEx2JQrf6wnVC0BMlIMV39
LGBaH2WZPQ8aOFvo8jIWwvhLPPuiNnr2zwnb0hr7xKHacr9k87uulbM3unhuVQ0e
fqxUv0wEP6O3SOciErjVQCpeZOSZv4AGqJSa/0UghsjGi1NCXZVaEA8RRFtkMocG
q+E376Jr1mzgzWrOzCheP0japm/VGs2wlCqKr7vOI82Hr/mK68r+r80YHK+0RFUD
OMn4AzscNebrTdAsLd48ffftIYvKZYNKS02aIzMXJt8DboGcCAqjTjdgSdWVijPb
whsdu2agZi+G+NTJ//v+6ToCAfrCplDfz+dBeFf6cpRZha9D4q276iJAlwNnpZUv
Vl7WG48fl6zlSTxRAMN5mCWg2ufWchaATc1o6AvxPEqQ73fXkvy+PM8aQFsNB5wF
iALGyB6IPPyhTEgKbmBCz3iuAZi+Qzf+pavYDw0dbGowfJHl+EyZWz7ZOhGy8ycY
keS/DWnwkcQDKn3Kgd3oLPU+P2KlJxGV02o9MSLErvNskcjkPFN0zWd3YEwfuNqM
s2SsXl84boCvKlyrSzHN7ncaS88cMUP1E89mx2r9tiXVk3KAQE5jFB4ZAXBVZdTh
06EOZturqtxDJquj9chFqoWbQDL810S6Z1kL1ydODIxD4pRpeJ6yUOx8lnqu/dHb
EYz4yYWooAsZYo/iaDoh+BI5t/wI2IPT4M0+V89cLwGYoSdGPrWda7uf/lWtX7UV
h12yd3T1tlCRBCjcN9gT9jWyPc5oO8cYAe8rs9afYENgu5bGqFmobWZYGC2XNMzR
VKgoEXVVyfRujABZeHdUfESQx7M+B6HIPw7pO7D7jO5fq2O68cOmP8trvFRhN02l
9zy9N2TUGx+oEpqlHE93M2O+PCC2OmXYX5CNnbtGyZt97X9kr8gY7WE1zV2McU5g
uCbOBWBGxl+enWIUqjQE14tHss4DL/+JLmwoUDxfcylNWkTWHH0/Hql7FQDxB3X+
Q1TNAnX5Bp4R4CTfotHAONWBz3IkQhdDJHNlUx5XyppvDM0/lPEokloPU2wqMc/h
BwEp5ahqRCyG110HVkGmjEX7SX6PAl4XnHeDOKARYQuePLzxfjTjusvaI/mP24oI
ZP+5KO5NxgULXajSicH+P3h/YQClbu09HJ2rklbtIjk+GlQ3xh65QbmmbrLTmQOG
pM5OUDGLqpmsetAzt4p2xsSEmQu86KDHxOV/dKUqlJ0olUSzSo1pCDn1OTcT8qnp
kHuRxghkjVLuwjuulDQ1nVD0c5EGLkHIHRzamORQrNnuq2JOe3gls4WM+ng3C58l
DWyr91RNnWxXztAwoD6DptqctdBpka3ur0Q0mK2xmINvH3m0EFyBHigzwpW07DNK
sGetaaef1Cm1kTNi8fFpuKM/KIHXV5F+XqXXGp2DeARrFON/TSCid1m2C+E2GvWJ
3wW1sM6Jf1zh+RPtA0Z9zMSNcPMzStqVKJt1hKQJQuVJ3DwxPVyXNN6+E4bAGTTY
dRdXQZMwRSwYq4NTVrvzKxLRiAxAdT0NfUoz+Zlxs3R2SZaUkFguqzASMiauHGkT
TZ8Bx8vp2wgpNXC0rFSuqtOusDH5XtroR99RCOmBzFifUXilaw60XhdwK99chCSB
jZta3L02oONMmW7egjZxyzYrNx9zRO0pca8fzURQa42qm7icmuMqRR8BnpLyKyR1
Hf0cg7MpcMhaRRKD0uNe/hAnmvkaZew2rF7KvjGV3AoPviF4GNt7OePo665WCFom
+PuUF/+bP9TMZckuJkrkEFeiY1ngcUNnG20M04ndMymSme/phmxRJBKvGD5Rd4EY
OnPIKrQK9ZnoYasHvs2JOxODCTtXjBElTwTQGatg94a6RB7UOnJSCHCuTTdCqUuG
/Qz02p6t6TWfYzUkdFeOM06Qq6mpbHYFARnLfz2CfPFiKkdGTd2Mbp5M2RAuQYut
BZf6LqcuApR9cf9mLg60fRQ+dK75q50+M9YH7toU7ZHl2fWFA0pv0JEwTbaT9nwb
lR/tvbq7+Qc6YusMB5q+LqJXRipxnghLpdAOb511Zse5O41GlGu0C64S6EJqp3r2
IqJOYS6u8L5eDL6L+PJVQ/ZXqdoaeuxuJ2Nd+0vmyXYU9q0QVBisMPQCvKqLSQlx
OZ/FgY/IWm3e3pWV5+5Gz7FbhUoxSe6LIxSgfNjCzQdfQlixgIpcOgeF6JFJ41rF
iu4WM0Issx05ZA7FZXETbV1Fkb5ERSK3BC9fqm7bPw9T9B6FpBXPUEJL8rkOhVpm
yXPXhFQGVvWw0KlTpMZ48qK5Z7Fgirq5hgdBnIuKtEE81yZrM2vE7aMF+0+kFbQo
fwMXtxhQ2qfpVRqq4zcibKc6JyaA9+dvoFA4zEpMb2Gi/jxM9PM2GtKd01JFZ04r
klsde8ZPqTsu0mJ/s0XLxQsikhMnhQYpl7s6VLUvKv8DAaPcZ8YTLLdBLnjEjGcL
JtRuM6qC2SjP/jD3pvBeHAqMyqevKESoLoAD2av+XF8K3/x3u0LHRruE0TEl9elU
v22t/wMU2vnp4anmrTo8YY1w0ytzADuXKU0LzsyVqio4xAKQotWDQ1dDBm2WplEB
INb8nzTpYiTJJKldWE+7af0RPenGNCkr7HmyGEpj1iFnhTiQLfz358eQa0yEIJfV
irsvbwZP5nO2r07NBlFZGUFWFzu9snZ+o8qyWYiQ7SQQO5NbXSENWrErmwycH80f
EZNtryEcads2fZWiT2KF68Ms0Z6Azq9wzs85mQ2ablSgeK/r/BghSTZpy1+bGTuW
avjoQRebotvTAd2uoQwT2EWDaOtl1hUIKJjLFaFCuWG6yiXB0jxoSycXqgxJZ3rN
h3Bp9Q8XQ1GB2bj6IfoCt7yRtukjrhFMJtvTz1krs5BJ22PpcGS5EKCGScVBV/pd
rwJRnyKHmR9Kzqr/8NBt3UsVV9PhF9RI+gXAI8Dbo13OetEghYTAlsQPLqF11gKy
dUsnVeKKZpuSUrDTfTpp43+1BmwyeFOcDftWDs9dh1h4Hi36hB1v6sLTUBxQHhBG
7tWRx9hv8cd2CZeYH8KksFNeF2bRhq1VQXdbu4yvxgy/bJav3LjAb+jD1EzZlkum
8gC1ndfzguegGwoG9WzNl4WggrXYsKWWqSCm2mMlk/tmaYPtSP6HKcJ4Ax4gTqNL
cyvJDydBbYBlsTuqOemBwP3HZp/7PyvD4kT6bz157Ej2pJ98k8rlOOFYr4/XCxEP
EHwEuNRsERDFeEpxoBMbH9sdboH1vKrqQkS6pemPOLG4fmXkq+8ICAgwc1dmOT00
LlWxTdyBNI0vszyfJknzTZbrhuf2eGTo4sBdMvId4OSw5Je9QBzSZyuMyACaq/9S
iRV1I1hhM/s052A0ZQ1L5mIXVtIeF7EPSTr/lgnryo+A9Z/nlEgx7LFujY5LLVex
727Z3NMh269VJog7IiScZ9yjhV8G+jKY335A8rrPKeiN3Ao5klIib49HLGoe8n+0
MYNEmBJ9PtnDGFm7bKoEc7PAfJwFlj7Rb58rLx9Yw0zoyKg85YUjr8PJNt991zUa
5H8XIADXUrKIgRRsryYT/SloWdnfArVTQaGMhyBwu64dHkFnFOMAF0DTxJkwV1wE
Hik8iDXRaCXQXYY8tuLlN6EjYEwnB4xN6FKqn7C7I3TTSwhRxlMpmrzbLRK4PKgO
oS3jaa9DLsiT+Bsy+d9IWpEUBw+Ntpu4+lCLDrlv7n6o8jMVVOH3vrV9W+VFYmQw
av9e8lcSmqdN/i9FQWiX0Hb1woxNMEp66+7Il3jVZGg3ODT5CsiqkjxoJTLPA+i1
FNQ92wNdtZrg8i/QqeJCdfJCFxh+4BArYF7PgWnvHJ8/aGIlHgMDGfDgQSMUPmoa
uwqxMkVAl3w2IA4lob8vb9U3DBFmsf4T/HWt+aRJobunwIzKsmkZCQq/gNAe3rDz
hVr8OIBJ0tcDM2m9BrbGKi4hMU4Q6yUOWdLkW3Hnqxz4WeBMEfxSJ+9SSBHkcNDR
1n7Zkl0gK+S3+bpMGLdxrghcL+ov1V3nVmrIJ948CjNDZKNfuZ4Udmua56V26a8I
TgC6ytjYeACya8oYD6OnrRaTAYrGOoi3HXDqoOpChOq3cmZGQFjW9Ij94TV3iEiX
5RfPlFrYefLRywXGtLiBITvKit9v3gCgM5Z/N9tlf6leQXSVcEzOtuXOL80jc6h9
h/DXerw/hHUyR+ttL0FNYcB1yPJTbuAyoBRnjkccKRJcq600qcx1YIMowXwhxvt6
1zjJUjxvCWTNTKVvuG/CkPjlmwMzX94BDIxWLfK7r8oj/EHNJFgyIJlm6TEdHZ/J
XY1wm0l7cF7dNeFdJOI0Jff3oM28KAoDBpg1PCicyeKMuAE6L8wTtw0BVvnLSuOQ
kTMA5RMWmq53AQ2DJw7TDxFKhBGY27xeXWvdP0DNf6MkX1rcdDWxMafeRkiDVY6f
Ui1iO/0w4LkIs3amjuLU9d/6w2vzk2OavAwq1Y7QiUXd+oHG6xfL+cZ6+937N2T2
CfPR3EIrhw1mdWhX8Ol7HFsDnT9kTwmtYZyZ79ABuKfpZgHcsm2qfmQFcm2k3cWl
5r9xno969V1W9UWUnRQvd5b/kZ8mETX+U8uq4xu5KLuTht1z1vi6LBM3pjHEO2Qw
lvGxhVnpZVD6V5cez6N3+Hrqqw+WMV30eKjk6ozvUT38KL3axibzjh7o651mvLXo
FcdZaUs/UNaRvDLDyoJ3Ohqg2P1cVNtqeI+NG1U8m3Wu+lIAjxtnoOWXkuffRRdz
qFAbJQOsxWTvWYij9ScTWP/zWNsX3qt4zX9QnyUhsjikM+b1EU93/5BhuxbPXIQo
RrEEhXvs4AA3odZ2g0zQebdcTjqNypEOlke/jcMctqi/Ss8f7lh1yqkAWXXD+/wi
Uc1O3L8Cq6dL3oEENC8HAA79vhyV52YNQmCyzjmq7skAcQGXc8pixa2ksCxONJx9
vWJYkZhmpuNkdt9BrPRKKLHvqOazP7ADUvqtw79DN0rUuaz9dHaB4jy0SxTHwN8E
7+AeQwIyCj45vNtZkdcesrto2KxX3cMa1+UEnnB+RxWtwEfH8zpfgGhrHP/p5nN3
iSgORfj73AAtUgADaeDJf/G/M1XrhcTazdNEezdaZbzXAgPn+lYONJcBFAHgEu0+
N9bsx8ew3G5/pb0QGTvMeC29EcnTuYFx12UuHMRw87q5M8FwahBaP082qAEZVcBi
XtIlmQvY5kfKMLsL0dhbEnkVWVnP4zUrR65oKQmnjFjHhZ6zGYPmPWg61kUlMUKe
nVCveB7rixKyaHpm/93/BgwqUzRMNdztWNPJB9pQZ6rQ7zRnmtoMLXQLpMX1oBxH
sWrktXNhctQEQF2CO5xdZilwF3JUbzPtD024dn9H07e05d6OmHuOeZelwNnIhpuM
0/XX4uum8Udh8k+Q/j7+obsdkSy9bMFIpZEmPoVUAFrD7PMi1qYrgzXHXwJquAta
s4Ktkx60kAzLdS//QMMnfPHfFT9SdwPfMn1RFXhzdkiWtFXj8oGKMVVXtLzWTxUF
cmB6ytPdX+pOlF51z5zbUX0WoVH9btN8BUtIGg/o8xxxYMdzZcmzCx4XFZCchKyF
QnNhlhPw0zfZjZy+4ScpnBJj7NEmp237Vo2QeTXtHXzHPoIlCq8+yr2J0DHPObKp
hXlQnciUBZHaemv1+kWeHq92uM9hotfZylvOOo8q7LZpVqcjnlQzDtzgB3cPpPTb
sb/NZmRAP7bVoqY6IyIo9TjXPN2wX7irPXOCZLj2F98A9dCbc0hj3CfyO6bPykUF
jcEbut3GVIZOjbHrdMkyfnXUL6TP4NkX/F3tgUHR9DUsIfnF4I2gSOdnlO0V9aV2
bP0Tw7SjOTlsG+P2ahm5PEW6oSthDpAKeOjHItMY7jAuRBUZ/DnEWFxwLs+5/G03
JK0LM0RUPm5XbgB6p1suZ3IHcMKUmXrVjat6V7pOnq1z4jPKG5Wag3sA0xOZgyuk
amQLplGy+hbI6Q/PXsBHGXPdD/7R/IKvVw288onOif3xMD2Tr3xRNb3iP+n3ouwH
hcq+N/XQPRGyE/0UQFQoBzG2B5sySXE1KXZ5ajhfWdtEMULggYVlkn9UU/ssS0Js
B++Hwa7pFnbEPYRiJcFXTxg59+fULWAWL9fZoL9y5Ra0ZVi1kjMa2bA46W/QToQ9
UADlkjePmJxz1JrHiNNauO60qiSQfkKuYjBbs3O4xslBR53eUaE7+9rnXui8IhlZ
ENocLkKcXhp+2WYFNk38bVOvsdSkXF017fh2FEGWXFpwiREJzkUmpzNXC7XQoa+n
K6S39yUzF2FJpYk7XrxEkWN9AkFpFWDUxk1Moz7GRLf1rgLl4hdYmHih7LbLeI3K
8jkQXd6/WrO4EVLvrHDJreZVTCRffUS2xm6t+/JeaT6sxkabZguCX+8V+nNnuH8V
ONLr5ThuvBl8TAIMQc8+X0KzGDSccEZlDvPThnwdsyUYfSDKqpBTdlxIpJiFc2CX
DSzBZGeO78xM0Q4lGhooxvW8t6Aet0FPaQ+siGpkcleX9UQYOu3DbEFp6uZkPijF
gaHqaoN2TKmJuG542INPkRZxR8bAcugPbrVm7XDRdciNjo9egBn6Knymavh/X3It
4zfN9phg0U9otTr8139LWblXnQ0SxiaVvzx7XrvdYUvLf4CuTG8yul8LVDbCfCAN
y2BQfbJnY0ajn7dhzpq7SSTSWUx470m8iaRsNDJhaXm7Wk/EnYJOvK3kBb0nNxq7
D07RJwvF3CLv7Jq4Jd0Oko8GgTQsg8ST/iSvtmaQMcTE24SUO875Lx5bMdnTxdBb
o+B5SNdbITxEzmFnGvGATTI4i0aHvyp8/Iv93SOO6SdrPihukv9up1DBRdAkyIBR
pAycEaplm8VTfqdfhhSGLBFIX6q//bEDITxJvGEa24NYNeiXeEEW/zkL4NFnnMNQ
fF9J2R6icZ16l2p3bF/+9yvc8uqR/lH2unwpBh/V2xS2qp8OprHR8V7zeR9Ag5/N
8c6WXdkrjvQ/eTlkxU1qjUi0KfWU1FP4ZFsUdxqxt8PMOHM/ju/2ABeKevWXXC9D
TxJ75Lqc8nRRqLd/+r+vGIxyVlxBeg+bgNI85o36kBPbHCHU1OmOW272yCpBvO32
3v7MeWFAdcFiKpD96Bwwexm39li97KSkughp6hCRmxjm0Tmdfhzgztrdp8HEguKS
9NZduKnxXiRX98zD3SF+PkkW1bjzMmW1voBVOhHId8IIoWUrTayOtatXzVjK32ax
fct+QvdtHvfeJqE8gy1sy+bNmzkMXka1FYTVWLahfbEivxIQ9sMnwkivOjnAAzR1
Fv4zblTNLw86+toVawt70p4bCx4os+OVOuiCaXfwem+FGwi0uW32wzfY6xqCrSeZ
1pmxChyqfVfG9Qqkn/S9xuaTLkzRpzajBLStKGRNlbH+/75SFm4AEvTpIkqp1Pw4
Fq49FcC7kVM2AMiXuih3yx+XBBfyCyZ1eJ3jQ7I+VoEpdloOaIEe3wgfFxelw7t8
i1vy7kjW1jtx1dSQcxGvp7Apk8AVcN9WWKvDiZrEi0w0qWotRVC+REIxXKdabQxT
K0/hEZcTfCaYAF/wEhz2hhblz6CIuUo1eGz4RN/B0D51WjuOae+NkjLZaQaZ/CRO
qocE5QfqCMNbppkN3M7PsMp4fRZRHm7DhBTLt53+C5Gu0y4tsGRGPN0hWxJzyZ1f
ucr5L1P31wN5/FswY9Ycl1Abv+WP+Xz1PAd/TFy3PyV7hcYA7L53D3yCXwJr96Aa
5cSF30VP0s6MvdsfzJp2ksyHnxSXHgbI3S1ia67h6ZhO+LKcoeMRJsC+YMcm5TQ9
eYROZ1ZoFS+VHvOxhGa0JRAuG0Mec3BLkzOTLPKEq/nuxQfqrNjZSTwuZVe/v20w
FQG9K9w5e6h+1m0M8tYyJhQUFghOV63XGzk1X2RJBdd+ZW8BDJAEF1+lBzTAOxXL
xrPtT05EYr61NHxvaeobsoc564ke5pYiRZaLSsKbeoRltbFhIRwS4U6dy5P57sJR
wclLZeMUi17spva09PCAWVIddsUrGa1eiJLvZowQqA2n19rm+jzqbDNmCngLjr1X
E1Y2mZig87lEJGhlM/4qtnNLnlAmy1Kq8Va4yGbmCDTJ3pKCr5w0VS1CWRdV+cvf
ZeOxPhmiCfP5fM3UpDRiCnH+qTX/HuYHnOmHo9UXJxS6+tq1ulGbn5suSZrYe6fx
xCLrgIJiUxHiSJtXYC6q6fSIz6jFmeO5Ekt3dswr6oussYDWUWnOOE854Bs3/6z6
Ug4jCDUgFeQISyL3+/RFAGaydorrKV8IiM6pnW4+uC7Pj2kOWrEFvm6mYpumjHsg
wtPlZFtHgjsElLjaQU6cff5mVoIiTOx1TdRsbBYpQIyJTP+7fcuQ6zJMMlNXrVpf
lqZsbzE7otDrc16bljOsXnqIq5ahp6/1t4Q6y6MeWU8InEoMpDEY3y27APuOsdfS
DAGAajq/1t43uk/6Gfdce3aL70nQSkdvRFAJpjx0GWKY1yInouKPTNb7f/CyRZFc
ilP9TvejPKKMPUQiKFDuoFRXafGO9DysZ4XCFPNP+kIXM0NyakeaAzGYaqskxGh2
KCIgcGbfB6XgVHlYMznfpfb50AGqHEiJbcrjOPNh9aIyd5ejaYGcciSxx3dRnnNr
wv4DM4NuzS8kSQQ2+Mkx7lEe6/38G7ssqa5kgdqzljRxEhA/erYZ26nmlUe6lCjK
yNY5PsveWVOEFORHe16xRi6tijFb9wLgCVuV9DTQ7/Tw26/5lIEU3ujpKAmY2wY9
EoMATJJf/h+NUKYP9RBq2z37P6JL62g+9lrsPQovx2cR5kNWT74uf7g5DFIBkKgn
5+WYoYSBOZBnXvspxwvFU1rsNW+/qz/WkISwb0RiNnIRjjWS4lhzFFdZVQE+WGtS
GZIYK56eiM9piTiF+l+iRTkEG6eAPhLqyobCrGmaxLuUm2yCdOe3qjTj3Qsm8kvD
BbUfWRy2okfzocayLivtfLmVOuM+IMvZSrTMTHxhiIM0F5gbPW4GoI5MVlFvOvDt
PJkRYqTelwwH4nrGoAvR8BqW433ckFS3CbGw5w7cb/WchyjQjR9+YqvFHo7yQga+
HbTxBATQG1K/1VyPUNIDAtjXroxxj9n8QvGGD1C0ChqdVEK5QVpj3sAewKB2A1K8
/mXd/lZP16Di0mQCkrKFWOtKDAYhsZ48/kXO803ychizEumRMlGpxT1nLeMZzjBi
KOUs8lLluLbLGGBuzYF4PcRYsscvQKyGsLSfJEDnwzhnvDuqO/wY63DS9I1l2vdL
1EnhqHHqX/1lyWkI3qZXjZndtZv/cJWkLE7kRDafPerYl+EZkX7rdVNoK0XwqUfW
tiWx+1M0K61WMnx2DCaYdX7qXZbKF23NEBjc0xZPiDVdeNUkojrew4Wi18vh6NFA
S92B2hYB5r8Cfygwqqn6HCcpT+nRN4mdPFVgY9RgYADDhPKpKV0DMSwnwtf5f684
GWWsdkQNeQN5yPjus/sJbvLQ8klCqXlRNB41c5vzRTq+TBkE2tP6kWpIUkLzZSCQ
y2HY63+/aVuVfaSeyu1M0qnHMPZlK1rCEs2U6hzyUa5CC82JjDu4SONSEqttysQF
pUNOv3PiIj6l2U4pBKYYqmnrkniFaA3FtWJnNJ1JjWe3gSsbsD25bbdxFwJ4C9n9
dpDmm6VxvBEtfBU9UDn8x/ZxP/88dUtkTofWwnLxd9gKvNfuyTQXRbZxcgp+D+Kb
bH3fVueMxRf3wHwrxAvbL5jS88xYZZdlE61lq4r85FIgqomrfUK3WtEFBnlPjgkX
uNowilyDJEEzXwXcA4+8HuBPDGOQq3iqb7SWxJrET6WL1CvjgTQIR2JAyTL1LCT4
UTgOgmDyCPCdNncHa8MV4xgMTFkK7ozcZbfCKsH6Jc64NIIsFFQ322ChfSmPTAsw
kNSbK0s86JyzFRSwdKCcP/QwcDafK7DETzaxDE2zrTix+iTyVyNyUJWjrF04IV55
Id/eoawgfdcUz2b6AjonX2OeL3/A6DCbpA9pq1hKVpl4zQbOMtGzb/3lfqGPrl7j
CueDkxOlaxcEJ/lCn/W8YnPFkOaYjehkE4pTGVS8CkB5dLBiPHLZ2LcK2QRmIDUL
jTObJmWtCLXfFq2j342uGw+Gz3s/+nxfU38BnUB5LO2Bv59limdx94er9HFXvzpj
yTpYh8egNLk9u5OwovZADJ0C54TQrREplUDwPkRqkREyn65fXF0YUGHNXiZJKKgZ
4RwimsJT1LYAx86WpH+ilGTY72FFRO6lfNTnOsFqBZHNT/3470DiJLxhnL/gi6Ka
vVNTSnSCUVCB1j384xKeHWxhCIhdAj77DZsafhtpBaBzEErVVAR8OMST4jCg+7yX
AmoBfytzLvJg2oQM+AusaR90gxxevNLX+fIaKAsnlIA5TpY4OeQ2uVrgPcH0oYqd
Mjo4Jl7ZIfiGH9+3gV9DXEnAZ4vSBfSPLT4vPIrGSPKtezxeN/Xs+wprBhNmhzyJ
BXhKGRA3ekkQ4+7yJCoF8oopmdTMG9sFEidyqtYNxKaF17prKFI8BPHLwC27zu0K
ir+XjSP2bRyROPvVU9B0kjkJlgJJ9CJsbWsFzgMIqQi+a7yniqoMCxBRIz/rQwCc
4yQMvgV8NVYkijs8KPBSTIwZggkTyCDQ1AyKqFebTQMni0OgZTp28bv/AxuAmngq
eLOdDLJES7j12rMPScBDSu7wjvugFVi2GbViMmLY+ZqzHcgwjR20Sxi2IgQ7Rt5g
g77Ubz4MKlszkouU2HWblMAxXXCgk5gnm1+PwCe1QyDmga9+xicAB0vX0GWLBzDE
Y8ZboNpfHJQ2+qk/RWp4x7UwD6kM/FdWFBcCUjA+l9jtcNCxq72Nres6OKxSlEd7
k5mB+5i0mWjUBdisv3fbXwZhgMuvV3I86UsJFK12WYhiMVbBH/evBbJSPf3NyT6u
OXzUzsK6YsIrHSykfjU+2F15LVt3BqCxXQGliW+ku93A6905ur69MKb6QOp7zKkz
Hb88lwliISybJ2qiKPpzHEIXWj2YK9qx3Sx91fPR8yQRUZB/FCeEofLeadbvrKBO
pX9h10F5Gsdm5btgdvLJimuCYarUVH9gT40IO2kRgjy41KXLYVUjc6z2yLobM6B7
1RNeGKYAFSEIb0RazmkXCap3Nm5L6AoufeYse6q63FCBUzd4P574ofDNKs401FiT
2Hyu5cNitXsWQTVvoaDO0bwIYGqGmzJrOBtFZjq6pVliCi8sFl8XhtmFCP1jwAxU
6xUTpUTjbrcgbvnH5TwDGRX8tSNVpw/5ODIpPOolIf1bqUaGcIQ84nZumErgdlCE
+s0y/W+P5M3fGTPpXt694ut4YRKbCx3l2r4PkW3kd0+Sx5Bfzc4KrF0NLLHhEyFR
hM8USTpesAWgz/M0i107BkxrOWyzmDNZQkQHONGJ8TY2eQLvMBs1hdqSQwaS+nJo
5+OmucGCsnQ6ZtnDF3yW2LSd4raOx8vRiMPfmmIUrZ843bwG9pVGvF1l0G1jshtl
DX5cI/zZG3u/K0SZ+ykM8Uu6ErnnWWO6BHFDhD8mpWK1NlcAd5clLIXN3QI9QyKh
J/ZQHxZ4lexmg5vsRjORErl4icOKpZ4Tm7vT24ePVbfpmGjfNzRRf7yvMzmNMXQJ
EM45VaG+K8g+ksiNWHsK0lo9nXY+mqNNpoA6mrLLu10z2UFBUgMPJGYMwPIAZskl
vosWQJZtLUjtUIASjy4M41TsyPu/+DbQtH9oFdiM9EP9TbeRdr+xtrtNIhVTta06
wS81XI9AW7iJ7BNrDqhCrbl4btsEEQ4nZF6Lep66GINln7F6hGFdcJhtGeSd4rm3
vYs21YmZmnPLRGbXu/UB8ZdkWcV8RFupfWrnqr1KVHl/tsv9Zc4cii0/qm59GyGJ
oqNjdCKD6E4hDhykZz9fiLdXHUQT+IkUrnpWw/AebNkT18avJXvRsh47x+niG5Hq
cjbOvR8pwFP7Rl7Q+gbdP2nM7S2LduQRfRZJO0qWxU3XB4zyPvNMdWHhSPDENnJw
3lATQe/Ida0x6HsNdNxriVel8IB54wl+Z8G9eLT2L9MbcXXLItaFtXWWLIpwRPjx
zaIb9HoD/u1qpzW3Ay4A/q0Hr7tnCoSCbsnwkJ8iDa3N6eWQWyt3EFDl+jaBI+CB
V7MsquUqLG6okFOBuzFjl8wAN22ZQS6YFUqHZqDqI5OcEErHnRVWcZInuTBfR40/
Le9q3zfSQMUFU72fZgVbyzlkdiznILWgD7VTN+h8/pvyMytZEVC/JZ4qn2Og1EPr
t/1ume0Sd8IZcIJ4KlyixoLDt0Rmpw6SDvVIqKCk1gh3VOpRc9QCT9bFudo0rYI/
SpUsogm8T2YdsRxSePxcqWodpoxR7qoMPT4gpagIFBJY17ZkEyIs9lbj8EKIa89o
lWFIuTcZq8r5GnzY5Q56P1cjMxaY2hitrkQYZcTnnzOCY7D7vJzDS3FAgnczshGT
YetupkITZSm4NfikJhotExpmhpZFKkjRInG+++uC0o5bV3ERB+f596SVtKTW8M1C
z/qc4cYX/herk07j0KvUZKx04VHEQIqtGCoHqRiz6b98exUSBgDHR6THUhhtrKQC
cPUsHCJ/3DRoWL/TEmbj80t8bEeTnfMroHjFGQ5701UHv/RdiiGP9z2itLdtnxQJ
rJA6Fmv08soqhNQ+R4Bte0DW4l3v5Fb73bJByRRV5amkBk2a7wzJaCSNwSUptO2K
JInNra2uJUBTwGD17PSw0euAS1d/yZdzAZCZXXl2HsJwkXtRbRWMoDGaMT8NEec+
BmTkxmmR8QzTLVql+wtQIcyQjgsqhU1iV3hFdhodK+w4ikHhcPM1C1qf5d8wJ8FT
wKk46Dx1+9xnQuTCAEQ7oXXKr9lCLxVckMImJLd8Dr0RVBuThdM9DHpcyMidhPGa
HN1JWyz9l/LaAAcl7q9jqjiuzEBXVYgUv6LW7BpUNvEJwtirPbU2TVAeDV2YU3PS
IM+KevGPCuG96jcATeUWd0e6mNvawLuwxrqNsewRlygW8zil6hjuCD1cSEe1zKbO
IClAAg8ZVGvWUYhpQeznCKuvjLbdX1Rg3Kb6cpJAE6CZbMEJf5HyFRS1If/QskGv
7h5MEP3Rm9x3Mk2PFEzw6VQTLc0F9gDlYL+itHdol7cx6VY0Q0NJNP/iG+ZlNnwh
EOMMiyh7JMHd3iT3hUcB5sPMen/foH0jNE8hxKopwz6F8+iTg+YdkFFIa3xmYwaJ
pwfQy48+4AA7CZwVKZeZHB66qirZzjeBXrLVBD/9VKqzN8+TDYL6Wgiir8vfyNL6
Psdwfe2YxZRNh1+TjvyGIQ1OaN9VLKOnoyLLoeXdTwUVthhcAlykTErLAv6rTr+B
NdGTqSBToxqEs90t7tJYVv3vuLNWCFzadIlPCDxs/nsCxx1DSg9yMbDQox5ipv7Z
FDTbw4L8/OVC5eTQMVCjZxRv9NIf7gPQh1GHLvnj+K2tigtOz7HSR33EM25uE1T3
DKoif9HVR0+rSdkCSVr7H6QIwTq7OdzT1iQpCNzqv8nk0JburinDhC/qNhL/t2Ur
DRL8irHU6k8/ndbmfvnI2aX5sy25qXjOaXgBs5JgYPBkeEUx04yVguXquEb0AsQW
REL4wCXd592kmjQDFgxHxZy2JmdNr1eXX+XEpr6//H17R02sgi0R+HNTfz3kxS2P
NKCmSdlpSKf7cfmi1/iNTkRbDQ2l7I2k+KuAbM46O+zWBHb31lF22f7BmM3ofggy
mmLJhFCNp8c+8g0o+0Qk13lnHyUx4yv70mE0yfpdaIKg9ST2ANRWxURRBoGwB4q8
v3nYgpQX7+RcyLfQGINedPkVlyRtJCczlyYpHpGgU34leUwR0x15Dpg1HOUuJKM+
E8yIg3hDlV7Rp6hsTq6QnmQtf474b38GZVUIfnC/WH4OkqjHPEIxiyg4GJRNuFS9
YUJv4lqRg/AiAXujFzEtsJfy2viHqJ2invvw2/rW3dTLmFiv6zPGvDck/8/MhUph
aO2DvyyBXvonXT2aWMZ96LzD0Rl+v8ZF09W1E18uLqPiLCaVKV25Gp15Wxe0LP1t
L/jSS0YOhy/srIzdrjksnM6NrC0Fw3VF0Mfa2fgtSkw6xWk2vqyEA0vgPXw43lnH
Jd1RArkhvUWu6+huQgq2vA1ljBZr3qKgN3zuvmOOoADS02WDTo+aCytKR3EqnHxS
y/W6QDDbhiVAeTsKziG3lJAXcKnDsxl2/8GVb0AkY5fpNheuXv7+1Sy+lt6iO9Pn
1tQncvcRLkLrmRcaXcmyiHEeX53XBxVuNHOt25hfOF+enauYb6jR1JrwELxku9rb
NF2UjQGHqbB0M1AcN2HiSa1t3B33tj69GEWdDXlgMCaHwfkZGzzjN8vGmYmLd0ir
3ygfRcAc06wJpxGqaOm+Zjei2y2fvGXtbLMPtOd5yKU5G6ohWsCR+wraQGzkN3Dz
PQ1UFyFID7xRPt8ra6/vjswuN2RZQu5IGKvuc0hmn9hYe1rYqbUPhB3MUj8fF5z4
SGCLqaStVASPtjqv3X4+1RYy2zniYCxfDM0h7yAhZPz1jvrGC4WRnumEl5l6eM9c
718XUhcwYCwhdR7KOkAoFzVTaR0YHKRSBD74lfEw5c2WX4mKPpR+uLlmfvWt1Ge9
/Vh9bzi8TkuJ15QPoJ/2esZeLxLLNYuKcF7S5xc4fNnVhHBu8yWGp5ja2qB5VGJV
kwzTRpy5R4zu/yVUcEfFQ4srRGMrNt/3VGmbNCZ6NHdcKqPGjAk3ViWAvY8/yEml
5zrgWxeqW6P2T65B7xcFK3Giiu5czDHQ1Je3CoRRbwL1h5sUbdbOzqgQA/59IQTK
5kLj/xmtmCtiGeevWKKHYkNudhL1AUUxAvbzmWX9Wk2/3l0o/l7KODKCUmS2XaoT
qM5wh6H+o/cHxkh6kfvrKT0TgbueVza7ErGGq+XKouYIkqvWHHByqWUBag1Rx7Hf
SUmqPYqMBvZckK/WJfak1gd/Ba0wvPLyA5TdYu00Q6gy9wlAaPcRpdx1Ce8vNiXK
ahBjTRo4mBnee6YK/W9eNFHD/qbCQMfcux+DCGOOXPZ3KXL7dVBvthX4z3WRz/KL
8gPB46Z2q9lb3pTNhP1Z0ldh3EUvyuLIqWA+BdthqjL5BX1cTRdsQrfoEa+hpaVK
z+iUNuaGAxKRhEyPNLKcqi5Sbbx5tdDiMaxE19XfnqKQGhtDvNAmErRNYFFWreLU
wdJwzh2VQAPpFIKBux4MUxjzGtZR3mbbbwmnsLd8ZB+ja0ZtnAVTncs434jo6euY
gbysS74UHgop1vq0XcOigviAQwY5n2LxZz4FpOK2RTRfS0VwoWeewllX0dtm1wfm
kZXpz9pRIpwX+6ze2FJXLmlRQYTwZUlDuE+qUOo7y2kAM3MMM/GX/kltMknNMKQO
SpNjesu3VuemKA0N9l/g65Cpk0r53OkkDoLCZteMftoXEmkiUr0JLek+U3ZKeOqK
u6jcWqhwPBmRE1B/Vd74ANcYimx/LCWMDPJdHIPhJh4i4LWPiNFhhrniYTLioQ5+
8t9tPnGXeiJSCC4kpv6f4dRbBdShd0ZMziDKS9WrEvT5ikT0XHcPVgaNM9ysJS9V
YzLGpTsdNx4+rUc/ZONAtmgJ+v/cz7Dzk2h05gSFjwHgAYKXQZoJS+t9YKOzBeVv
Rz35uu7OZLKVw9B0lAPx1hbaKOWLijQwcQ/xoLdoRgPe10dDui+p0Wd4sGg5mdhk
0xDFI/0Prmz+c9QzhrVf0IBjZxvA8HdYcJamXCZoQyVARUtcVVjSpk63MrQeZUG+
80B0CMo9X9SOMxeEWsuZ5M/rAlzg+MeojibHVp0FM9Smdp0YluzlSL8k7nw5Ccsm
GyX+ZrpIm28b3puh8CI4Le8wYfWSTe28+efKI3jXK/wWdWyRMIPR8bt0D+64rfVW
bPKYhpHbuyk5SoCyb5OZsa8h1PN4BYMzIPHBzFfjFlEy9Jxw/UxS/djRIKrbPoM0
g526KXMf+NUqfsqruwmXpbqb9f0n8aKat/6F1U6s98pUN0/z71h43tLeCxrWOUv9
RDhgNVecsUonqJliTn9TsurSnrBzCXmI4FOmvs3tmmsAfzGsBpwbPC8HKTTUphHW
CdcAFeBY1v5OAHCIVDkiqHKq6V1PZ+rnW6ljkQo1uunvgYI86qu+Yiq2DOk4t38h
ttsHnilCO4jQPUPIzwM53EOb9tRuIstig6rsHzqsTPEdHz0TrJZEBhgV08yHuTdB
YyhHYACqW6DxVBAyiInntdPQrKKCQro3hcTCU8wTY9gKWI4+yYxJKtkuMuRT3Olk
c7wbtRr5c949IPnH+RFXEdXg+vYEGYV57dI4HoXNgV2Y9E1MzKdNqThAWa2ixpMV
Pn82nXH3l6EaBTQHYbiicn+epfEe0ARejPMSsZHAKwRhV7GQifyM4HBMXcVnlvIQ
lEDoQSN5lpRp/XPI5B34dhT/9mOFkXLZy6QJ5RRg43zr6UlX/45irPVqMs8WfSex
Bfq1weGExUwssKsNCX5gXVxZuOZvFZFGPf40K2g4t3xe3iVZF7X0SLiMoAF+jDgE
QBs67Lk6pROLffV7rYgzEfa2ASc8LUtTvNxosVfoaxqATXaEYKNITz91V4oWmPin
vPOhbQ8NiR7O+0KmgSiPCDBzZDLPHxo3ZH/81qC6RuviqEOi+W2SgSWQ5EGsD8/Q
lfpWWIRHU5462CDG4sqG2bEX527EFoJrkTDahzw+oBbdqqqZejeurPGafA9wOPlB
Ul/ffWtUP7cF2Le5l2Sfng5pE4/usj38UMuBKNQj02taGYYr+00W64V9g2hPki71
+SUeThtI6Wc5EkHWt3MJnEBjnAwdEaYw4HneAc6iP4ze0z9knADp4U4y+eoLPPEC
rEjoDJ8/bmByDocxulXKJ733lfDcFHDtQCk+RTiyqfL09aL+thaWD4dlPRuNpETW
pfv9tbfJNm6uD0MEg7sBYsMZbn+yJ1zgOd7winZQL1Y9RHSRdZTh9Wa5hCcYs0WR
dDGSsDVyptnnHz9oT7a4DHXTX3fCYCg7F/2y0Mk7W6ufzVhPA63NVZACNKxFMUhA
fXg06OjxmGpYe1cYuHcepgj0v6KkU3mcGngW08c4zIYDnE6Z6EEgKuJ58Sg1bPar
coBihHoduqULIs1rGNZByWm/JPI36Md3IpV+QXnXAFGqRF7VFNU5lQtyTD7FOmEf
sxsax3LCgsR1iSNzsuEwxAYxpDgbeDLJZJ734YWP4xVKica1EBKve/3iV70kp1Na
dQkYIHBQXjenuK0f4sqitk6YvlOPq3wni2PDF2VsV+G+q5e9qbcc9rvAHvwsPnGm
vyLgJg+/iPbXg3IsBcha5fXziFPZTifszi231WLqPNTtxfoHUqqtI/LwGXUKmUSm
GU4A6uR9e1izWwe8dvfTSUrxt0AcEetJd4m1voBitmJJ+o3Hykhk8hRwLQ5ekXXX
z1XVHb+Me79/btFd4g7YfQ0yK+4qbov/VNtzPHnMZhaMZAi16vR4RBlbMJgAWLUu
1otpsIZ5UUo0DMQO9xFh8lExKgEd3XDY0J5488hQ2BLsrqLdWP7DQ3Ot5NmFLZaq
Ng3g2NW5bRz59aIZYyoTaYyfGzzw2mQcPNGUOIuqloPSMVXWAflllB1Zlc0ZVRWq
jVFOCvLNg4hy8Csxn/NMQbZ4IqRFBj9FlhdPQUuWlj4FinS+5ix6HNCiZljqOGJ/
k3KVYe86RrbJKCTIfiGLJsnqHkNz7qj3qo/n6AGVeio/btCHkLFanHIyjm1t7oc3
xdNTjW57jKoM8UHu1sz9uICDsvgvabiZTVUt/UaP6FWq9qf21Un6KyB7rXhFi2UX
trnsGlUV5fSl+9IOr6FxhYGeraAakvWe2Et0ArZDJmC3tZWptcBBKjY813JNa4YK
QCQbiv2ezeRSm5aJjW1uMC6mAkekJQW4dXwsq5QpvkrA1spx7eHuy7JK9E1Of9U6
L10q4vEB04qp28q7F4WNbvnojUlkMUoARJ62y17RxCEC43NFJHRyrMkR1eb9K4K9
7uGkEWwJmMYgXN/B7bW+sz59L3Th5lqlnymQHqVSxqD34x+SRjEVYpSz0VabzVYF
03apee5xPvRWHNpQJVXapSweH2XI8YmHNTtbCIDqsPF1z0mUJBb3DQ0D50CWd5jH
ZbNzviZ6Rz/E1PUAcr/IELV7B3uJCukpVwcH2Qo5o85SBSRXgfMa4lXiBnoKbOI+
pPLX2bSzMplNnjUcAk8OWsGO8cMJvJiD9uPGHDgdBx9DXU2ZgO+nDzKPrvk57GZB
k+Qc6XKxJHKqeQPE8DxRJn7z0FZYb3BZ4ovcS4w6EtT9IV9/rMSsnGRZqCbDlYpF
nQ4jR8CMCcqVKuI+7la7n6zsHE+nGzzM4OcxsaZ7TB1SAfk51fjp7vfbDUQbBD7n
RR2VznoBOU1YwQc1q9TfZUeOu+c/drQOqATIvCndMMeHYnCBtqBmojUKUA6bcggF
7HLRzwgby4b/CI9iTF7P8Hf/5pwuclv8v6LYE62mC2mO6bPaA9g3dZ79oamftK5v
3aP7ChphuLeeyR4wz7nY/97jHuSTJb14SA6F+WscDtLy4NiErnzpHPKsHPYkbHj8
jk2QaUqCTZ6BlxmnmamQR/lvZRJF1WSxNrFw89+uhMeh/5VmrE51OiQzW+nqyWcC
3FewIZg2kyC4pbjsA9c7jib8n1/uCLAqvrZMLZOOp0b/pIWUgI4TThbRYcU5pwld
Df/nO00JKOqNazZEKJjWIXNyqdbu+LRv7dY9uJCDL9HFQGKJSXyISbYuOWKZg6FH
EJ1VCKluA3Hc0yrFYsn8x3bnxy0ByLuzpl5TLcoWSQ6PEhSJUMN9IUMABKp9dChX
XF1TsHM+6UX4JPERMQ5eP0kx5YAar6+OhrJ+TdI0QLqpU3Y4wnpv9FnoAhPcdWWI
P3xVQDgL+gg15xv6uNqINEHTXQyGBZtbycy2Phg/aURjOV5Sy7CX6VzWE60E2EnC
qFnBRImhwRiOqy/J2Ub3AzyIxmRxDMppAJQJpkcZ9sLB7hV/q1qXDT3WasPJOu5I
1+Kdwp28Zip26NV9TfI7RsSw7jvuIEoLQ0axrVDDgT91wpZHkllJQ1aq+x/L1n6K
9yOlLcIsCMGiXasziKARtf+KeJVAzpQG2jU6CcU0BC8jU6YT8ym/VjRTGD8Mk6OV
qUOLfrk+aDHFTxb6SMaSEBecoLFoeTSbbZzHM5glPkZcGrDyG6mkp3+6Miax6c48
0MlkR1F/QU4ef91SCc8GQTJ7ocuGxKS/knZuQa+5OUs1BYKzMSIfggIwBQyBzCIQ
ZUNIuSxp8bGGLh99bwCHX4Q2yrUq0mWxY9HuO34qTZgXWoJ83maZeTCR29SbwTg+
0l+1826jobQodqonm17crkVRruHHpwMutKFksmZLm35kJ+xFgr7dNmWpvOlcrcB5
+aI9TeL+dQTnI2dtuSnZb/of0GCXkdJwtXT3kiPb9tCc7FVA1LaQ5qI35b3ihLxj
Xve1YjqQCE0HREZCUCCY/dYh1JvtWubwduj+AAvw61sH6Ygs7aS66svglriXXWEG
HxGYiC09NYn3K4oNF0KmUL3cMtihqyBt1IN6fA6YlM0759y4/olo6vA53604sCtF
qkpOwxLSSOOMLfZahPrkvq5vYco7Is3umIxFJlpLqsOhBa71Xe4wsreAAIHxCkcm
2t3kfgrSCGjsX1jqIFKAjDmWgR7l9FtXzYdVWeBupRHyO5L7cyqdI13xdZyI9Y8T
yJg+GFthJdDVm6G86oW39fvXQfd0Y3KNbgDDunJgg4ORQp4qr+NFsI2FXm4m8ViQ
F9OuSZhIVtFzqHvWbYGg17pzhmnIpu3kVAd6fwWou4vhk/N7j7XPKByncQfM84x+
3YRxC6Q12Q/u8saWWCbfYNGGUeROc8rEQpQnfkZw0CM6ocoedgoqFRpplHJ7ROex
K6DqPVuL0w4iu4LrsiqD3iMAlJAEmXBZT4aqEEz1EezafiQ1ZP9F2XmCH1qCon6Q
AZxLZV3o+5SB2z1Db+E2ySFQNGtYqq6JU6cUzAtpSG0MgH4mXwAPH2JFnOVHPbwE
z11rrX5yje3LquH/a8N6zH+TmFaNfNvTwlhmLzWXCOGTiAmJ0WZ+Hlw9ax5hLgLT
4lbwObbiguKcaPxwKy82+VLchzmfMTqO9Td3YLgig7dFNfwd9S3ne/9rNgDf7X4e
/e96E8WHJ2RPQUx/+GYZhnncKF9sYmz9eFp6PuqnBRHoJGX+F1JXRsSmCDlAQXTm
KnQwbrSyWYOxDU9tK7HkUjRWYUo5Wv+QVEn0RC8lQUjsQqHxFB1zAEYBCin7LBRF
H8kptDv5X2SN8cMJsB1+2/ctW2DblQUqDIDU/G2XWD3NDvrfKt7q34i6TH/Xb1s5
R7trl0Jupa33mpG6sDRLAAMI9JMoqE/BuLaX6IrtE//qBzTd8x+RKigbCIv+iQjH
uBWJzkZrcgT1J+KBP6d9kc33rI0aEHSyoyZvj94YE4Wt4kCOJdFTXJkanBYhYiJl
0IriWZoAnpmXSA8r5fgoAXcGsrydTU/hR42bwNlJwbkk/QIw8/a9a6VLpVVDgg6a
ySFa8XCQJMpnXQcEUMKGKitpazlDwcr00PDS5//A93n5GuFBh+L4IE0kijQvY0Ro
J4k09v9z3QliEJ5Oga0mi+xdK+ESCZkL0lBVwf4bDikymJCFjnnrWFXXAbX3N5QY
0T/M4Ft+G/yiSmq+9Tc5WZHq0xUs09RmNiTl5dmWctQjyXnzSHfSNuihnPNz2eoH
Spow/cK5XBkzXmxKEmS888nUEa8LL5Ni1fdDKxL7vYxFQuKEWzKawJJBf6yK/Wuv
7OkBdxz3Bw9qnqb5/55hJDIIR/4TeTPkOm9kZWAFzIzf5sdo50MSbUYgQ1AdqOfn
mYpClzkLZ9pBCwYioNLx7SWFDkRjyB737CHdR2kSwtHQzKmZE1RgbxZCMIyIk6hu
MLdeO30DiZny9sUy77KaORGat4owDir0f2L967I+OtYWFFl7ckt/3eSsz3yu49bA
4i4S1i2Mhj9Xe5Vd0fdl0uksg/ed9bhgkKofCw7maMOJyoDONU6Fhz3mXEwR2J1t
CjyeAqCy6ck8NKkwmNxRlAX+EGgOQqMJlN6ukK7uCV5afqpxtuG9lu8zGmZlGqdy
Ntj6NU77BrHvJdl4Nu4fr/Q0DoeTdvVXbB7qFK8NuVuMSvwtAYrkghEFSOmk+W9p
fJDZmHJYKzjccN9OiLAvvUBEby/XCYoCKy/wS41LeYn7NGFay8UMm6h88r8AHQal
jBuMAbNdVk/qDzqsaXvIw8IfY/zTfb7biM+CWzm/BK6oTHC6eoQslkRubaMGXF6q
gkd53eACLLJ/mOP8sPV+evY+EtsG8dD+zM9y1gSsvuOB/ZW1AMQsO5wLJehz52iU
Ny5/s4T4mwQnpV8S0BITpQyBcKifxZyz1/N8dxAA3WTRpeZDv4tPzEi5JiogsTxG
SpIR+c36zanc5uEhhywgyH41TJX4xkGXuDzeCF4G6ziLnxiT9XhKQ9g54QFjZdak
q4dpB/b+c1SRNXoVisD8Ai3kQI1h+MI6Ul+PrWSESlW8DN0OaQndhBai6q7n8Mm9
2BRuvmNkySTgcK+TWb6XiFmHE4gIxKz1rGU6q8lsps38ksfeJG4b3MCjvfXe4s50
hrIJAwWqZMnWpTIZi0YSKOZ+AVYDRy+jh2Nv0wReG/Y4FCk/cpZ7rWwDBIL2f6Qr
3DrqfRT694uVULVG2lDYck6v77+wc8Uc3UFnm4dKWS/V1hSCg3F7NKzOFgKSVLpj
Z9JzvlFEhY2crZ2d4KTKaSCx2uIaTsOuFpNXHXiHZBQfQDK+CAOYdnCLbiAAowa6
0YL6bY21eDus3g71RaTZTJUrVJrLQ3Wa75enE9uEP+W1cE3ki342HFkkwAJE7rVT
H8bj7766XDcY2804SH2LQ8BTaj+0GLiTaGYE9lsNXOGoGvZZp62pdkJiDfmr78ov
jRc/683MWU/eSgRZX06qasLv2bdY61xGLhWietAwNh8z+eE4leS66WTfP61plOgI
n+nfbGwKP8xOJJ4qYxbv/TqLGf6S0NXuIxuZYPk6MDEjxXFkxhMrhtlahS68cVTu
NSK2qQV/79woUAGx+l0S+Nsw9lR2v8i+KgQgwSzTaaE6Tfun3HuMP/t4JpU0zq2c
QbjP9kDLpcyhDGUXLHxvQjR9F+T5sVJlcvMkRuB3PEL0Uva7o2Akmi8jVtO6V4JJ
XcF73L8LXcKGRhsVHxpVHqqTRSQBm7INbS1eZWE3WXsFVdJ+1rxpvvZdFAdPjHXs
zv65sv+z2nzi4qTqu9VXZBx7H2g/xzBQJuSIig6jL50SOxiP2Bmk/CAyxrYud9+g
qIMDIZIrD1ywDyPuWITtASSs6FekOFg2iFmGa42m5jyJZfH6ayKCuC/GBnlrResu
zHvItDIdwCiK6ichHbPaAdtIRiWVcgXnucDsYQDWRcYxPDoerDGF2VM/eaToSBdN
FzfkS3mThpXnhiFm+9cjwSARAjDYl+ML/IKMGUYprDovIuUs7qdN7Cn1fG9lxxbY
kioY2g0bz1qlEi+1VSfp+RNudWDtPSThVGdwxQOrK8C85GVS4KX2OcJlCQmkDNFX
VKf30C0aDDw9lD8vBTnSkKY+iPmJ1rUqMXJ8r6PqMo36jKZ3us7wqfuIFrfEwSv+
azr25ZJAIEBOHODLWgnXpwm9lPE1DIppoI+dAXLTLdVuuG3UicqX7yI54ZUeDJz1
GvHhA6rq4odJVEGwCVRjurKIYvOr8oz/kwHvtRPgiYZjZ6xE8ldnvYjWA/7RelT8
CyD+hbZIbKgbcTBs5EGO6HQ6o2Ta8EGr3TT8+sFJOR/YXQupXQEZamFubTusgCnV
uXjn8I9e37ugkNlLpqt4OUypqc5KkjiRT5AOMQJUfMFDE4rui0MCT5xiMngFQc7F
FC4LZjnw03ccnoSEJxh/jl4UIu6mAWN8tmQYJ5z1awnZ1vFJwCzTRQ39DdLPAR5T
C1xgbFKzcEdRwzvKX/tGRHRrORFg0xmcfoMSdZaHDgpBXod7RY0SJf6fz6AwZKnJ
eR0vwI0kMXxKsOuhZT1+uWlqsrqzgLpSfG1V/UlurljWh0o19xi+l2XuDQ5isTEZ
KB4ZBTe3Sl0yVB3ZbHr/ocRRDDAbCXwxIhWFvvd2D6KgagSBnGrZEwz1mjqoNFq+
V8Ah/Cy7HvmWjw6/1CkemxOH8x+ZVH5i0Kg/J4rR1sST0YRtj1PTqeLqtTflgfaE
9gP9m/FkeK6nF0ZEMDGdHFZlnQf0BcRx3hmEtMCVmL5IHJTA+temTlETr7lyxr6F
+rmr4bNJ2ada83MBtg3vhCn8X3fW0uCYxsrAmKq6DlrlK8XnUIX8hXDro2nVwpj8
H6p5ULV2pIJJnlihpHOHRXosW0B34B6f4WsSe4m31cCgevgGFNryuaEN3gl5b+Uu
ZRnYQQYKIQRMOojWKU2QShPxBsMaAWoBhlaJyjzknQyjGyWTi02uJFvvS5Dv8KYM
wuhP8pLsIdnMpztggOlWZirtnqDKHGY8SRrTozaKO/AOmmJWQdMN7WOWamelm3nI
PrM9UZ9jRB70Aa2o0QjfDpm0U4ZNx0KH7WWb1R4ozWHnslxFTsEU8om68ukwFSYK
f28NvAz1xAfLLELXisXMR+27WxlqIXSzWqmViBW8gBj6DkloQu2fB5e7Y1fE8GF2
j7OlKZsOojW4QlzykbTMGkM8OI8sTw4WJpjd1MzhSUzqDJH2LV++PMzPiGqM3QQO
dhF4UXyKeO0vkkOoGaoKO1uqavz2hCgYauRc991OWDBbU3sKYy2fisdB8sg0+sXw
x52sGti2Kv5670sTkAP8GyWnuyhO+zjIaBeMWe6g9R1s+fUpXtQR/R6PDtYL2XaK
Q9SDGznK9+pA9N/6VPHFdE3/c/VdY1YxIE35I5KqSMFJRQFHK9dFrqNLQAkLU8RB
ILrKl1P1JyNlGg+8OdrhNVR/5arZ9qAkym4/IpM9mZf+UQ3sRPBfkH1hibQybS+D
CNhzpP++ouJn9xd10Z/jsAVc5DLNAVTlNYHqF6PAjXaYjiOlTTKDEWa3cPGm/16n
2D17gr8DDmqOtsu1LVs/VVkRm1vKdm44yflAeHkz1sqe3amfm7kgrA3GTU4U2aAL
/6JoytDwnJ4gxQXDllAVjSTHWNhplo63RG5lXoOJhPn0waaDuLpti8FGCtrV3C8U
9ts3YWkV6jSI6sQZaHFZFJi6HJ/9l0IkuGhTIvQEuJvZSA41FDWlddfCBGW4BlTq
2+TCa78fAeRJA5EtlpUHN34Gigf3ytSkjJE+mAzYQZwchCpEM/n5h/S3AzZGtjwu
Z/o5Zd+jwZ0/w+oxHByEaZRWbZ5YT1ZsgTHXsO3KTMwdqWwqs93ijKAW1hFGUinw
itbGWu3NPKUH3WnI5kle5ZgeEFnUPr8lpoEHutL4RBR+UDYGhyZKdza+DNDcTypV
+tN53KY4GPG1c+JcQO2zVZgUkaOgbLkuR8oqc9MtJQUq2O4rjsZpYawEpGjL7pUq
D+NDquQt8ZCDPAgzuoxEF9uTHSfRtbJgBe4+2wgbeABMaZH7Ld+YML/0tyHBuWXB
7CXTJ4NIoreqdiX25sKq0qyo10nvWxd3OXTIusOrv40jPnpN3e4BD4Q0hOGroa8/
Xxo3SCyg5Vz6qoO729ndGPbZXDJddnCnpyhYmCarsAVf0JEOiXInw7Olf36f3LrA
efou56TXou82wbE8z880ueQ2J/ITQv/Y3p55tBOSUzkkDP5nADy9p/7X3D6XvSLI
ltj7HuI3sDC0keHN5aWx9EwShJ2No2USKn5Z6PL4vrJd1EHSvWSlct6nWVF3Lku5
h7pP8pVVRlQmVlajoqEvlTQUVkpTTvKOrHXf2Co/OESDDByRg7NCsAG9B3d+SM74
eDgLQ1Ju50v0S+FcYnEGqxrHxMDwoeEITrmetuzFFsdvW/XcLFUynr2dNvKSbxtE
nDhces0oP2pPivJ6GlxZ/rHdUej9SwU1Mq78w1TVetez4+MT4O60P5WAMF//kRRG
npCtvRecKUptw5u7Ur/UMtFkVxOvBmOInms5vtCnZWZpOavkk8iKjOIZfoFEfi+k
r5CWRRFbC8s8y/DlzN+NMvsNqPTo+9dRTR0dfXqY1szM+VHdsHiroOYNMNBDItWh
c6Y75JBRmPjE4dwHaegPE6Cc5V7+dRUkkT2ev3VO0OJbm1TnPwJXgCLcIgKr4R9n
qMSqQwlUtG1TGj3Ki9UTfzsGqRG+rnPL5nVsXL0T3biJVNwMVv7S5LS19l+DeYqP
uHFKV72JAOs3kPjx69+hbcesZliZeuI8/76NdlctLc0VQf80J1nnP2K4VYcPR6y3
JLkJcAiexlg1orSL1jFMf+C/Q05NX22IzDNq9jRbnxaJKiIAFWSEwwKlvu2yKjP/
k6LQ7LHbiO3AGUlbm0vmP/Gs7V76n/8WyNRXj0fl39phcaFE81Z9MO6P6wcvT7kk
5Lfh8JEDasMa3LmgQDNRd61el5tNWzR9dmkrRCMrS40cmOt+ef2bq5eebcGO1z2P
o/y4mIEARnu1jf7ZO+cs2C3lDnpGEcMqGeyCt7hWTrNX6XV8k4LTZKq44+tuaiHD
6gODOZiR+d7hJNK/GTXcKNc54tqeA+GJRyhF6ra54TjNQufwI6SUx3QfPKSqmDH4
baGb8Pks3o3SmTUS65Shd/E4s47eFqEBxozHmvlSDHqixO9u7V4bJsz+MvM7F5Y5
CKeuaZXfyyAikgXnjJUTBpTEwPSKXmjy5Cv6nKLL2b4bHH+Wh9gqgNtQkTR2G3+4
VfF/gD1R5UrKTdi063Jj+MjBaK0sfiI3zKbC7g98qEg79La953GUKkXCDP+Nlh3b
97KpeNuZGILxNwaRNzaavnh7LRPRpSuVKr/ac8/Fe5TG3msGaOUYtPkM7rOsONE3
JvFWpLrG24sfmBTcaN6qQuiCAQifG6zV1Ui9f4RNTKaGYMpd+5VxlnvIjq9Pa2Pw
eCTGAL/k9VhggrUze+CdncI8TWQ+88F76Gx/Ws0W/ohdjcTDbYXnXtHyIK6esHKb
jr/JCQ34LFsfmYkap8rC2YUCvgEj395ZfxZjpO0NiO9nEeC6JnTceEYdmkJjc2y3
EHER97n3tej/OeR20qkC+4rxTGDWCKPeTgPNZufiXZMm7UJ2e5dacStU7lGRLGVG
P371Y+e4xR3W8vDhHrF2Yr9mLoVsC+8IYITyzHgmro73W5kwk5ABnzS1JpS1WUx0
VtgirCjVEmnR80OaLZ2thAW/FHgyDNuBIAGixMHcREwH3FHqtwSyjwl9zyo2aXSn
YzwTv3XkCLZznWFb3N/O9lOkpfdyE1DFQKNVB5Io8QkVkgbNqePhIIxMfxxRlVxg
tq3Fk9jakQRTAtAkQEZpKD1WdRnZUpcIoxSp5bayytcfVO/rrxO3EfwhV7bKkwkB
GnU45ixU1+11cb3MLUW66xM87Ro9QKImdTzYmonWRUP9DmbV0gZxKUHPfaQvaBI1
qgpTzztC3eg+yKH3hA6Oz2VjWGKQeU99rMiVnmaX94i4FmVhyMEZd+LUXFVpgN8J
A/HGlpPZD1ezYaOPaHmuJMzioCXjWkNjZy0EX4cWGQFMBSKBPYLalBFJ9WEEhujd
AuiV8wxtFnudci07KPrziapJUi0oNulgSBZXrTYE3Wq6oavjrow7j1mAkEspCDJ/
w64rPan65y/GNdtNi7p+rc8boPbAHdd1BDuP/KwYi6iJPHuT2DAH1h8JmytyvNSk
oAlCb/yKfpPMu30elb9zvk+PVf+BmeCHUeHdmukUjB1suKWGD8euwul4QEL/CKkB
ndlYgNdZ+bhKS6A2OwCjivnbxDZSXaVIeow0tIBDX9/OgyQuJfs8opVkVAje+JhM
pfvmidIbT97wmKbjrEvzZTWcIerFweYWP2y5aBil8I+r3KTEYd56wfuX6OKutKwE
0ASy8SoUbP5KiIExQ1D3CPgGOZmbCwo+O0oBryIctwRrZdGhwlk9TizRjbQdiCoS
IENyQdHol1rTyRydaJidBWGN6Jjjw6pZui3bJlEsT5TNVZ4IC8QK6thp7Fs0gg9W
RvNKzJtVAggNfTLW+crUlOTvbviTMhOLuHqsrljrUVnRf1StZtgBQWnZRtrZ2t6y
SfV/Yq6f7yU9arrDUQzB+zFrnajemdlSjfi9RU96Guq56YL18bIWbg3/n3HMN3gf
whZT0AvyiDOCyjf4057nwbzJQe34dvPqGUOBEa5ZIMmL9EPJZejl/2gDt+ChPSGW
/NPr26GKjgoqit3nyqVg600G5sYIAG1uiMV1MsaYqvtxVI/eQn38jvCGL9vUfuFj
0TA3S1Nu8R2SxGGQ0CEPkNIzDlpRDF27ndVJzCAAm4qDaV4jqhcQi8+2ueXux+Ms
nfGDCFhAepUOF35xpGuEgeNsYbOhPaKAyWGOTusNopwmmx/dmpSx5Sb4jBvQZABz
w6gvlDiHrZAFUzYa/tzmQdslyax8zFbCdeCrZDPcV98yOGqTgZ1KROYyRlBP4z/B
Iel2hTuQ0YNvKjDEAChJbVrW7t8WsLI9tb5/cwvxZftjqJrxbbleMhRYvltW5qdk
5OkT+elXnJDZ+GKNHuAOi7dIABzyg10wGPk766VoKGNiiTrhFn6qi1pbJDDtm2zJ
HjbWBt98oPQYOANnURqL31pnkDGHMJ+fIMBM5g8GfD0QBOdhUkVBsNppg6irfupZ
5wYU5LvRd0ArWqyaM3EuArOHORArxZhanDmU4qSRo7fCxMqoWJyvqEjbbI/Ctc/I
8npQp5q9sedARxQ4ltg4tyFGaikBen6D80pvbRz4nNl/0ZQflQ6ONUS32Zjh14di
6gLZrbS/C2ZrrwYwe3gKerIoOYR4xirI8KLkJJIWbpbkHYtKDPb4aMrgioXqBWQC
+f01LylPZnOvXONP2A8oN0vStMcTgfeTg3HFcF4/svSN4HU86PqHJ6srid+yWtcX
StMSK9ConI02ESn36DDMIcsmZjc6DxQVGjpzQwo3KhIk1mezxAcBxdcVSKakNDb2
BW+dOejXLp4lf8ZOj+Gc2fp9I10GKH/+wi6u5wBZJE+Fd6A8OLy+kzfr7ne8vubd
o1pQeyJoAnYBB2Hnd/VraiOWH2rH/HQn/Tw4idMhV6WPqWNUUeNq1YbVPntQU8w9
yx1Z46YJrMd0Jga+M5NTkrSIJSPNNVJzv25dWfLpKfT3GeTOjTcrikSQxt7tE1fG
zi+/9o4srPJZIYwfsisE9WpAyonWoyFGC+izdKzX7xFlHhbCaIyJcW3eRjiAind2
2S+CFs1UPvRegppoeE7dP7bwXz7a34uOWFn8QnwApJjecOz/PqhFr950gxI8OX8X
zEyfbud7jw7ipxa7nkO92p61xA5LlgOsQW4RtYQO3FHmzExLOVoAlmO0IiZeKQqm
C1FKMQnap7AMYx0IWjPKbpbP7gAwyUhF9eunk2kTknOmvW2xFJG8/ia18PJV5Ya6
zchOMn/KYPKb/Jv5yupodZr3lyMMRkeobbumYiBQnjwPQ9kZfYmX+Qi4epETtFw3
7WTYxeTCmCGFr6E3fPtEkQzPrHYRz9iCTA0bDGxrI4Lq+b9HodFO/2gJ78szyUl6
nFeu7SqJtc2IMhog8NvGcE5Wunjq8oJWGkTTeBPGcPwwzbdoIb6YX+/upNJ23CDo
KK2Xd20Ax39YGPD1rsqlxL3JHBUr68nudI2y3Q6fwa4WCaFABxHCpBXiP/6ZsekR
bifeVK1dwbPLajyMYEakDbJwjPRsPEo4gXrrwm3UF0s3rTa5Sel7Aiyx+CM6tWI8
jpsHJAjpfJ3zKzQsT0GxQxbGtXfODyXKU9/Bp5NE67X/4GGzVGVNInIYIbbQau3+
7HEpxo/i94ubdjThFTJ/cIVZ0a60MvvXod6VUPvB8pbqhE50VFvaKE4KHFGWS038
7/E4AASdhk5aMMgmiLRrIihlVbBbJj5WRfKq9IeEbyyiLVTS1HTypPW+sFbzunZs
jD1lMRRDBbvI+Bs7HZ8ZpU/XCJnMaDpkJkEPprtKqP2Go7HURuj7ZZjcdLQ4J7FU
5o/7ykfenjd9dE0zS9NakvS+ZKHgjTqULnpiyMgtXkXl2mgYeVamlTouq+9yp76J
6G0Lpt/eRR6A/emckF1c18+d1f4KrPikvFtRY5GLSgtImj4EpGq+KPmXfajHmD11
4auvHMLeLL77+VysxvaWaY1YLMsdQNhoyrsAezG/tLxAXOJAE3tNFsMv6fMdpAOz
Wtfg3r4LWaiT+wi9X9NYK0cQ/OUsMSWTN1+AO9ByTWHyeCDgEGECUxtMEP6vMh0g
0HEmtkkTin6//t9/L2TqzVFyOwcC+afktaMPSueiKMWjpNHmmR36X6E+TVFcE00Z
LSdbG5+x7q15isOaD2ki48sPuz6zOaJZsA7+netdU8YKJmeNAg3tVER3rQ1IBngc
QRDP/CSq1aN7WWBqZs+iNaz2L6TR+aF/1gEykNLzp+v3YzZ7/97HNhNzo/1XFm5G
jEzJTw3ru7ySdDv5eiJh7SrPx5OmYZKEtfqmxuFmoKvWi0R90n5O1zrdV04PTFxc
dH9xVCl044WG1xoOTEjOnH+BSx8g83zXplgesAG+UN19xvg4L0oHJz9wD8RGYLp6
KVNWMVfiAYYku7olGqFqa2gt/7KO0In6n+Hp+HowlLRNqPPRi7lLCU9PC0gixCp5
GiA+08K5FyP6WQR8joquNvwFWLuV1rql+A642RgRV0j7psZboWc9L5rwk1tFPxnN
/Kv2EXaEbqF1t2BZw1ZJsWIB36prfrIO/CUDy0/7426RmEoZwD7y38BT0NNCBIxZ
pNMcuIbtUxajNpdt5aGdXT1yBRIYAaX2OSsy5Y8FR1WOlMysoOSaN3vgiWcL2zLu
zFYnx/RyYOYpF3cShEds7Qb5o4VVxNs1lQ41K3ifqpNOJs1hqCaCEwP+TZMrNlJ7
N3LUQZ7mqE0O2qIL5cTGft3sxeRrqTL1nH47gXr0WF/hfCkUROSl2qa0dRnfuGcc
hoBOhf20H2arzYbuAWEZhCBZ6H6i0ns007MrTUhOcCPYtrGHw+TsRi/Gv76onj79
BGLVmESX/ixNAU5Q5xYlUXWXxOOB3ldBQD00lOjpFJLTACXzrh1MJLxe/6C8lyw1
CppUbrG/5Mzrjjlube0b+ROg2bhxQcuxw7DyabfW5FLowiOUKjWOBqMfTmJCye28
W5he+oLou1Wv+fOqbdx1VvlEQwrRbMaxiz6uPiHgpVaZxtolmWBB9e3dCbUialk0
Zjduhypubn2zXFRO4y1Akv2gizo2svFls5PHbeE8HMu4HfTVAz+tR02G1Qxk+L/0
lDvtl1LnPJ7/5CcZ0uVvlkRCPiFnvoHt/JzIGebAdKdaAFWaCUb0yiLqOKqe/y/J
w4Mct+o4emcYl45cX5chw8ja/OSUk5dhd/Uh30yRBkpGNwfUsNqzToKIGr1qJEgx
Kfd9tlAsydZVbsZM6d1DXd1lHY0te6lfi2oGPO9m+ael7dQiPBxlHq6572OFnAbZ
YQbrQ5cj9elF3UElqx0ZcSNegCFAIFMNDmLpYdVY3Lh5U9dpqJGtAZjoTQonawR3
xtguqIvyyO5cUv4S0a8hM2inpQ4GpUQoDBPZJ+v7bDmoAbbBvEBAwOGJh+Gg3THh
71gXcm/pX+KMB9ikC4j+qgvvW/80lXnvYCLGkdnElH9Ru1PDPIIoEf1LE4kHIV3w
zQVkqZHurdkjF2AtnJzB16svEOBgnw1wxvRJVtPCmK8/qOqbPimczQrpAq9KMAfL
VzwZmvpfPCSXkGX7g1nuUXkiVTZAEjQkEaFGAvu/v5OXnYXqz1kc0Dw8z5H8SUHl
DEmZeibqmAk1oF9ijtpwAaPRW8EY6qHplz1VcP3s1IoxCDOKv0Ui68M3YiqRe+do
Fc5vUucoCXzqHqxbV5JOi/BN9A0Sc5OutbXAUakK8N/Kxm88LujWpA9UvATVeIFQ
9fl8xJLNqoqdRYtCOI9AD31r7pNY7N6PlE4UZwF2sOZmvTQViVn3pb6STMhDLFUX
3Z8BkYQX1j4ycTkpRN+rxwIrAtBOUEgFM65PVtBRpldr2WHNzk3BflZ2uKS70SmA
RC6UvbTfprrfgI2ys2gjb1GLwuzOC3OT+6zEBTcXaaaZypgeGYTHyrwcg+tbKEai
t5C7RS2Hnb+jlgQjtdlv5XtsJzDFciIvsDbI77MFRXs9yjFdSW82mwXSX835j7N4
1cxu36FpnpcLkwPAgxM2maoFm/9BjcSKdoVlSqmfhZD7gLxLH4Ea8fwdc15hNZ0O
QIfHg1fF9L0dLEwQCsJCB5uxp1H7PcPj4nT5lbKoKs0/gLPtVUxqH8B1U5Tt+4hA
TneDvXTwyZSUeMiQNsz9xffSkZoyCw0sDT0G4HXkV9Y2eDeNJy9sRQ1r89HTEkNL
cwN3zyyaQ6riw4F9wQi0w5260Ff8GejbLfWRI4rMeScdIaRoduWMwlHfsdRrX5Ku
3T8jQei0IVHllxmixmoLLRzwoDMyCmjcxteLSFj4gQE0vT9QiILng8sgFBtEB5F2
OkR4W9gxTeajxZCM9D+DhYx734uO0RYDJ/0pAwFnLyZR4aLut+753yPj2/uP6VVN
oIUHne7udq8t1NrqSV7pKQMO/drx88nau8NxFuwF41auOexegS4El5YpUP9H0X9O
SJjI1nhw8nX/AbfBkFATAqOkB5ET76KQqnv8fYsGI6clO09QSvOjHaCZPPH42ynH
HqDtmtX6xcURWHwDn0ngRCa4xeXU8PDPel2mWgls20W7fZBEDvakj7i0IfAThMRv
jqzU6DqdOVeQV6lZygcSXAZpO+LsyaHODlCPeSWK1mOm0xTO60+ivK3INc3P0zOG
KuhMTxLz0/XD1TM+9ytQ60jpL7u6NHaTQDo7zQVtsaVuxR5hT2CGLFMso7tEEYSO
6O/Xthxkxbh2LeFQLgiYOtf+iJbZhoXW5Ok3GZg51SaDDdTJeU/9rRCEB/6dAyf4
SNjewVoytXU72LXjp2hv57L3p7lVg8riFp1S0OTrJRDpNEP2HtvaOihgQ4cpq5Rj
OI9pLebltxQUNxcxU5IMNcTVRJeDT9vLjCbjAned9wtIh7m7huki25dt+4ca0RtA
XUpDwknMRbnU553FSDWqfl8v+H7rhg0RFynix+PUxZ1kpIRgeaz6uRyuSsLZoJDy
X8hD1uJD5NjSNqmAsit9RnTRcNRupwyN76j+zniDu4aiM/ycqWBfR9cl+olCOAVT
+8kIr06C3tDjQNTC539P8SLywr7/q1MJiXekf/3t8wtC0txnblHaJzs2EyvskIuR
iaLHg9T+yK3FPNB/LSstLUZWEnZJe66Ts6ML5tKuGmzXTM3CnhDfSQdYJ/YM9RIW
RE10/Tc4Xh2rNBOgozRgX7ZC3jfHsQefGZHZPk5A+Hm3tU1IcLPnosAypdgzaQ+g
XjAwrabq/dM+3zSMIrgqzUNn1MqeXNxC63lM3m719ukk+xMq68YXAtbTK2Y65twg
4MjeZR2aHYm1SKjwOiSEQwiyVxytjO5KKR7Lt4rePtc2QOMKL8bJ0RcGw6A9FAcS
7SZlFWh9t5C9B3oUoNWL2nEEoxwhPOCSFm6GCV56QQN6qCwQZXXS4YyxgBewqNpL
m3KBF/R7u5JIch2b8fhoboWM2h+F6/u4BZCqcL8ILIhiWn/C5WwAfFt39ueaLVYB
ujMGp0xrf7JOsx2lTdpRGqHtzvttyqqfdudTk5Q2qEbqxIj0tt9gqz4VsqGNIwsQ
yuDCC5dMAg13t3ycqFcQtuEk0G4FBfZRDE5zYbaKJ5XUm6RI55m3rRzrqyS9H5ta
SFlHt9/+WzaywDc1F5krRLCc2dYBTiuVuUkMDuvQa/38+Fo734aSNDb2sLCkixmo
wEcvrTGdxlPE4kZCbVNw+Pjfxj8IieSYoxaKA81pR92F9RbB6YCqh1gaR8VT8ihM
kw0r1UlzoJUhdtn7X/9jxkEReG1THvbFsA4e6br9lYQNv/ayQrh/ViG3IZuvAsnq
yLflR/22mpeojdRxYbj7fFvK/EUnd+voPXt8nvx9Qp6DNZ/oY8zWkWF9n4GxJ3L/
FrHHrTWvaX7pJGiq1CnGNZaJMNJZKj4DEL66PAX0QYLn+LTUNEd8fAor3IK8NlwV
PCY0ufqXYhFAM312ICvb4oWrt+kHKhSK/sZDdlB1qx4YHpN7gft6DaHSvE0m52Gp
iI2B1uxogv03dRPXF0rTxCyTwH8cQfZ0fkOSR7cZPhzJ6RYHCjVAe6atCxHYVyEh
VCJhVWkxWpOSDCpsHeoCmo3FmgQG6veHoTz5UJt9XcQjLKYLsWB6PCO7pdObN5JE
VwTJyRuKzF0MPwUZB4csLVS0nMqKC9DA8Mh+IO/YAmW08AWtU3koWrAxCLlk2vcJ
WkThcekRPnjoe2mf9RpXo2ahHEeo1QwSCQPZeCPKrxkFapGdVz+bqJJUTNQNH4Wo
szy7MpZbW5q3Melh/DjNU4T2AJZSs8CWIw9/aJZCsx8fx/JbxVUWeJPBKHHxry2V
E0qg10hcdgIhaW9OpIvXRRnXIZ3GHTL4KkuIUSYdRY/mQcZ9Qgpeu4X9WeiahB4o
u7S1KSD6CLvV9n2ghi3VPoaBqxM6Sp5zf8wedSUbVcD+Fu1Yngj1iPJmmc9foJBV
J/xtRn+6sy5loR7uVaSpVGoyyAmrWJv5qolQX/KPJSIWGt7Kp6eKafVxfOHLT7Bs
L6k7U6wQ9xyEQeM0ehmRr1RatzcJbPgKXCRWrBkS7cgNSL7LD5GBJBwqQbL8S9kN
vCOIq/IGWXQW/cfFQ9Lf0PXUZ6OdUMtkTmjVpz5j2ttc/pINDSMtdO4Uc2XFZlRS
q4LfD1MB7CyeuHWNmwikQn5rePJCzyzFGN78yEqYDzenUiAnl41RZQbLgg5kWqGu
r7F33DksczzzwfSB/YYTLGEX/KNCCtDFQgePiz/gIffjm8m1lEq2WNkA6lD6Kppc
GC+0l0qLB2XpylAiKLf+63xm1R21BORXGR8uxURmqiFeI+vMHT/6mtlagzgLIfng
uIvpdAeQTZA05FUDRSRv7zxrg6J8JmBdha9D+ucgZ+U+k/DGjOTRD7UYKYqs1e6w
FNHGXkinpfUYGoJQ3qheL3srtRWp1jSz9MB5hTkbwszETScq3kuTTrYDvlm5KmNa
GfAQNqD54+u2s27PA/BgGF7WECHkbNDsxNmCH/b+sMK4MsSm1hoZNF1G/7HRg29X
7C2KkMOT2qQi4rezVnUT+IJhMaeIsK4m9JC7+TVsqDgdNVd2oDLgfiwR9KQPYEds
AYwMo3GjK9qcLm9KCXSJdQ3iLfsLo7BpAygNb3zJdTpXSlSNXyrm59ngt1XEWITV
wOX/kDe9YBeM6SMPWIaAbrDmEljKPwsOSnAL9Umn/4O4SxRvb29spIeg2kbR4jKl
mK8P+EIo6T6I0/0v2zUhgtg0A+TLLabusxplkV+PLS2xFGlqn+OkjhDT2um+tS1Z
HHV80fUKYlbA5+1DHHouQXS22QzKzGxnhDJhJ7izsN2O9U+0GqVjttZ4m9hOM/PI
Vjnw5qbadGqVkVOGII/D/Q+X0gktO9Zr4jp7F4az8+BdaDbQxebRpU9yO5D0AOL6
rqmpne1MbIeLvWuCnyS9AnoIaD3DfiFOMuV4Me9QGfIldQZBz4sX59yXY2gdKUU/
UcXwxyh3zy/o3xsuYq6DpIzkBPltJ1oSSYFnOHV4azXPbBNr4EhlmgCJlYRZeqM/
9soK1VoHAY32Wodl6O5743Vtm9Yd751ZTz4QOP6ik3hJFxg3oVB8+a5FF6u525tZ
5IQ62yAMxZAWEeq8DEU7wbniYEICDhnnFtX9dlPKpg/vRe8O15OK61kk5zmRPtx1
VvdJdCdVqlXre+7AeZAsUUmlEoSstAECNehqzTQStddPbeqTwRTjsxFRrcQdk2QU
oZ8H9V6YxW7YH8HgR4XPVGjgHeC5dXdQWTCSmoh2IBKe6LoGZZ3G+jWcEV4dmkIz
m+qaUiisZwMjzE/pY53/+mgX3ciqNJOGhkeKUUgL85hEN5JSk28s0ViVx+3D5sAf
S/kBUdFZqTOtBsA45CfwowLmviuLzsfk+Snsty+bef8ZAdxHFSEkv7KOKsAD8sHP
omoRnPIXHtMAqnfTW64vqOU6cESDfgoDB4EwJ9Qt3Z1sdiXplhiHwEF442pJ+d88
ddCPfdJWtPlrCGRGE604VvTCLr+mX/I2GZqMHhDpDsrY6QV/zS76ApG8GFP8s3GY
+Zg0+aI0uJbPgP9EXEE9tiBSJgd87zQ6IfYAY3DpNgpPRFz4ddelm9UzLg3V9f7o
AgHMu/GVbjUjPoRNP32IpmYL83+vfgr5hXl/Xz+jjWj5vl3JN2MTXDiKg0scVKWT
Qvq64nT5eH4K6+ijEayFw6/FZvl47zIHi9g45KwESGG6Fs9njT/UK2iyaMAKCRjb
+zQZ5LCn1TFiegCplutVmWSGkuXxsazfu8gaRMCcjjCUp/WcFMF2IK4XzP2bOFIH
WeIltXo/hwBL2c8pBhO8nZ5t0xpEvK/l6qZEJRGpI2m2wQ4QfLkiY51Nk+tMXtb2
QDHNYZnVYgui5z4fZ1Paj3cfhZRyIADt5kPuFOwfeDD6ZbXaxuQ4yX/5v87YjL/E
iwzqy+zhG6ihpjWz42khFzvL0dwvVXJ72r3bYBnSipSKsqjxaByUC+UDpGdL9jj8
RCHXyKKqfvYYy6/ohWx+DpmRpoQzJOtD44UbY4lxfci8B/iZOaFP02sPyogGByrt
BCxEb7590Tf6vY5D1nVfennqP4le0tkq6QKRjuTmS+slvex3u6W0u8MmX+RcWuE3
n6Hwor+/GDZRFDAMAgNHVjpa9mhNtrrw/boaO8zs1Sk+qH6NbGf0WMzunPZKtLmH
DkUWrBoGPWozDzeug+rf6m5fFNw5ASv2Eq6jeNlvnOICceAM8xAjwAC/+w6L4ICZ
Q9sU/Tvn2k4DdytJeHqBnea9dOhu1BXFSqBqjwbOfRkFv+NJlhEvgvfCw85UcVVX
jitcZ33wGpuKfX9rgztGh8eovxLYWurGBwXDwP67PgPwF1S6n0cneNiirrNKsx2z
EZ5v9OAFrETafUzaGX4wUTaXLLJGYX4bYhz3wUXzbR0o/8goCkgW+VSrTrAo+BOL
njiwIOa5KjZ5jkgbDBd0iXdGZA4HJDgbUlLUMiJTYDSPmrsTJnRvCqj+vzpzypSo
GCmxd529dL7ir3eKcnAR78eG2/hhRGTrzFFLbBO1e/oFK6zZXU5FSW2x5oApfveh
8JUCNs0l9NSTx66JNUNYLFXWWVwfHScUyWBKewFPde0HBo66mbEnPZpYxdyd8dZj
fClTCNj9JhZVFF4aL5eNU0OwxiVHWySeYBZ/GJDk9faVx1CE7XdmbW/z2SGr3tLE
f15r6r8gfzTkP6CdD7RcByXG0OkGVOtyW94pqHF+MwR+0e45b1kPIYCFfd/nILr4
C9HzJHrisBGehn2UbC9tUEDlgW9IyGXkSttzGLD5UZ1ovAD53mN+haAuvFzZkZ7M
w04pIfSxIcv31jMQJn1H0DDHFNvpqVT8e/4WxIjLGUR8RzsNU7r2zc2s97o5whHG
VAR5OjrLcqkniXT1enzziCodzKzSPRRN7p6CHPgOhfGR2jh6HdgHZLIja7K5enu6
mpmsrwAvg/7lSKTwiOnl6OVElcSRMbGtyTnw0lKLyySpKr8Me2KD1jTiMPlGsKOe
ietDJyN1xkLMV1CT+CzbS0J21kVGJsZNLlp7UOptZ4f4BGg0sCUXqlfRqskicJsl
urUCtlo0ZE9U8H8RtZGTneG5iAJt+2CdohkB0T4/4HVx1kpRd61OEdgB1K4BF1gn
VxTPf+fqmfbdWrFItY/M2Df2fR8eynlfHhO4cN+fqFSotC34IY8QSDmITFrVi6zj
/EAPZTgLJDWB/VhZ4ITUqSYjCtVIlKDLjtqEVCsOYzCGwp4uzsIaWWv2rwe/S3Ig
y/1p92ulTPtvwZsUrWisf2iubIOHUg2YQu5x011jHRQUCZFf2KOiO3IuVYpEf+yE
Glv/z3aFbPHFIORobTQ4Pmh5GqHyOh2MWxh/9uRME1/GqHvfrPI7TbJCWzSmTYJ3
LtcYNfU77k0Qafzx4O1Xl/E80k0LUuSd2ihhM4QCBW/SrhHn2cWMWloPZG0sSJtk
yD/kxNhz7yogcqrgJ80B5mVWlahyNj1MPs7sspIXNk13GU1+PzZcMAhIQU9RrTW1
Sae0yh4MkZefmQ2k2fwpLVeSLUMZ5xwtu6vXetyGDjbFHJ5Ch55/evUwbaPi4Crd
sg8V0JI48Adt5S07lvGPBzHvBV+7SL0a6fF9QvGZYICEelEQPZ8WB4874+Va1qUe
wIP1MhbwOFTSjvoYQT7pA3Qwf7+H9OlEM1VKg/lQgOTVj+vHtRCMaHJmcs6DoZUP
lZ5PQR2XsmzwbXFFJfn6EYn1jfDoCeRNpa8WZdBYIR+axNTd1kOErwWG24BfTKQK
NGI40zfOsm4H1/2zzgJdFo9aukvlswIE0sBttUJSo3r/PDU2q/T0V1QSnPIqryNe
3HV9CvOUdz5vJhDIMkXlyOy3JXBE04d3dwZOr+WctWFjwNqdTFhqNO0t37eizQEO
Eli82trpHCiFTQZkDMsbQ8bGHwhQrmDVLe8+OldcGOOZfsXrfB6TC4EOGld/kHrr
N4pPA0MqzEY+lBzyaP6eEj1cIh8KTHF0iu1VfH8xBPfa544BL5rXTILoKq3fPD4Z
vL8+uN/qBTYiZ2Q6j8l2zqD9ZxmnLYnmLsKiFtujftVw4QIjplhyt2WfypIvB44J
H2l0n3wL82LKSSDvDc+0wAcZlK7SR+YWMZJ/niY4fdjf11+jQV9vw5jOXa89jRNA
98vtbYWEa7n+NlCPIeNVJ7QMCqRaKsIzU8tr1VVcpsxrkZaZKEhXEJ9PRsnKCeU7
Kluz+2zgQWbaUhWqLTqdJ+qWrWGMz6hFeRDc/LJjcOUw74uwXoS6/MMsHucmN20L
6HbgccgfgGFGHCMEcwCG/MeNsf1LBXKOjM660xlstuDnx3lExeZYXqvWEB/nyMv/
nDKE+ieSo1X2GGJULSgzrwwshQ0CiF5lRag+4ts775+IdiptqZjGyPR+EYt+M646
yEG/6T6zd4+u5Qui29NszcUovLyAOF9yHbkt7lRbmnXkXd9WsVY90hnCDH0vwxTh
VkSWlUIJMukeliXiFbdI/EUgaiooYleDL03to+75xSyZATGAzUmGAgym61H4qW7z
Bs0rydLQqDOxD71zmFEBLRG/Zw5tMQzLKrCXidEoDgT0FK4tWHWGi/uJcIEe4HXS
C8otiJm7ciuYdNGvNr6o/Osa4jXYS/8Yn8nTQYxXLlt7tAOmBppdy6QfLc7585in
2jwtsZMGnp2vlTJBNyxcItMR2yCSwaprSVHHN1mqmh+BTQ0a7TqG8B3TL0eLn65v
u0am/rznrypI5S218OcdPcqzncNurk8xbvqaJS3RgWWqQGjiT2gG2dbJF/gyciSL
X0AFq1kcRkPmrOPH7I2rIjjEbfnHEZyKYeseAI9yxJlAl9PR+5f1lJozDjcou7iH
Ct11YBONFkB+mbnaBLCO1H9unS2W3JGwuz0Cpg+D9NzNMZBVUFW/fOwmjZfsEaNx
bUmAvxSdXV6Oc+9h2eJnfWzc3vooboY8pn0iJaSRI+jYqsdqCCQtOfOKfH4z8NCl
fCLBn4Lob9g3U17kCLUuVptVwLhvOpKeyOllf0KZvkiTXA4j6nfEXd0alTZuOgQD
llX9BuZJo+7b4uAO0SyENZrWLDKL3wQNoCCmiYjf1wMod4qoBfeZfMgD8Wn6wLl8
CzP8UvEDk/LzVqDNCWpUOeDc9HUxpfLomVS+xGHdlxcYiu9Gg7bNlgfIPR0XTzOT
SwdjkV5KlxAbRrP9g0ZrDEoJaJks21uPzRidYAmYaKFDj3sG9kbHrqyOKejN7icp
A+2vjrWW/nlwaw6EmnIq9NpEF39B73HG1Q2eC6xF7locgIcdgh18Rtp6eUzgF48Y
SmC4Mp1T5HDkwfq2Ujz/hO0F5JXB6uuKKP7lNxncAA9W0f5wYSMwZzjlk6f4KSpQ
HceZkd3FdhNAMP1igl72NzIgsOXiDfuXJxbbUplrMUwIwRfz2av+R8elOlimTgDZ
aj6tQumHE8+M+N4i5+ThsKJkcqKYTe93ClMv5rFlNiZpV3uma755ASwV3Bnh2iO8
iy+8PCmUat5RWr6evZixH/6NcB+gt4EB7eWlAgU+v9V34kj4314cgqT8KgyZITn2
D9Pw4OiBZNvIf58B4wt+kD8N8pC8e7LbNWhBzcMikIvC19ha/Xbm+qmQq9oJFgFe
jJFn3dmXxY/4U0HPbo94XfFzT2VV9/uFChtXdneP8/KYCFxo+WLJY6C2h5cEpEwR
ZdO9YoTUYC/jiGUE0I9+LT30Wq6NJWPmIKk8Hz+yp0/O+Ko6kdeYk1cYwBOq/0cR
KnmlwjMcTLAwn/CTzr+xYeGAuOm4K0XCyzaGAM1rReqvuI9Rd3p3/kj1+/1LFFQJ
T8cR2NMPSg4ZST3CaGYjk+fsqFKucwetiz/Qyi5hhE4mNxfhosISPTm1jjc99glQ
CXxsXX0hO9W3Q0x6YEaeq2WUlbZzjkYQq7m3AiFDrsWUoOnMmcIspHH/k/JKIy3A
BvXBU0UFFFe1FP1sd7lfgclrio6pgqYhjXcHiznCrZ2NO/y2WDDqY8zCq+P9AuFT
d+BRHbW9mgKk0igQe20GBivQTb/0sfuclaqR999ScMUVcsbk+4CfFQDkYISWZY+s
XvBKc2On3NqDOFvjA5AlwAL2sPW/7Mw0VZsozboJSlB1mu2qc/4xAHidTCJIl2ey
4imBF9X+nMpoTlU3rMbQROqfToYRsPu+ZT+gVR/DPBXiKnIE5uXsQsNtfjPC8ZcM
/+qelEPdEJsoiqumdyUDuD4oSsidLbX8dRfAEBwPHGmaubMVV5u/zceKlCrKwArs
lok830c/duCzWWw0wMyv3t3N2HwMaW2QuKzDJDQa/eLcXE6Yly2+HVmiEh8xXtdS
NJqbSXqUonP95VimR8HFSDrLFBkdj7nMARZ36zsqSZoMiU+fx+bG1avESi8Xm+I3
TbTaCOYGDfu83GUn8kKFVF8x96fGoMhrvWSHCbuEvkaLPp+tddTJLdTMGzwMVPLA
i7G+D5z+Z7EI8IdQkg7Eh7MjC6+JvGKDTbq4ykcuut5e1DbSiqLog/6Y/KJiUPhl
r+CZqdTxvd4UWMnoGIYSU8pn9OCHTu2GbBGQDoSJirWyUCjGJHf0ejXW/b06sMXb
AeVdH8AmnM+AKwEm5u0/De5VjypWXDdWTQ7k7N986trPmDoOzK6Qce/y9d5dmVXZ
rNAkwgHgF07Fl4ob60eFgu1b2xKoCD1CRhOYNF91Kk/N6JJKbfgFdOcZ2PzxGGkt
FRKsSwtVhL3zxYQn2Tzjm0Hyc1VvhBsC/kshhyNCpr8wTtF155riqD5TS7zLeoiN
C5XYY8f3nxgNGntLXJbq/Bv/zEVlW94UixmW+QnDgXO5Ktz1/lxggsfDn8WqO2m+
+iH3WVEutSQMljLFbDZTyE28laLBCSzAVftjW42X0AscyGGDCrrPKpC8PwwxhXf2
XFQDWxnj4SVsNM+q8RfjCDpLGxG0TJ53lkYUbO2/rKIDbUO8u+vmBysh5OFx+J5w
w04FyCxpYus4pXq6pViuwe/vz1n1tXzdERf0dAU98aFze7ek3TBThPZJmlD4bRKl
Grr5ByrvKg92TNi8/S+hTPABOmU2T7L4qc/MRy+3i07vp7bivq0izK3pkJfYdgC2
IRVWck/udvPEmozlVXgpI4punJKA8FoNJLhjlQUhdCF4n1dYhUebrGlJWq7mcmeY
g+3WplJRrJCoanPh1u4rpvFYXxN2jpv28N99ANT6YRWgFkSzK/YR+2Nx0dCBRThU
wLBOvh1lJOmcJxMn8TzbvHyEFuPbGRRfWUrR5iEHQZ4nbMvoqdQNShdrRvPA/m9v
VIJuZGPt0gnnxwx48qKcym5J/YJJqTl1UGx8P6ckuPzgemXiew/CYS2pPZKiVmHK
A+frbM8B6q/Ny6hJUWZ+8X7OZocTcjLk9gQT6vpUxA7HbmEfBemNZz1Hd6ZD04VT
/vjzXFZY7H6GB0xUUqRJJ57+GQ2EpdSwE/Xa6rYFvUC9ybDI4MVDgcYajjcPQS99
97784OfNDnq5EFNDMO+bBIzXFB976Rv8g/kCrZGmqG4wFlmo6gpUeCj4ce3bIWcZ
dfTiOSuTx8aKVQgRLqeWqr9tjYXl46LhOrzfZ5rV65bnTb7o6xzpa1m68F3q8zYC
aR9ZdEoHBxME6H4Bhp47F0t1X78a4CJ5dyt+4FTacpVE8ILtgEGVUs7zJ8/zHTtr
Md2/s6mKr4qx2oLu07sSLKHtOw5Fx3BGoODcNv9KOb07yVUjFtWUE92P8P5afEbY
hurILzj7RAsliWRU6VcdlK8DieBtaY5WvQBDK14DKj8LcnV21LFhKknArNSQRU6s
ST2kXdCmM/Sn416QNsZXK5xYn0CKf7mxf/ib49aqxeBpHBl56JrzU+SeoB2g/y6d
xU8mzn0sx6jCDkTNMH1pyJ9LLnXFmdxMFsrqOSW6pmCxRCHzoYtr/9M4GDM9BJn4
2XQhnt3PZHb2sDTCDJHP49LVKvOeJ9YdXwPW8IEGWWw60rkJWyknmyUHyleRMoNn
BmNLK8F6We9/9zZ46b7TrtXWgqeWvSi4j6Z8hpCPbRkyrBc7vQNIZm6+i8fgHvhD
rDPti6lxtXPq6enLgHUuiPHFJkOpJl85qKPdLoB0MSRH9fkV5XBhOLv8IIq1vd2Y
t6oRh3vFrXRXR5tv8PrK77SYlujklv/8MneNLcV64aiU5lv/bzxeh+JZrGRvpagN
CXfYt5M0ehuB6yJ2KnFzsA3CPDgCoVlxfNu3mf2srEeQgabvLZVqYGUgOoIdKc2D
Z/SKG4Lrae5zfXDoys3nrt4ugoKFvaaK+CKzwq+bf4XzaTGIu+sMVOpBd/RYt4fJ
y5C1VK1p5FKFhgLq6uDetsMEwVXe8z55VhzwAZ/a4C1h7ESUuL+0m8moP6suUpiG
rhTPdByff2enHm2dFjmYecQCqXzcSpMA6ZrBRWWYKckjMKwEye7mRgG2dR1vqoUw
Lnm/kLFrC9tnAurNUtwIP334KkUnRypglTXLa7W0HqrocyJ5nDlSlBAfoNGx15k/
RrXnP8by/e0Bvyb8MB3csonvyrX2M2VywwCvl+4jiJqnRGO9O60objdSRAe69Zy3
wBvD2QQilH1FoEu4pxQjeb7tt/aQrLfZJzO2YZ7ZVLEae/RHsJ8wRW1/NR5dfNGI
RqskJV0t9nCegLMCC4K/r+UDzD0Jq5XEAgK6m39gppwy2ObptrvA3G+o0w1uLuX2
F97K5mdzj/hgvGUPUfHpkFeExSmNvmR/QPLanv5QpvkaqkwS27uws0W23TGxBVN9
jw09mrqvC5+39pUhg7CT2NvAqYzUiT3c+PD+YYkQ0BmV2zq9zhMI4/XvA72mdvWx
E0OP4ThFFmYXnGpMbl9WeNItBSeeRBne6muIvo1Q9lOAD7xcquw0RFAuF+5OaGU1
M9x3u6UmnxfCJ/rHlexqeRHOQG60fKu8EnJF1tusz61skImwAfowfAj9aLLwdiPT
5xjxHdnt3uEbqa1em8RMSwzffvlvEkVLuM6ptUFyKKjZNd0+24Mjm6pVOOTZvN9f
K01NzGMLA8mQyMbSRNIBDVIAcFL2ATzpnd/ytveancgVUVx8nt8fSX+epP3xGDcf
/iXkt3in2l8uZkUG7YAtws6IQx4OIx9wneOqXbQmjuXoHhj2x474ZjaS2F9iICFM
UHbRHF4DE6aubzZNKltlCWvFeTh4ixIyOPm++EYbG1tU6eoU3ETb5BMrKLy6KNas
SoXezQoe1guqMV837WjhiGUTGyg8xMwR9NBK2EU4RjnrXeNAN2mQrl+He+w4Y1iY
hmAaJOOBXX4r3vND6Ks5zL2xzf0MKqgegdpgQbKnnvEf6NHf35rBDdkoBoG2EuQ9
bJO34ckQDvwoDfs6eDRezZNOj3mjXxvt6FpH0woh9DKnT/ZvuJJhmnXhg3wTu5O9
jbgHJDzTkt0tjmnMkECnpKmpvRNpc4r4QWTfgMinzdaaxteBdhsY44VsrDS6B8Vm
8oruLTjyxht0JYfB9MLsvxzpd/vy4i/nXsEDgSSq7+xQKGpuCsL4aD07WTHsQOK+
ds/5HBgiZxcuRHXwyTBYNnLLL0ZnRM0csVCL8kltN7fRGcGhDhMinp4irJe77ISh
IEWOOFgesZ6jKRghMespHFVrnkZnvI2FYkqm22wQHjuR0thMoxukwmVRGbh9Ifob
xYAc+zZkZ1EwYvi6qltrGeKDbXbQWkVqB4H2Yk1pnZlfEGhAdLFvGWOkB0FBbqbf
KM+TuvOmcCouam/So/1ftb4wpGOxUp5KQN1rwkg9W+rspN5R89okTzMc57GhWvFm
tqzI8d8jOh7GDYR5bX7f4iotXS31v2r/a3UaXlvQGmyJfzQ2NFPmKifZqXVF0pVT
ORoHUgghVGFNmjWyrc3vDwQ25a9TiE+mUR3xVmGYwBBRKy7AssYBM7fT+df0iRCE
TKtVrrpL7whR8xBzwf7cdOi4HO+Yk/Lwg11xgq0AUyYrSd5BA/kYgreEJBHu/gS5
soVs8OC38ptU6R55xecNuWTOZndI7xM3wuD9PlvYrghf3yLDIkOA9YY4ospGVqox
Zai2Rk0o3H//R+UCVOz9lUJE6gYFW2TH/5GzjoxJovcAsdTOmzVVnfAQWwHAMDf4
Mbcd2Jnz2gUb1uCfIrKhG6g7OpaaLhQlItRoc0hCK2E6wbzcIiF6wbsEHqDk9NYD
5VByviEVATX6c88/lLTTr7Pqfe8nbjHruYql2NhyMO6MwMGOGoMGtVoxmjNonhsA
ks6H6gmwSArN5Wt4eSXu09YwDQjPrO7TvbSYd7AGKcdVxbSxBH2+CPzo2d98V9U4
6uaB7cJoAe4H0/L8NrwzQIvW+n2Fp2AWA5jhGG1G5O/ePystCFS96MJhaSly1bR3
Qv6FqRkA3I2ccMS8/jPyRcHgKLzdXOPnIVIQkDSzSk8kb/1xx5RHy4xl9uX7zASB
vfof3YSE0jJSc/mkw/WNZ2RFEL5xx4OS7vWeXqxm3+9MLUIO13FKi674/HRc6xzj
OGnL7M2aoyD3LoBuoGmzoqe9/vRtIgg30Yr+I58JxA8odJoAKd6SL61T9aVBhJqm
6NmZIGGG3bKctt9HvGtahQuGhITiG1tPm41R3woGd0xtepqJEXzD/uqJPEXPffiQ
n0hjiVvQrs02MlE8jZZbb+n4thjEpDNT+h8I1yo+MBATSmlr9DE/Snq+0gok7Roz
CeCPWmfIyDAOA7xDVCNRRzND1tDo+DMbtgmozU3+E7+BU/jW+4CTSstzHUJBhMsH
xy4Jc+WiPBFeWoVFbmRjlFlFT2VnwG2W5W/9yxkb8QSW5iUzWSIq9KhbsduMLWmG
jPL/GOjq0i9EqVTg37I/mMrqzn5BiWwbIjzc5yzOamwVCglPZlaiauoxfLmoSkgT
bSeIYpT7LNg8Yu+cGNtM9joeRyzz4H64RBp8Fp+Rcwb3vPneBp/sLGgh3FjUvJw+
uyT1JwzJnBIiH//bmXN0ShEF2/Y+Z1nIY6Qd12Y+4QoACVTTJLauVcjHwnewOYYx
dAGZJ+wYA6W6FkE15MVneZZF1CZQDXrWCENPF7sTzQ+bcaYb8ll9J1O5evARv/pT
DvroCHPUNaOKpuSykZtgVVH5LExcnbSmcysM7PwUPrDfTjtCzFYTMgXkarM3SIZI
30ym1jCpYrVQxXLT+uRuRQNQ0RAvnOiutz2phbFCgQZDDRCdTM1nQe7ppuEe6QgO
KUlT7XENxdC8Semi3cBWXUGjO9+JU0GxqlrcX4nrGdthHGX9WpkWGMxYVD4/MfHU
PZpLUF5OQXjR0Qg7MdCdGA6R21V0TsJalOTtzlmbdmGjEr8TGxJNUUJrxgchKLsQ
oGbP4SKJAutGEiPecYzF12eLmZJqCYdyBG15SfTHn241nW7R+p2Dye4+lgeL77oh
zH4e2ttjGOxSAJ8aVZEL+RYrESQr3XVDLZnboGG28n8rVOJbcvrDapoJKc64xTPg
B314XKaFAA3JTdjycAWGhFTr7ep3u6CkdqP4HnuKp3DJFPmw8NqhTSPRBKI8Lua3
XsR+IztcdShePtn9Wr3mOwX2sdg4VoIhQYvPEv38CPcDjgz6vmV8PqQN7FqfXftU
Y7PBZSZRziSECgT/60mDBUgI0CVu22U6ZBT/bofNVMXt0KNTHjk+IY5aZNZhMeXC
TXLXEC21lJg7M/sdyc/Rz+GAfyNWmWSEoj59/zrv2zpKGZ9s7ENp9ooSEYAYDhYz
jvT0taXLwfeyMe/s/uDDnoadmDcFFFX6NqHaTIHeaEFL6vrt0Pzz3GY8H3/jlwaA
Qh+sbjogJOBk3GW66zyLF+S5kpBL2MP7iUSNIfhLSXzqC24v7AuHAcvRKT7xz5Jx
Dt5pSpTEJ9A/K8eTRavuPC+DSbeATCsUYzzRjehmCh0sd9CH5F9R0wkJL6YY7gDS
xu1+/nA2GHXEr74Ppt9h559zTaJ1GqzwywMdKegq2/HRNWeSO+8lgWbXC1lY2/o0
hvXCaNBt2b4ZHII9MQL6MGj3GbZNjTsEeJOA9tLTNQWECQ346V0RX14UBDhIrdfu
yhhvJdKhtN9yOL6F5QwgqhmVtB3Ip8cdSHZ7gaz/AekOH7FVthBI4TXjB6u+g7gt
uICJl1ovJkdBWg3RTQYIjxBPOCPMgMSrSO9vdKa+z2B3omIOIQetNBBE/3phYaMJ
NXxvnwX/SQBHJSXpq7MDZ2SNqo1IGglQlv0kfWhTx2bp9i6cbFUaBwn6yiMm08HE
71WR6tBYQmbi75zzGH5Y9OBIb0HMhB01PHK1Mb6o9S33SZQ2ZkSnR42Zx5y8rYSe
F6FRM7lZaejxxvSeYnOO73uRUWXZG4/rrlRmHVrRSq23ON9S1ZWzqSo1mtqdueDy
UTqfs9lgwJLuu/ff50gszbr9mV1ax0Se3Y1gShpTLvdPGCjT0DbkJFAeZqlZ2fK5
8/Wcqx8Nk7DSsrHCeDhhe/xHKQIP/I5RTB/Ea1e3c8VV7sYOgMwpPNXtiG7iB0Fc
QAZ0Jw2SYkssnJYJSmlDKrt6lcw8+iatqZ202ZAFBPDm3msg2XQl0EVjHXKMdjDF
KX0A070sBkIiLI2Qck9orPlbcJCSs8lGFPNIqIKjpxqCkI2+45EmINlitpMgzv8H
OIItD4ALO4Xwlmdl8qAoGN3JCnaxMMVnjxDV7GsSwsmCEH9LvrpfvuG2bKqNUiKx
EPA4/cq6XImctNGpJ3JEuKwnCE+WxMX2RdUn/reuIIHLxJXOYc3p+fhmGxkpJtGL
zwhcbEuwvauvE6oHRj8QOUN3VvSSZ1nKigduer/Aoiqkk/IYcX15X9hQNi7Eatx5
z27QGQT0IyCa4wOIu0D9+LTEGFXyNPANFYglJwURWtoe24AIM4tmeBHfzZsbOA9B
JC1Jjgo8smUymwgTbrMCUCVcj5tYJXDSZKUVn1Re1eHRGmmRu8Sjf7pjhwohZbxE
Bj0MCKQZHI22tUB5fHhSERI5bqbtFazXjyVdVRjdQh5ZcqS/BbiXj9df92d7TmIa
Daun/jmKiQ/bFlXT5+dbtOuqzdEJdIso5MoY3Rp0EUB3iQM4OwoME8ebwbQGFZtn
FWKmSWv424XhoVxavUR5xVSJUbxvB9mur8yGcUfyvGVH2NTNJ0s+vqh5LlsiBDfP
CR2BIALOGRm2McyB/9zFXZhtFW/N+cS864juEyz9ILmTNEpcr8M/s7Sx07HxfG2W
FFKO4An2vXSwRvJpz7727CVQ8pptMhptoEFBUDkyy4uNzmvo6s0gutU4j9qOPu2d
HO5mUQ2kqkAfZkFTyxhietsDd9aB1dHQsfxV+SCpgUDDyLkFL7o6P0PBjgD63p0c
/74sQLTx2sTWUvnhyInZJ6FsOBjsXmIV5M0ecwwI5pa5BjoIU2ti2BHcOI3NkR6c
HhcpDSu239+mPl1T7nLO5hEwewraUzoy5MVDLaBSCgWBo7rZ+hwpdU+5OifSLsP/
eev3L55z8LpmJ7NZJwKdCTI1rTgx+VWIq5F6MdP2WqzhQDrDCbWR1Am0Zceg9/2r
oeEyqb5+F/N8WM3jPgwoEvrKWG+CggbekEf9J3Dx2377ffhSIOkiuiQFrfv33Lnp
VreNXDL3sequV2LAlH1TwDprBT6cJT7h6Wvr4LyLmcf7IoqN+5G9mH+yzIE/5Tua
Q9opazqC0Eg9t3c+NM2rT9mMxi5n2qDKCazDDrs5/9PkhW8nXCPap6n3s2titL3S
Ej6NJ38Gnhxhii/7oD8VaOVO0YvUgE31eRjbO9DcpeiMe/kfi71wp64UP41l6fes
MMJTO+Q0Ua6o26GGJtb6sHTOky5FIU+PFM4jnhVes+3TjhMOokA9+7AZFqqZRsik
dQnQXXjn5Y1gpQ8oCZKWnshuMPSccKjHOdetFD41rkycc/qfuJKgV2XHXR/PCD8Q
4xjtdU5eSpsScrxbPzupC5mzyjBeLiETzVXDL0olrrgxl0qQXCmlDpgH+8gJToye
mMXeik3AwNoeZARkoMRb0QzRUOf+Oi3aV15ecvr47uIAJdzr5ILzeFqjbRr5kBMv
Pu4kZfa40IdNH9VRiulObG39beGXjV7vX3VD0/DJV2JYzKBn1kZSsA4nT1eWL1uV
wQJUzaYJPrBVT8AI6PAHu1NsxgqUhUYQzfS/qPW0Ya5YHFd8tIZqk1TTiR/OedN0
W0HjXWtvtdys2dgosyAcRjLM8rRDA12w6QD+t7HpqqpyG3bu10QlkGVZ2+1jy7n7
5mOYF4tGXs3V5PHFEEJROfDL1Lz6WEQV4XNgfyMM9lX1QdX6cqqVAy38BQOPUGdG
19vxyv9bh++fqLkTlw7WlAssqEv/K1GG4BJ/n86fPNh83v4xkvn59X+4KlZlqnlb
N8XngGV1pWms1sZG3aEE6wFv2J5vZU+CVkj4zhB4B0vwzCXU2hWcuWXRjT5w8RqB
Rd+05thD2Z6mz2kXoCs4b9ODeFrtLrrypL7viGdGWtaIM6ac985Cw/cCvyTN7V9j
qWt5Ag2cUObq3F1qkMZoLlWrV/wFqWzPJNxwBRu4gv/qganUXjhah/Jsua5bFzwY
WyQoUOT93HrD5TotjwmktvUPaL8e+CGCpfGRPGiMc4Qjgav/SgZJXkaRIpNPvXY0
e2BHSNvEfm0uk/A1dMMwyC7tnC3c0pIHxCyMhU2TqkN0jAL3YQyxX5JQstI1Q6OO
6kjVQ/j3nOG07Ash+YEmsKyFvqo4ut85Tq6pUZCuHzlrmMskbE7eRDQml/ASULeI
51m90bZGrfD5/NZn4wNSLBi/8IjQUHBsLDqLxjHbnTTjtzxGBrWlu6CPVvwYukdo
rH+OLmOGWFZhJEYOP6SxCuHFvBQTkQ0I07JFsFcPTzvhiTZ3nmWVyb4AFgJkYfix
MXD+MUtROlzaNsGbSWNU1xHxGT19xbm107OqvBf8vKF6ostz36wi4IpimQqb2vU1
Ig/USnSPFGCH9CGRNbTP+7bcyRTXeLV5T3pVbc4hroUDUHzUph9G6n15nIG6Akqm
b33A1RkLYdBXkP3W8OnQbN+JniP6fVv5w0VzTjUg8LR3Ud3j7M2+rkpKtkK7ET+1
EDe31bCTU0p7Y4LdWfHaRByMLSt9X/gX9QhHBXjYEQYs2e44ie58NeGFYwle/3tf
aFGVpFTkIlbCnCUE9gnVpPfcF49IkzvcUB/0fS5dRdXWWWBJciDdot8Fs76TKwwZ
J9o+ACyEpmEZWPLAl8AEuZenWygbZtQpfZgCkdziRlNyxjVMtjYx/ERZD1F89U9G
tnElQnWQNDqiLVvP9+xGnTqdmq3q+zgDa+offgkytw/LNRaC7z1wt+OkJFX5ju7x
IKWFtavsageJW3kumtjRG4JnTtaICNGbeL4gWM3pcI/GajUBdx3I9XORDmxOcpyc
0yjoJ3zaT7YyiChsQg2M2RDxC90GD1OF91uI/J1ZbxnpiMq6f/+4qxUNYIVfR5bF
d15Ccp+7eKTucvGyLIp3JH8OJIFFfybxkkL2UXbZ/3J4h22p7IQUQEPLllQixl8j
pnBP/S7TWpPZZmS1GavEPX8Of9gYXvMm6rqI0WmyYpuvujH8ACUYIFGo2ME8M/rN
vsl6/bk8qPieGbR74vHEVyna01x7Innttd49vymTJd9dF3t9qaEUfmjDP1dRzEUL
r2tYm73KPdOMCTLEJk0+DWSCen3QBH7ENL8bRDiu/jaSBjSPLdULRqesI6zLn1w4
exuDetAvQqxlkEj5ZE6uwVOH08eQY8RPzK7Pd4gi2AnNrwE8dGUHcyZ7Hwb4OEQZ
RuFIF6ou4dhmNy4kALsqqed5H2xgn0767GcXkUtx8frcQdkS0F6ZDpbRw6AM7xaC
KUELoneU5TNlsAEmzYMV5ELG7a3oHkyN1qYT320YOYKlI9VSJVhgk3flfLTwvJcn
CaoLpdVPnVv19Q1eHi8iivH3lzY5AnBdMOQsrA175UtjdmpcFOsyhS40X5F7R7vX
kn2NFT+7HyNpBJDGjugnvNhRBM4qELedmPL2dLlYMMH5DPNoQQS/1ShQ3OqYJpXO
Pr8xvXglD+DWaOsPslLBmJji+AxHYt603I/qhrUCZZtsSNQe8xpiy6zUp5PDzuB3
yUWr9qQZ5lRML6cVPj78Qytne/dC9ESPUZAliN3kqIo7eLP259ZsdPgCERwLgnvI
eXE/tDVG7xCxLTV69HwVTXYkqb6M+e6qHMW+I3k1EawCWjKqWZLb0R2Z2Hz+FPNR
xPqXjC7sToOlllElZ2038oqDROdKX96ZU5vAY7T/WEgsQBa7bRu8XNwf893+AeW4
Y/JLz9bnV3IiKI+mwp3c7fpKQSsWYe0s/6Ny24k8Ei939V/xOgSvNY92BROXlUuu
NiOLKeaenqrtlGcuih7CHCuB3vidtg8DQxfJmnIkhJzQYI3uqtrl3i8eqfG49uFb
U8CUnsK8jqtSi+9Co3H/iX+YmZ2nvH0CcbnV7PCPmOyc6Ig/4pGfALQz/Jrc/Y8r
drZacI29AMiQoTpFViwFXQ9UwWZV41EtcuMs3DvPWeW76ZqvSWC3gGwoQCjg37Jm
JGAmGK21T4IdvgQRQbF/AYUTosmHvEls0O8/nnabf9Hy7JVk/RqGsmwS0UYiQPIA
nGUGeg0yW6c2bV4v/vfbUNJoZ8nhhRO8XJRX70+iDhcXFd+/Ur1l3WKCrROiGLLd
07uO13QtQstyekDq51sCgdZ9631Z/XeF+oLqGY6D8b9//jB8EPW+HWX265Riu159
Wh6pCsO5DkZeuXkMF3AHPtBWCD6AJeqx27twauNAbwN33ZJGpOPLqRNcZPN9PsEH
8z9xfwUdBT7nW66hJdUQeLEgZ+qGaGxK/9pWG6CB8kv8AMxna2XKT6oInTCmDFFr
3dYWaSjNLOF76JZHlYWFKRLn7iWjk9k+nfleA0KvznHz6k3qdRzt7K9OHxeCBDwb
lzjV1ZD11XWKK63X78n/PSi6Mm81etE0nBfNMb4pE0DiwGbYr7Jm7h3SaepWyxPj
E7QoRKuzn613EDyZmfQ+Qfu8T/QEhSBWUdcWM2bzu+QOrm7N4vXZ0LoSN3RbHGj+
aY33I4WsGdQZbVsW9eHmn1O/Imb6gZEK4iA/RceK22EyNr6OJCq7QEm5wROSYhF3
TdpMGPZIN3KMFXGMDvcSldAll3Ha4upJ7MQ3YwShzwAVCKGoW2rZXST/DSLtlmlp
Rip1CmZnUZ+aN+oHQbVBIPjroes4TheYd9ybCzQn8OLor/2LNIbIB3zUnH7hHvjn
0zJftfFTmQ+v4LnjKEq1H0kcluNgek9/ZenIbIAznMJ+qQmzP2gCmOONgD3kRYMt
TCDeqGIkqf9apQgqSma52x3KVNfL/Ri+UCyYbIQ61eyt2C5xC0fnRJSqj4qw1WhC
0BwBIOUZ176+RLFijK01V9PUnIBI4dMif1CBwKher57xft+mUtkbCeONVDhyjCZj
rsB0VxQHhuP0k8De8amicEcuAOM3O/yBejf6jR24vOvxr8M/qNfmYlsJbK++tnjz
XyI3ah9YEqYbFgyfrLesRTRW4Lsdvjsx5BkQweta2weMg5OWn74n/IUV8JwVGKz8
uqN4txJMfJEW5KMb37mr9x8drD2eM6kRkVfg5PNebPP5cdhQs+4pmgSAlNrsMkHd
mRRUeECuhlXRFnSrXPNrUDHgLQt/K5p1lb5KoMZ/FMfrZAuaTFdTWQ5MOcDFjbY1
X0YuNE0tCrv5EcFY7ycew6vRBeGg094GHhxkspO8WL9Q2rw3PY5+HNV1WE0oVldX
fvgh226lWW93XDaC8pSrUJK7XrPeJwhZ8UVb5ZA4NY5C+ijtCUl01rpaPenZ6L7y
STp/eqAqsFQ+O+LUBfsBc5gUuRK9OEZ+6UHda/1THGpsiiqN7FBlPBHYncO+3a4Y
mNROdLPHFxab3FzrKl7mvxYnd99nRlZcgFpiHIwiaAnEo7N5tuJEKaQDMi/60ggP
c3Z07/aft49BSo0B9JaDjkhfcBakc8773dLmqbvmKKS6U7wM64zW2gNpjuH98gbm
9j3QNYHP+WcV34HgkTJHFBWRE4vWRjVDwXTXGv2xHt0aQMiKsy87MDka0TcRuuqF
/9XLi8GJ1OP002YQ+CtrBe++I/XP+YFY/N4SwDF16T/1hdbs/i0rIcxG4zZJ+xGK
nehs+h44O1lIEVx5ZEbQ2v1Nk5NKeHVG/fIVfUZpMkUiWfkxFZjQVmDJgy+4TZyM
xKNktGh/GxMLuSsbPvznT2bkVtIUlmMZMdckUVnXCiakwj/9zzZ1BuLsD2Dd0wWP
nriNR1ln00IbvSBifKPpWQg96eb/8mst++mMWchQYTTBzesQt/qATZYpB2HBIg9/
QInZ2T82hJvk8yAs137kD4qWhOvU0SERGYK3zoykfix/4HBX2e1FITC0pA/zTxme
ZFWE+06XwJ7TI+hZ2brVNAYL4rU4er+z1re0T2zfGGwds2B6mFcJ7ezdmeSP0qZx
3f5MT5eU5xZfDrJwA1JJfv1VGYiMnk2ex55VG1E8nm0mquHilE54S638dSOG/E4R
dwO0i11dnyw3KjXauZLGvYDpg59Wc/QUhMvacgONCJNEpIf43v2HDFttXoMMofzk
In4O5DfgaQOkZzxzXJnoS/Aor3LOyjb2fW0/4MXvQ1j1RGFl4ra68Lf5aq6gKVUD
MUIfmCG478sXSJ/y+cBn3sxc5xSTIH6kMFLNKJf0MfeypH7w7p4xH2q1uvUdFSAz
yQLKlau82MrFgGmM4f9W/1vJv24AimePNmKSLEbPxWpAX3VT1QUYIT2dx/qPnrH9
iRYHf/onRAWuBVKoVp629IFvGLi5ibNLik/g6ivt5+o87n9wTqTv83KHVqbyWTzi
Dgv7u5leksMFw7GMOjwkW9kxcpWg0+iyFypxOF64IcTLgKdiLrCNgw9T9taeer4w
QndUVfkBjQ2FhZXqTeU8qKS3Xv2NT1eDlnk5ZeWd7Mf+zfwEruy7gVwDbAU965KB
nkquRH/sbrBNrt8hazbj41FcwMqcCvJenMJin8jW+auJTkKDryoTwQZtB3pLBTV7
ddkI7mu6JezBRqK+YqNd7IF8lRiAOxBfFuOsJQWEpVpVHqgrmcNDpMGAn/x5siNZ
tAJCUncrtib+vLQc+NzYwg/fxwx8fnxNIfqCIJDrN78ADZCJOhyzo1xDKIiU/Xj2
btNuC2ByPwGLGB7OwvZHzy/qplu9o38+3Nh4lpNX1++U9bcI9dSM+0hMEKVCb0Z1
RaN4LQaiHA9PnE5V7PudC9Y14BdO52sxa46mLhyMdalRAaJSoNMweyC1d7eA/jIr
jO9ypmq+rE28LP38AbkHLm0Qe9TzKRrc8lYQkWblhl1JADznQnCSxR6IIrCSIgCl
u9AhLKg1g8asH43WshE1r9gzEhIGEAFR3KrzevqCy0QwMpEty0QY/vWUMEeEEU5o
yQpOd+AOFvduIQycUIKioUnnRiYAK8mWjpILrr1qx04dEDPYNDvWkNLPzewsHZSO
scBnjBf9n9Xjj5d7GdKaIuxZVicDJr+A8cG+uPKUejJriCx/D92Jh98CHBShFu2N
roPYxwr4cAomiUU7tkXMv87fzWR4HDoHMfveuVBEHBT0nj23qqaLfL9q+c7l5Eg6
sg983rXtFSKB/ax9Dednbfw6qbrc1EJsSRKZeFoOnQ4LY6ZOQgiDkzUC8Rj/7apZ
k+2OEfI0uPjPlHZGwAi3YpXtay0n3mCbEIMB407CJFxX9tcXqt/zUnKdkdm7bCPc
AY9caSazOmvoxGiRVcTdcXsu5lP2Ck3uNipVP89q8EiWDkHdXo3+URmjQzS7mCvz
VHi/M/3XGtQkRaeg1UPoytattZjQVZ7HSm7V6XFT4DeOuQtNd1pBSL3lTHEceG6R
amhHTALoa0n8iipRQptsDKENPXDRTCahjd+mYGF8loHv+4Z2nq7BCyH4Fasx4+8z
sMU9n23NKJJS1iq4hLn2l2Trh4NDxiHvmPPsAhZdfyvtUKu+WgO37Wuim5r7joaz
A1kb9Cm+mt3BLj6aGsSQDHBwjlYbiqm8ZkxoX72o7j24l1Lrbq0G2YcjiufkxwoS
2lU89p8QXB0UogxAC7xcmWkO78OnsAR2yYAm+sCqE3lrbMNHpQ8UXXBz5FWbzpEJ
lxC+t8Ay92uzapZzYajM+cMVQYlMoD2fh5Fsdc1avsEBX9kCgyoEwvvMAURNREgC
NsIHalLuIDuU+n3LKkvVOuJfXml2kseTD7ja4iAu6Q+zVEvY4TZJQBapA5kdFDT8
sOJS9KcBltAuEMVdXLF2CDrYd1RYJYGJdPmqxJNOwxPkP9OoHCPRn6QKAzY8izQ5
vPy2Cck7HL9elakb1ay75t67WBptJUcJzTbc3T8oO+9f4/AGCjhQVj2bIgtk1/3U
u2yqUaxSDxum7MKnhR6VOhzua8OQZbnxiM3KJTvlcb1GTcDaSOHoqq2k0c9Zm421
BsqrmStzYqgrJdcSAbWcRfp1sXB/tzv6jc8Dh/tNWSjqqPlkQwTuRCV+lHxKWKgH
ggHeD2JYPurcFX7MTTUmVKDDQx1QangKgeTtD9fXhp43iSvwYSNztSn3GDcapKub
cO4AkOnJS8ZbljHemeCIA8YM8sPkrj2AxMfgSUU75hV5DNFyn77e+1XQk6UdyYMr
fKeIILTDt2Ag2eHg4UiKbMreDhapuCYNRVSvrXEFfP2znKUuLbvZ8Nt+Ygchg1Sy
wsIMJe/oIECTox86f9ZmRPYMDcnq3GMuf9hA031XtvLyRcYhuKrO6R3AxoluLjq1
Z3Cxc7y1fNSvG1SvFht8oh/uS5+G84i9+Y+fkj4tzT6YHtTBAJk30EiG16MHg5rc
v2/aInWHONssXcgxhkbNfgSMVrPMCM2FR44N6fHlXecZZmDB4b0Prp+9oclIuf1F
XzRPiprmSNtximhO7csS9HAJMI6yxgWdd2GEVwJJInp7H0IrFxRqjq+ddik6jYcL
FtKgEP9IEhNbnFxgBnDtT0hxjDrOBixlhA2IdICJiEqR+EKDqRrulCkTt4mNS1jW
HLqMInlNTY06V3KHjmoUNSdhS77e0twhG4OS9OxyXZk4Ko5sM8VuHLIm/Ar9QF2R
Cyec2o0MQc9aPFQNwiDCEfGpzUupPDmW3SeskhnRIdWs3E9yyPtrLLozB0XKgwgm
n8xIF9egfa278gsskQD7yuC0sHCclQ+lvW3wnmqlvM4ShQBLeZZAUJfvq6CGi7QL
VOJDGzaP/ppclZulD+7v5oJR8SuFIujz8l9eAimzjk8QM+VG8YEPrs+361JvE5a6
Xky9lMQUPeSYnCpDYtjsOnrW00xiXR11aaneRHTcaB7KGIMYN0O06kFVBQLtqqUw
nBm7COdKpYpCzrw+F1aGAPt04akDcibczWznIpEMrJXlDc2p6LoNy21MwE+WRiLx
TGBLaNri+2x9JekDfGYtnHJ8CbOK+2EFmYUq2P3uXagLsSZv2WkTOmO8wyibeh+m
DnHivSvt1HxbBDM2USsFO6NjuByOIf0WrMSQf7AgIKB4gLIcxAYfTTsfJFhs8bZ8
PLN6JC0Y2zrW6kBIf4NkPnc/Vrxjoomp9DHCZcYnTTrtNY4AlCihhpXIZc/kuHjV
+UKEA83Hrs9v7vyf2P/kt14uLRlNQoqnAV63ElYmDDRQzHT796t4bUtzJ6x50bDg
hdsjMqiK8rNeGvh335sWvfUb1eDfGVKMcuF4Up9GAtY1wsdMDYq6VDO/FNfus48P
Q15pnxwD8iju6NR0S2hEc5+jeX7CSZnYtAyRI/DViZKc5AUTOM0+ZH8Mqd1VeKgj
AXOWK6EsXioC/O7aEfBPI8NTq1HMmZvkSYfxWQvkpjGRUJ2JoIIYB4Z4Uc6Rqdbw
v5cF1njMB01k27J2gW4x0j7Z1i93BK+Qu0fFNWuTFFC2Fk+bkTIi7wAVttINLSun
n93SR269+sqgOcEV59fF7p89nqHnGvYv4FauxIq3w1SNj1s6ewkqgvWoKrd3l9+h
NlZtJJlgzajvwKY8EGmn5Ar5Xk5XjCTmzfFUjnfP0l+7P9HLtGKrBZUq6kX9mnE1
6RSHzx1N+/GR8vC5GK2eJ1nj15qOPYYnwam5KCsDyIWP66S2vyxue72eOJ6qZkT/
1ensuUJp/un9TVvxro7G+e/m02kjHKC7HT//SXfVdObPLxAOJ2bHibp9oTwD81ET
YxBK1Z7oNavK+/H2XTUVAzslyfyJg1WuvHTiJT+HynB4ovDl0YKsfWQnUtbDVCGM
Swglinv5Ltf1ZOq5T/mueL5+I3DzggYd3L1PRrk5wmp0s7jNHcsuJPqBedfJL1mB
0jsG02KfrfWLYLIMf7hdzyZFhQePYtcrPmHNIeCKR41AWfmYuZCCJMxJvj6cJ+Jf
fxcJonEnMEJoVw9DOJypztuAh9ldx68bLbaSj9YZu2BNpdxG+eU8wBGhWUGtDkSv
9IUXu5mSuefSvxEfwoCOmqYUFHZ9ZAUWKYqqZNzAa3megmvZFlCM3Wrk7E6Mv7jq
CKl5uN3V11d10OEGoR6c1z7sdwp/pP6rJbZUC+ygIA07kuF/0JfhosypMtvtDYrN
mNjgV4kmwGNPUF0kJf6gtdoOqqI9rUvw5Djk/mhPsRWQ6Mhz744aQx+Dlpxq+p9i
5DOzHeooM7WxDPGId9HJDJ3v4wEe5ziew+zx6sbKzqm58AM8OppZ0NYJs18oAE2U
nLcn9wZmQZFQ1w9Uf/LZGSnukTbQnQBEJwUuq0tI3Rp7+AuXlPdH9izzd/cvamGo
OtuqmvgxfMJjRSRyjDOoyX6mxRUHQueaRH7MIjteYyEAb5fz7Bip6qx3Uxq+g0sV
2N1T07HBN93p6XeucFoCtwVJGaUyTPnfHVagbsJAc+rIU+Q7qJNqK1+T+DbXmzd4
IyEt4ArnzAHJafzHd0IW1OT2RFvVsGzXCU9nf1vspQDLS4zv+qD8v56xPzzLazhA
Kt/g5af1kU+hnn0/dST3qHu0MFf+Px1A3MtkWt24rjwceVJGSUoh8T7ND+U2+dK8
aDubtj3GEFO7xxvSGc4R+nc7eVMhxpW3nUD6yrwxrdMwJe0GBIFXu02YGoMvwoxF
NE/ngBK/VqbmGGB5uTpG0n8caqFB+z5NEuxR0zLZcHmWQTVWbX9CXOSwT992ftUR
iLJoalrfYo/y5AM4dGA1E1pPcJ3U8KZJ2W5ipI2k5xpdqIREoWj5V+RQ3U4ssTu8
5njigti2ACbPvI1GrDIl8KS0ToIG0ObO7zm+r7gsDBVHS1xZn/9Lnmysj4wnB9Dv
sN5fNuffYIevIucuBXt2RdpJ/sWL9h4F0oGCw953f6EX/Mor3+Xj9zwK9wsEWnLA
MYRNjFnWW4wUJyHnK6Lz6E1WpIRNFrr7tBukyhw+YMdBLJzIht6h66/7oZ4hIz4Z
b86Vh/GQ6ddBFsQLIRGohjiX6kzLSH9DSY5sDDGsPOR0zB7KTKbIzhdZa9jq2tJ3
BExATy6rWzC5J5m2aWQRgLNbIt0+Otd2/9WJfIWd1KYg+VS8TJBGmnRJ/kZp4WMK
CrXxfxluF7PORAo7DZUhPWNymlgSHMrnI7Qpl1jiTAO8TnJhLVtUVk0Nen5zYCdu
thr0YJs62ZUEP0sZI3JAqoQvEOFVGVe19/0C6X3D635W8bQfYTIaaur4nh+xnekC
V4PNW9W6VSmEHGKxsZPlkIRV/LsbLT/Uz5b1k24IgDPsfR3Oay+xYAsevEE6Lb64
OoUtkFa4lPBvZ2vTNZuPGSY/c/IZBG/Ql3kT+sic1j4O6+sJ/6RJdlTUmOIC/Ds/
B3XgQLcnfyuQ6l/3n0QZwtIX9MwG5inD6ySQwRqs/r1Bh5eSDOHWTBSahJUxorvj
AmSdvFi6S7eFHlY6tbUWrA3QQwI3CW4HlJQPDM7v1eG2y70yy5IV8KV8pRoZE5nZ
Z62PWl/d09c1CJ2oFZHkSjhFRS0LpYV35z6lFUU0PSm4IGRSfBe9k43f+VMNkOuJ
ysV274j83xdopVPXB4udBzaxl0IFAm9J02k9Fx27KQ3mAmmkBTFtgYD+DpW7gfl7
w1p9a7hp1eiXmMLLdHeNPYR30f5hVzEdJ3d8z622pabqa97KMQ/KfS+yX5TXphnA
v02Uh/t97cbhpbTvXXr5bqRcDP1QUNBAozpXm6bNMtIytYqF2SRBOJtD4BMkLjUI
XQDD/FfVUj+pVoog/ZEPwvJ/E/3knBfKaqABa67YJslCzGsXIbpYZn9niyYHwUn6
oxJYeCBkmWWwYn8JBkiHzzoe0GrZ98obgfrAcBOTi7K3sLF+72DGZBFoq08ZlhL2
gb4ccR1MGyfmcwNZC1MEuCNcwQh3bx2oaFM3Yk9+a/W+75hN4+qPjiwGIm2w7JTV
gJi4Rrz4lGQQL0l1bXq+r3LjdfTM8//NCi7SHIACJ3CkFjhrJH3d+Q0BQlyFvS+8
RSfLFXR2Wbk1bVsZq1iu8g9N/cTMfgDTNxaBopUkmjM3ECCBXlNIKKYa+TokxlWn
9CLnWT26PWGSARnPxiCPSFBXwh+D0h0J6j4i+Lzij36/HiL3fjGR8FM6W3Cwx4Lh
77sXOIcLlbqkSaLtPjveljc7jnxHNtnXQrgjAAsH0h7G2KjbTYPXsfkMBzIDw/Zu
d4/snCl8FyyV0UO1xVMpkMGCkc3xPBY/iNZVk8VkrGm+9XwpjoOAZJAaDVtktenk
a7p0uM6c0LRYJoESWbH0BvMUa1mDIRkMAF//Qsyd5uTTmzjj6OwSUOE/ONXQqsr8
NpOsqbz/xB2LiJAVRvBk6U5RB0pzBV9bJIR3X0rqNZ0b9GW1H/mSf5w1EL6VgpFL
gsxjdSlRgNt/C8N2bxLCma/+as3WbFsTzKYgiexy+z/dFLO9KPUTBgR9ZM51AeSF
8uCj3qTMZt/8sYq754ZW6nfAtVVFOgnHtzP6t6Wi6XsV0hdXOk+m8ZEmo5UcdDYC
aQbDPBVJteJZlLKzAwL3D0nOPKJBZsiKAgxz+G/m8URLuL2N5/IrLjvr5YmW54lt
V/6ZScGT+WLNuSMsW5kG+RxUJwigdrMzHpL5zkiehNv9Js4dc6nnPkZWtxfbewtc
GN1Ap6crX6aEa1GDSD3ypSRtGiZpjCxwerUftFUC2sjYLR7DvIhjI+MY5Eo9pVDj
zjpdaX2GZ1qWozAEm6QEplfwPHPeZ8gATqhTquOqKRYrgtMVz3JOXkokomWlN4qH
v6P8JEe1lyCXC4EpPdBVTqffR32q9vMblHrCGqIeEHiwRr0Q0FXRUVq3qOEhwIHS
PnQBklFWZUeaGNIw9rMFujgb0gbVIbyLyySr5QOa7DPoWU6c8T5c7dCcXgIHcUq0
xP7SYbAsIqaZZO1Dcx309Dz2Pi1dwfymZHr1MAUY7C6DPwdWQTcwYtNhRAT0WmQw
BTMV5lRDN7t6j5Ut4kI3pbGUP7RS0GdO9A2N5fAp24KbMgY1eqXPgszgZTNXnE68
iDxsDjtVLTV5IqYayhNbVTto1JvW4ndgQWwRYPFxqxyCZ6ymgbXekikUv/VJK8S9
GtlDgI+jgz13QucO3CDZBBZp+NngLajWYh7UXIhCApHXP5YiVF2IdwigF59Rk71t
4YJdhSJZGun2pUT+2ODmPcpq9Bn4YSnT1rgcZJckPu9Y8Dj7rahLkSfhu2U6Quga
a6MMLz+jfz7XhVUjmVbw47w0/UM20JhthHcdVisy9hDZCdobrKZ9sbjNZV5mTRxJ
z8fXbZXIV9WAD0+eap6pNyq6t8gxGdOTCksSBBZgxUEufUXLIvO/7kbGC1ttIL2x
6oZvl1oCWA4ulTl8YENRQnk4FuPovCL6ATbSN+ZVYl3puebX836tbn84uJv1DtCJ
GvKR6ekxeJCvvZob4dQruyKm8GyYLzefo/dMknEVqI5p62bKnwlnB3ZEh4gkQPzj
FqBBL/YD4SrYhosHcvuHkIiRc5b7G0seyP3eGkE7l1X7Qf0jircGRy6wH+4o85KA
deX2lNVj8Q1usQnnhY1UwqEJZEMxiQ3VE+Exg876+4Om7alG5udEf9buOToN7Ak1
bcbkIfa67rc6W+dGb0ja8VaDVvcLr1J+ROPIl2+xYWjlg9ZTuk83LL90ZmCCqiJQ
ezfp2/jnJYGiczgD2Xe0WIvHip9wulqheao6S6BoboZHdHZmtaqCYr9a61uikS2Q
ODUFm9PGoYg1/xKVYUy9Q5Cq3xo/6V0hfs21w01GEXoqwQVD9rsEN3oiCpQqNynI
kUk1iCaoTcWhBbtWnC1xdcP+sGMKg9yZsQksF5Bzy27rzrPFLUX1W/nXJX2+kt1h
f0s4rLwCKGB2dxnQJa6+RsZTWyyf8ZVkiiqHgDYbhYasO+ZOIaU/rkL6NupSKPmo
KzNyP/73Vi5k0lAbIKWJti0cegqO4xvwAVi5TmnV1bx7tS+IzETkYdJp/ugHzl3x
ATIoCmD3HD2LM7/RBv7OrrlSbKTvdxK490/wKtfFux3bL1BbC4ealPEoxntNWhp0
UvDcan0J6gysB28JVTlqpGi+kHWoFDzVAJW204o7MlHMK6iHkVOpis5kuj1TJ3Bl
9JufZFdznVJgSNshyepj/BN3eIgxgxRlnLWxftFLtQLvkDG0ZP+Qnsn4nvBcZvGq
Hr84vQRZ4QpNtuk++lwFJHs8Qyt9CDczA7ysRMWOXHvAJiRK8h8fgy6XWtHc3ajM
srXcnHZCs/ESdS8bWotk5YH9Zsl03dqkOkY8BJRBZ+DzcVkLwgbxUZWQ0Y/8dECb
MnepN5OU4HMK0dK88Dm/91kwnOQZW3+DTqpIou6n/wlNx4GA/XrGwoxHxzABQXof
ntFwTkUpHX7wpuO6ERoKdhw2hYYZbT5o8Nh/I4GWQo8JEoZwL/GirH35UHf+Vkfw
uIIXFMrh6gZr5y49lvCqcMeZarA4ZQz9BfxjVJr8BLw32Vw6Qa/8YoW2FvVAYy0v
FdCibQosA6qnUfP7gLJfZjtCx9wcioeu2STrjjjs4F9esIB16QZJo+J2JnxDUb8K
m7c8lZPRnSanH4CFvilFjt2HcmfKiO2wvmniD0pki5cAMDvz4+HMQxK7Q8F5ZTxm
AKryNGPbSnIw7r9fu/A5KF54/1XsPzH/4CLsnaSY6ws82BxjNIiw1OTy9G87jIKj
N2OkHz50o/uGNJACqP+eZlzS8hJrPRDyuYVSn4UT3qIhPjHCZHn1zfYJaOoVptib
LZwGnDR+2pNgDNI8RMiDlwDaSl7ZI1N6Lh6pR+TRQ4eiLciNDiF8P5TkYry7dAdR
yd5DQblXnaRal4ekvdK0rnWMC7Rqxy/C6h+H78NdEJtWftkJXpYyWni8Lj26MnQ+
HPaWrK8o9W5iv+vtnu2UtjJr2jr36IMEpVo8XSDAUttw1jB16KMz5hGdQELQJsiB
HxaWQeB/7Y7fxz8VxAzTXA1Uu75hgJpkr7ytKCy2z1pEBfbwpyYD+PPjkMPRnEHf
yKLSAGddv3j1ofQV1ITR481T8CjQ5bPuk1n8lGnqpYDuFuP7vvRLfHCtF/Fxb6Yu
OTQ6EgD/0gJ5oY5g/OPXP/4fUKZIfJn1t5CPj/n+W6teUv6ZL0OeEHhmwEudHz2n
tjSI6p53Jn8ccafzoIa/h8H3vbRQ5VZxvloaPubHSlfQYzHnZF5QOX8czKFof0ZW
aQ+uW/rs1fAO6Td1GqXgflvhCkTgeuTuvxtQPcIAyZiCfAtN+iILe+PhzXchBOPl
oPcMfurkUSz/ctocI5GCiWQU0r1Hy/ddGbtCjZEKnVr6mr6JN6nK/m+qa0WjMfVc
sHhXUXD7vsEbjvTnljMhzMXp67mymlnUBE0C1/FPLUIsseFxSFUXAiRhiJb5JWpw
LNYfcokaX9oYAL3MvlWqcMjASOZmuh8JaSw6JhQJu583E4YsJWiEGasBVhLEszzp
PydoW9Fbipxa8wxEHGhlSNgUl3w85C6VQ6P3ZhhnE5tgTnn+NtzCg1x1+u8bhstL
82gYHTJLrFwlXTglza1EGKJdgT9rtfBLNqB6fEmWTlQ8wx3aluiBVEKLW8L5nq0x
alLOGzCXQaA0ELN31ecr4wYkXsTgiQC0Nk0uAqoTImgwSmEe7GPUOatR6kCi1Eyy
4bpSMNAQQqgxDDtAY6PbRk3BNi074TBmUS4QXzEbR/2SGsLXa9aDtfrmh99GADdk
0pXGwLGD60TmYTTKk42sOy9q9qsKQsRfyWBDa7Az1dEN8qSSAAdgNscljxpVbbUl
IckYP01DE0E8DkyMRc5vxzJlkfwHygnAErTi7q0fs3ddv7RrpN49jwAtA4raRF4F
ec5yX1m2oN3PxF64h6vzYOgTZ4lX17WkaEdhcDY6FoGc6ypNzB6UAfPgfEonO1nP
4fGUlcPjYT3qT3XySSK5VfNutvyGWUlScDSVlMkNJym1M+7oD549ZwW/5jCGQkJk
gGnB30a8jSbcyW1zngoaNYsB+vFsGdUauAQcSWxkWfU1cFMkYP2K25nnRJQHZXir
2qNScjKVd4PhWA3cJ9jD298ZKpXoMVcg6wJkdLYfAfaIwFPmOh2UVpAzFsxabpzQ
AkfnofjSXyTPb2Wp5zN6LEgAYwz6zs76OdxZoKJ+PyvLzV7kjjRiQYRr3myD8qdR
dgBHA2COWSCJbGbVWoP0pXomIQwuyUTkMDGJI3GjBoGssQNiLqwoAt3akesW4c8v
sGs350OmEfH776S+zjFc2gUt63Q6x4pMYJcdOdZ3O2E7zzocy6NZIZQ1nZvj5f1m
h2wSFtmyecUNUYOnmhjhAiXjYpNdx36fVwDaxUM3KzF3dt5ytzzwekmqYNlTD+4S
xpnHRk8+h6dX7pKmJ7krtwXKiO44FMdkbcTjOjoNAGsxJinbNUW0Jdc9Bf1sotVj
YMctCSKyHQcIY+B8RLvamOocApOUOjyQ1tBWzjrV0xOO9I5Owypfh9tHkmd16Bos
xTHXKBCfEzSAZSe2EFL1MQkKqzpD4KNSWV96rQfwy114WvlbymPmINh1fuLtK8BY
HprMoQkrG5X0+dBnFJFdkFtS4k1f+/+93jDXhM/SlOP0g8lkRufEZ7qw/1vhi0uK
bUt0hxiKelfLh5K7uKTCHalw6v1dglXxkK8EXrOXvJfL08ZDAZPy0qvSHvA/Wkv6
2nmiLDw62n/zU/VT1zbeKWljI0z8li73AVmkJV4dkpJJE8ekvVKscymnuIYm1waH
jdXbP4TEyYkxYunI1Wm6kuiPj3TXb+NCeqQqtUdVJC/ydhX3PGAP9bGW+RpJbbdk
b21osunCUDgvXJ3sBjw8myPlrBCWnt3P0WtWyOFrOD5U1Z8Ct+6VtL34qorCRDQk
Sf+ykYNA935N2f3GkuT5qFvgBoeMz861SlXsvH/CNteuhc6rp+43AQBl0QuOGA9c
pAQAE+ANHyPufuX4T6+9foQSGXN/hq7KPLhgpQwiChrku6eE/vzoYiDcNrYeuzeT
Hv5N0G/nX5GkwbFLkOrs2zyBZd/X0K3jn1NLUqxjAefxKuLEPwbnNrcMa3gaZzIg
UAAO8ef5wKXhNAodS+K/H8n6E4h5YpzZ7UlbViv2gA69GS3uHIN4mbFOCCadHQz7
bJYsVysI3TEb48iOowf8SWjDl/fuTYl2f7ngwY2Lu4CVuoxKK26exfQbGbjO2In9
JzGOPan8zhOxdncLffzOHj2iV8m5x6rqtetCxxXm0+9TorUmLi9NdRk148Fc3msF
dhLcuXrIts92qyB0fZTZz/enp1qpj2OdN8qN4/Bt0YZUN5/Q/WKY4TU2aT5FJFY/
e6PJ9cH+98ABOu3nNb4KbRrzcX1pN7ZfGkYCJ4xQeHaQw4zJntFCQnfB6G1zvy+z
vC7nCv973XNJJI9h9qsl3E5rmDST1rERnpikqK6S+AL2WQ+l7M1rzFOIKtVl9cAD
sgHeALoR9Ob6enuTXRLJHDwZXwM1hk7KMMbKL2prFSd/QjfTUf0+fJ/hGXiZyret
dmeRLFnSD9mu388ci3jYj/rgmnNNhnYkr+UbtWtcoUbA8O139aKIwu5k2b0EAxOX
EYMINboMs07Jjja4u1/IvWjXag1iwrLJx85ZwgCL47C6Nqo8DezrQsohl+Pw5Nxm
6UQf4bLgu8PXNzwvGYtBUSG0wQ3PpfpVvBNbhcYYxysvrX49GHZ0wmavksvlbzAy
itD5jq8cPwz2ojzms3eVOJj0KLUawEmk/stFalKR6ssTJwkAidliBxdHXS+p8Elj
21HZ5VjuPnm0munWzipXbsmMIQ5ownTP6RLo/YCz+ByWEu3Rqx8yUfH5gGJ1R2P7
lQoK1m2CPBNKt7+hx0k/WDD6W39dCewala35s5vj09wxt/XtFRP+HrOB7Yyorojf
dB3JLDQu5Z0z62+Y8yEP6HlYGL1+oIdNJZQM+EhSYCBI+0P+hNd7RzC37KEGkRGW
9v0+iZ1GwYFEZWoTUEnTBCnIaxwWf6dvq3E58zgMT1033WZbVoODUVDDf2+MtDR2
0n9S4CWRzWukrP7wBXkxlLxmn7JFrf0VbpSzc5+9+EcBwrTuhxofj/cDC42OpfFp
0GgP3XqGqjk2gAl/VaEiBJIK+OPuadjy1GoCihN2i7MrFLa+wEnRnynqQfio41G4
6wktQiVi4lxhKM6QC23m4T530ag4Rq5fyOuAUzTImd5NJCo89BwJX0I5ZgDKfZKf
T7/EaJYxLwKtVhZZxv2+DCc1j3htQ0XlM4A55a8dd/KTR97C3TxGhnoRBCvAKp92
75a1fZLm0rhnUfnHUG2LXsXPUvVo8LaHKgude3uBThynWgop3/Zm2doPuepljvcV
Wc+hlL9Aue4PM2BLvt0FBdIIVRIcZZLQ92RrLDKKTUwFerkljVFvSwtmRwt7Xt7+
pS+tT0yGI9llqEequ0mKZ8w1mfzGPhYLkuYWOCxLvcukQ/gcixhZ5PTM5ZeaUd5+
e71XzKNBsa3Js9jvCqm9QpNR1p0DZ+MyaZp23TDVMbxADocRdxmzPpX8pdRS5/pY
tkwCNF2U0Xd05BrMEHRUJrL7/UH6uuTuCo2duLl0oK+iHH3BqFzOHW7Ql+U/xGQq
QpxjRa82nZNJwc5tAEZxbKwF+wxKdpUzIv1w5jdvUL95V5o9uUaWW0KwtFZCZB9s
ZMqVElDi34N2OFtseD63L8drJeTglsWLImLnYJoyFPqUJ28eWtmB2QbhkmpZ1y0E
ajKzUjdxiH0CdXUcAw/O8X8qqtVWRfDxD4N3bSTCX4fDR+9YBO0jJzVgrDXaaDo7
qy5ufN5UfblX+WW3oabhdwBCKdnDGiuD6zc5yl4JgZgKwv2lRukTWcWnYsJQ3Yur
AN2dciimkoWcnw9Ol6IZcHmN/GK1faph2ryYo4yRKGbuR2g5JxhXE4Z8D+jbmbSi
N4QnFiqGNKui01qIPFZVh4RsAd8ZAsKYK/5ITMnteDKKPEyEZlSx4l3tU2nmNI65
m2GyBtujxZKebzG/mcMawuSmqngUmzHClmqJn3CbSRAPNGQd51l+stYhtGosNr6G
4cISI97pS8MQ2+b8Iv0zNfVUVYftTWp1B49iLqnfHCYCfkRmk17OFMhzLFHVR382
8nPcstpuGh/MhelINURkbOyl5Ug6v6bm6C8M+MqwznkvmywVnDWEaPeahkMzBpxj
BtSgMhMyanykU47TxrZGwaTdLOF9rvuGGauEMdh95kT8phM8Hy5TjDbddlfU1psR
kZ+EyErPW4KzxCdJcgF9HhFlMQOlhDwFCoQc7vlLRkklStghytlTkwKng+LIeLtY
HgxBNw2Mt1KTHhxYPW0nV8uwUpSyxNIL55hV5oV2ufidQjtKhUzKHpo4upB2lX1p
PbwJ1aQz0j53qB1dDBWYwvsS3csb7F4CHNnpn+JD9HqbOrv2RHY4NgHY2Ods286T
332k2jrGo9bHnQwa+mQ9zoydJBsn4avG8MJPW3fSEOciFWCpXAORh6gEdlyh3YiZ
eLnqf2HNnNawijLTHTJF/4JCL7WfNkXB/DaJIJcdz21dCBOfw7ds5S6B4B37xt/e
LCen0U1kIwG+z91KGwNXqrTAJy9RkDbleSadRgpbe2QUqp7vFNxRYag63kMEhRwK
lgwg9jxFGR4nYklB+SXXo/Yc95itoDXNixaR8ofeCVXu0CFBVhsXMZ7UN/4T0UG+
4d3GbDbwmy7pWll8eYdguIa85t8/Pr4Ca5Q5nxeL5rljTvGO7zMhK6tjsLxePn2o
Wbvt2gg+IChB2XiM4q8R13wNUSKX3GaaoFqUKMguDDLq61ajZXrCu3p5pYEd/vSl
F7PrjkntWUTFfrDiN6DkJY7dhLn4tBHNX/xJOTUAa0BxNGjcU0y2DvdSr9dC/1E4
X+Xu8lJtNjrvBY2sOUBphr1fi2v0/AXVbodALkydSYjvWmlR4VFnhjB+E3a74AU0
8bJ08FyH5XteG0JkK8jkGdeW4SQ9BypJ47EyFBoYGYNruEvFm/L9d7CvYSJrt7mk
yHps9wlfhLix7EIFfMcc93CiwVlfmdhEJeTfEw7IX7IS1TLy8bsOW2EB/w2s1sJG
ZlrtRsGEFyv9IJl0pU6t7NDMrHlwHDbkX4QvEaEWUC0/NOlCHsHGMuTJzutcc2X6
KE/SfOxEvneQaPr5Pb0XVRv9hbYB5rzQnzy09TqW8WhQxsQWcwRpF84FC3rcAHGI
po81AeiCqtcND7Yf08bnMGXvAyTO+wL8ahj0Zx1Aorfx7l1359NV+Eu8oALoaheU
zrcXf6tfcNoZnsESYdMNIF4fwjD+russzKixSYI7qCC9hDwxme4FvHzxvnmjnozD
epO+5yqiqguaKZP+l27U6i44u6jZdGKR+v+SGeeA+7FV9hxvbyTdkBrXv71zJ3bH
ij66Bc+PQ7431r+B2IbUyW4GyMHWKZ7Yr5B3ZBwcLy0mq2sLs4EkklGosKXjtNYw
Vq5yuPee9LcnsXbsR4NJS3xxj+vgZYPkDctw73wgO93WSd+S1MVG0fv0Kdht+hOK
NUbIK0H616G6BC8WsIFqGe/FCr0GdL6di+xcb1vFGln2Xip9FfSGWidF7SJH28rn
3BUfs6c22fhvzWC+nDAYimIcqAtXo9NWN4KTwyO2kSx3pJfAMdUMSPcnMYbPZu2Y
F7R3iPDQfxhIdbA7fCAfa6eYqEs7eBZSUO5SmipaKiOHqN3cQOLzmB1XRQj6lJRR
+6Kp8z6jEaQlvvMEu54AzL2/5xN2NS31KiaY5wg1jxtx4EKeXUo8krW73dc9VdV1
fq0BhHcRLLzsaNmFdPscCHYa7ndo00mUtkpBxomK+Wy8wImTBt1m3KWKpPZiFz/G
KnzpPbi0vNJz7WupozzUBkLhIwecS0+3LlkRX1DQ8bywDygiNwJSgoc52iZ8Ktf/
60Bq9JJb1LAAyURBt3zdrO6y0l/kZyc5GsLZmxrwzejlUqpso7CUtfo4ZKU2bmNk
33H3W4M8GE0XC3okizPWTR1pmwx0zU6redF3oIopvFgBI+NPexQ/iCpBuSudmw9x
HlHN9XoG92oFI2vuZO3NPLYMUHj55DGErdgvyVppCtSbJV+rF9c5JQVBHQrZ1/Za
c7DTfu0NiyssrI/kgUB8vWiNyZVrgdOaKmRamRgqL35JC4BE+M00KNdjCi3yTr5b
1BvFYusrGe//blGRxIwVdGMlc4YebMyOJ7YDdn2R0296Kj/0140ae9heim9FT2Ha
U2ClzCZydXKpfPWV3ykIT8nYW2s3173IdMfG41CUgFbrXibpOrOXX0uTi5ajCqyB
rD7sdfLpRSAhVAVEhmyvpNXLG+2H9c92+ZvpQ9D6kbsRe6rubeCSvY8yatpRkV7+
EIXLGIsmvHOqd2QGB4zma4t7f/VwMUP/QsCNevfGc+MNUMi1q48NhVHSBRBQ1yu+
nWYBDRbkk+3MGS2w32MAlEa7x+3i3FuXaYBWBWLIeEeB9GraoCszDy/6AKR12CLA
HCyfQX1o1mc3Vze9WxVBHd2GTWiSzKJzfiPcbUvjNjtNn94bjonnOTlVYWUq+Ssb
ykcl+TVb3KeFjQTiT1q3LDgZ9Qksmln12X99PzgLV585MwWxPfEnZ4EnjkU3cky8
oqGwHtL3m8E6GxL+UZu1o4FyYAgld47Ld4ndhLQGhTGyb/XAT540lX6fVVB5LWRI
1eViSUC4ibZYqxQwFMy3cTD2ym+giqUqrJuvif7Pj8nceDNCCJ4tXSCrlMlmuWhn
7Th/H6tcGgZ9MeoMyMRiolk9P5tD0lwR7+ynFq/Em62TsyCBHo3aVXtcjO5OuzpU
cDAW8BsG1k0xWb7Od/Ao6rnIRuaeq23PXUDGpBBZaDGfgNyOTo1DRUGftSjInMwe
Of2etpKLEW+euhBp5z6PfmrwJLMTe+S2EGEdcEHrUIetiMICxxUNWXLKh2ZMm7l4
Gmlf6wiY+ghR9RyIZDaH4atSsRNVTMMNm/h7Z/Cv/Y4xjq40yCOdm2qr7K+eJqHU
9c8IlOY510oQ8TcCEHfeGAncbR/78vD3L1T6gflrwBYQ03lTywGUQPdZqQ1366oT
S9moOmTcGIZUkvHJIKLo6wcMAbzN18B8LDXhE1XnCTzM9H7McMfxTK0yOA54N2xG
Xqjs9MJlUj2OOShE0ZkCh31j/YHRN+l7xtpaLyzdPdwp2cbiOrH7tUsiBWwG3EXi
z4ygy8g4PhG/FPg7DjkrN8o7+pMNgoVrtULbULm6ZoXIpuPCHy2BKetPNQa9nnUi
woJHg27vl7HLVCPFBN/Q5y92Ik6viTXzvVkQXYLilp3a9RDzMvcER6EKdYVeyV+Q
DMdehSTiBqPYTZuuaI5hvBpzxq/iNHgJSRxypbQIJs8Hz/lpAuPB7wiCEeFmD/be
52yCBlWE9tInRX4eyPC4LAmNM/JqOIDiE4ztkbb81WVPl1Fu4y42w+FGAmcRsZid
8uxWMAYYUUZt1diHe7IB3PnEPrXhyq1fbPHtDfPlhqmEuEN/17hpIfvuxqoF1YNy
g9W4AvlPxvmnYjdusDjrqnxE22kah05B3qhPKBjbBW8Ao671idv1Nm3ZeutngR7J
STO2D6k2oGkQLJDkYjX2/qmhhedhFu7SSzwKn3TnylftxVk22lEwSJpNTphkdxSd
+AhpayIGvYNXJ3uCzM20Ce08/WLZQx8a9cBb+RL6ZNsa7FjbnD+/7Qi9BT95ziEf
NVv27lpTtni2prApkp+Aj9ZEagdtOtTPA9BQhTxxOHBPqsNtOrF8p6KUgjEKC5Pf
dTLUp4wM7AMthHd5XM3BBW4BZ8OToNE2cqjMjoqwHnI5QzTrP06lENwPcmL5G+ns
IRmnL1oQKMuOr3g+UqJ//JqaGHLlDkr/PLZdisTlARsBwookzYdGfiaCrqClqJmu
hU+O+rsyk23t5xCFj7obVRZKbpvW051EQEM6N4qVccOJ6xiOWBzpoSP3yCkumfhI
3mjhZo7htvQ2HbLcW/CcZT0QH1i8b/QxCzvbcJ5mDWLTLHi1J0o0ryGVXoCnYCbK
9cMak1VJ+kWHO02XVflqHflGFXBs3QCTVLKKL0oseYPG412MVrNlQr6T1D7bqhap
PiQ97glt+QoqF2/LfV2Cv9skappPHUm5Xa1VobC6k4Wpja0KrIvui/oAN+Vf/00i
gnUjkBV7NNVRcxbZ7c2nRfN1zPUkevrf3EDK85HR2AoglqL/p6oyXZtw7GwEjyIo
cBmf3QXy1ZxEo9FslD2zkENcjRAgzZJ4Qg22zo8UMoHFjs3S7k4ZIuKdiWQEFTcj
wziBerAT1PTQKGEfcnHbNSuWDTsu02wCeOq0QIpG8ApYvQPI+VHbzQ1AgFxjcI9G
uY8u4Sc1PTK6CrDdtHxFtLPQzCyUsJoKhoRqJXaxS/hsBJVXtM62gjPRi/LAfNlx
Sio8RCc9NK7wAm6ivmSUJuHbM/3S88l4mnMotuvb0QbPIUjmPMMrH2TLORJ6yzqc
mLDc8bB9LU8ZuRDkemgMTLxSgrzSl25gf0S4EBGR+2gTfFgSp/C5gipAMn/F01rI
Gtt39itaFUMZVkQ6CwfkN7/35yx5pu4nwALWXD643oR7j/uUTrGWbH9nodUwbUY1
m7BDeD/gTOieAkG+oHz7BKj/rEe3/YYNu7CeERcHcsOjNy4Ga3rk9VGtpB7DDd8e
A2yDj0RR5TY7YL8V62joayeHR2itdr0c7u9MG27TfTANyxg2kqJeVpR8UPXjDKlb
td5rQhcnOMjGhVhoxeTvgHavsfFM1ESSIXmAbcXyjvQnqJYNEZyvwTj4FuHM+rP0
jDpWDeopp2AIgBADOKZrzemWpENojV2F8wWFDQTnaojyN+zoVblCskcGJDeekHMt
QhAkN06FVGh+bMGB9BFLhvYonnTPNbSPu0sM2OTcJ+CR+ArMkmPJFJgMkop/swhF
1nnpQViuT4pShra5bJ0y3ahKTNL//rBryYrLCv9L1bB9zKvrYmqYGHYbKIkXA+QE
8r0hi3JCRtPq64yewvDentnt3lEQHjFVrsnMfgrYj6bOBnAUyH2sqQzq8SPeZoGY
J2oo6ydVk6IBQKscDtsdKhItgmIr7xszLYGfdS1YRgAO6U5ZcPt9XoTSBAUz1PpH
puRf5QgGZwnVryPHQnXqcbMVU0E4V+9ebi14i2Q1YqcvuHT2rDIrsKznsFkhHcMF
9ZJ1HhUpbthKByiuut8biYSjdxb3mulVvaJgfHMxn1pEACTFt6vilTfkALQietEi
pwS0IcisWUymn8GuHFGKDLQ4749c7kHoAVrLU82DYdP6WGGlx0a8A9MuOk7OuqU4
H9UP5BojwQ/b2TxC/Cwe70IaWo9XKT3mrz/b4AeFMjUZCWJ2IvcdaAYII6cnsg1b
SsyymKrRjsEL5QBjCMD7cPqLgugUlMC9+pgNdYWBp7ZOO2lTVYec5OWbhsL+kxAd
9zn41NRNdjt7m4GT46GPu0bPedviZQAJqTKX4OY5AYkMaSgM4hEFBpBgfnUCHrYc
ifQ9Wnz49olONc/w1Q8oGJmOO2IQNSycw3cRmD4rlc07wBqxvu89/hESxRGu+Lf7
fX/HwLlVpCBXxM9zIzQi80zEy/2YGyXRJJR7eLbFkjbfaU3MTeNTcedoOjHAbb/s
9+RwFwAALN4B9lxZOEXNDabrPupiWDcnEF9e64VlpExn/6mGXS7JIuHJYl2CLoMy
wpYH6al9RLBWDBgO/+3DYNVQ2KkTaFewlAFX9IlSNhAeOTLQQ/9FCaDUFg9Toe7O
7DgYvM5VSfH2svb5AS08C0oSc0EyO+ufI9LFCdmGF1svRPy4LfK7iVWdnhFwNowN
hmNVE7266PU3yerdQvY1fxge4rooFSMoteVx0SOSpiPhGPszY8C+IdXyZl4PdA2M
H7u+1zWZiN1zcQXsZR88SC9r2sJJlnYFtPxYqYpvtv67WKDUPFaugO55qvbS2j1k
nWZzNre93I3becpi6t1uAN60rfs4T5QGuU8/RV2aEL1Ui2skbWQDBwqUMjR95J7b
M0dD7XblKcdkttG/X5iGds7HpTgR4q8sYBzWHWCdqljS5FCR+JtFNfoALiLkcYL/
ODnAAKcC4Ebds2jElDwoDq3P6xet7SQVWSv2vJtAla3DBSLQbiq4RPB4UcgWNSSF
qoArr/B63MrHhYGSXTFzCJAy25xYoYj02g+MLBd0xy3eiX+SMTFSmF7tZeHQ7IjL
Bug/6YMhNQ+7zPXXu9GqmVuVDoLl8IedWI0p/TEzcBPtuPVwxFveY3phOin55ayo
aGTg6rVuz9zVbIXCWSCsRGG2J2iwrPVRcopS9IQ6mAqbrIucNU/acSXdOkckKHZj
alHUQFV9V7+E6YPBAw/VbhJUxpVudkwX58wi4VDtuZxzrfSh6QyCjGwwJUBFLVtS
jDtveAk5+YF9sN9PezTR+JKHlWfVhUVUQgX0qSQERAu+UDrKGlJvqKxa4XNlEooJ
eAb+PCK8fZ8v6JHhi3Fc+3nlFrHt28WwtOZPrvcygBHVX47wgljAR7mPLF9RBzH6
20UyGc8Dzq+B1EvNIPDB10rEoUpyRm+HU+AETGU4Ec9ShFPRHKBtVLUeNwUEW/gF
3V497lIJsS/WjPH4zzB05I8azs2eegVwOhq3wehdZ6RIohOpgmWLXsghAT6zX/6V
cUCheV11E9ZKu60o1pTnoN4rfhgmWiZswgy7X61PsP3ded1WWErfbp7ttkX2OF4M
I8NziDX75io0TEocHGQTuq3FxQZBUv8dYGgNBIooSo3mUgamCGh2p/vosS3gxLWw
w3SK8qHZNxyaY5pRq6Er4VFXcydMOj2cQQOsFX4uzvoW2H/6WCw4tgNzwf/jxLMI
H0utY/IB55/NsxQho/7uThQ60x2NHYnHAeDhJ/x3f9YLAqAwXGhOsDILubWhQYiU
JWMakYVNG61kgdqPZYdT5KXmSQN58X+a5KJlqIfN6oY9knT6VC0SBI0GiiDt0ILK
syPP0B8pNXghloBa+qu1iB2LwtCA9HE0Ds7h919lk6dvJb/qcip8MKfeLxrdNVgg
FACB+UMo/HsshjaidyH1UT+j1Am/rptcM9l8/9AJh5XJeOAJb4QmtKJhNisUymcd
r6GM/uVUW1lxYYT/2KFr5cntB46EC4hYqpfT6hKIVgEixRCvm6k4x6ZjINmD9qZK
dMXj2QR0ZTgtxS9X4VWxDAfWmCoPMYYHwnuQ4cgmb49tXStzfodBlTWFnpT8Ojs8
VsMtqhTMt2lhzm/dxqkDigf+pZVTsn/k8aHaF4dyHWMPmGbKjEIMs41C0MaHw//v
MgVZemq943lLgihFzFdoS98DISlek3zCj2qIqidFaD4I7Zh052S9Q+VJchK/vxjZ
sKf9q+Lu04uSOJTvdn3ie37BGN0IZtfhScJOapIBY58RbDeTneSa1wHzgzRMkBya
Wu/q3G+bJUBLAdnzBWWxPQ19eVx1010Wb8baTSjQaFxvZ8l6/GMXR2HwLDj/fk39
5JRlQAptBQbLwu8E7z6W7UBQg1QVZev8xWsM91X7uFD0mmSMG8iOvlvDixMw5Cnc
GfVYFqfWnXj1cdClt5rwJkpHvwxcnjDRdVl+uOLeo5Lpaz4u6nzd3kNkpOI6ADcy
eOhyVmSNfjcq5OsZrDXAH688zShmYiB4bUcfFB0Lz0/44bVJbsYHpOf7311jbf/P
q84Dd6Qr4m7PMOba8e3PROkaqcVQpj/lRD4DWRjXk7+E8FWVJdE1aim/p8F/LlB8
m806Ti4LpmTiCppkBuoujjJTsmSYvjnC/LMzKIFh8Wl8XHNY+pNZBzb+XCN+msqi
uJl9ZGV8+vsJ1IdRPugERwoU3pQQW1fJCLYnO40E9i3dlW8HE7pRgNp0RjoVoWyd
pq2WG1LpkDflAQidyMOv5/V60pt8Z7a45fBB6RtDn6Z0oN1UEf3E/DEGbCxsrRZc
IcgRhjwD4OLorX/DtWfCDiQA+3xlfmyumE3JxYJwFilf3hmGm9RtEDIrhMCKz8KX
2taONW2V/J3OPLtzZYdj/ugl/leG1gORSv24cIjo3Z4qlyigu6HpKA1HKcmRYT4g
3DzV+EuA3mYOPA1iyYwUM9dR+QBH8B9fXQ4AsYlZYSAuNFQFhVzXQOoO8ZnSDNLJ
tti36A9yUUbhdAqlkeXbPHA4pDVLsm+jUDSvUXfNmbYc55SwHPgKXFWugSDTSjuK
JcjkE5MTrEBM15ediOMRqE+4G9swcVLwSIBhvCPlzrZfZi+zPb0+uhpJ/aZmqzp8
fq3YkEz69k3hSC+hYWD6ubTQZmGcknj2m1xe7sMe/VPiL8jVK00HfrGTlYbUbhcf
Kxb8ldyJUTEyam96uFhKoQusGV9ebQRBChr7sBEcyy4DzIG+JVLuI/N2HPOoAg9e
OHyivRagAyiD0RfVXayp6zfwkNmFNLIeb1eYBxnDjSsn7kjA24s92ZylO0injNlI
0hCoBuNM5Zk10jzSZQ5d101qX0sMnk2MtYM0gmatsVyKNL3/QmjVKxKhYcEJfmn6
ER+iH373u9e8EiZszm77X9jVzhGOvvYRFMLKZIMe2q4FeTaM2QB+0OwZ4BEN7RID
F/i7kfIZixitxN7zvcGY2RBeP+dP9FGz+UIWqsCx6KItr5zuYDkTJMk+fWSS9qlo
Y9GV8Q1b5JGhQZktVc2FZmEGkK8zOHzQbKNm72Ukau3jzBf8HGUP+nuklTuYMg99
9LbsOdLjX0qPRchHKEisBvFCUyAh+LXxJu068npSvErM3pRFsx3fBb9PbKTzp6bs
AytK+4CtqYfMwiQt0CAePlx27tuLQFd0if5xA4BxMqMzQbRRnyZMVQeERbJ8Ourq
Z5Bxiv9pTQQJGI9mul6LydsQEgFMM/ngMvptfXJLXBRgMW0wQh+kHxjOPy6HpgjV
RhxZGn0Np+M9ICYNLKIqsF/cAp2JA9D3MIJ7KAgxRPH6EI/8SqLGNXzMkf1paYxa
8NaCp2JRWQ9oEpRx8qNxT+WuZ6ljLjjtKzxB7VouHTHAkhM/51h32nPEz0s34DgS
GAYexr/XSg5aGlkB6oxsq0p8vIC5w68XS+wtMRCmmd+tGQB178Sas9zzun5jTu46
d7qOrYbZLlb+J39cp7+bkqk/UUYae/a+m5Ex/0XoaTN5iXmrwdyjuH3LYVCzT5bF
lRPEMHlgUlD90vZXixWZ8/RBK9x7IFbP5Baerc9ooreGfARS6Gxr3PKE7iNo40Tx
8/qag6Hl7l0ytFQh2f5mmro5MLIdDs0VIxOPs5Wrc8sxNCh7S/HCurv6dnVQl1bN
m550SDaYEB5eX2Ogi3aU2b0kh9H+G8YfVdzRBNHFyHCarh9r2TkCb3BO1wEoy3/4
zllKii+tcCs3bchst7IjRbesafUDLlnAtb/DBpd5QGJUuq3x+60fn8K+ISBrYUxq
1qZ26AK3ElkkH8Kpg05pQBiTTydZST2sxgYitfh1B1c5PaqegeRlfCDmk6Zlcta6
5Mq+dUKpr7fE+dz0qWqlIpc1uuJi/RdEv+5mMRctPTrX5/Ld0Od/PP77oJWC9VIn
FkhC5WQokYMSqto19W1c9UQMHhXepZ7IlqaLDx/fyZl3nk0GtJLb/AqA/NPDp022
Yh/RFnMNw3ZgCh/RFpOFlCQ6R7PKC7iIs220aDrALfTUXm+AmAUGNbl+ymbo+833
EC9xTxpxetpPazIIOAcI9U1ZqNp3u1BFXr/YOOyvaptJPMQHv9u0CO4Bdxw/Ajys
a0f1kbcIcgrIJEOqZZnM9HCK+1V6+MjION85tXoBwZejzoA75Hut7UJD7axaovX9
qjCpPcSuVJkiTXsHr0PBsrkdUvHFxT+luieKuDRKURGnHsId5VNpUI93hJSYTaQn
9IX3nW7qdI4VpxeZzbeYTF3P3eUzcsdYNO1qXUMS1qDVNaRS6y6sq7/sl1rjMNC0
ftEVH+xDybxnUIcitSGEu/UFiYjm3YYNlJjd/bKT5b2NaA0qxPYYpRKregcvP9FY
cX9INgxp+MNRx7LG1Pt1WYc7O0AKNZ3osP9VBaqgsCQP9CEsYXjhYUO71HNWpSGz
XGQc7quC/TcOphiv/2erqKuCtTEfMayKzK5BGZ9qXnmromoR0jygf7jEoHegc2Yd
DCaT/nyE79oncPjmLFOCamtwtEKrqM7pFMp1rw7ARrPl/o5qxtxriDU6Ai5g7USg
bW5wHlSTUjlt/QCmSiRnyF2hyVC0T0ZtpC33Vre07879Bdb88AGnHD3LWS9SPCdN
3ONKPIEoN1uI0d6dyF0g+RiLf3pYH6zDD7RwMDGU4eoTxsb3vqR7LPaH8kXQIIPm
o8GsJa0fJtXM3BIdmpbTpzg24SpSrJEoan6rjwBjPgsMZXJsOTQJk5pPTpk1RxtN
lPbJkCaSrk9NKmu5H9cGupoVOOFYZtJ93i968KabIUTzYLZfIk1t3+X4mZdHUW1C
uD7yljJAyEWgeaUq7z0uWaiizaO4lLeT4CGo0Rk6E8i8L2O4zDvo8CA3brl5jwNG
HygYB6hBdbYaIOdvdH1WgdP7R3AJFRlZcLpjRwp0olYo8pJyNkpVnmweWZyvsF5b
7Q0NRNhgZ5n9t0D9bKZ8b4Kqeh9h7UfrXDGIuQtyV0OVvWCUBGVmCMSghZu3nnPb
J0vu6jhyYeQ5G7mSjxkaUYbrQYfHqu9izc1jC2O8wbyX6V9Lce5oLRbTmBeIligt
jZNJ7w3+ZHPSGlnR9Mb0dDDTwSgrMfZXT3Vi4nn+BYjOJ3i5We20F8WEBg1SYm9H
vjhnUxmB2H+HNwLciezb7o9rufGBnPgAPElU+lr1oA+2mMREXXuwdemAsCQOZdJN
VRDZLb9g0uTC75jaJC9Bn5zjwavKyFEFKMig0MGhnGRcT3iSnLo0tIljX4jM7Zmr
ff+3YEpw5QLTK9zRBACWbNFH/3q9RtWMaGVBN6A+AP6RuFjnyIxQIYqTDS01v3Gu
xBUj47cagsHoOmzpMxIR5tdFWlEdKs1SbOH/WIiJJseZW2nmMq1Ut2UqcA4RwLKr
wkl5jNo1OuH+FMO1MxATHurtmbSvcolyhMsaQPrWs3zk7gfEY6ylgXpAPdSn83aq
C0vuzGlti1wx9t0t6hojbiZs/qdb9JzH7NXZ0gw9y0MrhjrmJLT5QAYx6G/AJNQ2
osOvyaIoMHyCU3eK9YyWiuiqNP43f97r8ESQgxqz5UQmI8LBG0vKI+9AIqwySUhp
nxeUQyJEcpky6cVRC1TPEXKbiXpYm6k8cc6IkNxlPmOX7nr11DlgYORofXRGreoW
uOQ/FItCD+S5V+z+GGgFvxPjKrgvEmQRIhrAaOUJIlxuopQALEFPmzQg1HLiPdPP
ukdRQIRpCUGhAeUmK0zItnS9/47HXyJs6jDL4tEgmlHRUFahXmRVCkpw1Z88ThUF
xeSR7jxric18HRo02+eJejqsJkzRkb/pJHHoal8pxjsVIxGLX8dJ0mPJ8Ws/g0no
iAJdCB37RYkurRrEaVtcm/XuX6oJBE1s1reU9cATr1T9bjvUVxNqEhyGTcehUfFg
BsQIiS//qfKK2TQZAs88ETabflPvMwTQyfT4bWGuEP24zgWQhsy45ZIYaIy6Ctyj
phj+c+UbdCDBGte+11rCrcynK67vPvNS0rNJP/UXdp4pNPlRa/Zggih1SgIf03uF
ILdFeXxtqdnx0CSZpkiWxJRc9aOvt5oCnflALSdeGrsEq/hiefh8xnIIFnNhueX0
TmLoSoztO41hBICGnhuD+81OJFXzv70lJWpra/TqTc78jrmYHEc4TgJfSFekNtxR
L87pxPgHESjfLIfZtNgtpVv7itr3TJM81GErtD6/u1LX8xeSOovcbbWaJtB/w6MR
cA9FtE3R4kAuCAF3VSeSIcXy6ZDBaOpDL3B7uf7A5NOWeySfFbgMgUYSW4x4InLr
a98woGXyDFA1qmXW0LJrXzxvb+dHBSgnSk/sTdUcL+SC7hj7tKbzwhsiH2/yYv6X
OSbyNZuJ2CvWLcd9z4XAwf+lSOYTnM/kRmQinT54G6ijYGxFIZTyax7bIq2k5cJu
MRnWodg3qH57cwL+k82sZOyEZqzFu3n8Kd7A5N8YNAvaXcsJW55sZJnnn8s1d8uF
6zjvjHc9FtVYqeEEFdC2krOsnqd6jaBOh0+M8KlgsN2Dids+zY53nZoaPrfnssGv
ACuNSy2PELNDJD3NIrDlyOHex1w/LBpaguSmDfIipowl4MCeXQBcbekSuUeHCIAa
gaUBlJn0ESutv18GNgyqnfU1KoWH2dOHPJsHTih6Hwugmbj4kGALHkXRegYliKY5
FvCv0yiYDYoudpU8VNHm02GtdfeIooAvk7amg11e1dLq4q3UySVt1Q4Yg0CJhutN
jYhRUMbVuKsZWZEQR38CJsGrtrW/zpEuog7HF37K8+arb8/tlOJ6G41W8xscSRZ2
uyg/ZcvIxuUewVJOfzk+T0CjjP+JMFrxfqyyvvVVf1/KJQiT5CFMuwitIm+k5RPh
gVcXaGw9B4Acv4uFmYDOVy8Lw4g/vDaNYb7cSyhMFDMu20rhty9ADWhAEL0Gzh9H
VvUD72bXWdf5k/vLSEkBpXiFvCoHkVR3SX2JYLOQ2iAS8uFvckMpN7vApSLF121E
YyQSZFFshmCwoHO3UkWBImnIRXzjBpimkJd18zi5c4Q3aIW74pLo6cWyfseSxe/h
pkmvT6HPWjY5rlD+P+HAEwoyZV2yL+v/i20ug8XHjWj5TJbQ8vtVB/EnqjyHdSje
s6zC0AOl6ja6TJdLtn8/XJyGz0zB8QN+boHpoOv9au1tcMMh6rRx0E1tEZnqErmg
enkdOyAckIl6C+HgjblYYM9A1NG8Bq1qar3K43Cctvb/8+PdZiCbCqAxOZgQqrRP
+Lpaia5gEc7E8m0ONZyCtEEJ6uFNlqWllDVwykfnvqaInKZEQsACIj77SrA1oBJj
/jzE5HGs/FfSVNVmFDUo+a7sJN3PpABVsdfv1xfSB5kTjz7H+o7VPB+xlNGxHWgj
9uwlM2bC8Bd30hcbmCeRtd91kTO5GjRzrIzWoBSbrIc58zmsbiwHlSAsx5A+uCWD
sbcC+3n0T1XpVTnj5QeU2fQB/JoY0dyLKu7FClwG2QQF0grsqQDTbSlsCK/xRCRt
FVLY+LIYuhzUBRM6PuumUCIng9LG/llJhWJs/iTFP/a2sxRo+bY/NM1CjDZeIW0+
LVafrKjil3O8DZylWiXKdOATiJoYKGjKn90txKH0gsm/4oX9amD5N4BFgoMRxmos
IFZmj5EFElIBHRL39uqMgIQrefccfXxwV7/1mS7dp9UbEys+umxZVRx9yX+rdMYf
7feiy4M/iYdV8QHuy6ZSicdWtJLxUwfIq8JYoENMNVh+fVv/oro/cbb+8+6M/9zi
b5ChlvJEYRI1ADtCuYAcMHcbaN6XuiuSJLJTrF3wklXddF8RnL3PElKKbpHWpS41
Xbe8pgXqIGovXsnnSPjJ1I8K2galImSFZ5N9ZJJaV0nacy7aJqEwC/e4dWFzp1TW
duhc3RVdd4lZg6EqpD1grXHGiNcgn6JDUHrlckfdd0RzDEIh/RGrNZuoW3iKp8a9
12/LVSARouorbYLG22guljoB04/P06Lfef/RSRJ66TJvmqIw1UZcWg9GTYFLFWgc
s9V5WkVDjA6+0Qp8WewRji+tf0TuPn/zuinm/xGjWoA2g5XJ3e4uaKU8iIyegQdR
dh5//toRc3Z1G1zKScrHsmH3ZoixrEG6Tu1RCo85locr2m5mptIeoDp8LpkjM2Cx
8WnKQnIcnUk6bMhDFoUViSVt552yyt1y8u/04S+3/VDetXGQvkTWklf/yIavsW0T
RRw/It7Gu0mz3ki7+PbUEP1lmvE+8jjo0l4d5zzZkNKM14VhYQupTjcqQo12SNrO
NDOz/Wv1CJdRPB3W5B2YOx2nhxxqtRIEpVvaDm3jon+s4YFBUZHjY7DhuvNEMVOn
NuYlS8FLY+UyxkPZtfsPqBM4bBTu5mzCsk7KiWoGNFcdNGsBqzjxkg9pJa3T98y8
3vthMQwdZ1or8OQqMX74A04WuNHDPw0XPrh6iWO7ZJ3BmiUVyFYWkmQ+n8F9FBuf
FWX/cdz6p+EFWowBeI4UZOzVNTcqB9nlV6IvgJsd4+40njp42c+ZzcFr1B0RFzxH
m+OvTI3qdVLZoslymVtEttYXlxQMXT5lLwE2P4Is+BLCdK0K8kCYUKC3UT7xBMaI
qvCBcT7VQzKhcx70vC0IgDwBA6SLR8wFJ0a2hU19QZ0DfNRNaxssNlsOTdP/oh7s
sYK6FoC4wY6VHiM+wgYEx1cx1yxQMEAYP6x9bZdQEOcOelv2nyaF9PaBXkFJY2n8
J5baYoohSaSdqKOx0bU5IbRqJYjdyyAcLSx/aKpOtpMObkriizJ2DY0b3qvJ586F
1R6ZdUOZTEN2xCUrFs5EL6L4gKgRUoAqVs8DScCPIzo4jsFjIeob8PdeJU7LeALa
wA+9fMOKBiSlYbYRR0ytfRqffRZocOr7iZWVYfpxPIN5fcj0q+3m2H69Fb6XuTxs
nyb9AJSFcTsfCBJr0YIjvQEvT3jztp1cNP3DGxhzNac5VX96OJu2JKooQ2ACguRm
pgH+BS52aE8/2Su1nDfJMikfY44bVpKdUkVAOOzkcnxMhc+/uZQs7Fvc51nizySS
W3PL3qASt4Kol7YFFxGy0grtosrJIthen8PmLljYuVMCclj69DsSTlEbHQ02bjYO
T8tRx5hCbxuHuyZzg8lN0Wz4oT5ZakrHpoV5mwUnCdrpdcy0YE8SS801506a+NfZ
wygK0sa4Lv8WOZdH+JqAqJfwP5vM5fuAMh349ZpyGOmUn2zUyqmBn620kDFaBe/7
0SfCA4CviGiiqE8ZhZ4JFhJ/7KfCDuH7WWcI4jrcWWugB5wd4qken883L14aKTIT
7HkiLItjhzdFQCBbevzmH1hYid0putD0EFOwskDQMkOGxNfbEyrLGiiHv7jaD05p
J/wlq4uMGcqd5lA8LPofO+zgMclg2mbXDk4iP71qa9PK+CEsgUA84ii6TYyOveBM
NWtO1utAfxvJsD0C9o0XdXZJbnLjrIkrxnTjIllHlXCnTGQs/ap7cbTukasvbnYJ
OqNWzGuzxSRE0vSolzM0gvWmHC0ZZIvyBmkGrX1TcJ597UWK1nuY9hD1E26frwV1
fBwV+z2PGhc29SVjFhDSrpEu9ls7e7Ii7H4TzOIlvyGyJWkCvnl95gwzO03wyVQ1
OToQxzc45EU0KH0YDbw4TLqilJ+2JCGRuZbM4ly40P9CK8bXe6FRjunRsXQk4AZr
55gA03hGsk6HWzwwYBexQBZ2fE2en48j0Yal/DwRdZB4dXk0IVe6Ozo0faqSQAsz
Ex0uGLnS/+J3zaR9YQocfqA0wvoB5EIqe8TuFfWNgg2zlohUf3JirCB7HDbm5dEt
73KfhO54snUC8+8CSXafimZUDSSEfkE9NFVB4lQtT/PrTjXrj0r67RaIrqUV4sDV
ZI/bcwEpZQkr/IpGiqbXuXLhDy6nPt+1wRqFz0oWp43QoIzUJkuWMBnncJVwq6nj
eoVeCDyCKzpDvuTkMxwZbdE+4ent7EDWrWVAzIf4w34wlWC6zWnfMKzY0iaOFpr+
K3alZfeEKgjWuGXrVhirV1Dq9xO38WdlKr+3KNale2lGWuQJV/Bcqxq/zDm5tmym
gFsWRio+ITsNT+KYePV2krgzs7aG0ac+HgiL07m4Ny3eJvJaPukxYN8lig96eU6N
MyTgph7aJh5h4cKpUSOheBukprklZ4RqtRLtoSUERNu4RcfNfTvjdpo2uHe9D3ll
2Aih5nxRUHnbTvjVSV/8whNacFACB6sJugtjJJOYoh7AjyOUZjUP3YmWinxHct4J
GQQdzfS9gT6pzEfqoi7XsTGVwM3lRDvMs5esDzG1O/teERqBdLbN9bQlzhxPlN+F
ZO0haOCJlmqD1HmeSZwa0lF7VPV6nSsHvHl+NmcFGYPlL3PFGfftxLUB3KrZkH7E
t6RjTofUrIeJ+kFJZwBee4cgc4eITY22fbMrGmF/Nd1pGP58I+mVXMaZ/eSW6E2n
NWAVZKrbem6plMjbYZmzSxNkMolAucPrRImZiMP97tI/D/YSZbK9tUQwU5A9Zudp
mAzjlzEqbNUsc9sHmKIlQpydi/ysD5A7+53ZAhQADvAnZ10drSLWa958Bzwlsepw
2otO+Rcw327plEkO6bJUQG3MV9A7NRwQVr9whsYq3jUlVFM04Ic/OLnIzHmGRdca
yrtUwxVtnHlH+B2obV0FnbZMbM3o/iT4Gk+mUAzz4tq4hr5ct7mXOMCrrzR+Swsg
y3OPwwccbwcB0pfmM4ZGqGZi6hYJVsJENXHXHB7hl0uJhaSFoxkoLkrOfWZQ6SQN
TtppN4i8dacChMUyarUXhCQy1nBMSUiFEfTGHneuJ2Zl/PsTFelkQrVtfHF1pu8i
NxZRCq3ASXwataimNuPa79BBMAGVZXcx9SEY6Co07H3p/K/TCnUoDieWZbFw03ik
A0wEN8BBqpYEw9T8cFNIKSO/tDmu+ezcdxIIvE/Ev0IQZrcu3EZlz7y1TiQi7faL
IxUZfniFuKUR+TJ6LFCtfIRT+gxSgv8i8FyoBMghWHRgOyvt9wYO4zazeUEyT1qW
L1+Xynu5i96UJmPzlaUTCQZ1siHs6zcui6ZDsY++05UUQ3xBiSClWLSuoZtacaik
hgFOm4G0eCbENFKah8ZIc+83dHJxQpouWCdWn/L2gN42MLHaM3P3utvXgypTCX+i
8GH/AGIRlDe3Yki1X559jlzt8mKmLPFb3MZEyMqI3ZmrKVmEbcNhM2guToSfSdy7
PtOzKFh62AurQGXCYYqtO/py36ubZElKuo6ZO7uJPy4NMdmRCkmnW7ivE70TZDoT
HptJpy+7Fr4Z9ybxaBCpGOKLYio4/5e6oROhAgPDXaR1xeG4PTLgyEbRW9QRcnNA
PV+VWVr+A9gtMZyEd04ARLyUUbzhpEDkwzQ+xV/v+QBaINX9wpkE3ThvjxZpSe8/
6KitC9lvXoT6XFWbSYiQscduOEY0Zy6xcqgtswynAwkW+WN87xYP0txYhpPJgiFO
Uwq+kKnBbSpYJYEkqsLA2rdJGDVsa9jikxJO1pSTd+hG3HtGUNRucrK1ymulwwFN
O5ov//Y9u8ZnRwRicbnEN79OL6Pxoumi+l21OcXHpwKV35y0HK2dHRFp88CTKsRx
FFWjomY48subf4kdo0/gTViYKXxmsdsXqsqoIVL7CC9gT2h2aP6ZKlqtASIsrOAU
kBLTfzu8GuRYGhc4DlLlrLsZxvAJCqDoGz2zBG8LM68myaT/wrLlyejPNUo/l4A+
6wJ76IHQtsQQGxJjhmOldsOhBmZFVEt8F7BjPmZ6BYBE8WuxzUiCBbkVfL3SrnQc
QeMbK86cK/EBdJiOKPhklTPl/J8rLAlAb0lEbPQOgTI2NF2ywIMACg8v2cKR/mp3
mp7x3wXMDXoZf7AlQB8DTcqsSNtFLQ/Tu10h3I7IF75ZWPLwBYE3dTJAL4TCYsTZ
EXvV3k3CSy0hlP5vpnteFSIHJ5Mj64Exd2Fr17dWOAIkPc1DATtR6uvgmPkdxJ1O
BB3p3QemIPsKl1NGz0zb3mYglFiXMBdqvVd6bSdbaY8UrlRZd+7zdxaLAn/9Ne+L
A9IrZrIT04Mew7bJLcVOh9MNYZrEcIntR1qEg2ppmvoR3pwQhJYtioVgYt6VnMRc
8LE/Mt4NB94nmFCWaoXfCJbxvrWsVD/p5TNcOaOzZVjHMYpQ8dHWfVuGWmCcLCRX
SvBAPFBAtUJ6G1wWc835Dfu1AERZYUsiLyeQ+B/raEkyzZFGu9tR5Qv8PIj0SnC7
uJ61VzEIZVx/obJauQAc/pR4SJtoxkDMvOAp1av0JLXoPRPmG6MXuxyphjHLb/9o
rLZaYO/9QY2zRx6HCnjAleYpu89YPL5qXdgOtLkm3gGsj+qE0AHG0iaLjdZvgfJ3
VnT06GKcKR0lDA7f12Xr01QwBS9UysAOd0L9Bkjt3t5JJUd/+/CxfaZ8F4xHtXo7
xI8OLVKMK9XnPk/RM/e1k+JdiKpB9UnNFtr6LwOVI++D4xapvVMQDwMDfVHdWQqL
Rf/eT21h+oAfRSNDiT/uS9C9wjdNCbOZOhWaEMewGZKwq3pmNjiBegPygalNjN/J
uPrethKTR5oDpDufd5puSXAWc01HPYrImzAYYb/mfY2ienXJmkB0sHe3pI7vupIB
Ydwkzzw/1s5pZLTyPXXew//hqsnFlh7WaoGjsFN10jgFIj9m59JfcdV+1lmH0hfp
FmbvONAgMMXc1TFxhzkUqBsH8VHsbrtXkl6DJXsgzs7l5Pw+7ZhxGKGJnndat78o
QWNMTMXDrD9C8dc275/IdP3yG5fRjBYll35SVOJ03EvywZpPnGTinUmciRQIEIAm
m/i5uPP47WZTjekXwmWaKwNn/e2rI4FJcLbgy7ymErAORlt+H6JLA7EIJYa0AUmM
mkpCR6IptgltiZhGRXaiXsrBJuQAjcVmhHXOQsc7kvgdNmYb4iCCpnxZD72bAze6
u0VAK1xDnsfw8p5tXJvM9abmPKckqsB26TqdA9zK8uyHlMyxl8uBkLRmfKbIgyQJ
mMErBNxknGhVQ+gRaC5JfW8aZXToFybHPqJzUUJlgjcmHNXZU+eB+G6E0vZ1wshQ
hnObAIGb077F1nVp8Cvk30j+vXe8dgz9SeDGRU6GKntQfmx/A8CHkVETgnsmMZzf
O+bNF7PtV5kBg4jKvnr0jQkbwKZs/WxlqCuF8rOYLNVNT5yNYu5Rvd7dKV32tFLJ
n44f8IoA1mJdDTHIMbuSbQQ+iPIC2B7Zd5RTir/FwPtIRaDLVRxzDkR03PHxhOyY
JVvGBVH/MZ0uy/XYsZlDHUce8CjZTh0LrnIncHXfRO672ZxT0CHmlmyY7W3rcodG
4IJLu8PJWd3WLIWRPH0UlptFdaDfkzPZ51+os1EurB3SKRTMvx8OyuPEBUKy3cfX
Hw6x9jpPYvYnasr+CkyUxhAYHI4dwDXC7YA1DT9BLZwNgtWPcoofE8rz1pnqIpG2
dBQt/N1D9sg/m13z2ARtHk5RhDrYpk/u2+rHJiNxL3ijXek91Mixc3eoPc2I/iRo
iixLvCHhHvsJdkBxxI6WmEvbaI9K6Bf1bF74U/aR12YJuqeeUOwphm+USa0jCDbb
Z4NA00Vqj5Dj5M9sgnlt2sRwthX/4JFWNXVOqsFGuZ+D7NHxHOR6MJWpRJ1lbw1w
JaOfVAHeI7l88lirqqrTHbKZMT6hh34RfToP7Xrrsa/IP0v/h7oSZ15oH/q3LT84
gJPFhv4v0laT6Sq/3eL4UQ24He9Jn1gfdwYIjDx0rVI97RzgMabfQk0srbwCer3/
X51V+zHhL+MyZJn3z8sBayNLjZLW1UqZxPBgaftpNuHuB5VzIya/IJtRAXPnfN4N
XOZBktiXtj5IuJdQ1FYoZF4QXR6j3D6X5v70i/kIqZTdAd2W8Q+45Isf/jlQuzla
VZFM8DGqCJUlvMOGV1PrABjF8dzWx48dOXUSttQFt3FsrQJRjngxev0GsZo1SWYa
lwnWogi6MgU7ZcmyJusbbl3BKPPfWvEiCgXTGDFv9cruN6y4Ebfe+TQuOa0R7ZoR
DsTp0EIS/hmbJ9i2NMT43z4DGq0OpiuL3xjvjKNsRuxKCi6QRuhxBCasqfLqrLOc
LnEqxolEvXb59DckFh0XPURYbzkXMeO9d9f0jywjhRDnakpZ/kzrQROmwBZ+Ysf1
PIIdLRPCrl96XfGeRZRmJi7qItYo2T8cuNK/FRwHxv8eT7DDV14zGYpMGYZ9t1zb
xpTJB6x4HqWVKiKvm5v1GHfDurOQ8v0dHV/Mldoh++F5zrIrMOSOhnB27/aHA0ef
zcX7hxLSvLzlOIUr8nQcEq1izTC6fFQcwuONRwiq0M0DsUjiFB1SwhD28hv16u1Y
9RB3vWw3gYOEOt1TrYEnoljPJZjQE3R0t+Rn73dg44KoRKQV5sPd6A3OMof3TbnY
BsOF0NPC418qivRNIaquyB8vtQj3+df8DnIl1KsQJtyfgS76/kqS/aWqV2lM3M4D
WpB76GsSmXqIwL56e7/VABnoR9l0odQ0pRaQvWgV5sXvA4MCCmRyuqvl5mMXmsIS
ABhZErruiR23GioJyYxUZuBkLC836w7VmZJmRGfdV+wAV9WfGhRBL1kGW9zm2/SL
pxE+cmNkTfyp7ebdjIYWDC6/rUMAtmg7Id3KVvB6ixF20akXjlurxmO3kb1/3R7q
ppjm1Bwf/Ia65efhGhy0ti/TTw+7FGf+fZkmeXv8cWq016DMn7BfwQvIFY7nZArO
PV1rgzNlmYDaOKPi3bwoNJUkZzuu7uCi09l5rQX0YLcXt8xsJBDxO1vTEJc4lmNG
JlktSSG6joge0yqFhBGCzE3k0w7dfpXI/s57BlnlxNCC3MqdZc3h/sVa2og0STiM
DJ+T7xLQdrLmw7uof6Eu0JAQjGoG1rqH0JXjB4lkS+xYWvAqqrCM4uJRUq4sAAyr
QeeKDIcvsZdRiomWdCyi+hEhLp1bIcDgME/9JCdJrg61JpHshke9ijgRq7oAwI4W
FoH87mFv2QrMh/0wDirhlStDfrD3+8W/a0IT0GL9VkekWw/GXS1uvVIdMDEKYI4l
m6edz36a0vMO1Ip1z2dWp0MrAwVX99rYSYEMUZ+W04Dd0LISPSryTmS9Q67zztzf
O/XUNAFG+8BDeejyurrIua4fTGJ8mgqSF3pTs8DhAbNwZmZlx01N0jbj5jPbfZok
Tngjx0ikW4GMdo+shxYQ9HoPG7RT/g+Job0A74UKx/0nF/o1TN8C8/EG2j8UZWUC
9PpeFJyNvPO7UCIbCK0ml+VpMRv9sGk1+tI9EBeeJ1+KndSwm7iU/33/6Ux8WuHm
5fUTE7PDtGjx/znwaPi2K1bI/QioT05S+PRIke4VdlnHr3Xmi9LLWGoQutZKhzcc
d10e22F03qswxdIUSP3M9ONpToNDnZuQd3RxK506C7ypUSPd9f3OHtiztjxGeV5+
ahvn44W7jh456Ke1htFdYoMuOm+cPlFRHOIbT3YPtadKc4cVQHo/e130YUm2mcMf
iG+W6oYtp+QNFRtV2RCM+Ojg6VdjVNZOSrAHZEyEIY6BnbIvd57cUdkjD0QEUoGw
Z7Nav++mSr2eRU97MsX1YTac+hfWEKyALnIWcqGSvFO6Z0sWsei0iwWtl1KcXHCj
rnQdNpgbgJr2s4p69A7rsCTFxHGCy79AGXD5eyh38phV/F2ueGJwjOdoykNHn03s
olQTK5XhDGvhvkoqehBdzg1BwJnw30Rg/D2qMNbiB/g50pAM8XrHQNR6m0GeWtI7
bEiG7JOIxs2sKqDc2tA+fb6UZc6Se2LnPJ+1b3aWbFA14vgCj0mbsg4t8S7peDYY
VLrUUyQwGx6tVEu49Oaq9JSRNr+v945bhPhp4BQr/FZ5GrD6AH1tJEwSCzba6cSR
5mH87JEFuGexgz8e8NxK9bGNnmegtZGbD5KsZkjvZJ0CE9hJiUmRmnX/6xxqKPlc
OovH5GFRBQUrwFbNsEZ0Nrr3DfViApy1jyDjTg0Gs2B7dR134+Kg96i95Hx+XDWA
UHlRU7Ie/BvZRJpjRmLqB53JL3GVwTnf3f7Kc+Wz9pmQwXij6+Ka0ZTIHMlxLGVO
ZcYKDzHtypdpx1CafBAZaR0ESBFb2rj7PMc0SiY8XT2hI0GF8Ee7JQBRiM6vqU/0
hLV+aYhLCeiQiCK56jhqVr47AFr4MBv0p7rqQ3IBx/JzzNAsJJNCEJbZZ8DST/9T
eeSr2OKWywfJQ+1fTpEQBsgpAXPrw3ophnUuoA9asiUDjPdloibr5wlnZZOazXmp
VgPs4gpqtmPTDvfYjpqmhPfrYorKUVE9cZJ9KFWNVeYi05ercAI4tzLPR3UT8qAI
Cd5ix4nBE1VTz4lYh/RoHTBubHH3tZi+PNsxTkDVBJEb5a42eZtcBse3aSiJGje9
QOt+AcxYvachUOYPtrbK7haG5Nxc8PNtzS8qKE0g0y/TE4Oh9NzTqIvckJwFtx24
Gx2kODffD44sDxdvL70zyAlaUvvxjTZQYig7cjUsGcdLeIPjq3i9lt2EZyUOSC6A
CCPx40ckYeFh3mQDa3pzdpcOc51Z6k92yd/THX+6j9rsOx6n5upuiWXIAREfu85t
8dY0T/fRojzbmdLd00/XroYBmVqYcTH4HZNjXV6XPzoRwU4NBLNSYwp5crK70vXP
meyak90+w/jTTLH9QhUb9FMUcIj/1L1aA0euU/2pFIWada2T4fu2Ne8pW+vb5QXe
5VixGSHbI+MZC/OHihzDYM7+B4iOV6+3YE88EtaufekeQmFEXTOkIssU2jE2YDWo
YrjlKYa/ZV1ZzZPxyXutu+torGhMVZyYOSLeV6trEGnV+dP3kz8rO3xeE69RrlkC
+TQ2NA41EQSRPWck8Yj7CrCeaTFNP2dhgcmRmAVK1R6yDwHFqrPoXp7MkM3IHHrs
nApIpeuaBEAdVNSWrq250SvGAtJBJvUPWQ+bWyw6/nC7yqQPTbndLVwvrHjN1U6l
5PomR+BwPVGelBoGhNk44EF/GbOVcfImxa/Wef9ofUnrw6edVd1I/CTCRca2cKFI
PONT5tbQxRgohmDTCbiqXCgrlBozi4266SMBFG2veUi+nWYte8r+m0L8TkmwmoRt
3zMEQwDHczMluFwyqpLPe6nesUWJRd4qIoC9haKuTPtzCCsiJV4iEifOPxU6idMt
hPEzf8ACyl3zhsl6tHdIrcGTtvmaBWZ3gv/hlIlGRd0xYrMRnj0zmK15tLolZEBW
bSmCeFPaXnUYjrUDVBkmz4UwMg2fz2dku7kFBYit9gTGrgs7eh91hxncMA0efOI9
k5L65P82Z6heau7ghnfywWlYGdDPdqPHMXGJs1eXmBKtenaVPNkRJzO/r6NL3kG1
efk4tYTf6/tS5f0x/R/hP/waB9ArfPYQmnnRQVNUifuyYu83YOICoKZ3FuoDhgE6
86vYX9Odqj4znxyoRnnJvZyvXilYtJHSGF8C999Fwetli5U4gJiLkAMdRS0KPpLo
kbNMmXwKxaFxv9y+RkwfRJhQ3BRf09MGCgpcc+rU8TF38VH4kkuQYXJCmRMAeFsl
HSwHRNU6l7e1MHlgEOxFFqRz72Y6URizZsOYcoiGn1UxMEaF+N2dSKmeBpuighvz
IF0axWLGhuw/PMdwctQb6Eybg+hpcuW29S0tFdoWDyn+/ofQ91PBOgPFPd8pp6mg
r+B231Ml5RLu+4UNjVuACDwJVxeFvg0byzYy+IbHKbWn+2rd9OmxTh/2Ms6hremm
sZzNDwX1S+4yvPeX6MdNjCAawM7Z7/xQfdT6Rf1T6AOnaGuoP5TFd8F7b4vqHMKt
/JInKVjgTJuzVEdkiVXaYOBeMp8ugekRE8omrrUK5HgjeGg8nukCT/p31TeE4dAu
QYxxPWGEhm8gInsKk6aEA48AQNr6sH+h7uGUNG320oDwMb9Wp2VGE4ei329mYjd8
QNbbA14Ge+FCFmxMvCC66d1/bgD1rAnApPsOeXBObqoqurBTUI9YeYARULYDOyGw
Db1byeuhT8l9Da/m9deZxMvesUMaBJ5EtsCMDb2nZJmWUMdnknT2upTdqZSSYiBD
3DNQjbNl2AhyQNVwYsZ6kLiSmdPSs86GgtibjOqJ9PdKsQb4l/7JeMxZT8FZS85D
Ni28GgvrY9SRcabPIVFAydrNTSRyMcBEjo8rWarYJ+oa+AR7/Lf+qeyUTpzM6yOV
MW+x65IYHrdBgujcYrCaLq9cNmiQpuOg15OFX/3bAQI3YttGu4B8qmrtUvlKecTR
0+zZgzPkNCZTei0MDKsBbYbY/l5LOJg9Q6hOmpDFv9W9h85CsFbhtOwHkfbFcrsC
/gmWJKFW6sBLz39VTmrOn0M6Zki81wd4IzFebFrRhZULLfHFoM/E93+WDXUY3YZU
ppqGrTl7DCIPIb0vmJCZDEGRMvIiRpt0/8C04P5c4vL/Te07Ws2o+f0NcM2+Lo5M
6MMlkoFCCfmHzkYq7577aHxX6frHi+0KbytLNDKwYR3xO0yVLlMYRBI8gj6/AaIh
lOnT5d4YRUzjOv6qzQUtbg9ak4EEDEzoJ7Z05ADRpWNxiFCgSin7vtXIAFcdT1AU
IPyTRkTupMFiZQiBaOFTHvoeCpa3ekY0jyistlNyfm1H4mIuzES8b7PP5tPbzQdS
L6goiV0QqJrFvRMdZCu/KzM64f7YddR7wgKTfJbniUjY5Dm6EVafPsD8gSAVstkZ
dd6IJdpwCqOBxoaE+Xaf5Jig8fvv0Mu+DLQigoG+cZ7frUbKPgn7bhrADl5xCiZZ
GIiLg+WxOflJqYdAqgcSg3pI5J3bahdBBhqDDE3pLGo8OkieJIpkpBPunAT5ZF/D
qLcobuAi57kTXi2E4P5BJfscbkWuZh1MQKC4BJ4WnzdO66nV17VtT7u5LKwisdlq
Xas5FcFMChzPdImvM64O9W/62SSzl93qJjXtvcq1JhbZ9s7YgH5QND/nTlM1tBnH
BHDnabvSbYCxhWimRd+tj4vymhlpVIrCiw0YqIM3nIklGO39oH5HX4PBNyzAb6et
pmo0ETrkQd9vIingG5ZFiXsp3jRNypJCI1+uW5fh+eAxhKqOp6u3l4kC5K/Gbi5J
MjRvw/JCAFUUIPUf/1TsjQG7wrxJYwotoSORZo6ONhDhZI4iR+dmCzGQzRxmncbR
Lcnb1hHRoDlVfxgCkxZJHZCKj3PYfz2xff4lLgdnK2ySzE+UvfLqq5QmdAJZzsJK
BKq03Nnbu5Stmtw0BXBpiw94NgC0Yrz/89lszhFP2sB7hbKyh9r2jfakfV+867oB
RF0jdX6KWxNfmzDazFrQtu2h9AECrOVDGWkf4+d0VPU5Kp8W/GHxWmr3Hc3ViIIB
QIXakz+lQiB3AI/P6h9zsk5PCZS6wnDZM3Y6m9iQikb8hQEnqPfizmODFj8aPElg
8jzhm8vLxL616uv2XbGv7kfmwP6tjKU1Q4xXOlfhKqZgK/W3jwcHgLOY4T97Ourw
B5bsx5jhrhSgqJm1fwm6jSZFyWOnxjKH/o2quK7pSYAXD/nwsDj5DFBggFLn4K/h
1kGipeOZ5Opla6iKA3DkXo/MtS+zhsmrXSbS+jyy0+njIFvAOxwFz/OISeuHyBuy
L7K+hczP9wE8XdD6M0zqzpI7ZDc1ny7UCJVKAys4HoHlP79B4QYXXxR9rMbtSN5C
ltjTRUAwiNKP4bVjAmgAA2idbj5mKQi/xjutW/LCyGfwQYD9OGaM9VNyO8OrsWxc
sP2YW85aTZMwOYO+lHphMcEyOMxTke3l7uX3NeXT8TeWWs7H9rUpDcEl5nCX/Aoe
U0srPs9FCZ9M+e0D0XJfaL6TTefgluSKE4fGLvXjQYq9X9BZMlebvKBpi0Mc8u0i
MI8QUVraxy6U8shRClu973xD5Wjo8ozc3iNO53ga2TKAEVqr0bRAed0K7F/WELja
75jLMb6J+RHbJR30SZJEgkQfCeteyd2EDAWqTy1t/cHaGMK6pTBiFzIH7m94+fsg
w8cOHRsDMRJHtmCz0bYkRo3CMm/g0HsPImg1UT2FBAVhjZ88ZdHUmlhSbeEhIVD2
hmWgGY2lc8d2twEuZLFuB3c/gpBBbkDXw+EcpQ+F5aWr3c78XFA0MyVHFVfH+PM9
R0nlqRJEmo7aPfMCbJ4EC3meeu/ydB4Xeg5QwgNLGxA9BWivh7EpL6FsIjhegrpQ
RKxMNHpMmVoJOl63LyseCvFqwHiJttJrqwYcgBg8nKPmJ90iLmBYmXAJOW5NZvpK
rR5FB6yJw8nOf2c1/Z2j1BH2taDk+SzBklBFvGsRKnZ5yU5x7T5z09lVoxYVQijy
n3169+CqNCUi9fxHrqhpQSw58ehCoG3QqVqElwLbU+cPWRdrnt2Lv+l95cPju52S
bfT8nTCHwydPuDumJrQS6cn/6Erp0eKZlIQLVZ69mxLr4vEUyrVDrbw2RYn/mDLI
aCqMbTO0QJylR/rKMRjOixXcTfRhkdpq3nCMlUKF/UstBLYqyqnlZ0k+MdESxxQH
RjXhz2F2WSonl3ZDgOVKjNNa4DOd3b57qNFlmXP7blMHhPwgHEHGaWF8gNkss9US
cxdRjP5EpbiS/P9wvToIaYo7T5edvZn5osIvsMH6j8Ca+EenXlDyxu1SqyOa45R2
UlyZ4EoKa7IXH9MEEG6XGBbE8o/sDAOW9ZnOSbLnyYKYjwLAuegf3XaYXEQO7cam
0jbHjIyNksqI4eoJUBDriXZEHMmxHWVsOepL9cq94WxqAMx4buA0521C+0Io62gD
vUxCjeSum41EdH3e8VUzSlXfz9mYd7ZiS+VG7jX+mFJ0Ww/TYlryYzFIivNl9ROD
yiqaY9L0upZsjzdCdAcY4XhXz4UbgP5C4uwRzVSG1vYDaUGy+ZsDluyhtrPQBFj1
p/Ut5aNY3OqBVTESA3MZP3hAaJksoUjsous3YIlMy/qf3UgDLO5lcQ0vwaFEY57q
4MiEohTrojovxdiR+cQq7RotWhsRYDahhxme9Nu3B545VcoFsrEOpYQ2B50Fu/1A
7v0Ms+8Tr6ZK0YVty7DfLlaaTfv2kyBEgUP/s/9yG0xm1rOUdiTY+rsEyGb6btQO
ohSFqi09l+GiB42K7NZDZoPccBlcO47gBFUeGhLsMLZQoV4bwdnJsKzfwfrXEUie
8yvHA7betX2oFgy7T1i26d+y+qu6+iZslkllBq6rc8kqiePhRN2Yt9y1GQhPG36u
LLxtszpJHjXKftqeDCf54eJXI+llHdHn7TfYrmFF4z+7k3pG9m/Mml9YJi60YIo0
gQOP720AVKXGx40BWC+fwV9BOxsxQZ0eRUdKRrY4TMIcQ29qEHcCLQj9rQuaCZWO
vO2oh9LBvkyBnbP0EksfbzEBrfhy3snqbrnjwb3E2D4lRep2tSLGM3HLGBgj7AiL
rjChnsEhJaHg03ZW/0Ye2sGzrrTEakHw6lSXecRUKigNG6viVOV9SnIWodPhJPd0
I7N1foV28psu0FLFmFIUeAKHtZy1Bv7m36ivMzgT51dvi76Psf1FFSR255DIWLXz
EzfJPxhuofsdyhQrg4V6Kp/SvNo82O+GgOW3ETym+JLqUMZtC1tPwFwzM3hN0hTc
PzekqSLXO6HAs0e+kbx9ZlKMOGzXU8+S7MzuWfUZRlFx6K9UFRB9wGPuLoxwP+Cd
rqc2RDmy0HnMbwSKuFHhZEacG3uiduS4EX+gtemy8DruOIDve0hvwL2z9dXAqyg2
IBF4Gv5jiOLP0vyAIwdEsPfuuSssqbe0HRkr/n6r5pmITBfTQ7pwPVcJB9cB7rIk
Cp2p/kRljrbQnTXMH484veGeDMPisymeFlLwDXVEyx8uKqd+r9vsByd6QQpxNBhG
G5r/ctVTgzWNBTafVc7eIEc4HeEc5w+OhnEdaisMWx9SlOYXecIeYDLjYkNmVUuu
/djYf6mhxKcGqOHqw1q10iTiytYvduvJnGiuk/DvhkIZTTbKWBFmu5UU9/vDxRhj
ItYNNiz9pptnlaK0qlB9k2FBAiHyiToi/0Iqe4GlbKHqwzxyKzFRWeNxdNvfdpb/
EbbO4+nzBovTvKKlnU2k6yxv8q2ya5wYJqrjxpX+vFTJ61sREm/+gUVIeILrAu3+
wCT05D1M0XMSkWNUwVY91OAXwtybvLKA1b09SreRezcy/AWZ8gQpdD4OjAJEhvZH
Sy1Ux43+eiOQBQkdDKoPqhHCkEOL571d9rRh5+nY/G5/ApaSE6m5pQzX+ibIcGHE
VoDP8QxDAzKtLOm+ZXj9jhMWrgXtffcamSapXyrsutiKIJq8D/+zia53X7Nz/Tow
KnjGcx5qCytpIdrer7gMHU+yie/WE4FsUwddwlDlZ9JgUX8NvefGzsyosAVA0s6l
nrnP094OCUam5c0qkhiQvjl1L7dnJJ3Uguuf8yV9kUejDi4Tqki5OfxsHS1xA0Lg
Ok4YLMCslILomWzKWF0ZMBfOHmcAETPgnkzLZhYL89OaY+JTgyUySMRLRR5u0n+s
8UwWtYb053OXsm9lYMYD2YAYIvDVv2WdnPW/O7LLF6hIYwGHHWxT2uD3A4eKpBpL
xPU2SG7d5hCmoQvPvx7R7fMNzHDzlPySRzKuhKOOq2XoM3RsgDHIEz4K/qbnlTtS
v31Rd0M2VLEFSQm+NYqCDQsCk/+E/HldciMBpmNrJGBFVdQwij0Q+XErlVMhEeJ8
jJege2yJWHKZbMiJu9hB70TfOF061ZQDmtn0RZmO8eCzt8Pcfy4Jrgr9XEclwd2a
kDwEXcsg1Qvq978waGxfnOQvUcaJDQxAFUcTO00ZnGVOpGYtMHGi6d0m5C6coxwh
Rl9BttL1kGV+K5SAx81WCcngpW72y93/p3L+rPIuCxeww3ixxIGIKO4XaQ1vdaYs
VmaWEJpnaG6Fkotf+6BQcKYKjhbOWns5Hrdn2NMflRDdLT+s9Oqwr9Mwi9dxmvpg
jvQnkEhJ1SNgnrPJjc5Dsi3FpBWw7u06WuwtBLkOwwUktGTESWrdREQh7k9ZHhbI
vmPLxs79vTM9HdhTqIhRb+cHEW9va8W1c9MZ5ccHkEKxSP997V7lqzy7ut3b8Aju
bkO20Ng19fCFqyoOaMOH6+ws6liQlM/sJKV67v8YxPafWIsjlcWVtNcOff5zRqLO
+fAkFGC4lA9w1yVVM8MgLolMOLv5TjmWzvnPFay9NucyjZp7bO5Ki4PNpEfpfEjN
CQdVSWKbKZTr97ei2gy3sVwPUbPcaxOuB3p+xKsN7vXw/CGmIYVQ3inPJX4aOXlz
TvsSbDhWaxzes9yfjGqrWu/eCPZcGbR+o9w6ECT5HkxZTpo5vKv1V2WzrIBk5pvg
JIxlBkyXWUYXiy9YH4KFkzyPwxU7KHfQatb2KPAmv1B04+KPr9RvwNLibKxeGYGi
vR2xeSMnennbMyEBzs5cCH/x9G8F1CQ471lg1VlM9Be8BELA5n3wVyRBOXVwMww8
XoIQ4Vp2oCxixqexKeyQT+/+j1NUGwJM7l75NYyoNlaXdJVr66uDxQlCQCFprRRp
PboFQz8h+v/QLi9dHEGe9uG8t7FH2TfGTFrm0v+r+tpPPBv8Z1ZFdN9HT818EQa4
OwEuFHoxoor6ZzBcWkKdgA/oYMvCYTBEOsnatZAMT0dYzzYFa/0z6VGPznTMYdNh
sU1rd5WmQXRDirMR7tgy7rrc7WRZSUDlT/NdldnRjjGnqHKSnQDZe5RgTXu37N77
o1rBzq5iSqUZI+Ttab4aaeiSRKeFYEF/gmlIjxdiUTxDTHi7Aptz4REpIFUj9nFK
UK1c91MQ2ON7zi78DBM0TE1EDlquqVoNQcOW5Nw0Ipj+43639MFHCu0LQQCeAEf3
SnR7u1t8wrQWpceQN4tnetdSBhgIurbK0TEi1ZCA8yChJW4LYHsaOi/bD7kXfaTL
TS0pz32xbR/XA3eTjg2YHzgVL+kz20G4TBuTidN+YRjMOzsIBygGQ4EsDhu6bBcd
WMsodspabS3ZV2vK34e85N2q2udEy34ub6kMY8IsbKhoa+mLGNjGk6Idb6PeTPhX
sPnfn2Nj+/aH9fxgCnEjXk+Vpmv/xuS0caUgQV7a9TSsIMMdJHemAoB8PxKHV+7x
vGV0/HsccrjePyWs2mbFNAG72TLA6DlYyaHeRmZ0KVwAO+oiA9bpazuZH66JoQ3d
I99GXsj/d/APgpBVQzu4qM2dLtTq005JyLW/sDGuj6iM4r2VjafM+Rqn2T6eIPRO
NXuzIP8dMHJwAc7ED4Pj0TzKd5Nb1npsxJ187xGTjVW37p9kfTFQTMb+Y4yaCSsZ
MSV9iEjEBNTdzUa1sOmMDZzKXYAV10n/rIana1BwIavLaXA4h17cx5+g0+1TgUbq
LEqFq/NC7qcZuvzpha0h5r7FouGl7nkcVQTl4+PN2NCELLIsws34gq5kj083SNvI
WSwW7cvzxaBl0MKFAvm1dA6ZMPgQYHjy8yMLARikHyn0yWmcnaTtrVEXJXeOPp3d
+sd1tC+A4fECRT/xzNWX+OMdYc4CpSx51jSb+PcTsoDSOmkBwxXTy7GQW3fEKQWI
RsNSzP1ZDt9OS5MvBiulbXQRet+BPihBYydusBC7U6TlG4V9w2d2zUANFoVdrAQA
kq+j1Ra6KQujsNwaDSN5cqbEiLrUk3DF18n4xdzULQoTGfn8Nla4OttbvjB6o3By
IpVdZ21zDj0vs663gwgMdSMPO1ocFI1RZJsj6yR4vdlafWxQ71Rw0ckGlXsTBbfc
Ks7QRsjt7UXAhwutqsLgKE1Kg8gd+yW7HkzG4rtYN5eZsrnT5jKyjPjMoUR/uMWC
t5v5tMNFa/IMmEMEyuj51ybzM/Z6QZvTLFPP7dgtb1oBaYWzZCYg0y4VlnYLReMu
bxUOCfuameHCksbNntPKw0Uwu0sO8hDtblFmrRwye9emWygc4RWiqyP1WcnBYSsM
Lj3bP9ANIbKGULBxlRXMIfO6JteKod79IChOktZCse/W5YvhUh4zyCJD1Rdj7bdn
dtxM0xjaeAhYPwVa1AZeTcakkb27Xx9xBvm1daUisV6kFbGPHxom1nvfQj14/uk5
lVPtSeH0i/JaHbL31JkefZTaUJ0L2bXtLnG2qDZnJthKkG3qbr28m8DvaZRRH+g2
BPZD5kO5pSqfHNuM1xGQ3CAPtD2CDcwudAyw4vUoq8Nw8rH9CK+sIfzlxY/Vnw7E
TurkkFMHzfX54UXzMvKaV0yH/eB4jYoqXPDO+ZasU1faok6ocUMtbB9H1AcEhXiy
+q6PG6hmsAwE+LmQmbRtvbOPvwe+7d5NADJKjCLqsQKiNM9cUKGQS1AHK7LkvZfd
hy4vXHuYTMZ7DHC0N7PjIGj8mDs2/FHP1sGySBTAgfnikS+iwAqhWFqccwVNj6An
A9QLbHRCCjGR1krklMLppjOGwXbtcVANxkdGYx34s+gKB15iNc7agbzoAFWS8U9b
vfUsXQE2cjDmRI6v6oRuVWxaEPPf8D+X6NVxxRzaqjEB/1ywUbg11UQq2Uo1W1vU
Z1BPmqSaF750vxzbDpj8y1BJrZ0/rgz9b9zl9AHHOVTBsN4BE1VIki0Vjbv0u/ut
jVG2wWlMxc6oHAJOiXbczxf221hxDhIgpGyXKsaAdQLBpy8o+ATBc2wNKRY5dibK
L4ujETdld668P2kN2AnJklSWPiNw72dGLX6jjtOQMBTSFWLJ+w2QGL8j5dXAqHKN
UaUt+7bIv6/5kWyZCi9y2OSnajq6Qro392oCctoNBFgf3u4w2aDMfLW3NEtED4J3
zxDBPxQh5VfLMDCcpi47HJusbiHAB6PlOOg7fwGhxnlgxKC4nWinhJepKRmGF4X3
quNkaWh4teHVQFXHKkxxg9/eO6El0AHI1HSiCEUQdrKMmCgMpAOFHer0rZ6RP/OE
6QWzTI4dwK+bRqYPWk/7MlSLA1a+kC8iTGhHDuMkw86TGNybVZEdedWHFgGAPAYK
jeNkllh/m5CbU/20Q6txVVpTSyMqzwNqL7hsKZ5eo38M/OELT+FYi516yEnBzfai
s2kHeaBwMIXiQEGZhSOThLdBUkQQvKmRkDScanh4VQdDQHGRcwwHvFGWBFIDRGXV
NZkcrexzFiSP9x/LIZC/s05TuMfIf8M2qoihewAjr1hduiGewhjxCHUquXws0ysT
J32fWEqQxU7DVeha1isgAdmBbj6O98oMoACNHkePC9BiUW/tlTJQ1f7TeHxSN6zw
723jF5NOAdwJBxSpYxfFHsjmXybWTu0QaWXYBueI3RciNpyMEKqz9ZGT7REzfU6c
8xrgVv3oKWWGzSib146iXNC9HnlNEnum5KCF9CL0tiyuTNiZ4eC76BD644zqcbwp
pijixw11fTBKGxXrd3w9FI5HnfzbWSScSL8Uj6ZoWCljzaZurQkWP6mSvfECRaTl
kgwaIxmRQsMKRYf46ZpUtZgETX4gPHSRrWCpzZrHh7S51b8d0yAgUtL2ys+oYkHq
4dFPHnUNcFjMNTAHQGrmXakEvOgyxpnx5Qjn8VXOtd9xw6lMHaq+vG7fqX+QQ0uS
YtYZE+JnWM4QeNnZNUGSv62XuOO5+yZDxA1WGw253fpO5wBbqnbFzXWB7XazIujT
kc1JyIsomvL0+3YwbVcNyJJhvasC3TeZE8R/GZ6b4+ryCUCsM8ZjshumKlwq4+7z
6w7/XUQx64xnsUPlYkweBtttyOkLc97atTatGaoJaPPebpJD1Uv5y5vUj8YYBh3z
qyxAQ1GBFQ0kLRVh7Jie4ZzeggDEGj3npMPiCa4TaKcZkd6+fYfrNPO68KPps3rH
X/HX+n1TMl0sfQtVdRRbxN1GFOIANAJ0RX5xO6Epf5J1fz1+cmLDJm+QNK1m7SCI
IPJR9kSaH68IUvSeMwAGvpO5Ideh8aqCF2bh3JPsuOT6FN659nQbmp2ywTIzStZp
RRgQSIoDLKeIaWz0uz9FP1OQr4PlLMKYPv/MCVA7baBQ4Q+lXHafcqZPjo6JF4DS
Fu8vomEClXIFYhd3THAbrxczZ2+a7RZf7daS/ujp+YasEw9KxxAMtYWKFHG4p9WH
I//sgYz6M6VDn0Cls+Qp4NK9WTNEFYDg/O4MoEMyG5Ey1tumH9EWCtvnEKErNYiP
jexBLqd0Yo/w6ABYmUoyDk1B18+Pjrlr50ZaJd6k4yCJ0s5HbMkLSN2j1qCL7Eii
h3fdSErn8RE6Dy+4r/5FT60YpZ/NbriGsb3Vn9t+CSnTv3sZymD+Afn5l5k9lX7s
eJRm3PZs/5JocPf1bZfWLiF9vg2mVHaOTbpDQUKM5eEcCgrog1Bz7a7oQzghePNx
LqVNkPuZ9ZuKO/9jqLJFPHXyneh6SueNy87dZ0Tkv/Z0SdHtWpM4rza+NKHRG/pW
P4//hUGYj/K1pOIkneiW/ahoedqiywWdeTDXLmH/q48RoADglEUFN0pcxqdMMe6p
0jvM5QQ4vuzFpmIOG/sDWKQ9IV6l6YZwL2y5JEaE1pMncH1Nz+BbB00x8kSr2L+o
0kydWOWEtmV7MUOvjasnzRSwrclaJfZsMZw5NNenETJ5H/XDLgQag8RmHZA7vOO5
vnDQ7feMIbM7Hjc93lqK/pb0Uy5tWqDZkuh+hitvAhXcCdA+5cPAvoopY3mHfBsB
ppFe0bX3IxEMED7Iqk+C0KM/oHR/NVoTBwUeTXrEa6Li/AO5D2veqtWRD+afWRWz
XrxZKF5rNkl9BWEnjJy6m/dNuRg7tj8dVzPfTVBM0dzCTekw+AjWV65Cso+F9euD
mozSSW/CGypNKLww3HK9aCXCTUSFshhBWSar2l+3QuETCsLadJRyz3b84ZN6zutx
z/WZhRVw/5CqvqY5Lw2NDp1bl/3ibvbKNdSsWcxqDoUJ22Ulo7nML/dlET4r0NyY
rzNT5aCmDMG9jQmHEsZhOXorYJzhHnXJUuj9XcQ6pz+GO9erf0uiz8CfTQtH8exc
VESlbRcHhbEcUqRuLCOJng1sImLCJY0s3GuN2QR43d4zF68f1KBRxco1+LuhdMwu
uFxb3o6eZWl23C8yvCU38W7vwv0e9cO+iuORyunClWfYE1RPa5bmESma6I/HuN8m
XpU2v3yKXQ68C+sUV4DmYPB+dtyXkfuDK0mAbYl/1GOmzOEycvYxanTXzY5H8ONz
50PW61Yozrx8mvZ83kBjWn0JMbWJ5uJ+gKNbfVo1x2Xkkj115ZbwFQpa7NIw9INL
wdKtoCkky9yuGtTyAVL97gxb6nU0bbHPsZkXy7chQ7zdI8vtYQ0JDne9JXUH1i1Y
CcW3NvQ4UQjwMQhmfEWHsG3rDpc0gBAOXJsTlABSBfMbGxU0+ELn7GNV0pyLIU5L
7lkPWBI3LR5IjqpgO/QRmQ3liit9fhvh0taTBMSUsCKB9hhgvQ0ulEkV2XkVzz77
6f5clkk2KMgEi16Yyr1eJ8d/Hmw8r1rsZe3/a/0TMSd4qUtE3ZD3aGbq9P9OSMFT
fSiWcU3NGlSWK4Vtbdn9Ijlsd+D+1eaVdn0qTT6znyClz8F4IaG5zKSTMDCZrWp+
1RFAGaoWT20JWbAvF+DvOkz2iIQ0ZcC9V3XA2WdBLh5+SOGZtl2KNRUcyFO4+uIE
1xTQ9SZr+9HAslD51BEiMPxlr7eh0gDOngjLcSCbY1Iyq+RU/UVsSNdovFzSwCi8
GgcpFU80QCpNgDOVlLVZVyjYRyKWl3DL28xLNzHskqxvZ7hT4sLrdntIHjyp4uWB
M1acUGKaZ6iiUCqovhEW09YLP91xe70+mQp0mLN4KMhadtk8yKNrB9Fh2pM+Zn1S
e9n3uq3lutxcD9U0jYSV8AgfMmDlbjKF61SPSdySUP8mibYULsPtGnkyYB3e6Z2d
6m3XBo5f3nKAJPDWmeoQGaUEuVjcCOgF+q9kig6gIeApnBImyKoQZUiVI0IJvp1Y
lWSqfKhPj/NhLcJ0OvErroZC7WsV1vkutEpr8AP2ML4ojpeQw2K9DCxGuNXHjltA
1GCcbRpZra/zcpYyCHluJtDzVk/yDMvdVlj0bKQ1EJW9uuq6mzZyLpCAd4E6V7EQ
aYRWDCo4SM0nillbXgNmSM9BgskWFAAVa+6RpxBjJFh1IxCqfYPTp0DxZYNPCpQR
JpJX11SQ+dSDlHgKrR7yT3yre3hFv2o4MOGzCTD6+6QUwkC6nHe0DgnLwzvkt70t
Azvh5e867j3oQ8Be5m4//1XfVT1QyqqovOFnnP0tlWHR6/xSl7C8grCgWBZ43L1f
UYcJvO1ef9EgJBUF8OEHLIaAVBIDHF3kImQ49x3/125sLGxIhAawNTi86IzYn4L9
VQHqqQ5brobGKwkQKUPCHAlvmOZqRYYmmPpnffenJWee8UK+77Ooy1LFjwTwrX/D
c6Fz4r/SFvGKPbfL+W1PsYLlRs+Gq88tgybqwoJ4ARP+GBbin+5qBULdiqPzO0E6
G6zXGyN996+n5pcE6KAEVMk+ihkCiDtuinJ5saEVZZJURoKXJwO5HnMjdxyjGwnR
UgN+usIYJPMWjG2VpjTduo5E8KuMWVSpDkp/QyRR0Fc7UG4CABrnaGSBKXYTp3kh
b9cX6XwcHLOtMUICro/Imy1NmBmI3dLNzAl3bKmgw0q1ML8uorXbQsXa5rG6j0s6
WH9BubHKyh2NTot7xh8EASe1LjZ/5KezXJHayXTRUgmYmcxFoJ27+fbZFgNMt5+0
XJTqbPumbKetWTrsUNoDRDbn7zHfMg6MIRAk50wfA0Y+JdNdm+tTM8MrPtE9KQP1
AFav+0q3+Ym6FyQg5IcW+9EEFpjZBNr7rnim9JDQui/qkwNiHdFSfH1EbRqAVF+V
TYBQ6FsZDDgG2sFcbvPX3KVNhIUoTELfU6bb31e8Gy3Bia9k+h3TtkLXibRbjy/C
KM1jYnZvpcvtNoKbVC+0QGGLP6AiONFG9v/kzWkodcBEwzP5/kzV2a2aw27ucMMA
VajJT2sepNPTtR3E0Rb7icoEnWx2Lue2tSMLIsBpek86SWwxC2vj5a/UYIhPWv0E
2CZIQoMKkfCLHTMrCRvsdIUGbuVwo4l+XW8n4NWYCij8vWEM/zC20LcVWbNNnr7a
1SVQrlz4qBDypnI3/YmmQL2LqRhmEWDY+hqNzMQ4RBnnej9YKCv/puTyrAtb5NAU
lHhNMYdApNQIZc+iRwI8Jn7r3YnmZfslXCXjbHiYoIq0popIS3Y/CFLKxb6BdEwM
xu1I0swtd4Q7Z+jky5dG1pe2rjRsUmP5C4vuyDyrozyyTVpthLa1aVZmmqNFvwF0
QqaRliElx5cpUnLzM2ZtQh726auhaluHBnrky2HbkQP54sttdjthWawfRJJJWNWL
LKX/wEiiDvhLCDRdZM0fWi8opmE6eLQvrsJx6pc62PGte7cYd+ufUmnHWVUcZxIK
5zGYDW5JOvcFJMkTDEWOv1UAnJ311kvGZufE+lomkt5DjH7iI1wOzRqW0surAFaV
eeTIjDDsvS2RZGQM+2KByhKnc7af2wY5eJsQ+ZkatynjB+C9ir4SLOCtBukbavtu
MM9U410dLKdYQtp3oBRCIdrC0AVdkDhQeDQomtBzgZdRz7coVpUOCizH0ZuBJhnb
kY259czvJj4JH73iU+/PY9R3LgPxJM9k8qqDRqFR45IjhNu9XKSPrHGEHc7kbLOQ
51bukpeKePrTlnd+9qHQh8NB41nwU41ZbQh14rhzmadVmX+09S2bTlA5NSSZlqgd
5OI4lMcWReuyyXVrckqI2FBsNCK1MBkw86fXhB8+cz7k83yF+KzuW7DaIpn4L57U
vkNjoVHivgBNbko2ubWFFUlzeA+qL/sv0r7Q6ALjJoEhjiDVXSt0eHQjUT/nmKPY
hNn7/LLjq1F6nr7wSj+Q8F3fpcW5nLjjiPh0rywja19/lOPDPynHQfHWlNnA01mR
htwbZ4NXCxGzqVxlIF1Fi3/vkSK/tUpqd+arFrXVq+nn73AEBVmdjSQzVZMAbggr
zbtAoQrgFoWBNt2DKljrV3pDqrbP/yrQ+yxGGqrU95126ABGZaEQSjSn4cbxCnMV
qoMRjpfFxlAPq+w1NkA2SKRWCSvK68RG/c0GI2+j69BQvNzU5LSN5YmZ6kSMZ/F/
QTNnnVmdKeSbkWKLG7w/P6fZO/KyhToVcWXqF/Oqc6bbfDYxQ/qF6ZoOUKq+1k6g
CABgeExgj3/krQGiXr7R+hj2VjZJ091qimTBCIzxPfIBgisXIjmCuBNxF06DWwb/
/VMpB1lxXFpCrHtjRuNlPWyRsQY8nOUDV0PC+BEBYWXsAG1aUX0057n6Xiw4FZhK
R4FqpFbQKvb16zFajO8AN0CPIdihibgMePOkDbZTUpSxaEuzzzNbBpFc3cItSEGp
co/RILsyJN+aRf5fND/h1AtJQEgW/dlt/c2Q7AkLjYY9eyawgFB+CsxW9an/8Ykp
g/G287cFyIf/nbVv4P3HWbGN4BlssVsIVm9HG8aR8CTSLABt9o9bgJHbclKdpacJ
vKYowJ1uj1susoM9CUz/rDO5seKH+fsR0ho31pRNW5+IYGJCvfA8RTw8MKzi6/Uw
5gOwy2KSw8IoHf+B1puKSGDsNpX82nqmRnE1NztTUfo8SwSvxkMNvAvNS6zJPeUi
ldm5yoWeiIs1+IePhkNVBDL24Dtn97zHX+J7MTgPnuJYt4ADQs9ExSWsWyLJN6oe
PPwezM+0hzlA06HOD53ihcpYVP71zVaQokKbdI0hiW12hhn6ZXtzoisTqrZ9C7Wl
rCQmB4EM5nSxFBNPEftJohillBnpsqexhzOPw/hCkAeY7ME/iSGhjBeOmUe1qGw6
FQNJRTYiFqgvE0KIUQ/G3ici4CO3a63W7b9Zz6tXJEtTLYBkRyT/vRZD+CtsQha6
Pwvr7gY9e9h0ZpeL8uV749klXLmw7IjnfYSyJ+tT2tocIsSSOAXs0BZXxpDCvSbE
58pX0Ha3KkYEULoWyy5sYYqdqPmAeBkCPXeEfgPYPHDu39o/SwUzKj5ITTWN8VAZ
YJRTGA5oHizhZM5LNKRFFfMuGJdvGUa57dxIJ+r4MAH1jkk1WE90RiuUj/Kx7JyP
62whLVS0cPFlX6lHebdMoWX/Ve/dHTCkTYxy9Oa7Zu8dM5C+DWaVtfqEQi6sGRUB
t3FqhL7AnzLvkkq98gkas+e6QDc22YU3PkslpQqECAO2bsev8jPRSTaMjK4o24Sl
liiYw5Ygjmhim6lHzGiOX10WQRbnK98gAtQebOkjGhAEdvtlx9nbUeRXIDukF+gj
M20ijMh9evtQ8bt5Za34LyGahmHtAgVe5t6VmfxosTyE5aPYLVo7Gt4tb/mSThQ4
qt1cffy7wYE7kxcUWOmRSnQq9CX1cspDIGCKTSm+x+UvQoPl4auO0KUJCXBIeFAH
b5PO9FJOmkZJf5Y/6gwUfruArzJoKNPP+RFB/TSz4D9KXEtjYX6Vrqs+0jBPmVob
AO2d62XmH4ilOXBJq9gGfyMsTMW0+i6ztZi3U3QK2746zVFx2+091rCmU3T/eU9Z
g+UB+nBOK8BjzNmPUZQnYfUaokMqnJwvvqxmPAMr1PmT2EhYzbl9MkzRGlxeLZ33
ucvZvl9jOysDFAVfcFHqAWodobDRgeNFRYDk+DisU2lk02fWrlDum+SK4nHViBoH
xd+u7jsDbox+B15WQ3vUBClPIZWJgA1Ye31scEebS/wd4mgJmqIMCdT0bHKQEB86
gyQKQzPmLHH5pA+Be/CtU7E4JH7YLrLho6I/sxkTXoRAdnsZ9sF73HlStcd3B4Tt
IWrSPFcjF49ljG50nYCAH6YcDNMkJKxPRqo39eWQgsSS3K9unRw2mPd0Y4I6Fc1H
URdYNJVt8gYX+I7WP3nS9nIK9Bedd38/WzDO+BnFdSuorEbYL1toG/gH5L64XFHT
aJhtkp4em5XSEIu/4ZHGgAt4sPid7ZCZx6txt09ABkMaCW0vjZUzkZiHE81VptFO
YNS7b0uu3eFCxJUxKn58bW5w/mN4ii/SEzsP51igPew5odwKTskMlBYbHwFnsttp
MRlHRC1NUA+j2DWUVMfm+nw+yVNBvts7rsGdU/xRitibI9rHh9lLyMI/o5NsmIuk
wL9uSj0kqXJxIBpAi8BkEw/Z6oOI4JUu2yPT6gvLzzYFS1g4FoMiBeHHQC+g6vtd
U8/pSpbj2uagTf9nu3Vv9g+wxdqUUUxyFR6/XqqKclkTK4aCtWPUs1b+CwSGT0bI
LsS7N3cWygQci3NYxFoXbWsJffaWuxy62jLcmeYp4YolS8kVPPYsGUAwaFcamlrr
bEoBmNqNAK0mIDo1w/hlHwlGWpomQByxtT9QHasD5Ff4K3DJcPHbQm9ybxLiVABS
mspzcbNWgEVMG37ID+8SD+NSkH1EFU7u1ncE8HWmH/Ax/yVXIA4P8AHf56YF3t3E
TRAsq5n+3t75c6qMuMt1yzLiY4Rf3gYudKTJ9fh3Ef7KAvzg2I4//bp5vbF4pGf5
4ZFfOGk+L6NDKhKPe57FacNfk0RuJBM9WmpR9JHW/cM4ga44sEoavd1wfp1+vtWp
GMQFRxbrfWVnSqHtAp5aDwbBUEeVWyePjzsrOkgBh0yRvq5rles7ASOgAEVsiPc5
esw96ABL4jqExBtX/yD+bS5O7sTY6tU2WquJjDGHZuSm8LS22X+y+crrih1btuXG
iFmCvWzt2lJp5HqyS90oz6oe9BKtA1vXDm+NN7u8mvzuJG6oRleWUs18SqTWUF54
SgmOt7ezYxzBCWowYPuIh94i3RhotlM9UQuU/yFJbuZ5CRsXj8QPeBwzd2/U8O7L
M12rTLgYGl7dUYWQW0ZiSlkscUvh/gpQdZ7HzELHj0ijfq0yJ81h2VrUS7jWMY3d
cvK6qLKN4EM46B30CNf+Hs5QdCAMnts0rfgznnSmSl4j7Au0ZUwxJIqyhCnL7WM1
MrWIzA3YBglvSgmxDKKb5a0NXegK6MIyuA3gaUnYQpXiLtgXW/Pr2u8BAGQfDjhM
5c+smGRwRQM3IC8EJMomo+3g2GrInSLxP71rey8O8COOHLzYmW7kwzrr+eVJWBKT
4l01R3s4ORaQ89o5OuWFMw46LzA3G8b0mVkFfasIdspBpIMLBzX+Foube+Gw8QVD
E8/PQJxNgx1zzgPf0DZWDpB2VEA1wnfAtLp37rcPmiAMaqIHrEfO2gsrI6lq4a/k
ZsnI5fOiWIoIggEDZ0sZVatsNwi1ctQjMzQANAhFp4tgBEfOIGziBaaNWrwb2iku
yOv1ATxH8ioffQJT21nU58PDoKo7gO+OZUaEk0u43BnPSmie3zYCWDdvbjNFzvPT
ag4YOlM5gNwWx1f6T8dB0iVIcQv1Oo5moe4jSEcE3swJ2ArgOZr5UZBXlRxDjgjX
6oAzPZyHXKgn88Fc9KoD1L5MrjST0rrk4hvRUoWYKhLBIontQYiBs1D5mzic5tl1
9Qgal5vqXevMZC04xKwqBJgoxlxNlBfDIiSf8AT7uLZnNME8yK85fQUcyUJ9JVms
3t5woVoZWdgMNCp0y0avM0M/7XJwLMbMzzp17mCPZMqUSLqIMHQFhrcSIT9aD66U
+RiAHFADvFls5TeUZ7ptzxFz8A87QtPDJ460o+BDf+tc1z104XxW+acotMt2yH2f
eW6qQupj8YV10rrVwmFyvPsLFRgrXlUlynz5A13Jzy5MzCCOep/tggu9fM75lUba
/nq+6ly94rgDPcteHNNth0P+wGr9eD1ZrXRsh97r8aD37mEEQC2wBJ8NO/X8XKTS
dmC4MU8077DmEGc5XwAzR3H/lYUfS6ZcgPlQy0sQybbEbRCGoLD3+SMjnehGkpkx
l3ROmSY7O4CLcNAnN4h45/OpnKW3fejMvqnH8U6cM7OxNSZpAt2e9pnFPho+k99h
5zFxGRhxllt4OjYesNuqRc40iiof0Vr3hoP+0O1SCUg8zN3e4ixWbHi566OjtEJZ
R/Qeq/H7s3Ud3tvWLm8irc6bd3hr+SDTulj7VCbbEZcz688O87n4ERSytEfxWV2T
ED7opPRKTwTfEQ22MtQpZRUh3Vyfw3uB5Gofs3swG3plCOaceYVc2O5vcDyzk/IJ
tus8h2hI1ySXaAnXez5AnxYzHV9pCG1Lcb7pCdfh0/YO7rNU1dXWpJ+M82LWKR73
irCXxNrccYD5df8KmsSTkFlDbRwpOCTdXR+vqvFhI8fhSpWiahjpO1/LEe68h8mT
S/rYJmS+cZ4OiyYTcEbKQ+8Vn9I49u/1Cf4mxBrErtzmhb8xGu/zftVn3aBDpHSI
vOSk6AD/QGvdQ8pV4f7Wc1ZUy1wWmQJFir1+gy5k5ZZCwwo0/tPu39dnA17QedLP
hKr0CIUqBcvO4IYm3FV8yG+1r4PeFcopWGDKAEM0QoExaypc7ZXSTStVTzRLpe5T
X0oKMj/Uxny2d/+bAqRXB8bFTqA4KPKavLDp63XbcGfq/DVDdXCfs5AoSPIz5Ugx
7LS1aj5pMStYYasTIUGeVyVnL+GcGFdTggxC9o7hOLIfNdiauXauI8tbcOT1DQDF
A9xEVQTsLr7/2HVbf4kdPA8OxLF+VpwSN6bJhX3zdBLI5YtADMPTlrJRsc9/a60W
9hZLGQ3+bVWXfFgd6AFByFR5SIr/mdbqImnld5O9o3qkDxNZqKcYYE3RFC/DaZXH
XNktjoFEGX4Uqv4kZaeOUS3g7QKLSZrlzRWUqY04KniclNc5BcQxqSzIwM8/9HJg
+7Q6mR9aosob4Wof9lLmgnmQgZfFTJm+k5PJ6u6qIGSa+KaVZPFe4Sf1SYazrbmj
17zGHumQqfVXCKO3B1InzywsieAW40E896a08kbe+axkb5I7q58iQFbaExDBsBz3
9jqoK02BqhbfPLvKuPGCmjH6V2tofOPx4vx8BvroE06vMadTP9lOVGyPIiMq6dCZ
jTpH4GnwLWI2zNi3G7Y9CQPejQL1ZjX7Jh5tqkqNrBnMjxwGue5IXaCvz9oKugxy
viAH6dLNnRR4VT8XE8GLnV8Y9I7jOi1iDnJdB3Z5ZIwqgpMsQD+iZfdK/6IxHnzy
h1iBNKslNl1TWU4qcQb4221hfx/AhdmeOannmCHVC9v7AixxNQEdk6ihiYLrJP5V
zfDuwy28kYG7eGUPqata4ZzoXYkvRt9LSPEZKZrP44Ai9R+LCVaN2e+8nTWDMPZw
KDujH/jKh0OmuH28TLSPqhSx3MB/SN/X/HDTsyziiNHLbhi6UCEkyubzX2A1Fv6F
DeOcWpbDsfZEYMqD7TspukBuEAUEpYRp8s+NEroqIawT8HZUSOVEnJBh2VoW7QfW
J385nc9dpM1VxYyy3IAJ5tGwf3Iz08Ynt+PQmDbuHjdYUKu/GQPPTmDvt4SoG4DL
9SoZGBvbDtt7WYDCpTjrPhymAv3EaNzUfU83C9Upg4eSlDMq1/tQXhJowWxMFXjZ
9Co02u4iRAwG439SJxzmTchKNw1vfCJyabiKjngruNXf/48LK/hsGCvShEusrrIa
qRIo/ZVWlBGFSaq8CGxu6mxYdSGgbZZXyZreKYHlOxMy69PfSGwupR8WKDQ8fosR
kCGJW7zsdakQ3J/tWU2TQc7NhK18PQL6k4h3MbrVaOcg3G+eJx99v5oICdqHZnjI
l+u5EyRoeR03TUJLGsu45Wl6UOHVGgK/gmbY810hbOqdY9GuC22NIHbN2VXCu7lM
D/Tk48YOR3ui8qOjIMAauHcQFCir4s8JX+I9azmxmGPGN8G4zLZ8C1R3LuYB8AHQ
1aErLRMFspnBfLoTkoikKVKsaN9v+Qlng3AbSvQF8fIqPaphb0VryzpKbotHY+98
kpIIZqtILUpVWdcw9pe9ILuqtW057kQGKnrw4AKQWYqj3G3xt063EC8He04VXDLx
EMGnDvPjmlmKUAy5XREWtBUdhWm8Ynz+ct2nNTTYBiSuq7v2vOg+MPa3GKN+8+wr
XkUBghC8xK2MP36LlylhI7LBx+uu1fzmSnq029T3tXLWZBfN9kIdtF+UJb/rtqWs
fogzyEmxrignkvpl9wJQsYe8ArYnHtKG4lmvrNXpjfEc3ePq3JFxAra2tqhWKqyA
LtyU57zmE/pahddoyRE96Ha74aYnDmT1Taq26JVx43cHTATfErwm9LR9Dho4JH6c
I+DMW1PMMMnn8ie9lgoFW1qGXSi5JnWo+pz/IXanDTDKQSuGEro47x+Dst0rtn7g
jIzF6EC0Vc2PIYSb+zM0J4r5OC5XrMJdIfvOrD+lyAutsq2T+DEHu+nlUPaJE+1l
/h4v7rZBhgrO0BC0gh9LsOwxjSi2hZzK4s6WxS9pU4yFOhVCcpKr2Bhss5E0iODF
dYcbHecuPOeUt6teZ/+cd8v6kaRAkkJjZ4eGCrz0A1tA6HZz6zx3EdnMKPkK2quy
5gCTF4x2w0lKjqLbaeZmXtCH/qfh1u+ieQXJTryAfIdUQcSe91CuaqSLSBr+yK49
l0itRlzPfkOK+1ifhwRImhloO2DCbQbDt+pbJo5bwjnAb6yfj0Sux6BBQIBxTYVP
WoYzowVfGWyyt5qrTSD0dgfjYcO/P2QO5mE7coW0eWn/+MRiRQBb08gM20kYl4yI
+wRjLBj6WKj2r36hlIWHdg3KvPxKo+09F/K9PYqMziMsRT9wSj/f3ZcDLVGEBd0e
xaR+GsvfZwVghABLzmrPYH63o1T7WxpGH++DR0eJ1LqiYYXQFDQ83CApLlnDYLa/
UJ/wEetSJSFYZyaOqqlhBu51jBHK92YkoKYWScRkv57lTTEOA1fajmlsxUPpWR6v
QThg2HiqIeT5C8KgGLESISZQ/fB6K7CTZquZGtK6KzdOkFyTq0xa01FdYrGIc0V6
vwp8zFGNzhD4F/D0AOq4jU8wJEx8Dk9YA8o3DLJA/Y26nWMRCF9FefD2nvuo7qTm
XnU85wA16oC6UMrN7d9q7U+9GlZblQsQRBfnATeY2DROLi4QU988jt61V2CoilC+
KHMgWs24HtmigUXoFFoCqJ2b8RP+rvOxeN6hhZF8OhlrdFpy5Uw6dBp2JbYpPrK2
Efm8OfHqGLYq4/VvJYE+3gHXrb+rRQzM6wZydkO56McuGdcWhfIPvQGwX0erto5/
l+EK1jiLA/S5plFA1pU59SFNzsIIrLygUEfQm8oNwzsIumriuZLaGKgNfYIWOFqk
RxhyuNBJgvrlEt4TqAwTvla+fnXMk+LgRnmXKkwbMxCMtt6afmtuvWn+La1kg7nz
x1kvFKFvyvJWZJHlFIb8nm9rnNbWipU8X7W5DS7g8qp+0fQPKgko1iPbzwy/9Z3h
3C+cqlw52jczi1vfRFZSQjceHDM8ZmCZQObQxCXCTl7Vx7WZZKbf7G8ZMJthv0pz
Uqh5qvVlN2aVqF3Cp14XBNokokpGF60fv/cwtGvRI40icLgi4sT8ur5eu4GBjeSa
+B3DDGxwV+pPSGoRUqYKLujffL75oIeKYweZ6hMK78INb+Kfu8Tb7XCJA5C8Yemh
xRPoRdZKdn9c3qDjowBASmaxsrm4ZHGRKcZIiUi8vDJ9nl6az7R4tS5uLPYugODf
cxAEY8MrJqjlTaKsDoxr1g51WJeS+8GeWP7pXYDaB80iiuS8WSNHifa2ihYAGODx
dPCSTNIUL9Gjm9EQKXcJGhVfnKR+NRkiRFgLRIdrnjggm8oFjLaAR+EBRb8bVCtX
xt+C3wVk9g09Z7zG3QGGFL7ydNuk2lqcAb80FISXI0qP6wJqp5GKDXKFxOv1o5A/
qM/h0tnE6cG2GpSo+DMNv7lfRpRCaOq8IgHC71vbyoXcn5K3Opn6dUH3WuUahJI0
1HwUzwqdNWPgsubPYuqUMyKmtpWFDigpMbkGR1rgnvvx3Tb1+NNJTCLwwdFpSkmJ
6CSkSA/yUh7n0f/UEt/2FOb2T56/b8zaaju1EcaLzpxssYIZjMXH9EAb7SUkzQxe
j4oaRT/vbCTq2GDjNRyBH+99fE8L0qyKqdqwGygr8Ek094NAi9k5PXNxJp+oY3Xs
gyIUkbIUYOnG9i0L8NSXWibl8nK3bjYjo0bXhXmXRub5ifwV08ZjjaoJ6ljW6RnJ
OmvyeEW7ZDtCNAWbwXdKX6tFO/BrvrnCZT5W/Ejtt0CJcxfDMh2oK05gjWvO0gSg
1DQJIGVI8eznfQ8tVhb2jVJeUftRGZSg8aQTBaacaEPE1OJvko1RYuTDRObRek6A
j+YCSFfgzdH9zxAmuq9Oz2QxYRHOaQ0RXS+aIYwIjdqng2axlpJJ/Yus3kvjP7Cb
r/5rJtHDqOccb+4EakKi6Bx0KyfrHuCbsm+SI1+k2atu6uSVeR93zFH8DSOLFnd+
uFfQGCSFjV4l6glNE19jMzZJWvcMMkcpcL2/466UZzxJj0OwelG9fqFCO1ZpwLDz
ovILDrNGqmDbs4y32zrsjE2Stlqy2mUAu4wXkM8yLxu5adLdF9HDT2aNYkW/GKbX
yGnBgfSidtHDSTmmcyX80vjeSWWipN7NrAUQbmeidLI4lbGzRjpX12SeGdXD0eJq
qaWY1ltdCCJh4I4jHWVjm8v3B8W4Gekeks5Wf65blCC3FA9hHzmsAoWZQrslCKSw
+3PwfY12zmh0twJgxho1PgmtGCgLwJBvqsWYFpxix4BcWuX9kFkbR8pz25cYtXDA
9/RSUYEPalIGygwZ0yMa9CVj7U8SIP7OL3LxghFmK5JRs3e4P0gcEqmsO/gHvyTN
aadL9FDMcq48zGjLDtwE5CTXGwzib0BgbT3BivecasHIQT/f0xxlyzYGly33Q375
iURe4u9aZWIxturD1R6dxS/D04NH22z4OkPudBG7luJcK0ehvk0BlkGE9AiaYj31
E5jfyP0AJLUBJmcj/lTLJDlWqPrXDJ/iD4CJ5f8cHSYm6O1wzYvF7TwoXlmSKf/q
ncE3eYUYMyFGZCXFiyeHp3L9Y3+3EYGad7U2aUKw95k7tlZVOn4nuFuw5eJEY8Tx
2EInnyrbTbl2cW9KH0E+uqdarvDGjmv/hKwrlGcslualERUXkS08c0ASRJgTuxYM
gu+sctKxNqvZWi4URfqg9z/vZH8f2LR9yTe7jKYCF+0/LX0LRdnhf2l7Z4NvwW4F
0LUU3lNFi25YJopWyUj7ax2G8zWFmIyYIW2CJxo7uEhGh9J2uUABaSHSqMDw66NO
bFvsinaA2xNFzgZjQvUqvIv9O5EpVG9r023xxL3A2H32/16ZmmsU1x2Abh54G1Uw
GLeIaPxU3VtQZr8c+2fzIcafIAOrhz8N7R7EpHvPSIxIXcH010/wawVkdSE5600X
Mx5JwQRWV/lWOK0VYq+yjz8GX+VgzcPxOZAtqjFTwtdzu8EG2knKYo5ohlDiFtCn
IsQkQxVPNldXS5DSbgIKRK0yyoRrglgajWeuJLakoFckzJ3iR0eiN8KtLJz/99Pr
5Ll+vsuyNAPA2gKsDR0K2IbGc69+ji2zrktgeouvsJRnDqdgDqurVFeqYsns9hc9
FLLQ1UP+h8L4YQ75eVbcn8rhYy97mtkjoUWXUghTH4MHvdzNTVFhGibnZbx6NwoN
mQzk7mCByF1nBLPe0cuFj9YojadlEhsKZBFsIViZLhyZA4CdaLdDez0hZR2DYsHG
rZojuU1A0trIdrwSp4yef/8ec7g7K8Qc1TFJFY9cuESjoPoEXSkNLMC6tinf+BZU
6vGuJrA7JTSy3AK4Td9Rej55UzLwyBUSyWzKHVHe99WZ4bZ4axW2pXop2dHQTLRq
0T5r6R9BpSP58xKvpXRMf+RphgeXiX/JSxuj+HptZM+QAu/yjWyxmhldHpsqVvDm
d3ELmtesSv3Tn+QysxUiD0J5ExxaABacFur8WP5tQF2B4y0lIdpAY/iiFwzpz6Bi
mXokrHkfJAOL+FFPqVzB/DLVTg7Fdqq/zP85vsQ6Nzdxylx12nhXi6JX08/uyGF4
THE5UlA73R+OTvYAuoUbfckvtR3HGYf8hR5SkWD5xv10qcjZHusCoehm0ulR+eV1
w6NczK2H57hAQCS+/6FB0d+Ch31PrLFVLggCzzDu+z5fZgMqcin1+1qkoLrgy1g3
fVdwTR9RHdDCTnFH59LywawrJUAOeQMXMRz5ZSBuGXZ9CPOc0RN4XlnILWrss+Ln
6y4Whec4S+qfNx9VXcJ5AW1sQXMuCxHlsnwNaSbFpC/+GI76hTx97/kLisCXMtSu
yZ12z/irSBHQ6vgXcd8lcPutmY1+w2/coKxokf5Prl/okry7QlmBi3/XM2l4CM/L
dM07c5WedyFJghUICih4DpIIR1A3VXn9kfGJ9M+MwzwYa8q5wtrJrhfSXOwgNNQF
VV3LaDkc3OzzOdtdgvTKH/+nAJQmBItPCGzwaWoYtqCtcAJHx+u6/K1N2VL1b/uy
3oR6VTtoIeyswPotdRvWrB/V0NhQn+PqicpmE+eqV7XHV9RxZN3OT24YinbVqBFe
wwDSeqgbFnvRObqMPrSWaU9bvigIdo4YIiHXBa2yTmFCpWcHaKSN1fWBWQeeyp9U
yEuXVrXS6eBbagOJX+4pMuBFXd0jOrLcxrAJHEM/EFg94rZ9X/MOM9OCNxsuZrJA
2MqkevvhgwgElbXMZ5TtsF6I9Sk8T44lpqFPGy1nZfW8Fh+bUCic6Fia+tRBQOSN
gktzxdGBrCGgUl337UvePn/2ktMIIYwToFvvAzCYNtfQJoztXU7wksS2WAKBmlvL
BZ2u39J8L9x+Gi/jDAJd41FTwlRgbpQEHh+bQzJqqlLQgJSXNv7iV+760DGOL9sv
9fL0suN0LcGZQiMGkUqsuPPY98+AL7cuAbYlQ0h7AdDqASAlkZbORWOFt3WTLORv
vSXGIWwmoeXLzqUJYbFPbVLGAiRzZ5/oP2iOLOAptRPrywqG/eqV0uCzLpuc/ikC
PLMIDh71FYGiXOt/C21pZ3Aoqk9bw7eQw/HnPVJmV3GO7/l/umy7YHYG+3yDi3So
Mx7aU9K6PQjo4WnUGTLxtJ9VhvxTYftLJATGegTFRefzvHVfuufj23R0ssI59T+6
LHw7fTC++49KR5AmandT3T72ltEASfMazEanSng6AxcdvnXRtMocQ57YDm/5JvEZ
x2gn5u81kQxtWZBJqjGJuNPSL89A+IX6Xxv21o6P/LWL9UH8cZCOoMsjzPB/Jkc3
4h53XSeUTJ7e4nZIHNm62Yi2BKI3/xZJO7pmWTwiM+9icS6nFpcQBaBzyP7r3GF6
XwdKmDgQl1n2uql2SOyChDY0fMjsIjBJNo9OlB5xg6dsVpZtDJPMs0nrFE1aUWW1
Zb6sX18a/XsY2kWMuMcEcTYMCmCgI9WyNy5yronGIv3hdKtXFZ9Z/4gFm9iYJfXI
+oAJpQIA7XkkvHJMCClRlj8mfRtpOTtXpPIlOavd6DDTFxFQs/q9oEIAKAVs7E+M
GjcZbFrF8vyIRM0s8UjWokctszWzVMxEbWKHODiw3EEFK4YBkvzy5aA/Lhdy/JBi
j+IONjZ43hSDBdqu4rlLehEWNoudN6DNysUehmJ5uhP8omxyJBBnidfLe7d9sRXA
qei93icoQE2ovnq/XbIQ+2XSSMDb+g6Pg6405KE9uB70ze5cxhlDv+vRk6EjWYys
JQQK+z8CadT+X9qL1rCVb6jPuLJ5nfUmLMzxlv41XPN2uij0MYU3L6vgEIiNSl1Z
dVdMZNKVjJrymkQMfJl2TPYoBXRBNsZxvgd+2LGc0lkAyc9UugfODDiLOcLuma+B
+ld4okDdqwc9H9zhxCZXiAKXev8KG039RHhG70bPMB5vyyQ546+Vtw+IE4zqYpOw
80q/EKn4WdCYIFAyAzpWSV5yRFcWuB4XYpWSDfV4gIs56PhV33bLIQslv3swe4+d
c3JbaCQ0hH9iUDt4Divc8Q8MQo2QI7n++JLjYN22VaGAb0Y6HVXNIbKeiRyGaHoL
7SOtE3+DPcn7C056TPI4Y1t0UT0DzAVTvedxOLxJ6ANy2BI6+N4nlUldIzFU3FVh
jgowQ8UT+ejvE9eaZJL7N2VHe5X4NKCYtzUjWEdhq/jRwB8vipMuJfnhuy/IqpZ4
a18l/ZAzouRnQm1twSbUmdZMBif+VwlL480Jqq4BJzHZmtmvnWtHkTMWMIR0UpGg
Xngedr0MJgkdFwZCjIMf8RG8mRbKhkyf7/oDxAI8yfBQ73EfBGMXP1BU3prU6zT0
FgnHCIxyc1lvdiS4kZ9LlAns/2rhD04uOfWVNGhOAbHoBySlfD/jnDTrZ4hyhox6
dnI5weuf+aBXWgrZnpzAmmjBj8LZTBA7VnEJIrwagNFZLIhoRS5hXff5NN+EKBac
KixkQLabbtO0ZCvcqH29OH0zdp1d4jfUoj9sxIx1T9EmtCBkOYU/xDAgZuZ//bM8
KzcYNXVd/ilXD6GOaJqAEbVmguv8WylHHHDQEdCMiANkWSf8P0gD/kesNQ527Ysr
2SvMkBl7EOPLf7BIiFL5QbAfRqnF5GngBm6xK9B8kNgb8FBiEX9r4sSItse7LdLd
2g8HgwRj1+h3Eru6iZpGsIB4xadiuqoodv831ex10O4s8MGvuvy72XcrulDYccD3
neM49WcikkHw9p7g682xmLFk61gp2GZezO95jzBrLZH1dm7wDcVvDbEQ3jK+wObY
I48+3rNTap6dBbc4EH4TSYl5qT4ez7Xn9DTqmJDg6P3TvvTG3wv23LlsIeUXhNrg
0I7kvqLin1DdUPnTiVE7dRja9ddxPA1q+tWMmDPhbfN99axZ3OhCmOYVUUkDRXya
BdcXemxiCu12aPu8GpZ5gjmEDve87eLkzE9ZZny2FkE9FMQ9KRQnxH/dapK7ZfrA
6wtl5vqISa1VDEqCYQTL4/B0SujYPO1vi7J/xN/eLjRGqgrcAcfoqu+Rcgadbths
sea2sZc47+jZTrMJ+ZMSmqo/xUYiP3SyXHr+jbDILr5xf16Nytv+gDrZnG9N5+Uz
AYd9XhuEyak2iO2pplA25Gcvt4XmCYJbj6seDadsVnE/0twRjiBUunXihyt4Mb5Q
1KC8B/9Hpc4w8zwX+Sm4F8gwOJasL2TRVeTwTa1TtPq24pufgMV8Gt6Iq/hioy6v
h0w/uE9b0bSHDwrTDHNcbmPtvHV+FZ8sJeEBIZizLZtTep4keKiRdI1tses/qH0U
f4OaNUBiWDImm6BbWEXlfVLOJgDKBFtJ1OO0j8fd8iY1agZj3P41ozNWwS2XbJrD
Pa2PFuhx2nCy4G2ltNdLlwYTrQfih7dMsqEzGnD+i39XmmGD851/Oi/ilgV3vRI1
zTez20iwQalajfBEqcIvU3Ku447FBUybZC879Evf5svrPd8sEx3a0y9ah+/VXsrq
QtTDiQ1mgHaJ00boATSuG1A42W7iWiSQh7qcu7xzjb7P3O/B7y6Ph+h+jXpmhyRE
PgOgr4QNWcMLOLE4cQ1RAUiH0g6dnPkOI7TKGFCfqXz+BWBXOA5G4DctUuvidoN3
Yto++g+jtmYd5Ni/D6e3kYifa295yPNZYS5o90kbK0Nj/VlhKhUNNJIz+kVRBtjG
9AQ+ekwDxXNNQ/jBPB5E1bQFiDKkoFQHDPjoq37ijUgnHytfnCnI5UHjXRcD7Z1G
XFV4Gu0ipL9OWRZYMvMzQsWZY3dhn3AX+I3TC/JBpcRT5sTiH0/r/KV6MNTEfkrG
c8PzYjxvmT73EpM38qyNQA/mxcNxBJNn/Bwmb2NC+4J76P4ytNgxFqX0Wqv/DZH7
c4vwtmT/I58u/r8urthEg5yRUB0hXvqRvpG+r8PK5pNPcXC9HbZ9GdGPGRWnmjuX
AouBU+LDbuTt3Q2oDMN/368xZdBA/e9NU/sS5iTebSxoS6XNo/siDexNyA4d0RJY
bsaeq1vHqB93YLYmmd6wVsUXLA4DSjVvBHG0k0+fsTU5o9ggeW9Gcr52317cc7KV
mGZJTl2yOsm3/OW7vAjYGrBRaAbA6AFhBEHXrEkKM1zrw1ObJz4TrvEk6WTvT4ZL
mfIq/6dsY0rJy7YF0k5tVBfgmwNV+D38617k0Xgabz/Hr3j8M4YW3Q+65ZKJ70Ww
o1VFm+tFqjiZhVkYtypn1aVK4VVPSO6pwEBczYXwRTApyU4M1UAFfzbP7ld45ixQ
UzazlnyXbIjus9K5sbo1q5NgLRCIrFjNOr1+ymjKDC4g6uzbx6xj78rrxdpnH7+x
U4W39g0t6ai2tOINwZCLK6oFoqHkcRRuBGgPjr12zFKEDnZj/tBhaho1kK0ue8rE
h/LqtMHBIhHwyFbJmGrQG3ZOXZBweBZybrodCxQqB2WLncFZc/UHjvpq9H9S2q97
hVkJvT8HpeVBt+ZWY4ytLrqYqXO0DbWhGq6pApiqCmuGvbzDmVngrAS5D08qruNU
Z4sCl33wRRT08bOnbC+9BoTZm0qD3elJxwsDgrk4RQh+QKztSYbKuwyYHwi20WPc
iEFBDz4+cS077SfJM/XwSTMqmc2RS8QD18XeBCsrM0cQ0/t+4NfcCbh/4MTChNjc
lnm+M7nAfZKeofYVwWBQm+Q0n5OyAQXKbwcmznkviqy/GLctDK0uM7BaIm6VTo7Q
wWMAMM3hHsEpf+L0aVAdW+mO7CoOa+hisckixTvTYHLP4iOGqvkZxauDkXvnX/sU
ky5flyKD6GQldXTdECpkb5ZinhIaDcQN0i8RDZttjAHXKdnYBXBZWx2uF6nlzDL2
QJrUPh3DP2KHSvoDnVaHHaDkIqMNvjSCPOAEEZwdPYfXJdBJXGF9s5WSKFc/3ezG
v5jSzhqd+0o/BlE6M89jZO02Bkuiuadg+aXqs1umCtP/nkzOfpsJ49S+Bu3rXzda
NT2xPZ1jXPbbh6CW5vY3Z3EuES1X5E90alpVRRphox3iDeqeod02pGFyXkJkPGHx
dqcWYNNqQnrSn9irCClCecekGov7HgIPMIj4Rh7ssaFQ8EnJb4vx4aeHZVMntcrE
q9tF5+Utc/6RC7KDOxuGqb5nRIZrTXeQ5q0iekt3yMA5LLeQ3Tgvvd9o9OJPnNxx
BmzObLQQrYL/e9XohAqjvQgnQblR1Mo+sEJmlF37CmYOMbdDgWNf+g9jGWzMjQAz
Rsjl8XkxDRqVcEdHIlxlFniEer6gwYLClcG9yNzkvEVt89ffie5hJS887R7yd4ww
U1StlEpBOTOvuOfRe87s2KxHxAPo+ogFuI9kg5GF2LOTBGKByvwKK6JhqwZU0KmZ
EbI9cZdEmM3JIdFZPa72KcsKUgkxrCSDZrEXuMfR/t1JRYPwK0l0ali29PUl3aPU
LCX29Mb6ByYzWHECoWVDWStnQ98kHM0aWNxvvcLXUWhuSnSPAY3b/8DVYGhH+r7i
pMqxgZEnt3eGf4HKqMylIbRt+iB5k4vUBLxX49kth7XJ2IC0tLJAwbT9tJyhNo/z
JM/oC5K/bjZR0gU5euzDTBLXg+pb2IMFJendhtT5S5JLF2LnSzrTc6BKER7Wk3Lj
wLbijeSAf2NTz8AFb3Iu3av1WVhtv4fsxEj5e1acQeFmPSti9+NzKxY6bhIHKg5+
fjVzRmmjHa6cGLRcx/SA7j7I4g+4pO+cVHXdgo/9UVMYhK2Iv3FBlmhqcKEMRBm5
XCvcTN48nLuBqB+voLicbXVVYBHXEuGKhsCfJFeDoedbhP6lxIMsapFE2bAYHpod
FsVYzDF51xUy5PgDrSBOI74sEnvlUvhcwNMqM3FwTwuIfoxcMy/dZhLW5xjgZ2Kz
FDsTeszAva36BXDZPjT57Ywnqv3jmGFtiubgC+TQA2pC4QLGxIwfpWhbyzQr148b
tfTLs1NHLVmy/ziDAV4TywVIlzuL/k3fF2as12yzsYC5o9W+A8MjAPm06Dw5/YTm
CrbWL9A1od8j5Ej/PVB9DpP8pME2coC3Klb+Q6ZSTvZ+g8Rd41e+BcOLxtUFn86e
/LRwHud6qElc5TgIL6vFkxy0wqhURKLe7S8jjBOBYoTg2DHz20nk6gGEqN+KFzAO
TY6hySZKhC1mCd3MCDM0I28opEog2xJBatEz1t8YMH462C+jQgJG766IgI2DBr6U
vlkQjAAL4Mro1QodQWG3/jRAUeeHdTu9CNm+FeD/lHfI6/94aBz+ja8HuvN57Nnl
YoBNQ0+THQb1BnSeLyjy3DpkiqaTzcg6/3Rmjaj8cnAaNl6ifPzPwGzTVbwUb01A
ZKlAOpnWUYlH7Tw+RBhZUIN4/kO7n3hh/Ft8Mz2/1O/4uFVbYa/TYUxV0o/DxA0C
GTcoGZsOv1NZ1OPnPbfgEkh3QnPNB8nR3n178e2ZR9gUCqIB9tr1Pd65MeP5w6LU
rX3zuG/XGSAeU9um5cmS4JQoBIefxsAjZEusZbDxQmRxfLWXe0m39idciLwSxwvV
BmU+bFIT5Pzu3SWyc8UYVfkf6v4ekC1ixPdI4hB5MS3QC+T5BvZdywbRUnnPnyyI
1Hi0cznJOi/E3C1/DYq1Q7IyuAj2x2fswGvNEsFzt3Qj4uQweorGZWiWdm/FTxng
dRddkvETmmfd3/XO63P9Ki9qicNsALP9c0KK2Un8FwyIchZOTgM4v70ds/Qnlhzy
0pbUndWtYsfqUPg5B3N+ZRn0WDx0WImZl4CEdZIwOyCaxdQEv+DHBX3kFFod2DkS
ItuX7YIUmF3pHtvX6ANWvRiwXl2OoK7NBik/dEKhSYG66L6sIS50F/cFi+aCgDKG
bb/TAlrzGZ02svuUNIZsJjgKb5qdydFP0p3pDb32SIQCfGS0VoWD5pygK9DN9csj
gcdE8m0Y7dtNoO4xK8PgY0Xp7Ggiwu8/oOByh0ALJU9BfpxH9gUkKMxvJpLb0iYD
GQIquYDW4sZUbR6r0GkSyxBOaOtuWRkZpOZFw5kxC0EmOf3fcEbDLWv3XMp6MjQK
dePwLcHIYBeGexw0HGsVkbMInB9oEAgJlGDCa0AXFeysiBz4i1X166hZ/9inlsBc
VhZYwNm6y1Ga4dffI+r7TeUuYG5SADQcOKIwrwEbHR87cZoaTbcI+hiq20bo9DPB
spZOAu9qzEhRIRH+JBgjgEnNs6Vg1EWWia3QgfyXJBS08YJldScUPXeOATRVlBn7
dQrvTZ7Yl0qjD/CbIjMBpEQT/a3grzOCFevIAdbOktOYeqgIZmkC3Yk9j36laLxg
sIGO9lkVq5k4mjAlLhAz7jJNGXPjnuVrK5etH+EX2v7eSXfQ20+Owg5Lj8r2OpMy
n4TsYGhdItH621/BQwIuKRScipNw8DtnjY9FaAw4RbZFKg2OVNB7m/MFqQI6rXlC
Q6sEoUDnPNApk2ujXvRbI9mF9vPD4vCB2tEvnATxfnCfkYl5CDGS0UcXdbNuV5OZ
c/GvqFanHAqDEObzqRkK3fgf57URUq6Jq+gzgBfReE9lxkzfYJuwKvDx4ZW2Vs4N
G6uc02+1V7oSco3Ob5XP9r1A/1XPKtOzxr6txqTIPRzjHKexR2cVfGaHCvqrrlNK
IqwbsoCD4Ck/PgJsgHWuvlaZdV2RWb6Elug7g8CRGRvRxXB72mvUHl3tACSKWsk0
DJT66B1yLG4iV/IyYdpKPMYD/r5xPKYACrbIY33l+TVLXxeVX5qifg/Mf0BJTCSo
cPFQg+damyXoerhBUqiF5eNtM2XOFG7QpMu5bnWiprTDMF64Tvr22SEdjQVRLCIH
BiVHPkFiaUOb7zEdFcUjPW1eG0JYgJMQB6ZQtZ1WayPjOILaHZ58KmE4PGlBtwON
IslwQFDHSPVlj93l2hSalxB4n+35A0pqeRt0jjqWBESZ8ZUlw6Qd53F+380dem+V
dYDd3gPw3qYE61LHcBFbQh0DAahw1Pc6M8CAuOVhCH1bpI6RsGcRRlCeNYL7Y51I
fY1j7TtMM4mqOGgdYtVwKcrLft1Sh8+0eoPfAsYHyYrOuhf53eJ5dqkC8yIPtfAd
+F2RfSRt2jSSxpbO9rEz3zl7Ja5N6I7VL+kIvAmDnrrXQ/33IjfGQioygB9pRsCr
UMIDFVbyXkJcKUTEdNXSB5RZgRun6OE6lGVF0HqMJOxFX4iaNvDEQZqkUkgR0vTP
nGW1RuHO8J9hjkVpVN7hNRTH6rlYXUllGwtIbl3j1sI3KV9n2UhfeZ18hhcpoOy1
S5z9fZ4DRtSmjt09N8zUSjo4ddbake76F+ENJXK6tI3mMhkvbgkcGLmUBLcxw1XA
/QbgyTAqwzH/Eqz5Ov8ZcGry+cNwCjK+hBMyuU6+th19CRSGAFX2xZsSIfk5Ft9s
rkARAN5eiXFPteI8uC/lRYCJ2tF9llag2Ubasd0kDPgP0Z00VRhauroQYN4OU6GK
8AZ4iIUqxFpKYoGC+XX2RKdArnvNcFvkCp4evwXc9aOdqDEN1y8NpzuC9ixJKb0V
c2fx7ppn74TxR0LlYvONcSZY1/S+ravXnb5W9L5sxUcRDB+TY8u1OD/K5HopO+3M
CGU/R0qzQiObd+wo0tfHeTCTWkosbi9vo/otN/zqwEaEb1Js42cGRDv6Cdu3VOxV
pZQ3EmLnN+b99BfdE0m+ZR1wbJqKGw+zVJCqfzwnu84t+MeS3tX08qq0sNH/fyu5
WfkNeQOQioCbVrBXEMoRuQJIO37KQJUKTavn/YoFfrKGZWKKyrRCjYc95s7gQr4i
aOzrUcUbi1XAlNJVDq7l5dDydSlElWBSZfNfTnqQRi+0YzfsdNGRyP5PjoXmD644
Drzrm/8WBZ0CjPAYKFAvMEKwLVKhYdpigmdEY6LSZsKKtlrPuj8fIeMM8n1T0xPI
elTOCy2ubzwYPG72w4JjFXJAjFeQObPCqJAdfpDI7T6Wjio3Oeg/TlYHZenXaaAl
YYUSzXWtVTouFsT1nt8JnwFQljVnuPDR5EW4ULbYY5/Cm/3nkVjxqYizfiQq6vAL
0paNoCX3Wl4PBxZqYNQeq0k7R6jGqnvqXJS+EtV6TiGEDJCMT+qrqvFccd5RKWi2
1DKRCFVOA4ScSY2EkO2kNduh5daCUCYt+ykZuPsV7LhNaNQTsfiRq7m9dkjJXxR+
sy7Ieaktx1em+mIO/YAtirfZWm7F2dbQUnvGaHBrvQ9A0fZZKhpZyyD+Uivle4hn
X0nzTFbMj4BuXPIKlARN5PGS9+LAudTgNvk+IB4D6yy0F7UDn79W41i8dLLmx4OZ
w5SgB/iTneUBsMiadjnUcm26meofDlqaylnDPaAo39jhNANatXlX2C1f9TrcgRjV
aqxtQQMpm9h9Bzok31XY5HtcsO22AhfmqV1nL4p9Fe1ENeMlS1CpkagWs9ArZWq9
QJI2qLiLoigYrox4RHfP29idW8bOyX2nuut64pYqTFoJMkvBOtUiapIY8jU6oqB6
iIISd5Bn4aqn8eGBxNNPQO8zTfJzhMzy/cHo+3Upu4qonyvCjd02xhF4jcQFEiSj
QAgEQay/WQHrCfPLa4hV2as/ioTLKBeex6eoYKP4YZxzzm5v3rKF/JseDeWl8Mxx
j0Cp66zawJOk/6nYGX9+qzTGsqdy/yxHlhxPni5q60OpTsE7+dJUB1jF65VbFnLD
UkDMxt17wbfYq6oWTA5oYXeAlWspvmLqVXqKHvmu89xvTakA40f9P3AqMqZz7MOA
5lo9aVHFAo8uXC41vfHI4wubjTQHthgRHd9isgrDu9btndX/lgn0VEDYh80DntHV
YuN1qPLhzx0vckb4iuyAKd3RYhjtwHMMzTBpCOO91mmi2miu4CccJfNpT7DV1MMI
X1wsAOO7Ir2NLnooPardnPGY+SQ2wKiW0lzzjbXb+5CD6//ZGWnkyIyXr2Yn3jWh
DOs4t8+5uiIxj+p4coOWFcLDAkHzvAoxQ5Dl/S3/AvVD1viW1g+SrV2+RauDDm7+
aXIRPyg3Gag1Swzjgwd4eOLAqdpZ/lK37rL56C8OzLc9FuUxRnR/qNUfSz0/HU1l
tJscN13u3vOp3YaRs6u3LLTeXcCDFeEd/ZZ4vpALAIIEPNCJKVPMV6DMglX3AtxJ
WvPHvI0FsSmRgF/PgHyPY1Kgb9nWjFdDnz6fF1Vjs9m1yBG/U6OLgCCqtbtfNl4H
YnCebU6HnLjQNyZKROM6R12aemU/WCWp9kgVC4/f5dcHwxys9ziKdnxKYxnotRSR
StoXpA5HLjIV0OHOX882TX2lftZITSQhTZfzoo5NfeUDcvoSq4okLaIr11vu68eB
/N18ZUdsdV8+tmJKEUQTBecBlhjzRaVzy/m3/8oW5UGG3jg6n3Sd4KlG0IPcfJsF
aFnv9LIk4Fug7zFGNnNMSyU548FF3SOMlYw01p25meSKmF4VAgWroBszTRPUPocz
EqXKRVAFh8MyqkQB+QzozaSlgGVBwB8ahEzMWe+Nnw0PX+ertC4EWU1txrI9gKQt
P6Lh6tw9U3ImJUKZyVAJUB646oBsz2fvIFbyIj3IjLnziY3EF74YAO2tsH8GJPyn
8tx1nptP5W8oLuimbxDSUBnkb1Kg2/8LcpMp1bKrzZkooynBRuNGIqsxLi4OfBrH
7UInWYgixt4JSybZeu3OlSS+Kb2CWMsNt1/nVNN5HQ5lB/7QXotahTlsevZ6vJl0
GuH3/Uc422mk00LNTLBE4mySFne94eNjvnRdI9tZ8nNRCtiUMDeNX/HxYIqe43Bv
7uq02jD9ADajve05LoBR2owTX3+lNXZDAJ0zKnD6ZW7+Fl4NDFwWJ41NDw7HM5mn
Jzj71sknZx3G3KivFAxrMG6iwJnGDREwelDh1yMgDf5mjkA/mOUM1/nYOKOvCfRM
v3aIIRA+m0KY6IcROtQ/YfUsYkp4XiCQ5qgCER4+NtJnrJQ/X+XCsUhmRREFYbKk
u6C2/a03wSBqdhb3rhblqGca28hZNVYB8PRzQGc+D5mKn2RT3zjEZSKforp0mBDv
Ihu3b2nhkmC5HKGYNOwAsQ5Q5iV+a7QLCC0ickeLNZohaqw36BFRkIMB8LZ6SD7A
hWqA22DDyX49uBsvs7COOyI3BB+HsVtyEKIwAU4SOPGtg2KbbM3U3rFAbXLKLjlu
XRKavuzYs3gwpHPttzzguNzMaj52aMNWrftB7b1Bndy7hu6BM8+fBaAimlo9I7V8
UfVpCEbeHg5ifq5VTu778kjC7TJAzWPGzn5eDOWhWC1bNIZcF0v9jpUY5uAxAhaT
j6jLEvGqpy7s05skUpeKdR83u+h9zI0mdjrzO+p+YwlOYfPIvXXSvM+JvNuNO3+M
lXg6SRJVReRfXUUY6DVvzlj3I8iZvWtUQuY7GBAh1jlSZ0mK/8q9paAsx/nFJEWV
gA5enYmNuoDPUH9qpN3rK1+HWLa2oNkmojnNej2BF/OlJW+V7WbaZhAio50d06AE
91SrULaCEfEvd+P1yIhQnFW0+UV+6oDNyoMp2Efjk6m8UUvG+rDu83ZnADyNkFxk
sk6+6EevhCl1Q1gyI8vF3VCT/tQcRDdj0lW1sFUnVANpRC9klm8kt9pl2J4VFDFA
C7UuTQdx7OCUQRGbsY89TAhCB9HUe6QedUGIEMeTofJ+JSyrvSCLgWtyqR6Q5qQq
y7ZUC3aPfO75ytMIh8417eJaU1/oTJWYtQtjdLPjhBkm0AKkJBMrpkJQVJCvzMeW
KkrWxDD7oQYPTlPQZIxfw0LF51XpVg4vQscZKj3L316ODgt1r3ihwTDneL9s6gJ7
N8CUYDL60e81NbZyqog1aMF6VDKJQ0WemiMXXQh0eO35o3UuSeBn91beyhS0Bapc
VcznCDYOYml2bYB5z/sa6IsZ9X6DlWZAbRCfjVEPxbTHuPj9LGmRuURzfdfqewer
a8kTKEK72HNzjY0OwF4zR4RNDN+WZGLlXbFZihuq4OEcS+7nXrZaIp/qYRHekgRt
bZAdm7+7d+R8GwdWQ1cDSzHyKsD18hImX0G79Fvu/Jn1S/e5ccMox0T4xfPqBuMu
okxz9CfkzUcm0glwpn/1C+5az38bjY3/Usu63Q1sqsBrgTRkd4alRqagvQwUoWvn
FbyOiKgT5Ek9We++PLWJt/TL4qRtBMQ1DTTiAwXW7vbp+9V1Wpvc++Rh7gsKzLlh
uFLW+rXv+pT6RLvqZ8rDNCBLnBrfXcwbY+v0ovmAN5DIT5VlZlI721GDjyKgvjhI
8K5xTaQL+RSx1JUYDEuRshScxR3zwjIptOiq6N5C5DDJ17+tUE9FO/Cd3OD0jD/A
bLAFpqQlNw+o9CesrP8Vlz9bqeJBAbXlMFTF0RoNiledPxHJ8suD6QmCgIttEJau
nfBj1hCvASeXEiuufpNpK1Lo3pptDpDq+EaOQJxYaKUV5rfOmoEMV22kniMLsOuQ
CWvPQhrAfBH7ZjHVcL+1+yqmkAv6zCRS5KVWU3kZJu43ZyhyDJKDjutgmXe+fsUG
i9AzshvnKY0FQWJhAaz/m+SVBbwkloyCAMfEYRqrdPh0Kbh8A6c/S/dBZac8D99W
z/2CUHIhhGKOhKak9qSZfnWnKFwzcHC+vW+TpwGd8EEZPwn9Uevfl+ZvtRJCk2Fv
FjSMCbwfdz6/tc9b7YVMxknR4pRVgGG7qx90NG8gtLUj1QALzM+KjfWmhZ7nMLWM
DtWytSFp6qn3zz2wTM5OHnw9tTVJq/v9n5xhTh3XlHQV0w+MeFeFySTjPSM+X4cd
eMXr/pEHXr/rMYczFOOFxg+ns6H+fJAOns0E/P8yXwqjcGInDNV54VfKGtsp2kAV
tSrBJ2R9oSFDCJ321Vwiw3ESzNFl7cJRGzESGgAjkBgTzyZeOhum+9yTP73Yv+bG
8tlpen9hAPp2pGEC0+94XL1hdo82VzV8ywSY5XTmLhdc6LQ2bgYloidYtF1AOs6I
LIXPKY6vrr92gwNoKMsV7wXfwUhnL0qng9/KrAWH8n83ZVum0ZAiCKXXeQZ5guwC
WCdxggaWyqkFFoHMUFfgIz/lOLN8gIW/1sTDir8MtyE0pWHU8wihnLC7BPZvDWgp
rfj8jPEkG9BFwT2fM7ofLmTS+a6rHRZm7ywxk92Y127/LULm+XCgToTVKdrbi+sG
9JBUMs1nNWprIiPizJTjYF/bCBnT7oUeThnFUg78jzMOM/8tQZYQJpk1oqyGxThq
DA6QJ8680dy2WoZGrlmvSyNrbAY0KXSlgqA8zamqpcHT0XQ3zKBIRg+tQt1P//oy
hpBa/BK8jonmfIYYzUIYq7GHCMV7eW6SdzUxCJkixbj2NTkfEm62jH6xLe76pHDd
67IOSNlNDYw7dCamzdUAzedWCjni3tGoASrW881klj6ePUc5t9vL7nFJGDTgeXcn
ZKEG/N/2Hdm92hf7KdcxuOpp1lceCyX2+iCvusjwKCSt96BncaLxrAlPVdNGxGxX
NPTsbb0PJbmkZ7uz7w+okD0Fp8SIvzT5yCF68ggDYCmdOpMXqnu2q/FUqk0gxvSk
ZcYYdynX3UgJFJ8VZKdYchQoh2Op4ucRuGMl61ZumiclN6dnikxIZrlOLBi1rr08
hJ2YjASCFJT5YoEopNP4Gz5nFAxwjn/u8ScPlyCSykVUFBT21upJisG6sKwKNojs
cVRoWctQFtdi3nDQRs/yxAdq2OjsAu5kHCeJOTqZ67qZOCWRzxpBLxWStpUnUcf9
npGcXDEmHXH+Qx9cSTDoa57EVRca4EqidyMwgoRxPZylcAgGX1xL75h8B3tn8sCw
qal2wtdRg7ZvxqbUHY9UaIK6+NXt4gJS4aB406KY0tFBYJnPJGtRsyyNE6T3M2NF
aKVIabfaaPPEOz9yaMgLIvGTBxeRYvMXsWfird8siLKJv7mbgif4+M9MBWpMaCw+
AwK71dYN/6lRBu+ZhjYC217D/w8IhvnhL+Rlmnc1mwuIwYR8ewSmY+FxuEuYQacl
TwY0qVXzG42toIphW48SnPTopihAOob99Ji/aIL35+Az+Fny2I7OiWSVuTgW4L6p
2KGS2RsXi+YwvLaxvluANM+r3thJh6woAbQTJ8s1KFCczTd7yaWS1OGMSfRqtA0i
Q7MEdq/ydmuIo4LNlo5Gs3Ofw5mU/iuu5eC+eVN83wVJHC9UZy1aJtwCxSPmFep6
es3+6pvEo+XQBJDVzd+PuQYEE5YjMaSjnjrmq7Wa2n/XoVEwiFoJSExFHrxfyTkh
Qe5pfx9ndRS2497JzPuwwvAe4mLt6G7qDjUZ27+/xgqbJgjffEjdrubZaYOZrIOJ
HLHqBqA6hKBAPyvWEaIiCCN694DG92zDSeogbSSTzQnCUtdMOWFQ5rZ2ryopNdHI
Pib7EJgCbE2SaH1eR/9x7SDMDlAysP+AREGyTsxAycKseE3+mwmTCWB75hvAizYn
EfHDtam9CeBMDGKtkBIS9pARrXyxc7m+rohxqyBzrGnrq9P5bpzPz0eWgKL7p7ie
9iDP2Fwp0BaY/0j+SvtIXYpYQIUrr3x6I/OM2uYsKkFvJKBY4ZjTRlb/fhOiN46t
JJEi5jdY1UBhM4IFLrhiH4YbI/lP5PdXD9NUzJKiAvllIYcBT82LV8AEbrqEM9wv
QSnOEvn7O08MHB0J9xg6oZQtWh7odX3dF70OWUHOH4qwaY74VzsHk2jelrXsL1+/
WZ1/WToZIqQdvXW2tpLAGnKhJOA7YoF86JxGzxWnajo5J3ufbEweSaRq8tnI3ZMe
E0Uzg5ui70/WH78L1wCRpX66xmCfQxu7O2nHL4fEtjMiaasdoNpuE3UuxmUa5Utp
Lq2FsfuDniDCA7r9y8wx9HXZAg5CeJVcXVQdLcMF/Hyt7gc98fTFKqKOo2UPa9u3
wrI0y2tR8qSF8UB0h7qDkNqpOftnag5l2tHexbUqZHUEV+3jgHyKdsemdOw2z6Yd
Zbu+7vhpCibFP5nSMbdF1xOpWSbeuRA54jJMyJNhi2ir+M9ebJCSjP9wQxn30y0F
XniusdfR7z4PpXSY21JUMljDX/6M2Rdz3vjgWlyJLY3h7DUEaQq0lGkU5Vq4y/qq
ow/rQKz5Wy/+oqlzBBFT9T0MrM/5YinGcZtmpKGR8nsBOS6bMMMs4jJ+o7Cdob1y
V0fGgOeJJ8Rh4iNIHiCJNFwuivlNsE3OoZM8dYEDiLVp4H+7XP7rUqesZdyLkCat
fgpy6enO0COtUJKTI1ylx5xwVk0KVPg1qEueRhXFWLYv2U6AzV8IFjj7X/9jXjSV
FmV1YkxRr/QSOQZOjnJb4ZucUCYB6x+8Jgg4evTMQYbSMp2Pd/BcC2KtW57xnWlq
HNv0zsyjxhduYC8BpkKNn1bgpdQrifUkLsvEC2QeSFhnlAY67KX1IPLkg54cE6ET
eRI3EJevbo8QHnrGSrZAkB7oHhyejy1+Hpl5/vSqxqT6jABMjT0J7N/92PWdo8kM
1ZuLf1jswIAklrl/Nzq6KT5L0l5xzHCZgKdQDelpG3WPhJLoVwm80FZnE0hsFHtu
upxo/FJFqb/O5xwxCO1kCVjpDRoJjphMDTJQeXhk1ndO365E13nQ1nvMhXGx21sT
Z3UUN45sZk/1oWrVL6Xjcr9/C0feWLQTcZiHjiBNsDx5oV4DaJXuP2iTT/Q75Mz8
w2YAmpP7OKfuDbmcRd2zRzNMcFiZTfVrv2lQGKUZp7yOcZEGGUX6HBIm93A4Xwrc
pVQlpS/jcmtm8Vvn2A/v3DPTh/aoiW4uk6seWys/FLACc4uyvryzOl/YzhaneMT6
3Maw3iLAKDgLchgCG54PDa9LOjxrENmLbRLwS4ipGHQswRXdqts+OFUrN6diGrFM
qgBv8eH33pVZ/m41G5Itdcxkyf+YipRbXbwcixqjcG42GhelWR9xDRElgKvQyxyv
oBj4xNY+SOY8+2gETHQEgcU4dt/d2lMHcpRZ47azHLKB0EG9n/7oX6u1ALyX6R/j
jHHmGu4A2ycfTzK8RhUF+Cj73fAN5GwqdRx4T4Sai+wWiqJVm3iUVr/gzAj1Khv4
Z2OUe2hJBXd/rvDSGLd5lTe0b/Ec76kSd9kduEj0LhxLgwpEo1Zsxi6O8C40llb0
MICaBBw0JTT+fV6rEG2wn6BVXvEJ41lz2uLUFjS/c84Vd2J6XZNS7yAmnu4EH38X
jtKjSMpW1+FVsTE+LbeLjYYWLzZnpzA9lBBZmLH6lux4rezRn7T6fXG5/RxyaNL4
4oiFNCChHJ7UUamNXGQOkB8Gguvcd9kBmzI6hbKJJNvqO3IorhXQ2gLl2UBZDdrk
qFIc5BTOcO3h6JziF8ACdEpDfW+EJqTS3dycmc0FZZSJm9PLDvnTpSgH08M/wKPz
5WstnGwzcKhUeLFrcwN5Pn7+oCx/MbLQAmn0K/jtQH2OV6D27n35dBkHll1ROmK0
7oAyvusbtwLDT87IBkVUTqJMEu7OFLoYyF9LwoW2z/UPqK7R6BIHxia2w3jgT+v5
KgHNoiGvtaUpCoh6taMJwhkLXf6r8N/COrXBQr3Dv09lehsV3+JnqjdWYbqGfqxf
d1ALbEk6XUsrVlIRClMuQNrLUi3BzvyIlyDooom3E1f5r7phA2G5lWIknc8gnD5i
iGftV7pdMHrlQOikGvqCKEFMu3UZYIeoAXMKASk58IDKIsRBaIX7rDi2uaUZ1z/y
QaP/J7mQ5ARiDrp5HfRoK6bvYw9X6D2QxUOs3BFWFUjLGK2leqpFD4A/Lb4lYtTK
0rgSEt95IFB+wC7bvIQnowgsrDyV6wjhfuyFwC/KCvhg3Kn21Trfpi4xqSZH83Gb
HEhFuLdUYTkfHr8ymlXVQTfZ7H2DVTjN7kaVuxtqSUEccAvaK4IN22esZfSf3KRw
lrXZkXBCE8ePcIzwMT/MfwkfOQ5xV2qxQ9kk93KG9KJ1Y891U3atMbrvZnvo6o0K
BnoJRL9kfl8qfmHUc2dz5K+YqoydFL5c9yDxNdcKlkKGNtMzr/xtOzGko4sAM6z9
iyWBK4AGVN4Puud3XyiwWpcQWEDddQ6qAoT/jMz1Bd7p4OjBXtwoV7ZfNb0S5LpM
WCGFdpm3sBT6LxMFUdhHop1Wew5ldxaTzSUx2q5zA3szGrdLcobMOaoNZsipd4F7
IHD0qYWKsUBttsvL7DckB10TWxVr00B3hDFo0vv+JOk+MJ/xqLIrWIHt5O8b8y3V
crM0HxBAEuW06o3a0G/+st43nptuSkoU5ssEYefiLJs0MafcXwYBcmNbKo5mtPTI
cPo0CLZkYRhiYJ/F2GqC0nT1NPnl4BR04UEqB6yA936v4etAvdEWChmFC2aFrpbS
qf6JiSBCDZOz9D8TbIYUoEkqy6ZkJcrrNxUhJA+bRFp/oQm8N4pHMAjP+BTYCZJE
s++LUxbkX0vTE8PpYgSX9z4xoPRrDF7jhhgPXFVMXtSRGcrLHG73xu+D9vohV9Bj
JEJRRxGRRsHQyrQQ7xWdjY2cxTUmUcd9mErCbMIKNjnTrZH0NiIKWXXi1BxSyVOz
RTVmrUzwYgoKw/mE6ItbjkMgjWg4WWz8XBlshLHBO8c5KXlzdwroo+I6Kxj44YFR
zMS2qcyq4s6tguiEK2WvT7ak49kuCwkPP5flJJ5QAGvT+g4O42w9mvG2Jf3opT+j
WT0yFaFwWL/Ma/Kgp3HwKpgPOVW5R0XqH91f5GG2jXrY2sDQDgKI6HgfCLHgcEsm
HB6kb1SD0DIB5Ov0TudBpfchIZwOyS3V4c7U2WgiDQFHeiRBSQRfzBaWyHN1OLxg
Qe2Sqa8CYTc3tJ+VJWadvM/TyK0fMsh8IE57eol9mFx+OFiG5AxRLESzVKHN/PWn
RCCt4vTLeWQGBzVwVeFpwCKKv8ahvU65dKUbOY5IyGpYQT/UQ3EuuKfSfns/jqZK
iSN5h50a0zZKqOAh+QoArn2QvgtRlYvcNYTesO2DNzH2NW86m1GWZt0zlXH3w+2O
AkVVoTJb0Lcd4Zjx7TQYTR9UbOLyHuQ1SkmWM+vJiNbc3+b4aPbkfFbVcF1hc2Pl
l+ue1ECarBnpriUz0txpGo/LIAUg0Kjq3AJxcJ1nehp++VB3LyYOWNOn/EK8KZ6t
Ko965dq2btBd0Au7FPDWwTDsPWGAVVtXX8a15CAxWwZKb5OV9bCdFxmyYlBqP5YO
jveXaB0HQ8AYvI/DWvHBNyd/1nhq8YImMKEgcjWqh0IMXBKcruxfnA7jsZpVW0UQ
BQnUFSWjmZayFT3NxZME4MON+zbmSgA9kQaSr7/fV5HNvt12Af0inLCTK8vu7jiC
2icpcaxxMrI/rOXd4XkPbEPRqk4jLidbHkwQXPsAHNJjXeXmeXi+wEiu+t7FXhcp
w20tz8srU2Sv3VFcem6I9huRa57lhX2SVPxzORK01F0UoWGHv261SKLc4jqa/L2v
3UQk58aSIIYi3w3sP4BMYq2NYEoycWBkhpXa4uQ8BW8jb1EEv6CdhCIeJ5xVcGko
9qKzstOGN0yZKYfaR9JvY+VHLLTdsX9kpZpCAbTvTYbbYnSk4JAtZVPG58Tv9sUq
wiV3pEJsrCXtgZtswTqDIWPu88iiRoCvYVoKN4+EHsIRs4+xNTL+KNbhz07rZsUR
JQ9FIqDYDtt6OYvpt47nzTLf4xVE33oxD8+NRMZd8DjrOEO912OqGraqfbgwM3HK
lszl/nVNWLDIe30y5QICySBa5IOlGcfzte5ue/Cn2uPbEqwVoNzSTDpcBKco5SEb
YQMUHutdsXjegr8TTr+5mZ0PhxtwPQ/D7AA1KgamWv2PrOTDri8P4zkNaDai851B
ULeGZ2zXWxkMQjazeS8KOz8XC1uRMEuqaqDKRZBx2vqfwzCG6NtabhFjINgUG+6s
QnuX3sOjmE/kuqf5gxWj86lcE/5tM6Jys1q/HqmIzysMKGJ3hIYKieBV3W+vUqik
jEG8zcygHXFIgMuWmJbalKIeaSJer2wmjBXToo6VN4Bi04ZuUM3cEjr0YbLylQcK
XHqpE+sFgtSBXKy+91xjI2g3Tpj4pVAokRWYHjepECPKnUp5PVHBeobkB/sdABsw
Mhj23J2AKQn4IfJR4FWhkZm9m7X/sWbD2kfGhFytiIjWa7b3GpIFKPTf6+tgRt9I
7tM1v06rUKJjWmwy2nBTw8Wd8JvVXvp8aKzbZDSN1rVVHoghKWgTA3jU6B8xquR7
k7e0kA0Jji4QCVkrYk8KfZUMwb1U/wK9Kt4TW1ie45MVvEWC8dgRA9jdy0pmjoyZ
mzY3p8zvpmC68U5wFe1CP4Oyq06UOFP7/TexDgF/hFkXmt/+5lHwYwfAR2UGkJAv
Uthkbh0bI82oNCXjUXW8WxREJtJzc3rb0ih/FdOkeURMNQs427FIDfDkXkhhnZlF
uLtGu37uTBavu1WhrJqfc2lr9zz+d/cyJmuXMCoTfPrkwJrsuLfdYVLeE8S16AFK
dujVHcE50qYSTdz/sR6bG7F6Y3SbupQhspRTe3TjHuq/fuV4Co/5ypNgn30DG/ZW
BU2nHU6gLsAF86PKIjyUgZSgGW4Bf9HucgcgKiqsyiwLJKpE88APov0KUiDfWALU
lgkwwgYnA+7oouyr5ylvbSLfkZu9bW/xuB7Twm8jBMdKDParT/5imTWZPgS8TL3m
5nZuoeQbz9t6osae15TN7JquJZPTVdMudwIbypuKc5BizQlNfCMqAXVv3cFVGA3G
rqnEc70cYd3IyWVT+Rajt7Gq2p0cHR5i3zv2PukRB9Sh1C2MUHpnVscmf6wT4VMR
19q8DD6Qm/0HsrbhlIEjOOH6FJpypXAXkjmh+7K5lviz8RmSHN31GzD+8PrphRBZ
zHV5pZVk730hAD7WTyMFmrnnGfGmJvwrx73FFUdznP1eVM7rmaowBdDIWGJGZhaC
2/Ad79xDyieZuYitaEMV5wVovdhl/RtJlF8tSYrp9w2Fl1Ij4HtMNjZ4UBiwf9nC
CwkdJFJAffz+VUAFoXa+oDpuVd1DFA/eDwg6HoRX1UpAWEal5tcpWZQ2y9uEVn4T
kGK0Vvt/WFAgNtSI4TyPur539Zvo0jzQ5+tCPwfJLaMLJmhr7QdzsvGH6Sx/22fw
4lMmT3emhdfY4HJyXI1x4UN/ca/MusQS+hqmMoHZlhrCdU7a4xqjGaH1viHUra7i
bklqPCmkny3Clk2gEVjuWx+bqmlJuhqRPmjEEmsKj5vboZSFn0ia12vJnhtv4qpg
50q0BJAJ1pd3Sk6kDtgxeXlAkGExjglZxVYdz3hA0xWL+34ZXWLtqIk1soJA1BwT
BqC3hNSJnWr45shCyJbHXN0/8rzGIupIoPkGbIctKsPUd83iutDW+IteUhvtz3DZ
ipxv3/a/sNBn/t2FqBu2FAvmXBRJcNLSIUDI4SU20BhJ2Jd9lJG1pehL7z7XevH2
yD2gI4ad4vk/gRd5eQEOfCasTXH5mQMvNV3SxiqpfzUfJkozCnFUFP5tTVukDVEi
7LiDTMoW6dQe5vmnVN2DXQebjwTHXcXUDd/F1YCp4m/JTkwjKDPxS7+k9TBChtWL
1CW8MTfUvl1bpgbkm7h1gCFvFFN2XXQPkOkQAlk+kIJTkQkTQuXtFX+T5Z/YUC6E
QBqDnTCE3zk1rxQM4TXF1Vnx9rWX422OMA9bqpYNR/BhrFs4M1FPHzgwEamRoAQy
0A46SqBDLVBp5xviDEcHskpqwpHO53LBCL1f5+QOuYGfHAMD7pr8meB78xNDYy+y
/6MW7eBOnGmJ4doBPt6pH7Euqxr1AkqfJl15eTObnbqqZIJNUe6qsFvLtqhw5b7m
6+tg/Lqo8LzRytoO3+aWRD+p8wpAWHoIZDGIyhbIloRnPWU2AGvtJNEnzXbPu1Op
vd1AEcB8lgKGHPOr0QigYF8zBfl7DqLA73+SAe2cQqLVSPtAH+cm/99YyW7YV2C4
iuk/3frO9YYqPQilviApGv7eea/OdT9EDdEMrGU+BF3YzemAe4aHQiCg3boZ/5Tg
cKd5ZQpyDCP6YIQQ1WXIFe1S8q9uqAxHNwzDIkqIsA0xgK51YzWT4paLdI2nxtoL
Fw6mxQszcpmFUP+NpYTUGKCHpAG4mfEVI9kZQUcVBjBPSl82m80tNAWV5/izrGSs
gFQm6H49rCDya9QYyWnnRAsh/0Y6FFlNy0GDZEl8Edj2NmYKMZaq2Ll60efvhlzV
rwGGqGsb8gLHwosmhHBXBp+bK9uTpFRFaiHiUrpTZ8apl1XMJm+HI+WBdAlpv4Ze
qiDW7XB1ZpSXTKvKSegpBADJk3E0DfPFt74mIloxofUiaD4UnUvFhp7g1kG7kJ/Y
10gl1Cp+/1UZPlaFG0e0Uiq3e5ra/wF0wontOi+rGcDgWJTQGlnjQsWw/kcGX7Qe
Dp8MRjylh09TleckZ2nR1fiHqibKyX/UQ7vn/NvQZJSVJa5DZUmOZMatXmB0kH2p
TpILHt2vw8ezuHS59KlviAUvTAsD9cZiUY9/TDTEKHW3cas5nmlFOvPfVn4Womk/
pUQBLha0ZFAizmEjqQed/aYRi2lpGvCJhlxzlryx1z7nZT17E3dE2uMNK+PrTk78
JHBL3W13lwt61gNjvCyvFuJR388/SrNQJme5SD/i1Xqk3Hl2ZBOKfG5FdjKtnums
sQNaQrYJqBXpiTz31KismeznchTLmYHpk2hO9F2UDj9jy+99pON+UQnjK63uRSkk
hcU9x3w/C8n2aMPLdpt0N0gI5WcNIa/h+ZAb6lii5AEBtzUDQ6lsU8GNzt/8ecJG
vpi1zQJA3FjGUQtcqWXMi30XYnwKXM9r3SXU6XvEURcX0pdsLjmVE62Y77pQBeY3
CwIl8OS359EEwsNjj05ankeZsgfMuvRuFFFT7W6ltg/arCEOAw0sbj/6hYmocvZV
2lLK+90rLtgYWYZyo6kfDmzh3U/BS7orFqilfY60swIMpP4bO9SSUm/KMi/On86r
0TK/ybE9QC2hrPKMtIj1AErKoYZGARTSPl3oEgqVYFMtMh7ZsfVlG5PTK3xiDUHp
ECoyCezzV+RjIwHf6T4wR+LQkFiGULpNqtCpwPd7MKsKE5oeTMWeYQu0fWtfpvp7
Vy/IzN193fWMgCUiFnAAOsL1AH24t5IbJov1MhU630mVSNJfy5sXyQD3BBmwKx1R
qcwYcsCjOeyHLdYFsDWyWP7UIcDZCUwm61Q2gZ8GvGPVLFu19j0ZTGIwa73OMu0r
iDO3nX56uL2HHTwjQseey410EPMEMBqOt5/MzYlXyM/7fn7wFPXgp+cSlC0kvku0
f1iXSkHjP9dRB4RjAib5sA83xhnOCuLa0cwO5QBP5oWdxMBUU8YP6f4stkBMqW9V
kNOxOlMAxZhA5S0sj4dlpscrOydObqB12kn3abF3bXO4k8vZ21IKPy6CMRrrOcwg
SNqbq2XOEkJPzn7EcMnDu60K8t3bLq0V/k6c1nnbUOWj3LTcghS4W0RbMbEL3PWJ
zaL+oQwyrO2/XL/st13JNflNst2B0inNa3qs/dKk5zQM8j1sOEzQ0tI48d776l78
zonUSkjktpabkt857IrmWGvSqxMF0Xg5kTdmTpnnxPBjpae5BLKH581w1rmEXh65
P2n6vuf2Yru+G2TAmZ2iVxpSFXIMlGArOEA9w9PRYPN0P4LayTHivZI65GyCN6+w
5qJmknJxcbSM1IPtuJ2/thbIvinLbp85WDYDFWJW2LBgrp3dC/nIHKvL1pOzpETa
n9jSxf69inhmzzrEHrQmcdxU/EihNkYUi3ZFktc60Qken1mq5CZiZczqS4aaHgIw
6r5aHqTBQSsgdF7Y3rR5rfz8MSTUYzwWVCYMvsghb66niCgAQklOzKKwRTqOR7X4
jE8n62DvHDcI6Z0380C+WrgzCtmJf20jQFUU+m3vb8no/Eh9i3WE1ALZzoIgU1ZS
tnAt1jQXT6LjSSYj1A7BTselgVKBLPUbscQwj17JYS1CWR8jaYIMTR5eVWTeeKca
Uuk5tqviz27kkXFy6zxRfinxNf2CTP5/sArOBj/SBU/NFXlWrLNVp7sgtpO0dOQ5
fJynf5Gowxn7XhtwEOPNe622axO+yEvgKilYtqYgtIcfoOxNf2Nzc4qLmsiy7BUW
O6GKlPcLPzFYvpkip5LjOmEBBG0SGzpIhtnMh4IxssK/ajzJrpGupjXP9MQ0QOMI
XAIR/JuAVMQSNFh4N18Ew/xff91EQ6D9+S76kUAmXsuxpfbtDr50Eb6Us+9NgiLv
PUgh2z0Tdlzm2YgSnXbQ/HkXUmSxvPLahKZdU5If2E4pawepufN2Zs6ZmCpWcJ1p
KX7SXUWwBYqWkplagOCMem+zMZUQszma3YDRWttTfU/wJYZ8/1vAqCkQtFQbxFcY
hPN07pQMciZZRxDmvrWs5bKap1sjGP+B4S98/0BfLWZ8xYL56yHMNBTyr+AdCQjf
ovhdVvq+AdM8HY7oy3gyoDu9Nkdaa+Rb8ithtVfrz70YfLQbuk+RRohM6ZJbD5Er
bqUo+jLrx5hU6q+OfJRrPjgA6NdyG+13Jha2pheFz/ecAWj8wseE4fyafPxgI3Qz
IrH3R6YJoc11hvYmUbJ8/lueO87IQEfBBUrY0iVHRIDb80iW9qBa5IZQ5HMKCykT
cqYTzOaR+SLZUHR4phuI8O8wyjHmQQ6oUPTwMvWgZpyNvijbtVkBEesFJjFFbgX9
qQSLFTpSquQxOYl2F8dLAI9Gst92kNCTE3M4jrO+mYt204THVsUuoCg0W4VJGQhi
hhDCSzRfNlbbuaHrSqaAp0yNoBJIhesRWBvvM7V5h1bsrayyvZMmHt6z0Xi8hZah
h7Uuj0GxOlbUnoTyA52vsiDjEwSjdDKmVVSMCPHeEh3TCC4rXmxukayn/Md1bxwl
KChsBzM+6ZJcdqoDWGRGrE+DjnTBCxPweoT4jjoOJlCaKDCvlQ3wy4QPnwImiPf5
U/H8xWG3JEA6p1AGh0vBOpp2zcEFeWeCJcijopxzP4omSedZaNS+dLTymYKp7PG9
vSTWZNRA85eIuatnsYIgG/kTYQgN1D5Yk7BqwcxjJzl+3Qg7a2BJyHJxAnmoWVdx
GJs0sIsB1gTp+H99NydIqjL840xAS1O0GIPoox68p8phakSQFl+r0uA7sjjB7v5T
NLirPkJf1LuRKSQws5BkJhXXNVT74MfrF030hyeEMAceDIW5+TwNs+aoyT8ynx1k
Gtgm4o+PGmEOZ2c97gCN06vDoelsSf7gtO6BVVg1FMguMDl+vaCmLWkdwacvLb4u
bb7er9Q9GaLRO79xxS+UL6teEH3CS0NAvHWqEljPurOwUC4zpJChZ3Bg5SyrXfbF
lg/O4kYbIvfjZpK9nJBxzUomnqem1HWv2ml1l540VzYEK4Ohzva4zmjfAn3pHr2D
COxCeRdLJu3JSurtIc0w9NRbPaQHbOYWLDOx6oLX3QCSquK9YG4o8BTjB89H1ACj
nZ/H/jF1TRpJE+oW4/v+e7Qq8Ftsvh1Eix95G7yFBKupPQTJQfD4yPUlZkw8/O3B
UkrejLerSavkbN+bO6JLRakKIAdfEMGA6sbVm9idPsG/vYYVugh4eas9JGTxSmH9
0Iz6aPEtpnBuNbnE/THlAS9tD+5TEp8VcpWrmrCLbtmO+un9kmFhEsm0EyeYvWF2
RTtFZh5i9Dyvz6+1/aO3atwx4YtSkOMSsMsCRfUbaUSBXRPjCzr8AaGW3HHi1xkT
YVeenVIoXXChzGidZ4BeBUIB4cRbwXCNfC66JxCeWO8OxB2Luw8e6VglqtfsD+IG
leTC60nbmxHpN+zRU/kOqAjldcFH8UAOr4o78Nme/O4ildaeShsRjhw/tDPGV4mH
vjl6Xqpo5P/9HcLbgW2KJem/YeRON+jmXyZcoFR7QN8lrD/bQJi2GbaMfGa+B2OV
obbgJX/+82nsgMQ/yWtXqHESLK1/pdJ/Rh/2InYY+QYhjA2X3g/YksOItpsngB8z
FqAbX7jJ/qj/A5n4mRXnhKrQfTSPEcqYggdzwyyiua6zKCoukF9S9J9YCUk5p0/r
0SknUA72G6INXxA2tAWlfCkekHASKsxUCrpkyWRDZmtZJVRucuiP/ZbW2Es83O6N
GqoVorBEMa+htUWeYGjJj9UFdEyNTbYZDwrHJBnD7wf6CcVH+qP8AbdwpKBZoEuQ
q8rpiJK0+QxW40IVoJHNY6BHLaviVvJ7FwU8mfWXwjBkN/sM+ON1f8RLVmWq2KZO
GcaFkCe+B4w6Cpnlx9AZkuocRFOwHhqJ3NIRHqjPe6qrujTH+X+fDwIaVrLSudyN
z2htDlIl1MAZDJduRpIaMy5goawbpIXtW8NVUmQc0u/qbAcRa9mYFYR/aZnQri6Z
vsDOo/rBD4EGGZt6OHdaJSETR0i1zR16WC/smsdOYvJL/4arvoyi9dMa0xXCU2n7
PJzX8p/c29fqVFdJWqV0rs1WJ+Cq/FbibQ5ykFcxwE46Sx4FrIco5YyEiEzKeKP+
+SMW2j7naN+ypJoG0vqo13Fn7k3u9Zo57wSJpF0tThjwAHcq8Sxz64akVr5aAp+e
YN1R6Oxt0GeNG4JqEh7UoLFbzACTjG/UAX6Lsw4e/l+Rj0CuK5ggwpV565opeVGk
Lzqb4pmK7YySIQhP4BRLonufdnAzNMt7imzFD72SZKze/k0ES4Y/BVRif5205iL5
tm9IbzSLS8YMoiUxFBkm9rsC4prFa10TXA1/dpVYMWhAM2eDvpZ5mnq8Yh9eyXNi
FX6reaTTUKiY1ZvnzCVA1cQm1W7B1Hl+YMPwar6XoroFdKpuCmTUQg4MJ1BqcI67
k2Oovaa+n2Z5cmqodHzjPL4H5s8nFv8Xd0ENVg3E1Fqbj0XUymOx9jR9/ciISUYX
jalSC4g/kias7Iigjmm7HMf/fo0GFruGMdzsBERpfcbaxr7HfFkq8JUmdILnVnrT
di9OE8bYGx0VogE7lWKL8aMbZU0WJdwEw4j2OOf/gSdENijXxaOTE/dzq21d/Ykl
VoR5DkU18PAa/acxymVMFGfQ5lZHzYQd0YRy5ylM2LpEdOWWaSKV4q5awWHxsC0P
uI2KK8lG/vmx70CzuQni5ArJC3+xOcf+TrX9XA4pYsNirBqC6SBFWIRAKpQRAZhi
LlOohWyadZrSFkMwwPTljnImcfVctksNJqKXVPIphTBHXCNHxXHfBwG3tieLEQDA
g1LSNRPFKTRcFHC3eB6Wp+pPGWaeR/vad90q/TGZWD8a3ZKP2Z601NOZBmhV4ZVH
sDnx/GYj3CKLXMsF7GTFX4XErf5HUlxzj78RXsXvH8G7dYF+6uHpJ0CxQT/YqcZR
3EgN4ZWXpf/Ar3UPZjjbAlK9hcK8+8HJsBkT4ghq93IMLyAIS1Bb7urVK8FEfzpx
m08QJhz8I56X+zQblyKbby+WSJYXZhX6ENoiu1mrId3PxHt2xzOrE0UCxuuWljit
CrjeWgL+69MxvTcFQBZteQgs0LIpEbBHvT0JRoAZcwEO7OYeFOLs0cvZO4e59q4D
6ZPBl0uQG0/x2GuLraL7cSOwuW4URyS6d3an5AzcxzvlmETbYg1jQLv0aocuJNf0
5zpRnx4GmglWP96k95sAbXR0THIJYIGyq9pB8OLXQQXqVBe+Bx6SbrBEsaKpJCoq
ozO6SReKdd+k74WsJPKSOHLnHZRwdhty8hNNnH826dRA8HnY+ogCNSBy6MuPx3WP
gJZ4BsjnTK0l7TCwlrlqR1UDW6wB5yP/Jn4dsUVNPLxtY7pT7GWGm/xYNV9X8xal
cvS99Z7Khdp55lg/WkGT/GD5PpuuVlrcUW/zzdtjDzEuU+FC6q1WB5cjisRUlLV0
uGCxwWnqDm0cYlbhbblW2ZBq9fEjrrtQKxnJggGH/fKuDZkrYzWhCiU0TNfr6b2w
GFD130RLrykYKdL34W3LpLc8iO4mjRK+SKf4mgjXtSgIlPt8xv49vJ+jSPZCcXyz
yG3hfbTUt7NJUv+3KWtBoaDJBgHsLLb7NLRxeKC7K+Cw57mXO/XESS2P9HwJ6ofz
hAmFfSD16o7Ox0KUpScMmy35iZiO+rvi7ZLDSBd57wxt/za5RrQvYEp2azhh8UvJ
XjnCDZZaoXrv7dVpbtLeUMPBJUHYMOVEdAT1PY795EsaRY1f8ay5eQgdwMwqavsi
yGf7vv4igT70W6IRdM2SpW1+se7pLb6qPeKPJHw7Gdp6Q0Csq+8NIkNN0GnMDxZD
ow03FK3NnrrtXsRvNg8gJb/x3CIxirm958jyoxEW6AMJeGLY5ShgBoIbbEDBq41V
oQ+Pq45A0UtRbxA+zW9gSmvVUasup4Y6sdgciq9t2RxKkLVu+bC3EnXjjEFwHp+r
/1KjDHLKpdQZxfO/f2vrv0AHsMVJZHG+HuIiy7hKfa3+1O+Tce7ZQ3NdrP/yNGne
on41ef/ToCV6vqHFVrBkyOS33rCndQ3rbLnFm/fWSg5DWt2eccXPGEDNigKREN5L
Qb5Uq8804KaoJmsMsJWsNJkwg1YOhknbMYV6Wh4Gleflzp8lhWaDXYZO4wYFpnCY
cfipUZh4kNffvgy8A0syczJ4b1vT8iTG+A906K6ohfmP/cLJa0DCRGgoeNKvQDIj
62nxvoE2Sw6okaZBT+Mjb2OWGsf8RPZykBRYimTTc25QcQvS+B6pe3dtq4YZJqAu
oiSrjjCakJCSCRWVNvnarSdOsRpKBgn29lKa98rhjuBbcpusShHsQoWBvvFDnzMK
cacGsNOZwU+cxz/wgqbzni//uZx3owRQdEjQI3L/iflhZF1Juh/MqNh7XXpMXZdU
ylImGrsQOUcAHMA9X/rK5vHRTS5UpCtf/0nqGSk8WgGHNTckl4KDSdxiGBZiacLK
/E70oJDMCjPN8hzAeYOBG5j5TZQ4f5fPmTgKF5JcyZ4JJ2GHj/r51p01Vo1pSnXi
5HHehTeWGQy5UhLLxQI3+z6MWvyEI9SJ1xm76NIwTCevPPHFrU8HNliHNBiq4ohk
lIO6sZqJ/J4yKf95V30U1+ZIljApml51Qv20C+3ud2dLsy4HtkqUl7yNSQVv1I7d
ICn0Xhto1VVTlJMZn/TcLgP1qV9f84WX2KHF/Ky8mckTYWbHIjJQHAsF+dajYY7k
nn5LN11lFbqXIyLRNyRiIRyQEP86FsmPZYGfCMGfi8YuMoP/OWKsnmMWvvhMxoV6
00QriMGEZKk4xQbHPnX2xZJnz6stKx5Z6Snf+M8a9qJG2Oaw2NaDj3DM3PIC9Azs
x2cV76v1Yc0E9XwGmOWRW21SDqM94uaNmf7Mt74OgNSv1ubEEPk158m8kyECYZqy
6WzPO43UHEje2onOOqYC4zhxtHK952RSbMIGnMjz0WiUCNFOd4DvORJMMQK9ybUz
47+PoqXq+WKi6xlH/Gzgs2KRtcd4AGTMH26M7NQv6o/4j91+DOIQ8rZ585Ka1O1L
uuZX0hc826yLxJdGu2wjmbOtLwTbShj3wXpMRs2BwJC+lXX8vtYDf4yd4xrpaVsA
P3xu+1Ad3vqTb85GDCSjmaLUw5qlX/aX59b71B6F07E4jhzAg1XPITYg5bV5Nn0r
9JA6Po0ZVaNCthggjm9iQDjNU9Hc+9pjvh8G+0FvtJSmCmY9VLPWvtxpf9QJMNki
ytny5QZXGW4jhxeA+fBXYW3skkVEBOAoIOdDy1bsjjLm8VVTCtDtJ7AuNJ5Enr/Z
BnepYcGrHxUeirtRQkkAsSpficJ/tPhVfZy6cJ+tWhFUTK7tMeT21pV9Pw5W5mz2
1RcVZKBePgr6G6Ll723prd7rIuNcEdsExlsB4EZOhJDyCp/at0khA1IXeNENU8iX
eIMR46aSnH47H/VtP9XTHbkhfprObz76cBGq8O9hdnvOBdOPmuPZGPUMQsUGvzRA
rsEa+IGRi1b5WK79TVDBxfcmuL0U58qkFUB3NK181OUZNhOVXF8bi/FMl4LQG3EX
uiBBk8nsT087crMPPxM6snCHmwXdcQu5ObjYf9uLPHdUITBev3g2746Jppjh7JAv
dP87xcYa5EJcWqQCWdxwVhrjKj8oxilSuhBzeMxpvOFEGSTLulLXlwA6saGyHSUN
lduYh8aH8gBuaqC7pjwz9H3ZI9WY9yb7XV8CzCU/NWN3x8Vyf8Nzth4S3oX2Q9QA
Wa657EzZb+aV6URYdzLZuGPI8oPk7ID0L0SBf7n6aj3m3kTyq1Yqa7Xyz1eB5udg
ZiZ0X3JA7MQ6UpevORXNEVotlztZp/NT56vRt5R913CYCJ0B87OBnLhjsFFMN+VL
jpIUARdZS3Nb6L0bBSsTEuwPSUaMtij30FdWqle0BFKt0HkNv1cApwnUkT05gPkF
qUr4l+PSvRMEVPYC8mEA6CNM/nkTXmi0MdmOq6m8B4/MSc35QzdcWXhzGqQihS/c
915OjE7xCTJtVvnOhtbX3n8zOh/Lj+JiQA661YgyASLiw3ZIQp5/O8Hm+NUKSLqE
hb0zIYihK51AgmfvJHLZKOY0f72SF89QRKFXm5fPIRVtXAuXvT9cHvFyGev7mnl4
CuGC0HukVrr2LJgdcR2lC0By/uHe98flnnea8kFYDuZLv2QzzjiNJ4rChmbASqjj
fZ5sv3V4GKma8/1Nv+silXJ0dui2kL2qfTLd/5iDFWkoD2gBrF+T3aJN74jPhmrq
iKEVUvEBthPhJBEsIHbuytNYP7SLkWE6oTl3HisBNv2JWRyPP2fpZKyOZu9PJWce
5guROgEI/yiKW33AhtAv8QTr1eWiYq1QLZ8ZTUjqQamSRNEnSpBOlc3i/PwKfXS7
n8y+KAImBmIRl+5N7xQSzT5YOz6Wev03fC3vYMEbuLRyO34lpNctO8xmzDNtSRfB
mg5I6wdgLRMspSFnDThVcV8z003ptbPifw8M09Uc9LT3lL6epMYNKODb+1/nCQad
pHslZgeXHNW/dSiZryF2jtRLRVKVXcj6+esTKmIodZzXIZy9MHG3VlN3iww5HUXU
wTju3Sb+cH7G97RFhc6E3Ysx2OR5qoP940hnFq1gVxPW/Yo7ba2J6oNv75ZDqpWU
iDrKUo6eUY5YVQ7y3AWjcDhytqtuUoQtcRbonFqTS0azdgUE/uI+v7vO0alk39QV
gAqDLwpUaK4hfkzUcvPIvDjhxNgVu4LFPTwPj60d0FuGBpwPjvKzc64MejSBwOk3
8bCDHAMCCh4RXfO3QoqVZxR+zJiqQJRd9R5ty/E3z6OrB32hGKUNTyI+9L6rkP9g
fT+Knzc897VfSITfK1RSL2+vXeXrWoxUHelq4cPQKCwIVQhi9dTtezhmHdm3fWmz
BzciCK++55JE1Rckbh0q96BMFChKambtuY3HcwVIWY07zAoMlbeH/GDimnzKga7k
D0FPZs9N/c0irt+SdVsgvsXZ/ea8iXN6DB0LLX9zGPd7K5OkExw4rMYE0rz/XiF3
pl9PGujfJBCHe5CSvDIXlWBGOry5wZcIzhPaH0dm0do2LhF9dOnPodcSrQxAMqXZ
p/5qbkFyOF8zoK/W2am2dtBJ8a3rBexRNOuINvRKchD/tVPz2Vuu8t/TPD9MKVnL
iSQK+9UgpdiehY3RwFxnaKbpdTdCDYP5MYNjpkexWradeYcOqOy4ipOWpNW8sEgA
StMzU6prbVLx+/nQIRxL5EjzGVtk6vvo/ZRVZKce6QS8pW24SqxfwOz98u7mXZpr
tI99Qpvu1fLT2NbcseGA0DBVnQmnf6J5wJ717LyZjQPRNkQ6ZMcaF7/eIbX6Jx6a
g7N9rk0BtFWS/565do1eMfX0GCllQvnDcxv53mlzTPpVbdroTKGSNKceErOcANoK
h+1iBnmSr+uSwSA4LusefNeFqSXc98kVVBVbkSfUq612j6OJ+7Ht9ogUXBACnmb0
W8zmSImfn3EHoAHY6+Z8vm8l+qEBpYMRcYigy4HDNBsW2MqmjPgS6hzHK6I+9CnE
d0kj45c6x2uXQrLIjXKJV3V+LWMG3yK7rI+L/A+adZppoKC62MNye0HzVQ6m8sbT
dAno79dfHJ/lyDm4sebj5nGaRU7Iw45R4WCwUxNlfuY2uQLTey4bguYM48N4YdiQ
kOXAhqiQ/5+g7eM19rYHIebimUZ6LXwsZWwZSWrvvFA6sNKl5lcVYNkymnCAZgtG
ZxeDd0BtEJZXIGmu8DHt1p59nn7TA1yHNKudJ928y9YG8qjGexztSN7ynD22WA7Q
+V12QjCCeD0srZY6Opc2Za35TbL0bj5zU0+92kbqcqqhh5aqVo7e7CndiyrSmzxk
1u021fST3T8LvoLPr33jDGnztTfFYzE02n2cdjoUpd2vHNYkAzJlpdxRTwrTK7fd
BfFcH2MMDg0hn1k5LA0Ci8huhZgiEXBv9bzY7pAsQT/QcyBB7bhFkDUT0tRERqmb
XC/heXkYbLfhUX0zkRYh/gnWNCO74LnWNTk3ADhJ3dMhSeYBLiNqypVlsn7gEgt/
6UJEngnQro+vlqXmw8zKBWG1z2PGrx0ELHCq05xxKqGVu4+ctWji7pGwhs4AWhXg
wqLyKvb6/VoTqhpXBQmPcd8sSmtN1+MyzxrZO8VhcnzkcjXMu0UgyPnjBqA+tGRE
jSL8ppezgw4rDS+GL0X9HEzZtqL9+ZtqN+ijGCi+paHpT8biRKspr2tqFp2adSRn
CKFnDT9Bk/stqOMSnW3bzqXeMNEtVuho41g2s/r2jfyqqsaTWg2lrJ3JX/hErNmB
icHCTuryfgjUT0mU3JTcRiM6tBjjgg83hSf9N3b1QKQVRO60SZdOYHW+bcjNEi/Q
v/vietQUPInS1l6PKnGjjwlNiFgTlD1cmXo6XEJGWNxoNrFBoS9AaZsYYMx/+2zS
qDiqdYoWug4N1jUfX1TEjb4ea024NkpO6YzDwH2tND1Ah6cXMaY9gy8t+BTTX7KO
kMfqPqlPumwkBkKd7XTFY5GGlvyAz/aUzdzslh0IG3nt8/ZSbHmXlIAd7EuAEfkE
f4ThtqVFV89gLTiKW/7wPUh+RUqu5f50ondt2eGZwFWwMr/qTqf1TO41iwbG1vpO
vEyWsTzDAF3Bs2Vssxke7XNOsjiyKLIe5Il0O5FtcL8uqHq6N0dB+AXHAkGC1VJU
4knmWGP2iTwvsHi8cFS56VWOke8LTegEFGRW+68PXLncddFPAqPF7ukpTEgMEkNU
1bczdKkIwcYQJvUBdfvLENAycd3OblNeKEi3ad/I9ZKlKIj3h8jaII9HvHY/vAzB
DqsjnbFOqLBo2Epo3fAhrS8FybVCws+hPRS2RAsIzyWbGa5hP15ZiE92pH2YWFQ+
DdNZuUUIEaJE0Nj+903f3gl+d9/2Oh9S9PJb/htZ4fpebVlY430TuN8SToS2ZPO3
oypBTHP/TlI6UJkWroly2nl+Yg+uSukqmnFHL174l97p4c+O0kJhGgCGxeVs1bLV
9aV3O5teZ9RmcmYhTyu48+GyqOg51w7lTp30/d2Cv/Dcqix0hv+hkRlxAuF6vPMo
o9Jsqthen4NJLIQKkd4Jt41Hq6Jgve/wd768ezeAnNg6v0Gd0FTpflgIlwv03LLF
jOsIbm0L+U+A7xu7F616JIF+RpwVUXeO9mBTT3diThNcPfAhum6wSl3pXDT8GA4S
3QfAIk9tr+leduG+1oaH2TDoxNJYKcQYNrGNZBzyVklMJZV7uo3LFtGLVj8kzw6s
zDrDumWBWE+UPbSrIX/ACZBbZ+z34lCR9BEKNHdajdPlQcuBCru2TMShKnZD8XtV
hF7phQQm2VNOh0rOvmqKMY9RWEvvyq/dfhvzILQSgdsrW8xpiZrfxIlk2TlyAvw/
XOp9xRX4UTq9dZjgmt8d2iTIrv0ZE/1GOTPuBitYAcTsQ0cazwHsEgOJpd7/kGc/
xLUAEGnw6JhefO1AkVAxRclrSzQHJ2iGK70ViFUDZuFlmODf6+khlK0xOyIMIj8j
KsnfclYN0msNg9QSfOH99TNbX6NeR5HfqYuj/SbMYh5jY8eEpHFz7NzAW9aAfNJv
SiUjlrbpABFTjKVvWxPtPW1XeEuUg6PFQYMzQMxMVTEm7QUnZQ59Mr4DWbH3V3Hb
9caV4C0UYiNh7+eYNeDufb4VHCpUkRp3+aCDTokxgzZLyNQWg3ZLc2r9z7p7MmPg
69uMClvIMz2gu6fn99ktx9lCNz0fvpFx51eagscEQcafX3nsJF/xQ4sdOC41smj7
WyFzXBHOKpUQfGNjbH8T3qugptW2MO+qj0goNMwuVnti2c09g4njNdR8HnjmgnMK
ZFdKfB7Gs4zqTg2C4q7a/MILc+5oHdV1jL195OqzNG07nyw71pPM0gxUme9oKote
dVxmIloezEUaDHZZuVZ8rd7NXH3s7Ba68p2S+ACNifIu2nfjTehLnqtFgUfQwncR
jddosX8EHszLDl0sMzzD8K241aw5mJYGCeZaVYmZVvM+pDUBt2FCyhNZl9QWyI/0
6IrNhY8NODbGpU238bzoFZb/C0u1tAZW92qf6lCmTsFdaICQ8Ho+x2rGl+RXNM0l
L7zb7HPxbJKAEKsQdTmj50LEb9x1jqYMK8veIqbYHSLQ4Z+WNtKl1kJskFem12Yl
ItMNcta6ArNcNg3ogR18wzi8MhquwBx9/IwSuapPBF7eBqeTm5eKPO185M61UJy0
PT1ipQ4cJcKuGVwimqZ5LWuR8RVaYRtlY4d694hV8Oy9SSG0AulRR0UPgBMh5AnQ
o0tzFSs1Dw365C9Qp/yQnFs5zLHdQah5EXVdZIDytyIOrCqMlQnpo2Q8B/0wCChw
HWUqY+qeHsVuSJ7NHMF66aiwBJBHMYz5jEZdH1XuZiWcw4zHw5V8d5+oBMp1LO6I
dt9COffgVLsmZq0gLTtcaUFW4oq9WXFWybc8t7yaZRXm2UCubuzwqb4AzhAPYV+p
vs6WA8k/eSYXTWkxQ3+251OuE1H2roBT3j6+bwNj0yv+41F6uW4KXAZhpZedmYv2
ZYuKxYws6SU0CsXW8Y8kfqR5D/p4qC+jjLgngF6DONnAJj8BMMwsbIs4jr/vZBRt
kwHKtYd1aZ1BzvEUSTOi4RFLaBAx+97Z9m2uGcgsWXY/bLrydbv4hZZ5fZBBy0it
g+DmVm/O4sOJqR7ri77mw6XSbss4BcaerKWoJd/qb/GzugTEYZJQeqguOtbxz/oe
Or1KqdN/kcjsspUU9mBW8+gr0T0+mjBWZwFYBrrOGufN779ZdekNz+94I+Y6Vbwm
bqqSZSpGSNX0Y9Bq4AnijQakbP/TnBG4XOfBsQ5ckHBqMH7tyVAhN3t+hG/wAld5
FObUYB14yVFGoJCS+gHglAfp5n2LX2olhxjkka8PTT5Lj/CctEefnQ2ondXQUIg4
7BuCAHUEbzT6eh/6au5YA9yo6dbhU4XhA6zyHjMK0PtvWU88VRcaq4Og9o0JCrxZ
MjhJwy7gGlwhKemP7sCbNlz0Sbp/ghClryPHT6qI95wiV36LhNZkchd3adJ1r0jQ
Qr24Tqhu973/OgHtUWvDt/Zum06YtxbLQzEPdNI9wvpe+36bpLjFQaJvK2i9o6bj
qSTImOR4dhQ/uVvIy15SQNt+TIqYLMCeV8wUBtchaUKzM3QgLv9LdeWQt3kUQ7oG
6s9tBISl3AbmGT1j9cVF+/w/Qe+PEo/+38pIszj26U0wWtSXyDhQLTW8roa0cX+S
9MFbwR9GYsPaSr6zzulrxypCUz6zxzR9VxrQXyffPs7ZCubidVeS0LzMWFjY9bfC
bZ+McQwfvykDP16LZ4gVG1IM3svBMyh5ladv89svgwsH9W7W/ZMaNK0OlaROcUws
BzGUjHmhmDkhViAtqOheDOpFoCrflshw9Ju0tKed08gUUzqEalZ/dZ3zcUz5Mttm
uNeuUf/dInaSGpwG2YcALDiqjCVebHeRN0BAEo+Z+NwfL7I4YfekZMKu6u6MHs4q
RIUd7LsPUDU0tmT5id2hxY6FHsPMolsPz4XgSqFacJHb8LyIWmoiVWJ/c6hdt4yf
jP3uNr9nZqTi4f9z8DJ80mJ+kTZ+BS4itl5D+6tUmtaf/wnOm4GtATYKUWpqKEfy
AsAIAdBEEdrmJc5Fq0ejPY1NMhqaJHgG6iMcVcjNkuyaEYQmOhNpKoOpVpUwOvz5
fqYC+XFcDUli+HAb0zS771qcRIySJkY0PoQxlNB2E8phehDRKqdvBSMsWDj5mMPX
wPMoPlbTAhnHK2eucCh4TLXKLJe+uziCV8AXR9MTzv8/QzpXUkZETzYy5M1V+Vq7
jpcvhWtmsMbIqxOQp5wom/uAWLFZ0c9a7g/fWn4P6NhzD+wDJXMBPA6vrf7goEbC
AKOgCQSCun7gBH5suDDyiE5DcLDxXu6OdrZITkXi+NQETHfEPrDYYXYH7QcpKxSr
fpBiKX+2Wkf19GCWb9gPmJ6OZiLVn7CKQmYpsdhH3xuv5KFBXEAq4tyMcIUvgJsk
CWQAZDzAEhs0r1IOKr1f9Cl+jwpmF1/nJy/tN4i8N6pGyFIltcAlS8lZeiGOPand
O7USNJfw9me0iVmG3I4bNW2WfMEVKALvxHk6eXv3VltHqbZjDbD7BjteBUo4tmfI
kopJRH/K6iQ39ANnRQSEv4pov7F/qIuyaIlSr/Q2v/5tVP9dRQ/H6BEvy+Mj5VCq
C/WzcspbE9z0+us20/qs0S2CxsGVc5LajwAlW0FayrgtB21C38P/1VFYjh95aJpd
rW86JgDajoUrCPyGeiiJBiCsmfP+bpiORlq7TfaekTQc0cW4GFJ4ywKQULJ88e1c
M8X3DiZ/yQb1G9xc4uNVFzCkHggKDsLaSo4PkWpynSi5w+r6ATQKlI266aAFavFz
onbOagBUKatRF6y+yTD+HjzWHrHnVVDrnMBovoOf4nEK/FHbEDSGXikEAEXt8Ny2
K/QKYiunT2gek6Upx09VX/c7ObH3fB4X8bJDBHrXYlA/6Ku7YMb4XL+OawhjcYlH
RqAGcQCryn4LDFyXEUxzjzjSgPTHhY+dcONWImQUdwZFS0RF6bhmXwnJ7LrOWULN
X5902ycsVy41nwdqjcL3/9UZt2uVzJPYq7c6q6nwSvXG90MjerrotgS51oWKz3Vb
vJ5Ar75tpIhqKEVfJ7niBfC9ZIU0779IhQuhtuFYf76k2L98FJzzWhg3/NKNTjf9
q1x70SPDhNvKkLD6/sj3V1xSSP/Nfv8JSZFi+8zScKoi6BK8EaGjB1cgc9MwGsKy
wDVSyUc1FgxvcVp4/BAk6wj3dKRNoSK0Hx/uIf9oyd68Sjh8+6OZSHwvCVumcrLe
Ym9YlULdaOTOhZ1q13fgQZ9J8Bmtbt/f8sMIzB7eNXSdabQZXkDXJXSwdiTNTT+M
EhYHNsebvvaRODZUOmyy0P3JY5v8U3MZNloPK9IISM/zBiV/WGnvBOL91FrQUbSN
7XnCxUGq361c14ztFiiCSYcaXHyBNn87KajEArDgW74i5/sTQH1THaDqzDTntP6L
vSh/N2RZ8hYRLpsV9piULk8iQ3h0PrN9dxvIiriR/d4WfHPgK5VgzTMEjXDg3fe/
rlBLE0xtiOcqyT8OoEw7fQiDwgvzj0Nl4AyDO9/datZNZek82aC6PH3TdeNkQEsA
wynZarxEdGw+JtH0F4EDLBAccFhXZXdn+G1N2iPkidjzBG5kB2vHM4Ebx++v62q4
P5YW72d+dFkghmVe0vLqt/FaZE7zNmzhSC8m+br39VF/R+AhgB986SDzlEkzKqLs
IVAPs2V/RYzYQomwe275Vsy20PvgIm1zwg5vJAVSaoQyw0KnNyh1MLeC6O8ovVdv
/DgerNE0CAq0BKOKtTetoQDdM2PI5E4BTWZOc8mJmRNCjSX+gQlMD56Bg2hhnuQm
FJVOVevKlDEt4LRv9tlYk0mZSyyDJ0qer/G4FpEXCp+q92b61BOeBf0sHY98ZrcL
ErmAiwUYVsKw3bPU1VLVa71y8eoMvhFH7uHwUO5Sw8ajtUVtoCU+ASRBSCCHm9q3
vnbJ+uaJXxF3fuJ1OX7dO+L+C9NtYiy8QKRjc7S0CwZd9h059yaUJS4+7dZ0fQZv
EkRf2obBgXf/d7vnvDs5nt8EIrDlg5q9Zz+b+UWMynBifJaAq9PwVeSEcQup3VP7
+e03g0Kl+IL1U22UYQ0IWlNV6hhjP1t36xYh3LexSXrlgMWQQhY2VvoWDKI5n/KO
y1OTbNFKaNuQ/0yncptlcH0IAzyPV42rAzYsdqvkvbH2O1W8WZoYO0Jv96lsvL5z
3rBVyJshfXDJfeiKRApOZ33wuVLSe9GMK5CccjWbbVhrXM5YNFH/bFsq/KEG7QL0
TQY+YnrVu668lDm6o/W25HvFgfylsQVhAWWgqf5qOIJrRMO+dRf4aAByAKrnKWLs
LkZo8eoFIMd9KM1OITBsB4LpMSSXoywk2IwyYWjVUl2hYimbG1zv34u1ihOk4Ryd
JRNJ8kz2uSPOswEOAIriMPa8h8XdZYNwrSRhEqONIRLzYV25xPhq1yDOWFTrmAA+
CSdmgLWdk5xm9QU0eWfmNqpSFrajcwMOT54p8faX8shKWxsEIWRNI+iBqKwCS3pO
zbwsFH9RRExCn5McA2N2N/o/1e/oBTRn7MAF1Uj6vuTCPN4DsUAHhvxUhUuuViSW
r8K+KrNOBH58wVsAD4bf2Fbn2FUpqvghglgZQZWhZbp3kSdZISrZr7cCzm7DyS5+
zeS0JONc4lPuBMHXy8KIDcFMrDbVOlGjGTtWSTktMlyxLi4ppneGkFEi6242kC4W
UnYUmYbnQJ6JImF8D08SBOQJsuGi7Q0TjBHZjIESgjGfKWejkpJkjrxV/soemkio
OhoMpNhbz0dy4LVF1Odn0W0OQOacutXmh4k9xUtKIu6Y0J/q4m0vzYwqOnlVZyXJ
Hwyz04cT1yvIjkJLS/vMmlMP7ou72nv94tAv4N3H6KEwk7rdg1dXtDyjQNjarfMu
j9NlEXmXGq2ilkq6c8EFoczGiMaUIsqUKfVO0U4NDJ1cpXEC7dZNc18Bjt2fMn+t
5ReuOvQ/f5KjgsFhtiRLdYSx1JqIg/W4I1I6eHSa2I9uDtJgY+JiNCunosRLmvoH
7TzSweS+rl4pQmIb9x6z09xmInJJrc+UfmHcJ5CiQupNK9Us6uGyIXuy23PBnv4z
PbfQfOeBMxvKf4UXspAroHF4AzK/3wglg0prL4eEJOGptgNV+6NZDLIyA7lsGjbs
XdP2R5YR3UOpP4kPt5q/MBIjZMlhscSSMUbwnOs74VJQsikPqtnWjI8Zj8uqFWXf
nxdyhDQLWZf32T9wyhSb7b5s4o8S/HlhVdwGuoNwJH5Brjm5BLrzkwfXBxMKR3tx
lb83UfLe4R7KiMUMqx+zMlfOs3NnHn23Z2FfwTJML/8iIzUD/9B9DGxZOI6xdGgd
8EHXNMoLZnCayeWu3yyuDZGp86BoedYB21ZtmCgec8kfT/VgmNRuzbCDAWGyHfEH
6/PVbnZhvc3X1+BvEt3+eyNasYWKyuz8y9hsxVC2bn16wj5q3CdxmMeXQHKZxruO
2VnYaLtyrDoQpxNbBc0M+71bBIw52kg73MeqIc2Hrx0rVnT4djM2WcGn/5s1DU94
H3m635ttwoMR6p5UjLjvtA+s/cgLyES0iJNfoHiiftBxwpWllUHzlze1yXp+IqON
u0X4/irp0MKO6rVOAt/gC2I6on1q8aSl6DIZylqP73BNFKZZgGSRsaJ2vQt6z2Na
jm7ot1CMIjNxnv5FgOC5fdnlRcX4UYWb7GHS2qGMO71A2RrbnmF3e0rU+1A2IAcq
gunV1D1Pki9nFfbk1cN2MLicivOaA4IFMAVYvRohFtcckwSEbCgmTVuAVhf9FqCR
Tpcu1UFxhFqMrdRrXDIwW+ZRp1LYbSyL/xC82FX4peMY2EWbJ1vpEBJ9DJYdSIrp
RW7J1tejhbRTOVyxblFX1YK1Q8TKy42qogRdbgwk2ogFYHsdWpXkAajqmR1Ux46z
aKsrYmjmWBdjLhbg5V43230O/n8OH2rKguGO7DUPSv3a8XB1pHy6D5NeEQavZ+UW
kxyl2U04JN+H6Vl9yTVB79/SKqIgVB9LhVSUrgZZX9+dWyWKJG5dQ76A4bzpgyMv
DoLJbq1JZ+/IaG2r8IDgcH4h+18KVc5xNC3lGrR+qA4zYBcvK969D3lzBhpt79vi
YgnafX1qWDtknZRjAK9XXSYjDBU8tjDO1Ht6dyu6CymSBIxtv02D0WogbFI6bQ+4
rPXMf9uNojoSBDH4qNWVz36uwok+BjyY8v/hIk+g99m2nTDQyclEIW1ibmsy7Kuy
02Qi+5Y8fSK+mwp5W+fzfkx8uLXzrCQcU26LMdcr7hdJCw8j54lmHFvmWU9ie+7S
YYVZ2DNjGtygneu1QrlWvUz3gWcslZH9ConkzJ5J1Ky2dSvrY/uWcsr8pHYoc2ci
rWlD0TJU4xUcyuBn6IwiSyirwhY/EhyfibL/3aCZJvPF/JoCULybIEXdPKqNK2YY
iAoLIe829DyP+9KOn4IsM0gv5f6+NhjaOepUt1MpPUhJqBnsNO7812z/QwDAn85Q
ozRMNjs2USxxrOfvun0HG8TQ9IE0gPltzZOb3W3fb2m5C/1ceGH1l2jC8yk+usVa
t8ZFrstYrSzPSZvpcxb63xwJHo0glxh3vnKsOcuq5sXa9dxEP2CTC3XA0/MnDyk0
lYW/fyZzVeN4nrlRSDYCWUgLUYNxLasVdIpZHLNcUSqJ3kwf0whb16tbTL/zxREV
JQbqEGm8xtv1nwN6z7bcdLrUIT6BR5DP4cbC9RMDhz5DwnvlpO+a62Yf6BIMX6Fa
Eo19iDoQfx2WC+YjcP5LZohQxM1FE9eZjZ+pdb5vpuFMRU5y9Or1UiEJpiAVj/Qb
qST5tsEwR0bpKqjAUj2mHgyemMAfNk/NKD0e4Dz/Q4a3jBMMemY5UIlijasmOErj
IVTAY87j5Xh2dBNi/6Kwkl+EbDT/yC9mO+BMOiE55BGTJ7E0ZcFWMkHsja5wMfWj
JoVOMkFzVXt3mdOI2rRwXP/gQskOAfSt3LiDPGYdyswFxsW/zE94/XnIZjI6KwTD
80aqHtFwtwY8DPBQ9uE00hixrL5ifjoX5uOJOIvaKf9esnOTtscHEBDA8Z9dlihY
aGo1wPrysjAVa9et6aWxRNJtjZYNtj3cqGfHSbqYpZPJ8HXExxjgrr1px3UlLJQ6
v35V6ffYeGKF3NWhhdpUENT70WEbou0SF4YkRmq1oTWo/Fp1S/Ehw7NUPvVkj5T9
NgjfcN+jz3xeIB7kn91FyzRhgJ9cY4IYANxwxceo1ao8+i6XS4KrG0Oz7lq6VVeK
AF3Sv6/PUJ9T/In7jXiPnfKDukPhMBo4d5GQAQQFiw597SthGinLHtyW8UtbqFIh
IOr8FroIYO21dncDEyIEvgusmoVlp1hcBh+SpEbyU06ZuSRXT4OdMlwsu2GmcOjh
jcLcN9l2bnVX+2rj4yQqGpFBfXwPUmd0c4YhttKcnCnUj8+u1tVBY/pVTpGp7Rve
5u4FcE2MK56HAPdv2sDXzfGlSXzFAiLqL6CTDwJQrzwLCANSkZNW8aAtDRvWWj8k
BlafxxGari1GH80OOQ4v4OH6UQ1D3T5k4cEJq7ECPSEbcLE6iYITyw1tNgQeLRPZ
n/9o9E/wFD6KEzOG/nnWIkcnNelDoJp2ErteovNFAnft8Dgmjn65ofAGjnXmSfjh
+AnjpyWME/DzahXq1Q6bjqnU9XlRcGRl96I4t+R8GrAbrST4QsM+eGS3dgznIHhd
GmPwmRMAZPp67VFODdyQSOJb0fjgSlpZb90aUnMaQHwTZv8jt0hY9GuRFSLnmv6x
SxISZ0VMiFK+rqASyJun7rWDGd3clDijHkg9ha599/S18O+sh6nXQB78Mi3Qwhon
K5PUOwTixX5IRHzYwAbIJTOCiAe4ra2tI9bg1LZStEzfWeaGjJzRsu/RRJOH0YS5
ibYuSkVWOY+9YX/A6pTLe8dRlRuc/4SLuWYB3ztYrNhtYo33JYQxI5z/q+lKoXGK
1SIjhp9ox6FagWN6CmOcxVZXz8i5cuzKzYVj672NNoFmHi3ysDYfI9G5+aPmZ7q/
xJy1ID7Aa3isCK82sWmUHq/+6ERZVwVGkCSSH+GRkdegsJkFl3UU6c6pBy7/qvFv
WNgOsLmj7RL5uMUb3SbvOCbqSLdJ4ksYghdBfQXfsqeMpSsWCThZwjD/eFN0V3up
dATdQIM+hGl1adywoqPWxI/cB+xnaG09OTlf4iJk83n551Bh2YI5BwlSUgnVcYyA
XW26mGCZj3AUjKpieGThcNDhQot775nGl4nRwwdb/VnaAgUQy9hw3zKhHiq/eM20
VXajjEq+wFxXsWZawwtr/cbI+nOfuekUqf7/hXobJFjON28aAagrzw8psoVfwbP0
vzz0VZDZQ70fMoOxUWJBO4PThwnBFuw00AMWCCFFs4E+TSsVqY8Ia7FcFefl1ofw
jVoeGbHv2te6EbI1HPkPth0l624Q2dNBeNVmZ2BVIO2iAnW0LPARpvdsh3vBXmtN
3t9CnpTsNwA7QKn3Ex6G9UO3u690HrsKe9DmKYHpQjb8WKu2noTTZwTrmLmdBFr/
FajunX1iqbgmOo8jBFeiT3tDmWDDgPxfuXtxzEv1ysYWS+mBz0AAECqXaJT8dFGe
yPltRFTmyqlBCAtrs/HWs0PpEQ45i5jDFMqOUtBR5KW3aOiO2pq5rQZ8ulYiI8S9
Ererd5EoClgswLOD6JcNricCTA2t13jN84Ny7so+ZkHXf34YQ5x4sIUdfONOctBu
k0zrfxrUgm/Kxi5EgJA9j0cCZUtf4Z/Db6mxFLvEmeMr+yUbLj09pojcEEusn2M0
V/S4UQ7cQK8BJpDGS1rkWMLLHog868NKGF1bZppwlKuC7N3XZ8woa6vqG2I/xcaR
JpLsFlkgvfY99kf5S8aCP96A2ytSEuVmrwBJQSUqrRD9u6Amb7M/msbp0SFyaTUE
mztleQUqxHnNFFKCvt/nyh88tSvm2one5SAEEkIN0hMCH7K8EufwIk14H1aXnTz+
n+a5mYVkaoVxvw0RfWsiREsxcobm2c4GvN2VcCJJ1J/JC1oVMP5XjSXJIwygoTir
U/IKCiulpMOc9GN+9gyue2TL9nbgW3xS3XSS1WBa2d301FXTDZM7ic5GGuGxnpFJ
QI0bJp8TEkIGbMKvkXleXzr65pcM3/A38nwB6JripdTtzbzXHZn8Pjm+f8jyHFat
M/J2addHZ1fnid5REIG3VFrozlV/Vula/zEDh+6xX/lpJ70+8AvPe+nKjoKzlAim
cIjNJXpPEK/ZCA4HYQzMG6830ibnu0f1I6f7Bc/xUQGJUBApyL5H7+4JE/bvbnil
iajIk7ANW6a0oArAFJFAUnr4fgw6zK6mK0ITmho8AiLqeh7wmGJ0yKOjMmnXXKc5
UbPZ3d3/QYEHr85oceZREFwdM1FUAteoBlsJ7rpeM4b69JCneVULUa/PVTiNAmVB
HlVmKDbsuEx7DIT0rL2VbjOXjVTOCGtHJ2eFj+eVewEedf2EzfHSW2oDIp0nMN7r
ND5PAjz7CHWaPUQcr5oa19VClEXCTwBGwxK0aejXiF59gqHVjLMaeQ6hz45p/QT4
KwGM+t5qe4ybuPYJXUAqmhnTWCkcxAiHrMMHgR++KjE98Ls4hbaF4dxXLtGED9Vg
p2AGgyhc78XnAzb8mzWJezeec/K1SCHJ7uaVvhBzFDsQU7KBYb91zbSp5SI/scwR
CHzJREB2RckKzc9jwhCF96aLLP+QBUrIL4kcfIYh23cd8ZO6KjDAYi2D4dJSiEVq
vwGcRTpGYVpGjH/mF4qEGMoDbSgdaX5fYZUNyuSPueGsYr8P207gV2QzHE1OfLd4
c7ci6q2h3xTlQxyoeudop5nBvj+5ejFCbX117Z3A8JjM079HbzQ7KUW2Jw+6yFwY
u+DauIRE3V9/pIVm6G9gNh79HYz1XcMHr7rvcvXyA+jojNBoh/ndhfi4rd8hy5Hh
szk1iarzdw1FfLHW8qls/aieVmHUxUxMPt/SLAoQ7PoCZxzXC5zGgkLZuAkzURst
mltz5yy0avJJqkf9UEIGpQES7NEi4R5z7ERxU9attcHxI13AkDesS1Ly/PzESS7E
Ap60XZTWVcH8u/8YZmlxVpmKu2+X5nHHDVKOxOsz6TkU7qJpw7P9nVVl5HX0rSwI
7b+BI4SFAEVvtwiA7V6BuS73KEgNv2RxQTvJnHUEVYiDFfhx016P2vByi3GYIBBg
eC4mtrK0bam0MP01dv81Nqocd7GV/KdQLZB8QRGDH9oksIV8p18eQqQtQRZr4Mfc
ogrFWLTdv2TjtdC1a95GDpM8LVNp+DwVDf+DEoDsHAR/fvY1ylLr8C+0hRomu8v1
BltoSW94xFsa5edlavBJlJWHFlZtXPmw0V7vWpNCCjTrY54hkWQ+zmvSPJNywDIB
EataiBZeTRdbl1W/q7X3Tc2uatWQ/S3n2pO2rkJMDc2lisS1KqqHkObXYl0U3jr7
azjrYbfFLQC5f/q3FoB61KwnAjtDd5kEQjOPg5yfNTs1EzpsuScQgBbiRyfAO2+k
Rk/6qVQgUVBM6A5IQAP387ZIm/D5ya/+iuVupBCMzLy+lZaIGXZCkqRPb6X6+MfI
vdwpyf/xDE4EPL2+UasdWqmyobbyl87o9HNnYY5uf6RFnLIWayfPEsre0FkwWkaX
VHTTyP8IVTajfTp24zzBHTgVHRJOBacFsX3IsIrB1qJ7lMgE2rXw+kMAMMiYbo+9
bxbOEcUMi+8UKJBJyyT4yshk3InSIdwp01xbf5BzZJdN/gFyuUe2dSB8jR/UxaNx
AShaofq+FQNa8bXUriAHLwXIQsVQO4M6+i6utPKq6EgXZS/jb1mMWkbKnPLzXhK0
w37hlptWNRImTaA1oBCsnblYG5tPzguw1cfDmEGYe5xW6SNLcKBvg7Awn/yaqJXU
GjEl1ldzlysQBP2OMvBSr+bVQoUxOsD6M0yhxX4TDfT315HQlyI5QiCWOkgQPqw6
aENgbvMB21GA58hPdEFp8wCijvZ5VOQECpJQ6FXyJiO+4JxpXRUrIbcxdgZIJTyf
WxXNsvGBxykLn4isITetvd1MqlWaMgjPlNcjQefbOOmMkngRVAACpWxZDNC41D6u
N8hj1ffOXJ1KNShLIp0j/L56sPIzixDrFkac1d3V3YlnY528zgCkRs3q4boM8fxd
IA/bSwbM6OLY19Aaxf1NJ+0u2hiAP1C5mI0c4pzXiHVDsm+doEn/g4zToZ1Oysrc
hhNx5/gGNcr0jfzhMZw7dT4OK1HODwmrO0w4eWw+pBebHDNkTYU9f/x1dM3ZacP0
SyjEG5E6UoQyiZXK4Bvwsk9AlgBIj+iKu2Ypl5L5tng/cvrsJls5j9M0zR1fo5v6
fR00/LER84L2FmM+vKKFBlHA6fEc6n7kTK3SWXfdERZa6Qr0H7Tz2pvT5U4UX1TP
qpwYfTekKFe56pcE/aCh3UrVyhTSEaNVhVGKa1/iyjCMdrlZLaclIhAWQ8e576ci
0otZmzIeklCb2N4ISDt6VPH+4BO82NCWP6bzX6Nfzut6vvCC9ir3HOQG9+4NuJfs
rmvGWgCA/G5xDoD6G7/d6LMljiQ9Lce3alVV4mwnIZLWBIHWW9537iI1b8nuH2tW
ngWtUCF4NXpsC+kRA0+Km5fTCZEHX6rJJy50XtbdtPd8EiCho0aRq5gC53Te/joi
LZakS9P8dD/sDg5CkU1bAMFMz5k0BshUVvjjlQKfJYNL/6DWs8S0A4veFfmquPH8
195b7Ewlwgk463pMWWSx0Mw1AH922uP9QlykCM0yNP6AQ1WWJn1A+cIDEnWynY3H
esPrX2NM2zgCL4XvbCx3wZm4jGbbNPUcgS86H4LAy8BeAUYx0dWtE7kMPfu5UzUl
o87JjmHvkcvEYOMXJKr9srkiYtBLqcKgEObLUSbY/x3fb/bcjZz3G3S1h/mUfErq
IA7Ti0OIawNrpuuHB59IcU7ryZDrzeuPZfyZh3IP23/hfwXy35KdxtfrnRNjRijF
dEZJsU6rw+QXMoDRLTNeJSJDWfNJjXOzuuuXERXbWRAXMSPUDKyq4om06U42MShL
ncGPc02X0waUWuZsfKibu3inYfQDFE7xXKAMQwPY4z75uoP5Avf8LHLBMYiYBzpT
f+HwCZpLn561Z9ld+S8JW2raGmJ+sEUTzOtNTwQNC2GQBvjAlJUEZH8Y2uZuIi/w
GCAKDx1qDqiGuuVZP/89zh6DYZockSf6x7Q2jEdf5nVIGUZdV/6IzKG+6oAWckEf
l1xrapyqjGxWg95g3rtEifeHXnus4Pp/x12kBtPMpJ3I6ArAwSipjq97sAI6ayls
CDhfgEg4fUu3jX4WsKlNDrx8Oe9C89AC7OXopB/r9khl5C/JBY15mulUlSZwgG1T
kg/8QMA+6B3EssKrvVGzeWoK1Qm+Xq1nhccVBmvSaxPu5O6fByt8pCdXN2zgK7YC
ZdgZoLxDqbBBDE661MEK1PxUtCNf2DImsW4PteFUft6Pvlv4xIHbo3739mhtlP5W
GaRr6WfXee0HuOdJzm3JClijLbIyNV+3x3cWAsXySxPyotknu8njWDidaAPvI0QS
E1ReBzyoxZCm+x/z1AtJCVrX5uwItsPpz7F3p2Yo83lS+ilXWM4aIWUEEUmJYXE6
nTnaRVmIsTzCHYPUiqygvH8HdJ02NzdyF9BOZqtuhTciDmkTaVLxx+BUZBmvSBXK
sWuUMDv9A/9PfKQ7EcZFCViwKP5hkS8LVe050/e8P/zBfjxjY0K4YqARf7x2d0Av
BJ2bOMqTLrsL1E3+QZXQAhtYSgCgfc7MZSwGvGCElEubowhcTF1jMUKyCYMkZTYt
WQYowvVfzkc27jk79Fj9/UkSuZfcOHcl8urxJ2PG/fVJMGn4/EkRfNVb/C/u7MJf
Wb5mciGhprju1HUjPe193SZU9I20ChMTIylV4WQWcU7Ubn85mw3TA5cAk8C4dCLj
RyYjYZX5wfbhgDCWDlPmreKm+LRjufcuovFph1sYXOpSzJiNcb9vTNZ6CmRdEwLr
YaLfmMTcmnjMIC+dZp9IiR2HxXkPvHZ94588SAiYqP2zaS/dvnpNiebXPfjPS8RM
u2IrJurKabK3sp0tBWAJb2S9byKLojhRuY4gaOD/X3s8wuiL8iCqNTXNyc3JU6ra
EC+KU+Sa6NTD3m+YdA/zE2uPNKYVpeM74oWEEwiHJGQzppnQyjnwtDmKjDNrlrIb
INs8woQ0TrfB8R3becnzmxngx/QhxriWsmc0lwx4mq9oCLH7PoJKR7nAPdAnHNhx
4d2xpmCNP9qCBC7vFy0s0G+i8r6G4XzInjM4U2P3hYJ2zih7G2QIcxJtRXt99rC1
WRL77OIDA7GZYDNBaybsv+jhspecA6pQmFAu4aYzb8fNUGTCjiel0HAYHwx/htDh
DKlx2eulN7rndVb+UcxlN52lCJESxgbRqbC3tJ5zyH1hBPvLYH4y/PF9EWIys23+
ogikvo0Dt+k0umOd4kmz5u4PYlviIxH1D1Epcz0qsSz9enH/GZpowvVvHbX3Vlqz
g3e0NKPekKD/9OfQFFEdSJTdCM/CQAjwD23wV8VTJTBdS6TfmIUKV7koQxgULmJG
1RVDZ99Ad6+2lDrhn2WIZVWftoTTSn4b6ju+AXVFKki6g3/TTD6fpsWxQHKlPpmk
4zPsrich/S3N0fmBcUbcS7Oa9gstLt1fOH6fAw1UV1m8L7elePDNyaWrVPPM3AAK
X2Z4DKBKLmF4WokzsNPAZqyTwPpuKHHVVKycm6krc5cHepJusgdZN2ji5vvjcQ5E
PTUsjMsVOQyPuTCWinFYcyfES0chtceERrZhG0adD/wX8R1sdSiSgLiEYfJU1rJv
zL58wTOpDnDZsMcLjwJzXZNp/68ZZiuepAWFBMQo32z71x1Cfjwb+a9gffGZhxuF
4fdcDxKKxrYUV+VZX/TLKJ8Cpn11pU65nFRb+K62LcH3vdQXs0PF62vkYDlcvqM4
960AulxorAd4UXZcXR0K2VCxWFrImlMaOALIeo18OGmT7WCZojdq9HG0QKZrOckb
NFApLrR08SnCuMsR4ZcXQTZoJOkTdGyQHNO3FeC2Wvp3kDw67b1MxNLdn/h62gsB
MKtS4vh0i5gyL3DgeqzL9AUiXAc549/NbNhIZLOgp206GmC8+O5sUM0yz87e5lDs
Qjc/L809CD26jBrrDra9YkhW3aUPQLb2nUrLT3cn0mLXwjY7rcG2KuGzC1OgPSw5
cMuK4UjKOFaxt46UUIh3nY7uFiutQ6s6k9yVP/VtlsCxsyeGQIJgomcaOG2xOvpm
cefFx4DT+T7Iedrk96QAafgpnmkKooA4aKx8l9grtgJJYaSKmqZl3gF4bw3VREfJ
zMEH+F5IVY8dw0+VhQLaq6HI8gsDWu9rdg57RwH03gSv4ynBMf46P5luDe7nuM6r
fummNV7rkybTi+Yuaok8SYP1VHB45mJBUeH+znmNfjORXomviUjWl9IM9lnGWiCK
6lX+xgvy4tEGEMy04OuUF0QxOQKrWA2cfywM3N6Pb8mptQPRwJ/vPVVvB4NKtyug
1I2AoVGB26yxdCNa2/7LRmOExvUF6CuQpWhbbrp9jxHjr2sR5VIToPVMQYqnEnup
iYZxAUOb6TfhVRbejHGn/OA9oOObBPXzUG34T2n9Ug3o71+5ToKWEAshpNIEjlVW
pNrVufrQqs5Q5ITarE0h0qEAKvFELsV+genXNdbtDQ+KYAFvUeIHh3kI5fcSMeyE
qxhlVwHArAGmjkCpZ4+igqDh04zv/T9W866RJNb0vhWfYLznJR9N99j3H/loDG61
O939zERm/c/3qKUbucN6vJM5E3nNDtDGgSEDDgYpD6K9jjYNCeuvrlDBbsD1X8/8
aUfDv8+cA9aPYcIqfRpFgSv+V27arL0kenzA2Sk97MjrgAgOWQjDcMqA4DgLE8KO
MpE5l+z70PlY9oB5Ha7Af60pnf/qktQLSUNnkHdt74vlXXdMjchLN2E+7ftw9onh
dA7SbcXvvGu2LKfSzh0ckmnph461V28mkmWyqIwxqCsemT3z5Mf4cAIjwrqEzjDu
KQQUmK0RigrHi41p/isjzgdWa1pGSYL34EumSQO0olNtbfRyOFS/MkGdRF0Ir6G6
JtZc1vBxWWzILWag5QW+2U6GPpEZCVW8jxO6KiRjrO0frccWP4Vv/MLFCqHOblVD
QDZYXXxv/PGQpZvkotacSPsceRtBmKTqjAKKcr6bVfS3HYHcQZKIuaKapuJTlFGO
BBOn/xHRoSiN6ajwCShc6F40DX8xJIBi+Js6V62/3S5rvqLWGIghAQHUMU+AJJG9
BQMj0xDN2VTnUnvGObPbW/Y3tyoZ2KpcD9HiDQDyQg9tkgj2wcid9TlPr5IvJjax
nz7EtpSTST5kMzpKa2VuzK5PfrdcIBhY/FBrrmM4dlGh/02S9tHMuqRmT3x465zB
BWBJtPMablx1mOD624ZEbG0c2hJVMxhixyM01sb/Ev4GG7FvLZMbOJpGaKO5yGlG
chk7LdWPJbj91djnWCmVAR+LBufrWS4RuuimSV297owuHnNH0x0vWiSufyzM3ouz
E/2FscNaxSgWstZYWGZ1dEIVbvp1HXDKP44nXP3qWDizsyQKDgW2ODZkO6Fv8hf3
+Gml6ClO6YFDzBzWeDCrBVohvq/S7xc4qnVLig9Se+5/8PIQCKYNnbxOa+CbQ3AD
GvKrYgzJyBoF/6P624CCX+jvabQG1/inKiN5A0ftFPWPOgwJxBwYZ9rjSgJG2Wh1
a/1ewqmGCdNETgZiNI9XTQLNmwVl6g2igQsEl6ofYsoF/81stiuXlYbnpuHMzSGc
ZO+cqXvJp23U/JsQh6q5RJwQWAimO58gR3KI81n86v2meSd5IAI0ysNMySG7JJkw
/IBbiBHtkuDHy2Nvd9FkT0+/p6dkf9mH5mC0IP+H2gnwwTYBhliZ93ZyIr5KFN1D
bAKGTeCJ8bvUm+1YEELS61Zj/MhwsvfU12ROMZLvqgD4FmyqLREDPbFIk0DIrLLz
/vRLSQkt5Y2fAuoz+s68CldY2og84TmT8NeS6/iKKXIjuRNvY00Vw4esVVaHrbi8
08n1MANZmno6iz0+7f00MxqGMHhImB7czhfPWkdyUmrUOkAHmjB+JXGQnTFcFeht
5E3XRPSXZFKZZZuXpryBHQSJaCYBUqz4nFA2jXUhThfls8Zjr79X3doojVvng2lf
7wOCzXG8ECsoT4kXW0Rwy7DtRGVbedT22ACeGwE1EzDD6inJ/4yB2holRuT6PzDG
wFUR/W9f7VHwWqaqBo3j73xCHHSzKA2HF/ZzBSqie9slRNM6opWfhMsZ2OMPlhhf
kmEmy0lmCxLtLA+VpuGPQQI0UtWQ3jVMZL10vWBijip76OPa6stj5maX9Kqv9nEx
eL+fEfrNLaXeKrhg91sw2M2OiF35i8UlOsBq9nm6F7aTWRXv4vof0x8Od4+az3Qy
H0q+8WsDvqhJ9Nt4z4HsWtJZdDBItWmUlFShFjt0x32fpMt5+yGX/yY1dsDnTlk8
TxLOHO3Sn65EOPvEtMhZ88sjV1TjjSNDXSyz4puzKpTs8+BY/gPR57lH0r41YqaH
gcvA2+spkjODAGVttpDGJoVEQ23qxmrGV8GBWsxV7FcabgCMYcoxPLw36ePBPbGa
5VmE2j91VJNxbBEeYLz1QHAHXApZkAGhNvgks9kTA0Ngetqek3N7ua3Wb2543Zlj
QXPlXHcP8vTzN1ACJBemrYnBOlX1SJ+TU+E8lItx4YLPLm6twrAVj3qVzB3JR1do
19kt7k8TfJUtmXBEQzvos45M1UFU0u8VQCb5uSthogw7UYSQ8Q7qUU0u+7PAMSN/
U2I0/8Ku0y2Hh/Ip2Qy5bjK2qXs6+2FdjzZCYiKGk0m5kyzHboCkiJaMK+53vQ/r
1hlEcxz3IggLglg03acVoXDtVmrzCHvQ7BxvGJGOMhXdZC9C+HhnnI3UbdHzG9xi
LlP0L//cE74Ep904f7U68lZebMLC7EmMC+AaZvTWRcnOlzZUOqj+lm5ynM64dTs3
D9dFXO0EIqGXodo82EtTlsXtS8BXnYFmxIqt7IrHawq4+5nyd4oYJGPA0gj5Fx3J
kPSUwQAtXkXtFcmZ+AgZRnw+B7DAY+MxCuDcKIWJ9H6gGxqa9FQnMFleNfuO0V1+
TlI0xFiuGTwq6UUP66w/+7DACG4cuaU9yV9nClmwyRKnD/ZJOxmWKQfG1XBjapfw
7u2/xqqxvGG1yOEk4lD2uO4uQYDbA4gd8ApZO3+IrNtKCc9aF6Jjd3V/mY90laK5
0IFIxmJ2LQmv+tBSz08PHKBNEQyRUIR7gLPgDYsTgECX+KIbwl9nVOks4vvEUTQW
WHgneZ/QPMpd7IImyYAXh/a3y7oAWiJLHej7xXsLcwOy2E7mX3d+OznC3rcF4TPB
2ZHJ1s2ordK4aTbSDUDqH71SRUBnznkeMcj//lonR8VJLTM+bcP3MD8/SjLe924n
LyoxNk1OFjFX/8916U/wci16PKsqyHO9gJUP0rFqriMTNWqpUo/ZszQltYsfvpEt
zJ3GjH92a/7L0+de9lQpgZrIbp75oDOO/kMiaKre8EQJekgdzpHfypTqiFh7OEBk
AxyPWX670FJrU8YNsV1K00FfyWVuB+KgwjqdkJx1yytBOmbxeBbpY8DA9TiFKKb/
JxsHChU2jGX2yctmG8Y+HqllTv77GouV9MJyKNhm6C+5wdkoo6YGh612gUtQjktU
aK2g30VnxPI4was/tVKzKGyLSSM5MHCcpQReIOPMGISsz4jxG1cMT5M1JEu6ewBd
ebPzwaNjAH0HGHxu7dgi7AP9AylSfvry5ZlvKhaU7Al2HGki+ctN3utERZ25IVDG
rfriFqYRTkeFzjbK5w6ryQ1TU2w1usgZxzuiggofTlj9LewPrYTyzt/9r9SzuBRy
df7lwOg5kIYvYwwkfgb/2GVtzBONB3VaQsf5P+vKrLRgTfWH8BQdrOFq4Bu/LZP+
/axGJDDqzi0EziKmawqkam6YGNLdh30oYCDMzLaVmjP0hQocHjc/OjYELO4w6h2v
+Rq7OJ3UJAGn8Jb9Sbx/HQqsYYBPl0/ZXMl5O0a60dsSOfiIwmscE49yMs9ZKxWW
DZFIE0aPssV2YhbnOML1Fm5X0B4Hq9QqmyhCQhR9nQJkJERXdaTIZ677LunFjumy
SpRGtHNzyIpqiyftJi6cqLITo2vKWjOANBqjkElIt5fgWZUvXI696/8tmfZBfdEY
FCjE53uVaQDhvIoDWDkFKi9nisE6eyu/5szxjqoZ6jz3p4IW+XObO4DJxh8cwuxA
KT7l2pacWVOtMb1x4BV2FyS3b+jc9cNdKMDesdfPAF4NBTglH0vSbdOq4vx1BV72
p48KKEHB6KA4Hzd7+YEc6CusorefhFq3Ha5PNAHQcx5Z8IX7mt3vVYgYMJDGkIce
KclZ1ZaNNxRrJAxBDqBBRBwJonACk9Nmpu8ZBRBoxPG/33JHIZlDli/skUEU7Wgl
7MXSML2fFGj24aB0zNFpIkpxZVT2IqnUqA5lOcEuK9VZDvoREtWc2Ej8VbFrfEwr
eUjf7TExu6pqe1AJ5zvUc3JPVn/eszL3feSZr8PIpI1gh1jSJcxNOrxs/YK8yg04
XjgfRapvBLiKd3EP5bRmdFyy2E06BVPXchsfyYZUw470y1/248f+pa5MkPAEPCXb
IuU39slRWw37py/WNur3fM1NE5DwpOH4tyc7VslXZ8KJauw8jwNDSw7ABTNzD57z
Bc27L94kIuTcCZQkCc3BR0KkRHxjuK3fx9bN3HIgPI8P2i+vpbgQpOxMoZKmI+Xw
Aoo2ne0nL1OqessGFriLA3oNTGBjqrvIw/fwyQxnW1tb5XteYZOn+bLGIxl7BzD0
TTooHX1WSv4xW3YqQdP95beLlol7Xe0u9SEkf8psnO1IVGcXhw/NRuw0ZXeOYnob
GbSHraJv6R05R44jrsriL+6GWx3tBKjUlKqQ6kv9b/H2HHLJ1jaX3tawmA+ddp8W
Q3r4dCAIwZInk+kRgjylVBySGdgfkXc9C4rSeMdV4A5n+CYePOojUxTq6hmaHG1R
zYPqF33wioyClfxORjS3xrel2ncr1FKDzLWMAkWz5A859gjnPgo+2s1gvO6MOWsI
k0jf96jou/0pJlsKGhx89lARQUNsAEaC5BtqydSymNmXbYfwyCRXFHuSz2TiL2wY
olSTEhDgqcaqbdHW6ZSrcu3ATIEga4Jkk5XykHN4Ru/2cWA85NLhXnCybloxWJVz
cF0/D33gMDl7BbyuWJbuTEuM7WfooKIclbdGIIeNqaEefx7OnJeFJdn26ER0crNf
WzBLZvEO7jRqlwADngIK455tFNLtEkC4DmFwEInSKZPJwyPn7R2hqbnaAb/Nm9qH
mlQnlMtywvGNZcAlXHq4cTXrr3pILJIMn7vZSS+n6xFTo1b5aDiqzLH2BWY14Y45
kvBiLeVtnt7J8jiERZYi9eMtSmbbxhWLhgCkm6yvojJKT9+U4sVUP0dHw6BH4+45
TryrpX3MUTrsnySU304tu9j09SJ7//LhHDDBs3paVPUE/2cde2P6Rtet5UIvSVxE
4f6144Cp3H6lm3AGpLM/dVVu3naUAqvYNb0BVSQC96kni5ofssJyIUpQrbxIxltm
1XzhL5qBi6Nw2oFYqithtyEprhSUeSIRy52pqvOZq8VKozodpHBBwcHpC7TlMBGc
MEiW8iHDaNHkk507o50k8orHNzKRRc+ZunjzvHgPk6iZvCIdJeGQ9niLV5ohoLgN
klZw+aoOiNy+SWrZTcE1FaNz962ugfVfIEWoPlt/f+Ghv2q8nZUoCCy1uQ6BPOEr
qdbQF59UXgoQl0CevVKx1J+MPJGQIszyFwEh1MoaLVvj46hXJrLiYeaAdaeSXy3i
CFLSoJwkYnngdSqdBBgq+14a75xSKI/Z1zZfmLjPedNyz6oX+H2pyzdTJvdu1Sn0
/QxQNm7+JrKi86bLapL8JmwBATxtcwl8dYIRhl9Xx0PKiOKdZJHyWxk+ws2ss8nk
TYPX+y04W4G99mGOVp1oZLXi4IUTNkGMo2KBn73gw8ee389nX+xTBRV9d7AgIaSC
uvAagIU+JO6ew9oaWkmh2YZUjwr7zqg9k4C1Y7u34h3MgDENEl9SUcFcz4lFI2gZ
KSd7DpSgy9JrOVG+ndAxXbEMqq5ZwvcaomQcgSGoSUFoMyN5uWiPfa2iVvJ0D00l
4an8K0nU840jlQH7EBHXWRN3CFm6fPNJ0BvBlYkBGpGUCZPXDESOLhu0wU0acs/8
2jmM0pi8VHObq/vhvMCsAnJLFK8ptF18X/kQLsyqNk44ZaasLR95CawBSyrhrLql
V9VlKwh3Xcb/0cyMPtSqPF74PW9DWsq+nhddptKeMKMaXgqzhpl8T2cKzFI8P1dO
R+wPa7y4pOL4C7Ng8GFxPKBjSD7mLTU2BISfuPhQVNB0ZR0gT8PPjUbTnVZKxX6j
EyUOb1SfSasodhxQ45TzR2fqhkyrzx9q6jpa15zhBNyvMIvpN+TEerdhXTb8BZlN
hxWg0Sl3H/j4IT7Oa5fxMUo9nqZtd4ZE/8XY2meL/Z+gHFfDNTGJEzQp/hhGEe0q
HZokJuQpW1OjPuHKjXqEEk9e2Xau9AtiWFA163C4sPs1x1RS0xzEb+r2DsuBR/Yt
S2pFj2iWkQ4qAx9CClyqU7pXRylhICMIEyGoJjpmRbJclysxAGkdNgIGTnKso++J
qYA53/QTzKy9xEoFah+Lb+QrIZjhgN+ScecKYOoOeSBht04LS0/pScVW4TtB9L+Q
dU3yqLTL/k017qF0+uUtnUu4ZRCQLqhPvS5wF5UEFqVXFyR+Ldw/nVNRwL8f+ZJV
ApiijgIfwjgdLewaEXPOe7/12WzrhV8RM5eNwNs+wFXyuSTzw86e0WpVg/pNT5ro
FlVLjhCFrO9CxVxbp9ZaLvK1awlA1/tnAQA1NJFMjZ9tSJ3ExVAmD8ubDXutzuaJ
tBBSFR7Hl3xaWUP+qIgFlPWdFN+xFROvutTqqGr1asYJLMzs69Zfvw27ebfzB7OT
9uLeJIFAVRJgAqVI4q+qX4kClop5Q4t2uwm/cRjM+m72Kcr5vRC5W2WxKzsZeYm7
zGp0+xiRJ4YjUrn1Q6YQq6a4I41NPiOdhnIu2JrLNWM9m7veWcOQ2GTfkeyf3yiN
rS6o111ghz63eqGjXNYkRCN7ytJ8nniQIyjhJQi5PPduSwMIx2orbm+TUWAkKl3P
3Xr2H+CFke1HXSjxo6TtEOHcKg1oLLC9jk0hIh81lKctyMDx185X8JR8oLhkJThY
1Cf77IxS/FkhY6K9y9c+Ss6ztOfw8XHea5Gu/KUol56M3ImnW3aT7nflOD1tLLgw
YE9IgqQTviwupK6KSi2blQzX0N01ROK8h3r5YP8H0TZSNXFVe8DJNyuT+eLna4Tq
MI1RX4elFBbTCaxnorXkKueoJq8wrsvZNCWg7V28dW1RfPQFYBBjqJIZcjFv486F
saqLueJddBEVL/NN68pZnSd7/IFjrhLwlaWsB1qtrnZckvBGrUOXWRotoN/yh/97
R+3kx9ci1S4w37Jmq2f7I3j9279jSgQsCynoKJxwr4hqgun3m9fS1cg69HoIbGHI
K6mwDMtHbd5grzEhB0+SBwCelZz8mbc5iSh1EkDCOcU/lmnyT8qE/+1v6ct4+Dez
X1m5Ag9A57uX8P5PwE2ri/hG7tG/VklJaZcOKUy4SNGp8vY1GorWm/mD931nqRu2
Tm808C+r9hym5fiT57aqdpihF/a17x4o3Uys/buafuuun4toVCIVQCX4rwubni9p
0iRiXtzDzka+pYlktXIYRL4vZGMKHHXZkROF464I/dBps3ZSeWqj//YDlQdk+idk
hkUKnp7+T+R0l5ZheGcuYDyk4UYhOJhUvit4P5Q4D8kakv9qYlUwph3syKbRfOwf
+w1msi7MT/1AqtFLrTKEIbdzAcce1clcHGAdr8e7r782GFBP7gfFquQ2GrV0lNld
c8OReXuj/AvfJ4/MrTYYG2QCXGNrQ/BDKD9f0Yc5cK33+fMClohQyrghdIrK5129
HBu4RSX3CHsGg6LTt9/NLRW9Czz+UWqtm+YynRzjWuzE1Dwc+Fbj378t3z+APjHF
DuIKwCd6shUs9iykk68+kx6mHtuRuWLmtEzYfcQkBJDXl6AsL7w241JoDt/x3pmt
085WBvXUFAMDSmGSbxyjmVGkX1wL89J5ptM0bJlxf60FN67GCc4bM1dM2MceYSJr
P9EJcOPYZnvkZKqem/EGu+S3sXlxNRGrG0G5/3GYQkw7WSfEINOiSXOGHZ/d/v3n
zeT4ruvHj+HV4owjYnyoCwMNcRR6HCv/d1a2dN3+01Fee6nCi8luNaM46x6gwH7X
vZALPCT68jCLOyH6c26ADRHznM8bxEBPPk/Y8yLj4mOiAT9yx2obIcyJ6ha32Laf
OrNY5R105NxrUIRWhW3y70dufIMKqqjNNkreBm0W59wGUFL2g+QTisWFj/OV1/6W
Byskh/unoDEn8Sqn4Gk9/Hft2pbGTc8aykaQZS/PNU+GVzGz8P03Qm3VPnC3LYeU
ePj6vPpMXpoXQX70uWiAid0cUqhsrUTM+e9ZfNjDYYuaFHS/Y+dC2mcIdjTjYA7T
dOwwc0JvTQYG82yNxM1sFN2z0lQ7ei5eG/JQt5LrRx6odKIto20S6DgcMg1fBU58
bslCqw1SdVTIn2uS3CRLQAjn2agAPJCntxR9ayOiRIUQFWDgkAdUWh09soASv0XH
dn+3ZuIOUYZxHwGV9cEAmiLAuHAPblVNcSC5vogMxZi7fNpzLABne7pshpyDh4NQ
JfxPfVpJqkSdiLJBcOmYFdxNzKX4eD9DH+3vaA2A2Qy80UbVp2glHo9Be+ZEcwfk
kOpwKCcPb/OePyLdZKczH2NnvCZZrVKDRCsnCwtTZxLZDkK/plU5a4Gr9LmWD2Q2
uijVKoFUn/ADdhjoRvVXyZ039TqjjV1zEAQHiMCizIs/zC3XoYx+koDr7LGmKsXw
vjajN/W5Gldm70U18LBcI1i2SqhJtksXyxt4uBtRcTWzRPKljeutKdzhEJqTvZKo
d6iyNofNvKYPoMthwql6/DHHwQn/SY8ZoX/RDuoU2yD1rfaHnHnCLfbWvuGukKLu
s+bQvsRU1NJEAjrmMa0gzrrcoPnq8mG7exX5UDvauD/M15zpg4nKKuTDtIjG4wyY
AHJJTiVGYXtpDH8LHtlFdsTWL0aJd82SmFjj7f48IfNVer0wJsCrEf+5O4SY88cL
T3OjqttTo1WbkzTtyibx03+QCN3UWEvF7hqYVYRUJnGmRsDip32yfYMR7pt+KlLU
49AgBpiMD9Uw4qSdNUijUB7E5hGh3NDfZfnGYSE5UUW4szk/UFY0gQ/eaTVu5s8K
VToYbQz36UXrZyFMYC66BFFS3v8QtfOjdmD4P7++GvhaFtmHxnFk1+Zdih0Ael4W
G3tBiwvf6Yf29L3EALK6PSIVTRUaLQiRSyhjnHfQJ0P2SDjwLRaP/UY1ucnVhCbB
L/pI5XJm3XoQa3Pnaw9I1H/Yd3YmlIJ/oj2L3lnp6hxxfOGTLegCVfRuQqBoIcbB
6yImPfM0yw6RXLxRT7TsW4FVsyOgfWb3PiG51nOrRniqOWgpk6/VRRd/a4EGpxnv
nxLxvzBLYYCrDChIy9tarzxnGX6xuMCg9zEaSoYDLsRAZMIjRywjWC1iZ8MEsPZq
xFwypYRihBrVBETLGA1+9WZXv2fAzJVIDgAXvnd+/eRpYyYW2H6KNbZyJKVS7om1
soMTQVH3fK7/uM1nKMTsT+zNIfvJ+JaKZJfpA9D6jdCRhQxd7ii51UuxpshFgN8c
Ku+SGtslyC7fB+DlYZYu4uN3kcsFui4K7xSA1c+94YGojWMAQAfD7H4Wp9yEYYNf
nKdNgPoq2+YTXYU/DhTU2WhmeV5TiEausoLHnOgUesp0t281d7v44Tdqlj/ZVAd9
FagJ49Wvs4nwtXNiJhCYFOB1jsOnRAxIboIPMNOXdhyEujxSPf96Fg1T4tpJ3QmP
V1AesojObSbL95EN5tFA9X400Um4ObLnMbEMGQ8pByjM1j1b8Cuw43+dw/zDz/dc
Yr6TFjBl/VOa+K+7APz+b7u/u9t8gXNHhXxAtU9FBXWG9SDSjxe9GrZkP8xfipQi
9qzgJS9E+AhJhev2Yxnvm/VQagmSIxe3YWNFd/5K9kRwgIRJbBPvz08trFpj7yg5
pHaXOMthB1xxyh5P5g/mj0kjwD54OBlUElZYlFTwIGVwr7Ph6vwW6YDRTujF3Ndg
P+vu5JxYw8qLadmhXP+Bj0vtyceWUhFV3oAMC464XMt9RxkGvQ82fWVTuyvmKJPa
zfi3t0bQvORESlSuxO1ZQZv5olTmg7bBmSvYWBR9PE3Jiz8VOk0EFiDngf/TWGw5
azg0Sja61CI3OXA/k3tnVqXxATAEyAjbth9lDgd71ka8dgrn5w2pgDme/4xORKF4
Nm2hExgfBjiHzzlWRpBvpAe3Nz30IeRBMkjWlEJtiaDglVI4fqpodHUFL28f2a69
PSfwYGqoAP+d4ZBcqpYHWxwcXy3GN5wUH6EmmtT5BWJ9wWiKI7TSu6KYaaekMzx6
8VWCvW3Oihr5Oh3aKUwPLiPrrsBsICQIDoPrUA4tNFMm9IfU5RxLc8aXysCEIi1f
aWUUoaOhAJL0R7ekTWfX0YSmSQxb1/onAUdck6PTs/8qhtPHi5fAIw77P6Pba+/4
rDpFvbs8ad40ZxOmXhdBdUYfchCLAoTBbNGgkC9wDM3lv8wL1WB3Ss8YhEtrFQ9P
8TUiWwD5GqBBFGihMETiI535G1NIEpQfUPnqmWFGc+JW+VkBJ6xsudhL9KR1W5bi
Z/db1KZv8+HvR95b37vr5KRQEPV1y0n81rbIKnL1mCu97rGBQqR0gDlhWhjHZQey
AwoV28Lahsx1bMg+BlUo5gm+CpRlBSHLjpf72ElMQY5CwUJ31s3l7cb/lnxMxAsq
6xPHUV7Ic7vjGKJtYSUobM96syLO8nGzc5zkbX0mrceF0Q2jnoviOLW4WpKOD4Q+
Zq74is1pudRHFKJThs9zgSByqYHuvaovKkDmBgPRz7rihMakAVaCW0FOd8pEoVdO
NsyTRD0Qa5tvD1nLf9MyXjZ7Xbk91LALjqte8jv59EAm9/Et2SzHrazGqFw52UTq
BaWAlF/LB6CHp5HyJbrJwDDeSvgyQ0OFNiTzYd+1fl1JzEsX+/Vr9/t+4GNqhGeE
dXmbKUI7rWxqRsZ4T1a4txQVoWIQnPJkEXgkllqw7J0Z6B/p1ofD5LaPJUQ4323w
dKmnzlB3x9gcX2+95bEWfSxgxNojILXFjSeTjsIZahL4eRZYLoajCEwnDRVPLVkS
Yq+e2QnqBiuS7YTH6eiHOqsunHc2CYhnM59+zwaMtisM/bNhsoTVva1tl2lTvXUl
YhDN4VdSr85n41hCIevfFzOrISOF59r8BwBMxXLFdWKxQOmTjSvcwV+lFCuo0zml
4stTVW57ahznF1syi5pAsotIXk39o40iGk+WL1Yl9q3ISk1muRhTQpaQoFU0BZue
GxmIl339fdFyvIyPIrKhqz+bK9ByFpfeIwelU6qJYuSbiU7KHc1AQmQxJF3QMpyi
FigefGv0uQlEYSVW+/IFtEVyCIN0BHehQ3hbK3vJ/4nYZ0lotKlnAOF9MQivNUQt
lC0p2BblxPBEiGYjtBjacgg5YehYUckAYwJokEchm0W22+esvipPd6LhSCt4h8KA
Iuf3l7jwcN6TgQI49PisNRlA+VkjxVUTG5Wh5uES0p6RbRYvaRrAS6K1S5ANuyRL
536YTv4eUa73yZMTp8nO7At3/3Zrvm0TfwOuMWY6V5bzcJiqCNGZkebeheCdEu9d
7J+rwIBFbUXxtDARYRJvUkE5By9i5uFvWsHhHo5Kj7/uiRr4i5YXMLSLk6dqb3VB
7ggYzDlyWXO/X/aPK7vr9bgjJpzu5I9N0EBM5LivhpIAFQHW5grJs9iVOFN9JX+C
DDsR5UOhE225LNsCFTx4DRp8FkHEfL58g6+9Dare6hCFpLTQKv1H1rPTxM6W4xhz
LDeYL5TT7VLDgzLL1mnEsCFpXFuVZDKcktlK5K5vFgsc5HrO6LUqrjoLeTL4prc9
S3uX4zloVhOTDp5q2TLJZ+0vbdDalfuyAisdtiEUL1HMcWhTT6M1LOyjsYRJvjC8
KuUZUMSo1/LJHij/ZiC4ZL3HRGq194YL3wcnT2JpcCm/cR1rPPfU5p7GiuWfVwB8
OOdiUF6qgqvpJZcrjA6gxTYVCajBbcYOoELiH3IJ1iRgOfXxmCYUa67vg94t00A1
KOG8wzjiYu5nebUTHqMbCRanf1kbS6nzXuFwL37wn1UMj30h5pRJnaSHvfaDBtP6
xwMD+RoKlXjqjDflR/WzchvvM2A/5WV4MniBZzNhe9EhFsEYeMDoo2gozm7T2QF6
eqpG2T+gF4CiOb5RWXQogEfLf+x4xqdoUzEJ0U9skNSeqp+qGYshOnesVA8SuAX5
HxU6ynePcI2hHsQRLxPRWvPsBsj7lWzyoZRRSlwGvKl27hK7u1ykVLhERd3+8tLU
z9pkbfXttVL8CWLPzt3L43vIMTweNjcje49u2zv8/+3QmsYdkjWryFShL5MRhyGq
he09qSD63rgVstsuDO1YGo31P37084+QWlgU6ohBR5LyY5SvcHZaCLqe5fPOsiP3
LFFOMiLQVNWJ4tAexa5Fy+V59OADk9pVcImJKgQHtRPlmEW4wAL+Q4HXdHTYuTi5
GbZ/940gtrw+hBKH9Q5WMBOC73ZD1wBMLMHgCO9WiXjamGIQ42CW5Wt4BLUobgCH
BL9xB5PMx4Lv/tPdtdWOzArE0zq3GXK6COpZQ9YDhGFyQLExukUy8lwt3HOcRQhw
68Qsp5JwYKCKjsHY6+x3R1dTW6vm0xoHKs6PTQPD5XZ9F2UUMJJx6QzQtgPiPPEa
R7etVEmMA35agFsomlCSbCEPSrKxEee+eT+6Oa2/aoDuu9rvavF7dB4uKeRa7X7X
1CkNaNq/F8tFNt14jvCF7mnF8hY1dScF5DuY1Qw8yTdp4cDsOV6SrAs29h6jfjvt
eHdr0S4QZhehIrW4E0bAqkDZglRUhbMQXBmD4WYvxJZitbBkHhE/Ub3OtXFF0MnX
Ly30luWz8ZQHnuyIHnxzNiE0BWys8s1UtN708z+UXJ0U8mZcj4UVYFqectAeRAM8
NiNlRHKBhSd5JjcVMxP1oAE08MqvIG+tkpcT1mG9QmlL5FH3OtCotJ7I9AiBysCe
LsQnJ6ESXFc8UHVYBeoYperBpPFWsuVz17JE7CsZIkuqhk/UCUN2b+Fa4byiuIkh
6+Gryswv5L9ntrywRX3lPjPkBrvwmEUKgTfXiM4UpOLF8/XcKWbkAWMlZFqaYi1e
rjywlaa7RCnQbIyiKIvDuFQnQ3t1IhNH18hAlE3oItgLLB/XldIymQUk4kFpqSSo
8TBLjJtQ5hPIDkbktnu3Kk09PbPC4igMbN0KkRULk40RfTbYFbhFGbctpfvyvgcT
a+AGkUt9XMYhB8wj6dbtvmQ8so6JRs1tgJrjdWy1fpIRBVOq7CExbu7bKVaiHE1B
Jmrm0ReNK0pdRfy8QfwsqUQA0/rO6Zg9DaXLbpnKlBqC2Oyw4B9KynSXKS2LOfr8
PCIX6GsR8TCagpt5h3Vd/2o4pmmTPcFY3G/jbSKmBZiT6Ph2nBP3hDiRkZxfCngC
RUnSRb34oT/qi13QRaPAnFJf4yJ/m9dC1//DEWaU1hzAC7xG92+WURXxMOvZmZLZ
GfWDYaLAnsCBmTQcJyguOeP4rC2WmPNGw0fNS0oOflyZkQh+HKgHg4ZTjfh1MQlh
+WI2DKbs7nGtsYJc0C+/v6jj6TrElvfnBsu7I8RFTY6VFCb66bhCj95uSY13wUsk
SLj/W+12L3D4Gjn40JmGEVCRYRAsUiQ5gnlz44V+x4/jn8rWzgfOo/rxkeIizsPQ
HORTpPNP5DbZet1reMFwHXmgw1rt1g7KMfWJw4VyjGxp4VVWGPk/SYI0/Xpp/71v
26XZK4Oz4rBLSsxvmnamAoMVJrDCDOdXO7S69d6O/vOJ5KdDTQls8lRPvANciHIy
8JNfUSc+kbxfgOrPF2ZVl333OVTW4uLWYk1f9QATBegSfiD1R3IZF8hWBJYW+KBy
SiJbcErNmgBUWFjceoXXSlU2CHaRrdP92AUJJ9FPtvwFR4degIbR1F9QJHgFnjhd
VXw2X6g+O0bRoaOYO6Lr/Ni0rVOngmFRxL0dOYXbX+QupKfkR4514lHmFSwNrkMX
1f0BjWCm2nbH4tyf/036r8gzxsq5CaHlSMrV65oijboYey15IneWl3qn9K/2ObkA
hPYVAQBs21RF8dWyiuUci+qN4svvi4Yj0KZuKS8cyETMWG/WkLBFdj9W4mn4+/I0
L8NaavVVpnrqACxiRRnawmlgRKh1/rPBiY9nMFJ69E8yj4hABtkPDTW/55DzOpAK
6Fyui0AW2L1HyktDswXDmVDvsGPYRR846rn48tvvZlynXcTtwxtsOPkbvGtGsb1O
xPhgZO/ysfoapj3uqOjHfQQGTJ+y2vJuDTGNgV70euU8AaDUyAoYx6EMOglWMPZ5
eqKMOjJdzCR2q7QlyyQIgppY97WdqRZC3qJgqJ7jWhapoPvOCwV1EYxB24OHD8h1
1HmMviw9qJ4rHEYcqeuZJSw0jjQQDOhe8D7BVJNVnYpeJVAC06O2GSHoxYSXccYU
D1c7mwS7uTAZ8bNkv4mKB+yJWjzc80o4/r7tamboG3wBKnGLIoHHlkGWB41v1t5G
ntF8FuJ7n+y7lePCvdTf8eB/SfMtxAr/or7yIQaMpQY13WdrjKyVNGplSGK/8e5/
+829A6D36w4NIcuYNu+f1Nr/jjL0hLL4l2zD02SUOt226sw+ICwsGPzSyk+cCFV6
+ixFPX4S9AXNT+B0e3FkwGqleKF6aZSSwbm87bbPYgUV4DgJy5Z96EjmLrVTvUA6
e05R+bO+YJvOE4rbNhOn7TYTZZjmGUAYotGEphKsqaSD42NF2OXOr6t4Fz8rupy6
9IKAeT21X3wqCL8ovskeiVgGc2nkOq3G6SpOQKNe0C5vGNrshCSjGFPrZoA8vRmg
IByjP8pRttTKMJL3HUmUZRV6JyIp9q8Ywe0cSVdF4yjHhG4WQNchyUppCJJLipJI
vsBx8wCZmKrF3N5yMYJ29KOREZRuKeQFr2hRqh3F+iIGCA+wdKbgKCnraG7eFEQg
MEH/tXq+ASBNDegFTkzgl3NdObmryuw4+Ri/e/NQ5qFf3lnIgVUlQZwJC7H58RE/
EBN7G6YWzUlCdkX3dRgc4rrrKfe+8ydKho9KFi6VddoAYBLqzauneo2KFCbTXufV
556ZR8eIS1uHaebl976lD2htU87yaVM01AvEleRpngbltNj61vKXkjHXqb+WJRAW
fm8we1d20OeV7Hz3ir1Bb+8VgtJ1MPsEP5QpP1tCMsScOfOdyZZfoAAfihotcSSn
133nBQ4OxhAwesIB16Ot+Nt1uvmjHXpnaaSo5bjnTZth7y2kkEddXCStR2L+n37O
cQNRWmvzEZf823j/yWRlBndfbJNcyNNl2ncgUvbExfBcaTYyc0ak8IsgcYjh2P6r
pviHHOCF6pdkrukJXonWDQfOD7AVSrMcRaiPtQmAS6jJgMym4rP7kbW8Z2WpqXZJ
JkbLQFmPwcbSDpJUWwsJjLNIMWq1CnesawPPuGcvjoI9uFGkL5k/rG5njTTLhK1B
MHCUQaaD8bHnalTVV1zYGj4pK6upDkyr2SEGPYqjsEAqr0+owXZgJyScMVXRrPSt
aqSAEE4wWYJnJVmhz4QVmAf9XxnwfBp+klxdG6dvxiRuVj5RBdPexUBtNfDTbD/f
RRrB52lIpFehN5oiIOGLrxDmUAoWu49fg6iPWWZzRsuJP4pHH7zcuPGEMVzZaI4V
rRk1DrW2rh0T9FBsGzstHAWSi9VZxT6+S5Kelb3mQx7007XMGNW4uHMo1K+j4Ktg
n94pWSdqAJPx2N/UeVrxXDpIHUxRHgUNMXZ8hoDkczPpV1j3xFAlRdN9z5rUzX5H
c0vryuarH/oodq82t9E0V6cjaBOE52pJmgyUkNoQ/fmeeYpIWf7lEf5VzJrQYXPM
qT6DTaw9vJYbanT/lv3SwISsiFXcoyfNwBKebHVKjfBVHksE+k8jDFq0pVi+b5kH
QrJEA+p9v8a6JQgzh/Tuip4i9tFVLwf5kEbHt5hAvMqdr/ff2kC2Jmadf5iCUc25
QsxqOHsPOUXwiJFMbs1c6pc7uDv+6Jl2gnXGS0f5Z2ZG2KNwP2aovSuXdapco/Ms
CNbSr2KwumF2uvh+C2HZmzLXCu8JJCvn/vNBUJLzoTeSmSsj65O0DfBmupU1Egtn
KMbwlsYTynNri0FVa5jr8MQ97VxyGfWOFs3um13rFyXYXKye4KrUdqElO1AmoBG1
HP9kCBlU2g9/9GhYlVldxx9ifL9038KjsjdNHmhPKy6/MuX4wgDLKbo84ie0WfFv
CPlB8j/vHIj6o0khQuERHOQcb3FSyaWs59iKvPu3NhEiLiCAZRly4+YFi8iWF2hx
dFTDB5ANkAuWeTwoIFzCqEAn8a35xvVJW2ZtLSNhHoCmp2M49YKgkeVVAaqrCEGH
jRQNaAC/Jdnn4MccTbXFss5SoL/y/cYtDiKu5OHDg2BR/Kl6S+22ZT5b31p/1/tB
GLugpnpX7hou7T++64EvX4IEvmkBPHj1cw0FJDB0J5KW+WwR9JoR58jSKfislkJZ
Iy0JqJxefTD/8QGh9ucUlDQ+xQ6PdpXalGYttL4Ol9/4PCbyU3Xvun5WoQisv2t+
PK2VkZ4mECTbP65iX6D5LLCzBcl79f/xCugqw72cAFal4p+t9szN3ccH8pj3XAsW
tojZ99PCEoDjkG1/PIFoY+R+VcKxQhH+7WaozVODso08eC4qUNL3UQLpVHiCLC8K
hL0HmdrQecPtxB8RHq+1dt4hNKric4PJajlnsPXFkinBPbjWOUpbqVXWhbqVPMkp
rXxKLgEmGLlGGwqp8DcHwWoZxYsTgF7bx8dVEhv+bfdHM2NWlt8Yil6l4OWW8W78
7zeeVhPb1E9GgTATilDinfeO5Ryd+y1vEHe3aonD24K8VkrL/Y3FfeHk3pCUFdEE
s6sLkRu337gKj9BNe3EY89BSb94uC0kzc7j42Aa/kZ9M/bkb7uMx69usaud5tPtu
jyP9jNQeaOzoG69RBt89xTyH30om1lyHUn8SF3dMsF7Wfaq8hb8g9PJF18fiEj9C
BjNPTDBME1pFzXB6bHOdc9hJAvzS+a4wMSb+CLLp2cf8c1UYCi0DlksCf5s2y2K0
jP2wuzcD2JJNNaevqSifQqhx1KOh/wp6+Ovi81XMmIXOoe08mkvWRXLIRWXch9xx
OJ7NEeN26Sem1oghsCTsbBpWHhedNIz7Z/np+q4aW7gpdX9OWBLhnn32Iz9/YIVG
/m2tSPMPq6Ae4diIo6nUTlibiQyQxkjxC4buUb9fXzn+jvOASUerunGiXvSb4gG5
zLUKfpGL5nLhWgL6Jpr8iMvqk0Gorfp73D8GzMAlAVtaPlYzMWSjZ+f6zH1t3NHt
zKiQRdr8jXyrdBDCnJk1tkKVOdyN6jyZRkLrCP9vOXI3uFeRdy4ms6Xvnz3+T56T
YOxxNxwTYFF7yRhTACMhwz6Ff2MNpb52ILvP5K9jvRvAq7MnRIF+BKGpHXtiWVSr
IP9/cqkunAYvQ1NWSD2XHAg5VCVmkXdDJBmj5HNs2DjVxRuB06hI5r92VwK88vc7
nuwo0hrOoABQ+R+u+e4qiwnQJMjorx+I4RkZG6LPN8gAQ1UbUKmuAJMbbileoQBd
XKk4csCygwH8kvVR3FFO+3bCiI+KDUr3hvtkWItQm+70HJe6zxj4b3T6yl5yFV2g
ikYsoTAcZ5O7BakUukpqDB0A8/s8sdST/WYh8S0CZ1A1agdug//UWMqLpbtGtMdW
S3Ir+/Jb2P05pRLxEmoIZBIt2ONdDDIXdwMfuXVw6/DRc81Cjg47Jjq1bFjlqdB2
jRBsC7aaHy1l3h0vYEnty7/RLurSYKaCPBUny+6gJeRjyqfSgF7QlrHem+X3GTaU
o4uUW5PQTQYTVihWX49Ad7C/+orLCjcAsySYyDXy4J/BeLBLqusJeN5/r0nVK+b3
GABZEha1FNvO+wzInFA8/a5lqpWr419o4QY6xfsUMXaJgeJ7IDNT5kxKJ9JT40Ll
4JzY3+QkAohadBJrugzlkOlgBUVmRS9bQ1lSWkw1sTyOAsREXYXaUiPf+IAqTwJP
dcOA3ZsjBwdNF34GSTSWzNTGQOnIxFdikWhCJZunqOTEvLZJRJ6/a7aZGC5KQGWK
dBvp12cApo6WOjtsDf3DfxeqCEdk4mn/8VVVWAqm2xbUOatcbMiuokczHQU35Wsy
iyno6vbDsp2ZlxAyFYW6/iPBvAs6mCeor0NzQVFJvdrmFSr/+iS9k6NrMbvi17bG
DUEyvEjNVplSjRk0ZZLuB/PBRcX8Rrqw8wIQS4hYTVgaG/gtgU0WAGPi7RWOo0V3
5dBoYjBTQTVprwJvxRk2u03OPU/u6JYGgae5ZXQ08CLpkQReClA2Gw6JPMjISm/6
7cWp08HT7mstMp+ZmMmtU7Oven+Sv20AaflfBZ/ewqsSFptJ5lO+AVENcggF4MVf
wlMhGBMJW9xo6fL2HPomFOqNIUbD/kNo6L7v623PDabbKsw61Wa40Qz6arjYJbYJ
v/LBo1blPnxKc0MeQ3UNuiPrRMsBTZayTM2Ron2NHYNds2IXmfJCepAph9e60WyD
L/ltDwY6t39kFzNlYLhzefaswZG9T9hbtsQQFp+BJ+fKRVic3bVhjRRlh8yBTYPo
nXBJ5lvd2DA3GVvldtPTKo4LjQf0GxO8ZG+82u+mU/EcEDNMOSZU53rRFJ9NGSnA
Dp8Z+RQAX6LDtmMKCkvSP0QxIqHbh72z2oOMcRJTg+HjIJeHbBYC4vDIYvZV8hox
RRKflWZAhEV2F++guGWunq56Tz4M11U7Mm7jqSxqoca1GOTKd8WJr2rFCVFLmECc
iq6LQNBFLc7hx6h0UP4VMOTi32zoihDsGXuNi0iqWKfXk9zOSqw72JETkmuPM/HI
DJl3tehb8bIsOfaqkaFAfzQkXFglBHtW6YzFvmJSkue3sG3tAL6usYe7uWvyc/pt
DuEDAIvMFGhJVJnK1bqsh+er227oxo1Ch12z5inT5SRtFJ9TCYNW+WLYaJZn5HUJ
aJtBy1Jzt0NvI8RTh1zzkCq0ZT6sGhe/gnL8JuXUXWkbwb5csNKbULebraeEpmG1
xL3LB5Vrkh7i4HBvdS2AWjy8e2eXpn6HBIX9u7yv2jUT1hwQpqELD0oVkW8nbBC5
+TgmXz0AmPm1qMWcD7eC3UIEipomAHWdCUeLks+pVXiPQWmSt+LsXESCqHEml3yW
w8kQoROcm3T+hfaCAxVhxAI/AXzrgaVihfswakSokQQpKBr/e+chnFOMwiF9TUmT
4aAYB46l9Ap1vA5UiCFzvvbR2P8YKn5zfbfJVParUj9wrN2f6JXB6gxIyYs3jPoH
imQ1gm3LjA5zWOdKa9l528HenRtgJJI6nVnAdl9phD+LITvcLDUZEdUGemXTNE8P
pZC8xkYgbuzMsBH56e/VwScVjy9Ite7dl9FNBC9ITghbdfpR1Vcw0aq2K2eBu4+b
RpiGuHVDK0ue2CH/DX2RJS17TMMfaLNgEaL5pHRILwpnttWY2ntokkwsfGuzHa1F
P98g2+ISdYqiD5wETfBVQCVtlrGdIJSzA4wsVknz1Djok91YSNG0YDVxG4MpEsei
8W/WC/bVElpJ9VI2VlWeL7+D92JHxdjrp/5RgNzJshzaPK1MAAkrkfq/q+xXAJ67
X9ar6b6EbpaWRh33AAUew1MDSpD4Kcx/becciChPMfNjZ6dLtuZR6xCe9pvx6U3n
GEvlmDzsbecE22UBTaIGsvtGGBV40ocVMJttSEwSW5a7qTlPboRc9tDyvKE/wrsc
qF9QVBxdcxPZstIET5ps26vufKfwKJLJcIdBgEGhwnx//nsZVMgm3a11/hLO3gEu
9y/Cv3swlTRTNCUsMX05NpcjbMpB+hcSyE1xCFTpSusZXndG/hxc88oDzkb3pTNp
wp6+KwGX6+MD2j27D9CAw9DHzvQ2KK6pQ6tZ812s702rvS4G0p4TQqMLXKxDHkSR
AP2omfPqulwec8E27HapzY/1kTajaHBxAUnfq9NP37VdWzmOfZ37MeiZY1bAIyFK
mZD/x8sJSZ+eAKsACahkNIlDmQhvjpjGQ/I4UM1Gk7ZgY9miSQTeT1Zx0mbvOBEg
/hYPmHR1Xsnuit7saf6MDCCu+rIWcGGsQW504DfFzojLim17SK3dNB7MBmBRvh7A
bmGBtylpieohcw5+4N7XnGrUX/EjPkeKt1xMe+Bx9HOOS0je2b8x4OdERVcIsg+Z
JGfXSJgBxrRaIZ4e+5lxLf6sGCYEKYBWbPhVKgbhKkT8ZrQ1unlEMDZ1pYsc+FYX
7+x1sBQF0m37QX+9xkNLYIZLRhZAxMhi2CSJVhmmz6QkmtYkmTsc/O4FAeTbDW9T
kuczrbnTYjVPffDmqNNSeWXsiT8vZLTbqSWYyEidx7zPh3bSKLrmHvC3lMTYtKaH
ud+/Jgzr2DN4CGmYim5EA7yq67JUOJh2Y4KLSoGHe817ZLPlC3fi0jbR3XqrxQ88
HGEs96DZ1EIfjrZ49aoACehyJd/Uh0dOGOPMkwTjGnEQGsOjLwY6x7FQB9KpaNW6
EbXLe6HcIfUIlWvxXOO5tICLXGkTPCjlbJPw9Xy5Yx4UskF/lxnNX16ZxRGu9paG
cSIUCdL5q+UVx6T5UTqnugh5OYpKiSJ1OHgRboeB5VrZrbsTtSKXiZkpGXppj2zV
Fe3PL4JmxIcGKDXFqVRt6vMwz3Ap1GM3rW4xEeA655fxYLfzWWu+O/tAUuUjF/Hp
EyzGiSgZvR1YATxjW543apO9OT+iP0nSS2zWws8tXdvU2mD88EjHy0WQNoall2XP
XbG0CV4dGwQ2uRJkTxE/K8XO7KXw+obR7BwU34o5U7ddxD6mOXyYZRMD0m1zBjp0
v/ADdFUpkIOKcvezx72JbE/C8RGawnvwh6I2FY0VWIFkfs/RI47kxY4cBAbpPAYR
wUL+a4fknpH84MTgisomWz1Edkul+RvTYxGyVtQAh8weymrQv489AHqMjYToWwdX
eOPI6hv3HREzcAK5sxPHJiuE5T60vQ7ypaVLduwGzrnQR0NDk70tPKfOeQDR5Pmf
7Anvmeze46dpGTGyHIFdPu82GxQEw6A1CTjQGqUOaRtnDdPUnIWJ03flPeEW7Y73
QgEBAhmMXJNzA2YSQosmCsnRdSy0dk7Opbx2K1jCen0vYW1Vuaw84YGDbkx3+k74
cG10n9Rrzf9r+SbKBNqdLdOs6TL+l5YtCY4BUYyQXMhfAYTSOuSI+JfIgfQLl+1W
V+PiZI0pL5ta1ZQVXr5EkR18vuxgcr+8taVq1YASsOevtibZkaTVS/pzo+7sPWbj
7N4oTaEprXmx/nCwD+FmZ+cwmfHh2AGkeBnCFQuFJCYhhTiGy/Vdv4EuyqxMM71X
BSuwVgLFuKYI0XYVfH5xfikELH7Pkcn32096BUJgZIbIMMk10jovpfXXO+84iC6S
1eXmyFDV5VIWZlKJi79OICgbqnT2HTcxkedDKzodMi7gaJ2U2f7H+l5oxRknOP3s
SY/0YqMJkg/aLPSPlm2XXfUqZCJIlqXlGny0wKXulk7KplCgfRFWyQ7ltkSVjBdY
r0gooKZJ6VKMuf2WBEzFqkahjUIpedqPgW/377m2/nmD5MB1jH3uvvNGb8oORnvP
TbphcQg0b7LqbbEYKzn31ezpl9EXGh0bLY+iEOVT/M5HI/xSyLIeG+Em8nZ4LfTh
7QMjB7WK5UpsWHRyCbfE/xHH7RJMV1MFbtdvM5DFOZYpkNnTQIGsa7rRcXXZD5Oh
0qCNBxsSVeh9CQ5foNDKl1cHHwpoh04XDTXYUgMlnsBPzV2b5FSm8hrrFBKdiccS
412xIZPiZx+/uQIKD/aE1mJfZ4nozURGvglrHzIyBxFOWDmZlTrV30pSz5vXRv5t
lxGBCICghzroMRybVVpmZv4Du5FHXXHkFamXZVEHTsYvyljogGTT2AmN4CkiVeKh
koRy9UaNFqNixFJ1TQ7z7JA08S2txYAPt9ioaSytmKJ4Tb2YwLBWsb6MBw0gMWRU
PjR3MUmgRNsB3yVx3hD7r6JlblzwIMJ+9i3wEW4pdTqsi8u26DVZ4O0BAeRz/AhU
n5haSLqT8TpQdZOZa77u9M1eJp5j51LiQJWFn7vpwXdNipB/o+xoQDOmAv31OlMr
GKNyLuxM+g5CzvCA31vtaRGE5e+cX0UZ7ZmYBpg8G5vJYwO+MS/Vs8BptsqqyXGs
CdqfQBMA4jIJTnmxI4jpCJPGNFb7sbbjcCiALCnbMmEsqdVE4y/aVC/16urhfU0s
GLm/3x2VG137rcgTY5ZftOkIkhBC80dXmfRsZusA5sc4iTscwFzy/GxRHRCcYt17
EEfmc09H0qz1Ye2EnMIEz3s7FKEfebyrwJMFF5A7H+5WUv1+fm5M5xf0RQoIScSf
MEMcgC3756zZ0D6jpPkC2PCmCTDJTn1aQakkOUSO9+ESTy7NbpB6HnrRkuNsnb+L
+Suh5g12puGul8ihbMUC5irpNUOpTfUmnHZ9/yaoTXhlkAlwn0pw9NN3VB75hP9u
NCYiWvWUmdcOCl/dlAYA0+QXZsS0P+IL6aqPFvnBaqL5YkrWTWp1CsaSz+zUoHge
6XojVBfui5gbv0XKMVXNhIX+N7wsV4vkXn26g7pkh2mUxEg97as/IxdHZfE2n4Mo
7n3pvL3wX8X45wqzoYxB9yBWqs5x9XmR6AiXNujx5I9aiuatDSnRxiQV9PgaGnZe
yH5LhBHAmCGlpaj0vSasePYO/LqBmMUKBT7Jn4uY4IeVrshY2Ks0DRHLs0g8/2Re
9+CZlEuXVcDcEMXyCgQip2coB9JDz1NYaLZjl/iPAskdQ0j2rt4iTCjmhz6yTCMR
mNTDXtvlt90Jt1t4TsEUZrwFjcTL8VhGXn3+r2+KWrrHNN4c7aLZycXAEUGEsF1F
8yLNCAClvY5SObTAtIjlIAnDcyVP9ATDjYRgmxDMWZ96G8irGY4PGYy4AfAkWziZ
siWFcBTgp19yqfWUevwi2RbxnYJww8xbFnmm30IewWVhKx4Iz4/+FZUJK47V200D
1lUS31K7VhyyhO004XrBNeep7KHZv7eX/6RR1+ouZvmVL/3WIvbwCRFTh3sYHbS2
SFcHxesq1x0BS4Dawt8MxPencgfxQcsw5LjDxNR9e/eZ1HCBNLx6teGoMt1bgFw5
OuBHQ4h4o69wwJ10es1LrWV+Dj14SFdDtRYWYE+BCg9/C89vMkDGbuiV3jGg2OtN
YGxagFThFa0abbIBPlxDkPoQmx3AjyMBl0+jX8c96SQDuccdRTMK5bV/ROaQJGdD
zcd1E/OXsYQSNv2grnuxuNWtrl+A5KIky0CGu2NM2kvP5X4UAWWC6FE2kf4mIx20
4gAFz1p7SS3p+TUHajFpKo5kUs2HhbufeYUHjepGyTkxPRxMw94ADD2NYhvis95t
i/Z+67an4Tt8HrWdOJjhzbKi9tU2nciPc+H0KKt53/i8PyL5ceRPn0RYZKx3o5MN
PfS1bA83EGCZ6ijwuq0cVoiRZl/NzEaP23L08YXCrV4EXzM8ejgdTVS+LiVWSi81
Zko3W0iD6P6Jltg1jJN8G0o76aHmiU4yvxKWSsxwDAqUiJrUkVIsqM4AsQ/3iOVH
tDDOakCZ16a3t5QRk3OOM3YPKwOXq7WLSQoP/iSj+yscE5E44LRmgUVa0FMvq7fO
K7A/yah9tDZdEuX9IprNBOWwy+tCDFhdYqP5V7XKD/mhJk9xdje1oaO1betKjzMn
sId8pt905NxKaUFnc4xFVH5PhTeWVKS67ljnbakauDwLxKXbe/9Bo+2b3mWlv04w
NvgElSomgonsxO0AXJOJlztuCDOjeY/COg024ANy5qGfOVupmdiktGiFJzyqwYL/
YWP/FzoUu/zeCf84Sq38ByjbpEtfrpKLiV5V2DqXCIg1+pQhKVOlKuBXqrzc8PRX
uxaprhj002PffaH3AjhdXWin+Hbpzrhw6iRmdXZfW4c7876gY8yVnZbLPb2S/76s
YQc67bCgXmS0W1uDb27iE4b180l7awQKz43PTm6wfgYy3Mzkb/f6/0zWxzRLPhsL
vb+vcwzUrSp9lek450w+1Fhs20hzZoxI8sVOHn1Qw+uV9IyvhPdL9ifS3Jgp4AcK
MlnDzXfI89aJXdiogEWBxWFuKEJtHU4iMEbvWW00eXQuB5imhMBbTXOem5n64FRp
taJpJWWWyFkMA8IDtmFwUQwyrAvi2ci8hyh7CJ2DemQWqmpDEv7+6zkcpxoh5U+L
Bg2xOMDC9YIDYV4wRyqLC4O6bvyd59dJWs+d9DBG75AurKyPmtq2ksoNZuaDIbZt
uBb7XE+HDqptTCl6L7T2PidIEr+7Ph21iU4Z/ZXoMBHc4bicfoPjqXXOf01O81zv
yr2Q1v5+uQG6OFV9oLaVT0mp8ll5Gp2ybGk29kVMe12GcwJXJIg0yX3l0M1bxYNr
u58Q9gFY0wbo7anDDLb2b3Q0YJD8iDWHlkNanm1offdygG2sCqunak1DkFTvinkW
RyjvVHvVtGrTMA3QjFyoQhl93D5ujvUu7v96hnCaC8FhExl1AHLDBJMIdnGfb5jl
Jn5gaefqqGyF2zd1zzI6N+9GveBYBTJrg0HWFfgSL801bl9Bb+XiLOf0D4fag+dt
SmHWuc/R1w9dwREFNLzu801z0pw/T7d1w90QbBxWL/1P4qXDRvdNARem22FurvGH
CAMD3GiIlqWOQsbv/NP61NOMQ5BlFB9WAson38zjfF6UZEkAMW/VJdnmD3s5dXiF
ktWUHrpO65YXqDVm2/VoA/sHwbxpvWAHnrre2w1EM9fIt+pJH59X+CU+Cpz6Fys2
qRblIyEp8p38BrikoZj6s1Q94qDxnoYTuQaAvnXpzV4NVQZUX+XN31gZ++j4rIQd
H/jGmiRb3ueEwhzw+eXnef6qPBoRCQWDMAN4XWDrOaYPHV2hjQRYN/7TvEknQrTi
kJOGaezOkhhrDFpDzF6hTAvYI6qmVX3udiarMLMerlQkIJ+dGyYJT7gShaikV2Iu
tLUYrlEE9LXgKc6tlXNugf3IEWheJFzV6jJoQ854TrDxkVpjeD8BntW4vN6VqCVo
upShoxij8T6vlCeJgsdyNKnW6JybeGJb7Gt+3ClA1ffBFWAEtye+hzpB7uWZCIWf
wvKs9YoVE6YPFWx1mpeuUqFq9xwqhVfKXfEPbQBHXOJuqazaJeID9ZB7J0lXuL1T
ShA+izMNoCvECGQwE9AowRQV9xwWVXE/LBJwcCzQVslMTEcswHtliq4M8DXh3A6p
0VJI+rWZXx9Gb0PP/OJnjGyHOOOxbiFnyxpBEDcVir4MrU5QLzLvXM/FDg1A1WQP
FAynAuF8xF1oMQPKc7jgA/sT0jin7GPGTbTAxACGPB2OvrDEZHJchE01bIx94Jok
7rJEFtgCjyM1vO/FC7anmUwPx0LHetMId+WPU5b2p5BJDCXHDyA9FwoxDxSBsw+M
tvyptJXlof9xElv89ZSKNfEXntRUpl9CRE38q3oP4X6ZOSCebcdV7CGnAhKPx/Go
X85rt9es/1wVEd/aaNFidrSRMgujTFGfI/YwX6FzVxM9Crwv+L54tglHRsTmNAuc
P9v1A0GjLf7GmKU/PPH8ELUUtHgAHCHEWpOhiDfRq4C6Od/PfrbttWSF9xJ1lLJy
AGhs4X0K/BqqY5c3rUC5LFJ/fesWTV785Au4KF6XbX+C4UwlNauZZIFJbKTXqQBx
0wELdD299XrL3Nz8uaDAlp+eD8xKtHokjYfwNMalNuMG210++KHh+vEitWdtdo8Y
L78U2NtH12lHTtEBZltiOlmvbYk0tP2xrSCaWESCa1DToHuZobNFzE4RXesKGXz7
AD8P8Ouf9FU+JFczQM1wt2Es8xNZGRcG+7MlnY74oik/ZrdEa8njh7vQKwlN8YcN
jhL29hPjCmOhmVkRDDE111SSLyYcYyIJ60/cebmfWHpUWVny1pVNebNcYG0QdikW
1viDxljgl6WQA0Q/OcfU/oPHtyF4eE46CrU93zFGF0ChhBfhC3CixCIuXw75N0d8
C1K5Q58fxLzrSmJp3L93wFpK05muXZkE946FKYQhmPj+W4t+cX0wdeuQXpYFpkA+
xagRt2diyuRUyqzHxxICKrFt4jbG5OZ4dSVmrGjy9sttWTSIIb8TNWuQaa/ve1/M
pgkjT1JqEvkNy/e8NYvviSXbdIvwIHytrBtFQjvoPC6F5E5qohtb7pH/M+iANmju
nwPzSBFOMatVs1utCNMypocxCeKWNxGYSbx8wupuHYBGbH1y8pcLoRNf56wkrhYV
U16UhgCsuL4fbv40zEe86f7n0+VAhK/983v5uyqcfn0tk71L3ZdXQy9ZiqURxb0t
34epTMSDaBvgOSjJPPx0MYOzXASj5HN3iPHiuP3VZICcwDKCeYMBlrgE32/IexX4
OF2bf1wfwgI+CpIY8ByAEXfI1aFQf+DgvSf8ZfjXcGEuDbDn1Vz+tYg7PfkOKvPn
IHxLOpmN28vePgkrlPRNQcYYTeiHXN+Gna0GM+0BuuKTKgZSWiM4sjb+XFRnXpc1
lPjtn6QCYMrnPF+lvV5wWdkLYEwmG0vQQLHEaDFS9ZoY+wwCJAgSvdDqXw/jQ1gn
BaWuTuofPDvBUvxBSmIbnovac0bwQJwino/mQ6qxlAhy8K1xee9TNS3ofEaqUjcm
0cRrncyzBknTNbMzSpttRCWt7qzisNDok++3Fdv9qyb8gkiYoPqr9ZsY8PA/DvMs
9lwRll+1qnjPiC1zTS1jgYvkYCiEB1XvKFkA9zOcJgZ4QGszBGMQcLW6HnJioIC3
Owp71hfiXb2XvUNdRJ8790L6oylGLEOQSbp9v+QDVUdEr51s/Ok20hhq022URis3
DM2Nw6sKk123pUVRZuIgLXiYvsxMFQyEuilNc1ndo6GpQaVsllNg2NxK/GBR3LuT
cdkqO9N9If+1AgsYHF8a4fK/UgsR6v1VPDSmIKFSvoeDsr8ZNpeWDTxauoJ6QXAh
UlycA/b+KSswVa+u/NiJYNIZr3shO2Vudi6j6wnpNC+27ZOLUDfV6ebWVAfOBCq/
Lbbi3xsgeNG3FP4WTFrsJDhm8Pm3LAyb7JhgVGgw06/U5ECBZ63uf0SKqZK7mx5G
rb1K+m2pNqattbIbD35Bisc16/n4LpTeaz3oAgmvVtn2RPxNPK3PuY432F1oYZjm
xrI9AscqInlzG8ZrlaNPiEtodQdRlpBx1LnL4NKujFJ2Amd02t5t3pbAEgem9s1+
2HdjAoyssT4iQXwcUpdDeVVexNvZmqsl0o/dbxExcVRMgpALUJzU6K4SZjO8pJ75
J2yeGl6Es2nZWmmmhKPznQoqDemRGzBd1BlUhEktaDEUXaRytLe/WkDCEndycvdJ
dwtRUPpo+rS0R3tuhivGbcY4eMcuCpjGwCCkJw7g8jvbTr0z0VBp1S0RxMj/2G4I
00gUcyLWlwu1GqmyZoPTC5GIyl/UV4rsXqDB3nrO9+Teubi1EGMzgK7+NN/T3rYe
exxo0SRdGepg5cpHaOX7qjHmc6cXYO3yAvRQlj9oaoOOlBvIfO8fndk33B0SaqoM
vsjkcqVog4TtBFnRd26U5wITla3vLFbhyVdhquKVR9zJ43HzeBxT1iJ0xdoNrJNO
YSrBKCg+HLAgTvJlYHsTabsrnq5nEux6VVu4ICZXtFHWoqDsebLVTRfLPF0U6i04
9fbxsk1Q9Wk9JgXLnfaOQIQP/eAVOW8hO6NycCe/y+JuaLWV9E5d2dnQLe+jVzGN
34BxSrMhymq91dbvqPqrs7UAwR5IjsE5c1qD8NBWvxDJj+oZwhaY+OVy4YxL9Cu8
1TPmIJUVhZGlaw45WE+morEWR1u6LaVEKTGxTq6k6OBz7rNRr9+S3ra16laavzFg
w4pUQbHO9Q+/45Bq3+8lE56jhwFnvBDL8VJtogSWFJ/oVBhKy8kgABPrtA0g61Zu
OVSPBf4xhLhmFGOkx8BmaP8q8IF3LK/Rby5eHp18vBQi+72wAJlkpjKm2AWXVexr
JI/TevhyUp4Ti4xbf4uQ26j4ZtaEVNO71j09neSLIBv9RE2k9dqRAziaZbOzR4+w
7CWdpfmO05yNDL/tOyMfuA+elMrBEEw8RHl04G0RZwQnF03FA0fwaC+ybUwxitwI
jQZ19WBDIDCzaiK0P6OcJO3Ah6MME9AMYiwyffQ3f4/4/4JSvWTWgZwfoxR1yQws
XCAdOQ/4f6LymkD2I8rdUafudiFqUNUlmAtYEo+7GSMVPS8x4IlN0xuAEY0XPxm8
TAMBV0+mZy/K/xGTfrpRNF1NIlsZiTWuLQr3FNPykTpV4dzr1UqPvgFsii3HIpgy
zClZNIDqAgsdYQsxqycN6J9/nvqnLlW4gH7rxz+SN5oVSkhtFhcMVYg6zgCVxRz7
t4ybc+N4qUzB7WgQnSo8OhgMXdKl7RjFaoLI88XKxT/YDjCrJbsfkzok4+QvDHKE
8pFnnt0uH+o97Pq/DYhv/R9P2NaQoM/StseBlXxfn/cye+Zz5rr+tB1XkQObqLmc
D3eQiYJ4TygJgD+c6iwz8rE/KuD3R0eI9MKnspC3cFa5Z9FyfOve+Xv+hbiJlUs1
tf5d/tWc1kGO50IO83bqvSaJlvbfoK6mwX3mkR0WNmXjBdPLJ6HCECVIk6Yv/N6+
Ywbxs5nRSVqtlqUkg7YGrN/u0LeLb7UvcuN77h21bweGv7x6EDcHei++Ej1NI/8b
ircd7uFoKJYP2LN7UE83alkOVzC7k2Lseui+HDnlWkv+XeB5aLBWTkMdzSuNsbOb
3yFWAj3wwSgYE9DZoLceyDqLfO5ySU1j7zevqDz4IWdK2997S7A15GfQPGzKiLCh
vUjfB+D8CBlqHlyj4/BycwQUaI7v7FGHTcmKyT2EH2e8CcJ4tri9GJl6MPW2nBxM
QMtbSzIIdbTQ4hxEYZ4h2mFoV9Rr69ssq+/fVXIzTvW06PdRmHQV2J04sV0LNW7/
7iYPcNu/1NcYaNyofB/rEa1gVjezXI/Cz9IpWF3n2N9cEfCUUV3WquNtg+/Tkq/u
ABYbkcfZWzk/BCGEW66JxDKLyITsLqouDXr41WM78ZkD82VPRd+9OxkC0q5wwogg
lSmAP38cY9QpKJS0UuyD9N2OxMYWD/54MlKqZK0M0kQFl08utr1tT6VLQ4fHyrYK
fiSnTMWsZTZVZBPi1AwZw4Ge6OvIueEQjQ3Nr2BrakFJ7iDwG0x0CDypYnFBp+44
ruNo20a/UeRz2Xs4jVjpRri4Ymj2K6BAkQGYQs3EA6aZFu7vCQllrqcgdB9NNKlM
nIpD5VfIdek3cTZ5eIN/Ly1+gsEGHrtjeByxtqGEED4P+dFGi79MlRDmvZtQ1l9B
Bui8qJa4iotGNmcPrXA/C3iilriE2WZtfTJEyPNl7u+gsal81sFaazhICZjxtwZA
VCjkkFA0TMshKu3pIcmInY6we24ILarTSdnjSq74tjv/geqBbkAlDktWqGXVo9Hh
SeUr7ykaxxja7WW9Q7gnQ/o1lpzZ/YJijOMHmwz3HoxwPppYBEZu5S27a4OAUkgP
WombdB+O2QBLl1zwxB1Ur0n5zlvZ5o7B85Uj5iuJCeczVIekfdbMIJB5RZ7JvYpz
ceFYf3t2K5DaTHhXEB/Dvk0tQuc4D3zDMHAXscPFYbZX69qsgpvXPy8KuQw+EFfG
kwHCikLHHqLycQcWmiREjUcdyWl685GaHCigVz+7QfAc/YTErYYVlD0k5BfH1Fm0
sfwb3vd+aszD2d6iYEQGDm86gq91o7vEBpZ+mewv0OI26fSJBfRqIowlua46EQIC
HvZtWhAtF1kamf3hWhf0g6VNcAuhD8wbvgKak06RP9y1WaqtOXAqLsg+JKL+qDle
kPIeRs4rGtjc+3hNS4WAPXm9DHRtznoNNR/pqR7yKqZetr6iMAH58c8/dtk/sEzz
/1fm8ocC0T5WV3tPFkOW4qUpD///+qI17fQIabGXA+2/7uDcbNNyzfB9uVtIVDKi
NotaSVEoNjAd1gVDBYv3KmVAYegooPiuwg9zTfxRwg1zQ7FBzwmXfsYTJeLV1gmV
OxS+V+CNieuwZBIpA4M4fdTWw1cHed+FJe0g/CoRiDfZYWFItSwdEySqeKDeLaDw
C6LoWENHpdsqglzrTo2cB4Vlhod8kQJdtal12i0axas5/l3xi87MWfPNx5jkyJ9N
EjT2i0N+KgsG32Upy5/ILCy2BL8FQGSXD8oShPRIZUzT7lWfCN+b3F4x0qDeMzH9
AbiRKy5VqPs/QOWR0Huadl29i91cC77JLB79UBJhODiXX8zrkJDiLRBJwDbQld2d
eu+0MbLOSD+BIItWQpLFcI6jWEOzTpa/MhLSyPaSw0VZpahPNGgCWwl3sjWF3Fq6
m+A7BsJfZXNd2B+43b9FpOBV3LzGjBvnn9gQq1Y9gdTOJbe41mSL8vnQQ9KLmCmB
pEJTrO+B5EaQnkTk5hjoio5cWhCdZQyEgIRrhO7DcBo5/vBrydvJOdctIkQWhgfQ
UEHcTSyw9hq9ZTXJcTyryhSc20Yl+H6F815UN55MK9rpTXx09myVqG5sPn1Qnlw3
iP8Vt6nOzN0uXwM6DhHb6WOLB6aer2ofpS/B9YDdAKjzfXAPyfQf1r4elBwiy/GS
AFQdIKGlIjBfvn9PD1q/GnLUCfYukYyzE6sBGscQ0Owf/Wga6tSIckcxtFEXL1Tp
7RzdXjGJtQi1FMgRYObPmcDmbNv/DR9ZcOAEZ5Sts7TR2LxX/fc2QsFC2aHGQSxW
R3XAuRPDUz2hb7i5kFYRRP36ChiMAXoli6YpB+16Pe6JfBVwx+6CTc8X198K26oU
ULCd38HW5ViZUWbvvnYZUR0cHjU9Kk/ej6YC8iV+nxkaqYM2PzXoabub/UPFD4DH
HVTLXyTAGDzBEidWazh+DrcAyXbB4aAJG5h6PX2MHICWluyhp0KAj4pbmazCFZGH
gglHtStFgFjcVHubAnBPmuFs+aTwnJHhBxNy+FArOfWvFjiRoMyxoJZ8iIv6tP8m
/y36tJB4CCvY0jM0isl0frbpMfcHb0OklLRMyeLHIl3Hlg6mdPXpSJ9bYqdZwub2
6h7DsO6ssPD5DwZuwWT7eTZeZewiSrauH9JaOm+yM5dqGJim9LIiBYGXsUjRFjC6
Reeq5we9M3GFt7TustQ9UgakcB3uynFTzxx0bTcY7s1N3omSFATs25Hlu7AHv+tl
NeOpuALg0g5graqUU1BNTmikT9FNh73nZBRWvD6B8ZbjXJ3e0dzvVaCq5DlJAsoh
wUlFPpY/998q1lvjv3TYyVruQW29qKhCyQBdEVPIuKmiXimfVjWX3KkUcvvSR1W+
PujbqESVU/Bv1QonUaXOiOtKcVTRHkGMQf4EK7o9BRnxCmYs4WA1BuZacxgfdtPW
T6AlS+IB9khL4CghixV1XgE0/rVVgU0GFoHm9UivXlTDE8o51svJo3xsrzs49B1e
VrqxzzZQdBwBiSrEr40dxJa6Urd2fC7LC3oigpWGQe07MW9A1LGO392HlM3uvIHr
AIziNbyFpMzqMk0P3WzJRm4YcqHYAW/PbWXhAQVP9BIwiH+TgL8W9PqBPgy1YaUO
b1viNN7ppv/hHT6KZxsO67MpJmWI3oBG50oxe+1wpdx/+mEfDxIabGHggFiC4gXs
yv1+b2mN9+4TodvkIrLwGxmCg+WG2wkpu0PlqG3jFO2634L78NL+PH0lcolf6LeX
YdN7aBYPHXskQUc5RzXElT9rD6oUnmsN4WOdIQWvnj65qIf7dOawHyJyjoVMzAg/
K/V/H0WUhBf/NTrUAncsww/hfroxIlRy9Mb3QFlqMdIZ+9eE1fSVnzCIVRIeib29
6pbX991D3lqvIcQXQu997I0xTigqVf3Mfa9yRIDWFgId+h6nCqdjN9TQCq8Zx+nr
J0nN4rIkZnqyZzL5B3r+1+duue9AEIKT+/X6nVN8fyHOGcvDQq0yvatnPRUCQl5L
NVXWeQ77KrTOdVPGvfHMOUQSaRk5cA0uXQ5h0lDVXCGa6nFg6VrLhxsuDQoY79O4
mRYUAIxZ/J/AZ2txF8tRzqddqK/fJ/2y3MDLQ0WAvaHyhmo/NgEfaP/GLROUKUoj
cukZTmvp3Z05tJoelot5eh9Gf35VvV0rEvSod0BnViD3u8dpv0TmddzujU8SCRIV
MjKFdktDdeZvm4jBK3fCTHeDGs0RDG29ZzoZ9JPqQ54guI/SyuSN77WIs69vZp+H
6V/0qHrAtecVBdBhihRyXoP/6Vu+M2m3s/ikAfqgbOYZbPvTp60mBl/iEOvMTwLj
3yZWeWVM1ajLkA69T4E4Sq95lasKCktdRNIUBydDZkR7zceFahlA9eMsh8pq9P73
hP97LY3uSuMQc8i1vZOIDzFyyS2k4koOdSNmWU9h9x9ShuvEIMqnlV7DMSDpmmK3
q2VAXJ/D/Pzi5UtPYCxy4MTwi7XrcKysFoVbvS0diPAQ38aBuQGC5m9ccigPj3fZ
g6z4htMnk1k1Mael50+T7g0NB9I9ImKhOxcz9iTk3cUThtpU0l9cpx+CuxLWLHxd
UpeoN3bdXLPwDbFLeLYgD825cgSiEnAqw7Pu3qeJLqfusjonRZAPi1Q/x2LSNsWi
RvnrtdhPAB/7Y25/tJSXCgs7i/hKtlQP3055+X9H2qwUmob/rHrqk8Rm1f7dfpcc
joSB/BSae6uTiWje94Lvm9l5AgCM70HUaLXuy2p/mZlzRwLN1EXtHPrf8WUCN9QV
bPqF5HxCwuIZcM9b8EWrhjzArCk79oNtrqPQ+7/76hJwYwzNYbVxTFyqQIVcFLDW
ZLLvdTFkfpIQ7aARocMpofmHn3g+qxYfpUEavOAStPHS3UGJ85UdzGo0JUvLlbOi
Actlupdl5uf/0MzZTmZUD2uKaAyQfg/aegdCCvs4vhoae9joz7HFykbW/JL2LL/b
K/a6vOrwt5jrgv3tA61PP61IKff7vW2X5HPrh+ak3ZHJ6zf64JYXSrrpZqDhi7i4
hsK0IQj3i9OKEnn4z7hH9nS4Z0tidIIjdtrFkTWAlqnPPKyyCbelQJ9fllBUAIJX
NBveKUMXcAd9b2dYfeYuyOK2NstTq1KaukOFtqxJjiFBrGdvgnY3tXwHOdVLgrXu
B1etJeQFvkqAbAmIV0WpbvoDu0PHYMw2KBFtUna59lrpcR1eg3i3DcoL7TZn91Ab
mWY395J7EYXCbO2pzNO/u6T8VpMqrCG/E5gPMfQ1MP/we3u9684xhSfDxE2df4U6
v15lyXZxYCwD8yURrtPAri6pOOy5KvLiMzZHk69qOO7ifzFeXtTVYPJc8OEvdci2
ZLawoZR1w23qStiTK1iIkw94nbySVGAi3kPKspnjPJzFd+xrpteP0C1Gpy+soEzz
bWqhSMztBSTouOZwYTyy9rwrEiQxq8bPdu72IOT49NMERZRu4sUzxrIz2ygnoXUF
TrxHrWIOUfXeoMu+HpkaO96asRmGSUOsDd3Ll/rZ0T8yxhFk/cNAaE80Jk5EYqFJ
Fw7F/wGieYywyEHtrlU1knsFweb3s6Nc+H1OKt2lSs8WS+/iBrulvknFIz+aXJBi
A6Eve86BLu50MjxhqNe33n+MVlN97+nuZRnMPVhi3xd5z7E2iDW3XlVRewDKFGMg
3LgMAWPLzx4tyEJMZR6TrypHX6mrfwPj7n5aEm0tcVM7++l/3L21nrtyfwHk9iNg
6ZWJ727HmOvbsZ8jmJ0wNWpA8De/hVgoEGiGd5nyrzU83mVUWYe1TySAgg5814a4
PGZGcNTK8ULPRr30nuNPC2Xd9h0yvgfmPYNIxEeRFiNJzaLVd9tBbkybY/YYEPAB
hvexRYdA6G3kfTBZ7oWBxObi4yiMKtNafJWVq2pNYgaPDigRuuNb1MZyNps1928R
ILCMVnOxQqJLAcRgLXSxTNwHyQjrXc9MU4vBlbvN1lsrevDj5CUurVJvBA33M6yw
kIe6WAdQ0Bicg+yNaYrF0gaDQIidtoOcUh6WRoPPZVXYDqdDEuJZLS+/AzZISkGx
gep4urDhQYq1rRSaGQgPc5uyoxxPU5J0wOsEDTjNRlxDGurRGXb439e2+I+E+lyh
+9RFQx25HTdHekFe5jKcd1f8qdeNjKy5s3NkFJWtPu3qNcc5T2q0rhk3UYA49r5f
SjUb1gXE62BG3ecXjpEP8rXZQ0o1xIsW3X1TNioZMrteaf4knaEK+7YrtyoPRJlD
t0y6yWkXbnlgmvkFEWSZLDhFEzf8h3QD5zo1+iI+y64lFX7kdOFmliMaJYDzb3x0
iJY6qaXgXK40fuyx8yg7FiRE5AAzHAnt8F+I5JI4QMMyH9jSn/zjJNZWq9ZqJnna
OBC3o+iIov9FazHnMSlUKhC0DwSNk8wizqHg+jvEnUCFJcOJmsMNEYpYR9QTnYU0
LJ4uE1KbcgWbTnKDQjDK7fmsFkELAlCWZ0zziLnhOQjw9pL8amE4t/juKUPU+8p9
kJSe6P6c2VX7F2W1suO5viTeGTsFAplistuIu9pP1s+mXIG2P22uJlpM06Mvi38a
oq0nHDZgI6CJMj232wmWFX+QvqGhYmBXNolYOMkuvfBSHlGEPLCHvFZn4LipeZgr
3MMUwYJsAK75vYGp/og4cWWNWf8c/ll1DtIUXjVMTsx/rtf5qZHMCAi3Nlsxmzyy
CBiiHGCyj+dTb6xvldwBfT2BTsAQaodvykvZHYrgfuM0OXvu0fkUBzQawo6IhDP6
G1Itx4BiomMK+mIqcnmOKLKQdBZ8LZYH9IbWAcRFyH2lND5WjYL1DGPZokdN54Ra
5nj4Grs+DKNnsYyS+YOm9XJJLTRjZwK/ALkcPCKThfN2nbggShOppi+75QN7+ffM
o7ZjboiOAIxrHr8hfE9n6EMdTBY2pz6yDNM2VY1fgOvD4TzbucSChrtNFr7JsstX
rKLC5VC2k5g1KwFeyaYRxEf2O3AzRO7DG/1bLDd0r/GdRxbWGlHFmPRbQj4pmpHk
SLb4GW+tj/s6Z7uTMLYU8spBDeW5tPJrHNuQfm0k8QP+WNjOGjBGTeTD/cqN4oCg
jU//xsOie1QLGVNTzIXhcrxY7B989ZO53WEu3IZIPWvgcw4gJdMmL6MZzYmHRvOO
L7RxfXBmoZLAB6s1fhb/ukQG06LYokVGjTK6/WBq+DSP6Q4INQmfSHtb1u8FtnfY
KrhoxAPIgClmVCTU72nepV+ry2GjKNwd/6pdUitTPvTL8Ell0ERmj9Ioz19CBFfw
Own7oqcIr6avZpj42tTPMgWdz3slX39YTzjJAfoTNzrAdFnhJX1loHAUBb1SVteW
Sy7DdPPzjTjdTaLb2zur9JEyEZqK2rvkyHxWpfVSVg0uGT4os4ptzWePDACmMU7O
ktxiCtD6e5CUL/YoeVsmf91e1SndTDZ/wKvoqAMPyJY2gQ8r8QrYE/y2d+Z0HGIw
4yh1ZZSYHUYE304uVJ3st63PDMnnJpU/pAcWd9tcxcaiZKMpejZg5IDRMWq4b3gf
ZTpRG8vZN2SlizKNcABJ7UvqU6BGIYPToZvfJc0vzw9tkVafnppJFUmfijrpB9sK
x+PTCcA6gDfMLl0HBE9tfX7dC3sgvuZ5FAaY6ew8wbUhlBxoNEVvIfNgGIole30E
hCtvZzjo3KEcHWrF8RSe7ZMRIOBd0OKMLfCyCqjL6pgNbfqBeZjRoVB3cZSFoeQU
TZkMzOHz5CiyuIuYmfrVZ/eCzke0Wx4B+56NvQfN+46HGERbCzTP33ACsnljUDkT
wFaIVgBI1TF8l3U5RUXo19OZoT5YCq3/h2D3CtYbe0YTUBt3BAIWRJSL+n0MXJQg
w4BcfcwMCX5cNTcrWiRC4fPOME6iAkvRMqm5sVQJXA10o1efxqulDxUin4D57NWY
9kwhZDf8pWlABzDeAEbBJAHNk/ho7dsj7NTSRvR/dlxnGJQ+aTIHxvbirCfEO/wH
GOrZv4Hg5jR2OaduUNi+VP2PWXolR+nSM7Bkapa751wduFX/JF8dpF8Qnm8d4E5/
F+N3aWCzVmfbn2GOcZu/XSUqn4Dc1nuxBVfl/+Ml3SL3oN6rQ0pY80cLi2Pty5ld
pg03B+lUvXJbrYWW655o7an4rp9/oMSYpC7RLWXJarvzntj+iAp+tZlxeDDUlEr9
021tO2z8fTYaGJedvZjqYuwNML+Lm3PiIknNyGEVewnO4nT36IgxYbtMSazh+2pp
z3BC8xubxXPFVCTQcIplKxMmdbaft6lckWZWt0MoJ4gJXJaPnu1Jfez4sS+US6aq
E+qzdqgv/f+mQJkgd7skS2NCWd0M5uztrZMfegf46j/JcdfU378xoj9BCded5RXm
rDk/JGebLM6KUAfnhn/iUI6YKbrWuaSqqR8zcHpgA2NbUz03UNS2tTR9dCtgAHs4
1Mqi23BebYP9bhOLyqlF/2TtrGt9xrLqM8vPD2HuCrN7IORknJhdlDg0QNOaRPs7
BszCY/raIjZgzqBPJRlxwJoTsrsL4oMkdoVHugZlr7CU99FyjBzMU3wb5liNrmCw
liYmqQzKVLuJ9HJleG2/Oc9vurHrDbP5KpqDortaUs32LHGSYvQgnHDb6STqT8bF
DpOfeTOwndoeyn+XjdWvV3nrqj0nLYFez+Z39dNlAf8rKhdTPAYh0AEnCzRUn/4C
nwhLRvmOkpXvIf9GMTi9kULv/B3wyTFer6HyUXU2qmAetEso+8xbWpJSgMAon3ok
QPSVFVjrJDa2auiZ6dTB8YJF+sAJRdkY8ykSqJsj8P9fs/AmV49pwSScr4vQI+Xw
bQ+v4kpt4wHHoAwh6cnm4+jNiWLrJiGJha+sDPQhXrXGsCmgGmXGW7++HddAr3zb
UUI7Lj9sXmSAnh9pQULQb/SBerk/Kd+fR8N2SJW3Hn/z8YRonHvmhEBzjJdI5J8c
rcgdYQx5JqeySORMTpUfauTrKQMcVeJOxh1HC0S85jT5KuahQNqTEusx2LxWt828
AsvuYW4B1/yWoCHdXhw3m5go3WpPDgPZV4fv9WCGmq0glA0dV+0KVxhM+KhiTTIu
bcG9eO+MeKl205kbUhf+t5YwwUOmy2V8kw8ldx2RuaMraJfuLRqgXwqDnOO1Z9go
B0PMcLA1rsb5IUKp5Y25IZFE3oiB/0qZl2QTKgcyxQ8ywIoBr6f6Lwesdgp2Hzkc
zWleRnWWgpGmzZ9GvSpjE9l12KGIzJhgi4Oer5Jjl7qW12+dGiCeag+kfUKOFLPZ
ZIppwwRs8mAUqearMuW7Cw2wlwMHZbbxObajlRhiUoydJmDd4LvySPGS3XsEGNsI
DSCbu+Q3bc9EvN39mnAS1eFiCN36CctuQ/jph6jPj9VmeqS1qbHGmIQ3e//bvKqw
NZk76V67eCkC+iDB3zzFKA/S48FaSnUaDj5vfExhE/gtwatZT8hELSY62Nm2LW1h
QdoKs6yx/zGxSoJ63LBftx4vyLnPGfV+skGj+txFrIXbIl+lTpwkF7rrXGaEqZxo
4lVGBCwE4kKXURUTQHovAGjm0lmIWS97Kqxs7CCiu4yA9V8rbRawUXiqgZR1Yx1X
P06ctPBEHJhL81FW/iI/alsqmnEZfrIhsiFebHWr9oI0jQhOQdY7BvOMzqvKRcWu
g7jOwyLLqEyfT7fnufbFYRAwMIPn6E8fYc4LsN9XulobWLRe+ydroeQFRa+ugB2K
eWNxKumPsedjtKFtE4pV1zFZvLIzSPHNosUQS8W6vUxZUqBY+JkpAHzxMsjb73+F
4hse1VAMb2tJyG8OMKr+OZ4hJmPsLkWuKWhkllRWOUawEPZqfgEGGg4TSEirwRVp
6ryxaJRIm1VIQlbexlv3Clg3Y7b9agD8cuJcOx+lLDK1wPNFZ4Zj1RlVW2uZbkA5
iZABsgvNkElH8TK3H44eeg3KWIMIWMVUSeutKUXKL8FVjBLvSZBg83AH6fWusocU
wHTlea9OQu+8aWoWD2SqA7KJyJBbv3/qtvO3gkk6iFzLXXmcGkhv9BGJfSfZ57+G
jdV95jtUbPFwWUbOPlqHQE+mlwHCNV1ZEhuG4l3P1NnNjuBbHRShKkxWQD5+EW4y
kJ5gfeOWNf7pj8/by//tSGmlRjaogs85gZuAiT7glKGfGQEUyxNBjENQuy2of8R/
Kr1rOmaMn/5VuGCjGya2iZEyqsYcttal2eLzAq4ppGrDCdB7E+pJNc/fx1e1rKvf
zBpfbFKNswn++aAX+Y5n0qh/HyloQ5oB2rsgNtwvXRO/XrWLm+B/zdAr1U8xYFxU
xOsUJGCtg9E9Z9wvVnm5RkqlfEbETsOlxn7GxOhImxzcYUoTIWX2RRxnzV2dFSli
opzq9CS84cW0l5DsBHK5f3Gder4ixgqwfeezE8T+8xhaZYkqq50fhGULxyihOo0M
8ocOKNYqMNH5bMVMuSsmaoyi8MMywLHdah+nAZfn9+eSCTKpf5rjM9d/80PzyzNt
flh/BRUtcvbZZ6vzHdg4eDZpM+W4heocsI7piL7mXNnspnFlO/Z/sxP+rYFV6Vri
w2zYGmswRDQmzWtCVoGrN6QPhSGH8zCYqJJsUsrBdVHoY9Uznjlm/0CwMJHLZMfD
4EVKQE9plW8VUHx/K0MmKCyTfCZSFT9M/SnJiP4TaqZEtBXkatY0R+jHegZ1Fybq
Mwqe8Ep0z2AYJLBZdQNcThStlbyR9R2HjT9G0bCCBenHo43LAkWLCzvwVIWTFzKs
F6Us+ZHWN3C1lS3HYu/Q7l0IKL+VMC+z0KvhyVO7L3MJl24eaPTDRus4LxCn74o4
kfL5PtNXk/gs/ufsyJgAKrBLfC4sxa6xmQD5y9xMIYmP+BEsAgDvGNdV1VD9h0Bh
uptAu3n0LSyuVp86D3+VCWmSYrJ8878Ymw6Ci9wabFAm4my8wcqh0udenyisllLT
dYTEFfZp8jR/3U8Im/CV3qud0uwc8HSBL9+qBYAR3B5nDqkr9SIi6Uei2R+7I1nn
O6XNLFkObHwYlGZGJQW6yuVNCqEvsfPeg4DUKQ920yqrHybNEIVzw2WLi/y2T9Jm
QSUsIeOth+5XxKe+Ag4RqkMs782Ky279vzRIUJ0WNiBwcrE8k6IMe+scjjpLQzCQ
L7L16oVAlwrp+5ZnXvhy8UkJxHGDckuvwbVLnh+n1yR3FYKmfwnQCcA4b9yU6hob
18dEv/45VbFlse7lkqfD2G9tYw34E0riEVnFohDr5tJ3Xp91QkjNxZf4RTziN7KM
tRzFwNLHSNapmJg1yv1SD3TDdp/ZtXvRIw0AA3z0UrFdFqQ0tYMt4QiY5BhGavbR
wKKxjI3tI35QUPROXm83dBYzfd9+CccAQsELvMgflsx2OSKBeVQvoNCXMPSy+pKr
PcMMlzJweMGy0wsG7P+uDedDy7OxoOmpojMD+mqpma+RdylqTTdReYhrH8jEgXBW
EpOn8U3Oq6+gxAqDAmxrsBcj7rlNt/lq4O03b/HldCQp72nzEdVB6FCANLgIl7SV
qITHbcUkCCew8Y9ece1GSTOLV/9SdtMPXa63b9wuweqQFJK+vSoU2A4ytMchVTwg
Kf1qmyWh6nN9L1I6arQvEVT1Jtlu7s7uLgUnSnDiUfGK31CrAuj87Nb7gX6YAetY
XOyczI2O0fPGFi74lsqKCkBZUojn3vsaq9Qv0dy/BV7TMuBo4nfRPoMI18+vC8vD
HUvxlfRooF+12JMO5DFtvujiIQHiTVQarCQOP2ApeJvWg9ocTHZeXEKQmC1b5VmO
gD/qoHn/su2je0S7mPkNxKMkkAu5ZJGa00V/gpHcgQDBxwNAog9uKw183bU5Ibzg
P7jO6MFegs2P+LX6raYaU/JyKzJ5kr9P+4RoovA6Tt6SLozZH0tPsXC2BXuqHxNz
DdjRJ+Lmb/bWGYBvFq3HdQGygt9j1nYykDc05w+cGYkrNfFFimHVNojw6akTM++F
OyAqfgzxsZ2Lcq6ZYumqLGPLiJ8WgO431GVzD29fTSDrfHvtd856agOcxM5w7GgP
+1HiEe5RLNY/uxHtz/spmuMOKtPMDZMF1p0GuJQe1YSFw6I8Hx1j9GxJfU76mO4i
AgX1/69LbHlXhjLjSBj9bbBejdcPX9c+8lisIYg/sRPArvsmA6Y/ENIrVwWOvfhR
72ef36k2WCvtOZM1Z2fBQf1sZjMpkwrjEttd1DnrCYSAuy0J15szc9QfSlpsT+5r
saVcLCtn5muPfDpFTbk/YRu0KMbjWBtakJmJWwTa/7EO6vmerebbh5qkTavleWJX
FbqY3MGWgTKFT5mBD+UhjCFD+LY5CLeW6x+h+lbFo2llvkUfCJBVzAci5+oyZea9
ah2z6NXHRAF5712vQJo2LMyQqQiZdZhORVHiRAsGddGQ/4NUcHHBEKO9qd1opCnz
WmVWe81lJURv80otCnuwZEvSw40+UJHyAsqf3qlAN1cC8PVDIxCkxLY0+3NjVyMD
BiPCpylypz3mqT8L55WJ4uwfh87ieq0ZTGAKzN3ASN4lIZYgbpoaJ3H0x4fDNB/3
Q9S13PbDsOQrvrq9/4aTw8g9ZZBm9u8hz9sxDRmKboCuvqcg2Yznhvwt5dvNz8vn
kd1DTk6CVudpD7Cze244UZKNaNsCV2P9wXqRu6MCTMFJDOrYnptW7njfD2MyLtLE
Nn1mMUMyi/ewfV3EpK6xAXM6oRgrCfDMHcXIUBleKs0WLXi2XMcbHo2Ry5qKhNyM
VgyYSBCHnJuDTy76MDRaCHItP99ILbYwZNN66Ijjq9n5R04ak2pfAfc1LPQGjkVi
4V79FH3eEm0tKsJ50rVOKpDSgIqu4R/IiOmT8wPvEuYfx/AY+XRGhIBmGKU49aDk
Xv9SkGPYNUjEKoDePktovzl4KarBJyctxSkGew1/sMOaovt/R2urTQBC02pgsvI+
u6jTs/5pEIt57h95XVNdFkyU2cVM+aYfBDpXXq2IQpWtiVQ3bXCgIL8o0JyLaLZ6
q+U77m39G7NMrXcWptkMykJigi9mGCsyzI+waRHOA9PXtw0T74TsUz12dnmQAUMR
bjp234FRUBsIDL61QskfiznjdR/MbYGftOGlrrETOP5qXew5vI9XziSo3aVtq0wt
PBHPDoMUMtzbeMP7I4KHGdhKp64A4j+JxuF3zOzH9G0B9iICAbgwXpIp+xW35V7z
IgSSvmeZCLRfL646rWhgVIBuAc3772rkb62515R3ZXRCFuWK+hKPosiMtxA28Odd
ba27mArF/iW0gAiqI9orRD9M9XguLcpy+rG4i2u0ejiUO/DTKqKlfjvHWIfNLvrC
nMsb5nd5/mXoGPoQuudeyti8I8Mc40mVp5GadGl6D7CRNrYi4p1bq19gsYxoT8XV
tzVppPox9P4KSOrLNJA9PZvo4dW0JrMc17QjW7eff3pXP57TSdPrSEJmRQdGl4nw
DGEX3IcUK1XS61sCiEGF1rbq88RrDg4Xm0MNEnAHNRlFPwCbCXm9I5DifrZuIibZ
/n4y15avA7DNhTt46iR1nC0f/uGh07NX/gZxhUryNNQDP616q9beY3Oc8A3oJGKA
RXJmtHly2WekotT8LF/1OusSEGNqgAl7GBC+P8mLWjTUypHhV0eS2sai8Er+N+nX
FC7N7QnneiPk5nDsk4bapLkOrcVHBJfi6O993zi2pk1kd/A8gsPDJ1m697u41O8X
078xQcu7wPt1PbAfcnUQv1Wzy6kKfnvvZG7AbAB1iHtS5izSzm7PRrIkfu4ZhFOU
muITy+hMp1F4NPECUWU7+V6CuTfgnSjCmoiC2oL4CMao72Dl4FWn6C3M7c3CrK3z
0xRfBv9DShtCLiGC0VJ1nXG2HcIsS2aNhO/wLqwT+42V979sltYcwUQpVh6UxOa4
0lLBD5J9U3TX80IxR46O4V9ZVXVpO8XHwG69T/P7ohYCdlZoUNEjtwOjAn7zy0yT
8VJoBiOtU1orpBIs/aXE77/DcT8h34nmv7Q7306BLiUPDiv45W1pwcWBCv1eXarb
LcLsILHNTlXfxex0xjFTrEMRvCYSFr95raP3ggvrZErAeLBN78d3Z1sJWg0KV3xO
KHYmuzyGlR6ljOjoP6ZGNMbCszp91UOAUGhSbcXuucljhzXESK74C/DMRDeqqOA8
QiKr0yjuzpnEjQy0u3isjaXxRvUXCmesb0Ekta70twvCeiQyU4wUpKH7MyM1zJQ3
UzQfr0iy/I7++JkiqpQtJW92ttmDuxKkwZ7IErayRcQntMFpjgzN8zb4LVgj4HvP
BCYIzzUKKDIPi8IbgmxjPhFtly8ujBYpNT6Sy/9aq7BwjVNgKGyDgs1aI1TmQnlF
IH8po2z6xehIZ/9EMErY0VLaQhRyCV1Mm3mqeCnlMjygSXmtKHfPsWLr255bxXZK
zCOymEYLxC4GYRxYcGR7X1nmEamCVTx5WWpE5jrknOGIzxS/SFIxdt28OGY4NqMs
c5HITbSI6PwUCuSz1ftIyxbXBcY3cGvFSd5QPG0+aPqDs84/JzG1YGXNIc1FiHCC
nm21VoLsCzNQkvljiiWabvTzuFv6p3McJpyadX5liDAk+dewVYaKkqKOnWRnVwLn
iZPCKXL5tOBK+F4mvgRpMWYQJARTeSPpwAdO6igJjwQDIR1tUq1LDDVJkqsB7b0n
I+52QAWAGflK7e+wULOKJHeg//4NxaCq3hOo0jvzQyTQOXHUP6na1xkGuCectbyq
JjCmI10/L9zUt1tB3g4Ehux3BMqQ2Sg/InIOSLtkDgFxh7/zRJj3xft16zXhmoDp
Kj5Pu8ZEn/L9z07rotAXD8EYIvpyEaM9EaXqokgLDDsAnmq1ki1nBzexTL35pIuv
+FgDUtpSaxUrAzKUdURm+OeccfNvv33LAmO3EbXbL+anPUoAMVMeUODQfKQiz4f1
KYH5nI9nDT0rWmS9Y/UQ8ruhSgBDOi/0BgSWjvDBcT6kaKqIHbap3QreEzf4j2Pu
fbqMqC9gwb1G9eqSD7NNT1T6xS5WyMmdSfXc+VEB6FSNCqiFFoUVp2LVR61dKAP6
aS3Kuyw7QRescD9JD1YxkhFG2ozBQvZq0I1pSKHfn3Cs9+7t5MjLFCJU8sc+f1WR
WphgIeHHqIgsagZKnxHCNmkkfIJrMMUdLBKwQnsBKQsVSW7JLTQA75bFhRsBr3uZ
4NeGBpvMinMl3byNYUgHWugk47je5HUp7HpEfM/IXUS7iCXdYVosL2+9ZeGVYNda
CdaRZ7F9fgRI8rFoQNJrVO1g4GHNrIlG2tS7h80NDU+NXvdgVwS1u8/McAXm16rU
6l6sOLnt2vVJTpDkkgbw9NTOWTOu1gFXWpLGJlp9cm9zCObd8ClITHvIwGL8+Pxy
YKSrqvqFATm6GT0JiGc3cFZi90KwBO7Gzgfrpg+jD6Z2g4TM8xkxmcD+s9E+9J+h
aQ/YTJCxAsu4QUknB12VfW3hNvzxsga4fu/5rcSTVLbhixvKuetjUkX+WynmqdOt
tS133WQbGj7jvKS7QMOLjaPm1V2/W3eXiybr/3ZLaJW5Cp6RUKP+T+hiyLQ/JbSu
ldOchCU/2zRl8L9cKGhf2sJQ4ZAnDLsSK6Ysizl8Suj05xKcpgnPR4gv1BpqQOv/
7TMFh8qVRkRaQMXotDUSfVPN7o4wtGmPZjE2CDHv/cKiVG/VeXt5zWi6gfLa97DC
4NyH/KWJZGUVyhjAjtHj2lsKoRXbaaydbsgSzK48sUwjR5/YVt4gbXqoU07XWy41
ydh+/5FwxgtgbpL6KpkI6/f9eiZcIhN5zln/pAx+Ef+4yr8YQ2tjtHJnXmBES1W7
NcfHMc+P95rWkP/W9xySCaOnfJwoRQ9IjJqi+gSF4XCiFvXlE+nLTc5UjiHKCCzG
mTnA7hAk5+r3R8gXx9i6+8FrXC9vn91iV8H5o4hg2hS5rnd0qMfW1lRghxh0zf3N
Ci17gDftjmssNymMKjAC8Ktv5JG91e8kNMapRfKYdXIWmfG0vuBxkwAjtKNPQFpj
fCSAC7ie8dIl+k79oISVxph38sBoJT/DFcLu8WFoQ8ALum+nQxKNz8sgQsC72Z1n
4tSH2r07ufzbpe2S7AdHqwSt6GRRfFgrj1dPheszdq3YzIIbjtf+wblKaMwUOemg
fDwhlshrlFR3iyHexmbcf90F/jn3sC7t+jKm5UMEJ1fr5yb85DxHrCyLB38hbcpU
mLybn+ejLczfBaUK/ZJK9VFBHutgJOfc5SvensAPflj5ObdrvSasHgXlQdhrMFTW
P4GQpKdobbIjqFqJdpHxXZ9ckArL735MnCLk5kZP8PggZwrSTIEH6gFyGgpSsQaO
L0t/M7rVYS+GMMTru5cdpQaenBT1Fcy2gwvinpCYpjH/GCyARySw6An/VakkKL+P
caLwSCnWXsc6BLsGA2G+x682oUEj5Eb14Uu+rQldAQW9YrAg42gCPQ0maXSvcxyo
azHwoIEHoZC+1klIHT8x7/Ruij/e/pGEjAGDO/Wv0c3G2ZA/4wJBCq+d6uKqItD+
fXFAgNTxKK5vbzJSZ0xcNNY0at366M/woDeTSzKwsWG35GH3B5EdyCUGlphTLybJ
W8/YKyHfmOZDdKGweSq0fWEuk+MWJZYFs9ttNKMkgVs1omag2N7aebZRWvzmYNl9
NGq0pkKes91g9OScc6RInJeZjfENsvwb8vR5lRqESEkOGSGVkwOMIWkjuwH+VWg4
rLpgC+OyWsxRW7H0KPailGw74ZSxTC2Y2TOO1DYjGo1Y3dKprYwa4KI6jvORQKaO
XXRBmUI+tq+S1X63DrarCvRT7jR+Pc1X72TL2P1F+NBt9L6s5XVDllp68lQmG5nj
wkjkj9SoBmjS8rOMVKo38KiM/LzFFN1azTabyvZSaWRhXbD89D4HoVtxmCIJChO7
3I2rVw9taC2HGm/M9X2+J3NUFv4yiIi3YMHlFL3wYhEWtrRrrWYhZKdefnhwVhDz
7x2v7TBfJ0/6DaCHfBbM3k7iwOjV328ZlROexkRPQiyoXQ2X5u7MHe0Hi6tLJDEU
1sneNj7Tp+flWhIrKVfPltNac0+D+nAyL1/U/kNfGZEBn34i0eFzrRUi6l1WVDQw
bLVsvyzH6yFkABvjs6SWaCagl8Tsz6j+hh10XP8mB9t+WYAENFWNgfvEMImTAhsq
AahEQJ9V1LEqL/mCSVPUjXggk/vy8r8wciTsbwgZNVVWxBnjRuucV215I499txGB
pi93q0ZHCuBW/lEWkB1R6Q6GqkupRwyRM2C4FJvljFrhczSTgDlCerh6tyRXUlnI
SmrJAody/7K0I7xKrb/BUZ3Qq1jfVFXIYewSTzuzo5aXglaR7wMVIecZ9oYAawxo
dNbFc0ciEjS7QgCdu7d8UC2qP6f4fYJH+mabrCPVWaBtg7ZWx5QSxZKfQLXjwZwn
Ru7bsKIZlTUnBXA8wkiDvKL6UteRUx4bDXx2FB7+gUCyBY99FSQTrtQYR4gHssOy
GiXS9kDolfhpkeesDK70C1iPnnFum0rT8mfocHdcMLSPdjDa8Y4/3lchFhDVMKzN
YOSOVl0cKq3DH178R9t2OykTWKGapspqAzBzAaOXTSY3dlgy/ahIagyHRaIlVels
/6Mg+OfCbseyMEu3OMnCrljJS79/+iQuAb6B+NhJp3r8nhMNTZ+LP8ssmDpGsQE/
SATdeDlCdwnn3nI5FW3kGdL4Fj6j8Kz/xJRFZAcOV2r947arqtFNB/ub06N85uOx
wyOVTNnnvB9f52KZEyiCC/GlXSQn0xlr+QKBMytQgTCyCK42dHvSQMVcygixZO9t
5MBWWaWKYHuXiDiq9Y10oYIKA7CBEXoQrcuyKzzQoivZgFT6dgOjqY1q4e33GUtN
EslnPC8cQEJgtuyb24rNIrr4DGxWmoRYsRDHeNgh/9yVHsJ0fAWXkznDw5tkJRB4
54tkteX1boVFHV0qJ1eY8eah+e8rZZ5sVOy4l3RfHMFEgITDcQjnzL3ddiY+d9Hr
8u8d2OSHP9gIWKeN0jZNvf7bGBG6nuYGgmqeRYElTEekBzGkTHIkT/xcEngVKho3
++rwF8qQ8owa9rc8FOhK8XsktPcn09nmiq/1kkEALPrvJBj70p7uKnBkVoBYyNah
Ej+l2g1HEVS58gTgQH9nFNPNmTEXSBCqKbVYV76degZBjGafqnWi272mlDrAQGnO
QtT2I4LBCZ/JE1L7LpnJ5bme/sPapf8Gw+QURWVPgVLDL705w6wqE4yZydZz1483
dsR8dTMW5ria92ouW8Is3+K56vJm0CKYX5jZoLcHgvH+j/k8i2xo3J4XRWDbxh+i
6EkgvW8apKIb94FHjtw+5egm+zzJsIAtLd5MH+BQsLKt+9A3or7N+AwC00i+Pfjj
DyMGUiw5gYUnYdFhcDKhRYGfo9syPKt8HsNAOdOSH/UKsrT1ofFduM7Agh0iPdJm
o+Epypld5ClC85iH36wz0y5Eqsc3iZBeuHX8Gy3Svn7nR47Doibgqa2xunSmmcOS
VEK3DMvV20t7Udlz6SX3PEQlC7mM8LHIZYMApKxnijXZS0syjYPzSbKSvb9MTlWI
Jg9RPi1o1Od7AK/Dwr5Cb3BjGG8ivEjAoXMOffugT6FPVVz2aH2D46KAtmcGcOvP
ghjBCoasGTD9sOKD+PNPauVa7v29p/1UI/y2o49lPuwp/hhS2/HtEt93IISpmjcM
O3y+5yHybs7QTHqei6siLvQsvbnewMu8520YYCkW7HVwfHhnqcCUZq5NUT51jF0H
20JvQ+vwpIUUX3krg/BNQ6aSwm/kECwycxUCjGxqh1Y74f3HmHW6GJPW9G8cqzD+
eUkl63jLGrubyrwx4c0asUgcmTm3I6TaESdYhf98MbBKveVaYP0FRC9KrVr0iEDl
7x4f0MPxwF2lGprqbSj9OdZv7P6KbIB5XLGzREnpA6jEM8rcJxIbiOHsLaQeXtfB
0z5ddqs+ACVTqhHmtWaPR6exsR0SFQSvj3dG6RtIDe1jSWgchP6PRCVpI4LLeamP
etPJ6bBmi8r+C0UtCnTIgT1Div6ik2SyrKiLSRQT359xEqfv5KDiS2V8jbORw7oU
5kQkFII5j0tzJ5QU+UUTak7dvqqV8urHr3QGgqoyEPJN0M8eK2e93Acx788N78jH
QGnuA9lVjXTwI8aZzL0zM0scY1FjmEaqxkFsFE+R5wywp2if6zd+JQJLZU07fWYv
dUAMezKhL9ez2Vw4HYVf+gRvSDqQSVia6OPWdmIbNik6xkHeFN30xZ9b1I0J7yZo
TN5pVn1jD+2gXOGf+lp+CRrJeHITLK5tSDD5sH55sCfwpi32VROUsBVLJzuDp5v4
gV6rSKBg4Id+8/Egc8Zk4m9rXKLFSTgI72QS0IdqokZ9Q3DwvQ7fPtnjn3VZVW+H
BooLSaG0wsoer3QHJRDFY6/8GS3URbMx3S+pI0mBSADH30LEOjSEE1G8afmQcbTF
L+nI00NHWTkwMsS3zN/4E49dxTyvHvPKQWKILnQFO8fOzaGuqsRVR5FQot22imi/
d7Ig5Qkpz9eOroyUW1TrYnu8jjLcGWrZrCuSYKnnJtM004O4E+/MhVSsP8AJwM/O
LnhjgYE+HhfAmSFnl0jRyicN0poragjvRiuwvgSDzqi5xdPQy7bkc5xlP+/HTAJf
Iv0yevLYy5DcBxu/dzDh+QIym66+v9gLloo/XaJTcBJB9LMw2blrLfBT/T07NcwJ
/JQHanxJImxke1EJqV8Ytkt7uiL97TnSuFpT/Xzmhyr+4AQA4qkNAvhweTw9+DTd
qHXtpNqpHsrX9qhH/S+BaA/4iuSn781uswzr6qAuhNzqMiMM8RmE1MfthtVxlcg4
GlvhIGgvC9VJA1dWT0w0khYnzqMlDYNYOCJXgNx0+LT3Z18f2BNKxfaK/ZJXdt1a
I8xZzr/M6pXfpqVu8PO0bd1odCyDizWBKXNsfzlZL6Y91GaX6RmmIpLHXSBAgqGp
SMOQc/HxPQwixVCLMnPO5kK8/6QkhbR6Gr71V6WEOSwi85g3sW0itq6pi54wC3ce
JrOp6UDYQT9O9CNhLHAp2o4OTjv7+J0hCvZySFVk+LGybKSrGdv1Ak+8yogdA+IU
dc3g5Xvh1jf+XDzsAy8pZ4NEmOG/3vGLgrtFLigBsgAb9VYQ+k/F5s23mWjKON8e
X51s+uaTI3LmIMXkuyajl+F6Ycf8zN1b+wBevla1xiMP+5SaaYvP+BBlmnVPGJp+
MpWw/4pk/xE5pEQdO+NoVgGoe7mprXX62VXwCLWmHO/yRM5y3vFLmUvdSmkG+dez
ir3ihse/0U08p4z42zhklVMQRawuIQZjgXgB3wbn9NqVTedm93cSC8XbM1eumk9R
1uw1r0RvRgD6wcb5K57XS4nO9fADha67l3Hqtix5ShpHPw0jytyUiuAYp4UMhVAM
aDbAJ0kCe3TgyrYyysTOOCiX38oXbOBsNxa1l8D2BTCFvBR3Ejjn7VK7bgekiraK
JEcQ8i3SMgDDhnCIBjI+N90x9z8sdwJ4Dmd6A54OGT72Tq0XTcPN+mN+CVNhTyyG
ADA4VALVXahLF7pIZgIXH/83i7lLZS4nwoHPFsfY1DMEb0sofknqCt2VjVMP9ps8
rZa2OnVq/sDSa+Wa0ahqCRSffNa1ucCo7MTO5j9v2TuE4AU+QOuKa2L9C3LLY5tS
rtYrCh4SzoFCFHpBQH+tqy6nup8WffOJowgzzYGWqHJU+8NLpOY+ytHojSF3U9Nm
bGyq7hyiD9HZyhIvh6DJJLjfTR8R4l3xldW6cCGIxf3ikI49OBKHdAcSTwzsk1Ft
DidcCLf2TwfZCjaGsLSQL62nOG3zl93hxVjbHU+uPnVT8SpwE3LT34HsgoQw0XVq
z1gBrf3T8frmfi0+yTz86qUqpW6xkfceREr3OTGoNtIv62dXMZj0u+z4it4W5Uph
JVfC445jVYEHP4jExX2hqOMj1Ld/S1PzxmnKPW69RCBHjVUNwOiOw8WdfMXgnnOZ
ymji1a3sVlwsdajBQy+FWGI/4ubrJqxn3pw+TFrIVKI3XcBkNCP9XHmUhlwD8EDU
wJktFX5H+04JQyqm4VwT1TEEYW3N3efE58H0M7IzkBqKFlvvNdnnim8DPFBEHF5+
Bj9VzgRmp9M0GYcs9zqjlZXarvXeu2Q80GO2foW9my8Yu9dG86PKs07XW5fir7OB
VuYcnSYuFwkk1rGMooEw41u0xW/RTOsjHTWr3z8a8KeccefG/c25QZGQAzkD93Q4
+yJrJUFPJnnUANmfposYaUJz3zZLXqXTCM68Hc8/WQzlQq3QJpWr035VMrCKq8gc
UHXzS9VhuGPnrAF2cOPwXv6n2UUswy9Q9uXtbOUx53SRPFiU/v1OWzd6sw8XGBdH
w/86K3ow48eTm2QnWhMdCgmBEHuNA5+NaUXL6hyDaiVFAQGH/6z87PeiptxI0J51
a/DhkUz8t/rmZD4xCGATb1EkUDo5t83f0M2/mfJhQbMM03tpDsvyGmUNdVtSTszo
+wcrlrrtASgE+/SlK2yRt/8Dth4+d2ZIuPOgVlp8t+r8KnWH31Y/zNp7NTwtQSDK
Z1fOcNU71FFvFWI1diZAJH6gzX7ki6SegDGX0qFKhMyWdKh6Cnw5Xo6l3n+mJFyo
EdEOLFZml0n+CAq+RKQz0TFY1dR+9ZIz8oOvjHC/HdLL0TPkBfN7GYtHLJCU+SZX
nE+W+b4jVqyZgyYWlZU6Fgp3PstegC7iOY/KOc9tn7w7yt8tGnRK10SuiAP8EacB
ahtDp+vHxwUXWLK/UcQEWfIqNivKSYH4QyjeeOCax+JRM7IGMtmphXOsqk7TvoKd
zkgXOWe1LECmrb3hFmOFP5rRwiir/fnj25VrYJhB72KsPWnlzg1AikfqMk8FhLtV
USOVcu95fHPY/9bUjg038SOMh5yzTpbO5UJ8o4slFn7TB2ZJEIuEL7laMfgIzLD7
K5BJxe2u3A1ArL8TWHMgm+fl2rEwIyafZ6mJvDUrt05sBVnKGVmOO9sR0D5X/ST7
1hHCRRh/cp3FiddcQx8GtzO9ru4/tNsxSn43NucKTYv0SDAxCLSSKtFgrIsWmueR
YVUjFBH8YZHJZqlXYUYoQifeSg5LMXF4nBe40HcioXHEIDxbEyybiPgTynr3T6Q+
6zevlu+za6zyCDEH7p751gFBVnneWzMZaebp6Lg5Dko7DAe4372xCm4MuE2kpjRD
2jlo029CLg8drzAm0a5rJ7O+i5Gf5qkx7KQ002/5wLYlKBbuuuXUk37Azb+2A7iw
uzSmUpa3KkMUJusdixtSdFbWY4c+FoRcHes0dLjHVV8DAY9q0zf3BjhCUg9d//DM
iclJqYAnfaJY+heSAh/GwsuI1AnE9tYsn8lvug97KNGvgM36L6IU/cmhIGIJBYQD
fCcctBByj76WC/Yk4ktU7jHEX6e8XY2nLbWT1e3F68i+pTw2eTmf+LC1HZbhkc1d
QChr+11mdUPYlvLQ33adyHI2g3xq64+fRAP9r5IjFpIU/UFtdA++JtaYkJZg2+t8
2zQN3J/xLD3vDamhGwzY7cHmUfzx4jPE4RR2JD/CJhmQkY5ybBGkTCq8JKw2NYWY
gNrmOXKGGJlhhkqxxioBpdmnQBVvtHRznpGgSxA9MIOLdnuTlLEQA0YNbFrnbmfg
+3ZzjBGXQ4drwGDhO5yagFdFUm+q6WsRM18hjYF7RvFLpddG4QiBdG7NsdJlqfA9
E2AKPPndeb+DflwIo4XmRBCYQUokByUWYNhlCYZzsI6Jyd+nCPYEIQU2q3sITdvC
I2qqKbgSIMHy572Dz6npHllUu8CNT5FAcvAy6F1mAfFc0BWYduuH9+AXtUUv0J9l
4Q7Rz1o2wRVNj0DsMN2vlzq6Cm/fHNWPpXyltIUEWbW/2n8SsUa4cCDrVyPC9jJF
BAFqIKdqDjDlQaP6qf0j19CRdERAs/kL/igQuy4tT48uwgADKo/bJ0i7VCCQw7hz
igr+Crqpt9I7SJi8t7z19HJ3hBDeqEtNZNzyUDEBDjxuqe3pHxbAoGvvk1lkIsHX
Rl5cFm5jvOi48ldWgrC7RAfUYEfoqglEmmucGyK+YmHg+7axKo1g604LKBaTobRv
A3X3EErJm1x1eoBwNiIDUPPgSkX1AW7d/O+v4lTvXUqOlbP00KCeJFozaCqlqK1d
uOkumxYUZQOqRK9wFNAn2cd37mdDxxITy4lAL1RTTwy7GGQTdruP7SxRJSor1Psj
75ATbJxgrmvPcG/F/aaF7pIy9JZlVvUlOfkH5x40ffhvddL4Y5PiSNs2Xm9wM+Y0
nTXzX5PoVpV5q5qh82SyFP/rcPS4VXdKGlqCDrQzm3q2E1Lhl71QOPHQ5E1DVMBZ
dFtZ1RYGgsTsKFK+hKRmeiedHmyhmb4WxUfkUepbT/1N4og1ypkCu77LGC93a9XK
de1qBdGgxpHodYEa3pJKdYcj9PZirEGqRJMf9cPsVOUnNW132WA40IIcRslilGZ2
mQr4rePFhPIT9O5UQLaf6A2eTKEYbsQAc/ZNx7Vq3wlH5IoXqDXMYyR5Lq+Kktk0
1LUoYEKGuR2B6bj+PgAQIg5wsVN8eSXMR4aWRPNDuafGC1ZOYu6+rPhQZHM1ndVh
cxO6Soiwx7PXghcYvquah+HmK+oimIR02JIej/EkPwdzm3WNI5uOgzzzPuQ54aQ4
hyp/KycISNyPNBvEmFwE3d91VOuvYfBqAXb/bdsP5f2D5xWcEV8NXUw4WA78e3YO
f7yILBvjbgK4GUvvkV97ocI/lydERspteBgRJg0XKibAydPHwuIH7YieCg+TvPuK
DYxEK0ExPtP9BeOgCWjbR3Wwf72d4REwM2Os01BxFwNr+v6nMu4ruqk0pU4Muffo
Q7v4AcNGyOE7UMmVEBWhcUrfLkDc7hGilPUPiazEFWuyD6tGLUAGDHXnRAvdAngl
XEpQDxQE1rL35vg6KZ1A5fXsy8ONP0HK0T0Zg3pHz/qeK9hdfOjnjzdNwNEQp2wh
vYoO+uYeahlqemrIs+UWluoJL+FxooJqGmFbTAUUhXFXPwBEy8tqsg4HcCydrYEB
2bb0cUFTyBH32kCjp+2H719mva8ZwYkCPUeJ1Gh3Z+pXSJU2tBB4ITvBWhu6DgyI
eCLHlDwHoFypAZwUSlJtktwrAXsSHe6pKdT1MYuzaYv3jUvb6xhcUDlaxikgFVVf
+Jp5oeURQ6c3U2jnVauKTBF4tDkJdYvh6iHNaxNwcXfJnNPDJvhLubHj8Y32zrKP
OWTjkNeE9+Lw4A3/c18BqbOc+GVJ4MFkc/xtCKP2aSsLuqodetq5/XtGvY8VWn7N
l3WnTzQchZ7KLEMR9tf3/V9D6cQiLI1Yen31S2yIr3uEv/Ps6mHE62rzEGoarykQ
LDv/jCq9fIVeObM7SgBLFG+p2PevMk6BC6+4QH+SXQcEdn8huW0nj9RoOrj6MmhE
EDEj6Pghu0WvTHdnegm2yuCF2U8tQG9NwINSiRd5czjDQg0sCnOFU4p5OitPdbVt
22IWNcwq0zpLMv3Si4CMMF5rmZLi0pxU7DztpoYacE4HF/Yk1USqHPmJXcITusT7
op3nM/naRvBchSSTlUEe7wXxlNx4+dqy+nMlUv5+I7rKEsqDW+EuVx/RLwxxd2qr
TAlWWdE4zPTomA3lf7U+tjJ+UFRVvkM7a8IZqSjcfVsw/fPMBLsfs4C11Bo+6nVx
CeplikRc0NjxRr8dYwA5aDwOZz2zvg9p8hItfMfKg0w7lcE/u1S7iyqxLXHzV7Kh
W336jiRxk01O4bJTYInFuVIP6U8hXxh7cQrAhUri8tkbjg8PZ+XL3RornVM5mKs5
w4y31zmNh+aqOrRg94n1hfztJV+hj6bDEDzcq8aCm9pLBmEBAbaFMGVJqjKBgLrG
08m7MCRXnxxAW3N5LOamy6EPo7jK81uObX8W9PkCz2L3WhD2G+bAmBIf7C7VTxkk
ZSeCX8PxCw2tOCCJvFkQF4Voibv9RKW7EtxGcQp7RpMskz+daSceiwWiHkrBbNnR
tDSyJRtgSqbxrserEyV3FyPq8dG28pAU52YTqKW4mPFM22NN+jEuxVRNncWHBHm6
xS3NBQOpUhZgeqS1OAsxX0fy4bonnz0f9A9hLjdZCki3Hf2A5mZ2cLddH+PAqu/K
Ds+R53GNabTM0kJP4wPrbNsWxaJdTYH0m7DjH6WlGGJz4ELwhGqbalMG/9ZNcHUs
rvb121Kprcsofyt36saVjAmv687eb83j+ES/R9uF7seQ0oO1dKeb43ftusQHgfm/
8MT0aust4hL6CJRi3yAQZba1Ib/+AD44R0z0V3SglQEL/rSb+hMivF+WGUb9Y7M4
aqY08hl9h+a0+yG2oo5SlRyco/tstKMVt+IF/Sx1K+3n2t5FD6AgJR73Kf4pU0uW
cFpt6NCzKOYAbYxv7rK+E364vs5NAjnklSA9HBhetG8sbnd+FuzK4bnarwvInurw
o4qxNIqKqRLLqkJnyFUPnLtiIg3evgts5O87NI1W83Q0hulY3shAdFBFOQm0AtDt
hNZmTT8roID9pHUyxxKz3xXNjfm4rVKrkNXHJPhv+MmwghDQMLAu6xYnshLVRdYi
e1pJ26uXVIsmgKKH5l83Eq/Cbl7Mybamr4WwJk2OeI8DGEJ915SGcCrn4hy0Wi44
s6EXTD7LBWv0DPKUH+T9oVtwjGaIzpziLujbpZfCudlsgf1p147HYOG8eHRAXU2P
gWAX2VSb+YV3qAiD4ZbtdHQp9VjH5lkP3TFMDESjiDR73bvLa1acM7cf4H8pJp73
IB3ERuAeo+YkVvyPXewpI4xGCPSu1+zrFemt7oAZydyo9G7BTLNYKvVOiuPUEFdt
gZTc1vh+hgv17gDtbyrgT60LIHm+7EDEDGozm4QfdgI7snT8V9Aq4ytRMQGjZigS
nGopS1gfzM8tHjuuOAh5nmAXriceaZjOgSPKgWfQhYJa6dMTxVE0Y2guIf2pqTBL
t+Z/9aKNE9NHWqnsPkVJDrPnF7L5/M/I4AP2CpB4ATDRgdEcDrIQ3aKjAzl6BGDq
brataqMtQpEhMyNAUg6X5tS5EFeXcq7nYzOblhlabPb+2swCok8UMuvb+cjFZGJE
Q7J08IhM62qxgdYolj5fg+D6JSYDyJ9j9w4aZKwCpKZp8QWb0ypIXWQf+H8Hdjy8
j2Lw01HlyAmyf6b1g99wOqX3tvmUku1LatpFfaxvPjrn0YfqeCOjGaHRGVWciLDC
k1AseMk4O6kfpuuvcuNDcaz+QYqt2oTIrRE/Qxigjf7WsSxAzi3eU5SV8R995qFD
BRStKont0KBTCIwjFSgyzCDeicEb9Aw1BuhPRjgnflqArzN425Z04qUUi06FMMi9
7xa7gtJEKBQPoK6LaWyZ57NK/jJjaHP0jnRyO+z/bNk9f1VxXeDHn11GNP0Brz3e
5aMCPWvLCABZzL3RdOYZcSpWV5tRQPeemHYHEK3Mcaozny48+/BDCdGsp6qwxldT
mmHd4UpIxxUTMMGXh0uQCWt5R+Q78lyc0m2QQQf4x5Pr1vxvAETdYUu5+Del4Dyi
WzNsnzWAAiN0PEfxzIx25jiZI2Mqsd3p0iR9BMdA6yBlDVWK5LhlD8Mm53OK2Mqh
lVe3Ka+J1QsOTFVuo/qeTKTIXAEkyfGYeP5jJiVixqslAV7a449wRosLBuh2bzOy
tS7w424zEE8zUoVENjEmLe+rBcpjX9tuBNxdGP7lmvjK88z9S4kKIPOX0856DTeI
B8e0icIB6fIbbyQl7ZeluSYGCSi5gv1p13alG8Cj/nuBAEIKx18/hVd4Tv/XjBtr
S9SPwm4gB6ZTVRgi/VlIj1sp8opA92vA929Gfsh1Ijdt98y+Wh5gQJ6NUaDsPCWe
malyVcmMjdfPpUrhnhwqGUnLNJATeqS44FM/9XKeb/zW6ursQOAJrfcEQT+xLrmm
sMZdOg9s1oRy6LbKP+iviIth5LxGQtGbjWYaw22VmXupQ8q/1wYskePYtA1sCyuT
RV+u/M6YJp31jMvzsjoSXaqhLYM4INyGu9U/8OB1By2rchlzUySI15VTmNR0HnwX
um2dTeOWyOevD61uZujO9O8nqE5moPmBmQXiDjkggOYwNVqdzMDBFRh7uh6Vgrzd
3AEN4p7RD4hQn0V5iLopPn4KLlKwED+PrVrzARzXkhj7bEVj4To/FM90q2D0vB5d
M7Gtm0Gmz4A9irJGuBsx0+KkkO4CxsFB9VUNZ3nnzfTArCoBoOZyT82kKibEtJ3c
LDGmo/QoxUjEBbpHRYeR9BzoqFzp3nUijo8OgEoK4ppZBIsHpJjZN2eHc+g3azzF
qBmJvwSVJTJsOeAldlU6KazHHqbz7TRH3yvqGQOajW4LDW1l+2W+GwgAmEk7kPGK
xGFXep2d6O+D4ojYYnJKM//O2WjxhM3FZk5xKjOybaA9PbzSKr/16puY6qjWaWYm
K5u0iZlgBlsLM97LX7GCDwPuvmbQ9Uc11qaDt22GMijT4pF+9kt9rE8L1VkXhzfA
9VU9DY+bNbDYmcGfOUi9dOE3oDmtzp/C3/5J8XT5wl1Op1ORf6ewK8WZI4+N9Avd
XKt0WnyqpZIdl1x1UHfv41hcW1OdPfGhvDmCNICZhsGt72GwdYJVa0MzATgz+9Rt
XYsXAqh4s28Bk5KibyTxlR5TLJhPaH+4zO2EzZA9BTFf8R/5pxbVPdkofmNDJApL
3MwAcHlh6RJlpSHa/OE15G8nVJZjQ8KQ+soLyeVOVJl7mpaiDDiqtIP+Ib5b3n85
H10AthYU7T4kpMM1lLmwjng7YKNCWnN4v+e5guws4X+pxTiO6RxLcwkMt3U3qlOc
gFVwnhekwuea4UksyvNF6GHDg8imXVk8H3XFzEE3cfzcCdMZAHx+pKyHB9wAnHe1
9fiZqwZ8591KM4GHXbSl298HIkr7Nbx4iPj3aQnzEdWVTYc7NubTMlp+beEzbR2n
wSOzyF3wOxDN4tyu3t/aoYxE5KfdIVy2V9UOOr5LuMAeT5wdhRtBIoNQh0qzCdUH
zYmxMfBUflPNBAKNHUBzSi+6FsIQtH5kfFzX1CCKJLCJfMdfZH2Skvau7vqA3z+y
aJk8W7GyvVw0s8aW0ZiYrqQQEmkGcHl0GI2S+/8H2902nS43xVXUnpDhHwoDL9cb
GrHaB+4KlFEdBmEs4AmS2P80jwvaEefS/JzmjYpZNh5y6pkg0dVFO9Pf7ws4d7zE
5xU8wHzq6k1Vx1nnEmwzYtxNrOEjWNJKrbCHqZi+oEsqsCRIq53ZhsiCreejybzQ
RXnN2/b1S9F6hXLii23zm2AdPPxDDJTHYRbQ+JUQ4mCWAg7dpg+WBHWLQdjLFMS3
9hsdhuTizd6O3eNsSbQ0AsOdhoaYdwVjtA2X8JDiWv3Noiac5hUxHUFqHe2Ob+k9
VGehOTF+h6qreG4P1mxc6PAE3Lxao1bVNer7VI29FjdevgIog9y/l7YvjDGifmor
DhAyVTARQka4iNnVS2pnq+6LQC+Y+vrgn5ac+zUPYxvR5jC3VdN7Ql1k3AjttZn5
Htf6/t1UzrjLl9qZklfnSW1zUn/9ubOtsNGNPyGt53cLesI17hDuBONLn7llAgdD
0geMGMHw2a7Mv7I2fLrp6wyqW/bx80hIBkYv7eDpbQmKaryeLuq7+xV+0CZstNE5
WjOLSuMWDRUnsUvurSi0uXkM8YgbDWz1HgqjpyWJl21202oHueQ1QgP1p4/S03Wp
7Y3El5j4HHJ9mXgen1QPNzdCd46a7u4W4a4Fxc2a9rVZVin6EdmR/cUdRr0RCqbA
kq07+kMAaZamlzdO1ouERmFEQDSJu6yealz9ySYBorcdCfgF3Yc/Lgqibg1CxvY4
COyI9ilN5SLBQVdDWXkyWk/3nwmKrbUkQMP4UXjYesjGNN5o+9AxOCRmoOHXAEog
ewabfI1Lj51jHhcDl4qVWWYzszPEh6daFgkWhFUqQfGrAHIiy0MYqj7KnK6RZ3WA
apd6aBOFMUktRQyBe6p8u1pK5VGkmXYmgoz+djPRUlVqG7iaT6XWHcLUHjX6Zq5I
joVOsTzViUK01Ghe4wyFWW2JXqmkO58QTxMOPzBb7nEKgrXtZay8Af3ODLE9yJVK
RivvPcNd9DZ7Jhhm45/nprUnqaYv+iwmGHeRXo88nM0U7QSDUf0jo71lt1o5cfCF
Jvz89e3/7AQRcLF3F1gqnFZhLMeSD3XXakJk2sE7rPUlgnmHGQeTiT1fAB41aMgI
4jlDt9kkN59BTr3kK3fQUU/xPRC3GempyF+YskEOjoUPLr3mxgRSj3PmxoOCybyg
GknLJqKfOQfyXDAGXTUB/L5L004RgM5RjnjxuTWjvYPT276tqZOnH5X2exuMHm01
EGfX491As455cmVoS0rUk6geIVhc+k0glsTlTcFZ/cI2ILFPELPTFtZ6e4RWhU8n
iPfz6o+Lmz74GB5XkJWuyVv+rmpoydp9rmoGT+G9ME3epISalF821esbZCCjyFKl
xIeudr/VrbbmAxolpm3K6K6PKC+7j1sGUJ+k9IltBl6+XtJrVamG4aOOLl607EB3
7qNDMyZnKDkQngdqfNT0+uhC5u0ujtB+3jU5Q1+8R4Cf00OD4tm4G1CI2QclwLeL
K6QasW27SNzUtXGOarEHOP4HNOssBWoxvbvRM1Ehd7gZAzU+TwP49L8lIkeR6QP3
BhN+IsCGHk1Q5rQuT8Q0x5nxl1NWfvPS0ylX0Pnpe8NGIDqxfGHo1i7u761NP+eT
sTDgXGBy5ERFyi5RRhHX+ZxWhpV+K/NlttB02QicZPOvro2kq/o0md4mvQ6PuYFl
J4rNzyR02jlWz7NGXyXHlbbE1lrBxSxwM+k+BDk3MDk4nePAzsU38m3Y8MmAuUmq
zxCOY7v944XlllRtrs9vxCCTaru3xYGfh619udwf5H8cH3EwYwrZnJLxmZEuHEQ+
4O9XIfCtvwmzGDB+RTqbxdac2x3aCe0U6/GkxHYpI8zyFLDU4WldVxKTalepCkxs
3ER7L3MXMuTblM859lGPjaFLRYQeOolgqwoVnoIo6uYiaEX/nrqYsCMcuscGiyjP
cAeUl/VKQjYHr53ex02ijZ+rsHXnVWtajbAmGJDH8twXdRBQpqJO6flh8wYDlYJe
qCSzPEF7X+5PMoMAr74ObT2KEcRZ3CKWuvehCEmiFkrtOwtzrREz0aVpIPj/PutU
du7Bh1yDyoHwbM5bhCsZt/hKMluNzDFHyf72iwZ+JoqRoI8o1be4LaCIwfQfyPfC
DGLx/95OZc3B5zD+rYuwP3JyN1SYfyWA1N1R7vLqGM4jzJencI2vtfFQlQohjQRf
HViiiQVhk7tDBdCJOmHLjcH7102jlSOgXXbAEWPNcN3/PD8ReTRtQLQwgucscPjJ
HA1QWq/orxK8SEx6pJYtYq1skaJ976dosA7HOxOPeKSqwNV1/SL1PSFuNsGgY8xQ
KXekV2xV9a0ZK5CIxQt80stKzilEfVGDr1On2uWXRWqC0UdbzO9NMJ+/1LcU2KPj
Bvy39sntVZ+XYPYdxNBFMNlpIlrKiJ6UkT+NdWkVNjBnRgaz01muH6IwNjXsdXKu
DhIbe34UUI/Caqi9YBeyciFESjHXD9lwz15YfUeG2yAcG2uOHsH9W35chI9BxAkz
O/obPwYmqfJehbrbKtslFTss4k9H5bCe63HbahAEnc7fbHR9lzW+vkGBZa7hw8QR
Fm3nidubIlA/j2cMegK2xXBSVTBkkl+Gm3d4HOxBF35qp69QU7EeE+6pdl9yVW0e
o8qNXN7Tk9vS5sMjX1/8HjqlU6OglcZCblo1nWh6UtuOEbU8+cOj9b/A4HlyzXMp
Omxsu6CrpcJdJCvWQ71Wd7zRjHH83SElLBmUTGYt12FEVnqtQuOKtlbUQIB5ZjU4
xzD55Be4UdGgEQstfHC2EC7iQTLQW94yDhisWLNrh2qNy/iIohfdxKCMdH6TEaXG
Z6/QFnT1H2sTRpwnWRigwkAqDQ9AQkeAlF0Z56yNATeACf/vMXnXzBSlTwyQiywt
jRurOPtmYq2ceOGsaPT/djuTNrGnKi0zGHKlV6R05qaG5X+ZJjSsQEzJ8wkYoxnQ
ybdl2/06/dAhJNidYl5EWUmwUelc00l3yLBGdCsXs8YSlZP9/XN45wxwS3FGW63l
ok3N8OnuG/iwjdGyjXcQSi4IOiJrGNStGLB89kWhWYdSH5BrRisw8/pM8D0rQKpp
sxb0FHKMV6O5eBjtD8587hcv7uza0aQ4njM20Rlg8QXBtnncar4K8NEkt4wd7h/q
tGR+ohPvdEpMcnQWf/fxotMNsndAaAvIWrLxujVu8ckuAQrVZIxB2ugz5Y+DcySV
In8HyHSD6fIxOg8zwRbgCx2aXPxDhPCyVha6V2KuIDlI8RVUWHVjDbIMTCXGKLGm
ZeeAixyQlJz8mA/BbWvQeDpEtAx9mNusQiCO4LTd8aLT5B2XDFnymHStfdZCEWWJ
0yk5x44vKxoTE/zGGZEQ+kblEaWarUtMCYYflh9MeL24JhZLWYZy4SqjSmxjxiRE
d7kYz1iv3oKNrLpyCL8qIf6uU7YBcNRnIDqeUNvy9+ECXlXekYdpqjmq6a6S26WW
+JPU9hWMgtVnA9OC8ZobgbueXKrQkQpkoL57wjHQhBk9vi6XusyXekkxnc2szOLj
4qRUbR8M1Eb4BcoOIvW8FuIMMZxvorFlxrp7rk0dQmTnBBh5Hvn065j+6SQV2coK
O92mybRH6pcjWzPxzTD3Rn9RNx7GP83p+uTDSQ8k1nVHuAKCKXrIGYHDHYdxfKWt
lXihKygv9VzClt0fwGZIlSFRFAaXy56xdJ3oej9cJAYMo1IdsfnooDOP7Nt2Fdhj
Mj/DLs8pFbraK17hga1LRNCuD4LERDNuWJGV1o7KyOVs9JwHUsvts3uZleobHZSa
ggjBny8My/xyM3oMnVPdZcU8IP3ZHtnZezVS21x5q1+KPtKhlbOcalEa51sz75P0
ygFY7WPUBJFJDAw1K8/vbgTDTXMq8/KiXJdAexBURpx8XpS4vLcmOiIAdmczGBfq
CHqRfyQnI0dCIb66J1JsFo4A4cvA+cPHsVYf5QpS8S20LDWYyulYjdK2nZ1SPoXH
fSA/8uUs1WYd2SoW22A49I4Tom57m3mXrrWkocfB3bMx39lkuJZTErzHXGVceM35
eICNumbauy3xpK8MkhmwOdpvCzByz04yx8CsawkC/wJ1oQryB8uk+bKEjaxeWS0b
PEHO9ndQ+cNHpx4ZrgVGJ1gB8uDKt+eVsVWxQ0G/v7NhFLR9zQMQOCgKIfaUu/Jt
7fheNGpLZSy2sHbmM2B26JsUTUHvQosnpftK/hUFLz/po5lEzRCF63EhdFDBi3N6
NLmH4is4JD19c3VgPSAFfUK29k/2Bju4L0F+9wOryX2u7J63L9BI7AoaNkeoLejg
O3Eg03p8P44CCHaVwZWSep/H0H6dNdeyzCQY/AWxFSsJWRAZlrJsD/pABP0hXTl3
6oymZ3AVTApzpqTdTJAsJcg9aWG/XT6HECfMfIIwmyIJWjiJLvzDYil5gK59p5XK
t7azzoejA6Fd4ESOVQSiCqTkp6ZP98urQxNXPcreGdoz1PcfL0jPy+PKa0R6c/bf
3gmS1MvZPKabTWjmIfj22GNE1LiwtmXpMhkuFvMjEccj/BGmsNJdvxqdtb8YIb6S
EfZHBD77dCqwAvl3E+pdVzB360x6thNy9ilFG40+a6eGLei5gZMxHc3p1AR87SNY
inRv5mbIh4tTCVY4K4ULkMo9bpLpS0OnLgjhluh7NAe8NhU2I86inrVZHObeDEHh
z/0vHAbXTuY6BsKeVXUYlgXJwUxgnbx4dyG/IHgFMXux0QyPsLFfymu1IkXXMnjr
nTS6zl3iaJXMsy1NULc4e1GZWpkaUppsPgX51Z0i4WiGisZA3353RaN/eEThqyM4
xNFcGuc5L9qVw2LrWboas0EYrfzJQ9xbAdW6kx5520i8cgd7qsm4kCw4dnUTz63d
5hwkcH7zYTS+5ZpdxQHDCSU9sPWGIewmz8/+FEdVmC3P9JgPZJY4EZIvYZABjK8R
OGBoXaF64XH+vj5A1Vfz4FLKJyS2ZSwfF4xyODsEeGpgo+WDd3uOF9ZoerHGUfzz
YyU+PzKFmAgoiPGOpOSr0Bd6q8SSvPgw7F5ngXTF/z4fyLzeMsTpdHzd7XIlGZ1g
T/y8TbzfaZ6fhwyAdDtgSCrHjmGI/103uyOq36w//k+0cOlwgz+qm5L35fYQ5rzt
dnk9LKWlerNzXirSJkFbJnOIKys+EemoUwN47nU5lfVoVJZPkWCj5i2f1m6/Ijfv
V6IPP9hX/W9PA4VmUx8pgsjNXzJEd+peLJ71bgHo1yvod2shuC6WkQ/4YBl7IYCL
qhQwZET0WurKptddYWhYT3inHtEZRR4qY7UOmOwZyR6UqnmFZBf/eBe3R5YJoyEw
FjJiyMKZf1y/nv6aso4p+XjfgzaJWqT6jPO6IZAdISi+d05J0jogvDrptCzBiH+o
VCeYppPaO/M/wfdiBGHLtGoqsgEBqvgZ70CISJyhHWaOYv94ef/bds3JhtaAmzmR
wbvfTUxoxiUPUjaZlFl0Q57c5LWfvQfETAKd1LjY8kAvYCTqkfyztXNDP+VQU0d1
tI1NrQXNJDN4fOcPJLKbp/ux++1gAdIcsI82vfhdIo/N4T5diPmZxqzbXtTE65+N
zw+ZGJaGVhpGSuBUC9yZoj2X/sfApiT3iVPxVnOfQA5jzRvlC0UizI1OYVgI2y2c
ExL/zs8Z8zXlgJFZ+6/7wqcGwULWP9Ahsy455BAGIJKApiwKs5GXfL0jbxOzQLpw
2Zuomd8H47OonYVGnxGQ6hBgoPpKFSrG6jkqZ2/+efMGdb5x0R6/BY3yHjSVBZz0
rqI1C/RoUDLFEsUPUNPaVml72PyeGK03HmpLJjiBcn1wRH+6oDDroxC4sNiNd/rD
SMUs4n+GgCst6TEOrplOQONSavurVqOQbFUYn2ekbo8TrP0ksPtFszG3+jvMFFN7
hTfQN8hEv6gM8AURH8tYZvnz/PtNQu2X7cQACFV9ixcHNB13mzmwSSwVo1nuaTGI
ll6eIhPUCXxSVIOnFK6PohZFInFoIsrBrAO0cWTbBN1iREDyVpbl3Koo/NJmH/G2
e87Kf2aXve+ZcAlqzv4SzJvagfGrD2UCP7KtMjMVNu/P65DGJthzlNBrLU/hCv2U
rHyHYKVtU/+WqOXtWVxRCpnI0d3Abdbne5jY7Ij1IWKQnQ3tEjkwlveKl79v5dM5
4Wj0U0XIcll+SQZYG67UhvHqKFwYcFbe+xtHShmjvC/Pf9MeM54/nBjyFtuI4SM/
cfANsKCF6JG/+TEFIZ4KGb+ZG2eCUMAraOrqxRWEBRpiMbxhtZSBNoPT8g9NhnbE
bq0nd+FRUwImYSGB7pl0KBwpVcHRdOO4nY7TYjKMpFM6M/duvg7ponGgTytj+cXL
0rcIo+PpfscVxY7xw/nh0a9BN4E/fWipbmO8E+ol1TOeYweTnM+SVaKoGdZU+UPD
my8TTcSi3CmIWKxboqxYMfnZhCeLQkUgOgrQXtv7dNmxnyZErHl37AoQkW/q3/Fw
mvQTPZPgQMGJo3s6XEmErDGhrPEqyeKII8XJ6tZXNV/qb5Us7mvktyxW7o5brJ/B
P5Aw1UiuRW53dQ0xmKGH+9GZ7Zo5rV3WlGlQzDh5Vm4W/u8HuI5JGnFEExE+u3iv
6i1iTHrlD3wSseB4KyAiR/dWwtu8MMQziI90zMfNsMTBV3lSfqM86J8IKJBR8hhO
kpzwiFDbpyNKQLKPtrika4pzSF6waYlChzTiPZer6K2sau5+qRIRsrar6RgC5daU
gnBYOUq4ZdcstzDr6xjefOwIH7OYCLxaseVH/oCl10Sz/jjRXXKmlkydZYx5wIXz
ZS+h3K/zseIj/Qq39jgYlv+volhKSlglv3wdqrOwOpWTeRK17YVs4AXLcLKlE6og
G8FRuq+puhZ75oqCn+8iOLWy4kSiOaTVMfdrHHSZq6fd79wWmOXxzra0lhcXL+re
5QLq25Bf59ibGbJMVqElhrzvJ4HWcsLNx3z6hsIe8R5y9Wwh6+e7HjfM9gUMZHAh
a33fQmdVvGzX4ICm2yb0UmodT860FYtdaULjyXNfum+PSnm0Yh00Hey6n6HXZwoY
t47J066Vc0ml+1qkZOTdofYFMQ0fVcsHMBZ4EpvpV2DVqDUwvTOPRGUHy+K5qYLE
ggRMBUuicJB0UHOmVe6d14URintiOIPjYNcz3GDmYzOpSy+iMSEqAD3Kv61qp7OI
opvVesGf3aMKH8QCR+w2oy0ZQM9J1rw4qjCD1D7bbqZoSJvoc7/eMHpxoh78r7pg
99xoJ8ZDG8tT3QJBVioJ1Qyc+RZI9+AEGMtoNMuKriuDYKw9SgyOlHvArZVlgJ3C
4JEWOpH8yeOrmrz7+UFsmEkNOvCW6BAYt2+Q1LBofjl5xKq8lJeuZq1Jy0bfIg5N
FC3b9B9x+Li2AZoVSrqYsbe4dmXrKpQcDRPcPJERObTgL7JHj2nkdf6Juu8VFaD0
7UvrndV3cdgqj3i2i92L+Hz26MYPSmjc4XgyHeye7yLT0qCQqdwkVcUKMKJxPQ7d
k9jrL+8RNJNM2krDW3E5ES4MIe7T0tD+C2JJxgXHXc/HQAC2v/PQQuGrdSZEL4J7
vDDfs12flGfetWBqYH3q0DGMldEp0D5Kk7uU3ffEQyAKbS/Q/zJHqYoZi3qQyqfa
CWhqsP1DrCtifUW3Xdu6krCUmg5RepXcTvGlnr830LdYmcj5o1LMhVZQdG2uIgac
pEjYEIkI4IZFaI5/LY4BkRafy44TxB/B3ymvIrPwmXF+Zq0kihniwGPwhrr5yrBN
qqrFsScgeM+qK5cv/0QE92aYCJsjZV3FO8ODJF8RVxhc2sHoTxH4qbJ/izeKZMtf
b3/JSNkDzbBaVgamnFmzqwThgzlYQjNh0UM52mc5t0oPJ9/sN6ZoD4AFHP8FiNBI
m2KnD7RgpSeSo2OnIzuObxdmw858GVKz4d4rhlfCH4EwphrmVT5OpfkrJe4TSfD3
AcJI2jQLKELQ07ELPrBZCu0FuEdm4Bgi3LMZ2Yp2k2v89I/S0yDxOeBPqzCLtikb
vgPPK6QqiIVFcopT7T024n4yWO6W+kF1mOwysvU5b2c1oXs/lsX+jN8nxZyGixE2
57z5UAu6rQYx/erT/GU8pPA6k+n7aMpyJJqjYR6sjxfqYHQpSMQrXIQs/SUoKN/L
DfBvt9YkJ9VbPDmaVwQDHJyC5eXvOYWB3bMsDdAqI7EUxtDv5ui3W4y7OG7t/cQu
RAcLi56IhyGqHZqooDHlz48Yax77XhjRR4cIbCBMeSj6uoN23QumH82n+07KHv29
K3fnLlwogNsVo1xmCHlnaZ6Zlo6E7slbNBvuEANR2X08TohVbZWrPaBXvWfg6WIX
QGKaM7RW7Q3vYR0avex/bEKB9jDOZLMlHV3HNiKVUvyzTRI+iXM0rHCxWxeQchv8
sLN1Kh3jURIebGy/qzsYVO+IlpDpROZHy7GvtuCwkwQf7YiCzKFEnFSf+ODfvu26
x35zYp9eFhU/3lIedyVVqcWG/V6jRnL7x+YuOmQ9W+7pMaGiO3A0ZoevfKQ2FyKO
RlJO7JzP+SUwmhAfab8Zuv0pkLC+qNyZj2rM1KgBn/vTFBgLSjqp16reBt3CI9Hm
EMcM3DR/wJg68ZQFJck2NSOKg8qkaljyaPSybPOYkvNtzh07mteLKbqIhl7STWtX
L0ba3HpE+PhFClMMmkVLpeW3RKb/jWDiOB2cvhek1p9sSHZr+JCoz9S8AIV2mX72
JUUu5YhDmEyzHNKKnwthiCboY0UXuOs0tbWtQB4KG/J/5XKl/ES1U5ISc/6TyuLX
WTQ9DjDQ+r6gHD+Id0CYdSYRhrAhKWxvGPMYVi6SXRlJ2nQuh1YqARjb8tXiO3q7
4h6pXey/uUHMyJECyxlmswLhTYYpc+GzcSNnJ0qvlWZefbZQmSI5tBtyGZOCrLlF
EkMkeEk3oXPIsKPOgxq1nQVkNrzjsbkcEzzmtER+b8ND6oTA1Dj8RQlf0pL5H1Jo
7dTcC8v4rxqKFCXNFlQNSxyjRdczBwPUn6VmuVGO6hFA5cBW7BcffVz3PV4/yDqg
nfqAF+RnlNNt1dC7V0ewt6eNBtw+atlcWZvA59qafwdV7nygVwzpp+oTRhaJfPoN
eQULFiVbtOrvJc6qM7fhnaSnMo6AgexS6HBjK2Uj8GNIzHs4kjE0iPVT4/GUiaks
nbVJnoXZ0TvbxE+4drkPQJGUYS2DXKfTlosHHR9k4g40yMAtg/ocFzVHykMdkWQZ
dJz+W5a8LL3+owQ6MKdkttfZxMiqkbzS0bKa6B0gWPzaN5tfG0eOOR6yLoyKWfAn
kOw1kwaYt8sGfAC3FxuiLZb2ocxrplfXIM3EwvarzMemA6tjq3AnsMd0YDyiOhCn
2p0GdmD2Snj4cNQ/Z4CLd+QJdIbuIPfINLd05dircqMBJ6iB6i9YuHg2ETBWFbes
qdDDTsQo/4SFxZMeBuqR3pOF9L0+3b3uYROP3GG/g5lv9nQmd+weWN/Ucc7VfNmX
yb+fcTg9bxYsn4CAn5+ln5RpL44mFPJxhnX1N62jKHaGk5QwZxeKaROYkC3EocMY
/gv8MC+2q6JvF8ApKMLUEp9kY0z1UeViZN7Uwg1w+y5a50x/Fb7T3dFeHuPM+dLd
VMAuS9S6Ex92W+9TCzRtcQNtebZl/DwwW8rTQUKNcN/PcgKHvvaBifg59Do3///G
+yXmlXwOk2cTG9sI+pgLBD058KPtV7EuJg8FPyoRFE4k4a6J7l/BxWtxYR8T2AkO
z8XAtXJC+u+Mt6Q0SZVDQO1vjN7TIvFB00rMQTBsHaVwHDEsYVRbgVOljm+6VIsT
K2iQaBtktqnogY2ln+7TSWmXl7PIVDyHd79SooC9WPQPX993H8fkHVkEI2ijx7wj
fOopHnDoy90XV21bmrhRO9998j4QVzJniaPm0LfSMdiRmpidupZ95mliZ9KC5OzP
Cq2ne1E/O+aR7ILsuUgTWx57NzOkr8yWPtOUUJvKBNxq7jLDpTelpPqno+TctQk7
WlNwFNTFvTJ67zv8D0BwYn9g1YK/jGjaJC4UzKb8XxxBjtPWPqvHiUm2+Yi2iOt2
Ske2XN/1JXPH2nqLu4LlAsEd82vGlkQdHlUXWZD1VfPqKujnbefdCd/Cndv6k9YN
5n/HH4s/CS5/tCeUG48BXIeSQPtmvukDcvjC8DxFj8Sg84KWH08lfupyzp0xyPjj
agdwBQIHsYgoWiqRqZOUt+SeSRf0Wj65ZrpPFzOrQKcAKnNS6jkKTffzU/mDuyXM
lqXKK0kUTvzOtcUJr/6/ONeJ4QRHOEBOPdaywwjGx0vTFseQa0glnWdwrUENP4Gb
thK89/U6lM83vGS9kSjuURoqFOhQM4VccmMIRX+05svuWXRi3PQy24GenVsD/0zF
nznCrcqPy4c+vuGg33Mooxx8fAh+k6+P3MJxfInEj3cPBOiI6WHMh9qTP3GUzW0N
rh9JgBOYpHN558G/oj3VDpnKImznSp7X8vXvLkg2VFRA2o6Hg4swvF2vvVh8yU3N
xA2cbA3wcJmkivSNug4Zf4XR5e6DupPXLV6VNqRih3FzdCHafDuW1JTNiwGqjlT6
9ZEUMHOuMnnIrlWBMIvTMcXHlb9avVRlMWHZk1XQ3N27dFR5iadyBYU5MXBtCnyb
oeZiYaWfgdCd+9hnOIYbAze8DLNkzkNA7x2RdkH7yrDSw10/fB0fCpmN7BERCsiX
X+hs1RiFlAhNzxSHyzJ2pxEgDSrxer4fWDlvhLlJjiIxeRqG82/aB1olPKyzEl5b
J8BcZgrNZFyl+Zx5IVqgE+ZRFCfTQVsr6hjDViOfj7t6GQR5vgIKxPQh8MuLUFzV
mCe48PlTf1ipNRcLlVWttcayJ/SU+EfOAs02ixosrnB3tKLw/GRrckFrox0y33nC
5uyBBsQMvqOJHgrgXwu4TclL6U0Hz04rlrqTNkeX8zkyrq6hBQwD7OFddyVuRSPt
0Ai5zMV3PuovXptj4xK7yPnvckwvLbHBWthWkQCGgkfMwCS1e78wo5AZrk++JeMm
FkDSNHqMILJyrkpM6MbwPd39ihBfzjCI+KDIwqvQiVTuE05lqTyVsrF9xyj5KQ22
FEyv/cypHCk4tVmKI+ixQvRTQWjZ1JUra4xMHRV+MpUrYLlf5+rKmnEoH14y+PZ8
sQjKIoileOOhuEzKhBwMIyeg88xjHoZACOT+ddyIJr9/xXrBiRcqB0rEd/Lq/FWg
o5KZlqFW/iXM06hlWJyXHPAt6tFP22SVdi3Q3Vdw2zf1lcoxOlmPwP5vnlOb9VfV
ML34AUR5uRbi156mKCAYUNdVyTxpuufTgyCNXUarOSISxegSLpaPOi2aCK0l4Z/A
FvEGfjIl9/lcJPHP19gsUWQFxY5QuWQw1UvRwf/rv/Md9b8aqZn8yIKYLqBXE9vh
zsYKC9qE6x9Z0A2DwSsd2mwK0NoVSDHoM68UBxRARThQsvo6bgTDX4OLglHk+kH7
KhD1z+ACHeeQ89FlMTvQEs33/WHMR3DLZUsGaN4kha4McWXSXzoKQO6XD9q1QKiG
ioG0bVx42V4c+RtEWmNgoFkCeo8OpCa0yZ5kUfvHdJfKyZ7o4FWaPA2xCZQlEIry
lHvnP8NwUjnxueS6Wgcoq57HY+3fOt/M5SrW01fD1B4uWIn8ET4K5/5hlv1vPLbq
Tne3OM9NQacUOQFaEJl+3BjsJWOhiSuRp7gvF1O1564KaG3yGzkwIboOu2vaLlqn
7f6/DTzL3fTKh6GZvKa4VW5RgXuLE17WJf0WcIr93Cq5KXN+5HV12YifwnPMrUtE
nMPAkg1SphUEY8zKtFXTxHfW5PuG9rl7s5zaH7yKDwiuhgJbwFUKsVx3aPBeOKch
QqBKnnJ8lFaKpI913Mp+HtknB8Mz8Pcz9nnA8U4MLFP6ff3XtEvJQRwzWoAvxrbg
S+vj7/PLEqRmiQCQ8U9mDkFNI/UbZXA2+xXxnNLSr27aP6nU/YH3lS6ZjHW73ceZ
Gcb4NwZTvacXzeWfvpj6Yal+O1291uec9OpYUepSoUhC/j8znh08sWeO2nN10pb1
J5EAalytGWkc6eIO3SYceZiTJCNkt+M7cXzoGNFLkniaRfL5uFQNBkTyd1z0/3Jd
NfGlz4jRjWGR4SQfLKsDfNqz2oLRlvPzltRsjOnfwv+hQ6mDznjuhVbiYPYoyySf
wo2OIByr1ro0f+ZKVyedcH+clxaR7gCFslIxmd9uXBLg5E9nflwGDErB7ae4e4eH
MWcdpauBC23u0TD3jYDp/gYd27o7uPFYP7Yt+U89bFUiigA7ZwuIZVu96RNKfQI0
qFWwenGidKcz4brMZghHDwdkR1cA7nDxfW3QQCc+F7jqbr1hmxwldMCOXMZENzvj
+y1Ji0e3pWDMxAdnEDiI4CAODDkxPdJXIuYMZp2KR0+lZWIJ6P5tSwMYGOidLt6R
3TDtYztzuwp5KFaLI0Y5OSWVyZgy/rAAMMwY1lcgnIJPd36ZLLmL2SqUMAKv3F8j
3ysoAprGaBxWPGgKquaF8A9Y7C5DGxWTmxDwZC/uh6rvGegVQFGi8RCmQISj0/m5
tHGIsiDtuvvIpZSgn4vfMKRy7IYIB3f7+xDBrQjYfXrQzjlu7z4EIkk6038wCrFY
vKJ0CPhh4VHLtgkrz9xu/O/FPl+ntwxjf4M8s2Lwgi7s3eKVUWD9lp9PrDbV3aqZ
/HzyRQQbsGCIZ7mcBGxies35TW2pztGZCSIxZwaFmpc3UGtu1tJbtlJhkx8SzLxI
6wbOfPn0ZwomJe3xqQ3fKvtSuHgPW7WAStMN6MymS5R5hwMq6Zh/K7YNPMmTbsdq
zRjmVYfSEYt6V1M0s9Ey824VSZK9uW9p8Qweqpnm6YAnIIV3LrQTnpD02K2TgZbc
vd0aZZHDroSII6UJEC2xLTPDjZ1syAtmSItd1XOyAj5OWBOb+LTgK1NRsMwAhLSa
un/5nTO1F9Kfoe4+SJqwWYfcxC9sj2Ec+qy2JfaLEq4N7H86kG2UWkdNQhiD1o1U
tyS8AzCq4nlwZpXZLWLrecnEJ4nzUAJ1jwmxrrHjYd9RfZzubt7i1zFz5pP/o1cU
Xmxdw4fH44xD4b+P+xSo5eFDC/KwAkZZVtWaGXOzpOCao2vFdjaezL/H3f3QzEJO
JAjICKLtI4X6U+uMgGoen2HOfNiSQjDTPH7XzK5/AMG/yaRJiKxK+2XPKvkDuzJr
4oF010l4K9DWI+IxXrWplbBV/aw0kBJokRWqP0I0PhlgoWu/RJSy2OqFXRZ4feed
NmPNPZEUMLiaRLx0jsMpPwUuQ0bCXeIBwlYe+BOCerKU0TCGPB9hHUVBW1FmwbUk
JQbTI4/YSkbNWd+8yraXvW17IKcMR9mOcJOGv8xEFIytjxAZkr8SN4WECJF1llgg
2+t8z5uVepmmR64N9ZCih0M92ba58eLGm7ycsYuoJVWpyGmkDhzmlnyzzeIuVoQD
fkyTgLaN2D/146t8eBEA154CkkTYqETPBkvuUz4uYML8sLT9f7dvLtECY+kHuUTX
cltzneqZAd7b2hGND6ueWp4mE7vvr8b9wbQcSiXxE0c+FqmefR3VfSfAr6HiGLL3
8ZBa4sJqRyjQsAyrMzWT8LjeUEzQQW4LAE/hU2O+g2vT+R8J1zVKEjXDNE2gjWfd
H60nfPbwOfwpAVErD7awZuSxLH0BLXuMi8FMAwNQSC/KFQMFt9wr0WrvDt+GRTkw
bWDI5sbPa7ibYhppZyGQmDbuMN9JLNU0Dz8EzaV1FNvrQcBHndM/RLpRLPzv6MO3
279+QJsU3ly/Mv3pjyBWOm56cRHDJYPUEPm1wJdrtTjy65KE/n5DwZ4MEkVksLlL
j+KYhWSvYUUVfelZrAP71O+a4VM4XXrii8rFJc+NyYJtGejy1HIkf6gCLd8U0oLz
+Smzup6JnXzmC/HM71YKONAjbQGoreEWruugEPWkFAEvl1obdYn+o7Q463OgJiE6
cIEHBr6qgk0DRlhxckMiXdSsok+IL2kYSHgAyQyrv9HCWS97BzWEixNJDcocx8Tr
U/McPqvdAbuiBQXvUeBAnOEHuCcqLKHAav1x56eeI4bhqQT9JcMwwxrzghPBtgOA
XDU9lIE4dcM1LHhC61CoZWTVZtgnW9EgGajIuvi2qLTJ0kIOm+tDv4bRiBrlmE28
OGDfeKXIgUYOviO6DMqklcjXeOHozc36AedTOopw52FsPc4T+XVSflMbrV6x27PY
zkSONVz5rV28GwVzsFJJO2iJ/96mxZPYTXNCMYAHxbm7xCWobW1ocZya6JeR8oEY
5LueZPm8FgcuH/vHxS1m3cFhcEh8EW87mlcumyOgcdTfIUnKV675OXDRPxe8OBGL
0paqnSqt7w5dqPswGf2qPThWMLfXerF7DQHaJT5tkLXLz22DKNtIHq2KJVnAIzC5
ibW4O6t4elzcRCkoUlaL56lqtG7s2zSeH4Om6sZqajQRL8PseuiUJzOmyzMA/diQ
+ImU/+gxNTzTe9Qp7TYhuKbCNgomZR6Gnipw5HvT58n69Ao9aay+aKHafW63GRhB
YMZHcDOAq+r4J1tD6tj6ldYKti/b5o1GIclXs+apFFnHTK8kr9smmj9yEuPzxz1M
hpxO7RfoC/hQZuLDQpmkuDYq1b4syFbDvtDZH+ejBPA5h95rx4+nToyHY7bLLM//
3Vh82tq9A2z5oBVRT62IJX6/YMZONR3k7ExeBzxPcBDobormuJMhRur2PL36cC3H
0W7Q1t1OnB+uv5Vfz5es3w7pXhTU8RGXonPTtPl374PDUQy/yNEF3/OAJr6mBkR8
r7bDZsQyHaBnjoU0Wsz+aMuXqvLA4MbB9EQaEcXGmMgMhfqKEXSj1z1+QGCUykZX
M/Oy6YQZE58jR4/dNNMCqEgPBP5LlFS4N47F/XgUMP//E3K7/wz9jFTaTyHiA2T1
Zz/7jtJisWjEHC59GX7fy3542b/s8JCS3oSJU0BsVIwR+ViKmHHu4kcsPws3gtnZ
4DzAwz5V1xUElfLea6lBRIW9CHKT6Y6hjsVzeT5KSUQOCPuUHifPeXPdBOJ6rDOr
R607bo8tQE33Ugfbgi7CRt0jUbaXn8aQoFpOWuW5m3WWczd5jvbJHlhJeavQQ6uo
GETgCKCFdKdwp0Y/T+71Ymo4mQO+wOhnem2Y2WUMTZQVlaRR7khM0YPt/yGkiDQO
mEMuMkZXIQQu5v7eKlKT6L+N2q/GCciX8bTVsa0bAfCrStBHOlrK6+s1sK8EerQC
7NF3LfvKYsb15FAqK42ZSBzXn8s9UCF/mu66s/ym7tEMTFCg5o9Fuznn5Yl36T3+
RFh8LWpTJ4gLDP6hKhMnJxNt3l2HvOAw7GUFqYSKjNqYT2tKYiK9g73WkwzhNVTl
7JIOAg1es8WF5mgs081DilrsrsFI8+YMcJAEn31rYUKVBbbL7ugEAApbl+jleLv/
0fTHh7W/2JV2uyGZYH2N+xl1/K/X/eVi1rqIf8JHlxZH7vKviuv18gvAdFXj9d76
3ZfEobO+6nqOCAYgUdJwF/gkI0sLI7gi+g9MMhkjpsyGdfVloAzwmjpFfp+vStn1
aZMSkp8Bwn7VEXD3SHuRS8T7MzQXe+cbVX7D9NBOkofwX6zqP0gNYSScHt6iYnay
EdwkGKCJAhXLf/m+7hVvHMuYNN8f7JalMFr+4ChTMYeRWD2WzGv010/WiGJCwvBW
lfD3/dphPtOybKxjeXZOog9DXKhj4Vf4LQsIp+4fV/EwiUBsK+psJOvtTc+KGmVD
TkUv6bGa1JiT3Cwoo+gBqagAxvMhCsG9G10CazhzgG8ncoxYIWueKDOvRijB0CkL
SbKly67kfXDsIBwnXziH+bt+qz38X4NzW8L6R8wIFueN+0sLgj6cZ6wVyCL+h2CW
9LQxfVXqSo4QAENZSHRTZoHHwbZOkDEqMZ75I+DtVAAnQDVS+VvBuZfxQMS5XPot
N4ECnM1l5Nx6/GyHxehfJNJn+fQ3tZofjFEKY0BngJe+fWMyo250OsH/L50D1Mbr
KsiFKg5njZ7x4/uJzIM8XtBk1Btq0F/hnGXBxSNi5jAedpWPJF0UoshhTzopbRED
rLhu03/HWGi3NgWiFw6rSyU3D9524Z9XiuNhsf0G/w3+k+wnca5u4FaFwGWG1IgM
bO2WCsbGPor+o9ip2wFn7rG4mr6/KCo8bNvQtWYKaUAPbxZG1/uzn+rmF4DmC0Cg
NafyPcZ9Wa8NwlM1BG5F0KxtSSAHi225kkhIB0ktCymneuJN/Y3HAY+QrAZ+4Weu
m/RKGuqiV/GLd/XH1FMYx84OZV+i0g6SOIzKNKndWD3wpt2HPkMTWK0KPmENOS7k
vdwUb/xFbVdU0wTbiKq/oZGxTBKUKjIWjgyWo4UwJrQkoX/K2JyLMl3SxzjgksBd
hlqd8ALTNLuwSvWIVsb3CZxQwbdRaEKiPNmca/h7xZaZtawhSl2mZ3GL66RAzRhj
26uSq4UCTZs+Qb32zvMvYZiRACXaA/opRFb2nnREIQuBD0I9YrnbdW9ZfEtlofog
ciDKPt81lobdbr20/LUMCHG3CwX5cv+xWXC66ylDqtt2Yt/Y2+AgKoEIkyn0rZz8
FxTrOqkybDkxFjj8vFZihVBlHDuKsxTBmPmY32jHVdogwrRnZk46VyAqhNkYh1WS
346e+aqlrQeePW+hut2WT8+z5WQHaRYk8HM/UQksTpsfRXghVQeMXUcWXwRbuCIt
kSXDcK8bBfxwZC4UzsAYNaV/NTp8527NXelg6d93OHjQU0oxNnOWUkZiuupm44Vx
8yiWQEcUNZ0BMuCup44v3QJIKcGNHfntPPA5R6poWU5gOkLZIVBV7CmNjTC3ZPnh
sF5EYxJVzlhx9grK1BuMZs/c2VwxcHOaDeUC67tHmMf9eV4h39zIg1ZmRtX4Y07F
br4bM8NUKMNuDS7oYU+9PU2pCowcM5tHEMqfoKFY9YpyKCf8/oUi6gOuRhJYx2tX
A0CtujRILcCKkRCsV0Z4TepETyVhuFnQtcAP4yKTqlrtcK+Izp8e6SGVGwgP5HjT
w1nCdECuIsJQ/uVIH5bTdyMZ793u5vKdNJGcGhwS9xug37vFc9rSrpig5eucMJD/
AZw54EaBRIBl6ny8JbAW6Ua0iuLjdfyhkj1YPfNJN963zA3PS/KnDGTooy/R76V1
HXI8QBiJ1Dvv6SvGEpOUGU1PxebIy+GGrR9nKoFSq/HtAMhqXoJ/GOam/L9zpppX
P4HGKbhvhzM7r7R6hEfn5HRXz4JiT+c0j0WC100tRV0hdYUqs/Yq3lQ0NYPGEsDO
+r8irrdZCszWKMgQ/8K1KdQVrecWq8oW0dc/QKbpwJpUpJCrsIVgWs4LJlhR+at5
a8py2HVuPXuH5/gl2Z+Y5sW6E3vZhqA/UMlp67o+wxK61T4t1QP3r//FyDYWOCaq
WnwvJX9AUxTxe/EcbdBCkn9oJySKieR66AWzxESNlXQMDE6yPsob4v2d9Qq0eqHq
R5P4jif5aBJkFmH4EgZHENZiiJADWN1ka7xb09x63LURXoQPPoccdQgHNXda36L6
8blg8qDrtAjtlXevt5cKrwpWaZ5yS+ZY1PABR1HJF2V8gKIwVApiO6OTsOSnGY6O
ZFnFW2RODrMEhM4U1p66gYIbsoKkyfTwAiOvbyKiAhRy65jzdNcpJRixjhF150FP
kAbp2wHXlQFDpbCeLvn0cw9cWv+GPW0O7kS+UGC/4BGYUwlUQFe9JmX9qWMqL9Nf
a2J1EmPuwbmBc39UATXH95DIzxd3aIeKPNrZUzJuGnwb5/wrbc+251o5dWsUSWk5
GoavcEfdXV+5WAhwXeEZVOZJDjrUm1t49UspLsPPVqeHPYwSYxHkup1IEVyt/3kc
E9eEbfGy/xZp/P5tPLx+m74ogOu4L0ACOg6mxWOKcJgH7lHqTCMpsuU9hEwL5qve
4vPRRQ7CEsXioHt9D0wx7b9SCZXyjYKrMMUR5hdZYVCP396XigrOKE5AX/dIHZlf
Wp7JihApPKvPjCIgKy+R/pAqQi9/q6QcOZrhWEHCVyyusMt9M9/ij36nOMpyTV4/
Hv8hGlfeDUFKvw+l/91t5dVE5OXOlJq3m1H/FwiXP4AHHeDyZFDt9a6l4OG2GrrW
c2/E6+1xAr0pQcxvWJUqARqDIvVY8K+oV6VMXoxxCMK7sn4LoLuj1tW5YRlHdC7T
keYNEShhvkD2EwMeKGDM+/kZlYfU4Rxywr1QPbj6mhErf/Tfa78iUP2V9NRZIiNa
ab+44g26hD2tN55VR1WGU1cIZ5/4Xflfq/T7DSW1/BqqjFyLW73mzdG5Sgl2vQ2Y
RL9zGx+01t6gFZHFUKE/++KNTTkweephRl7gKZx+HoxzAjxgNCyAfN9elvO1Tw1h
LxCCIay2vgACibFb5Ii5y1aLezRGBhx708qa73ssNPxtlbNciMjS77hhHK+lHueN
TBki03Qd7z2PmfQhcASoHeKxePIvrd1KGRLXeRYcUmi1wv4Z94sjTIQE5aDJlQYK
Kmf96BuALSf5Gm3vd+mwqkwrd8/XYE4aBhaJOb8h/B4xzfEg4mktweYSeWOe44Wd
URGG1sXlMyv3sBnJQjA16Hz7+F5CneC1uUmuNbfDCoX5k0hop/sFhe8PBP/UuXWj
8vvtVy6qKzh9F/FhpyUUZu4lvj7/banDRZe7DXsRCxZzvpmJ34uShiwYe7Ej6fEr
+fxVnVSMYO4jGAE+tjXg7PonDZwyF1piF7zgsXlcPWWcYVfA2B16I1K/2DGvCtpe
+0xmjX5v0ZpJEECZfPHgLqXtWuz6sTqtClK1QjmeDpw2HDeAmo+7I43x+n/hfOMy
WEljLUf3S6es8bTJ0jKH1AImsTGmbYgPqExvrslqx7WEkbMwsG68Jj0gnjZH37i6
Ovvr5KQqE/bFerbC2IVwHl8mtjg5ZDYqeZttkItpkypN7jh+gv9ytrHNXCpMDsCg
DISdTsgjmUttjIsG/UFLrfhEq3sP/oSa4LrP7UXBew0ijbbEzeBiZ6fnrhuHfbs+
/DIXxajgKEsZ7oyVG/Ryour4o/JvdEbVaSepdyaInzPk4hAS7VftpMn70/u0Wiqb
zG66Hu/DUPwg3xIA1VoYWMDFN2Z5GahE3le1aYvAHSOkLYjQD232PsANSaXankWr
+csHqTGboxGZePxAUbzJVEUFNc4juXJXs60lypu6lNymK/lfBs5qw3V6MyuEbzmv
nXVmPxDIPWtaWJ4cCwkXNjgMXpbX6FQwAlcZ6jbRwae3FvSLwYcetsqAqAB1X/rP
J3YyrOF56qoaYOL1IyZa6Cv1RdiNDQq1sawhYVvX/4lKQDyZZwgMaKcKGT81gObn
MALPCZMlzBc9M3Int+/bgHVgt62Dbx/sUf2UOrt7ECvyx6LeKhBtGENv0f1j2/KX
nhTTdb82UOBghxqRUpm3bHd6jGlCI68lLPEaTf78ll9mQ5ahYf64F2kp90NIoUUr
Rh5XUcIMG2j/J5szkj1lUlQ6xuQLLXQ21UFbRpQ+VNObWe7ghpzoc774SeIUqlJ/
/WSBIC2OzJFFwoxAhS7hA7AuDM5VeJhmeZFNXZd8EQ4O0fIJhftDPa3dniNNSHW7
ZOOEOQ2aAYgyK7MIegZ4+/oaoO47Aby4OQCLiaHiDT25G1/IgRX+MmZPjhGKby6+
fi8py2hL7pZYuAtowgRrDSLXM+wsVdDPYEeWkGV+6JMkMQHL+FOC7CSooGRLDHP+
KULTOxfxMBqE4dzizOCAzIgdpdRysfqlZmUvk4anOh8S8mEUOpqrsbrg2eupPzde
j7vRFKaX+j0++zJbMgE5mWNhv1UmqDfSVZSw0WFeV52CmMcpdBdwspq+fJZR2o2l
8ZCwXipu3u2Pdyit15R2TgUKI/LWZzTbD7BPj8vdW2c6wjpWZ0I/VEX4r3CBltgG
52PRlgCn7/eUSR7S9Zg56ehwvU2geYQT2ytMOOkUhKUg/kWvrJ2V85YAPh1ykwp0
/569UW710CKiSySCBEoYbxCNRQkRnxfgAV+wBrQ/WBxyy6mESR2L3V2eLQErhbL0
pEoRVKW2FXZEBffO58drbMFGbuDgTUzdnfQuZmZ4Je9xci0tmCXE2c7MHCLm1sUo
w5BB5SuouHTU0TRZ5wmPjkredqCnrKUtWFboRAJVqJRoy0Rn1i2cOMaF3mQJ0lmi
i5Ip+HcACL3YDu3GsP40cevywRJJ8TLJuafkjpmQx7Fx3ee04E8Neh6jhC70w7O2
oyDQx4aa/SpFgvPfgbkLSZ/z5c3pyaCaCssYa2FUf4OgqGENlzNLBLKebvsgVEpW
1TTAQK72483WuFR76wnjgJyGz/ya9QN1xMo5w91o78XUyJ58D3SjRIBHUo++Q/SV
YcAlPhM6H8ASAfK/8X7xrCjUTdnOAcRgb+sB88+BrEEsNmW5abYCe0icVaXhxAbB
Wets5ZnSCebG8IHWrAtv1zP0xVdpSVmyJvLOVPNeOc98nLpOhJt/qlRGLr+8kZ9R
fsAVJbGbgutYWItWm+lg/3hzKMfYDCsYfZBwCK3xFvN6LUIw01SK2d9Wm/0v+Rul
YhGF7wySuhoSGPCf5lQIvQF8ICF3UFktJPI9+jm0EBjsp8VDtQ0BX9l/lX6S56Td
LuzH/p/J9w3dPrfldlJQx5Fy9TIkQG9xMUJa4suEjJYhwaN5gdgQxUhcbhM96h7v
bT4Tp+hIDa2xnpieqV6HlxEoDWcZ7F6oAOp6zoSc5DMfyUHDyljIZEuMs+18c2ZS
jrWt1pzRk8qegYhhZRaP4VSaRd20w+hWQoIEOlR0eo4RCvJqzd6oILzKPBZ5sJ9H
u4ogeqGK/eqBE+8DV8shdhhzk469DtSAi68iFE1Hq29CfGAIqTqleB3pXtn3oAUv
DKrQIAWtH6itV2tVldF+jZBQEFpnFVexOAeP6EVwtMWrj2dazry1nuLISNeOwzU1
6s35D3Y3p0VuZZ05aI588TE7IdhBI2UWBKQen3h+5SrPStjc7TPh9BwSBDgvvEHd
9+uLlVbvP4kb5iCraR1AKR9eaeSisx0vLkijxbo2bfdqpDloL9L1MBQVyG8RRFKX
88GqiPAPIp4dRfSpMLczED0BwF6PkYGkJDUuSkQJqZQY5LC5iIx38CAW12RhzG8Q
Kf2tlfyBrL5on0ZQL6h+XmmbeWenZstadYP5qaVIYZZkuc66HCHC4Ug/sq6iVCbp
fK4mY4TEAESN8NFLPB3LK3JHd4PzIt13sttz7oYuYHotB4P7H5r4VKVu9AUauJ9f
YwP/dYuhgGjZnpv1vTPrVtsrvJVQCi928DgYE4miuXzBmuATPZsxQKIG5/Dd8rjp
JCELru8AYFdWmAONlZO8X1eBSk0OxUuCTpg63U6WKv28JDR8ZjlbMudU1FG5AFpE
d214OH0LcHUuGBQ5u6CZffYBWi7z7lCwoLxUBznXcEXlpQnXXwFBAZ3yXNaIDdvE
Uuti0qRzixfWh0i7QjcBAMyeehtOmcWPA4/8JXQxGR372+SAI6FDoJ/Dw4IgfvN3
F03QOYv5HxrXEN7mZ7Y2hI8WIFd6Oh7VbO82PzibgyUlt34vG8LanKOKVWzHXpDe
doKwCNGwqkN0wmcRRJcchTuTdKKnnKnqjfgpFQhTfRcyFy+/9Yr7ISwIlGHUYfsP
16V4QFxODXDlnQquOJ7JBULrHuTDFFUshgITrXs9WgSHOeBEzKlMmSOOKFP44Ogv
ylpiwnyCjMDQPuwk0wZfr2WZiYiKAq5f6/JfFNwp0xiYFHEi7EDEA5ph9IQsfMHs
GblV6xdt9r9k0OpECRszmCNaWFPyYFIKfug1CNb0zHMMkMcoe8t9IO/A/jZIIzox
uBkhEmb6BInUP/+HPYxuqRnBiSGbUML9x21hapP2go2tTaZUFNmO0A8OL9ln6xLq
Hfi3eiq3nsFMWEDUOirj3LBXRDfHZ1wRlJSThN4xPDjmL6GTjqcTBlJopmGS7PQD
/KMBWZxoFsplxvuubcWabxTsc1O3oZ8H+iWrsTA3Mv74K5dqA4dQSUlBkVdi9PGo
yI8VvLzuedo6YcNIn3IIcjjMrAYz103POO7OudSdw/Rk03ysXiNulrJuWP1kF9zr
6x05h5IoHpebZTzg828QJ+K8yqDqpJ2BlhklExtnMGobD7K7PIWTfXUaKDxkdFO8
CcGgbSGqp9LkAoRIQ3yEamVXIfBmxH7kFoUOJI5nRNPJEAZWj+HRpp+0SXViqPno
UABquU7kJ+NIhwnGq/BLgvWUX5qONVheGu/8vAOLFo5t1YjzcjvaVFkzLp/tiN8V
VNMvTPnVR8pve7vrZgNss4aU4kZQLWXJpjupU/jndK1MDc3rM/jX0xoBuJ95rl9u
2k111gg0QXZ0TiYA7CMXRS4o7pGIO5plB6cdzvpzL1mkQUgCliMFwaSz1NjxyJOH
4J4LsdFlncPVgX+tNA4Azi1RB8b7MDxLSIe6yHuUFdQfQmqA3aEasx1aVqUUxWMH
7Zpyx6M0OCkjK8cY42b5boF3vt64Q/9x3Kc5T8XeMTosObQSyG0N/6cVb+Idfdjy
ySPYOyfp0Y2xnt8ftheoj6LOqgVVlt0Eh1hSXIqZQDnmcC8w4lvW8eV1hPb3Injr
OMqzNqbgQD0/ql8ZVb5zqb+/P407hYpYky8sy9oLAdVRJ2eCTISFsnPdB+lwzaWD
Y8GCEb3kR5hSCVZFr7pTpJpZcit1OcToYr9rnVSOyg415bSegqRW5TfHBhibekMm
ctVChpj0CKauRqR/rbzjiwnCOq6QJWbWo1Xw2IQ47NPF3EX3j/8LTyu56fuWEIyf
ed2l/ZYDhsv7Of9OyqauwBwTNtmMQcYETmAq/phJ6QZ4MT8rm2c4dErK83pS7llb
5+gqMNJNWozgKX12DI4SihP8Bj7STwGckMOvFUwuN6N7o0VwVzvsIPyKfLL6NlQk
r/ZMlkXxltlw95rdJHIaLSmPTq8Yjx48ALLNPsFEy8OYwuhchRV/YCCiCTgznRp5
aZ2iiOAR6YUzm/QFGJ1+0V5Q0qyfqzDPSMyveqLeWNWVm0XBmcfSnOcKCQVeWpIi
W8s04XBIu8cGXAG9lgBCz1iK3UJTeLAwg9EHyP3PQyhBZY6LWYCfe14/Y3Qy0/tG
+uGodzmc1+5o4D+akDJCSlfj1n0gZnsbl8Mxz8Rtwj2dNos42fLUbShlW47ssEus
s8pW8Ud14DgQroKADhfPKgsDzlHtj23dLKFwO76Izx4ePqdjW+qwJFHW7ktDdWbP
Z1HVZjEd/lRxQ4LEUnVRcWIxqFMwYw9Nc+TGXQQfNTbc7h+4vq2dXuAaryRfRPwS
vN8l7yX1wiWBYc2V+CrZ0FpaZuMbCsuUmJWR/GPS0JhzrDdqn7AJfgm73XM3HL4M
SITWxYx60lQJnS5VDqB/4sgI5J46WNw0IdOu2B+3bXag3If+B/eUShmYWU3dQO3x
zmJmiEsFTFh2aBsuQoqXHPEkvjIas2uufGSOLQkQNvr/o52lSOffFLEiMn/p5LiX
LTKugjhq3vi/7a+HEm8+Lb+fJT27RfHP8zZI12d6T8UeW4aBSHvHTNZXMHqLwZ0K
wFHEwg/VfPzICpHDBUCUGyg/+0kYS5sdh5SyajxDi7VgDWJAe2N6x02IVZhAH7ct
YQOU5HiLQugoZtaJy6/Za71dFRro2M4DbugDwwlpSJJZAtJVNAPZHl4SNDcjzmpB
Ehcobtdcw0iaffB+WyQJ7eldcwneJsHA6NCELVcOFmlqVgWzbdTzq9JzSv/1zUNA
KyffwrQvWzD/lJXt/N8TT0kuWiDQN6kV1MhHqDeMuKGHxWCZ9YFeCCCudVu3E+R4
H2bLXercPi2JacmTIJtD3z8HMKq+9hoiEhsfmFhJ0H8brTDTSGT8Ci4+dL6u4F9i
+8jOX4toNdjOsshK06dLMH4PsPp2hyMnne8oT+r319aHuE0Bc6c6R795GdxgYrAX
Qi7WTKTNyMbEsghdq2jvdHubxkAiXeKWKrobp6rSAsiWJV6xezIIgtfI6YI2RSRL
UhxkA23CPoI/zbPpRcTc/lIjTDcfXl+CLGKFZh6lDrM2uHio/i4ndwKwcrlh2eDa
szPQaNMhjR5K/LARd7i4Cd506hvBWjHtKykm+P9anxSLlHjYhuzoUE3/ZxrpJHFI
juelNbtM2FPdEUvH5OfYPY80+490sMg2cZF7m0XqqfFzKVWqgsF9s5ksbIbRAWpA
eEy6OEG82+4T2QOw18DDZccCQFR2MPuazSLXA4zBF5WNRveX4Mat5DTm+3DM4qIN
9xqDJ+aMwVDkqVFIlseViqNacZ7F77Efxab78cvSvDXLgBc7g1pwBg12GHhyxJtK
VK8RTiLeq3CIPqu/M7Z9cXVJSjHj2Hf5ZRlkbklCf9BTZh6UX4q+SVoQ/khPoziB
k0pSV07KZni2yLip64CWwoSS6sUTpWMYnAehyuAm9pksUBASlLiWn06C/2ZFrz9X
C9abakyJFghR3YU2cL1t36bq232qrCzw/Ps7FQzZ7FUdXESL5pobH7dHn5hqfRPW
/JrDp4zcV3tEXJYxSA+qVWFCBu3DAHu8qaZ4BsdggYzriPxT6nPP3GbRJ+e4hqCS
Nl7lT+Lf2bdciym/ey2MJ9lcHhyyissjulIQMCl88IFjPHISftsaGEIbuLfIwtEz
S6xuA4g+DwYfl9vMtJ18c3bpv5Hmje0N7AawcPtz4WUxL8wl/8VmJ9vvjaVjN+GJ
CdvlXrThAnrMmi3rGsHuxp0TQyj2mLkA0VrGGsKydOTdsGFbCGhfKcxVt4lhgjQd
LU2S0nq8PjLwM9k3hJ27gZmiFoa9Jkg6vRLAJGoPxsVxFwYg3UXppOC0ZVkfQIch
G1qavqj5ihYmk6BbW3pBUYOiFb5JeT6nrNALFtn0EDN9/QidoTo4BpLPU9vmFv2L
ArkD44ZEkUaTa+VXROn26OchgoF0B7jNmfCq63sIE90Vvypxr7pYsTWwhRnc7yja
Ks9+/EppSR8HabFZVhDO8dezxFrP9deBuOzJV5yapjryxlFB6NtUuW40JcURa7fZ
2yKNxweTrrx4m5ITdrmMDIyXVp/ZFxYtz7+KBv9Jp4BIuh5BpjKBzcLMb6dw7gLp
0JJ4o4FgTetJxcEtMn8hPXszlsGk46PHdSr9F+h9S2frMfGAnQMxMIBG07fMOQ63
4g7y0Ja8mpoB5BqVaF8XQE9Ph+fwg8RPllDbK2TO9A4VFUIN86I8FKSgJFEHC3+6
JMPwxg+1cFx5r+L87mUCqS/CMrd9RUPvtYfbgcTjjMCdnXtik+AaA4B42hcuqesv
rckDTFdXBwj3ar2DvBdniPVOB2+EecHFl3xtfalvXbV3kOHHXgWScAPMbHVqJZXY
DA2rG43q0+MO9qViWBiuYRxvQ3gjpIgQSXfFDU58mmw75UxcAg3zUZawWvclVM7u
aXAVkC9FKMLA+N6eHsJTwA286CZ9ip6/EUTJePQjzLvowy+S/r3OwVs8CpnMGp7Q
d55kFDlMWKzsILZXXUeM1K4DOodi1cMfl1pe513YopU35KTzPCn6DC1ucdkXctuE
GGFDJoIaV1aiZnLnPcKf/2kWMP9NKmKG3CfEJ+iMYcTPYo8XmKaLoachF9PbuOjP
QzUZsB44w2Iace/Y9tev7q6n85dZNJtNf7bPsZru6JfVUDdIYHwvSY6d9WW8iw3N
ix55XhSEeUUZAOA/U8W+zRSiXiHa2xiMMZrTOWXW7mBHlH10IrdRThMyOSUKkuYw
+THw+lE0G2xDV1V04CBkSDn50+D5IEDUmwpOHnFf9Q7Or7dFpc7SMKJvxDIeS1To
lu+/c6RKx+l2pHxwiiM+tSWgqSmt1LaVPSA8x504JGbZGDg6y4V1goEq6+WHpcUo
NaErnTPovzuWmXaLFBpmJnN4QN4syCe8W018ODaaEosaz/gLPzbwJ62KuCKe5EVT
9KyZASdtND9ugR9Zfx2wRgu3GLeTgwpfNL3PTUo8srcQzMI1E1m1s13s4TJzrmGj
Z0sa9lQ4904bPJNs+gVW6RdwPfMODA3S7geRjLGcvowxZTGvRJ3AUXRu9Qv0XTkB
hq+Fhe+IvInnMpP2zVFoTaH3iLWIO1BuQwYW/84GCwpqdApE9UQRdPeS641hY7rB
cSDjCgQbaNYq1J8xnQ7ga/v72fgONfyp57k54Eszl5P2I2ji1iOYwdDnBkp5Uflu
T7tOk5oq6UWW/oXjIAbIvxn0ehWX4mO2DgjDwYdQRP1dTIQj0wvVMjIms/B8jyCC
WJ+KkZQ2Vg4ltqu1K5p9HH/q5PH8GF3DDv+Lccr32FelGStx/M7JZZPvrlK6cDn+
Im6lSjWgaOBOd0xj/uJmliq7LncBVoq7s2vRUGq8Ci1npUhaOBAy4YjvVg+eGtWF
BBmxovohaqGx/EAmiFfe2dZqfabCJ8HYxgPFcOUcOlVhltcXb4KSwLuqg/Hbai2T
HoXPIivJ6Opf0zfTOkK6aFzj6nhCazRjGsL5FDfCM0fYzjOwEFAqunKtzF0M1CS3
d3fRkpS2gELjAD+36q1LwuNsTun4OoNsoTsYhoZeHYGmmG14mzjeZ2FFtt1BJ+Ju
se6sQ+JdrFH0ixzSoKZ4b4P7v4KrgonJfwOZji0Zu2kMztW6ivHx+4ktDVVjllj+
//RlkcMzWSFM++0OEVYvuqaYpPFEpxaHu28LBCIHk49KSmqGY9jWxjrWmcFtnI/j
dRDkEt6Zz8jeg1F0/0T5BXGKAjOsEx6cs66zMKXolM7Bb4odcw4dikDRrqMNNa/E
Om7/lVnZZHe2Tw3Ql//kPdEAj9ZzDKyvkehG91SlWzvkZYIjo7cHASXPwoSyXhXN
SIq2wGoKUOG1zgMki83JlIAVDcBYcSeAaeenNCymtiIQjU+jQ4prhTFn7le5tNtS
dU6IxGP0C+htZYBS4hCfM7xcuvft0B2JqIz/UKLpLLnp/t4To7Z3Zcm1hJcKGqjL
Nliuib389qz7lVlmsywtQeq45NApU4r04p1pNFk8Q3Ae5dxJSYhtbrdMaltxwol8
FHydSsnl92/kjs9s1LAtflI6WO2XNpcEoAd7h8y0RYrp0A5+a81667DTjB03JDYw
JiPgPJ6RTgwKdMyU3KbGqqtOBuD+Yb5MJwptwpfEBXbXhXaCFNUT5wFAWFPBux5E
ECJKWumjIblP4kYYXIRmmymWnvlQg+9EvlwqP3iWjfgVYlik0RcyO0GGEDA+sAmU
jCK6M4X9pEMjtTCZYlIkBKkIZvdQ+88mGfHvJofNIV4of4LKZs90zDzx1Sa33bUF
+sy3IKneZQ23nEncb+eL0Ix/71CiRpD8Tya2Mv7vErjc/6f0gU7hz14EFsnYdimf
SRSq56E/KpiTC1HEAJ5LzWCB8RUUSDCdchDk2JAW5vrnBnkeucrYFudMzpyORl9M
pxyGq7QMtxOpM3waRZE7lCE1b2nmZT9C5ON6X/KxRixrJTYfEQfcmYlWHcknrDlX
3S1fOrocA9Pjfz/xkjvD14ZUOnpVNS3Gpq5iw4qeRpWzouJVxSAgyRvfnEeBpKKQ
DfH4Jkl7d0C7g2uhhKnsgjFEIs7zNKtvGNb+uAhJu8xvPK8d3qvf8Cw+/FOqseSI
5DYGDPd3/xlMA7XoZMK4ed2MQSUyrbKiX3UcO7nrqkIGl1i/6KtUR75jrH1UtaOv
kEBksSJ5zVciUOHX0vlqVm1jXbnZwKOuRK4VI/Neyk4d80hpPstjAEel9zDrcN70
WBDBqDyTwlXSfhbsX0lOlUeuOhPaSifwuYuZAImKqa60OrGeARy8mRy8+CUyXfNo
Qfb49aYMsjBnq1yIQlxIY0KfXw6IyLQ8MJCEXUNMBiFcylo4JttO0At3Yz19v+bJ
po/iY4xfHl6XX0JpqOejYs+sByWCOpQX0ztBaOs9naLfe75xR3leFpf2RqcQJwzt
4MUEOD8vK5oB2+2vAjhPzSCO29yZ2UFo9ZO7ueGc19ugGm4bIj4vgjM9bb2IUFGo
7KiFi4Ju+4XeWKgV4gbBa6FocYUIacYKy/3xSAuqfpcKwT4mB4NRuoRJ5wlO0sXp
Q/CRGQf5ubAHkknYiRbOVcdR+179Uv7JofNcGm8iSe0bFP0JkO0xCFLscryzBjO8
QaSd1q2LO6t6AL7gc9yqcfszJAx7Y6ahgiwmvHbMgnZn2yHx2w79ZScSEu6srbEh
E43l1o4IlaR/KPNMb3MbewQ8AAVcQVcTMgsvROB9vYElJ978RYz8FnzOKnKEaGVI
Et496xrb10gcBZ8dqlSQ803EThVEJC619CG75bqwrWWaaew8ONuEEeFt4jrvTRc0
GmI7DdbvW5K3SUQ+2MpUIWA9YvD8E/I9Z4gzwi6AOWGCnWup9yefglcxLTOsgrOa
HLlTkeyze4jE4T8Ee4igBeEjFhOiYTsTUvaJy6jnapfDlGP17FzyCQjBhrsNk5qc
hVcWZ1nZuHV6QzsjqKWhBac9d4wX+Q4A2lwVpG2fxD/v1aL8t1b8TzFTHiB9Yf4t
w2K2MdL1rw1cDzULeuyPQwlbP9LVUhDL2kAANies6kmY873LIel/gMLaFZtYwcy2
Bc/xB8nW26EMhOkTDx2GPth78ZD7NVmmskf4NKoCok6M3Df1+sB0KuvafX/Q+bpC
fhGkfjHSrj76Gt62V8WPE5NvSukuBlKyiILNk0ia3f2AOqi97G7vv0YfTiIsjjPo
eEnQZrSkMg9tG8pDwbPIjYLaEHFQjhQkaErKuDM+GB+EhyEAe3qEw3qHm1YHkYrp
oTUidVBvfcp1nL7iLWv8dTBff2zco6UT3vJ1lE+ucbSGbiRU5pMaI4YzCYvTRsIk
S/W3SN8FCxzV9rG8VPNbNE5hRueSw+VOwsjbBZ5p9gnHR+vy6UZ6QqMV3Z5zhOCo
ReeAuIBMXmPEGHFRXi/Whez/DAcA0amtTZCpQrCiPRyIIlOoV5pFwhS+t545DQxd
kbv2fjKi0QP+TZLAQh0ZbpZ14W+1cOXEkk1bYjMdDsRNAmzUwOxjXuqcw24cHIrb
XwRv/rt5+39WMlGzTklfRzYB+/wG3/EdL506E0LQIQDEL7DESsBLG8x0KZltfzfq
5nqEEuAqkfNjU+CHqmY76JXdUgFCNW1+/Yq2x0EIsJGh6qk30uZwjaS7iJdMbtqT
yqEM/pcY4qS5xsKHd3G7wJARJwI9xta55jDBRapVPYjMd5xaC221u7JMRuyB/BoB
lhuF0vq6ZONvy1KnBh+YsCLXwSkUp0mGZXyqtynsRQy4f9YSfi9yba+zyaaxdsOx
DMIU63k++BDMHqBsZDH5cgmsd5oldEUsgUZ5F6kalhgsAnt0YRNctTVomVxFcT7z
TvXMajNLQclHOpkpyzuCURje6ZNC4VnFqu9wFtALCJ19AlZNjSvD3FQJyQvzYeTf
XvsNBtIrOKh7dGJ5v5DlmDrmvRtjreej7LQmDWwD8AYXnbTXSXfix0/kCclRWYeb
AfMJfl6EWb0OA/Jgw1ZyWqkhmXZNYmxSv1NwJWiUP5nvOkVcRUp14yFB7+K4vlnj
Ta3YslgDRLi005rnfI1RgTJ3ytrvLq+guUDCJYoExelGBQoIz2s0AOy/6J1PuOOg
wYiY/v2E+f1lViq24Q5RNAusXmPwALyrqJqu6U09opDNnjyP6WJdcNl/QGyS0bib
qr8DQowJOfjILyC/zbskRq9JcqZYt9OUMUiEERl540RSKe/HVv9+7n2rCi8kteMk
e6JJ1JS1g5tLNs9N77lfLRP8aUX07GeEpK/b7LsJk34D0gu9NU/geGFoRFZH/U3C
T8KPHipLglFueW9GTNN9geG7VynsZLftMa2M0LKf0rmzgytW3fGyzi/lh7SrnPLP
NgHYVUXC04e2N8yPfuiY+mkNeqa9XQ702JL8rqcb45alvqRVTrMhqwEEvC9owcz/
A7GMSe57IypEF0juYLwverd5CF9XSuJxtmrnPh2zPjGg5CAb/4V+MSpRyIGRcjV0
Zcy8GEEpduzGmncRgQHiQHmWl/7EZGG4PFbWV6LNL8UNSKpUwZH6UYR+JAEyehs6
NcPx+DpcJZQQQ6LjJy1Fr41FxuXJ8E2k7H9oKtv7Y1lNkw8N/9/4+BU+iyDeJfAA
9YwMqq8CHlO4w7nbL3d/wtqhHXGkkt2LAEJnfYo2B0/sYQ/IIqR/DkrC0Lb8SJOO
Y73N+s+MAnxOiUqyfxvcGVKTAVkpOjh+nsBFeVMf0Q3scc/KKrHcyREv40CMt8pb
W2JrmXC+CaQzaX59y1vjKdtvpjqvRLPb+ZuTP6itTw/H5jrLHwSF7x1BP7s+mNo5
fKCe13qX6XlsRh8AD8M/rbj3MDvQWmY2MEQVXk7VWdmuXmnW8XX/t1rOuq/LDxiB
jUHQtGmZ2zXKRAGCnSNqXBRsAuPYEOxuRZguFIbZVHRPiQ2KDrcDslBHdsbHOCvj
KJpdG+DsUWutB+8J41nM651C+z4MIwL9rQUu7DS8d6B+jcbUqu1Sozv0ezG2Ljpb
21PobJ9tfB+e0OW+Bqtzfw6ByC8bjs2LRfwmkzuGjQl2CE72uwlPuymiBManAlnx
lvQBXHYNr+I+9kivSjx3yR3aZ8c7VW6g+FMF9Jo64c2BKLkegF9cqKhEBbX7bubV
jQn/qhdrX07emMmQluW14uVpAQRgzDo//w1l90EbGx3zOyZ1GAI5YM7w6gO+UHhO
u3Zl6htqanQARVaT5NiBJ3OnI/ONFWCwDIHxA/sk8q2I/WfzMR8ePhy6p/BvMWqT
REeEdwp3EP9GeX+y+9L+tL7iMfdVFvuSvbPZ52ReN8JaeWvp4ClLl5NoIw0kxPkV
xnC0alPY3p0V5mU+lGAqd+6lQ39HtBy+Ph9F3Ajt63YgUcvK4V2+FECTBpXYcERf
+B19qt4FIiThbPs4Qbdh1SGIzDJnl3xg1C8Xys02nBnL40Qogs8XRkrDO3CTLlqA
fHBzPVe/pQTm2Yl5C9hmP4UOzahqEcDAG6K3magHMCMZ8HCamC5VpjCl7feoRmGo
B4ZkrAT/eQ+IRBmIDbTdWz4jZ2bYkvoKG5umsyAgVeOPk6QJzWr7chIgSU4BtD/O
1yw4ahlaQ+eH4T52gWSW7Jf6IlFANUzwEuYZ8lpsiuMwkIHonN6fQ2RGNUxCHHQu
2GdH9o2KSkqIlQCZ9pqJ+gxe6aAD2IL0dIRQDnQh5MD7LQ6mm8NBMXKIy0UDv+2T
dDCXQotVSNjp9tO3sdJKgtm0fETTfULO4NPF/pt84P/AYpmt3fIL8NEnLos+Nm/H
OfLf3NdkXAj2ecYZe5lVGFlJTJ3+TAFJv3mCdJI/iJ8q6vLP7HVsEL7QJyKIoPbc
Wah0+HkCSCdcziuB2u5mm4l3AfzMMmYPCbnoN90Wz2RsZ/VQelnepWqqbjA9l0bT
vnnzlO8SQx9PCxWRTB2mpdW7og6EhSy4JXveXoxyymLn5l60IXmYjdpYgbR+iXp6
SPVNU6WLRm82bfTHjgdDuuIcblIhuPu6qyQZVc4Ysc8/OwPdav1SY9NeFnljlxnj
L0eqQCks0U/SGjWxhBMlOI5jk79rYKQEZCeqxAVZUqPPApGj157xYC8zujrk+tnD
Zupg7iCBSd0wmorTqxiJgjapsFQjzbPdx/T7+x+SJYInj5wnAq7Otnc7UmFqj1d2
W2B067mOewzc8V3ZAC3rMn9crBqipSCwrNHSv6o/YkM6OdtbuQFBgWVGypfhNZFi
C7InIcatIlYcIXM+tCpo4hLzLGupmETunSq5zvjK+BhCATe+6SE3IC4BWKK+F3S9
QkljKmvJBHNimTuVTPk2e9RnuRuOmOdYiW1AQkkoZ3cbPlk0tFTXMss2FqiwCb17
Tmsu5WFAh4SvLngL6UoLX/239MHcu7YBpYlgMCF6XL/+YU+6oQ6CyJkG093XhRXi
8VCbCmkRuC28jHgpcTRsYwsIbjcSnfyAsVQd5163efLR0yZ7+GPm5FcT8h8gtfpj
tvm6/JdVySw1YLNzlRUCOzHsjc+/+UtguA9dR85V890dfRYaPiLInalagJt5f9Fm
FJ+PIc0oencgXm5d4SsV9bmqIPSS2F3jNO5EObrBQH1zXc7jF/BZEtaQ8YugjLNJ
sYjz3AADhRyQU9Bg8M4bws7ucHZh85B2sDAfTi2IzoAwQhREr1YWTs2C7kX6KcQS
PIQWaKJ5Zcw/rgNU/f6PPn83AwsRDPyytBaooGT2fYBcDSa3W816c4EtR3zsnGeK
Q412EhwS3CrbDD0L3XEAhe7T5Jhwwey/53KDLR2NeJaF052/kA8bFWdfxsUczdZI
t/w1woI2lSqM78cQ8bdnJ/i6P06e26l0siL6CBKtyDyaZvQ+CUGhdqo+cdScDqmk
ddi8+a8pGN8fG6ShGiFOcw25kNI1D5S2VrUB4bv4kAz3f523dxA7YeJfRCHRjB+7
TBiHV6cI/IS6gzDPIfZeJKiHY2NPs7D7z0a6mo3LzZB3ahPm/kUxfEiMwe/ZCNjv
L1FxQMVdboHBTFGShnWbHk6xJX7/zM2/pfX8Gsa3HTv/Eyiv31HwM8sdSks6+NVy
iWVZ1yE+Gevsxc4+Xw4g6WIONslDgS7wjlXZ1GIXhakKii487o7fDtALSEQAeYqj
s5cUZdqO/eCyfwEmMHZWAeRmMgjVxcKi4A6gnrJjGXBP/ao9J7epJr+QszZLqezz
5gL4tdxAOpu+SRHSvxmtGICFo/QuOoV+tYdBzbp/ZwAyv0Ih+EIBr665nNoM9C0z
alPTGt1tbDJkg9F2+gO+y8n/9Rs9uRGRT1dutDRhOt1N6EfLWLq8YC8sOnbfi2O1
PVOkGkO8ZKTFITnxxA+IVwwZIRF4Lr6AMw4Kx3i5dstCkw1Gle6XzpvC4y7sgeiC
ZF3clNyE0TUuCnD9ZD4kLfSR/P+i3dnLMRpub73hWl2Y0Alp9Sy2OSpzuMO3bUD6
83gJpD/0qkebl6Mfrpp3bHi1gI6xVSEJC9AqLUXpw8ZfC/qBm4pmKSCIWKKu6EcT
ylsOkD5QSq6vCN3uX2d8bOxTZVFS5ugisL8nG7WnQugkObkMmki9n7G1XlHAvUCd
LNQcpii3BhHlUCu5CVuYenxPiyv+hpIdd33/GUg8Ed/AHzGDc0UMAjTzWU4NQaEr
EDlPbmi8vMAuzD3J7DfNfTDqdC/Ul1hJhY9ybEfP15H6CODAFR5mrcQzZ1eqsB/W
8xPoV6bq2ezCQE/VF6mfhmc7SRtsUZnei3w5SYWwOOC9oA3l9FPbITVwwFD0CQRD
RHjupKPXIZsiROJ9ZqlRxkVPYIYOgcq5o+QPBmZ8aXwXpjyBMSJdsGmW4uJI12UE
tXtNwh93irOJKy91uWz+mQo1O7yGIfgKaE6uVSs4Tk8webg6nfzMSzgMRil5svXy
SEQHUTvm/NOSCraJREk44HkEMzrQl1dXD59gSzcWgBG+KvjOisnHPtc47YyljTBB
7cENlUQcsyvzKy5aOiQu5ZyhLSaStOiq8bhrTqzxvWgmlaSyRROcPwPqyBGDZpRK
MGa+diP5sj1te2cix977NpXrS23688URxTt7t22WuvSnjdm/+hSWtM71Jwy72qXe
fhbbKCirQVfYRKLTe9BXBmCcz2hnCZ5vlFVapstgI9r/fGbSr/eMr7aSt3bquuoB
qpeADQYxM+L66KdzntndezCDc33V3ZGYzTAT065/D5ftNuVGdqJego4cxQCGq+b8
iv90BPQaVNAQHCzq04kWGM4jretqrcu0djIonQLnfUYLcWkfrhaYi6a45NAxb94d
PTx+w2NHiyHjvX8Uek3guJqETzw1SOBNYa0Q9R+57sqbeDDxyrgQntF356xVmcEO
IQUjr45EiqDlOqpSJsDgBNJ7YlpVwcbJbD22VPPsa7/YexCNPhZsxliRE4qw5tk/
z6SiiSNxR5gZsaJLqfopZ08kzGTU1ABBJ9GWzaS9M/L8zMb3j50ps57LXiycaTBi
r2dDHoI063GZoKevxilmxSi1v4XREdTywwbGlFxgdfSqYg9KHhZe5Bn3CV4bNizW
JOV1hhD0fDDT9kieR+3LzjCgVqqBYtCBNH5ouFHzhG8dgrzHhd+41dQrhW3GljPz
lKjYcn/Q7wSKz4CIs/vhufZGMQw2/1GsFG7fBQT8rM+qB/xn6FqitoIwl78tgmDG
9+AwTvIOv3ot0HRD8S72sI7mtKXl9P5uLvbxJkyrFGEGfWOWpJC8eubzVH5KwRY8
J0Qo4ZGJOjyZDQqi60CbZTYI9KOoboQyB6/VamgdH4H0yWDoUxRJer3PMRRkAP16
3xr0iOz2qI2AElzogjJ67Na6BPunuzIroIHrS6fvZTklm+KQncqaDI4aJUMN7Qhc
Fp1edUdSJNE/oei45YXCBNd6Fpmmx5vBwgdpBsejQqRDB7hRIqxi4O3Po3V4Lyep
9/qQ7+krZzauaR8tu+Y6yoboIPE8hyaljDgV+VxBTkgtNOBCiaAw1uJiTPPqxo7q
TKik92/onuNoFLZRooFOO6u7wJbtgieaU4JI1KtJDMPafm7UljbwK7xAS5bkP3XB
6qfj/Qo0M2XcERRHQr16dgYGIDggfGqjPeOrkUbjxZeqBYIVJG+rVkbwuzkV6xGn
JADU8/Ha1eZdLQjYEcN7IPw212dwOPEs0k+zg9I1o1Fo7nnGcwcVSp6dXoJyJ7eI
DtSyvUkmXQuDX3zd/Se+h3jnTofzOlxrbwWtJykSw0T80MSucfcKwTOsPBMzFFWw
ecInKjRvoXjjnQL4KdRvD2XXpxpJs6cYWzNNnj+05NB8X15nh12XLNay735xAyCb
bIcjnECigVcHvvnuIILhTK/wB+NM6dC26FxQ7HmnNalmjMWMBonHmKlWB8FN2+fv
P4rJqI+U6ZIuDVUz0UMyaQW7fDUO5LltW2DeuPwXeJfoFHSlkSYY4VXU3LbkupB4
8mzdhTBvrQrYONppXmzaXgl6Vm1jcdbADMtU0/XruhRyvqv6chy7/y5WZqVH+QIz
kmO1aLvdUqEsusp4RGzM97brGVRbcFxWEvzUAOHdtZ0drtlPnTqXh/beN3nH+Y8D
RHo1mM1AW8omqTD20HB5zDt940MpZ7LrQr7ydPbKP8dlrTRp06YULo6jf882BWdo
VZ8lLf3WTXty2rQ/7ZPVAWmc1btYJivVQ8OKRp2mYy3fUBX6rXcdo4LxPahom5Il
UMTyUHzta3u6WR3vVREI3wzSMNWfcRh0pZgx+Hz0ABGvP20hVqw/+mkh47D9dzHE
sS7FMY+Yp2NqyW9cKYdrphrrBfOjyPMWQXeP4r79S8EDZEr/dqnPh6m3k6RCbpwQ
IglQYfHT8beGW2GouNTYWGpL9FfQgRzviKHbdfd2sq7cu8NnYU1RTIntBHJbvxBH
XJQjla3kyjGQKKtXjV0Glxfj17fwlcRLCq3mpinLyu5Ndu10j2deeb9w8JV6KwPi
1nNLf4qc4NYaI0U2TdYB9zN0a4G2UR8LGV3o3+q5wv2qeLLNdQ/dLRRXq1cizLlh
BxDELb2qWVPadpSR3ciE13ilBOlgC+WqU96YBCHBIhBAkZ6GOQvyxDBnc9VZ81m5
tpx1Xj57oR8j1KS3KWTXZbEF/RqQnaCvXMbeebgdvpRtYXZOcyUv26gBKtkVijPR
IFw6xaxhyR355vT4E72pQYF0XbnyN0jTBS58pOMD16QT/yh7R05b8nmSN1NGbS15
9FNfvJjo2CIDmtd/JuOng4twzl+Gdmc6fHqb9yqnsT0be/eTQPVqL+Cc1afxd0c/
U8t8V5wzo49tjM3buL1cUYwN5v/n72UuEzZoE7z8TPfmXCZT4ICRf462/ch2xOP0
H+k6p9//sOPPVJv7CrF1oKQSCHdiFAO/XoNN5NcAdxKKBtlvePwHD5+dDQxo+N4h
1GhwX732Q1SnRpmIjrWAfghWn0OaFAPkYPa0CR7uoDev0GrEB3ijJBac6G/nUabj
D5A2W7IWDkjdYorhoTOlqg1iCJxRAPlVSvB8vLi5wGiDfrlqQtWLnmTER3R8G9yU
Zc4ARnwabrws1GiAWHtuX/TyCBT7cqFxy1zHBsWtLduOmd39bBQc5A/pAT9veILc
bipcmop1Z9+H1a1k8EzwL1d8YwkhojQwGfqXBNNEXa6S0v1YNqZukNdiX4/gnFsY
dgRHW+0SeS3hVstFNc/Ig4ZqGiWyPyFa3A4dCFz2am4VSOddajUqtJpcl1l9IxfN
NgyuNfN7QMUZLi0MTFTIC5/Y7vaZodNLE+mitioKssVUzPsx8wsNja3z9GuMugQx
y0e4iV4l62UMaCajMKHzaiRHrvTeUjzEul+ygKWxnNCom9OTmnHac7hrHrIBH21L
uM0pky1iVn8x+ZMpYClwx2DywiOkXCo7lAAOqopB+CDFr/oOqsrbs9+2BvFUECpq
/A73W/44d0f/Ji32cGn35Mx6VRXKLo3K4mI3GOdMDdiJtbfmwVyDvKprwt9/mD3m
URj87O0sqyQbjvbMa+h3r79azvaJZUZusXyqLS1jrp0DT35e4LZ3vgJU4aqIhDKs
I5RpaRyhxt1IKtv6y8/H2Q/T3Zr0Kb4tVJ1PdZhmHiETzDHJSMphkWcCxpsOTPpL
Jcsedcq41CSyZgQiM7G0yJPms8ent5IOLkPocEmSy+r1rrFTOeq6DcOQInneZFzi
qngQAVVqLUzxqS9v9PCAh1aGUNEJXHLhGT26LcnteJARfLJ8DtO8H6OxKzsaY6bx
fHzMBpmSVsorGwm/MR0gbyQs7tHvLe2pyQ3XCRhKIpGDJy5YGQH7scUTp9uwWeDx
tM3cX/8OgYxAM/Elp5Pi4uuefB2PAnnrlXbHPB2izXC0Xiaa2sVmZ19rHT1xZTQA
BtYyCjzptjw9Z7wyXgennHkNfBPzBUvhGhFG2ARI3Z4ntUP4X6XZYaSFBfKJcN9M
MDvbw1Hy6d2kVIJpuuaK6jxpVahA0hHI9D2Nq70gssb+zHzkiAbAV44IVfFCyE7/
1H0Ye17xPCmBjYzqExvnZ4/lzHAfFdFvzQ+fxEwkLa5wFtKBZ/EHN/fymk9+cHO1
SgpOTVexfJpG0P+D/UoPaWzhoJcl+Z1+Nd9wgmJLjKsxR4jReeEpvrt6DvSFKfxJ
fA0YE6TFxzLQRoJoVtIhtaVcZjU0paacYVtqYfFDNBqcgHbnxOu8mqy6Zn1sfA10
nFoOXTi8EGdq+0CX43tQn5/gUTyTXLPz4btKnL1vLybjyN7PvZQjcgMbwUlCRJVE
9/TH3hwPRX4Q77k/Xu+UgKRxZ4zZuioQQKJgpugE8WCr+P7b4SCEAtbS9Yamoxfv
roeGfsKnNUp1v07Edln1LOUtVx4h2LT+ZV5f0lfcmFZ6b6W7jKXGuP+1LRZ5HDgZ
uwJp8XCq2VO/3DIIafkk0J7uVVxeYWWDlQarBcsePvDwiOaDrzm7GIU2AFxNW8ja
xEpfo4YTGcONSMv0beXu70WUVem7+yQGgK44V/rF5SLgkXinGo/oEtKHnc2zL5Je
hbLhKH14kvfe+vyHYk47AZ1DG1fJNbhs5gRou2P/6f6DCX017kv/9YAnVkAE+UcO
/QpY7Gvw4xZKs229TNOLGL1u9RQgIrRmJ0PgmJ1Au9HhsJcyvaS8owXyzmsQSn7G
jmacPZVXM38/114WnMBZFP45r6plrg5BWKiZfS3sX5J8xCmbmhohuSpqAmQ18zRZ
wLQSHEhm9YLzLlg3MNPgl4knXsIw7iBZ+3cdd2jna7DxOBJh0TLk17RBbwf+ezrK
h/Pm0DT6zTGeUOUbUxuwyEgH76v1JEV/NXspR/LP5Yy8QkRwg0Qs+4lGFHoWmWac
6sdvWH17cHDhRDvIBoP4ryGO5a/Zz62eOeU18k2BJzhAtXJ1B4k5qVTZDMehaeQb
z6E9Cj1pz3n3AuuxThK+VvfinPe9kZFKLGy0R5HbQINWusnnraCaBuH+ntmgFyUp
t8ZHokhboYGkduN0NwN2Ksq+Jm/Z/rDE5I4zgk0TTDhvPuY65PDFdETeAo+4xuoS
XWfoagOSQGIafK6Va2B/JYPE9IPfwNCW0hDmge0HvPS6bgBLrCqZ4RQAQXyUcSUC
af13xHzGyK4ACHkdAfXZlumZjKGNbaB9r+j3kTohZZwm856ANB24Ot5Ynscg1Rzx
bg0+7PRmY+3L1Sw32YsNkujNK05MddGSXfenrA5TJinOScTsiAvnwqLb2AVOABXh
mGTEmPtVPMee+x8znydJmZnVsd8I3AekVntQdkC9ygvWdCkZgH6TSaQErQAibwhL
n5aHw3LbzKkBPZRre/07rlesp4xKJEmaSTKuP050D7atZyHw+T7nxuZh1GHib6hn
KlJCmh+a5o22NJhtY8mPXhN6ojP4TO7wgvpXI+0F58A2XEwOLJXGVTTqC1x8+UcK
dPRSPszkEqUYjT/IhBrzWpiQTPEnDkly7PKUQZDxU+ojm0H0eA1mt+Azw1Z9eyOO
3DbwTJvEG6uPeoA85r9F+leJ1CKq+n7hrmuMWxKhOdqPRol4saAU+YiZNwvTOSN2
5xH7vv4qfAjT7sZtTsnpI7MiLiNubAtJhFiCrgn4t/7ORNOYramSm7KHYD47SiPM
40ByDTTjrpmViKUph03lVCAsD61rbZr9Mlw5hjuyxWjx8yJReuKnMmqpZSZfAUbX
zwifKzMTxEE4bz5IBi+0AenZsHA5xAhv/6PUvzlvYX1Hs5CtGzOFDvR3VkPFtQPI
hm05ruZZuZDxDZ5lB7Lj4c+X0ECcmOSDSZQ1xIbHuhlMMAZeUXZzBJHv2gwk/k3x
bGlvvaQ92q1odU1TGMxlfzESUWrjpRo+cenFZZTPPVdePQ1cbEVPtLCNrmLPbpvA
UPGUtI+AcHx4lzS4T3I8BPsxkmOK+0kELo5cpcwDhFGOPyqrWQxtXo7XIpPLFVRZ
pIta0OIyAtRlxaC5VswP5u6W1Uy96iomVExzoOHvi4+lbIhP21PrHSamLiZqpO6i
HhgjovugESUqVN47U6oxz6jS9/IzbynNyv4v4z8/wnZmZ20WneuIuxDcrKSFoCS5
MprDVwKxl8fae+Ffesqh8JqOzSTwqZthRx9J5X7tB3eH/YotCNH6aicbBrl3mudB
9DXzhYJNPcLs/W4lb09OsmjaqomwV8dHC4mt5shqyphwyudDCU062RLkwtw4jzYR
hUB4jYoICM+D1nQtTCWGs7N1JBamkXYZAD+k8ITMn9n8tw9RqftrKqusSLpQ3WNt
+n9CWDtjchAGRzFAA6L/tBRMMcsnrqzt7Rsp1CZl4EGIgCtPMyNhPEZAlBqL2iZv
Fav7jkmlAyhnJABxTsem2jSsTyhklyEgC/2T1zTlZjHq6BO5ibYfzLb749oBOYHJ
k+e77Iq8zt2L1m5A5qcBupFL1a0YRGxUN2TASonAuoXSlz5a6kPrJs+x4gi7TFgW
vaT9F1pebpbk0NMy0BJGdXUYZj5YUxKesDkWsgjFT1hJeXHOVV3jNuBjpJ+YnN+u
tZwx5en9i+ha2VYyxEYYjim6EurEjDRVPRpPOJgIjIU3t/xLVckVMeW8QotoLSr+
cfPOca9aRIvUIMf6ul0S0lV/OTmUGyN1bI6AKX4NkWPkQrGSPaNiY56bH2YGnfJ2
nZqlozgFQ2BbzozC+UAAd15ATgO3OEOq2Mclq9gVErcxq6vGZz7qxdw7wEybk7sl
PnDLriOSXRJ7dxG6pi4UOv1ZYA/qB4e/zvBCVpEUqAET4W+sisXDQdsJizQ2xg8R
6L23igH5P2ATjcY0EGLF1yOkcahaDyMhNDX2z+u57uYTXbUBA3SoJ4uN5VqeaVDW
kDXX9HIf8ZrOTa2kNTouHceyG11FtV291xYvtkaIC45pbUo0NxO8WB7g8eJvRcJS
hfi4WV4/A1p683M0aDLcR26G9MAFmnVrKi1IaM5zc0MUxQB2TeDKzdpbaRseUgFW
Iu4IUmr0jBwYRzhXx7/+90xgT432mVh5lSTjQd+Yrrujnpn246Pg/2WlTAcFe81b
/RsAcDs/TMTtEUsWuOpgkQNas8wt7hx8vJci9Q7h8QxT9ejDIbnTFtyTXb7A7dCA
6I1GSRQeZHvPaRelijf8a1Sb6TP2ymTMLER5QL5vWQ/1zLvdpp+l7abxnzvlBgfX
HqLSamHXC+81xqatDdRzyYyG4yIwxp96aMr6wSoBix1iIEZJaOK8T9Aihi6dLsbt
3OXngylrZSXkd2VhCnxZu+OQ3DoC850g6R7JguQt20jlpIG/mc0S38sDPpV/uuwu
9fAUNkcCzwapg0fbyVPoUrUBCQQ5jz1kQdUPxSHR2IsX2hGpFYLh5PKMlecVU2Aq
dD2/ub2xb/SSPtE/idYhl2z4FLJFu33LIsP9dER/S2qKJ247FOLGBo3SLqmOUhS7
mwFeHFFYbyCSgKbzIvuKv7Z/5XpCNNaTec5wVJabPauo1lgwhiN4N/achKR7aCck
6Tr5t51Qa+gdRGp2eIIP5WnYPUi+z7opXN+ZqrAIZR6dCv55fO2Fs5gulh+ua3c2
re/OSpJfgfO2Z9tjDyII00tb31tlue4pvRZeZUb8MEZkX8K0MVpo5JT31Ippiy81
3XP2wYiSWEPrXQrgIIPbBZtGcWUoM8x33v04BJUz6UJSaMx9Mdy8scrUX9l4QzyS
WHwPyA9yTqGYWwatE3XZBiP9sQAhwIXEUQmOCGJevs96i4awb1CgSCNoVnBLEn8q
rnDO0IZygnt5TCSHMZke1Y9b3p6Ec2QIs5I3VnGvnaRxNOn8GYubw1+dO992R84O
zuYZP4uLUFIURLaqmE/3GiwfonHsNsELmxUv7nY1lCkqxnSYMtVI0a2FAKe6dvLL
HAAWONd9x+3Z42KhWL/8RiNnCO6isxGx+i/wDDzWrZyr7L5ZUHKrvwCczEh63woY
5YCSTtlMJxiiNJwFRP0spHwS9oZmajQs7nqHc2LeEG0e8aBjLCQFBdblms1Sxif3
NcszyFi5iZX7j1xPNB+35hCF/Ql/Me3nmrEC0IedhIcrAk1L+Hpd0S6eazZ/2Er1
cfIUp+ahLHjVlitePVQgVD4UviXypyzmsbcGXtmEIHeOKQSHmH8N5PUX8ExyM/fp
zkV0WxAFMnTw2DTewF7PHwIc7AWOkNCU1USwG9DNUSG0vp7OCUqbE5YXeytQ4lcY
Z43FJ7owvReXqneC1k23FnexQJbcokQQcYA1lXO90NXVcK87HV8WuDegJVsZik1Q
hACXsLY8T2Mb1sD/tcYafXrn1LIwpvkZahW2isnFrh5FNud9udDv8CjhOM+KYbAr
ulaRKAeJ0aEWjBtrdX2ik9TvJ0ytpD2hdzDFNJ619zDB1M6Y+8XCoUkLfr3Dwj/o
Hc9MYh9Jc3Uep+h5Lsya8P/n6A7MBi2tvJQXW9AtQ8S/rUGXOYKQylTNSi3qXYKC
ibClMfIy3TF/PbkBHVvsVFSlT8zHm2bzzE4sV2dctuTBagjieuJKcHoJ447cHgAp
aQhwrhaHenBW6HU5WTQ2xdF8g/qi68CHCmfj8aCu4yWrbHJM31AyXf5TGB8CZIse
udM/RUeK2jNlcqCQmlxzUenA5QJrHJRSxUtIJnNqB4mh8W5D01tLYHup6a99o0AG
sfytcobUd1Z80zxD7j11WcConwCFumNXbxCdM+AkVYC5hhiKiApTvGvzNUuElQjh
Lg1Ou4Xmd3YnM0I7rCuwiWeEWgFX870gf8BOew8zTuvfHEXFPNl563cgFxtKOwO+
lu+9j+z4+BvX10CDn0S46C3gvJ+EwDt0uKd58ADb8G8KiYulARPBLByFeqxhFYNW
Ro430RfDMLtyhPULHpzfiE9Mg2bdTHXpCmwZW/ZuTB8LwgeCdbcF5mtGITfaYY1U
ydEjrIUul7/RrzNJ55lEkUwV59d5DZR3pqOFT/17xQOB4WVpV2gMkd8TBBBcBHmx
rmf/JD3ji+vRYhn6BUlHM0FL/y5Xo+Ecvqe6AjLZc0VLBVkp6ryrppTdlDhXJ0Ow
DZ66M11PWHmSPsQebCeJP0UHrLrAk+kGCMedxPtQroDOR3XlQNMPOxFU5bkm0hpH
uOYXRAy/1/pE141FdDETLDTAe7nQZbmvconiiO1vVZN3e9xkjg21g+GkRHAk6APJ
Yyn6nCzSLNx8Jhp3XsOndfhdnR41TCH8qeSq8DfzQmo6JmkeWBXvaWQTMEEM1qb4
K6e7vSGIXeIdhTV2ddYYmbJ45tqxJ5Z9WoGC67Jm0ylCRDTOjOZL0ONy+2+Sl5As
VI3QcaGd3QagO9DhIgGAH45wfMPRkDaBrunkBmnLNgL8ZXJFs/rV6pBXTnw5LW+k
MfyKxcTlyJzFgd0zBL+L4fmjL18w9oEACUMzVFR8f050PNd//dGhgYUXPXKmecJ2
S6INGP7qnULT7vcxdPpzPOLS4DGHwIu1AIeICN/NEsdwUIb+AADK8krJwQI3/RyQ
r2RKVyivBCPJl1EDE34Av2LkiQha8giJerzoXlkQpitIJEepiMzHO3/r3DAVXKG1
PyOM32CY8q2s9g5bcFwAURplL47UPrpP/GsSOQZG3qRdmSYF9l+Nnbndsw0qSxn/
ySrCY5yMvYjKl1vD7ygJp3q9wyjmDYzhfGd4be6QxrxQzXhFLCXaUWSsRei8sgRz
RJVLsVS7N4gAuKePyGLQm1q44Kd/kurPAX9/byk/orG79CUAbDaBfWw+UJjnwj58
R7wejVu5+Nzd4GBtRVXYwJAB/WFBtf3UCnhTUolLF+0s0SH+EFBH6Mb8iB90J/af
1VKanZmloeB2ap20e4oA4JfUkHlRL2CK8adb6CdMMn4xPdPUNIe/iSmLBb/jJRTl
t+K9zWpBDi2IIeimpsw5Hl64Z44y6jXHvO+NZaBhmj7NjEDbnE5SMqt1JMuht3E5
T/vjHRuFFt4DP2i6yWtS/1kQRBQRdScHb39cj8uEI7Bm0JBc4BKM+OlPqrqQFBhj
giDDbDTmM/4Qn1qWeUrpFi03yC+H3c9F1sSgTDCurgwrUVlnNWx+ybw7ymVrX+1t
o9bkwZmdveKYB25/5rUMhWAYb5umNs5/SNZYR4enYuZgX5inVCqBJ5aRJ2RVKY37
Ny5gs2ftRhTa2vAnnjrCENAYNb4kQDhMANVZJRwJiN+3sio/xzZU+/CDtvbujycH
ppKXcPJnKA4keMXiUejgcRYIhstvtSLIvZmNzS430ujhODF0FhtpNMV1nZVSaV/t
mrWzR4w1CL8vkha2Do47m+q+ViAFoXr7BjTrzVmJ9BsgwH0EDLlT6BdDzcMaMCTZ
NOKjmw/mnwPrlareItKqd5Zx7HkEhy2L6N5Qw+joeDp36FmzNmjzomBEcmgjY165
pw/acAyjNUK38iSoXQl0YuxxP/T16buqz1nSpxVWPXu3zzIbjUTGYhrqN/PEEE+w
uiZikJMplA/2tIAr2Zf6fwjRaV3ozV9Xj086oqL73AL9WIgNqGYSbzSdnU9HWUri
QTRkQkgR0bfibm45Bp/raeHV7WMwJ0s+oqXEUPPY3eLWxKH2EJ+KizjYOgnsX5bQ
N2mxkYyywhD13dMJHOvGmF/LKoFOqe7Fj88TiopB8tJxUpD8jhodo73ZMSMQWQvE
IUY9uYF7CHxZK50UyngNblDG+4kHD5iY3oyLRIhyjvdO/2s9P6EexLHQLfzYvA8J
kfU2uMJbXVKq//S6QI3fWB7QqEfbRHgIcUDUO/IhEQwS81BKreSiuJv0zc+ZTm5Z
5IzdpoBcTm3giPUcfuC2DpEAmkYOcCUE2fHP0bS/ocDWE9GlA6z0nbc8Pcf82Fro
VjRaS8jSUuIoz8yJQmg4cOScPIGbK8ZfjuWDu9CG4UBC1sTUNSR6p+6AdpsxyygO
1614xxSYBSx5HQUjwKg9zQcfbTpbnSFImsJ0CIS9TZqCC1y3WhiBGxnd/nVY/qox
xw8cDc0yrqQXXWauaca7wVCD5/ft+bfvpnknIlYvNgAOzEyjxIljSwWLMpBrvyaZ
627BujhRJ+N8mgjdJZX59HwdcpbOgyrpIj70ZJLuSHs6vmdweVYUnZKAHfBAPM66
RpPGq6k7wMgEgjLvR4qnKqdpV3CrDKVMY854WdnfDyxGwDlXadPkP3llxG00IVJg
ZyTwHrHHP52bt4Tj52H1y7qD5mJEL93/MDDtxYPWqI7AjDAH8YsXISkWcWmsT4Yz
JLbUkunkS0+VkRjv9dTi4mgeaA00Y/Q8Mnhh7wkOloEjKPy3QAhDDy2oRn6BoJBd
nIBJQpZMCLEwRYMzykQbNx0Ql9AUdDM6GMhL7+PoMeyTOc5Z6RCYvm1n3paqehNb
hG6hejttPRSgqXpk7540XtnJDZ9nT6E7v/hXkHAn2xfYwhNhn70/gGowNpcKAac4
o0qGuk5sQpZ/8DJUAtKzu0A1NL+ZNvxIUwkrQ7Yl3JQlBDPGRcTYWoFTshGlRn0y
90BeNGC4ykv8h3Yyd16LmT5H0jJoKAVxJsvA8pga94biT4y3yyOSg2O/N7ZlWTF1
Kns4OFsX3BXy9x+uzKsjyFSMxxifVsEhKpggYY6DmXE2gaQABXOQE6u94EYCkpMg
M106xa7US/8F2cAa1VtK+b8CtU9aR+adfFUrCn+ifEdguHLcQuZt+s9l9c+NQ8HF
XisV/hWTJrrEyHyR4kBwNzwECosi+Yk1bKUkFAtyExg+7VfUh3IQERggxcfaIR5x
nusvJVrbawLlKStxBk5wgk7fZCRjPcWJIdt7Ej3ggh/Z6ZuNZnBq9ganYVatBGkq
AVkBgj1VD7SxvTaanRVbZbIMqxxTqNYWpZlEHcl89t2Aksa8Zz/WY4+1duxDiyQU
zfua0vCkmsknl5MQerBqFwCLzOsJ1Y/rHWyrY1+TVL7txJAIkICYuqp31VG+DdBA
hr12QxavW4OAb/U/WRW3+2gOKXDrvkXYURtsls2fqKsMPFvEm0qm7afpvatlKUAk
jIhsmLrYnYo0FnPUQXGqG9YpzfujJvAD3SmjdyqSrzf7XANW8QN5tc/XGVMIIs0f
9uGnXhrg+8wVPcqdwgBHNxoS/0ti3jaYganAD2FjW5M2JgxF4jWBbGhMCdSJVL9q
U1K5zMmU3BbCTaGtj47TvsDxXnACO2u+y19I06YxodywpNfIjro2jhnJKnbuFsvt
1MpWpsDlwyy5BdurqTf9IDmmWwyag+CDY6hmu9/TH9zXWGycoi9KJMSB0LOghvUp
FcM8WWQAHvhCJuA9McB9FvoqkCd0z/BNcAzkQiO2epYkiBudQTZPTIRjAQm0wwEk
RbqxkBXioJO7mXvljEiCwJKqiDS0jQm26GTtaQLihycle32f935YT9DEBppWmX5X
u1zjJA3gzwZcYakFt9H3CFELgsUFylJPemDnaWyfIkxM72Nmj25yR+3N0MYBVWGx
uWQejFZ3lhfy0R/eqS65qE+zm8Ed1In0sFjp1ompf5tSDT5/Opbh8rv3sdnSR92T
7yLn8ak5KC7/oN+4NqezhUYV6ciBsKyxNjFB/8WYQK5klOj4nAXJ2Nt4mXgE/B9N
agq0ea/7NpuyYFdO9Sj6CtRl4JcfsH/khiJHBn4tnCXU/SV0H8cIbgaildPniEt2
I8JrKTHthgjp6pQBdNzBsK0eGv7c6v5/umTN8eVjkZ47fi+t8+YQmoNubWcPT8zj
kfJ8v0TzVtoyDArInRGxho3Tu1i2kj1tcQdK1DYcc9i1Qalo/jfyGlQdBFRUIkUn
uLbqnicpoNiMtbGj2rg7G5tuqrohPEABquVesmpyfqpkGFjD1cnp6ODCk7cwcHCT
l46H9D45s2nM3Rh/UWnRWBcwfCGM7M5TTe3khaimWi8LcJk+wag+x4lb3N+ViqWW
rqbmNSWM6qkCWl3zc4UFjHp66R34oBrCMqpEzcAaBY7AAH5FYh59/8D63jUgRM8H
/FFN0rynGQYz0pnt+Q2tCCJJNMA3dQOTIr78Uo0dvlfzHUJKD92G12tTidqAq/oq
CcaurQkuvJYsRZKViY0SVKOPsNTjRHTUXsHNAQtcXalblqT7ZW4JgqS29eypKJNu
btsduM6XTNUZbN5d0O1P+GN+LXF6Imn/TJ0zfBWLk0vCWvOtnAHDkKpKj+5PK6Yz
vuPU1dulvdJLmutJRMrQKd/JmiDfwH0bQkn1opowaHQAAxzevWZfsFRuXmxuYQDZ
nQKVCAHzW784EeAh2bB1UpyHSsMDsG4ws/iuqdvXXQ6d6T7MRKC1DxmNim6rZ2IB
Al03zQcENbn0DpEcGy8UOi4xsf3uJJ7yw32pLRa93cLGxE5ZPEaAQuPQAVWTPZPW
Sf52vXNTp0slAdS1chr8EqNciKxlsutEb4GgOwqjq8H5rs8LhJS8tOsJqhpEsyks
o7QjsMlb0H1UvLvG2/WTCMVar6C7RbYoqxYRxH3PXQ5zdi9lf90cpous+VCUuZgy
L7SJ5FIl6pkUKre3lM1vBEURDhLJjRxrwmWZzy2BS4GgoWZGnwVwplC5XGrXCszE
myCvbbmqzrSreb+hpYk2hT6uPwGxeacXICMhY8ZyQcNxy29bW0ukvzD6cIwF1qjZ
+q5gEYK9VF/ulGPtwURoR20bGDzr//265HKG+iM2sCWG4bO11FIh1N/A25jwP4oN
RpLNNs6nrOs3j1HmYOS8+0wJStUiyX8Qw4pSqGbEulGB68CnkbrdikK6VgDfxday
JKqMXTprTGXDrp7wqgTgV69shPLlKp8mwuW+BLF+eeiZHLBLCF1v4rN50H05l+5L
1tCrUPAq5n/N+ocCNrjCLrNHlC5w3viv6IChvzuSpsMty0slggQqBu+E+qqZFIvI
vsOoqV4KKaY8lwV2IdfyDnNCaMsFLlwZbAz/24EqG2sgesxLlRx4WEXOgrMYP9h1
VJmyLuI0n3x5Ad7uvkG58A1VOgqItSMby5hqJqgJTXrcR1BboDCSRkfdhZcI9/Iz
oVieH5lMUImUmzItIgfHDrTlIE3EKBZpZb4fe396OJT9bJaU7IXHOVRkhrZblApF
uTX4LhjZ4DBaujPEF6hDmfepuFuk4A9R9mz0ia7lVlaJ1E5BXNhkHEv2J984P9Wa
6Y6cUq8/K/b/U4j1ZP0ykS+A1lUJrqwNc72iHG8G1I1sbmuLPtW3P3eOd1xwuXmT
8w4Js7ogBY/O5BiWVViRAHrcCzZ0xpNuBwRrfKvYh79cHjjDfJRzQkQsSQGYTKPK
Zy3o18aFEm50BqWKI53r3rQNbm36/OL5FstQXWNc3FPw2hpbjXU/RJnWGsiX8/Ea
s6G9oEddNbc6ptWhyJwrIbnGVsbjPstUDiMoT6dSK060XGYQtQFe/lbJFb7/zWOP
zdTwsGcw20IOHPXMV6IBQmM0Tu8Ls9x8DLg3OoF3d7x3TsmRHBHRBq1ZgZLMzpPB
SZa1+olSB5TcECOr2rH8X9mutRfGMfyJ2NTSX5FeQkZn+oe2kjC3hPuvSJRle6yF
fGIdQ1gCfhpvOnAqXKku14KsAHrFav3jtz4+u39qxpKcJANiT0WIJD9FygeySn6K
Yn98YLKYJZ8TK9cGGw4k+IK9YdWPAZY9JfQ+vIbEf0gChk+hDe7RO9+EB5cSfQsd
9FG+MrASxda1i8PZCwEW+SEt/LGADPfzK6hvJu7nJNW1RXVBs0b2W4bKzFb43xRW
pSUOt1YEoFO4LaoDtf+iZqzf7jspgamzcgCpeb7eIyY5DLcnkq+ANitwD2UkxOOF
+tR/Z7WE0+4aNvt7B3ByXeHKDEcedInjC42UZ9MnGRNTzwIeH0GyaUydPnFVeg3w
YUWZcVnK27MSpwPY+RWyJtNzir7n5wDeudEyi43G0UxDOQfyNVA8nsxiURoQUUQi
H2EVHZeGtKOYca5z0RF3K2eKeerneNSzh9Ba2T6e4irmDC8kOGpmEbhSYEgdk9Vh
b+bq2F5oOdJ/T4cPjS65HEenYtNfZkX3GjpzeesrxGvTLgsRCGNBf/H1n4dFAdPr
MPMz+dhug+obPh4Cw48dFV35Hlfy2Sf0wgzaYQ+W2q+hDG37NbUAKGw7Coi0+Fe7
j9pfMASOOHjaO+xggYCZvTVH9hxlTN8BGmX6UDV4VKtoM+/mhPmLB95oMd36UNML
AtSdCgCLwVUHuVSCa2o7lfwY0EhiNfrvs7lei3tjb42wjJpcBrSV24BOF3DsoBIR
v5KaxKyV++UlMwrv57vBFIYQVPPUsDa2lpri7C8UGiRP9cmXA8xWb/Bqb0IQtpcT
bXiD/2nbtOwEFS1fU6NrWpt01oNFKCx87CQw95bVj3gPeX3+nz0u7+f4jysR1O2o
XBWzKsViBuj8R/9MtavfXA/DjsG/cp56QIh49Sy5V8DSSCHVmY+LNE//rl+7zbIM
uojNl3rNcWhwCmzFpZaxo2JfUhXYp1Yb4Ff2P6TIoNVaeehpSH82p7rG/PK4BYc/
91yqbXw7Nsoe5oQWURbp0Wm1Tjf22mVskPf2wH9SEG1TaHO43pA7nToiW/ce9Toz
1appLjUpoG6Wg6ui0AKAiXc0PHIafrjzM/LAXUfmD361fMOx4uriYhGi9Gnubp7S
wETgiRHtgKI5nSPIb1yaA1VCbWzxtIhEtRSADwO+sqoPDD9+cS6BRwAwzOaX4kbH
TmFDJsoCC7ndpNxMrIoteNDbrfyqoGI96F1x9dHrYsKL1aPnauex7YzkNg96i/z3
pd6SaJLldEGOn6yrQjNAqinLhGK/xfPG1BxyfDF4jjSA0zblYShNzS6dIO/ceL0x
4W/B0lAdIrm4rzKS9mFgXGVj8hJKPEnRRsJNTGdivcFqh2qS5pvPx29VrfenkVaD
EveH1LaoW6EzcBEUkq/Q+9I6MNyKyV2Bvf2WX/QN8Z/wGJVB+C7lMLe6Sgn/9KJr
in20ZPGwxCW7dAZY6tbdqAc+dQq+XEEJ+qCOD8l55wrBOnnw4KGvuZB0jFfMMFfB
+LyIxp9dWiy42Z2dSw9xUiCZXwuP3w9t5fFudFbEHUPIefWM2UWJ7v9aby36oQLl
69SaW1bCJK3vMgk8j9A7DecMLHFTBWeNWgASiZLsnKXVBJWYfD2fMmpJ2Sti8Txv
UfbYHjj+GIQMWSfCWogfB+0L1u7cc24eHONqqrBLWBdV0HFApHsirD6p4mOnXB1h
WP/VXm8q9qIZn1rXbM2KFen1cwgMa757Q4oXCKNR3kWshPDUJwTAZcyJFN5EZ+wk
s1gaELjXmDvwka322AMlDQmq6JK9+QrIsUkJRtOg+ORPBU3AdEa0dgxk22nTzSv8
QZ+yBnPwOag6ls4q9uSO3+mxGNJVPiPnup21HtAa/ki0x6Ir1MdPm2/YHSpeGZtM
MPbFLSpqImxaUQAJyfNi4irf6ZSveV3kJwlgsibqOpoi3cPuth6R19H95W9J9iQ7
rItQQmp5tandjO6X0tVfpDktCY/3+BDS5/0wqyc9JWgxFKai5hZHP28vaxVRYUWQ
XiEoG9G2ecX8kHkw8J8F9p3od9U6bWkpESqmI809nHO2XwTb7aGHPbG+btbPMt/I
83bxOiR3cTFcx2CNhUTMOgcWYQDA7opkYhmuoD1WZmtIQrHFgMQtd9MhuPIswcJl
Wi+mNTO8+h1KK8xzxjeuMis3oF5Ax2F7NdplZhxuLe7doj6QOAZW2YZkVLu1xwYz
rmj8I3nWSVcvU5kjVQq4UdBkbwr/3EmGlOr8ZPLUy50FU20F8FTOmrO2SarsjLYK
s/Q9wG3a1Z3ZFYbpNFvyv0zgqlD0IgRGUkS8TfyPoWFTQjN7vG9TN/Fw330PYHRf
1VK94gvRxVH4+3Ynb84yeAf99fsQ1BcDmUJPGG96mlIvr+pwv5wBtf0ao1evfxm8
lZh6NXvTZigvCmf/tBzHE4YBG6mpg+ysF9+XLPIgRrRNFgyvLW3bk/b4LNou2bLa
Ik2HEGBLjpfj0VOMlg+6NQLazw1uy9Qj36t7fL+nFnWamGwuZ19cmdrRypwGp2vK
ZZiwZbCW282TIE/06o7pmcJbLP7eiSmfgNUrgLbkuYVCXo+GUWPnlRbSbnFb+JoS
KOMClSjDyxtmVl+utZM568ih9p2y/cwLG7V19riKa4jLO4eUsSFTLWGgMIzx3uOj
kLFY67KCmdHN1ZF62ZVQQ0OJa95CxG3bpWOi1fXbVgTRhKPp272IK3kQ8e2tcrbW
tHsVDGxenIt/wXaZxzQ9b2838a6wlMlFTz4V+t+6fDFY07AxvVubHXxDDDJYFNW3
i//YnF+kujiuXDNFDZSCYgEsycR1CIAvRktOhlJxZVEIf1Mc0VxRmSDEnfOGG5oY
mJ6j1rrs+jw/kep6KUpiROHhve5K/yBrZqBTfSRWHoO3rLJruS+I+OOM6A6rDPUM
LUHetCtHnz2Y7rRDIpD/bI+bnd5bbEPs2dwNxbKyEylOUPjRJ8S3wIvhNXkGTMhV
lsHC+nhqdyClLpqN21GhZc4OPSCzBazTGxDGNadW3xk5w7mwC6f+rB1ntpBHy61l
p7srxuf6oGCzcljWB7r39mj9eL8lY1sOzTsywhd8ZizPxYBjbCG2CvurZUYTedSF
DVVndw/0B0CoPk87GicKn2GAy1K5fjx6vo7Vxpo3A5Yq+jqbMPFOiknTpN9CRE1L
/GinTEPCSV2hD8BoaB6SvpijEz/ehG28WvMRnioeOFiadLRKkwB86ldMCEsHX1jv
bhPL6tvWs8WTaiCFCkJek03D/KYngc01W7JWmDat0TNrISsvFwNoRcZMWBjKgRGM
5EJtQ9c6kVrDK8CyGUg6F5myK2ZNUF8LUVqQ30wR2HryvwSYVB5HNnCPSLtG73aQ
cNbP/A+m8Dgjh1z6tQqRPLUQnXVBgbRgdYy/Uw/UrE87/1RRTLur3mSx7ASmFep+
+jey61wbXfzMP1+shdUsBD1ktjPjc5n6im2Q+CmaSzUhBuys7BMrRwRDoqfxCS9X
MNjJXVxvDsupn+hOLI1ssazEo9m1LlExrFAnSOmi2hqVwagjKVeTWszxy1JhZpXL
+7zQtyeOCtSLiR95l8BY55Lv7AE/KVx1CxohRCeMeYXg0USEQpa+YU3OsuPpETgi
LATdjurPsVcUlrTw4E84EzjvYwVE6peT6rKmW3dVo+JbWbIDF+YRGrLcG+XmFHho
lSJtc+zREQPeiXw0bCHz4Zcd5WI4YtHb8pORwnoSb6fqWj+vD7NbeKFSC8B6a3jx
b4szLBf/O0yW4xlD7owiXQTvTKLHUN2hEihqYurFpzS72YDDA5JkPTRbdNksU1UL
1OFWlrPVu6eVxRJQUj9/CJnNyVyN+jHl9qzgFPbwZ6/n3mgFS+JkBhfHXcQl4fJA
TAmx+Mlmtqg7LARIk8mBQUqNCdj12xRofnPwjE+Y07tyBHpWHT2QHKwvBMdeMNzr
x/Tvn2CphsaMAo9DijGPHfq1po4olFiNk89PlcWIbkKkt6GuMpS/hZtlgZD+2lEB
1/hpLF/Ar6cbz5xToROiUi1HSeEC0ThKD0tK9k8OX7ZEqr9aFAdwUmkKmfLB+3uB
0S4//sj+w3pR/bThW2iN5wjr7aOs4BAFhrPIkexzkK3LzfYFW5u0gTbCmaAu0kYy
DT3t/TWcJS9HVVAFTecbqgheEHpjmhf6tsUTd6ZzQqI5i+L2B61sejWutUaMh7/F
4SO/ktFVrYdhACZZblDfSeb/cG3Jb6I1lZdikbyJBYZC8XkU7Uph6Heg4SEVClOs
jfrKLiHoP11y8S2S0WUY3RvU+vaCcmi3fYal6k+vc62e6iay5BFrOQwsyrWqc64r
I2sYX5uWgRVu8rEPEOBpXAvG8sAbjz2ItdYn/nKbKywS06hBtIHvWMDS4F57E1AD
oE8iqjrJn9hG8nV9QyWws5mOsyMqCjCrq+m+LxTh+vaPAl276if39X708HWItjfV
X4lI+oSdIsfcfzZLz/1RP3uxIe0jInZZZ9/F2TWB07XYgfDoAzOGfq5851ucBaYj
R15uzzoX2dxOmhkLNSudWX09BW7AqBWEvemjMJ30zeIWbl3hHLAMyQd3cSnF5Gvf
65NpOi6ox8udLdXfaLFOmueVBPiuGCXk5etaUbryYEei4GZVZ56NQ+/HoD+JRbtT
So+YLAobAZZpB4XdlKfwKt8NgSYDahp1a1FUNoSIxJ8p3xLzTTipgtalIV0hcgI9
HJcrwutPoX9piuMWIjIiKwGPA2EwwaofeVts/eot1aqsrGdwP9CDhUlFc1/iWH7j
VrxRT6K9mx2aYn4zP8sOFo+hyglH4W+fvG00dr7g3tERrDMBmWPrJeS8w/2OBey2
0P1pv3BM5BU+sUF+0x26/rT7onVYp2RIW8S2aMu2RaY+MSCZtTOSf3AcvrvTYvPm
jzCd9MqoL9aFkNySw7hbgXVB7WkU0EpIWmP4XVOydfdFK3IynkFBJXYb8SMBD6x6
2/QC9T9aCSzbsy22ESq2/ZdJTxUSdhYAmjTVXxWjonuboLUAzLuVaUtebkIvb5BD
LXxbQjaZYEUQwIurrVlJSEJlmvq3ixt3xbyKhTn9MPdPgns2bI+VzdkOIvS0/3FS
tuY6d4q/q1wU48C1YwVJo4ifcGl1ZAYosb0D/IPPqfOoWT+6IAf755l8DAZTgG0a
oGKBu82XK93kNWtuIs2E2BcovK+VLV9Ckau3A85IUR4mzmhClUtjWyqntM131UeX
XpU+4Kn9/GBbYPE/LlbbtDSvXzovEkwNaI1xOOoAC2awzgRwkVl76Gt/W9yOF8Ci
X9j8Ihnb/m4Q0g+Jt2NGRJ1S9uM6GujpoPxsmrKL4Nppcben5052AQULDh1Wtzx5
1PpKDl86KRpNAwDndcq9EXQ3DZNlH298ecbmCZd1fnPKakFPAli8STB7N2ugWV1K
6S9R1cHQBX+fzHFkqCf4ZRl2kTD7uUo/pg+0tbrCRr6tL+Sjr8Xz+8Eywf7v2f19
2rvwrYrD6f68fSbpYMJkYtEbwm7SlLxGkrYXsGdbrcoC6FlTU2QKM3V0K//2OJFo
UHa3Qq2vIjRDzTCCRY+nYuxs2siXFK1TNnD0G6F7qXuqR7rbKTR8fOFPF2OjKVpP
GoRH32oRAZkcZzs90Dt+8F2Aw88h6FhzyCohczLNfemUStvD1kEc0vEx7DmwzfOX
A40wL9Pc9rLnzlHHMmRmqaL9GmSHnSFQt4ijhlrvLvymbia0qFZ/vunFwu9AM/J7
UHgpqNc7Z7Vp1SOzqolAuBmng+hvxoyt/rJJBhgX5BibxHeW7t9bF3wUmfhO7lsJ
8ysAx1Jb/GbNqivphUEbaMklwNOdVf5TkkxT1YmpPPI5L9MaadO+U4jqdOIS3sME
eImOf0jRlD9rr3qceO4BXsSc3/CoaVHXoL4LwYlsyNgMyaQcGWZ/y0CaFfTzIepQ
hmBF30qgDXMAY/y7gWjp/dTak9XSvh9XnippJblJINGp9rCh71sh8YcY6kk8+fkG
6LYQpbn5qjNdCVySg5CGPHKnKjmFlGp+Gs6Jih+jaq80rmng+ocR7mt+kUbgI8LS
S1m8wD2PeV0L2BjnalwAfhI9bwclqxL7aNIKqV6CZ5TI7pvJwycSGvYty4QWSDua
dzCqw1TVLCGLw+HshDpie8v7yHr2bRMzDylZZmAmZz/F04upu3cC5FFTRmjg9UUe
6vwG36IKuLJqCiJfysM6QaHbMFChq1kLXyeODUXiN+RyBaUq86Ww46gndALaBirX
Z7Y4PJvz2YHp99mryk5KI9WaGk0fuL7dSwWoX/ipeN0COQnsGcUsWu8XEAj/kIiK
j+t4768G4JSXQYdp5l2Dt1HA73ySw44lShieNJVxKmxRF+l+pmunsOQOK+oCAqfV
bZWrDDEAN5WHx3rGKfYjrplYvQMh1L1JAMOrBGIC9wcqnVFATzNZA3j3h2TqavrY
v7ilvu4bUxxbeXeBtNHwTvLfYG+R4hllUNIL7Qt1JsSa5joeT5xhxfo+LTVZ9D4B
lwOXv5TNAicuzYppMjvs8oj1blfE52CsHogm3kVFdUtQXm28uYPN4FzJ/k0GASPp
LcFb8z92sAZc0xL+XJoKmt6qRvukSo1/BYvbMDqcFeB0T0dEgJ53DCbuhl3sK8ib
kKVEjjasEgJej6daM7X5lTWQfvGAXKT7lz0yTSNLFZWkDRjhBzI6Blh60dW4klXh
hoq6caxee6UYT2suRm4ihBL35b5F/Wafc3xEBJyjo7dSXWAIMROxPP69N0mzXmg7
jlz+CpxT7AW/2Bv1Pt5FTWHnbpGPu2t5Fwt9BXHZlL+SRNNduW7laiSB0D8SBG4n
C5tySuenBZQBdMPpZvkIPzfkB9bsMJUSPmWVTXvJdFjw/KLfQXu0lXBYng/ejomD
CyChQlloqv8+Eamyx/dRtwhhHNInPAHRAFzzC8UzCF8hlEPXheo/oSzoCjuK43gK
kkSkHMRu6ETSu518pHtbjOqLTRxj56wV3PXSe2wdaNBSgN+1ud2jJ1tPaofq5xF8
cns+W4wAV5GbCd/fl0qch/nGa6zNJ2Kn5clw7943CsO0sTYElEvb3PdVpZ6eoXsp
e3HyGZIeyI0kHaHor0NUb1FJSDSUXfuSogjvtIpV92m5HoEIXwgcyc+jitrkNP/z
xzYwa09/f+7r9IDj2bjrsMatxRj4xc+2NCQpsQr4p6zSlldLH8ICoifgDltJCXhS
bIPDgpS5qfd4ALuT7h5fHZ2puLnozDJGLAzPCNy3GTiAfoWuVPXyamS5sn12sT8W
M4vmsBqM1iiiPThg8ixxR/UmEAE6BMVtXYYmc8pM+s/eAtWokYtUNan2oZymxwXC
W0aZmniFj3kkOOx9RT7CXWxt4eAIalB3lH7Re9QEejDn3NknM0lVZSJqDPDBOU7j
BwwwfKEnlugBs05kqyUwCaIf1MlL0LyPP2lOFPBWM6Ml8BvarfQRU/yecN2PGZXC
ICwEfXYMfB5AtSqbBw3lRrXsD1NObE+BH4EV8RiF/qTCEmYU/gJVYo98Q+mvUHqG
g8lS3SNFrwmXSNDcWFtfUQM4sKZXp8MTnkdDin/7XWAO/4aTpzPv/YS3hRdN7n+B
Y4SS771GtAIAp2J7uoDnPLU+30wcKDzk/Q4bExA3YpsVOEljIooFD8tdSNhaNZPp
ovTmKV7hLS5NJaNNzWxgFqfBgnBQ4y4PgczUlNwdEev1Zj28lZcrhv0AHLmxHUqq
QllMs6sGGt2dtuhQ15HT/CsfkFkY8PwFJNWFyNL0Zzvf46JeWs2A7vXTdY2FB0UI
NzEs4hSIDqT9C1NoaAPp8MT49Me2iGClgK7fbXYYt5aLCbFHHxy81Id5xw4DXJSL
2DCgydvXB9JI8tFOL8JXo5IcLE9P+A0i8EertX6r7nf0zNTkOzbPMHWjW7gwXqJm
EVHe0fwSvivmjG8iitEv73szgsIPjuLFKL2Ycf8cJJFiYQ8MI/LUbcmmXE2AYr30
FF82+G2TD6jOYuVKvUPFXm2bBxuhtCe9zLFCDFmr76EJYSD735WjfKQ082d59q6a
eN1UPII2CNcLGyavM40+DsT+t4FPNCOyYPGFxnnhznT6fsigD8DLlUCCpdd0j+i6
yBEi46rOohcap9k5jyOz3yvSTaJfz1u+IKejjm49oCwr3veTauhtn8siquYm48zE
7vKrejMSYD7ts1Yg+02zbzSYfKVkSvZRPhg1CJeLY38BowGLa0Mv4ZCB8VnH7IiK
db5RxIRrOs97fm3Nrd8L7UJlHX1D9/i0FcMvu9FxgPyml3zlsrINqm7wwWIZKC7y
5cnaKaMwNMjFzzAqRZI2mQffGfA3lUSbgLwe+uMq6l4HQKtPoxVKchPNd+DO6jGR
/SHrIG/23e8VgomozUkZHAFzy1MJF6kNSBlM2fyRwcRsID7yH+h2hqTPpoSDKMxy
p5sgu0IN/AWcC1Vun8/+9aorXGmqnSx1G/R+W/QXwpUtgtQhIxh5CxUgVPaVz6W6
4gFA6PrqwSzcSb0lE9/UNZbtcl6qN68Cv7MNiFZx/738+Y2V0+I7FmK2WMMxk+Uq
ZRAbRh9h5mUn6nQROZZyAJU/RsKVi1dNU6COFfJhi8ouewXLmRiZRasBDqCYBmmt
jkV8h4piZvjokGXiay16tJnLPrFUVQMkZ2hZdO7ZLGFw7Tn+7k4KrkQVswjkUlJF
DAH592xRwzibWvB5km0mocevxUNFS3LQj+gyyegGhz7mgQwxTAwjjKRhKVuia2H5
ntbtkDgayC0/WH2TuxcV/jqikNOgvmccxy/NJguF0vP1UEc4Iae+sempVEKq7uod
XFi9vKO4RVsBrrABahEUzKDLklH0sLqk6aYoVn3hOMRD2Q5lHGe3UO4FKAB4+UQK
3I8b3XRtdrZJvNASI3vSBmrE1r9sANMT5kjhirsy1dOuYQlTR2SgS0RAkfKjp/4C
fWvlUjFYK9xKqPfZofqCWUvwuqVyrJtzZ/avxK9XHyafXHtR1TOUx05VbLDzA4Ay
tMDCxqOQIJP+/HsfhibfDAvD1qAxR1jwzfhk8pUq9MiypGJyp/kvKC4U2EJYdBaV
OgU7O6uAr7DUEqRW+EN6AS/poHgM2qproG158ySPNu+AzaIHYhUDPA0UxsbEVzGw
bJIYIRiZ+vbsS510W0ka2YPEbd4z8j2JhzSZ0gBGP2zSM2Yw+WUnoRGJp2GPyUZv
9jkLXlTPWep+qD6x/l+Dc1PDvOkMI/HmQ8hbXu7le6lyd8kjVGGFt8SJKb5TV2KQ
Sj0Vn07UfY+gcVX9vHa6GGl43xZJ4u2G1Cm1k5OnP5KO8bxniy1BmNtwYGzpb2m2
arCJ3VKEB9OLgBEMAd4glU7MP3tTXcoVLQ7kJb7Ax4lFcgeGXqFzqfJeeFhydU0u
RYOvSUFMPRLq9BbMxXs1b3JVCnJKRV4kS1SVCb/t50gBwtCgmsnW5m0TIt7oKuIu
Pv6HaBcQD/xnYNThMLJZlqXnNMVCCrbpz/L2pBDT238Ox5xVg3aRkfDP0goJwPo2
5cJCa23NF8uwfngURv5eJF6u2zCNsHC1pEi7WdU7OL2EauGEHkusdRDZPf/titw1
ctK27qH093Irr9abXapxpf2PTujqtDKKK3/4L9b7aVw1nvdDTQQvQkCAyzNdCIqm
LoI8drKTYDCYorcCSZHmf1fYAnhK3/WcW4gLVPFlQrTehyRnQ2e8WC0RFOii5Bza
QE391g66iut5m3xQR8wxcZWMrcXSl0hE/Cdqd8bhLumiggIanWa8nTCg40SvD2j/
oGhj/04wMHyt6AiUDWBWu1ZLKv7AEFBfIGz1BX90ilkE86H133cxZTIuyrQkLX+c
uXZLtpYwozFTRWPjNwmbWUgYK+W2KcSfCKIYzR7+hPBgONYpd/Ka+HCq6PzVEpOw
q8KmvOf59qefuFCPaRjh520E9XI6GTLsZkNHsv/1+KGllO+YmUEKDDZgB0sz4SX5
YDyzvM2EE7mT5PRj5tNb6A+Jb66LOCX3lwndD7OghW4g77Zlxt3fJ2lLwW9Hl3i1
SAYFuug07ulCutG0xS5szGDW11fCKwvhIB+k2iFOmehDSPHob8sCMQvcjAqpCr0L
ZbscuGW3+qFxqq5d7HFRUgkAjAO1UUczZroAwQOAwkjlM1o+i8Uvgt/4fwkl26Do
DqBPFkcEMF/O9RbUnhal+F5LcwNjJffd9uYXQX9zFdKR1eIOGDgQtw5lYrh466FD
zDxF5HbCpMP5XlyQKhdljHBEZjzwz186n81wMAHB/Kmqpf86ce8AdxezFiHGHXTb
uAY9+4Ug2zu9Cg7L83isEDlfXx9EuI9x8Im8xT78ECGM31q4y8oyKMChyy0bAZPt
yrD9pYk7XzkhUNlqS3DcUcaYT8AInyQYwYCzRBJIuGIKMuVkNZeYbCr2C20Ivvyl
CycpkhNKjITaboMWRb2Z/z8TCwOUcMsuVhbfpb1XNBI/TCQ795FSoullk2V6Hk9v
j9HpnqKHvix3Kn7lbzBp2f8sK0v7rtcdhiZ/f71ab00FgHtiEwDMaupdCJUAhit9
dRbSYS4rNSrs8keQXvZNg+ux1rOwEZMxlwqpOM/DlG5CUDV0Cv+DbSfDBSpgCI5+
moq3DxQHbUOhhfCvWyztCdXjq9gdHnV/vXBgbj+qZU7GtOaak2h6pidmyQNO8pSw
PT+kRGfGidmEMzo06Mnw3EH+w1BBsh2BMP780Nc6EfPZuMaKL2wMstWgeRDqh3Ma
Er2HDlvxFMCGfGrITfFr/o2Al9VYapcN8BVfzF3XGQdQ9OKfiPzv7wOhPuxC93Mb
tUyROv1Fgd1pHnloCAcHX5UEgBuBMlrP73eIRaBOzVDEK5PXzT1ttgUXFAPOW/4A
SIRoUC1u3GiP/ArbHvwLCtfVysektrWyN9JsM2sw78WNT0om53GQ7n085DRkrs/K
aNrbqLdUgH9kSytZ/jpZVVCVb6QzMqueoKOghwh1WKp3U7NpV9+TWnoYb9YMBrXQ
BkSme5uKN+QyVdvxC41MkDz6DKLwV9VwQXU9XmGD8I1mdir+ZzfTyHrhverl3+3L
C5zJsduTUWiEPOAzLR1cDqbkS18is+WPiGv7zNjLTDxIMw0faR5F+XHfdImLIFL4
yJM7Zq+iPn3Owt7a8yYOA32VmfRf2aAfsb31bNAWDgpiWkHpQCUClyI71hWDRp6a
Oyi3fx0S8kW35i8mOUdDHA4tgmT9FfpHWeFjRx/8R9J+d+zPR55rb5zuUS3TCznl
yiokJ4ARuIxEuIzBPwxxpNcapbamvs30fWMKMSqjCJiduAra++TJZ/wTQ/nKO17M
2gRl9NHJ1JqAqzgV8PdqZXqnkn7AHbiH8jZ6uwSbR7q6hZ4yU5p8qaR3vh6dV4mf
6EzeA5ES80ocmVMdJgfFoej79JCRU4T3CLHVhd+2GDm5WMXXlEXTsTrJLW6FNVKm
YPa0sCDPPTxFozfGw78BjZiO7LjtVeN4/s2hS9Kq8rIJKrr3GdohpsSPmS5eIa7g
376PNvzeqLJwb0hkIl7jd8NuXobICVLcDrIhhwVY/AGYVt0T/7gWh8jmtchLpGNS
IUslqJu2MUY8HK1u79N5WR6DLXMKP+XFtzx3wDDCgUb5d2AHQdiBB77uBMmhxmeW
3kNXYVzXJVZ+9UIUi2mkpaT4JsltBX//hNHCFJtl6rAokf3fnRx4QMbrlJR7MTO1
hm9y9TNvCUhjhP5XSC5TVYI+XwTp6EN8jy7gRja3yZw3mUuEwyoZFnyBmqw4kQrK
LQeHq3Qb8dxQ2SbGOtR5ompil20c6AfcfY95jGeP+oUDN1YUhN6x+jU/gtj9wbq8
qYPvkTAUgBHdqAF1K9cISITOGrdZC9JlMgevhhUXSOZDhRpPgzOosdJJnDKyHsEp
I1BeKFd2/QwNyQI040jpfWaB+1RzQTnq/CmJxTJSkIGmrQDauxie8NR+B7Hz1Bac
bOCS7m1s/ugQUzXtZQd6gex7Atb6piiu4chOUw29CQA4bcnSG9A1IpF2D9+wr217
ITkbV/CRPJsFTGN74MRtZhoohr3aIoZ5Lom9TR5hoIaCnObZRTnQje08jV5WjKQL
VDfimFHoU/7du5iGiFvnQZlCfSAC8JznGZfsxPgYsfBhJDkyGlvzsQc9QDZlQkxo
IHx6bANfE1UYC1AtkprvM0NFIwr8eiWOcf87c8Gw8PHgRfMaOD71O5fKte0GKcY+
GSULu2pVuEwzrVqL+3TfIW+xSPpoPguK4xxiowpwTqZYNmPiTpE4S9RrWf8qUi/0
oxgTOOjm8Ef3Gz5U8WcfNdxmIa/Ecfz47sx4daLrN9bHZKOZj7zIfEXQheVLC+EA
tkTtwg793Z76Z9f3oqlYguChLiKdg2yL4k37Mb6PmzKAht7qNimQxq3zIuA+n9Iu
HeEmuU9rRfgHIzfuYCenysUDeZNow5RD93jLxGl8oW8VU/j/KTE1/LmUeMcQSosK
cRc5l0s5KDBEfByfCf5aJ7eshzFX/2VFfXO8k5QrUde7hEtc13nrgcRD2HVJEgqr
D1EH2m79VEJ8y7yxvbWkJMSu+IYnUpHVgbVACgWKCOPI3r6xyD63XSrFhgqYx6Kz
CzXaz6Tl2VLYBFHupN8POzH8nNsqHPo/tjgr3CYQi12QFlAt8S0wyJ2nAfr3OAyw
75f2Vw8dyawKo+dYbIa6I6Wcc6Y6QViVe6tI5as7rWpwn89wv2/X0eiazVaZZTwz
ok1Nza04UQLlWiFTEbFNBsyfAFKcb2auXQqICug13xkBsnClvb0FhtpUPlgz2xo1
fT+CMWSasP6CETIsySL77szTyBy+du5Aw26b350GnmkBA+GuUaITo7YmoQePeZ7S
BCyUHp4pabNZ8OwIxzQ+Aug4RXoprLwqmlbIlIkF0cX+my+Uw/Q1wYP4IofIDtY0
D+gD4Z9UFGf0kj0RgV56YQAgo/dGboHT17IDooeiwN5ETa5ZWPt5no7I7fYyghxj
C6wHfG5UkGscDurAN7oqaCHTf+f2wX8BI9TeikI9SjaVaPSXv8YSxPdPnq9D5hC6
qqZ2AowBZvi1K/HFIJwgNZnfmYy6+xIVjp6v9r9Gxh0YWnihLzmvivEbLS6UzqQV
gN7cQCH2OdjMVcgrO4lvmCvAqs8QeSjDOApZYRIjL3elbo8fwCifcsToOIUNCVzN
7EhrJfxT1TbX7QYBWoCD48SBUc4BhdcHZ0DjvK6nZnuhPRKfIZqeyOkJMFnaMoIU
+5pLCrW3MHjvtxjxH66fYonC6g2NBRq5aSOAuFxRGsogequWje9eXb7HEVJy7QFb
tRTc/C3OH6cxL8N+tnhDxwym3adVeXdCtdJ1vmvEskildXjYqfrardcRBG2iBWbE
BtiIyvrCK45uGdNEEMMyt932Ey2riHyPLACvu8c6kGM8lDEt6SxJjYXBTklXWxd4
U9TRbMPjQXwSq2APYup9lM9SbbPY3Qcmetk/qdRVYzR7R7HmjbZG4AJ01vWoortC
kWYXdWXmmCcKOpW1ihv/V3J2itwGkiRi2tM8hONWzpFNUtkKDYksPQHq55s3/nWb
tsyKAKLeUsAv5vjscvGKRsknXpCusnc0hh6idTMuV5hryrXliKeAL6Yj4N1uCJaP
Wq2oBokjnsCJn0jAT1DLmCHz7otNylbYCqTXmEMUKWzt8MkSVm0bw2sTpJlt+YA3
BINWP5ygUSxidt0q5BQRKY5wmLbbeDeimhrNYEr2sjDXF1uiZ5la5drMGb18rUDe
kgeCg3Xp0s2ZmPyh0xrJejhDPWjNYjtNNmS2cHk5/Su1+fPQLpar0o2EXtXLFtIs
08B/fol9decGwOVjMv/sHF+hedBZHhgnhhRR0pXLatgVusODiyeBFug1oiuHddaK
eP5bGJZSegm7Z5LyDdr6aYKjahHKl1hGepaYHPG+42pkdncGp7na/KY/acAE9EtP
4wvVxhx0AEXpTMRJWG86N4sNoKvAhivIUF0fgRtKwb49AqiGLDwc/EOIjZgIaRgG
bwAHZ/SZRZBU02XTq9p06qDnhHXTlsedfQ8BVc0QpdbxLOcMrGbyX6Y37mfvwUx4
P4Da5xzLR+QSBtTRxIgpEkBVfigMIJu8KXhaDRpS+VLOp7/cNH7jRycOAuPLXPXb
MDnPFwedSwReweu4BEQdzMqbhdVZGTTblK8IhExN/Va4SP8fKdN/4kW6h0Ycs8mK
+yl+NMrY8x9XWrb5If/eXK2k6vYfWaRU0RwB/9SPKMLhxeFVrL3cGN1UcG1PnqH9
dvZH8aev/oiDajYAAfUTjaDRFZ7hM6hr5zS+HxaeBWR4oGuff7HnOztYxtk4wUle
8ishszk8rooVsfoZXYNLay/ijXYIpPhTxTxfYYgcIKbReALJ2wca1vY7mBZ2gB+y
uLa9Kny4qczNkaj3pkcV9tFhm+zyArb4VKtjswA3kqArraxTZ4e8EXcfJjOI5CqP
A/pt4HE36CsJTQZpME94wP3/ioM08/7/pFxKqCx32ZKi7ulqK5pMEwR/OY/Qj27p
l+0hs4094KKNSqyyxxdVNg7zbdw0nhXhzUHhLp1Eh3RP/x7BhAHWhAOTaatQForK
OvSdJ+m98huDLSs/JTV6oYSMAYduUSal8HZNwXiUJwDelAwCGG9Jje93Wjt7wxC7
U+4koG1HnHNs378/Ex5dC3GlJRyoMQjlgLRCCdTz3QBSMYynJ/QfL9RqNtedvEzj
drOZs1jzneO8Q/2TkN9yA4J3KUCp3s2zD2i7rdpBD7qUVsF+PDRa3xGp/8cg8bZN
I7dx504+8psWPtlnqCq3fx7YQ8KVi9ZluFvddsAVUz0gGSLU9gfZg+lkz2WisNPz
3opLS8Si3s8NLUFsu03bu2ANJBHXI0Ij0Y6Br/sHQT9vblVu71rzdT1IhWBkm6ja
SgMPP7s3GDaQ8q1+CiTAlYevYuK/iFSDeUUbW4ThAz+3nqvfD6/JkA7otETUK253
KYPbPCTInWJgQ8pVNVLvSolrjLCxrwIX52fbPU+VhuHgkU6xASThbMbxBTMspfI3
QSVQcGsEpnSbce9QNDAvRc5/oFi5+2GsYfRLFcB9lwFEl1qGk+i8ImvRYjW8NTdB
X3VcSYnlCCF5cqyMRn8E4cZvIw2S+MvUmz5bp9+HqgUZ7M8w92E9wVSGNy/K5cj3
qGgi+g2AKNSTCp9fRTPS00HzDkfvIWkr+AOQCa5nwvFlwlnqkdHSgheyQ6uRXdGq
MVKh+es6QiqAnMuaSU3t0exXvmMQQk772FdxbwO2V816D/DcOErdQs4EhHlpQRUd
2i8QZS+XyWBvsVu0fIUZTZDxTk/x0CQcrm1Um2v+eKvX9whGS0DCKVw+8MmOpIzF
DHjSteKrRPf3d8/XD6GkFrXKvQI9T2ACShHYEZHNQp/7vuknkzODbXzwnJstdn6W
z/Pz5kykNn4XQXJncB4EvufxPrLLhp/zHhbhuVe1N8L06otlzGwZE5i8Kw52q7Xs
+3LFgyjR0u7kTS0dKgxYpSiveFpaWC5dhCpmYfHTj6pzkMEhPCOr3T7ETjNGXXZu
+ud47/t4pQ4ISzv1vEC6uzLF299fDQ96mLyKD7ti+tFv+iUw2NEpT/pRwmpEisLF
27alDFM3qEp9cUKFxEtV8D6/sO2a9Ntg2owDIiRpNe7ker66KcnpwZi2vtCR+Tbc
trQzfeKE5w/8tlYqB1cqF9dtrESNiu23biY9UZ0Egkok/cHsQ1dF7BMovdGGDdDE
PlBr5uXU7s6lpChz0vA/TjZg+/TGd+uGpLmFetTaffsq1eg8DtZHAFTHpNLebwK9
qWYuhMOGHHOo8+IIGrl3e55K1w/GBoMxtVRLQUtvEEypZ6F6K0c/ZnOnUKrRT1aO
ju0UfaNMeoVfze8IvwZoc28m39yJohOeT2qo21uGSLj+VL5wScMyQbj20hsjQzJu
3A6KvRWKteddAwg3WpDgid4PrffordeUfRwRfqsHOhCRSdNqXVnqmfa01w4au0Li
jbAk9YbrOx5o0HUzhs8qwBg87iMPSkmRDPdcIQ9RS6E6ibvFQ2aIpOTPQuEtbUmA
9gzmTYiWkAYgyNxNBa3hw2gEm9t0VNxKsMhOsch5KM0lXxE7W/hEFbScbhsqoCGP
iG0rs1R1I9Qwhoo1sT511gXpXfLQwanSJkJpwjyt5ALwceBvCTOOXD0wcY0mI2G7
AUkHijI8TknEbJnWCWsi+4CDLiUjoFXwPDsdgedeq3TfR39RTBA/mpCAgvT8MA7D
KJgmFoQPCur0lhpw63hwtExAr4rOtCSf/0f7m/Q2lKl7aItbuqG1Mf9Mkr7xT/w3
LWzoBvP8UMNHda6nv69u8zsZh/lJoXJMwczlaVFedzjc864jt1CM6ynIDMu2JsEu
NEcM0aURgEmlPNHjFzQ3OknLihACeRYtFeuM178hczY8qoBGecFdRni+K79Zw8/F
c48K40iLgQAfLvxIggUqUXHDMv5YnTWW9HCtLQMsO0qvh9+iHCIFIrQu3+iBtOfd
DYMAmJpMrK9RA7B/MtTQGTxvDul6zQvFX5nH2UyzDw2kkLdGfj7BAaLhbr7JeKPb
T+TClMZSdMKRWiQY7+458gxdBO/iASkEI2zsynZPhuGMcQvRS9rs+9rsv9Uc9L48
e3x3UNzgR7aB290Oj9jiQLOiAZrR83B6JQXDZJaViJnpw8UaQpXggLfkexWHpNNg
ZBUIVM7q3al7uvj8Yzf9/D5hHhTA/ylCAcHSwj0pg9t56S9jXNdEcFpgpQAjtVzm
bzIlV6NkQzCGxggJ4CHygRoCoYsacw4JTrslNUjbna99B1UJP+oTGnPj32kmmonC
rJQegOtGG6G9oTslrKkLolcLMhDsKkZ4vNAALLYODPrL0bcvjUYkvYWzUSJxNOsc
HKIJ9YTou+ub8wKD6/weeDwEGxfX4+NotEWozY5HmzR5Er+LpYu7armZox5ck+xS
LvV4biOS1+fBJ2237vWwlIZbq3wFFkSw4cKsc3yEmCsYjnbPsku+6BoTrZD3q6PH
d1HtxQ7DZYd1SgAQoNT9smZhNULiR5r/SgFBa45LsrIZYTi9Mu0zOk9AVxdXUZ/G
pQPPAYPHco4JX5cImmTozIiHeWTraKn351+jtWlJP8MS0mfQaAjzkEfclKRwayQN
iL0f4kBzoMs/h7idE3b4Usp0ERvEb8GlMAQSG+5Lnqb2adpDN6ZyX1Wv9pb7R4Ri
aFtbTBg6m/SrcQqQoWmaGI04Tmnz5Hco1QvBpzziY5oHdChnknkUIXrTmwrox5YX
iwL47NRE9JMRj1dtPmtxPLJUopi8VxxKKiPT6MlNWLFbdZGeqLigaFpny+vp+6bp
mTwEd8mIwTlewnvNIg31Y3dO9vNpkP8yEqYaG8McpW92XHs7XlyNzzPmWicy7pah
l3klQ113UaJt65NRtJFuKa/i/hz3XGRra0DqsfNamfEk8wGnoOc/BLNeOosgS9Tq
RtWnoP5f68LVeyg47fYnYoO4X8ucnRBhF5afOhT13sEILTpYZ+xM8jqKGRHPPM+a
696/Z0kcCWRTqj82+psjSKVUA8fJib+TtjU6TemkcbEI3T4YkkCPKLeJ7yRi7Ml6
y1HqmAgFtwHD+mMTHqpVYlXkrkIJWbpPOveiN4Gy46VNuWRs4NFmqORyc8Vh5YwD
iMYilI1dM/zOP15yacUZ1McKIBLKToHto6DNZSJRDLko40Bjd73G6tBu3tNOyOYQ
BgTt4MjqH5V0K0ZM5AhVrovwE8BEYDe7WeBFmK097LAtNdhL2Ip8P/ZaeSXMbB9o
1d8Xgzo0qzhV2m6I2miKhLuY44583l1SEuvMkzneidTuWhba4DMHKrJ4k+dCzSJ1
MjCgv0AV/H+lP4TVqJwxnoWpg1Utu3dsqM9vX3VlG0pq6p1A2vYyh3CUvK1Fi0Xr
ISW4iTx+uk4Zz8w5BDYZGol/JORYBIKJWW/jCEycRzGeA5mQeX1/WnvlsW0vXjh3
FSjA2UX74dp5uMylkz4IiNiLBBsKJiGpkOOeVKq2JhlV92/+FvdWk+uWA4v+OnJv
ylSx94fNkgFHooFC/DHDGhNnI+M8TS6eVUYDrkdSh0TsqRj7JnAz9y+/4ko9oKgK
kRgsZQ8A0D4Q76k83qLJ8Ka33AN2HbAiPBVWHK3ubih63HEVXMM0BFydrIWJmJb7
+XJuaFxndgwnQRlTnkcqGqtvY8APd0I7Kp2rLsTVpNu3/4VYByrv5ETxWtqfkNRj
C1d7O4XuPa+62pxrf9DmT5llkoCBJI5gruSusE1ZncIW1cWkXXr7w8+qZAelbCeP
eTaoKMd92YJGv+RAFvO/jngooeKFhsXjPdmU9HWKdNZMlvluzJa8iSxxkCb9s0Z1
0rH68YZOSGYrx56phT6iN+qj4ZTYkDZbsjdgHckS7wiKTlTqV+k7ZYN5ooJfrWOF
QckCzUO0zZa3UV80gEKhCqO7RqEB2k6yFSdSGskkvvZe7Pr10uH+ME52GeaN9v2p
c+yhpcZ++Klkj3Y+F4WLVsjtvsJsCPICPoSH0ySB4qX7uYm7J7e5YX7Av0xE7Jt8
TE3sW1Jw2OyxnFFgGeOTti8U+U0GoSEz1PkmP/xhzlw5/UVsssnWpFCCT/7tFR5p
SM9csh1kvZSVJED9boKi0pdO3FxqO4YMFuwIbzfTH3ZcL6iyBXfLBf5tsSOLJ+/4
POcddKzLt6K+Ho+zEiGKnuQWfmRwbh+GXO4SziuDKwmY1DAo8DmRKQlU4yo7KvjH
Ni1Hk7D0Lnm1lLBYx3erBnB3mr3jJJIDF+7qdmMxQlxb/hZbLZ4Iiz6VNzvBAx1U
wTR0P1f4yU3DpICvrEdzyRO5qRQ3t3SGIgLuGITDDwYWJmq6a5i3DgNRqns1OVDK
hiNskjiFfsO34JFRixnoEKC9hG0r/i3ki0EpjuNLgA6+apju8d/Cw13DuSN8S6DO
7Yly3oNftdJm+IItmcRJuUPgYkViZDXJWiLjhPad9s4bvU1n0M9UVxXnyasu+bCZ
e48s6CAAMmTFAJCkA42E8o1DmFiaZXbfERPon1xnY/JzUzsFyQRSuTmsMzVjm26y
14KKgkAyLWrBE/hb8JtgglsPJXBdcIXH5AqtWdIwX03k7KZiq1G/FDgsKSjljvJ+
qgS0YRFLl1coGcP95Jc8TJ6vNS86LInImtOb3KULXe1uW3gWidCOdpyjrFKxJr9E
0Kc2gyPtqC6DqvyR5RO+Q7TbiPxInee9LQZxe5Y2O7y5PzxEEEg9VFa+PpOWiLp3
YcjWoN8QKNr7ZuCSuoLOjQjcYM65lTKnDx5AVwbtjojiN84Lm+GEcuOZNUO+ZBbx
QPOZctQCUQjcmJFZZ9FV4DnLaTkSDZzCUhca7B87X99gxx7NIl9hTO5GUZXVPLQl
BA9h1gELqt9ct2jYogFktiNm1NhZmQ1f5SCZe8pHX176CimYzt+lvvOmVyZmUdwU
LPqjsexNj3Yjq50WEoE6IGm7v65GSX+kr/UQvuYqlShu3z6Y/bekUCCeYHMb7BFc
46GELS/vsW7Ap8Bt2yVdZPghmYS4D6IYNpphjKJpVOT4o1SFp3RxFU8heIgJ9sWk
P5H5zykC1IyyPO0kgR3OhfJ2I1mhDHHerqtF6zK0uKcIMaQr+CaKjdFTjBrvUWYG
2ebHvos3WL7UlHL8xUJVV8MQmyjCrTQ+lW1nBUY7sC7rdpSWgjs+Z3Ecnjxbp8gM
qUqIXsBMgs/Jz6OQQHULNL5INbrI3DXyjTXrmVJdIi0sMhO3G5z6W0Yw4GsBf6xH
dsSYyfKU1IqI9i0V8Mz9X+FwgJDSKFHvnU8TCvY/tiBCUsKYUDFjglSUIJE5tgef
Vcg+WaEpoNVksXVCymgAA5dQLn6eDf9wEB/vwIR2LibNm7PfRqLBTf65PLDlcq7U
t624RqDXqsa7XCicMJdWPYXssKCp1cacAUe1fRSxMKMAJeesCtau+6ncabzxCnJ0
Ib2ZEIhoWWyR1NCjjWY7jJQkH1s0PwMnkmrF/zRArNS3imiJcQUCRa/bQdJ2gN86
9zCxfvsl5T98j8cmLituIK29O4/dnSjzu+DJLTspePlAOe0DrAfDrtZmTqCvqdKA
IPHtnXTqI3N7HjlNU1knjcsWPltGXRMNkxnSBZTBif3LpQ49p/HiMQ/hVCHIRFJI
zNQ3Zawntf3AaKRJT3mFwh5ck7l2EY2ThOHjGYw1sJuVx1CRKIgA1L1TgY8EWVn4
cqQIe/Uh50V/0g+NVhC+hZ/S+EkChwrwv6ZZWlVJ47NG7LpbGukZVWLppjh9DB8W
P3VymqdNYyUXgBczsTmGyLKuKCqx0raaXVxqPPXsQH5taMCdf4o0OmXLihST7N+o
vnNUswHp2e6sst6agw5agehjW/6BIkIf2sdN68kk7A8wIoHSi6OpVo3nuEgrjuBg
i3QlvbWqF21XplRVG/uvqK+3aDcT48HBnxlUR+A0cAfRdClUUixDK6mT7HDLmrhc
OGwquNiEpQ19C83ZgNgkGi6dHOdf46ILIyeiKh6jDZtitJVtsT32g9jlUo1O27Wq
ojhBL1E8ejObqW4PhnQibrO1/t5/1kMcwnNTvDw0gbbKU9R5WurYNS5tUbTR4RSQ
9ZZrLYPrCZi5VsG9MtwXPASk0UUthw0p+xIdFP0h26DzF+G7diw1fSfJmjS4XuYt
FLomfcO9sUi25A2Xs84LOs2Oae9FEkMGm87dzt9RJQ1sCr0nH5XvhRGAAswbU4gl
7rwrtFUJkzh1dJlKgw78N3wfegPHF5qAswE4yQhtOJfwbzQihQnLwiRTymuz24VB
41JnAI1McGszr0s5+VAxbIzOFJOdLjQYQE47/QIcxg4QY9lIIpz7zMeKgQSgS7aY
3X6GIo4uhIC69aiH2YLdZ4ZYHrgoBBPDqZ56YR0Ud5oy5bDy2ORYzb9ruC/NaplW
tzjMtrkqCHIyEA9Vws1IleEscD7+bRlasYcAo6sjZu3WNKfLYmOpe1RElXj6vPhO
P4tsZz50zUMfRHX9WotmqtetEClozHhVT4kY7b8gRtGQV9Cf6xOfemGiFr5edLrZ
ZVYYhQLrPpmKTSjYiPYrg2tHXnqLm0IxwjlVPQ/2j1yMS6ltpuJZSw6/auAnVkXH
SAVxoCd4y1IeblYLKJzvxUPQ8x/CdTSxIb40XchRSXRN5ebHX/vXX4YjSova3At5
QVMgpB7Gf38AFM4Mo/eSs6TXNHiztDXkHrfZcAab1UBTlhGxT2eQDJ/qojBbZT/5
aLuFDV25v6Bmv2vh3nkHDMF7G95GMtcWGT7BufG4cyNvV3fd/QwfCHAVCJ1zO4I2
CEcPXqbOjSh5McE6Mg+V/njtRLAzW2Sdra4CLj2k2Sgf1+4x1u7zMobmjVTRU4rw
MIVInwf1cL2FQzk/JTZ+esHOSdDY14M5Cg9jRjpU08Mn2NXCDLcT/NyCwKdOkpNl
K1Q08FspUaNqajJ1ezHvRGFEfEJUYs5ZCt5MDqh7chu4ZXHN1quy4HAh+6yU1/wG
+kdRVwd4kcl1eRpj4reOEuX2BU2+AYT5dZ6i4bx1DQ2gsnAsgTYNbbendkwEg9G7
8LZKc1dtGNfUxTdp8FeXclzBottHZk/MEZW/+wnEQuD+oo7amZAu/lp5ow0ct+Kq
UMW7MzSA9YEd0bzEypHTemBh2P+ssip8MPVH1D/I1biYNXwSa89CSWwDNAYLMQLf
RdcuKjUZwGvd4nWgyzGD/7Llasgjyd8eGO6Q3Po32Xtg3UPGij4yXIEYp45I6W+L
d2T2VR/oGdFYzNcZMPZ3xRtRtD+mLat9GBKdhzuaFJBPRf/9fKpu9DeTz/Jin86x
nwuqk6CkmDdO1Hzquk0q6jnLf2a2lf14GAJOsTzVQFUfiQi+HHBuUCL61dIyGrJ3
fofXH177ZVIHjH53fnl5jLyWo/9sYf2vLOgfV5ZLE4gP3j9p+K/u/1RMoRGF9N9E
fsIFczren7oTKqBwSyJF7OPhXtOyVymcXKOKeFo6K1M74iygB9/Gmnl8y5OIlIvA
ms+Lbn/Lf3o9os7D7CWyyVIKm8Y0jyJTJxFeCUusoX3eDyxe5y2YfpbXiHqAQFgn
i/2rrjawcrcUBfs2Ybmm6GkjBUy0l8eCkku4pSLLWKEKKpE7D0yW1rj2j4iNPxdh
Ir6JF48qjzaGwDk+NTm1f6qXfTUWUrEktsFRh9BlIhScoTbRMjItJl3fAMifc3WD
43fG3GeyocytT0GJfjPAFDXeUHymgqBiUA0K0ttXSmoHGIytvW33AVV5sNGk124H
aNXmonHidIIkw2kTkpGJxqkIaKYXuWzGKU2Joo5E1lwC6LZFJV2i4BDYo3VVex8M
N7Am1J3Omw/uJJ2dfSpfJYLQ0/NwZtlt+8dlc8us1c/2wZDrcJVo6EerhwkezQuM
0hz7LE0GVuqLrTUoP2vUAXySe9zlGpV+TcZXWFdqpODM2ILgwShKBjWZXtEPB6lL
nFnF4G7cCSHdvHd4gH3xmDD8yD+eVenkqSkuEncnN5jdt5cGgYXLt+Oxf53hfeCI
xOMItmB13q9Ho3vuJhiBub++LeoAoyU/WgFttEtTdlz4PVLIO8K6rQFyfAU4EEDv
9vC9S0rOpSHqD6mcjdATTgT+/iUKK01/zW2aobvfj5eZmtyB75qD8BT2Jn/hsZnQ
I5CeYpZuuj0gOSOS2Q1XRYzwZPgWWyiJQ6CuVC8B47Ud2lUHGjGGpy19hFYO7+nR
auXguqEoG7iSWOPPp//XG5xvCPVrU4STR63Xj5L96Da5QK+NlDiS7XJu5ydYRujm
+dupHBxHnuhMk0NiUjI7E/+8QSbEaLue8HLxnw+vca8ecsmYL/ATqEbA0H/on4wQ
Rs06rnultPkGkd22vvxC5r+TlhE0U1vN8LAz0uxP591Q6ukDRVaD71g73PyKubxs
NRH4unppz8y4aJyW/6B4psX0RHuFPWCYnLFrzuChnO6FyWRh/tfYgaxiRqklG4Bj
x9xJdI0WG7gjtsuF9wyc2R6VFr6VSLB8NLGqMbd+utM4UIjmfcxYBMKn/PoDDtCa
obettSO68kNZTWXg0JLgTMfAsqGTsllIwZs1SAHrJiXCBPi7drTvDosx8SWurugJ
yf/jhET8bo1IL5lUneSeZMwlQl6pdmn3ZxpIXaIJ3J2CjEZSpvmH3EjF4jYaoySL
R2BGfNQmNO7UcGcStevhOekFdAGrCFIMC7b4F+ILUc72QiV2FVQC9zOLiKqDk6JK
EcaIKfiyFfdG1SdcR1paxj2PMb7R4ZV6XEOqb7frcwIcg/PHfzwIqjMe12cvSikU
vHnLqJ4LUU6vDbhgJpAsa2CBFV5WaH2vkakQUV2lkI8mVCL6eGI05I8wQdW7fUig
btfkUphs5O3IPBvtwMoRuuQ4xrsrzLOMLUF5q6thiM+YVcCjL4UhsvGalL0mLS6y
Fwr/PYDq+v1TxqHEsqM7bbhA53AI6TDCQ2UMZ8+e/OynJdPYswWtCDu15G8KBtfT
rKwwM42MTezhz59WV7G2RY8AQ8diU4hmw8prBZO/76Je1BZLVq2n2dFxX9BjvfET
c2mMQX2qP67oKObzGQGMS52GG+AxD8W3vWwB8tZBlD9jzF6bjrMteOW4ZeMLRxV7
9ukEDiFdTSSHAcBrl6/sptf67i49zbkFQLJHsvMw2ZWOT0EUf9oO4Ijhx4K+Q6l0
5wiLtDSefq8S/CHN4iBnaxrMoqb7a4RtKKvpK7kPZHDCXUTaKGR0Vn1Ps2H2wyar
yfCi0GuWpfwFg3xnytltgXFx7X9MbfnhKo/48KDunXpyNF/FFCeRQBwnE/OoG277
A920qKit4ibqB3B83oHB75Prglp3Wo+6OineD51ZpNpxfu5zEetwCQZrrlMl+heN
RFK5Gq3PA1u874+kOQ/6HlJka3u7DtgDARL5tVm/gjnVa6zh2cUkkvoL06qzNnMx
DsiCsRVunbR2GIDgODl/RWQvRaemW7UyZsS8g6MXbcxFSvgss455E+jaRMgHc8Ud
QwICKeeqs2+3hng3xk0qSz2A1aHcKcXqYlTQpZcU2+HKbF8clW15alPrYrTCxEaB
SWMWRzItb+5O8wmid0CZqqVbF9R5h38khjsXOzZFS0aP92JVanssEzY779WxhtNx
M/QjD2yvtCYLV/BwYqe/TWs260aZ+6oZ1CmTLIZwQcAkXz/9bHtWQp75cTX/gZ6U
EjmJmyjPEOHolR4kNXG7cCzr7XxwO7pkxHcs06zZ4oKC0k3v6zxR5gmq2BEKQmby
MroFOz5kkDaI+ZLoTPiMx3TTvMHeOgjXqJF0lmbL7e1/BCVmM7qMj3QePVtxn+Jd
KmalUGSwQI504+ESAjXUokeji6wxdHJjyTS72PVfDncy198a/krFaoJQLrhzn1XL
hK6/zYTxU8FCCZa52iYKSV+Iq6VnWC4dvxddAKvbXuo62aJwKgv0xQOmC4wIMMWF
oeF6IVpAyHBZO650yCMoBP6ajNBAHdaNSDF/EEsZmb7rwM9rcOtJFuUOAdfrrfVJ
Zf5M9CJ8QwgfSlP+tGjou8b92/+d38nft4kAY3CaTa1a41t60TIsgkk+oD42gWDh
XowfCUBTcTd/tyx7qaaDMYqqDu38aWLRwUYNsW/i3cO7F+Zgu+K+EF+0mGjHyhXF
vTKDH8gAtCcYmpEyUHyNhS0zfwUS6dPfDx0JvSjuEDkQrR9W1gUWDDS9G27DAj9T
tvYH7X64Jc6dCAM9tX1073fdfE3izx6Rtr8cGhkfJuErhYbZvrGwj47xwL7rFOiD
xYoQ27yPgEtHDsoOJpYl7Mc9GtIQv8jQTCiUWzrnL6hxvc5uOMwcZ8grOd7t+9pT
OwldzuE5C3kjufNsotMDJYZ7pNERf5UKWk+UjEFy8hh4IWzzp/dSnn+BQklwU+Gi
Dsd6m2Pe4WZXEPACD8u4uuIkUfFrCupjQruy3F/eCUIJ+GsOtmJRbt1KdP0Jo9Ri
O8hQ763KkEP8VCzcBXnS0Nr+uLW+UCyzBRigrCo7EN/vg43enECJqCx/KcAqL1ia
rAAIoCPsKy+enZrTqAX1NwEU+PNqGjYZCFWkQy3aImZrh+3vpTHMz3tGYMDKoomi
Dqne7U0Iir6yZfO2Bbj5plp6hjHnq4VxjCK5NzxMQ32Se4VKSsnCPnYObEqD7KTc
bu59O4Lqw3NUEVMn+3uZRLXubdhkHEIdu5AJ0LZVPjLBrZFbqV2Ar406GCHFeFe6
16hXqWWpcYQ3tpftUydgu78xZmBeBjIHK/nQFxDCf0EdiNOih2nbYtrslUhB8/82
UQa7bzLlBif181VfZh2idthBEq+lNj0M7I++uHCS6w+BQeYOzQR/L9Tb7gYQx03n
tV/+YxjuK6o4N6/u4k8MnENUgXyb3o0/xbY1susdr0Nj34bm8XTkrJq50/FjLK+x
//rtuLilQMj9i0GHpoYbdt46RxqOtD+tyfUz20EDh7CGnX4I10/kW1U5LUIwkPpV
4CjSyYInOQbv06kXoU39T33dMoWOXo2OgwMnTbYFNkwn+DrNLFSyCUd9jLocQ4+7
wzNL0fWnfWn+H/RB0spXyNmC6eG2npwBhfoZTmJ+WPi/ZTpa+6HcuS8CXsc/BJQJ
6iTjqTyCzduOxANuiHsD0tJxum6eqmMgOg6e5AIksoKiMAJq/KIiFbLA+7SOT/v1
vCkIUce4ljq9s6Y1WQ1rcvtNdntQ0NQz3fZ+f0dstybbSqNd9O/3AhJpUmFth5PJ
NKVEXmoL1UrPExMa7KJGkil68kFG3HKqU1lfG3bqQFxEV81y4ezyGrUSZBLmfOsC
qhTCmxKIFU/NMH+5bFp1ScHf2SSazKkNXLDpErdaCw4IK9fwQxyj1g68PqpTzvDq
B7rK9J4qoEgtccleoVfYxas6kXd0V97YXalZIVaXnLZLDbhQrQcKz++YNiDTK9Xp
BM0f2aR5iehD3arZVGETbabDu5/Z871A9uHV1slI7W/2+j8CvqqTQSNlK8fguycf
he0bG+IDP88whBYvwp6aQcH3f+t2GNY72DquXYOHHGOocENiaw8ukVz7YMQn+l2+
cohywMA+UzdTgWjCTlyN3+pCUMPmD60ko0Tsb2ibZA5ZzS8JsCKqQdo1pXf49Qvq
Qmyi3xxCJMYa+eWItMQa/qEaZAjrrBI2q9HNuZUZpvFxFGa1sCkbNeeQ9ixgFQrn
kyH3EX5K85LBT+i+jqCbZFCrjzUamIKusnH9LR901UMcnZgRVmNnBJCIFJXzxlCr
bb4jqZ3ly6FcnDLRGEi+kkNaJk0am9v3xNr2r9cZVnR9YmJO9WGWGkhKpmh3UM4L
9h/pAoGHgSaib52ze8rTWwkgOghTKtTaxtChSzmUzlJ8KgEfhwE4rMvSs4rVP37s
Qwe+VztkCapamtv0YESwRDv/gPeft8igroXw8HsUDF14ulxVmlXVonUV9ICsGwSY
7xqsfBdmPQwDzaXr9gMU7ztoUo1spdVi8KpgRfnSMzJK44UwFAIFxUHPZIyN2t7b
TdkdlwT0tPwgqFITeDsEAGBSnn6SLw2HxN1pukvtK/J9m3L8r8B0bTPZa1LFSw2a
4TwOUYdmLSn2Lpveo2jgFjo7ddfum8kBKt7M+feawzNC37Fdt5az2jixElN9I+uV
Wd7jn8jW8j8R6bDGFGXMhVSrec2sSrcOmAXFU7dp2G7/3U7aIMH/fLyr429fzyal
aMiBzkLLb5Rj4l8B2PjpPishFP8qA/e/sQLd9/8c24VgZ5dNX79Cbf3Nyup4xK4L
Goq0JscI/o/2RgrUOc40i2Gq4GvtwltwBiLeO+Orj3zj96nV8e5f/ywqU/A6BxFy
pAnRFAoqctVir/8l4nMupbnF7+r9LDRSqaQTW3Mr6+wkRKmPdTKXc9rSXCAWmQ6Q
roV72b566msvXhsQxfG5GvpxbkVIusNI4ApaWveGdCad5QLwuXSFkC9kyF9kXleM
whqvXkNkforViXXOyZuTlTGUHZo5+48vIMM0kFA5VkqRua9AmiBo6h3ulih2GJdH
WRL8AOJIfjQH1573yM5myrHdQ6Q9XWY/eoJMqVOuRmmg3quRwDSMaGsZ1DvpacDD
GyAbXXSp91mI2w6vD9N4se7XNPONu5DZV0/TWd/vAKbrRnxwgpur8yNDcsVp15+b
9B48Uw2nylJXkCJLimfMN3Hk6Fvb1mw3cL5x9BTKgYmTx5QoSACwBfB54FzDaaW6
G9N71YPV2qpJCUdy9/WJ1rWr7Nn71A3Ynxvgc3OUOiR/R8kylqw6bYmXDs3RgGf5
KoHpyK9tWnJv2cRy4JNFd8GcB+nwqt+agIvoJXMj5L7dyGG5oW81c12Q5kyyDWhk
CE7N7rlxOAmBcaqfIPFPrtI6tXJjSXY+cywgQiTiLpEjWvnG6z1hUa3l5TtV/0iZ
SFCc+EXq3CDS7UdLVZknZPXKvqQ5tQsodksVGJzEBfdHxrwQR7NI100k9RbVd4PJ
OgluHLlUcQrkcERgvEki38luxm2GrlpjtfrtscvY44KLkpvkHz00XLKvwPXjd7Dw
mOTyris4WOZJnFVos8JB7BUiH0r8NahSPLM0d8rGRd69v689nxXlre4vcTqzyuiW
Iu+X3iyaxtIBpxl74NwOgahsZqKupBfNSNdUAAhi+yFlzk9lzOYpyGXheKoRNvWw
v9F9z/zWjuO9FmZI/qNUV/AwVgNRMXXoZhGPKQQbpDrE64+nP1mMbO0h3DerYZZg
LSUldy7i6jEbqdMNlfzp/R7IKHBCnkllMpWHbGainLm3GQWnWPMqd5STxUYel+9W
6Tz1hhSGlBXsmUzve3VUE+DCFB3/Vw1DWUDGIjSjbibiJ9Luv2HBa1BTUlq+5/VQ
bIOqtvEks1u6OdtT78ZbC330wfdXQ8CLMFpUM+/5C60u7t7CINI6R5QEe+SJDxuC
nXoj+en8h6ULUrE5wwsiYSzPVmJOvWFssl4brhFGhTOHRRBv8PNFIKMr1zIVDIhy
fIbmXotyifiFkzwerbN1LBWtmMlCIpmsORFhpr65IEpp6nht62/4Iq60TMdZzrO1
r0ta88ZT2R3MMzFl8pgBmoTKl5+UfTYAL1vqa/44G1dYMwUvDD6cahHr+CSHKCv5
egZvs42ipD+DdDCKSNU5hdfQ/GMUeRRjVfs963JrmW+sgrjSh5iXThz0TRpw//cf
TK7bFa3yephO13EmNiYd2gvYx5fVIYI6RW59yESF85R/+7huYpXWNkwshxtAr9zF
SjAt9ZtUkm0Sf7gdcQBv9A0vlIAmCXwYFAnr2I06SxOEZphNJm6FMhGkYW7DmikU
iN3zYbLhGWDJ4ZkO3hs7F14weDU9g1T9T82oTktb99eOiM4Sj4plnHFhihKVFaJa
o0m23pH9OOfwZITCJ2t9+lWumitG9KFq44KVQiVXvV8xkuPeKLAcP1kYMXMT+FYI
XzZ0JnKSqHS5WZTB2jEEYoddknm8AHsf3fNULi/Zh7yIasESigvrj1iAtdhD8ETV
EsJacoSwvw3bo02Y7locncZnbeObuNbS3PZ5ACU/Ozfxh6mXEy/F0lnRxs6UKzfU
c/R8m0Oq/b/ytp4xYmrangOqk7HtoCt1yF9d+M1B4l3A7LHMIFWLWe/zzccYQIb8
1s7lgoNQvzJ3eRCQnAzxTkygO6d+fnghKxCMzTaD9UXG0CO6lDSd+kNtqgEtgToD
ddFJS6+jozU/5iBDx5zO6MVAPU3a1l41cmi3HBg5vk2hSnLD4T5Ghd0csNxRSGNF
eYNRAbn6NNY9Q96lEdDsBPtvWruDX23mhjGT9wO8GwYKKrjICWcwbh7enLDZYSJP
/J0l6ZC9KNUV/3phh8j9peo9Gv1VSZUPJ4vRT+L3w/uKWq7f+qAV42jd71C44MnS
uO/EnhCkaDMZLY/dIFnJDLbmgBHKiZxOynAX/S3nc1zb9r7NECno9yHsvkXoZ+Z6
PlyF8Ppz0I2wsCW8HafrEVoqa3AynYiZGjxY+qOrd/nzyTLHA+V0iNEuHDSTtfu2
ZAfdmvcrivVswuLCRN5jicxsHoJT2DBR5pesBLezOPM0K8o0afpX5O0l8QMV21ws
ABvfiQFO2IT+NcC+F0zF+fqznvDmO1d+/aYtNWTdgl7SNjgPswWMapKOybNVjNG4
fP2CKVePnVY6umTy9OICJmIX+7kAbwz6LhiID/uxA7zB+ELa0OnjLWsmQsRTamu8
dlo9yPoRY/H7EIsPS0eGgIw/EGE+hcih0gzJ3JEvfXiUkaEtYRSxnqvcOM2NVbfm
sQsRUpHM+4vW/i1RC5JK56kzquDvGTv7puxpNa822FaPe/rUErCWc6bkTLK4Q4Vi
JBzelGOfVlYzhEtPS0BW6YqQA4Qx9TA6f6FQj4swOAYH6PpTSz9HwJyLKMHzj0qQ
ASHeNEQ/x1B9BTUbnnFqggPoYiQDDjmILTsS+FvA74iJNX+YOEqoKxyC356GXYyU
95KE4fdNjlW0ldTJVYBNw8mXySpyQWM4ZXUCXVWpL7cxBOCZ7BlWGd91JVuppX55
Mq31oIV2cw4ix3hqXw0DtieFfcVAfGugXNBuyVBTlbILbPAWHudnLCrC7Dh4I7OP
I58l0MJajU38aOQpWWq33oaUFzHlTM7wgzNMTsIIAt8ifdwtMY36v58SwGrEIcQQ
Mb7/l4WDW7yiYvZMUHBemm9Dzt8jkuyWaVO6tQIyRATZuUz8aUozf+k9iLvDVm/g
cdgjh3z9qLBJjz0Efp2vH6HgfGZyOtYFNsaarmUoSF0G88nSHdi5rWR+gdssbj9Z
4HPFYyqPFqMtYpa065nfApsMoxhC5gB02oV1NuEukoXfD0nCF8Nenun+u+bCLStc
ndivlZIF30QmUYjtf7HxRlHEjkP7KueJXcYAPpsZmjGWHjMcMHbCPxinBur1DLpv
R3ImxzMHCiXYMSZx0D8Dm9QS2FCIU6KWPjqrToCtFhk2wuz/2USgBwAIU6JK12EX
+8+ns8SeSLQ4OtA53fsvIjXuuZJ++MnGMLbeUa8vtvPFFLlTNgNroyJT8dcc0f6X
e24s0dUUBCozwgB+KtYdASGaPptfP+1Dz4Y+A1H4L+sv5r40FX5dAKSQG1jX/oWs
Z+MBS+iFrb9fkRCdPCQV7buP+eQjfih7swPQsItGNcBxEHNJlHXMUGT7PU9XviwP
r+DaAxVLtIes+ZCJO3Vtit49B61uzFFHaVsCeBx2O0xwkFyP4D5QrAje3+j00BO2
5JtQZMNFgaY1aoTxa0xl/93x4IIzChTSBUwvyCuDJ8XE6g9xW7TgeDuSwj3RvcKQ
menCcQRkgCN11EaB3vwyp6CrIbBEsN5V5UK7mywaMAje57/1lD33vKXdzzdJYmP1
BA9SOKcbta/vAsC12XP5KnmlyyRQl99DshKRNeaG2DHBZQ5YeTITMcyC+59UxMTx
3+xSShSB/pW5ggEExOH89L24mSRqXWc52Eof8x9ilOCyDhCyaeWQTFDVfNXbdL8q
MVmMmvFung3k4gSsrpc/6bY3ayPIrmW4mAcUdWDAA9VL7F1b++P0nWe7Zkw2kJ60
DXjyY1r2W4GdWt9npBHco4YU+DgxPVFVeGDmO2vBqVLJgPM1v8Dwi0FoEENnP0kt
TRqDSAoOkXe40rlVcOB+k7unArluSeJKZdFUjeRRD/do366De+meKRgcVz2WclWo
Oa0XoyvFZAeN3wltpWZkYdITZfCcUwP0fYyrCsMyz34C0xXW2eF/v69MzCtgKk3r
K9FwukVg5heCfTNNkFaziCLV7h6HaPq1s+morTqJ58YGjmgojzW+4Bm9lA3LB5dQ
oUomQ1XorRLGF8HSr+AlnWddHyyCEyvLoLFrW29N7g3wiGzpq9AOyVsCxFfUDrri
UYYTOcQ1AVt8IbPSSnAR7EVWOwGlq8Xem32Q+n/aCWlToMO/ym6MmtXalTUufrhe
jM0AnyEw/eS+K3+A2kBbOf8t9YxR7F37IuAnh1r1oACuLUMoilcDgZMxGlTWvGEB
H70zjliYKNzvseZrQmdac4L55orWffdCnmWwYkS/L2zmPCZj+9omjcxObv2an1h5
WXXqajgBkVobndhADcIfHpbol4rl/lHw9MEYWpGSRBtQychq/FTJX8Mty+c0B1BW
oT0oC1JqQgZdmnM4E79+RFxotWFfTK+RMaIF5MbB6+hvGWonmlOWNr2c4rZB+nsc
g+LB0tanYoMF9y67xwomxn2xUaew2IMs+U9Saia4N4k0vSIzFS6MtLuok1UxyTiP
4Bkk0bnQ4PxF/DaWSNRiPaIKr72p5MALTXUUQF/Hde8NzMCxKfnGaqHJ/7ZD0ZCN
2HvxVNIyjLDdM+y+yCEsNelB/lffQ99E8XrXo3rrVOomjIPu7TJ4LEsR2zGGEGLR
aLbF/oSr3N8HMLE5n02AAlnKVSwbv+PGH/eAwsm+tLQsjuJo+hoOiGFRzbMJ2pob
RYj2u+vP8rNXvSRPOvwTVOXK6dkNBCZnvXUlvj2aV/wlHVb256H4cNuv0cD8RA8O
GX/AyQdc1sYt7s37Nfbcq0fsHE14RvfrGZVgKZ9ptGeTSCL0h/PPm6+NbEMuGWEh
GeDwAmbP9G0AB2xds08xhyyj8iEE5nAmTGb88fhe5nJMj35gIgwLYc9y8Uv+LGIe
J3pmCkwnbdfjTRVF3LcelE29RPEM4oZ5gex0+voqhj1Ziv2ez65Gp9EalcsTkheA
nbcDu585/IY9sG6rL/0SNVkU1NYFgxMzwtapVIgVk4b+nU6V7GbLBYuffym3AVE+
SNVx7zVC5IqH7TZMzLQK4clffyWloB+XRERcsWGblHx/lNddJoVdL3EAwlbR4xTD
qJt5rSWAOvuBDyA1SULnfGO8VvnzE2oSY/yxVN1EiD1+RaVYi1w2ATv5IKx/CktB
hc3myHYTZN380JKZTeYGDeDG/Ciu+k+5dhxuv8gDcK6CrarqU38sJATpdXEI6x5N
2MkzZv+Nd0LjFvJAb8asuBIHCybNofO9ZVJmhKB40kwjYd+g4pHbQ32iiz37p2Yk
wTccpaBqe0c64aKH8qLd9T+c61Kr78pjU8Q60CWreSolUrzNsgM0AMSBoyctbxFs
Yp4/H/26Anp1xx/SVdkxocFCeOszTCTH+qaCwrG2ec2vuFoN7X9JA46yn+KUHgbG
Inns0U7BHRuQWKoXbp7tvSSfytd9V7DOZK3DG8rA7VlwKiI7+5c9aPREjpnR5to4
8kPLUQuloUInGSwzjRKCkdRMbG8BqXvXXR7GXxIe3eqcVmAIY6VwdUWVAa3WdyOM
Za1zhQcCLO+Gsx8MHEsaoeKyPweuMmnwopcjTXEoN9womz7r6Dwp6vZ+Vgy+FsjN
7bLVIPFSj1Bd8bWWUOTK9maf2nWPQJWEq79kZTYkQp27OcraOiLXLrxvuu/gAfmE
ceQgYjAMy4Pn508rWDw3AxuYXqV+Oy5sB9mbmt//+cX2nX5Q7Wg0VdoG569v7Twb
Pc58cGHuqPrum3hUoIGJHDFIZpDtbe/UnBhAtTkxYOSJblh24i1f7cX1ZmshWA8Z
Q5XIS8f4Nta6veh9lyOm7QJk004YasTN3B9StU6HHcFkGyBk/zXuV9Wj8eQSEef2
OANQuPBmq7oC8TR3LJj4QQ3O6cPp7cWo/FP5+m3BhqgGWHR+ZRvonvJ5tZfMNgIE
GiVdFUty5RJHEtMzbtaNfhy4gFTUTv+A0iFFkIdiTgpzGuJ3+jgjfQOOIcwqviB+
Jy6+ZJ8vzaBV080FIR3+ODK4UJfFi3VjtnC9iWlSwijgEgvXK1WTZ9iYZeYauAAt
vCOZCzzkxp2xQ7JF0LKgzu0sB50aGthJwMOEj8etLWlkAlK8ygyZDp68wfrpTUrd
Oi0kDrloat38E9WcxyTCRWPQgKN9elxc5g3bNGUWE3khuK+0N1oVem29fvEeRr6J
PrCO7EfW/c9iv2PYw9fr70CDrjfbIkqk2xs3hxzEH+rsNAyDAGbVRkeYGYtq+4nn
v5Wya3HSYEAR5ha6fJb6doHoJObt0PUTLIV/jMoKXgXLYa8xWAi1n7Gg8AyFd/TD
WxFpC65ebIHDKalSFrs4UlXuAwRy+s4aJDSJv4FlZdwL9F37p0STitvCTLjeRG6e
MGr2jGzPdU3/ahE8+Li4rokiDW4DNWcR+/KCPdTAfWW6Nc/6s+cv6EELfU+bQeXQ
Za6LbXyxDr7qcZMG3plq0GnraIRYjeAFbbQG3ft1fvAs+0rs5l27e/GtlzcXYPnQ
x5FRIUX1fw0nET18l7V4MI8NffdKXWvvkuA9WH2fCXMsz1cO94dl78qiRsthOva9
RB1hwNdYVo4HOZWIZlpv4HeKqYA4eHvLWD87SoLs56pNgTfaZJChmUlB1J3NFwdC
xbDmUFbegV7Ti+27JwLAFYgNO+xrGybJVP7sdsmiSU1Pb6/J5RQE6XXn5ldgtF0b
5J4c1o3ELtVclVThg/0LI77Vz7JhQLXGWuO4SglWDlSng/Vxo6H9n92dE6NhWWms
iHQU8a3j1cGt0G+6Tolmi6EO3JYpfWjQ9qHVjCm8Pac4AyavjZ997mduRmsKhQ/A
81gTcc7mCdfCYHZFwArjeQfNy55IT+WlbP0sW3iEkzc6TQvZU4L7fUvM89ICICXF
y7TaBMOn22oVmtw+gGScvYEa05SOwblPTBPbtftT9mdt6woIKtCHFbHDlX14VJou
mkLqTug6BlH1XcIP8VcwuqGWyc18Kz21qER5Ur2rx0838SQeV9/9tsq34Zkd/aM2
o7PGmmfb3QqrfVYkRyj4iRmd5UYpUngo9EBBCPpmtB23J2dc8Hh6A6j+KMTyQ6Na
kWhZYrsMUSJEygKwHQ3/tx+XPzVZq3LhD3hGSTLUawRrNguvTRHtcEfLjQaBdPTa
pbctwH4+5xBzj9LaiXLOxbVE/ezK7MUnSvT8LotIwYGn2KnBTqttenF5FpkCf3IX
rBwQvUSUxkstjmnFDWblklSNucBHsFU3AN8jzh9HhaFGcnwcgAsuAZusUVIVfQsM
3DGEY/ystfBnryK8qRHHmplFo6ZsGz62PLjOjbazWGteeXw7VAneUNH41y6Yg88E
BFJ5FR4ohXZL/P6NGlY2axc9BhY3bE+aAR4Mr7wq87+TrnsdQW8w/M8rGjFlnaeV
xQKoDiZhcfB29+gAyGpA+wKEHxhq6VC6BwyEk4jA9OynAD4AdO45+YC3zEj6TpzI
3szE5wrYJFoEYXOjI57Z8MidM0OawrC7YfRVHwkle8mXUnqufrTwJmEXbcEZcEO9
tVb4xZ9wXkZo0s+N2Pve7JEx6VM7cP67JNoan9bg8Eia5+LrBnuGYDR65YlIxQHR
R//pRjdctdY4Hmldo0aPNAWrmFSiXh2Bs4yOseVTX2hReHLlT1sDhnUQGACgqJPR
p7xWB/3qUkYZkdntpVocL8h5CuSPv5po3cceT4E+8y+r6W77y38jXqMhtHCyx+c5
ckRhfkGapFcRjBQlSagS1ma19cR5fMtGmEJdhs8QNwGpjUzm5eZCrHpObhf5bEyy
CIGrTDiQT8PjqFUOvMFBfJocRTAXZ6aOn9AnE/ORRQ9XL2RuJzs+Fzp/2FIMiB+/
MsE2eMR9HqKFI8rkG43r6AOKaqPG4TPhUrQU4atR3SVMXkwZqXws8lijmmm+fcNX
QggVASiE4R8nay8fgn47sZYZpwrpnHLAmC6lWmog8w0d+g7aTjAasckt5hsTwFop
l1lsTIOsenzx8FTbVausLDdsMAgqbeK2b1athblPoQK8xBQ2HGpIAtei4q4VIXNs
KXEl+LRJYB6dMf961FJM1mOw5XcZx2edwYHIC3ttTXGZKEZ1L8n/QaMZhDuCq/qq
k1dV7wQHKSsTUzVQVzf2tM9g4dN5PcpJa7zEURxzA8u0zCCpuhwzFu+buGswSI4w
zYcmKlnhNEdtLaFZSdbM17JhujngWmN6iogPV37aVoYSntNsQbKDMjQI3R0QRnaW
mqX9fBhOVFCjMv8dA3KUTmvlgxxdpucbK2CtbybZmsYPOY5Tt1F3Pb+ca91vEOaj
GsL9jS+t9CnkGVftcp1aKAzWMSiuLxV1Ouq54gnVEWSM8LNbozBMNL+84QDx0uUm
U4i8A+igvAoL11qLCZQeFhFYNN25nVhEWcJpmNvfWyIK9jFBypARAY/ogzXxi13L
Fm2g4C8levqo5IsWhb1VV7K2prgLmzHWto3pwtKarwpZ2MdMciJGXhDOTXIg3Y5Z
K+wJ02qc7+xmIR1zL8NNMS0ZXlR9AodOmTqxMaddn6M7L89p1ZfFaJsWRkBJeyJW
2BrL7rBOW8QvmyADSKTVQwS0hhdjdyJgypNB6wh2qLt+VhyyaATibPAwXVLJucTY
dXp8xYjabn0H3ef4AOnZrsM+Z0sSMi+e1gKt9c81tDf7eN1GKz/8z4BoOyqr3Iq7
hdI78b1CCDONUF1B9zM6c844zePZA5NO5BJFrZ9m7vElO9f6l2y9gjiGUS+ycN/Z
vM6RZLfOP+j5gdi4hTBoHbBwteyc6NKADEFwy2LAeK00R3/lHLzHuA1Fv4QCVHmS
EhU3Okewl7U1IrEdSDpX/1wIl9IOb42Wh24g9x0TilANVLCJ0h7b6onEuxw+shys
hw3jn9YcTvtMiFrJRgUq6ijgzaWbuyk/NvblICA+KM+fsa6lEI/nmF3kYVBl+Dlj
m2KjXbaG4eNWz9SmSx0ILzyB6ziWQz5th9Jkl3lZc5A1qzl4ZKNsQ/IQ6Zpjkd13
PIGWfBXA228joeOrn0CAer6upNaWVWQTuhKJzNCC0qPsjh6dNdJlHkN6jeTxkCqp
ebg05OpXA+cv276s99K9AzyoORMn+BS2PCltJA2QbIOjfMH8MA5LajSJ7nzdfYUV
gLhhrNecDmGAh+S1qmg89Sr1U4I7Tu02YOjRtNWX/GxnbojeDpQLoWdTk5l7xwtj
5jS5oExGheWuCMFhMKX+achbc+kBBtHnYqTguRAtm0V/Qb0WNkx3UeijCBEAKZWt
nX5tVBL/hdY/5DowI3WIzNequATdhrTWpaCbZyoUx8cqtuFb8hBb+A/LzCqxXUYO
mf9YKYB1OdjXp8/Znt+b+yf5VXA3ulnbf7gdrOJYSzltkBkIlWKpEqkYn7VTej7p
uLF2NoXZSGwjejLYrcFeBzUEpaLPvKfUkhv7Dbi+YBrfwL2J0chbGZ+K+9RXlWgV
RQEGTOmcUrllNMSa3UPoysH5xFFoPJ4SyQ9bwwwfr9x8EkG1Mekknbz6LF+dsckt
2nuC8XMfZL2C/ZZLLRs1BsmMj6cwCNRcvm/Oj8vHzz+ib1cAOSaOdTGKfDldGmBK
dPmUGfeIc4MzXGNDNlMsuJPacGd+L3DaAGnl7S+eMv+AXy3uD7xxsuxmPCUuLR70
1XHwiskTlsYCZ85ldYn3E9iUekiEUeMCg8nP1bXnXJ4ZQcwwgYQELk5ddh3NbLDP
JacCeCSC/tRYsPinHz+1Nxzcs1CjFrB58LpQ+5W1KBGaoPU/DOUtqJdmoUEFEkKB
m0WMcwSjZFU+D8wAF4jvCzAifMCQzWIQmEGYsFPUAbeWKHkSf0nksdFA2Whm77hF
00sv1qQB/9eMF2sQ/RW3eZOXb3FZKwNjVVGivAdixuzpuS4/VyoE1Foly8K6ln61
dzOok7ZYvlSA1ES95GU74pr6WReYjcRtbpudRVf4FOfuOv+DqyIcjUwcmMOO21BY
4Y5eSQu2AkOvO2bc69yoGtiIRJJ9YOsmvF8BBKaCu98crJknOy61vCVJSvDMmqHe
x+aAW6HZ4TaDz6T1v5yEa+47MjPopIiJIHGuCV3MTqcW2fVxoMlKUa+JNS4caYeq
LGbp45loOLX42SJhOdAKukt1JRfqUX9myQlNpD1lLv6utxq0qSNVUdLuYlI0plNM
k2mrYsmy1YINRN/5UA3iP6DP2n/YqhYcP4Jq+scrLDGfT5DoX0lY7xKwi3SIX3IZ
fIlKJTmhYIV8g6TR8QkGObdGNqUOYQqgfUj3qa9uuy2QSqJFyS073qlHv1SVEs+a
vxuYm3td/iNr0Fvrbb9c/qUXFukyF/UqJvtSKflm+eRQpW8KJMYE2UhKctavQMob
kwNSDWqapXfbQm408yoYdMA5o7NRkjiC5MjversmRDTpoF5HYyk58NuMMpdzvu9h
eTTqhIqb1ojFhq4G0Ku60P80OLRaDRlyVxOomvXUQuZmr03ML1vE2khZUkLAzLCo
UAekMZhR5Gt0WKYY8Geg/1gWOy5VIFqdhbx11WzQGHeWeZcUf8I4YPGsxLhm7hF9
NcK8jY30+TxJa/QWuCtRzdM7RURaenhGLQs9ZVlE1ZW13vc27rZrlTqzxicnH1AK
bvvTvKMebYZUj+RNZeMfZriR/ZSy7ElZOwR0HEjV/sI/RLor11TzrOB0wPiHlh73
GIp7xnV9xr/w14BwK2Rf3ij+er7Gds/BY/LtuX4OfWREzaTp4zRalU15vZcvxrAv
sY0arrCMu5LCXxm/54egV7kGoDXNPR+VD15Sxv8wcAhXljVWFySTRBEMhBBuFYCW
pK5bst0yZSJnnf1X18PfNDX88eizt44OmaZe2usbPBncQeLO49LqNIqIJgruyYLc
pkuvz2kXmm9z+iRado377LmcvEmhRwKGzHk4Qh+Gss6B7Bxk7L0HIqiC4jWFamuN
0YgTuffG3IOa6YTYITI2H0UNhISh+FjAg+Ro7HdoLRrJtaIqNXtHD4XuJvsni5pu
vmaZ/DfIg5zJn1wxR99xlmsUBrdpacf223MXvs50AiD3kDAlb9scFvQqgBSacs9B
7+/RzVLvbsP5BpL5cUdEO+bNT/DM5YnTlkogHMXpLUywQfCInwzbeXbnLunCW0lQ
9y3D6GQMa4dWNpfv0WzCNc9FJHfuD3fALHHyv1f7wcBR00/Y85x7kxRm6GRcqwJc
oTHDrskmg4NchZ0I39HkpNHaBIzBVc9gZv8RWPOC4bFili2LmzUL0vSeBhYfM4z3
hOzLc+1fcVJIhJZxsq++oS4zkE/os2SIowccTJMKjSWqX8/XpPUJ3GuyW/SpsT3u
8asHnl1EaDb7XWtxyeN+9cPkSJ9vJ5/Wg14B3R2wXndHGKEa4T+70jtCdBrgeA3w
WFgylULSd07bya/eaAXrf5ViYQlkNyp30pR9wpBDMo0cYYfs/3XPfVtW+DcHQj20
bRMQ+WYoKgoW3g0hMZPRAjh4Y9bPD4bkOmoPitbFulJb9tAhi8pPHay8zo/O5frG
dEg7hs/w1RAcFLJ16i4LnhqZaF/Ad6/kt0ZWkiXvtQIb4Vm5OO9bT5G8naUWLelM
iT5QCwjAqjPA2xCMqbFSWuGIowvNim53aFITF51vYXn3F8QDdwIhA87V2nlhrNfO
SEr1OJz2DNBEh1UgPL0kfyNRnr2YONWFvrABHpxvFrj6y/LZNPEQNwrDfBYTowo8
6vpcCj8tzuRRPsReGOWsL+X3e19N9uG17Un+ScoRc3AzWicFOgvj253FzjqD+eB/
8n+mroybh+spD91bsDLpK7MGAWXexRdq4ZA/yhgdOD6XLMav0woc1RrOYp4q8KqM
q8XclCd9V0BjLMgBIapeo15JqYwO+qNolsdNip8FGFqz/QKZJi05l/6Nq8wCR8KY
imNg9Yx7aIaH6K5AjJFxrMaXl4gn4aY05TUxOIetZHz4MQRI3Gp89niJEIU6RiV/
7x0Ej9/r6YhV67BeCfhkczNzWp7MNLRyhkQsbJ2+D7s63GpKj+adQaHtZ+xaputc
t200J2ytAFVAENkZSwUcC89pnjyuDpnfT9o8ka2Gs74F7SiQpdqB7v4sDy/9+OV9
tRj+yHtnCcdjlhgfm6SBAlSR/OD6l7yfcRKKvUu/czBi2oUZh4fZcE1r2T+JrQu9
uLD60/uMpeYooetQmxHZdyzPFKCBK57fcl20nq4RJSRAIQSVCNffYQlK27bwz59h
qSS9tcZjVPCwvDlgDBjRHGgqKCOglTUX9k6rl/vHh1guGtzNsRQeuyIWTK1J630O
pfGvyYL84uG/zYPqHoHCq9aLvSyo/uwBCOtW9nepkX51neUcpH84aTGLMC0TbZmW
mM2a8B5g6fyX8+QYsWwBG18LvrjMsvXaj3j2Ormo0bQmbSpY9IzuINncRxz//XlM
J6VUJIloHgIh8xS+lc/NfDzm+4mP2IS0Hdg2ROmmmZazRbzl0K/7mJ2mhAhjHkSj
Q7L4MiRqzGsKL/4PucWKRiE4k/zEkOxMb7nilC7z+TsOhfIl6EUtAz2mrAihvC+y
FZr0gP3/XJKmQiiXBnoRPmgH2WQ2FCPQhbn7xFIOxP78jQYCNvZTYgGcBk9uIbW8
aYFvnci4/GhqMEtsDuvKXbIPuHf3W22+chM3UeehPyZH9p5ZjvKwuMZeLadCjQHM
WJVD6S1cT1rJDTCUgbNGEEaCE44PFrSxIuM42BklyPkbLznZOG3RCamxKznN/wsO
D5S6/f1Xwy8nQkUIHttXRuXvaK73eaPVjeCp2CVx8lUvxj34b8R7h+S80qXrxGHb
US7mqPV8X7Z1K9eiFwyTAKUj0WHqyvOtKXJFOaFuQ0wJMLwyQ0fzu/qrVOwRJUIf
30ESjT31XgVU4mitGXkfAjjyGaRfpE/RMURGm5U+CK/SrdSzc4eJ3wCqu2Xo+aIp
4Z+Msfe+fU875BH4mQA4KrGY83D/mW/275qRehV9vjQ1DhUd+FBFFzZvUlKs7lJ2
rj0oqUkEW/u8yWqEH6jGXT2YpHWZ1wa6P7KMIshSD2VYA5ZjJiS6t0qYpe7nNmay
UwPHwYPQI1AeBlBMYXJx32Fl98nYQeveumyyeQxj8bFtPEqZrkRhwiQvBjxyw+Ge
sXKVDwRGbpAfTJctuWaflhJ5DEeAEDrDSIR1PZ+FGtrQfOP2X3Pz+icFkkB6fLGu
CX/iYC8CnwXWF8uD/c8YrMtKvOJXAZMepe30xDVWuCC6i3Q+MUPyzXzk2pgcEZ9J
bU11JdF9DuUoASTOa6zd9BJkUZxyWJL67wDcS7L9oYsfwsI+R/e4WjfCTllIqKF3
wKdAtIM+08Y2Jzb+F0jo/26xpeA5PmK6XiItLAOZEXtl640S3Oe13gXlBuXqu6xN
XabJLVqAROB+fpv0yTY8Ki86FoqqSStTPFy+C8eHaoNR1TvU6+7xbZNZZl9uO1Jb
yfJVEPVxEt1q9LUKHD07V1IZNrU/D3iHjHSlhPscIX5bpgo2LbZaiHmk3iEGrdKi
ZsY+WAcBU5puXvdTgPnqosirP5TlwrJkn+XAIL+BYziiN4IgfkEI43HLEbZQfQvK
1IVSvnl/pOAd8DUmhoZv3TLl94yTdO7MLGkrXuDyhKGONRSGvkTj7Rrw/IONwID5
MQQAS7wUG5v8ERHpuiBFej6WCfQtebL1zeG8yyntwdqa+fhf2M7vWhXHmFgrWNNM
OPdktFz8xShOLi5Mpb5fziM9mjtJKqIxBTZgAwiIyop2EaxmKGSD1l65B72FHIsG
YaX4DV/l+I2XUNAD5Y8qNNwu2I8B9uSilXLU5zW4lzLG4VF7AAKMOE/fjja+WpNx
JpmdbtJFjMf98MgN3w+ATPUIMmdwNaNb0PF+ZklBjh4FPNUj2HgjvcL3BBbIJge4
weLDu24aWr13ZlX/reXMZr3s+HgQ8ZM2P2YxLu7mde0oSN/y2nI0DGQ2B9XeUr8T
vSvZgcskRnuyhaOYQKQwwcBZUE1GsnxACaf51ueYOMXXyH8IidJFUe+emuGqeF1B
CSGjm1V8DO2hKAEO1TJeEc/wZdG+5GhR9YEtP+YFS6tN8I8WbhIPJz9LrntsbQeQ
LOPW4aHka6Wm/fuaGkUuBoEb/I0EjcheZTTydjlKNLfv6jBvnjJ1W8AWotu8RiMM
FPBOZLSwESRBzIwU8kYnjtBwMi7+TpFE/fYDhiVciEpuYgFZ6LAo/7e/kaSSOVWc
cTZQ733Hgz/I24bDGjlxLvAxhZ0yQhGiatshoGxulEUj/O+HLA6QIzcDYFb0vb8v
pYWzVR8eUX1GYKj6iMp78CXCJVoT7lJVFM+53BVPLpPcw7VOD8dYvuqt8lAnXB9X
KkXqIIcmM/gBgpDyD2RAEyO+HSoLBWkJH8BAV5cDgEpQU0aKZ/Zo+tbmCqoPFvHg
QwMFrBpv3v3pmOYAsJK8NQeAc7ljRZIR9PPd/9Df7y8vWsMfQqpQrXC4yiOuXWw0
qJqd0WkJguPDSsOqi5QORlbaFR2t4eaTtfxPfzvKkyBwIb61jqK8tA5I0PAnPgGa
A7DJ4s1LLK/3lHBHReT3h3S1sujw0UNfuRKmQg/OXrqy9YAK7Os/bVYqqaWdtWud
+9S0++6Su207me2Yd2vGDTEJd9ZUNRn9rQPqkgEpiGTAjIZXzYBZuOtNtFwrzup6
UgkLUidGyTJ0fnmq5iy/2c9s1Caya0iJVkr+o9kQ5UptVRlbqT1clXxnQ6otqYt7
gyxCQFT1VM9Tkx7eP6qmHGIYYDuywu2XzNTgmi+scIoHTleGtTVKN2Hnc1SN5OdR
WJjH1uzN7PWkZlK49nRR6M9Zwvo61TFi90iRUN/Hi8WGq1355EChjOgyVpC7dpLb
Rq8/JUJ/sctWKOKFLkJIi3R/eTvjSdm9DdAtRUS+R6gd2jP1q7/KQn0TkNBxYwNI
+sB/hnKTz55KKvHBiSF+4Hs+mT6J0PgmHsI772+AZY9LHKAWJrjIFLFAZuOfR8op
/mwLmE8X9bfx89ntkBbUw2Bkw6IuKCS2bNUmh1hImA6ZFkmbYWsQlv40IMH07VAo
7YNVhB6bVBuRJzKvM/yFTqQI8JJ+wOdMl2KPhji42Fy4P/gRxNwyMvUeOEMiIOCU
Gh6tihWYS6m1zZvVqvND7mp6Q7fI2WBOtQI9RgnOpxtzP9xN2xj6NvkxEg4lTFIb
oT6RycRvthXINY56QLvQwXdgzLrWVuC+nOOmRyHuYmtuZFoVdhU3l5dO6JedPTTE
E4qdfk6d33ZIgIN4BlIlQGUwRqViT//ESBi5PyXnLLP9IhBBqXZ/vir7BI6c8Lr3
OOAZBtzWmgKHqW0JGGD6au7AK02vs3nXGFvDKrGSUGQaLXLz7JSwbcbvDBtnn4A2
oYz+IY70uoPVJO4UVjjJpsFNPRkPPnwZUgB3SQZs4Vu2jOD8A2nNXwYFefw6mHpX
XlQwaLdlKCGbG6zKBX2z0UJpZkpXtnNX1QL6Jk/MuilE4LQKzMpFKdeIh9cIeKYf
2xjFCuPNbamGxYPMUoY3AEGRgAvkQ0TI4xPyRBQiMQO9Rykd9aaNX5DZZ4u9wi+m
kb3cP/b+RIRXRoG8YplW3PNpxkmHDzp0lVi5NhaqKIyJ0aUnlCJ4eRmQa/yvCG6S
zBexTjdMomQ1bmJGdIdGtbyhsPH53cX7USz8yx2V/YSn6kj0CFkPP60sGBRVVYGd
4K6MshJeMS5O/LCo8KYI1zBQVorrM7nQFDYO3AjlWt1I6HFiGcMKTOd7+m5O3vZa
XybCcIt1xAgQgXQTaQLrMv3IfdyhG/uug/6ItDpsnyJ/WUh0qEyB5gb4N0wjyjJl
LDsa1etX6V0oMsxgL9zDm+OPrp+bp5Prp5dae3aDQnArj06GDTCN0qjKPwXoJRqC
l1DJ6YCdgyh4L+H/JtaplOBPmXvlXPUjP71cVdU+0/49hjy2CNGnVNVsrBfPSrzt
TDFtJtdz3xY1x16Rb3sKa4925ogG7KzdyANUUHCE/GSe/Bw+ym8jj6T3y+cAy8f7
nJU6itMnDIH+ARyDls5QB6S/cLs72iCU+Gf5a0GjF+N19si3rpsX0Za4bixx7jii
bbo1MEU5MNY7hoIb6nXUa7QtfnGTV/pJahcHhyt8cjw96GMYhqSpbQ+SmZAGUtjz
vwRel/eu9M46PWx1Vx1CT/uI08YhpR0tzf5pfpf4c1bpS0aCl0h9yn/NaQ6NoCsX
3rUVUIjPDumt2jBDPC8XgPk2GW1Rsusr1/6xznmRMvB8empj3vZe78CtRkecBRnC
qzr0kQncJeDNxj5qBggHMziNrX4uHeCsRvlK7Q1OFQL1kK8nj8BOPV6YyDdlTRef
qXnwNhj9eKmeX9D2igTGEitvlc8YI91dNG+6K+odkuCaYrwhP75EnJNA6KH0R9iZ
1kJNxFZyZLvsoyxd2UGVzJkmFkY7078FYbJYUYHhStXPA8UjXL4DI5NEH9RmMg0N
rxZunZYHK9oV3EAbduGopCm6GChjA6SepQxZMxA37tutWhc5pkViSwbiY/Jj4v5s
4dA+mEHKT1wUGhcUyn218yNg9m3Jq/HPtgYmxoyCIIe+yPj9jI+BJV/8mrdRgdvM
bKJUIy6BtDgFHNa5vAdD0CMUHViaS0zYerxAwHvCnAXGCFWxi/NNxnj5HnxfVCN8
qdWkUxmBlsqMS8bIV5TgbKrOVjQrTi2RTmiU2dOycgs0IHc9p2ZIYK8ih1TsVPRm
I86FDtx/EMfv/AAVwKWLqHr99Vfsqo9Mlt5JjGaGm5AC/K+2QgwN1DpvY9oTfll3
0PYLpm/0etOlY4mU5pAvcjSvdo5u5UreysTyiM56ov0/v4eBwEURu5ozJ+k3InVp
7rs+WMvNfXVS+wJt/3LkKDp05iRAA+1wmLkvTiATaxjOTaVAAp/qeWPIfhAJ4ku4
xZZZSStOQjD6dvNPQpL60Vw7DsLaUjESXX+uUn6vfMhLM1LYgMdg5vhmeIEZKvi2
dDtFETJlLL5XpI5Z2TPH5V2bPiCIcdAESuelZrI4qODff1vTKOLHohPcnrmI3hWt
VMlMn7tIeiBd88XtbwXywNuE/R5jw78O0wmBpeW2BF90WkiK/kNJu0LJw3PQrUXm
5zC+Jn1M8HTV/VvIRCrLVPQO1i1O8sl3VCPuPKDtf4t8R7Qo4OL2yVcNGLIwMHG6
WC+6DjFxyH7EICtT/uxboFOGr+zjlX/PaOzSBSt+M1AiOSoYdeLufiI8qNn0BO6A
KSy6tIv2sBpxAolfBtDqCItkpo8RrGed/r8YrbnEJI0+gxASB1J92MqvdbRZSBsg
PQ+X0ayinJwa+X199uhxf2UfX8NXrwzC+PTKi9ZcbfNFM6FfkTGoydcNifVOm8/s
LtWN3mz1sC+899ktF+ue2Cgd11oeJLCDK7SFpHiqk1UGXTtc9qZWeCczfr1YBROn
a9gcSkrM/lMrcmFkWcX90YtpJC4LX1CNpXJ3oOWCNZ7maqMLAFKxNujvql5fXukL
C3VSuKLW6TiNg/7kzKIEi2DD7FzgaCQ7g6xMsmmR580XetB6Tx3laV6cUhqpbHO1
oKHPZdq4dRs2yG4979uplVT+eEWzBdGdoZf6s4OYZOKPctqqgNkVuNOFBgEi+ET2
xkEElELffbhjQKV3BGSee1TMZVo28gwFibN6lpYNFTCV6Biy4nFNgg5Il6HJQF1H
vN1d2Hv3/H1Hzfmntf3nBZ1rKmvCLe1U2LimuugcTNASenc7d70vaPsmDGBNotX0
0IWXhxPUuXrep+nnP38Tj65VYV1+aw/qrUGIzfW0d1wFJ6H9olnQMEDtfAQ33LCJ
+JOZPOm9tGdKOIlKM9ZmNBdQxTcgviuRZgzfcsHKt6GAwngwQo2dcI4+z1Dq8DLL
Xz+GiXD/iLjNzcwpzfKTDxzmC/yHnzX6SMtTD6qNstg5dhSMW7my9c9nhJS1Ngen
+TV+SKT1ZLxHxM2UQFMznEdnCSUoMU4mXH/+d6tC0tOAzJNz2cLwPyhnhvaMlmGo
UajpiBP8/hPj+n1ulzr5vchkIFWtRYVhBpZpbFazuNQTpSpK2Nw0b0IjHk6fM3zl
9MyafWXPLAsaWuk+dJAyqQUgf+I8ouiZQL7Z1QR+ImLjKOui2zbQxSkXssScGxwV
fzmdIqZrrMbl3grFXoquR/Hlz8aUOdspnPC5e0JTUczHp1pHX7ruUeuNnCfhRo39
J2S4tLIeWw6dA2gjx91ls8qQ2bGUCwFUocsLQ6oTmhuimfiSec9bQqyonChSC9iE
g2ZkbZOiBT0dkLfR3IPu21XIjJH5SWv0iHZa95Flh7ztZH7qf1af04NuCo+V62rN
8Z0SyjPoUJPiLuj5PyrFc4KSJkPABpx81KY/V9MmE7jLhIHZsRlik3FIaF6U3+sL
4sKvj0saaB1uKUkVVufYnd0Zv/aOKtnZ3aNyeBYahf35oKCvJjr4basOEBSzXevM
Gylhkhev7dtAwxG7X8TVp97xcXjS7ZHKv38mplbp60StHzn8ZZ7H51Fw6C2UXnkt
+GvJaqE2d6ftr8C28TLarPf4gKywQO4JyV/yvDB8wJbBfyrf/80wt/P2awQRYC6P
1vO5a/czpS2kGOO9HsP0E1iJDZ7i/J1v3VYHQcDKUSmFRZx1JbLdF+zq5WAvZLRS
0Yq8q584zZcg+VSFNF8ZstL+LB/WMZ5P30Sfs+UsprXlhAwopBhYvT0qSvuyVTqJ
Xu1R+3o6D0cq9Ci6ulso3y2oV847hc0WVOkldz36UwZaOVfaK3j/VzzRE/EqFEtj
xiBgM2qf7yRwn/VaUd5j83othJ09IkkZLpUTga5gf+iUhvL1wIJ7er+QBU1qzXxg
pXuc8DULqNKAxOA05yPMa2ZIfulwiNhb5SCrsY5zFwq2pEpSQkIWfdGjHG57HJO4
gn9QaXxK5Q7E/ewIiMukzSBDso07RB+7hB248+JnXqJ0vnto0nqfKsaxH8k0bnlr
cJXLvEWWjUy58Ft90gXUKZCZ4i8GJ61JHgdCDINBRO4Q2B/aiNQrQqIIHHBVNL+d
zrAX/r7Zoeckx+dU+ay2euwUNAdxW8slp9T2xwCqaDD/BFay6yRdrgafyr5WhF26
GgsJPUFeCV67Sm0bpsuaiWUpdUslL+lLkzzfvLQreyQiVDvcflUsHFpNgSVZVUIb
1w14FssqvW6GF5c8yjUUMyJ8ENWsY4VtIRsM3zj9ypWBStMBzCxyJExElrW7+lCo
Zv8QKw/SrDvMgcPgOA0cNs81BCW596ybCmrM7ZWDjwqlkRSwSfJ6ZG5qh7XN+zKs
N8P7Hd7EaCbF3IItrppNiWUSvPUp7oTqSW5TsbuWWt9zFx6MQ/ghgERk8Scbn6kQ
gwXUIfcgdB3H+UCiNiR1GSvNAxvdqBsdXAFMnu1SV//QnAvaq6Med+ARanKo8KmP
QLgsGN8fp9IYmCjjVG/kdKkVo0Hvmp14Z6tlUqXr4IEyaQ5bwezlAONfGluk6xsq
+G7KR7GywHZhgJxZ0pMnjGWw1GIeCy5FAhapkyGS5fYI01qU3MS0o3CcP6zrx+0L
v88FxEB1H2FStAFUS4d6LfCo5GvzvBcdfOMLX3wxSRhYcGHjCy0dpSnWM2IMquFr
mqvqv+2xMTJ9GwWdm+0juL7BwjbS2WnG+GrMEix7ZjGofOwHZC9mg27jFc155zMN
ews7aqKtsMrmWIyuM6GdT63OsM8KcIBLtQDD80Baa45aFRZnwi7VYW3IEyREi2sg
UnH5nLLdoofOuPv1eqGvY/V5fBJhRW4XhiKfACoiw61TY2m4gPZQbCe7OKSP5IoG
jQh7i2mSlsrD3tooSfmt6nZ4A5aflKUeAsJXRQ6MtoOsqUOTKkT+uJd0FbUyazmE
pfe+CUCE7Ii/Y2xWXI+V9u391L5lW71Ef65hkk0a4/ZTnD0vf71mlgl8LZtUL8yn
oSp+Hbl7kdIjoNQBYABnD/9TIWgWEG1NigTRLe0tBRkReZ7lc9N5vWcNjcUbOGk3
RoK1hw4WLKh7vJBoEJrjr+PJzQYV7skaK9HP5MfTT9VOP7v1rD1RiM/kNWkl3KzF
D7ogT2SUsG3dobBGi5iKdDVrTDiYWsEAaT5K0R7Ey4VGhK2XGnBuNjDn9Fot9ZCH
ZKQ5Mzor7wKX/5jnNlDfcCEkD6PKPrVyXyznHRFbEP53MTs/b+iMGYBUncnA6pKO
sZdDlRA+IuRsGPqdDBTktbdBKZp6tBakn6oyvskzMwBwNms+61jYhuU29LFlyIH5
yvTfJhjiBKHGQztatEBtxZ6LrX0T/UCKD7Ek66+/E+RsgaakjGTco7boUInFXHTP
v5TxBlFUGXuxgAEZSzz3c18DlARqsxUkj2EmaerK+sUGEZLhTeOceesZZ1vLNdat
MjpI9s0XSajHIwjECHLoCY3IuXJhWJnQBF0qKPJhzi9YxFjd0IIDi9mI0lkOMBQT
CdMNWBPu9tlBJIn9ovBNfEgkX4wOiYU3iHnH76zWYLXGWisrjWsSiSVl5kQ7s528
/f8idh+mJWZDkMFAHzIlDNK50kK0p83gQKIZo+DDsSsIeECTADUvkI3+6VvlmKdL
5xTZWoOWmSGmsF/hQ11IyiGH0Jp+H3Qre9HIohlegNWXNUGP9VKwuLIYt0x/D3QW
Sy5qTV51nMj9Qhc1DGKWWAIk5luecRc9R/d7HR06Vg2FFQ72qatwTJds7vt2FguE
OgC+FhnOQ4gfD7kn8DfDMPCqlmcxEyUVkerEtO1AwpBSs99s3VryPjMMdvFY0eze
fptB36qVCeq6Fs2WRta2Bdx5z8O6sODebuSokOHI94WJtd4bFHsggpPrIU7f3bXx
QtYbZv1gBk8qYs9s3xqubIITOf+GjOUNsA0Z8aXMEkl25J3RdaHwKQo/VJ59TUXE
K+yeo0O2lFL/r7oluS7aj2lU7ZUfH115rBPidfC7bVC9/8ewArqZV4laiNQ1V3l8
fbw4+QUnJyS7wwebGS8/5HJs8RIHWj2Fdy1oSS01+mTp454lV7WTzxfCvaQ2Qdqw
9TVQwRnOF7r29lKiO0Q+1BGM9yTCM6b17VwPD+0U25y1tQp83KixnHw1Mpvo6ddF
9nse9EgD/PpngVX4yBGPF/1u21YMS1/d9p6WBrtKboO9xaqz7yNYeKYt7CZ0x9qw
WuXPnkQWedzFa7ANJclizPgkR4WKv5GLyGf1ha2LjNMutZrjtTWgPKrVOXdcbAdL
5eaub583lZr93JgVgzp2Aga21VbIJc1ACQ01oZ5ygvT9lwZ9pkYsZfVVhklJr3np
RJDMJDEtDT4A2CCiQwfsMr0o8aGvjfobN+mvEhVZf0/dpzno2fCQyqdC7ULrGmpk
CgWG43OYciQ4OBC2wpGxhbKS53LGOKgZVqKLPpMuvS27e7QLnYtFOtk1OgtLwaU8
dEeUZczYGT2R3uOJO3gWovQvqRRvh0gspR7COUdGV2tcRS3KMt63JfVal/fmlX9e
xZfJZI223mmUkJhG5mIJj4iHT4XqNCTIYqoCSYt3gduNYPJ+EhkjL7C9juCt6nXj
H0IvluVzpyXEsENX39PHl9LU0i5X2PAoHLGGshD6Xe01uIOX/FjlBoyk9MlVb8KL
Vv95BTNzi7qcv/KOgtseru1pJB4pqiy95zHwj7Zos8tG9bZHQ7Ay5Rr21DC2OFx/
uc42zyspuvVvvKLAgP/ITrcisv8wJcEBXDu5MIUgDfHbKijyNLlkn41AX7abO+ny
Htc2p8m3L/v50yFklF/xBYWohlfhO3LD5orwiq2Ji0+TWIIQeKCSaIjryOF7JOCp
LyREmDgz4LlliCGrLnmPPa9aCdzieTGU5iJ9C+jr91+d5w1GxKCHJRDpUxL5TLjb
5RI1Qsr5srGZxEp40NBCrm7R0vQ7kgv9lPzU57TcA031Dt6f8DGrwQ8JbJcTrgMs
90nhDe8x3ZFU4vd5zeOQH/uWRImuoRJsBDWVQwGAYpPWcZ3aJEi31o3EDy3PsfFV
frBOk96UxZN3ezuFVle4BoDhf+DS4MbhcIDEPvnoDiLaJJqDwCIGAiOvz+m0ShIY
A7dtrcrzv6OuHIu7wfR9TtugyZpV+GSsdcNKUaU174M4y0+GzmCORn3mU/JI2yCW
602ul8NEVnutkIDW+nS5/dxvI73LKI4xbem3WdiS3wgBUwNo6CiZD+vfBYzXXl3B
Q0vUb/RXq0d5QJbPqTBlgMj+/YDif8m+gkhM4butxA557pm4AnO9WUEd8PdCT8Kw
IBdD8mIBtIItO6tg/ImRQmU70Rs/WOCgkcArGjs9cYLuKwZS5kN4bRmZ6Dxu/LeZ
f+4x5G6PFBg1/SKaE/KKQwgydgYIedNl7gQiG5awb0kk2HRv5+rEjCg7TClngfUL
RW123MtBqPjYbaHcBEBfMycMU8aVBcl4mJ2JVfVnaH+CjB4hY99mudlVyzQD9BQD
mYhlObkF7LPK+pWNjFqdJ1b89RAsuaEWVWXRSDiCHP8qogLbqMcNjp+hCWW7CUpR
GlO+8KLc2YVrZnijPrrGNS4nNOqtbK7PXjZ2uG0dLncIzkxvCpmpcBtNZc56s5kO
1yj0TRwuDjphIy9/t5JPoaAtgzo051ViV8ha+wz9tuFBHoSP8rGUZiN4sq7tkGSF
LBT3abM0ReMowsYI6htPWD1fC3mDOwURtQTQeXdbz43+s2qNqw+m2rL2o/jWBHuU
C3Y4TXMStNHfhIfa9Kz+hJ9XqkfxSOaPYSo4b/UT44Yk5B6JaoQ1ECx0GOx3Wgwu
z3+TzQUaUzxuMBrDFM6SCWaCC9iOlFCgom6CGRWoY/2OOZAPtdJ4+nASE0YU080g
EyunR/k5t/qNk6odMI4n4rn5lJkOEybJUBUWLG83T3GRUCl+B2toIiPOUwsHuVgi
9mTmobrVz0oQqh0Uky3lrka35221AsqYQFZJk9Nqzinit8MH+BStnrJSALzbDInR
veXsRsZzKcPwdqh0pH799qBVPuoP7tPDh8MeOFS8W52olKD8xmKhOPS2Qa/m6gYp
chzHU6VgSstm54GQpOxkCzOtKCIcSR+EQ2VjU+bLCx3zH/gD4XswXamrkM9MpyT+
DlcLkQMvNXia5ktFkqaH1aL+RtZHjkPZL33h4+/lG0yDC7KkZWTLQ7vFjjFARljP
SFPx6/fBci1XvEqCXZxiNErbT18mJYbvIiepxbYKF6yYSWRE3i+1bq7Wts2Hshqw
NGKalEUhcZF5d8/i2en0PUbVwiKH1prqMLuzuY2wyLD62hn/liIJKGd/2zl/HqBF
f2+bY/95LKy5FGmCYERHkM9wyU+EyMDZc7W1yJZ64f1ZGolrE0jNDUJ1AzlTNWKO
DzeDr1yiZ5l60DYS3R4CK/KGOqGJM5TjyUdKupnC2vIwGP6MPn9jntmYFMZrloBY
PBnBukB2hvWbbLdnpKO5fIUIiyt87wp+5xGYZ+yud7KIjxcfxmFFgycl9wYl6+ZR
4reM9nTnMQsW1t82o7AwxQKS/mc+w8q/Grmvwf/xZz1zloreWwrGRn+NyD9VEt9F
WkFa7sBPa36hMuQHOMq9gHoVvLnzkUaVdnuZoNh04GSQYntcLzwI5j3Jl8nwtxUm
e3rE1lWRAmggjLkJro6Ucq2RXhEPvVfNMqO9ZtjhxifdRWeDj0icweSxRmqDdqGO
bapzKdUG8fxZ5ZfAvmrjxjaOL5i6uH0065QSrHRMUC2wLAMDlWDGi9JExyIWuJkl
6hmdG07WlXoWu7AYj0y616yAAvwioiI4ngSEYuMdfLhGfxZNN4X2BvCpVp7pyzTc
SiIE9bP+LpynvgYMncOQVy5QY+B0d4IEaqEPWA3bVn5TSS927bJSXHBLOHR2GKJG
j+Ng8QvEShEE6RdI8rrSJpiVCjzOQcyryJNJpzKJzjsWRslKJCwIL4ShXTZgF5vT
k7P35jj+zXl7lfecXv/n0s67lqkEfVY9BOYQ6XYO0krKMTEgae9xG1I2BmIfTjT+
npt9ahM64VGEvp3PDhBFq3jb7no3vPhwmkaBpZbpJBnsyTRENhYpS1mYgI8gM7fF
8XCfm4hEgwGmpJ82QPQszSz4NdCqgpBGR+1Qod4Q5U5E769ECQEVmgL4Tc85P/Fx
Sy5Ft875aWbKiNby52Oc686yVFNqMQOfkfLt6BMD+5Xh+/9C0psQC1mBHpo89fQu
+RHhheBPqkUx/JXL2iqsGMhWy4lho6gQTu9S4CuA4fjRpG2VNakeLWbhYUKquV6Q
er1XVn72dGLOTgKqZOwJ+FqfUeqM5InS7uduEpp517fENrylGcjCs3bnGXQSl6EW
J+59GF4VziCU4TkZJSywvhBrVTQh33Kn+OoxbPrpeeQbjhwCH3ttmeiUT2hbUEMy
9xeLwnhvBjOGW1DRaYfw2/3d0rhYyPhOsc8QYrmocYcZyO6SrA778hvb0ZFrSIRr
ZY3xbhmJ4/72KS9jGHpY/C5a+vGxvsd14VHY74BJcl9Dy1DtLq7S9wO4lLqPqq0/
oH3vH9nzUYYt5Z8+ot0yuMspl6Y40PrCJ39+4TGZzPI919n1E5CNJmCU7uZv0v5Q
YQZyyKgME/O2YyXpgY34vl9vDfmXOBy05svTWBnWGvcGk56pIGFkX1RiB5lU0fFP
s3vZKmKTk2nCanpigiN0yxqfrYCS74Pw4khnyV4dclHvVg0A/bmqKnHafmmV7M/j
bP5+PlYSndY7Tqn8dc8cPSEWEkRwPmbVULJ99Xal2D29L5GSRwX68WZQYTpJE2ta
v8XqZEaplB0gMv1glEbkxka2M3vnblBVY+liF+6Ws5Us0yL1t/lKu6DkcreZqYR+
E14BfRhNmgY3h9TS6CAeXBiFEdPBlYaTN0wKknEH/M6PP50Bl/GdqvLFU4KVBIA7
n6IgsTWpmXTKBzJivUcuPHx/6hjzAnwttKdBW7tUCup5gSC/qX6XlaRZId5imOR1
lEe5FhtDPdV6SGMDc0Nq0aScwOeAHO5fP4CfuPyMYATvZPnui1Ai6JZnQY8S8GDf
zZct4ECwW+IUTM/J8TtFJ2mLWHKUDrQdztUIFPtu6fjukEdnfJi/H5RX6oytsuRA
pFsOREugnSj8Y5ynMS02rS9tLj0qynCUUIARSPKQOtGSSDt0wWBebp14s7UXnQlo
oIpXSCnSU6fgUyOyxNgQ/bPNUvJadD8U7+WkkjePCIySP358dDtPFStvp3ndalS3
hAaxor09YYmxB0mpnb4zzMBsuUal+Izlj4jS3qiajX6j3Brn2ReevlO5eMHAXW/d
Ul1MR7MgPuYwcgqlA+3d9oVDxsZnmz2D24F6vOL5SSNbFDBjwDbs18H7pY7hmnwK
du7IaQx/xuzMVDZdvh9/ccpOPZwwnJCEV906+fd4MMh4bnx9Ir7cOBj+VlT/s76+
6FaJkNQHcRqM/Nbn8gSPtGbdFkSnfBwVALgYYztZNBo+8jAtSlL4Df0y3x8m6eB8
1kHaP/M18fOZ9RhoXM36scWylYkE3ae25eJQobjFYCuzxTm7uzd7CDakOQDdzK7j
iDnDr9nV2ymPdC2FYjkNjgHh0gdJNxpJCCZLLzHaC++EB/nJ5rIzKe+sYf3mfzol
t+mCsvyTBPnYtL6ncsJL23fM+RbTOSMiLeTSvvdIW/few6bf+H2YtwwNj7gMqoSp
lSKkXK9rtTCEPd3zJnbhOYwj6DKN8dE7rs7Qde9BiIVGgUiWqspS1LXcYoUgymqS
QfDJiEqug0GF2iubDf0EVcyV2bUxCbI3+x3uYlaZxBOybwkMaUNNZa6/GQ8whHa7
AEOWq5j1V9sk9biDdiVXnBK7gAXykjOdAhwGpmNiFN8zolFkLLDitVvC/EWKzkvH
tRlqbwqcw0MmVTMk6t2Wqf3Ejkl6CDlYLzbuzj4p7lYyBQqY3D9e/2UMTfYNVCRy
2Q/YQNjVU2laSs9KI5n8VGSy6ZoFE8EcrDQvJgOC2pIXeEpkcSgZoytVxhl3cAVW
+XnAVhA0CqUklqfYEyx2JrM9yp/2r4qwEKknr4hiyOT/WOXpTsllDeM88MLtXi5r
dBRV0P6D4rYMhn01kVWM2f5FXfQJjJonRzXMd8KHVSRXHXFmCKeOcS3ilNj+/mWX
lFJjH0eFWauteYPH0GJQKDZgwXjsyhPmnTpKaaLr5cfL+07B9DvaSXhvPjDNRBzu
N9zp7NtdllleEacBVrXA4UF2tgxZS1FwnuWaFNSa9GXfuHUfq2xs4k+ecLPaffEs
yYNiiPp9k2aIaq2Y7xsf7R7SNoPyV4hH6O+Cn5tj6Z20elowgGl0+RAcEMmkJaEB
IVFY8Qsl6OiG0ioamfiqQCYOld8gTo8zYxi9svd6KCMCi9CwPi0bOTokB8n9W5YA
k0uOd3COcmIFa7OCAM2rlFA5MpNG7UmlPRIYdd8bgACZwBpbyfiP19Ogra6kT5g3
KRP9Tsmlpf22LbTJjJE+yA9VtJDyTp5Mv1Xx9dgLXdRK8D8Dy79wNg6aIzbSp5gP
JH2Dxhu6kGsg/cIKrpZQ/8/lpZoMGif3OfJCpSfwTOmOxBK/FveEoATNydWqW6zd
j70zOq0UOCGV5r8w7UTvrGWkX3sFBnr/Yzd6oqYIq6rSUcgvgVMPasUiNGOi/YBA
I4N4MQCCThYZqNZWjwFfB3Vq7MaMZ843oRYV0spV6seYilrFURxo5rgOop40gvOo
ePANo/QqrowlEhSOgT9wxAHVPpQVO7MriDhI8CQQlpAASe42740xZ7ffgwh94lNf
xpZTJHBXnBhgGvaLiLuIvm5DfWjf4lyP1zvk/O1LBFb5caFc1NUaHvpGC3n31q7O
jSCPU4t1BBze+jtlS2af4ZL3kpg52P+Xsus8k3l9uvIxZCQ6plfPa9guJDpo8p6R
ygo3fYrTCMXkqD9fcn+CvqyKFQn2P0PBCZ1HEE51w4yvix+PvOHRKV7T3QcCkAW2
gbKKjF+DLUwvVXCZOAG5EstEgkimHznvuSCAIY7S9h2JsyPVo+J/sT5a0KN/lvMd
JFpzdmddcDT9PzqBuPq5jYN/Ffn+Ls3xRb61dUYL708a98UC1fDTibVGtRr8+UvI
cvXo0q700N7gCNLKVr0BFMpY9s3GQWXpA6SJk2dD1kyTHaWPaUtiLye3pQQ9cheR
31m2c6ywhdF6juNO7TajP9NfiR78gcPDEmj0RnSLYa2VfNrq+Z23wCsehcCgwksg
KfrT7DMUKFDPXaCFWKhd9t/SHMGFsxCY4CJoNffbzTmDxvPIVw8vs5cmwrtiNJuN
Ot2OB2qfBgWB0tg7sAXWWob8kFN8paks7uk4D2A6MwuZXXcSGLxIPlCWzrAIuW9v
bWg3tqecVoaV1rFwlKjJowsJ6qfq1OCxrZn2RIFppnHaWqyp+JhxRwdjHl9ANfvJ
wdI5UUWmUe7kXq67qnFmDTKaR2KkFgUSE1qnkre7NnvoZlvc5dpdMcN0j1XEIHsJ
H/oEPl7fluGJlyGjVyzfckg5iWOYLgmd87bNXkSXSouyxns7WVM5Lu//ZPoa4QR5
jgbhtcxD+o6M8+6Gsyey1hsMvW1CZCKB8K1B0Csk+tEg5nh/Kx1vlk3e2hESuYSp
5yj2VgIGMJwrYPZrptlOeLW7Mm8UBHERvqEB8gtFa1Ru1VDVEF1oj0IiAtxAiQoD
zF6o62ontDsH28IoI8SFYzj/L3qCzV9XsOrXJbBAfYfTCS7HCAJ1OftKfajNp5mZ
HKpm61DZRCWNF+Fm29M7+EV2Dw0b01nNjsVRBHEocV2ihwSAwjuQBBeqyTFJIDOm
xQYYsp3gPF12wKkeRcBDK+KECpeZgYAZFhOOXs4fkH1QT7eGnZwfUqAWtobZbPNK
JHKGFuxAUdCs6lD98c4CNDZLq0kXv+jCliRuRCANi6pel5p4nVqYPWzU8JCUCQX0
WOUPZxc0k+kYYhHB8S15vuWW6dJPbbnT5lkm9cV/NFUfY6qoi8vuBWv9V0yiRCLN
IyiyKmAKSkjMmF39d73314GZ8iXRtg3+ewwMecDfz+wf8TMgEugycNNU/sic0kx9
kPC44dmYU/7W4aZatiec+kXlDOIjTtfFV07bsLVPWHpIJU7deBSTdCMvjN/H0p7y
Dc3Z+fTykl6R3lAFE7XxOdzH36Iz7n2Rt8jR9CdhARjwSorZOqeePnmduXHY8We8
zGF7e67LDz7XoooCoZcld2EUvyv4rH+KuZiSU6Lb9p63U+UYnF1uSSwjn4DQdR/X
qaZytqR7z1C1Ia5SRtl/hYI9FKBf/T1rKdCFXNttSR+qSPpsYM1Qbn7DZIOmHSF7
Z+XQrclFBxD33VZ96Z6pNbdsZS6BQdXYdySsDwwoaiTmm0GyyDAldM7vEvT5zuod
+UbTSMN7UMhwyNquwq44yCGyS8ZI//auM9FLKtlgX3BOE5f829fXna+gSstGiDa6
MV+UsY7KkO4YjVYh/arPgfO86+ZN3ruUUpCxeTqTwtEHRgd6Rf57nTrUENb18ui9
puW/3IScLc3TDGWcsyviFln8utBZ444AylVJVPtgF6r86d6U4s1OGGaTDX44NNnF
0zkNXNSAiAGMXtmE6fLqACY7dKbK+uV/K+u8nxjUmkLsGhE6yLg3cr4l+rPBSt7f
YMJZfxZHRfqvSlpdmkknPNZUIPMWoWsHrfz08+S4I4E/ZlY9vTMjaFQLZYZaxHFz
QI3IKucsdIgZFYZYVEGN+FnRYe3E0FN5s9yTchKTu54oIl4anoNK/KRzS8czIrfd
THwgpnDErV1dTL0nu4CcRgCSls/1id5Ts5Mr2enx4XrUiWkQZjG1eFSovq6xSMEM
ZqpyS/B5URLjd7fvLR3kFGDco8UBtsaQXW9duqVUQPsLTjFWYL6p+uefWnGrH3pM
qOkBueBie75OiwGSXgQNZ/2RFZkoEVWsyd1rHVRCm/cR700jcJGcszltzFhH5Tun
ADGIhL84frVQBoI5AGw8jiTn6jl6dH9T+ju47r7Jm3rLW38VDl5FQXTIg2Dh43LF
mePEgtiv48vM1G2zG04+ab5UBOP8e2MTwZyPhVlaoRZ0vH9JEPfs+4eRT4NgHgh3
JyMX4Sl/qz6aEpLFk/rs8qwkswLTRxhmTouCJutiz0N6YrUFZYo4lTsIHHnW4spT
kHsHM+isJE/WTUpzQeGacgh1wUzerRQORQZK4XS4+O5GRIWp2qfGqICIvN+keBZd
HUQPPkbhGD3HCaTwTPAWWstSOqaDTeGkaSslaTyjV6FMyzqKD3zVXHmDx5daFNhn
gn7OMxeDatCv7PR7JyRtT6zvwYBs+Yc7qusIH0sV5POY4S/xHxFA9QlJgO3yFydZ
0PuMbfjuRH+kQwRFc9dqu1VQyt3NBNLdNwMojIty6YFnapXoXI/08UGXV/F6BdNI
bNda3dFUfihbS7o+iac0plUFk7onKP4fqzkiv1Y7OzkDcBDC4UTMuWThoAlcLkay
iWoEvI+COaCCaDguIV+pNVDj0rmyV00uUlgymljRZf+M1KBItkwtyxwkJvBBBXpm
SR/VoDHN/2magsBnxPVVgbpND0D3me84piKuvMsPC9tC7Q6jqBkne2NSknb/9i3a
FzXKbe3v+JtV6TD4aLzsahVGaVbjOXaXc1CL1BdfINW+76CntWrl+hd5PaUfX1XM
3B0v5Rq09e4Huw3F6mTlCPpMTas7FnyJfsoNsUC1JrEL2J8rCzKVb+sPUMRLUvOI
UcA/U65mPC8RbamuSPBGi1KyPMBj/K+Zvym6KFTGmSRuZBYUQpvbFaX8SIBGoYnT
FRGjLGEyGDUYIiAE9py3hh76zByg2VmQUS2HYXaOj14I/38sRNuoKK7QDSEV9rOx
9HeP44K/k0TPUYQO9ParDScKv/MvKTHyGtcBSoL1SzSiUmlOUkR8GuPjDZslfXcV
q5gfZvLxdPe9uGLyCTO87xb8cwjfvu7d8yGIyYOvQP51mrcNMLKn8BLNGQ/2wpQk
NaCRhNFQwhSd3gnz09Cp2fkSXeZIuit4af19pID1O+RLuuTo6loXSBOBN82dGWnH
aEiYTfn4jiImM/uTvYTrM9nhNMB7qDgco5anDqBR5kbx6ub+Th8/m8E45LBp/XCr
nMT4Zi9183kNv05wgX/q1bBft5I5/RgWkBczog03L75jabWi2Iip2OjM1HwMZ2y5
PtWuacu4HQdFHSV3Mg2frbCxHeYnx5ofjZU23tMIfA9zf1ALngyEj5NHadPs87Qu
Mx0BiNlH/+Pzmbm74m5l4vGHnthce9VMiEKgYrR/tZPjmDInmKoczc41OYWgpQfk
dqDACErjWrxkmGp9LDSe5DJw9eMtD1d04adBWGX5ezlVTC02SHEcGJQlCYD2VDIf
t24l56c1QWzQ3p7bo7B5qJGfG/a2Sat87yH2rKdwrIV3LU8QxikXACYasuKlr9C3
ixe15tL6ApFKmEVv5GoN1RExnZWbHDy7hTqi/OteVfRztCoqYBVAlxhkecTM2JTN
LXBcI+jlkcghx9YO2SujNTGIo1U04rX4Dxwo3PnI4Q93GTAosKKfDNhTt6GCxgwZ
u9uKOOWxoThKAh4fcCEhm+4ZpPbnvjcyOdUrCN2EiQl1+dO++J0t8aK/oElgT/7f
sXPDSm26dkihQe/wXUr41mkfxvx8pmBzgor6DpDeJmGAFP37OBVBIwSWOOad6+QQ
LryGSe0gGPMvTSLMfQBsKacgCKWY0ZNROBaOhr4AXxrYaGOVJb0aYndGixJgivZn
hW85Z6ygMSwRvoQQbvGymJxaOezdxlOzhuSzJATEn4eGb+DNDOJES+xCvevx1w2t
/3RexYWDm95XsmFrtweG43HrOLB15GW4xIQmA4ffIiLmj1JTyTkN2S9jTTYi4rBK
Ocj9upRSrTIUs+JIp1V1p4CwK0YttuAfAzowvE6uxP/iaSN7CI1MaDlVOqtvrVD2
NOb/y9OaNSEgFfd7igMxZh+V0TjZmhaFeEwv2Xd7WzLdz6l5Ah22zMaUuKTLzYnL
62z04crpaPD1V9yxkSS4+UpcWZjtxmZfWzRXAvad3JEWGSJ6XTBV/aZWy02l6WPS
V3NGT8IugyLY7Cwr3FJxdl17UuwfP0v8GW1isKsH8hc8Fw6ZTcrhwh1uytNjGzyI
WWQEbZfocFloSuNy4ftQbPgik/yD1YovV74ULM+20K0/gO8ZA46RuzBdABzOP38l
e9dzTOGFneQbfzuiCcYrrsu02q72ZBeYY4e/i+AYoN5KgRDLQMxug0IGbPLJLV7m
nNq821e0Ul+55BfVezOi6nJ1NfAHRpOyZY+NauPIAfyS+57TKcjec8RYgZ5FO5gN
BdB2US7TsQkGS8aKuM2LlvwqMTe/5cgGF0GQqzh8V9x9YPYQUikXizYHMXG9DUcM
jqcHunxrVg75aLzrxKjxBqqfyBkfK+odvK+/pgTpdhEMQGa6SMaG32ppHzcmph1M
y+OgHhO+x5MlsiV0H+ByJNkeDZjznt+KpFu5hQ0wPZdWJ0U0W0Zj4ejaP6wFfDvI
TqZpzBe7VxcjwLBW/v0sHfFy3EgZoGvDA2yj1S5vidwdpY1sp/Fk1p2hPmBIqLFQ
QU1mA8Xe+GNICZ3JK7R1jFK+MtbcRK7woYP0wX9qc+gCYf5ZhwW+qxjVYSzmL3oe
pgZpQE6+LkcMa1vJ+gLdDqcq+niQjoestiR3m77acRI5T0SvlcgN64iytKzis78o
xmUDlUJ2cC9D8e3Yqj4OSNCBbf6zxjIDVsEjAf0u9Bmj6/ReOojrkAC7zW21gJrv
3+HzQIbQf3s+K4QP84OGkMM/UlmYpG2UOhrqHl6PTEhOVxWyviNy5xMaXsxI30UY
VGwou1HYk1kaCR0HdNZmjqpBQCUHsbokzOoqZe8XRWmr5IQxBeoiJApLerUVYMnP
v+djxLS99XmvOBMfqMFF4rVYciwTJvj27EZMj5gYbX/OOH67K8l+s9yslZYbIVGD
RByN0nkhKoI2SiRb+SHOzxqwibdT493uL+jmEqpHDXB4tBnjgIN7uK/0sZvtEJ2v
nDjRVzOKPGIng7muAsNABdu3b6wJpPHxM+i5uttHhIFmx65ppt8z3XREwka3WMj3
03pdT42tnyDGzO8Keya2XQBHMywRTR7NIlxHxSRXQCUW3VVAHsPlFjh6KB9UIrXM
D7EotV/fO1P9s7wwfncjHMs9pKbWRQJxS17JCDSCSazmF44g1+UE8YsCobVWIE1J
B+9Hl+Rz2qD+PNDsTX1+cDT6CCouLPeiRdYrY8nO1h0DH27oz510vv/+FykRPsMk
eWKpzsgeEVJG1PBnTlrLtOF7sSZXRywokCNNKeRD+62rCnrT0UFtE8qldHrnIBe9
cBbfC60WZNMSkRWXvDA+9BCaVSOK4WQKxkD51YiHyKVHjMOa/3NDxOTPBKt22YQG
SwA0UCmz1ezPJCzB+wFoLvgIdKejKKXMq1BSDo8pCR44wH7t3ApymyiIWZlMyOsM
+Mckw5pmBpMCoXpNte+1Dzgk6FdyzJZTEYuf0UGmfJMHkDS+llz2d/x/3ny3bO9f
j7WbLhn9KotTfwCpAaUhvQdRb7AfiPNr4BtFEyRiI18zZ5G2YMN6GKHHXZUDBjVm
jYeCGNumtBr35bjLM9uStMdpl9ZDj0Uoa63kF7C8dUDH5L4SOLzm9pUBUl5zz7iT
ip1eqiU2nQhG7I3IJT8tim5lAVK4iBxKIZR9EEFLZdDLvKG82w5EQmcu+nKPnUV9
TQu20M8zPqTcP6ulshofXWoJDCtDFurzfGqaQ2JlfoepkFFebXkPWJ0zTTLWT5V6
TWFTVgH1z/G9elGQkfno8fv9zskjx+BdqZonebW7ZMJbs2P0Tw52klVEnuZYZ6ov
PYTxONoDbLFnat5u0LTRxHDmqz4jMntXvGbC9V3Ho8b51DIDqqAW8spXDPatmULQ
sxaIO7Ue20equ0l8SDQ+OfMvHKSt59rxNcSK5aaGVw5yGjhN91bqenHb1agjtGKK
HFfflerMv6Nir45ctARnAjwqNAWSSn/U/YOSZ+tmoj5WHOte5ZYJwMjAPgySs2wJ
5x8Perq8I+fNxC2sWFhy6l57UjjBW3oPP/ssNgS0WYRKHGR6qelg9YCILjBFtcgF
8UcR4OO2As4IErb/Hq4IU8vQphDglDskBVga+JipVIKHiL+dTPrKKqhS6WOEjdRZ
E835/wjznYfPajFjsHZld/kfpCX7YYRq6u5MaSzEKbGwCQ3QQG7/w7OJADXJa/H9
kmzdoaG4IrxO8YaAUTG8bUMVF/QJspoEPDudHr73ejdKoFV7O5TNrWlnhFILMETt
Nt0UCHq/lbSLyDsnx68pLu/bwUEVKiUYC0T0tcZ9J40qP5teCnUNj4RZUixS82hZ
bQqGrM+Z2Aw4e2brjqTrKQjwo/MwAwKBOx5GOugyRoolO1ZZ4BR2GYUtzO6zAMMg
Mixq+68G4HZ6FZKUMrF88JOAtNMSx0SrwVPM59foNI5GItFU6EX6054e4y/aKOJl
XkisD1o09p/HjbwtQKhXwIc0G6v2RfLMFo+KeK2FevyBbmgNNi60WhIcAyajSC5U
MVVAWIJqj8FmRa8w/5vDDyj7LFV6LJw7Akvzh5PJHYMRKQSfS/VWgx2Bhq0OYC8u
gJUNWiaP+pIrRcTmKs7s0jkVFBe+vTSGwEJK9vg+a4fP6PIMj5PrYielba1z9FNZ
yY8Z/xLJYwD4x4aU2gM7ZKblG0EyeOS+YZuvTCu9QQKzbkcEQLk/lyHgAHqxRWH9
61Uvdu+SrXFtOMPFMEmRXOgxjjxgOmrIo7S82XIIctFZoWlVls3/nl1vOJvMbepL
4jZzmks3PuaPvll+2d2AEvfMJuCSmP83vLSoGS7C+WRoRCbbppzfUnuAZilKUbUH
NJJWRgpHTtqcf5m9WRoqD5GW93wd2TShYWavanzJbhcWL7NsfjNq1790urQat4Qu
uMnlB3zo0x5FC23xNi8isgmaV+Tzf5X6Gdq/+BUcgdaC0MAi0CsB1aKtiHbJRLwZ
qJmrrU6hcCZXOcFiRnrk+CCT7Um1aAy6sVvPOdrmxxhtnpcoXrXMsM1eveneTipR
Lhjd1h5i3fZAmOHpVd/rpESqGDgVPW0FDihY6DDpgSP/TluYDqbmLtpyz8GW/mv1
7JHZzFAtgZgfC5cETDOM3CkAuaMS90i6hFrSckOxQd0qHNpQWFHnPPa2tFUFYLE7
i/rqlMI0fsAC3essV3KB/yc0kibFHfbNMNadD5fnElOLPG7oE5rV9rOAg5Zu4JuD
p2hA8hOe1ABz+NoEKsLQJXRokxW6RTDGw/hW7YMFQpg9YAdKqsPFz3bgaEu867Qr
y93bdXvgLuyP9x7TZ+REDEnhlYFqkQYebq3faXWO0nsP8ffw/uumB1WX5BLdyBCh
o3lTngjp5n9hPvxKYzMnezZ3CsPTlbARD/GEc5stxDX0be54+l3MvNRgDX7+GOY9
3nkKYyL/kV/iBOksJ2pn8q2xW8cHDWuptC21NoBZm0KAbg+I6doKqWTkJsgDaqJ1
hiq+m1/yMePW4JG5S9AjcrMwkrnjJrwDDHJU8yJtSHpcjHpss5x7m3Wnw4qa7fVD
K3zIsRUFpTJRgPYZ7HC9NM/pFf+e4+0NSABbn9LjyQRcSd8d0IN6yfGJQmI4YubN
6vydNPI2KNL4b/YFm+z2RSYzQYzqaEvaaYkCt91qtdScel63PyU+a7Wk/0EovNtJ
4z27Hk0D5O6jB4iMpip4reLGbvKu2glILSxpV9Q8dowAFkkbv8Mn8Ly2RUD0t8Lg
loKSYUAlLNj+AycHGQsQfCLlEtj7qhilUmzv1TaNMtByZ9M8++/iJmBXNH9XVNSO
esBCPX/9cnHvaXNXlhdzmiDhWQD0F2kw3lTm4ecHa0kjFzfYRDmX/xXPRi7Tp73L
bNNYYHWRpbSRGgK5lfAnGxFkuy3mxHBen99thsc+njBYOsOHVfYttalXAnSq+iBM
4X6XNJOmqeFdE1IHkrPxolpVjV4dymYLeqLFGWc34SnuNp3K3MIULafIs9pMIHjL
4gdhIxq8KyF6AjRDeIXF2ap2JsjICXjrHKxBiJF+3lk8a6hJ5qQroKK+UlgL8cUR
ghcfpCutEMDsyEqGIlXCxfBnBCoMbuPl9XT4T+DRDomle0uoY7fFYuaTLUK8yP79
I0V3jHpeKNgge7a3EdxN5BmKIPse1HI2S9TUjo44LYOFhRNtVvEZqaAuMG1240Ym
pDI3ykZqk/ALy/SLhtAFliCm4Ya82G4eVAh9und8iegIzagqzG1/eITbNf58HXU9
wj5xQAi193KotYwHKLYupNfvr6CMBS0k2o/j14MTnE6n7hNXJ4ghVF7JsyN4dR6V
mmfTWcGuqV8jZ4csX5CEX3ULdD6S+XBX1XvsXClfFNwfQv71Uze1DFl0L+oNN1k0
9mCFJgTVHydNjPQXsnAJWoK6LacsBnA+gcHvhe6zFbN7e4O/VOmOdj51d+Iodsw2
jX4mqPZ8Hjvfis2QUg+GTpTG/hCwgOtLUiDIBUu4VqYaAM9Uunul6ecB46MuVy0C
PgKtcdb8rMRLS1ePVSpMlOQGwLx7a6gY5VGWruKdkPYc9Dntd/xBBZ8GWhwsJWaX
Wto6QDovw1xGUFWBVZeXrz2Xmr3v7Qdf9jfv08uMJqMT+hCEe3bx9OHDAXRYYh3I
pcL/Y0+YMZObDOqRu+Ow3tZAEjIi4cRsHe3a/C/hBq97y0AsX/DXsmkgSd3owA/b
i5d6wdAdZINaBGDpZN4MFL9bgLmJ0vmRwT4TGj3hfSXK8G8+jSjptCNKcKi3RiK9
wSmhOiEYm62/ZXCaN24FzFcBYobMCeGC9Rp16q1tSdpXRoxmraM3fXFa9WA0R8dL
AhU7rmyUfFZvJh8hCccZeXa+b2OSngnEe6HA/NY49D+MZt+FENylKFxitiwDhUUW
iLxIg5djqNuMXOUcyPk/s80VMf1QhG51x8qXI/Rc+ygD4k/Nu1QUwz4/kXfkuJy7
l61RsQIoCZuMu8Hqy7tvlE/uvP0ladwpBW6mdw/OWOflCh/c6a0nGbE5k1iC9+vY
/aUsuu1L6t3Z62Nzobco2S9oNJVJf2jkteKXvfI3j31ECEY2N/XOhjpT06s/WfoK
3gY2pHbOwjLWonxuv6H91wMxuvuQqTZVgPF80+z97GWBuly9xRHB45a7ZPEvkHrh
KQMg7dR4iZzgD6VdOcLzseH3VK6GPP9gUziIaQM5zJsEDyk0C9JSAboI6yJ/RrrI
4r4WeFdKW9NbfeFT/IsfE+3pr8x5l0rz5FKnMX3CyHVGZznQti2cxQZFnb4x3t2C
yXl7BHUdPDFGYwEouf11P1zU9VHIenh38d32DatdjulrUSA7T84zVOQxUdCejX3Z
qFr9Vq9UpMY/KYGxv8oIAzHiUOM4KaBkj8xlZAKPsTyXl7sfrwvS/MkyKYPKuYUu
rJnx5IM1+SZ+iH1Naxs9EdDvEtv/CY81i+SPZL/r/+YXUCUUptcc8RK1EAWh3+rZ
BjthbNJSNRF4vHeSXI/gwTbXTqS9bfrrxK7DxEF8ZL6R4a6rvSFcpRxdi92KZ15h
kGZEjnFsjPgfWvWBd9rK0/6lCHE8OPU2A21v4adE3dy5YCWxG/QK8ccuP2eeXDDH
EJn+Brjoyx9Z6uegQJ7H/VP92YxcxsqL4MCboHFifNsFkzcFC6M/EVhhENVPQC1W
0eoaYBZsPoCgAcmX9pGh+sRLLpWOTGk76jk8FaEwBdzI2ISYE44stXm7hTV8eCJ1
ZUiZr8uq2AB2vOah9fgTBDzsbvgBw+hq8oMC79MVbTs4/ntixVK+2nU2P5doQkaP
mUgJPByybsb78DKbevYca4t0tp09SJXfxhWsaNsS8Lm1K8ac+LSIPUmju7kOboZg
BKydbuvYFot+VQ39MHU6xAy02wkhuxXo0+C1NPVwIML4ESeWADLxAhuM3/hM25UU
JcdT1beoCfLJVGBofHgmSXS2d1yL1vtaxHGs2F/JRuBAThKYc1i/Kxd9xM9OgW8s
a5OXj2hubthEaIk5hB3v2YOAqgcYByFs+5NbFbqcwLYJmIk5QNo/BU3nHHQ2ftSO
XHU4JT3PoI9h7YvZPDBMWgE1slC8qfm8za5bo25zv33f0gjRGGOOoDMBpiKOx2Xg
/duyoAs2a4RgKuU1OpbkmOUqvmkMnyFcU/qH8cyKmyOnqZx+nl2n5MkzjdMUYsPf
mfwibcZaxZbnUhYVRDRAvoPIWIHu6I1+hWsb62iQCVZ1engaMkXyq2EtWtg7+9Bb
4LJeVa0qeuibELinlFpa3YfGNIF7QRucmbS1QXpJ1af3Cy1qy/XdSys+v18YTAd0
1N0zkSF+6usacogNOOs0VATFiF2QdXZ47D/RknBbXCmmR7mcDKycRUeesB/FbMB/
2PMQvxbHObGtokgD4UufFvokI08LW5GHISJIeLH4ul9D/YRCcjIAl2tQJ7UIlJIn
VaiHsm8L5k9AV3vpwtOhUKfPzrZYQRnPhBuLIkha3IgGrcSEsVkPdtOgLPrU1ZPt
cWHcidQE7Uex1I4v4IXJHnLQmujrnSkCG25n2WibOsuIRju5qFYoX7pusxOIWYeD
+RVWA6HjLb+KgqK/Rt5ph321um0GBzw8TB2KbLgNzzdYiismz+MvtvUruNO4TSrP
tKCo4hS90+o4vF/0B5gGrM3vJsiNGFSdZbkZfNKkLst2m+U1/pcVCRTtPxQBt15X
GmWqrASM2yT+IACwlIxOrmLjJYw+FVP6ECT7xORlnTSjpYAUxxI/dT3KnWp8dJUk
PiT/SxjXXrJX4qcR6kruSQ9dALf8ty9GTg9ye2ICJyqe/6bbJONS0F/c2t51njg7
OqpX+f2CdKAk20Gnd+Wyls0QiRdag+BK3BkCCCFCH9BeuWckhOqWvMFJrWz6NsHH
xP333zZIb8oeT5OPitw4SEdPy4HYt/Xgo3WfvpASzHo9alm+FdbNowx+iBfPD1X+
gUMpso1gbVEyJRrnCcW0xLw/01+VM5GLxEhOQuZjdhMv4oVlXcpXdIGaG4eAr+Kh
oMwbGsxcHZ5u+mA/R0DLXp5v62qf6FT6xuoioF3UcQsJnwen3jc9uk49pqGFrjTq
lKMtVrkWzhsSMzVV+0/OGNHT7Bxy467j1VB9P/EvufjU9+/R9Lx9WgrY3n7+JuHe
NAz7MIH+OmIgQrb8tWsev2jBPH9mPbmNFxbQQnn370KDiHKnuSUoMeqnSLN1iV7w
1kqPCLSvcivla9sfLbIda98ZVQLvNGOjwz7y75/HPvFgN1eBBgNZUEyDYtWP4HAU
1bNU7SdHvD6q8mIQuNtBxCcISxjYw+WqZP/PUgMNy2QtEe2Rq1A4L62/9MegZWBd
b+aCGGdprcc2Z07wntas3D4a46EY5N8dpmDUOkdjvoPmJaPehhHDrSAHJ1OsCdsR
jdprj3gbhOfMTFWsyLLAc8rBNWZEnbOcc2oZkIY49G2t78Tl37zYFRtYO7vpwJL3
NvwP/KMQr//y+24TEkPzvLGc+mb6KDtvU3171K6ltX0c4MQEffZasmB63+erxg0u
0Nw1tsTfZepPJP1fgKQbk8Uy+4Q6OXSPHbd6XT3LMu6HQSUtgxHlcBuiNII4B0vj
gkv7AABhX/OeiBEYr5aCBhxXHDAiVXyOz4qhYc/06t/syT/hXcJ2olOxPZDZG6E7
kd0K0p9f1FqRCNbkQyCR2HekGtIw5O6MWaF7w0OXSTvP8TwTkzQr3Bj3ms8Droi6
YxWcsqWYmuUOKJiC76nXsPeXpTi2Q/tQ5OyRcmyq5CccTt2OMnanNGkgAGkiOvUC
IWX8/dVBAFIg9qBk4Sdeb/GLds0QHW9ZcWHroM0fm7+ymWl89ObMVW9qWY41g+rq
yZXjcB+B5L0AkC3TeGS5a7pK74s/smT2lgYrjjuC0KgLRSz7s9MpPxzaNhPiVng1
npxDHMl/LZez3w+WzJUHU/7i24OJ9vXTo21+Bp1h+1lXNz3/JWFmmSQ0KkucpmRk
prcvpuRxeSJMZhUbbhCgPbPHaKjdRqj65veMWXh0weaKvlCh6jIRYHFuvfcSbc0N
dDSByTS+UZNRTEF+p9ESWD8fHiVUkGJCJi4UXcIbtKUqB6YpS9Zao5dUcSLSUKSL
oc2gx0d4Ub46AEpNQCKaRMiXettkqwse+jDl+/aDh4NcLh2yYEIN0cb+CP2zCtOt
Cj27Bc1PXb+3DTr+zY7S4seRBpRBzquEdv2T5WP9J3wt9GScfQ5SMtzonYVEnfrj
hhnKIsvijWn1/ZWY1yblSQTFVZLWXDcJBgEDmlLxs1idWF49zSmMWMn5i3HyaKEe
oVfgJiGkJFEdZLWWFJOYElxKChM/P7b/4o1rTNDE8wRykInXUZnXKV1SamNKf+0C
K0oTvW7O+/PfHhYGBpfZGW5HWDD+0YfUtSuO3DQMuCeuv9+k0YP8qNaaePMdeUQB
BjoKmF9ICU/0J+FTiWzYlhWtiixm5wV7iKbmwpkTpUCrx0PZSP0uxiP723Gm1J1W
9e5iJj/+3D6wXdYzJobjPVe8j1oCT+Za2KTIuzLZ2M+nbRO4UQSaC2z0daI2lzac
byc1Li+0bz1i0tkvPFZmMwea7svz3pEXX00/oAfZ1061YXPOriy7ueRpCajZeuXP
m29xwIesi/3b2YHRoUPu4xqS9EwnwOtJe4F7Tt3/k2tlQQV3L+j5SXFrJzp04bzD
e6usISOA0TIimtBe0ohomtZ2PtoQO7QBUBamjxfJVkbvNxO2OZSnLWveCXmoU+ep
ArrcC1TLBjTudW1kV7aupVOAqe/+2fImm4D4TG0Bq/2aZp00+8e0aCqBd6rf/RGg
XL3QN8HDn9I9cT5pIGnjSiOZRjeRHEzU9Q3k4T9h2uMBuzsbiW3giLU7pgvbjJTt
LebwsUZoxqpWEaw3D6VClucDyGKOGqGcoV0YaE743cBs4kj8+TKSX9zRGxwsWhnI
2m0NzemXdkDyyjcd64DSscA9n/EuScRn0HcWZbqa1bz+xdJ5LW8TNcqllwuiYLzU
BObYKNtZnO0TklCSKxBBzaXfNk2tEnitz6nsKyYQ7P8+iCSrLC/nVXAWgn4QJaso
dqebx1fVprOSOvpN3xFPMrq3CpvP/JLUkNSqvMWX4zy06ZjsYFmjr5tEUiX1x9Db
r0LGxPrv+Aa/1Mw2u/A+uGtADVni9edqg/fQ/jtBf0wxWITuv8WbNmo9lWnqtV6S
wxnjjSPrRsobnUkA4NvK75unzYzFSz+XFtSQ5pTsIty2n5S5cRrUOI+HAmZIrbXH
Yp2bAa2TyUgzpluiUg64HK245Ie2gcsQ21bpWAjSI1iprJ7aFslMygF70Lqm62fT
96Wb1y9VqTalYK4Gp56FMHVy+WbVifycHVEZtxudpu+elMUqDSUBlJ5AhOJI+IN7
Z1lk/Whn5asujVKfOUgGBIafwqFW/XniTPjarmSa1FBL9TippYNTYKuQAXouyXlD
H31JFQRH7Ei6tzfmTV8RiFmkgkhjgmKXcxxXHLTacnyBMeNRyopS9qjm4HRhJL+L
FNq8KkmeNRFMIona+EeCwqPcZlEyVkYyXMTrKMzL4HF9K8RqabiT1pa8GX8OJe6u
JnbgjyQN4mnzZ86V2aWfXP+Eq058K+z32PoboaVCoEX4V0UL+OaHqcut1ryzUS41
tlAD+0cy1S+eVHsAI6NC8q89TqPc11xJKEIZX5BcG7gGvaplGZYJ/5N+1xzyIVGB
PAcVOxGdkDqAoMyS1ZZ+yz5Vstv3ll2CNAQjERXPhPzbyVgd0VwM0SDeC1xoH5ZB
7UmNCcvmSU/mDGXVO1XtUp0QsoXzlibeXpNspGRn0d4ll8fRxP6XM5D7PLJRP30E
sE+HLvpuf2J4noX4lSK71viJgn3B5Byiq1eJyeshHvseXvoktYhTzdD48OT1fTn5
s/kr5X2vGW3jN0K5X0uix/eLCjaywFS/DlMuKl8UfvwIJoMCxMHwvajjD6s5TdzS
vV5isEZfxGpjJSPJBbUi9jJ9C8lxSFmWDu1hRzT7dE/dqqp9MlV3Ep+GeeDzigym
TDvFIaT4P/Xo7QeeR/RlSZUrBKEvfFGEyVBAqfGzVOHUvxEADKEm80QvPTW+21t+
xgj4U2NBc9PA6zwaWXmhMv5xsV3OMpXk/yayl8O/aduJeoEHn+sOqx1EQqC58Uyd
ct1wXcfrtD2yJnLF1IScFV4kzPYxS257fyHJDMFCcXMl74BVQinyERiItpfwXtUU
MPR3y0i1c+QSXr9PUAFg5MEvGrSZP055GmPTDaOwUrhPkjLkQhQB+pek5WU9bPPA
38F8cGFCUcFdIE3pMI7AeqaNkUMISWJMnAErTweCdfb9ezzYB5Zw+C1G5Zmz0ri/
ikOo/ff/sgblfO1e7wCZpVQ/iPebhsRJ6EsXK9HTmpqMcNtrIvMUm3XUCGl4JRKR
Gb5wSOrmQluewWZMNMLZW28np/JZpT8PRaNssjk8FUGdyudDKzM9d96XaYMxrZyD
v+dMqCrIETY6uygiK69WqBaBzZTVsVqQECiDVJHi/f/mvwJbKQ0f8/WjlPTvUsXm
6HnOP2RliZzLVPFG8INCoxLkQZw0grN1pydHbxnIAJdkBvciMUbfZDqYbara9cpq
ivjydGsXpZ2E+sQJqQg+T2kbWWxekeMXusObb+3tiUt7C/Lal0YQ3WzxmRNqY3i2
sgnx1/5Wl8ye0R6nxeNBp4vFH26ZGeWM9+f8XtUsDhSxF4rNHL2nHN4Hv0QC6LvY
gawHWWefvn9IKqh0mGyvkL124jp6BgVs0k8GlF/2y8A0rpSoGUPihh0a5/8afGjd
6fDKKu0dqQRTFgXfB6IZt9EAG5NbwEtsH+NQ0/79dC35S8XMqpxVaicRnCJfEZZl
IOZ4vgPK8MGuOIOCjT0UiSZKl059RkvF4n8g8BIkr61fcG6FVbH1t5GZKiqHai3i
Gg4Vyw9sjamJOxFifbbCDmu4f72Zw264cXuerWerfA1OhEG1kcEodQges9J9iFVE
c9JZa0VARqyXQRNAVwAgiiD9bMcyz1gT5uDTv+vFkYkK//LltMByq2lR2oY0IQI+
PASSDN1AMLG2VoePcQfgPKP9IntjGHZNjmQg0UnysjPyAVyTrHZEED4+FIo+6xVU
AEprvPFh8ZFkUCdEmYndS0R5kr06C/VIlmd4q4Mgc5SZpnFU3gvBdIpnk/Pj6YM3
3X9gs7HBUvJf1zrOXKqaP2UQrG5Tay7VhxxLXDeARlwFFjrEJLbisaNyhEUKPar3
3K4EVvd7CM8Zi1CuwzAA/OySV+fr+PS2gG/2HARYlhzVMeJ5xhOe/yh+L4juNGJv
YuXmu+IbwlH72AM8FxIMh70sZ8IvLWVfi3gjdeZ0l0AMzzGg4H2p8hGkNPgLcuMT
+jFR9BvAtQuRWhJ9qIAMDFgAewg9m9MY4pXY6uc+nTqfaJdKDo9nAckQPcD/gZC2
3HMsBb7YhVYfNK0pg26r+aZLRae5FQzS5xs52oU7fme2XH9cyudgTbRDZXlfnU6x
dKYDhrhIorvYDs2WOdQhq5M+28CDnGnTtJoHCu2TWF4JHeqAJewxJ3gOM0vpre19
lcozD4WEytNzx6jZ76/Ov4/WwOhwqQ6wp9mcZ1Y9egbu9OL/cfFyo8YqYpgAAhKE
WzExmQtdwQ3g9Ip8Cqiw6QJ+MmJ2KsvQ/fkhQXQ47gFOOu1O7lHFs/1ZFWdfKTOS
sEmStUpZtbc6w8ZPETCpqQWlWCwvJsNS+cArys1NmN2+1G5oj0t9P+GCPkoBEi7C
sxWs5UDMJmw/zlG8nZlho2pjSE/i2iQkyJlPTV2h4gKah9gyvcGFZhsQwkxK1MDa
mfwfN2qyrYQVDgD0yPPF3lejTbdsvsVquFv5wZzJH5zSJpIYW7V++RsSS0J194Wb
O4h2VEhbFtZtdrkRVyFNbUTnS95eaNcZst715ooJUJATJ5lRVBcqA6VXHNnRAQ7H
cztxHtA6dDSXT3tLdBtqYtgur2ULB4oK0ixVJkwhmM1wrzS6sKpaG/iOF/gJlCXs
+fZejOCIQgvSXXY6O2EisC8f2pYjd2eGuPsC5dMGPiNUGiT2Xlp4b9KtBefrLDWi
T3a4Es8IzxiUic2aklmzqbplXm/LpsbrBCuDCG2i06za95cX+9mUURzJN1psxPum
mwxeS+DP2lBd+PsIvs9cXJtJAVa7QnGD1UptzfYkQeMnhm7v2pDvH0FmoNgk8Z9e
Xz/pjeEy374pB53DcsT68hXrt+39K2DbiBipfgKDdYxsuWkmexpdszq9RtzEQldB
/sak9W4IHiTxCPeF35Tdkh7LIlerLREC+At6zjnaBkym79kG4tIO15moKB2ctXVY
YXYqHlr8WrlizSRpOrcEN2kIFvOlQ/dKIn7u0r6dPIzw6QcqeIawupk96410aIVO
Pv1gaWkJlZF7t3MC4R4ZQrV+vjyEPb3GM+USHX3CVuOaMoFYwSXPacpf0orK8NRb
QRyfwUuRVR4YvPEUTLbY7TtPrbJx/LKHPQQ8J2+4ssT60Ajc+M4cbhN4Yc9kR+29
hs8mk2Hkh5eOdhorWtU83+DCeqiQ7ukabSb0U4keVfb8Gh6HZzNQg+m48A//vGOi
O9A9ldJ1bk6CSPjQz8iGr1ymrAu2uCYe0A7ynSW+QjHqZz78TB+uTSV8GBKeItN3
p2qhLEyMhW1mseJRY/Uhg7OVxE9il1REtg17fts8o9C3u5AwDfTTWRYmgrDM3I+V
I5jNmB9v1TEZFUvWsNr5JMM3CEs99c1lENpQMhtMLA2CUzW5oHc8ZTy/KJasPV51
35EYSGo7N1Tc60yygp+6O2y4iziRRTal3Fzy3SrOPPXoCoVRdCXSZkXVn+08wzxQ
t6vF6ZvTGUViEVG9P9JD0bAkMHujG0sOEJjZE+5IJ0fX7uzCIdkn196D5OrO1wAC
PrjQwaxt0LEP+sQk3/viyjcTq9HXdqP2J11gaUz2ZanQJHttYnI8hJpVDFZhXrJS
e+V6roiTuthMdreMP0seRSveiLVkvHpK4PE6CFqA4OBCPHCzQC0uwTVyrDrv7N+/
SCHtwV6mOYthiBAbqOZGIzDZ0+2q5/EMoT/54RFkYuGBrhmvmj8yZD6iooIOqmNX
pjVrk1RuxUaho3BIpBMvS137pxxYtiX6kuhqvIeO0lW4tChc5FlhD4WCOoWsKLRD
mMN6UjjiMs8EYEX5iD8pDiYNzYE3PVsg2+v4iMfd43gITTylzURIOYlJ255029PP
9X89Rp9Z8FiRR16DArtSpV8sLyz9eyxOc3hrdnrl/d6sGS6a5VGsLP8Jd7yHt5zQ
Y6YKEYRzAzUeSOT8/T/7Ahuw2g7x1+n1cA4D1Yu0LMuraQJQBFinoL/u8HB7bMlh
CvDiDp9zjaHakOERH4cXCGiMTx46nrYGSvUJXWTM8gS3LMo7wygTKDfd+oQxMWio
JLu/D6mQ6Wn7bzdfNuS0rThIVZiB1lb+mkePeFB+pj2pRAy40ZfoHZjzSqAbMVob
H/dOoeNh9wvZlrw05ozOedgfdzpQqJkjbcJHl2iUR7VBNWUdshTNJ+OCUxyMMp1D
tUropnXLIBxMbhzsMv9w00+FltECA4Ts7T9JveQ+576yFTSZRLOM2O96NAtnw0Or
tm1Pu+++OAi8xXl93eWsiFZAYJUqkcRkmgoY2wv20xEXtYct3cWnX4H5pCri3igJ
TcnY0RThOFX6MoxwEYvK3mlPVIoif2yzt+OREzrdK3BB2S0q03x8Mg7VACbdore0
gQdbh0Fmo5TNNHfnRHePqcuFnIMmYXuIqEK3qlmXvHINpdTc/xh0VVx4snDUscxu
4DGRaa9dhMlE7de0OGjVnMH/JWhYS78qZQMqDwMcpjeTYS+tWtT9iOnsX8w0W45k
Brk4Xh2T/ps5x7fwDNInwsd1OBGlbk6x0ajVNi4sYEOrPVDH8HT79CdUq3iGt8jT
X9qX/+tmzzCyESf5zqHKrWhS6S5aL4rV24tScFz7Xd5b1OOIb1NsqW6shccDy/6P
xib1zi4DBGvNWs8r5DogiLYKtMmLGH8zr7SXSAj1P/mnOlNxXQQkMsNWv4X3u2D+
d0xdeLnXBgUhGbxkxQUExVCjsNi9r26ragqTkpI/NwIVslrCeNWHd/1t3c3tvXfl
iPRpE+90lTKKkLa2/RgbPr/7D98S+lA15WBZ14GCLMYMXz09e16IfKPJytCdZGo6
ja3u9t/ZbXfeq9J7dvR8OpagQsRQRDzeeGiF/FW8OyKFDd4UMxb5h4myAx213GuA
j4h+gAzfS2qfZiDnzfBKN06UMR66HyBcot5t4ne3lIsA2WUjeaKuvv3nQgwYJ5kd
7sFoAaTrBg94akrRZbuHererAFStQujqePK75txtphRfNnV7P/X36wFpb2DEsZZQ
FxI7MG5Upyah/Q20JZ8eGKP9dysSfgFrhf0LXEHLNvR7NR5nFmcOfExNWeuAgFB0
FRUNkhUatiKRsHFHoJ5R9AXOkzZCygTHF3gtV7Q5jsqVcWDbRePDRWaTft0MyrOn
jVwtrs/VgYBalXY41xtoU2TFYyARMApIqm3VEXAntaWBGdRv2ZGoB/ZJk/1+ZmSD
ZfXFYsmlIExhW8DEtlBqaIyPxW/q5hAek7EsOXVRb0YApE6QMRzzWGLb4zfIqGpB
j+Hbm5ZE/p3ut4eTSd+vM5rLv1Mxh5zwitXzigmUFl3dS8YDY/8gVE05VRQgBo79
LiTmY/yLWA1nl2pBCsM5QkXCe/kkE2VkIwhDXV//MRJ2o68D+uOHIq5JaIoMuF7g
3ZRF07YW8jSm0/mZOZcbbTeRLozdReuh0HO8foJ1lY9Iet3SFTSH4Z/obQK02PPy
sHXA33evuKO2ACFINCWIR/K2kCpE/5sTrfSwAnBvXvmQL0EJr8paDgNppjwI99Ac
C/zvAFBZOg67jDFd4uTicMmmJqWm2de+AYi2AFVrhjkV2j6j9cqYg3a000TM388P
tdzoSmQs6CEaBDet3DT44dZ9NEFz2RFqbS3o/noVHGc4Fxb2LxaNrfh4CUybjdO9
3ANhmS5v0UEUWb1YtG9gFM1vQoeGT7+CDsgMkKTgjcU/V1UMS3l2YDt79u1ne4Ua
cRQE97ozq5JOYWweOmCSDGsB3dws+oGO+N3EIHgBrIWRQpL89AW5BKmXH2Y3rmaC
JDVQiMUJMEaYdKv6wl5dhHPe4ERYynHsotNsPyQhVNQp/VT5Vk35a8P6RBXBew1q
BUjNYlVkeYUnTivRewkscmipy1q1JzXO55iFN0f2ET6Tnk1T/ItQFLBxc4gcFizI
63grSvJ28ute/6TQ+PyAO0JhWX+sxy/OqO9KkNgB8ILxPxPRTjE2p0K6hCaOmi8A
OybVTiYzNvGfkqGdWh9qi8KTcEraa8rxvdvlzYtmboN3qS0GDvxyiIGVZhfyczbH
Wf0MOHjOb4Cw3TGUD0KPCi/HuiGYdebzAhw/o/I/XqvLi6b2p0DARt5sDUq+J5UB
s0N/p6rQIVxH8LwrSBmXst1hYNDrL1SKvKA/OW7u3Fw60HMiCGR27aLZpmXju7Nz
8UA9aGLanijqqUsYv+mbkrM2DMo4dE6MB/PW+NLtbp9XNtyu84XMq2LKTP3wO097
Uspb0GWHf8QKQFPTEXddwialpWpWfjq88SeinZwBo3fRTTFTDG1q/Oiphu4HD84w
e0yFLek2OXyucEPDpZLwuYiwlxXtMuRMY4lmj19+LgksSrbdpzZjXtXVRIS4TPZH
oH1I83Toc1x7nBeVWOwArIOKxSKbYEpLFWykQlfeKd2WrhOJvcIOVkQR7vEMDujT
fgQf4kjurhrR/Du7joq3dGA1x8p+bJcgWXStv/OsjKM38abvXNNhf3PG8BDARWwk
6Kj4jAOnCTsiMdQBwX3fHKVsABfVPHZf7SAL92O8N777YGxUOmVEhmra4VPB26jc
5zeo/Lp+PFxT1qIQxeXkvrDDx1vRk2RdZBbDceaoFE7JublsyIULgd/m4QjrWkYe
ic5dveYSKrNYGbK4DElcZ3bjGFGw7XGVuhReWanJVIKntuqpF8K669o0d1E/FenH
54Q+RXgtdkxsuIzHpsIPtsZk6NbKvFUqFhCSRfGuIcnvs1FD1yuo44i78WSTuFUK
KN9uV3Eb/xd+ylUOR8qxL2tvYk0PkSOsbHZV+tUYl1Z77j9YDBGw9oqjnqkJzdY1
+DP5z6j6BpZBfqukJZg79PdnHnh1B3OpEfYgi9ptcmPtQJa75WT4mrtdgMgk5ee8
NGaUcCIBC4UTqeejg/ITsF101pxQCXqBpU3TaF2jpQQXctKIJnyjoiapBRQqdwfb
CSq/jchFQoMcEZsuF0c4E2+WD05h+JVihR6VjAwD/GXiXtlpw/OLpmgN/bjPiXZr
1VJ5I4HdYg2vj+6vPJaKspBto9Hz+e0nyv0m7UatBjWAsVsJ80TlnVTTUzcPmfeB
0wSWKcdlIhc4TtyAV+PEi7NoWL7fT7hv42sHjfmAWKsC45vyCM1eRGcebQrCC1UX
WiFTM/SGdOhjpoqg2W9TdfqeY48uq8E7XecJpDjkuS6F4/znBoLrks2Sy23GeKkQ
0MuoU333/sSkBFib/rG6Stegb73YMujc0xofXAqTQNmezjvUGfGtvsHsrPCVWmSR
0EfNcJPH1cm+rMRUzEzLNSWlvfkQrsoSh/p6Sft6sWSdAb7a+oSTgLF1gbG2Y7gp
ZjKEJkaEvIpxrHg27vZY0QGnnevCIO7gnZLjExg6NCx/pULs316ciMsikS8tfUpW
16lB0TZyuVZnMjQN5TM8oXXgnj5RkhRJyaV8HRuu2ZAHP9XepQeMkkaB0tcr8sT6
XnJHshrJ4wsysozJcD9f5Bf842ar8e7BBmN9wKd82bnfJyBAUPr0OqRO4NvMBJEB
6FHzeHn/iZ9ypleYNHQnXETdDn1uE8zWm3kXo+HSipDayW62koNI1T7kXIfx8iFU
nb/4GLKMfODNUB+8TGlbfghRxNx0sJzb67pP6Fb2ebrm80Yiusyh1RZq198GTmIx
txruceJa2O64EgaJEf09RHCkvIR21nWbF4IWzsB20yCzN9653R28lkfHypcrKmn3
RRfueE24jGoongOn5gKNS+Uoqx55Br27cqWhiMn+9g0cZXdMbc/2G/q0wd8rRbi6
SzMwhGXoQWXMiXgUOjfmsX+y0AlFVG5AeXlbbYQ/WtfJLngqDmhMH0oXTrW+bJhR
jfvSFUWxMmkMhT7QYNJOmCxWVXwJmELr7F/HPmucHJqP0Y2bWX6r0f2+8914Eukb
AnvmpTNCA9xrNYmQl+vd73XaY/TbJwFddgzLvWHMXeSWiKf8WZDKsGvH1hfuOfXb
aqo7RFmBTobisccTw/3mrFXlU4QyItXvQIe3WRDY/L++UWx2gpjePHCivJ7cibmE
kFcL8tQ587YOenoXNvm6Y/5sktxrsNXO44aHd108qx8TbVsstk1vr6I0C+c98ZEn
hCaqm+nO4CFZCabScbCrF/v6X1Cf8RK5B9yenk6VCiERJBaDFFrFdsRhZOCcUMFK
VERT5y3aXjJzA6xyAssiiqVXc+5W6QZb/biVOEiNlFOIg7iiEcJqjtqh7TXcCwwc
NTzCTwcSx4MMRLHKevij7dVN4fAV2mrz+kd7sUdOf+o1AwqCdPZJWBISVFRGiJeK
YPx4QSbp+Fq5mMSL1LI25KAlVn0GdGA5d9su5TYOIWB+I/fOhhHS4Rv+SX/s2ByT
kHykLDrFuwq0Br3Oit/hHF934AQ3NRRumkKjqYg/wRPWUl3LyOTmwtVR5oFsAsXX
pjzdn8Eg0PGoGRnb7CPkyrF/tkqmXhaJBidvwsSFo6jll8FG9Y7o7ncNJbMFSlHN
5dibtBKNvTzx6PWhW4rDSQCuKJRAt++EX0GtjTQmaQwLC+ciNpxxwmzT5l+Ibmtt
1tvgJdrDT0QoKn3JzkdKqljAQ5DtrgIua/et5z68bhXJGQOfm+a9G8ZcolF5zxxc
FRNl+FzxSsjN4dmPOi2E0Ng7hGjiT2sMA4aCRZsszMrUFqcaSjXk00fhM3i26cF2
Juh5t35c7heXDMmJ2eYKtCK9go1cKMm1TFBMU0aT4qkNM/R7cHnqjpVOvTlG/N05
Wqab+AdgNh/Krd4suHzpyM1QNXOWKNPd59Dui2b92T5vplXQSLDTZYtwbZUL6V1A
cPyWaA7Vh9yi3xpnGQpA7q1HFDX8ZL2huj4JNDqOYIymFI27gAgsmWNg2MDr3Uge
NUifysxQU0+lUxps8u1DT6FynbJ9m6FTtxIy45JtsFsPNAwT3Rhmsuo0kk2LMSgu
o3n6NDhgli0ary6fcsm5A8m5ISDzfLyzSQ++apFUEH5XlrdW/cn8DwFzR0NWJsPo
BbysZPsf+V0CaHFJdJwBTtXLkmG1zQeAV7qJOdZJzh9RrnIC1jCke1L++lBMGqRF
06vboSUIB5djtISlD8NZ5TNe/zN8sNww9M80V/Lw8MJo1afAM44Al6NTnIvyOiEI
4cezHnI9RC+X4IDAq7PlbhiIPIiW8TtdFvHua4oy3VqiNxvhCW95ZP2Nf/HKFHWe
LpmenSl05B6/u4dH5zsCzpdKylLAX3BJiU8b2a1tIOrIK4V97ELO04vehmYNBv53
EQjIermGyf2cH9VaigUf5DOqQ1wcCF1Eiizgx4QrQ5ADNZVvZacs4YlVji5l1RAb
TeY98H9XLsUAvXW+7g4BUK5n42jzHgd/hQneE2jNB8g1Oj1vZxspiB7uj7b6AUNv
7Czq/Ec7HzmYRjKEnGyJGfGfYM3TLA3zmnJjaLagEOvOM18Uc7OzYCeCwnCVACuv
DVF8Gg/r4CaLAgTUaH49hhkxeRBy0UBjfc3j748x4sFaSZJK74Sosr22+Q+dl+2N
uXv/BiU3Vb3+NLHPQR0doFDLqL2PryoGaJQ5QnXT3XPIMu8fd7zzlLLrol1I5PCm
a1lbBxOsj1310NHTQ62gWfqjorhPrlP9Fg3Cml1W3azD8mx2ZyrLcKu4+QVIJs5K
hRigylsf3J8rQpNaYtzc/saSG9utV2Pge0WPR8S3I6r5ky5wqH05wfmVSGnbWe/3
2/qSVaWVx+aT6+y2ssYQSrsGzlsU7AhltydLolxv3dQsbsd8BX94CBjypb+/44Rk
bT8sS1oCqcW+2NZU9q8n4u7YLWaNRMqpTGBS7wt1XlqAvokS2oCW1AhTqF13sdGd
0o7exCTNum5MsxvYmM9E35BLpcJq2bpVsUIL4elNm6ZXBKCOBpfTAPU4yZTyZ3z2
F+Njugz7ZTZwxZHQJGBr1XZ/qjzQPv0Iw0XG3L0GUgfEO4DYynWtzewLNrF81idr
MPc8hib2L/udRp10zMM4MQ9stGi8Y7NQJV07Cjk2lVju2wtJO5hd0vIjyB46RXJA
jXtSZ3dqeAPQeoaZkepa5LeSG0T60KgTuCkVBm7pDq2nyqPe0+ZZqeGxNQvzT2EN
V8i/ZhTaClGV8liMG24NWNcbSKSIcAWtWcm28gHWX+Zv+va5EX8GgodBacJdj0rV
im9e9q1sMxKQ2mUfUE/SGnl1OOtX/unymBvy0iFhTNRGxVXWxpAILIS6eW6F+tgJ
Kzu4/gxr6x89S6TK50pX0GRe8yZlwkzv4Esq4Bd7rKfEyRmSI9hcENnV1/TUyAJ3
spYmiKCTyxkX67Z1qwODI6vcaizCh2y482jYhZsSBej5vkPvwgeMAwHu9L3tf9tE
PgElNK+zbx558wax6y7yw3ssre3LxCdpnYzzlsq5IN6+ueIh7rorpWzFe1WZpM2y
I3bR1Qa+ycfY8/AttucGJt33fTLfWko+FP+jlVY8YKSrbAh5U9IFDAYVSYobCJEH
FcN1bpS1WK/YgS3arFJinR75ishy6t9luQF/OfR01b9GYI6UNeHYFPJKu+Utd3H+
m/5AVyfMnc703gyeYu3b5627hsqNI/OnMuJFOvlk8B+oV4Nke+96tZY9Kd0iBluU
ELnRhv03txFN8jMdyTsfNxhH1isrvsl08awpdBWCkHFFtbEMCaNVyyu8CES2vOu+
SQxovndpYiOk3r1NJKuR4IGN9inSGY/RSVrGG2JHEIV/0P24JOPoMudUWePbxQ9/
rzRCBi7CEjjWurZk/pJfLeecHicow/6ytrVvsjHkgRdFFpIUzQKUVNqlvpA5FwlF
GmncsS41wW0S12TFKokdqVr8PoEfzqKmi/Dlh/WeEtC5K8fnHxhv/mvDBwVZJLpm
xSA7CpH/IfGvz5+MtgrnzWU/VqFcWeF7xiNiq1kMyvChOPNsHyJdwyELIW9kn++y
2AFR0BIy4fpBilquLwttAxsPgbwT7caIuxK42ikU3x6TUMoXX/vlXqnRFhr8bbEz
/bIv9FXY7rV3XoRbDPIFKX+T27MwrJCinDnTtrUBQY11KSs+l2AjLQKDIr7H4xTx
vO+JWY5Z9RNaX1CsAZLbeFXzEzQcKldkrOnkng1B92Le+HAtUNN6VGmSpUXQUKNK
4PchXLrSe9RxB3BfVFYduPLafWnN06yqV4oBqLBSIDndTJweuCdd5N5BlnUgu39x
zqr7ryslzLWI0B96FoHPLI06SrdjeotU86vswn84E7KeNKcLIGD60BWyVGgaRfh9
2sXZxZkgKXmHbMGw8mjmBSkiE+sIgk7ObAq0iDBUamR6Ml7cTzzLIFeKYQU7vULV
sLKepYthILtOBu3eea6hzpLhSPjMTESM+RSc2urK1MfpbGm3ZLSWHzAK3H24V6GF
3Tf8zicDzeR3FjMTufBPsf6kcU8+zZ4rJ+fq0fwUMyvnFIt6njgIwgGR5+YOJIud
MzFHm3WxHY2uFOucbaYtHQl6/jXJo0fCprK0M4wZsqacKq6FleSId/Wsus/nOWlE
BXcP6CIsK4GWbY1Q6EgPEXoFVduLarEbaApasXX+pf07EZsIiXDADnAfKiFK9wN/
o2cCs2GGu0dSIVt/JwxdUp3s3h+keGAvT9iYZ1VcS9p+uR914aWOtkiKGiFwUU42
aFHL935FwmfKUpcf9WF/YvLMScA5JXVYhB9wRS1ZONnw+bORBzc16zjhBOF4ajf6
mSnlLMKAF29Y8IvOae0iC1sB4kfOv6Ue/0HL1nJvoPInGgtMnsD6XPRa0IhFDVfV
i3waNjg/wt1TQ0KtvwvkFe8S1P4lzZJOxdMWvpWnm22l6vPHyAD2mTjUSntjwS6M
xBQ3D+gtM9aJUTqeJ368MLi9RMxzX/ZvtdXGINeNe/s5u8zp6UO46mwt21ryXZ2w
KawYDNnGzpflYUnzhR3kSn4A3s0/1zh4s4gkCi9gyTvcuabOgCtGRfeLbtwiyemV
h99yvs5bAgd7FsUUAU95KJhUFLfcz1fzxP33uAarg0MWTVUZVpiNFUPc8DsexYGr
EgB/ci+Plxje5FNaYNT5l/ZEKw6MZbXhiW/1sBAfAJMJXrRdemFod4yXgZdpC6Lk
BkBB1WSoszw19+JnZXv6gKJ0f/v59DG0gsfSR23iGDRPvrVeLwtsQzIacurIE/EM
rinWnKt5ZwSQ23B+LHEbR/mjjnjN4kigYoUG7MwEcG1l57NkNODyCAFhonfFOqZL
cDRWmOOMRefcY0Dk27UCfoqlZF984pzHBLJqVce26NzMLWCLdwcCHG5cRjtVlQ0R
nsYP1UVra+g4N6C6Uaha+FXodt5cTJJXAygeLSp1g7Vq0qETTHtIyEP4G5pxLJcX
QOKZ9SK2k/sRMM6UqvtJDAy+X3OlNriTmFBDQqTSO9XT+otUZiqM75QT/8lup3na
qWzfkzoBu8MzCR+hkpUXIL7QQqt0jvjMMNFm39IEq9QTdZXJYYmEudTxaDwcD9nm
0TD4yqsU6CvdSrgOuL8f6faB35SPZ8tNVXSyjUG7Pj/K/gXbGFq0STkTa1OsQgr+
vUiyEAQUhhBmmCYXDB/1FXxIPHoltg7j+oeBXb8SwVLD8Auc7x9E8hx9T49iumnJ
4W1mJfWpmBQ1CVqkQJwTUBynHa7aTJIPH3a0hgEfXYe8NMStSea1xI2/Kzr6WXPz
o7J1EnOCikrmtdP6M8q73QYWqunY5U35hhMR5iyBtFn1B/nnJvmFkKU1GxbCatEI
k2VaZRaRXapZleEulUHZ4Im+oi60NcmONHbHwJeWwhaSkNUf6LsJI5t1euiyovQh
PpBlki5Rjc414UXehhnQ4O99AY96xYinSZ31OINNfHuta2Mla6iVOqysCNCgDVwb
C9gf37PJxNYPl0Y7u7/9vD7Gb56axwb0PT5zjAeySuS0Uzvk5kvG9o3dNPPC04Za
xbSsuErA3+66qA137kiN72tew4gx1OGYlSU8/IlNpram+uuYb6J9xRvu1zokuBTW
V+TmuRupO7R+4Q6x+qBOVhMr/CSiHnrFpMnO5tsRYMpA9y6leVv376ozQtSCv0NU
f7l/HAEAHO1GDXnU1rhQHYqhCyY5pEJSNXWdEGoFk9+Y5tAWEGmZK52d69IIomQw
9aEgMvlUBI+gu7kPbR07vgaJYv9a10AvMIafDMaWE57tsi8VyKg9vnLxMd0FYBwb
rrXRh7CdrpkznpwrJIVlWuQVGIJuYMzGzOi0Khuu6RNN1oH6/dekB1iyv6IkFk6G
6sry1T/q9pBfaYlb80O5Uzi1BHfcCgkiVEmdLMsjLjUbEqVlYPAOBNyrDt5Ih0RM
YuQVFbkqtr8OZPYPX02+1OGaM/en+QvU1japYh+ZGbX5gCqHC1xkXhv4egnCn2uI
E09MWNsjU0y101NWjPsvPELChSQ6+0o9RHOuY+0zpmp/3IDRu31NiecRgnBqRC0r
bxd1/fcwxBe3RlkdblfyeomX+7jwvlzy6tSE+7it5YIhl7DBjRpdQjHUcOvTixiv
0NFX9nmBvhX5VdE5XxD/UKwrLFOZH4l/JcjK743FXXYQA8wCPUmhEVLIiwwAqpQ8
tRpcjh/g69P3UeInXAqe87QOsGmqQbTVbKgVcqy3rkfdtSxs/E4TLHioIYQ0hgHl
57sB2YBEyfOgIutTPk0HRxmPbcnA9wku05bgaT+mO9vc34JJ4xnmEzKcxtaaZUnm
23u2x8TNVqNIMbmwWdWmRo8l1yZLqQa4ArzQn2BOzsTfOyulYpw9Y3chc/DRABVK
4u7HYR6qK1m9JR/saozIG1+jYK20QgkyQU6dA/ed/1VCUSe2g4qhCnJ732wQP8Qx
CFOis6UUq9LkPc10uNhgknBfAm30UtTevtgNXzlo2gaRfZ42MKV3GFQezb+773J7
wxF8tukO9cwzrmF9ro4/dmX0Cur54sIJxQUhcIsbQxyviRyeVffALvuK8w16RkmP
PLMlz3l8YbGAvOtn1Tcm3hJMwt5tYwC0R7rjGAy1mdIFJK/WDS8EF746poII0IX4
fXUvRJGQLscNsC6u0WqCbf/oWQo7j9uETWcTJnq+zL1rvmLr2b+la2m1DggEr8ir
eA4bak97xdl/mE1ARJSRLGJeDYbnBoRezMOs62ty+ZDglColXcwtxLpmxsH/Rkjl
r0rdDsC+bsJkirKTtuzDWQTBiMDpfxuXP6TT5Aj1/ETIetofaf0GYwAEC2ZedVN/
9h8O6DSmSzf+A5X0xHtCsELXMRcJKLb0cFc7aodzWNze/y4C2Obp66zh6PrXgknp
860ihDnSyDejNCCZpSoh1dx4Nb/otk15/vaYSOYpaVs/fkyeOjzKthVjXzSk4Rmp
Ncq+U1ce/pELq815Q4rgZ9qPJFiDoJUTuTDEHo4ptTfXww0Ber9I5G5WFp/QSfIM
s3A2LCsk3HQ0FvxK9TofDi0gjiY6GY4RiEVNAtijmhmeMkibeTzE4FeaJn5SlhMQ
M7JldSHdKNDDmmCm94JFzcra4q5kB3dyUFRUGPfQUwHIjoA35/UzktcL7+HSbcTq
OR2uNmxMh6Cab4cb/lsagjJ9jiDgQ1Q8dMrzdmP7cz8tYhJknBQvQcAC0lbxDhk+
nNxzCAnK9roO98LIQZgllZmap+9vlvgrLXcL324BJXmYiEwErSJh1izVIIwmvwOB
EIgB4qbiBY016cA5CaztjP79snS4KaODpea7NW0c1z4imrAJBzWoOEdiTNjihXaq
6ztIZoG16tVjpBZtdHivrBSUSGbzXJi6aYbfAp/eZYVl419H5ZNK1TAXk82eepDu
tt+vuXft8N+F68RrFRwnR/aFwqmaz9O5sb7xeq4jmbD3mSSgYmg9Qg7VymxQeLS6
Kb7kaosWQt6Mt5XW8XzfAYZRQqR9iqtT4IwBzIiK7TjVAczGdaIM60bD1NlXSLND
ZWAfbdE+kUdSc41Rf1ffv5wXf4e0oy1g5vsjG7cuSbv6+prfjyeTZWHCXo1e4qVz
ac2yX5T3AFOK9/a3hXRsfwhKmSbNcsswv60kW4XtwZpw2lw3ftM3rxmz/ajoEPwl
yaX++UF1TvKUny5KRAXQVsP677+jrrkZB50vf/8r+K6Zs715BYDFpl9JXUz4Bk83
yC9KWT1kNmkuYGX2nY2aMTcD1te15BhtiBmqO+GCftjmnrLVVObWbrQh1Q024u+Z
h4y1dx3eX0u2SYKLKNHvspItbDAL8lbDzaoOWvYvelGFrFZyQIkzOh3nbQ6ITM16
Wqt4s69ztLjjpGMAjHFJnCn4v0oellZtWPH1y0oxUpEkg9P6a/tE1tq/ofibet0g
4rfrFZWKrcV5FaExkKW0H/AiV2qIAJxbUN65llOh9k/6fyMy01cZMbxdlCUSKoXE
GULo3ZWymq5gHuLoDun6CBBnm5ohhUuK1iFeiACTv0sW39pGZDIyettah1mpKKuG
/s3Ja4LIga/eioBWEtRB9MPmqs90eDmUoB69yoUS4JFjoa7n8+34z/IDWEfC7ZGf
xWtrzGNQa9ax7Q3cj/kOlg5yh60XxdGDvQrjluUcf/aUGtviOIySspYCaM9Kd5ut
9aSOF9oiV6qUHK0Y6wH4Eg/sKptFQlyXCCDRR18caPtpx4xQHSSbOOqpxagBDpcS
sD9llVPqTyGNhfbUzHglq1LMfRorHGyBB3E5OIWzajYuKnPepgeR8QCwCb1nb9Ol
Kuq/tmb8Wndi2PsKrmwSQTVNDANTSbpzbh+CL6V0D/3gR05HCdgS4EqRv+Yh75eJ
R2Ltsu7Fb4gJxBRe2Lx0CSVEclLK6JtXmjs214pOsFOACqBhRY0j6IRnK1q5tMKi
EeH320CxUl3o7i/+7G8ln/qr8cnLxVjPKL0kMv97YsKOUBUQsqZXBM0dtm89cplc
y4lcT8sX6+P+EoAnqG65HFMTVHH+RQIFmBTnZjjq4aUN4el0aUELI/js5GYseKVW
0+vpbdZ++wEVG2sZPpbJhJhF+F63s2Iv4ZlFHavfjjHe895ZZKLPs7fjAdCaXYA8
GAgb4ErTxc8+AAK+fnN+5VfntGBSA9nSZhEY18HsiX5qGMhKQaGPf3BAJ7RR9lGA
cxT3yePfsKwCbA0+OOkGKvcZaGfZVX95Pw+9hmapPado8MI82P7Wm8uTY8Dz1QKN
yf7OUjMwxgtHp+LXLmDxz3kbgQV+6xmbj5Hd+NAA3YQzDxwqdWjMye1oM6hhKYHO
VxTppPcGPvD7yx7Hq5jPSyGKKojDwA1JcMpDEM3SS2ffcXUW4sr3J1CsHNsxtZXV
uzXn0xx6MwR/ahsR+fhS1kFcJDyGgoiZIB0tGDeCa27mTwE83cwhqCd1/54lnSEl
DdJPzNdt04vx6uVLEgTFy7Bj2wFxj+AGenND1JYRH8UCGQd88uL9OpGe2UaMm0xa
du6xeUbNHILMuTsds1j3GQD4utmhuUHXpgTFhxeMdM9DRj9IFrBY2turxhTIhD8S
pAcVDR7S5w3+upJDs03GCZH63oXpJzbmgnpYNTdXNtqXC2ut758D0rBou5KLHf2b
wO+ITWEg3+xt2Po8Frk1aykofA9JykvGwzKgO4P2/Z0hiIUr5dNaT92UFT8HHoUq
0wqv7Cfvm0TO2ABSioiPhv3MEc/tF3AsPB2p2QjEwSqIcZAzbfCMgoL6SuybPo+H
9lPH6ZIjCzitLaScyflYdRCzSyERwWj2F2eIVGmReCrnDcXwqcrGVGeq/l4ZuTDf
zvAwO8Y7o1MThCqDrDezjfY3aksjkxse97PqltFLgj4ETnmT28SNnapA2fXbPi0j
SffWlTfHqXfmVef9xUO9S6nw5ev2giR5feZHCJdf4XVRLHowS87iVnTKixiSRKB/
mPnWiWxDqPkICwEm9IJ6jdwDY3ok5Z30Tv/Ed6MK9iHzlaYjxXdY70Qgs98kXZDb
+vrr75BboRfElLacgBnzr5U/sUP8tWDpOK1KLymlCu1s6KdYmk3gq+79uGIJBpDt
at6mZ+yJTv14YgBbSqfWHEZiEx8DOcalR+SGH+ja79wxQOjH/G6Yv9hutx/tNWs8
vqQILVV30RIEuCMn27DWLEsoLmPgpBP9yAIXtUA03ickSOBzUNAWYDzSNnw1fJNY
mMLMBzxqysukEf7aBBsLJ3kEEM63nCRTplBuIRH+45Tvz77zTFfVJgRnweGaHdJo
osZJ0HNRBeDc+nTD6jaw+ds9GC7k/o3tEANQgzGeKyRZGN5KnCYB6/JSaradswvN
3AJLGvNe/qMU/N3/PPgqrcSHIBEnnq/DeVXclxepdER9vfhKqXvpshJDMYrJUjHC
yCkxvGn/MUGsqWNHAD9jMJ60Aw+w3F25Xstg3XdtzeE/duq6+nDwh2fI29ovBcc8
qC8XOtWFT+nywuikBxgg/5kfNJtCd29Rfvm27/KyvOeAV7bPRXtAZ6cdHoGY2vbB
16Bo48vb2rwOWAAhjv8JU5BTWoEFOY94Pw3YB5+/ZoL6pMO/5Qk4OXfflES2UHnJ
bzVs6h6xnRMmUcO4hb0rcp3x5KiuuF7Wy5AuqBHac5+Tgubvl3uYTOONVq6078H5
VCf8sj4Vv5k+rVklWA8F50XLvFFXSdh2SCwsyBUPStv7we/Fh16qDtkw2uxDW6M6
XIAnGyOOXfvZg6HT6JMElYbrtIk1B7Ot946PeONakmUK+CZvuGApBpay1qYJxAGq
slaYoLykBqM8yVtsxq+yvpG8c4guAv8Y2ALLBGe+YnWvTE7rCVlJkxayCSbpmGBp
WteasT9mxPnp2MMFswrgCs7MzOYaqf7K/zT6eb+sgg4/eNlawK/5M1/IrppItYa3
Q12PknR2TZdt0U5vWJcjn4/6iJPhTatG5O3twGwLZTCfZCeH8ydV/u/gEV800Sg7
4y1WC9v8Rd2k87g0iiU24N/mQYYdHB20ac11g47Dq2YrRxuk7UhLNKd+GfWFuLUx
3mJIvYf3+yZuPD8CCIa5Mz+7EHJ/HG/Hn9YLOlfG+lJ0vNe6XK6QYlI+LCWYMKft
+15miGRb6clxcrygUwstmt/wF4/Tyfg6bJc3xyGQAzEThp3cSaVYD7QfsGIXR3qm
pGQ5drOro31S579lv6sLtXV+zpHJQAc6T5sDyUET5O2mNHG7QX1yAVRtaCBTrKHK
dOyDiRx1SVt0klSPBBjt56ujgCNFCxoePobmbsv5F44r1K67ABx5r9rLNZnF2BK7
S0xK9s6Qg0yUGyAQR49kGx/Y9QnD8skZZvWYlQrmprqghyEr+h+g6HUq6RrOwDk3
6gSCeqDrcbnXXQnFajbk5q1eij/YuedEpOm0+WtaGaxTdalhyIYcHOlZ2uQOeBuC
H5MrssQzXkUMaRY0XQBMLU978/ZNapfo7KYdL7ymq4CiW7AiCBl+pWCr4yooRrr3
8vuxwhCoWpBAF14GOasWBZbBYXzBY8feEbKgoQ++O1GwHJbuR12iBAzNslTItXnT
Bm5jg33wi//xiP7jXsnUPuU+i8C9IygqzzlwxJb52A3RsNoHWY4+GvaKjQQ0ry2a
POfHednz5uJd8/+KAwK/qUwNQnKO6FB9jADM43SNt/ysgMYAI8M6Y5zLkYKga0nT
bEerSJ2Ba6VzK+MKyp/rEzw0H1Q49iJNeZvg3v6W2s1BMGCXjrnq3HYRXRygIQEm
MRqfo5k8He7/OjZC9sRi0kMEX7U2qVmZoUxAFB2HethegtnowPEqThwhAMezvNNS
2Kr8SKvbnDZL3JON7oA2GynQwSRlo2nyvcco2+Ve9Lqkg7s1aV0HMgTm36MOK2LQ
bJpcHGKPJXcguetfg+WDrhblV7ZIG/sH9Hol9qMrt/W0FKnF5NJEwAs/FcpS5IMu
dH2SAxYMgLAqwPaWn6ixGSAUC151tPCFSRnYeHNMyB3Pg1ytfn+ExytlhvBf/WfR
Gyhuamu6Bbx6BvSbv1L+XbceYmrUXKR0s/ZngL3bY9D0P0KMQ9oiTbsnpHfXiKfv
0Kh1P1ZWRN1aqHwu2Qfe6V3JBHjivjdi1oe+aSDDydf1Zpj7PjCyLDfJFSZObl52
gUSGONGA24ETrYSoxWO9/QUXCEOM91vgaa1TP6ETuxFgm8QnatEBtf3umWzw4c9H
mVPJn+HEY8YkDjR6itM1l3hyoaYO8s9DOp+jLXOwPUNQBfZLg3EzfrQeHh97xy5r
hFnJkDCw6ja3c1Nd5MyoFNvJZXdKfGB5R4rclwkBrc6XeWwkmlf1NmIy6wVKruUK
eMpFBWwixtu9ULNqKB8MGOMNp5s+ZXod4gnCeLl8yD/cdglSYUI8L4Ou7idhkv6P
patHQjSnIGL5NyyO3LNFnip6DV65t0o7vioA26R/YNG1weO0jrAhr4hnFz7Ot7pF
TEnavIyrrFJQASRVN1d2GBhLxB3FHUWGRRmH6uwX9bojb/iz/odXinDU0W5MnEfi
WYVA2Jt1qeetlUYcmMBlal+/Za1hA9eWtUwwcRNInMU7u3bQeSlJp6rqUKPoJXsO
ERhIJ4iQpCt+1ox73IXdCx3TCgeFsf0tcb4bqdQAz702tK4uQCpYeUn+JYC6ARad
wfFV6dJcZR+/u14/QXiGh+yfiTIpJkR+LP4twh8RHBd+pE7/MijV8QG7bTzOuboJ
R8rlgSmvJYdNMFjLQZQN4U3Uw1WIkC1atbcJBIfz9BMQxhkcHsWgy5WG4LfS9jBo
Ks10JJ5yqje/xbosvry+EZ8whaIKjgeNN5ihVKsj2XUi6OhjXXCmhK42cuT5DYRa
tit6TiToR3a1wAll2v54Z8xbtCBlM7UGxaCDJgrCXaAg5QBGaKq0Z13mfimI9RJZ
y4o1WoplvOqnk0txjW/RkkP7p4OBsvPPVrPi58j1xldtOJCgYmqena51hccK2MRx
Bi9dWbcxMq0HAE555VtfPBo9CIgFTvU8h+YwUCWbsr1FN6yf9ZNVFH6fAlt5EVoj
85Y8GVd0PSHBjsaaxhGYOVw70busUqa6qZbytDn69s7lSoFjlUMFH4mPKB8wmXo0
ku4UKNpE7WH5ODDjeGUYwLTWKVRY1vCLSoWWyiHgWGYkhl4m23QZ73AWRe7hc4pG
TWXic/nCZsH07dzZGtXhunLkWNPSW5hLKi3zNuscWAJp1TOZSyMtajjF79PFiQ6Z
EDyP5vAsY/DOltXAKIbsyTHsnq9LGVGbug3Da7WBycwIY6Y9MTChMAyejeEq2my+
7rbSg9y7cgSsa6t+fEcI0+qAyvK5d/WsBBE1tg0xj2leyYY/1dSrp7jWosS2yyMf
Wgv5w+zY9kxYWmoeWBhEQEXZ+uYQeV5ynwH28Oh5OrLGWwYvZPW5NMS+SCX/JNWj
Jg4IyH+3q/lL+HZnv9WTMLUx40vyf96i4T4404IEPG1M3n/wQ+zxrxX1Ozz+0GIQ
OLt3RdEtgZwrIGrmxCq8S1ecdsm0S+ScremwFpbUeiYi/7COZLihACAoXOsYqLLw
OF110lzMFHHEVOrRs0rdNeOhJF9Umf3031ny7WTuKq7DwXo33+XJg/JbMg/dqoMH
HsZwig5+Jse3roTx0FpHqYFzFxFMYrl+QOcOYX/JJiSSwqPZ3thyIkCHqrkcTvZy
HQ3BoNSxjEO83A2V54i2ZdCzaRBrsJjMhFgbGCbmC5BjaRr9zz0+x0Nrvq49aMJE
9xdRpSq4nu3CTOQ4Q4Pk8U1fNmlA9WEZLSA8AGrxrMFH4dEYc7rIsq5yyWROfcoi
p5+qXyvoJJEKlEBNucrufB+nifFTXj4gUKuCihoK6vxEAkNIrd12uyvbOyOT8UWA
U48N4j+CMp5jytVpNYOYmnpINVifM8vp1VxUVy5vXad9hw9/Z0R+kO8g3pV62REn
DU3ECVhJX3htZcsoIXKLQ9CbTfGFY4RIkU48Itpxj/OflvgBzVp3TTjIepUgBiyi
xQAbC/5+DYGR42v+XprTBH4SojPgzNzYasUl1aIUbKcoxWuK7zRAoufeskHHTCnA
4brSIyt+/e+kmnTc49yaoS8eWFwgBiH0rA+y82btVurX2iT2OLyIFtbPWd9d3C+Q
A++pLth7yzZRvNWHDgq4dDlLURRig76oHcOzbM6mHzCZGyjZtzQWnAkqLRoT8Q5I
NWRFx4Nf4cl7CqnKAsNOBtPhfA8xOr7uX04vgltiYsIKB5p4r19r4Q8z2fXuqhqU
IsgCBkk6zH6ZPcpUE4+fImhg6TWlyLVs+5NKepAf4ynDxQUokLIu5qVAO7SycreM
lsRW7kbbgcbkgj35HvQqfmbxWpAEP6exV5wKWYAVA88tl3rXJMr6/8XAAg8APHYx
i8oxUIXe6QyFw0+4fcv67BnUVciHX5Z2dxqR5IgS+JTD/mfgRp/x0mTWOUZ0euj/
OIRNZtk6Lg2pjXMSM9xFD1xlXIxDqdWNpbER+qbmlwywUJJVt/S+A2xVXb+x7juT
yTaJOicqRZlzBrEgFttfYTZuEUyjiKB6rwKiRmXrAvzAtQkGWk+U2HKr5qKSYBag
H6UJWzcAE1QMhhCtYmM4cpZatpmr3dqP2ypUCOlawzRVFEYxOcbImL3BtvWONywR
ivccK564Fd4XlEaLtED7stgEWeGQoF7CleN+hz393hmNZLLU8KSI2mXCbCRBOE4P
rPHWswJkKkVlDQ4cXUVMpSaLNj6IISrWgkAiUrno27KrxvmqEHLxBHsT5DZWA9G3
Hpkn0aExY0v+glcA5/uJE+gaFmbrUne5mMnJVawiYQ3RVmC0ui4Lz/BFbv/qTKCn
sdJWUvJpeKrWhciqCPUxJDAPzwe+fk63PNwKmZl2w4MKGZRyMJlT1Szgzz6kY8Jt
3KFCruJ1yY1NjWazZugaLNFIGjKjDcInGQ6iXBDREjyM/gL6eu0v/E7Nlf46eh58
1hq0gOo2d7tIqtJwiDlUX7gnBD4NwkZq3KHEfGUKvwP478jDk3F0CKWYBTPrISmY
DLz+8VLMs19u4kpkO1dwBcSzMkaab7R7IWKy4heHP9Ys+V9BuOdsaWrV9u3g2MZZ
2HzNGREoe+72tTJKxTCXd4FG1QmgkdBEe3qPrFuHDPnKmkyPOKqgjm1gpOkmSb7j
ewIPs1JO0X2M7br235WIHeel1x6h0n3qgaerSijJKoLr4aJgOkWRQco3VPw+1FFn
SvTvJqf/tt573Km+70x+hUsrbI8PJa/yRq3dlL7lbc9xFaC/vt3W2+AnICBYmJsi
+WN/geLwHx+DDcxSY6V5hY2Dsay4emzn51OvfK4podtADwLKvNAjtGsufDz6rZyk
B64x1i2q53iZSGwBDqZIY9SrgEAcfNDMsci5CqYgWBRvIftKMGvlBPMoyzBi4bX6
1bHlK8AKmsedjJwOy6cQfgScwbi98BAbhCTbyFS6Jrl76y/QQZFzMFTjqnKJ/JIh
enVX9mxItUX29jj7NVePpDXxP5YieAkeahBCDvdrCzrV5JLZIeWH3wlsfNbaLd4S
lzpf8gcyJJy8KxsWMv3CbmrvAvZiCtQ2L3hCzsaz6k7QAdH1xqVbxl4uQb2TC7VD
+iZb4y28hUiZPiaZ8p85ne7iBsTakKuDNmVo8VnrCpchygcjEr2MCKMGC5nB0Tlz
9RFyhPTVB9hW/gPH87Q/qfDbUFgD7T4cJ7csqIKntXu5Yo6L1EuXBQmoSaVr33V4
2sDj81sS1CGLvcwwuKbvT4hnworSxcyiUPR4PDU0m2X5cjHhRhtzlpAZxoQtDyaP
KtGqpqHm3C2MlKrFey/SQvXWQw03VtlHfXK9MEmFjqkX4H2FQAQDKEwInUK9F4dQ
8Yae1EjnqCcOG/Z85fADRFcdRWraoD8LPY1FZl8SwBHnus5bQu6X4+kR74aJ7G5U
1WVHkyGdHHlTjGjaz8N1RYhohNMHgMz4QAqW5yxoY3tFunUj4G7AapWiPrXQJ07V
LdpItzwC1fs1ztK4nRiLkbHlfq+bPhSIzqC+JA63C2DDh6eyV6yUsbuwZvvvoqNP
JZRQ67iMz3EWM5rLQ6rek5LlfFeXJ/8p2PPJh91Oh2ujE2cGK6sSd9Yp4JboQWbz
vniV04+8XNzCTo62f79H+FUtk5iSQwVr5P7rQnAH/tYcT5LCU6W1wJwIKoX4KQrT
jt373EFDVa92l79OltiG2ccLDTDhJi98/yowprDkXkc5mNLIvkxSaCq9baKrgnIO
rU2Ri06ZsNqS8Zf9tLYwM1G7hBArxdkIhwgbxcTMYHWhEw9DlEVbZK3RDe8/CbBg
HUUsBaIWoAyR++r1CMFxyJWBDBkhj5V2y3dKufMrFQAZX4jBIZpvvMRpJSWIk6XU
DO1QUT2yvxlqZMjcVYdvrbJcQd7Cm0WC2s1eyCHscv6Sw+aER1LlcMtKyd3NrYup
GvXfMAIp+Y26MvOS1g7RrVYHjeTNxNUAPuVGxJi7B/Pj3I63peb8pkEvI7JTs8ZM
Mei+9ww4Ufk+eFZzlDR005V0hGYwFCTPNI0zqrmx2apsPzgx+QAymFtT9lGfhGYY
OG9aGgdPkeRR+xWTzDHCIao0fkZr+MPr+MiYLZh/Y39/8lU3wNLo3V+Ip0oMMeHY
PBEA+gY2+hP9pG6EpTyuMEwlWFk3Khn9w1wpkz0bJ2A447+llP2Bhjr2Y6a81ZvV
+saqNd/7+3jIuXY9orYTqWWhSXrGTssHGnZYivgrURTg8xM0iqFLCLt4d6wBcMDo
I5BJqNsJRSH15tB8JNeopDAN6Vjcdk+VJ8BcuxXsjJ9AkQc5eXaLIU3fXP23EkzY
4h2J4TTx3dX4MYNNeF2ar/l4ktjt7w5k2Oxm3XKWNDKL6y+jZY2Gy/P53vB4TDqi
csPZ8NNu30YcP6WznkH2h65Ah3Fu+L/2IEfJyCCLWSfm61Bt0ESUNHXEmRYLjTWO
d9U87cBUpvWa/aUDaWii1yv2PdMCorVWMImHXP2xfFD8rD0/qy2nUX1gbDy3O4JU
cT4P1crJyKFzZ4JmpKZccK+g1Fi2SnjmaEjASn8aWzVglGfJozmNCdGsIHBtxFUA
CgDAUCmFtSIwUtXmEt1B/tDfiO8PuV4tmWXgQV6xT52Rx7SXqVhRO0lk4UiCDaEa
E6GHjfZ6sgBbB3gmy/E/Be67MGHYNxudf9czBZm1eqGiZXUoxIiXCuKRT6TpVhtO
IbsRNaMQ3sEGVhWX69CpU/jTj7wgU4vvLHDFGVck0OHmA0eeqovfySn6h78/tfdx
sFS66f9QBm0OgHAUZdWzvF63lmIekbCS8pdk8wixYnIp+hhTzWo/N8rk9gtNLRpj
whkp+UVZmrhAVuc007t42eQax1eE6jpsHCbIvOoZdEJ1I+Y+LVusennT+rPINLTo
T5kLq4yKijFvB9q4Nle/Mubbpocz63a6nV+K3T/qmeGB3tyJ5oS1z1tuPdkLPbbb
5xGXZSkxYIHKukLXZgtWxgnXN+X3xRsn8Bbuw4sCqlwWvliA7l88xWQd4qspAK8R
8xv33Ew+0thh/3mbQ6iotFJVEzVCESFY8CeB7kx4+dLRWFydCp4XKGXjjS4F/tGs
AhbMeSNufSPWCxD6IZ0uvbicC4nQXpfE+itVtLXz3VYXuiW2dbwxSiihXJYQoQS9
A7It3CzSfltzvWxfnraUPyPaGuBDzTRv8KUwso7ysaNwqkBndKOS17pbiuiy6RwB
j1sV2rSO3iyG0v41svJGvi3GGyfp8Dc/PgBrEMC2mM3BXSv2cOm/fo8ZcmNggu3/
BC6iOkycoo+9lchpTae8rOFo3XvcZdo47d1TsBaSPyECBauyYM5eWNqX9vHOv+2D
tEDgdtEZUFxU+fDZ2iXyx/VGb08EO4fUBFkGeITxuClNBXI1Slq2ZRCYenrVIBqa
dXK17Bvo19Hs+EaCFAwjcGzmJ/5oKw4ppZbTnGXD3is/J63UP/72iq5aP2i97f5O
ZOxB/zwx3+GQTZWCRWzrBodBi7KazOMqWlXx+GE+u8WortaAMjoDNtdPEVWSOWyd
wVlOwpY0SpH78MctAuHSiabSh4MPPpggghElAsLd+p5xpq2P7jouLJN7+49cCge8
Vg8rzcfQ7kk/1+xCWXFLH89p52EjO4Bmuvbfmo6SZ1ZHQ5WY+jm2gImvfn9zbvD1
aTUKKx62UTBGjTzGVq2mbHicYW8iX1B3Zt4Al6GUsfxud8f+CsfSXMRObjH8pnNh
cn7yoaUcsNdlTbLRFVb6q83emt8m1RMd8abogWhgUtvs9/V66gaoSK7WpiT5e1be
f0XOevqMFrDII566JgkcBBynHoRKO7hqm/0mOH9XnsbA/9u1rbVFiTcPxc6lYKff
S7tpNQQwN1RvxZjoxzOYlt4pxBUMYKlDMc0m1sDkLgUodq0BGbawUQIWOz+HL8sH
lZ/AU06iZpRmohkZrmiv4SdwN4Mbr9DMCNmZ3DGfP9guT4PLnE1wQMIiTrlC9UWJ
0PMxVBQAEC6OA0PfcTz1sQ75oF9dpAyVbSEQsEcgeGK8gz/Ot/hw7CSRybbrthwo
4D616kjvACElWIKYiHNtMDLBD+HGS3f6kSwUzLmEcixJGPcfX3YlOPWesJAQe8HM
WKFpw06tUDgulkJ4qfwJGHV/a2QKURzhZNsjg9VspzvVpM6qeoQhK4pGeQvI2inl
ONE4vw6AJ3GOds1QrFYvaX8AakBeCohNBsUGuO8tpZlbTZd/whIeALNORPwtIGfJ
NsNR3h1eyCCuSDY8+z5feB7dtjFYmDnr1GNWDONOTc+lD9R/jrIBgMhSXbaVObpy
pZdVOvWSyaKlr0x07haTAHoVNNJGtBK/+Pxb+CPTpFvIkCLr22l3sqQJLNcF9tV0
mkGyYPicf1Uy/rnYeFF/XtL/9iiQNG066QfaQ1gPLGjMbLsNnMsUfAu4dYgTWtyy
1vTV/12hSk2VJmZpVYch8AxSc8Hh0mz7bja4JzjK1yrqninMtIuIWEy04dYdsfxB
1ZeJ/JoupgB6GbuxExdgt0SOjBRhRrFNkxYq4l5+AxGv6e8EtIEs21850eVT9tQx
DeY/dqvrnnXbUsUs7rsFkbsr23IKTw8MBS7dqENlhgjIoImUOqoiB8G4db3MPNex
Wqlc6K9EWvVvxNbN5qJxH6pVZ/osaP/7ic+ljU+dZmq3jvvhmFSG+wJRKlnXPaYC
kdGinDRqtPciVhL79sidGXcCFnELk/rtIujdjZqhU0sPckbrmiIHENhU9msoB9p8
1uJy3atSAGZhmyO+zw0Fl+ctwMCe5/lSW1famA/DleISLLg20yXPHeQUT12hd9M+
Gc/x+rROl/qq/GKFs90R1pagsKGgWlxQM1AK5l4SHuUfLwBGrFcjOOcKfv+EFuJh
mBtushaUOiyr+q4qE+7zPgB0FwaOalqpvTcJv0FPOcAGnNW1HAPjS+8xaCxvoR68
cNeIs+ukEW6wxaZGSc/nChKjwJ1kcqPoWbbqaITdngl4uIP2Lsl+4SUPSJ/l/3Jn
QY7DYKvF05AtoNU+BpmqkMtiTGt2OhlWP47xTVC7A6Nq7h0G4cD4hzNUKZJ97uJ/
LHfRjsMn/Md9k8Pgm60YP29EO3FlFNbfWBxEc1q+16Yu20ijGV4gdNxDP7UAWqlS
8ybviY5UTgUGH560o7q/GkwHGwo1Yinn2upKIqYTDIMvQhPvZSagyiDia3dnipY7
UHuCvJX0tc5kXDYC2F/4ofzOwS5TgsTZHpbkjgqkBKijJrlcipljhK+i9dlHcWG1
1m+pEb1csYmiHME19kQOr2qaIUCEtOqBd/HxUC1m8Pn4Id58eiYN4Y8xEgJrpikp
fRx7tN0Lca2WkZUqDmwHeZxdilQchFK0R/6bCEr6zTS/vKRy+URGzA92SLXQcB6d
1q7as+dIpGSfXd8BtmX6Vn8iT0tS/Y3aZcGzqTX3Hxa8x0PjfEJEwslem6ScxTgY
2Zjtud3LL5XPfei4ODMynknIOuhaIQ3bkyiRT403pxrQxwizT2FcnqDerpPUUvSr
uxLmjA2mHMPAsIv44S5UnEHWaKLlZP/kK7DUu4d1UUgym48fiKJFTWujXZCEQfKP
ilgW35O/jDk9GHJ/kaw1cGqdu7Y8mFtiaDAk+MTglJBvdR63zCwzFVZclO5lDIYh
JZhELYnEgoeBoGFKjfKwuqiYLIvqbHaZIPYkUBOjLoyH92zRVgeHZNf4SIrsF5K7
4msCh2evDLXpGzuIuZLmMenzYD8el0p/fjQVmZFxpdgrRtBzI8wQutqCZx51KoVd
YgiDqExaCxfeWgBVGw2F5cTb2Ngo311l+IEbX4uV5HL2/YyTsP9+0ISwFNZ3xwEY
eqtYfWnoFrKfH2yC4lyfrJJtTWd5f5/eeLkOlUVCVose8SzciYgclLexLAW5I/8T
hT0bR1QHi1Px2Uj/48VmRXRBtlJfjRAKCalln4IU5WOmjm8Z50IZd82OzU8eryhe
gIZ45RXzfI41HaDbDB4EAStmNjwSO0Vt1StpcXU8wWsgrTxy2yJDooA5MeZWN9rk
y+HIhvj7MWNraxenVmiKX7Zqj7vgeXLvw+oOnu6YBDRHiP/DkUTN4yRzSlNmu/VX
ObxEL2h8LyBJZMoJHUi0tCBsVy/iN+PDYoEMKxZfNUdQl8eLznYXk6Jd1+ec+xt7
ey2eVuvM+03eaZ6G+rtLqNMOY+yIcaDwr+SMyQZlRaC+4rEKOJLUednXMrsobeEj
OvXO/oyubbAN9v3C+6W8d6kGWCi/7z2I8rTolPdMttXpJNxNwsyUMNTxrSmODloS
ICI4/IbtFpkkRZcyNW5IkXNI7SOTtBfjH5iC4hXDULpMzxLPbTr4wzacCHJxdscE
nnGE6W4Sm3ZvK1Of6rGVq6CT80QY/X2ygqMR6kvazD23epJsoNOTX+RMniwJV9o3
Bl12w6JUhlO90ZD9oHL4D9hS5rEYp0VxEcFeoRUhIwSyO8+Ca0104ttohh1ihc+M
Pfr3BEunVkPcY4pu8hKx+FOz1YQ/sFrcVOCdZiwK0x5scQU35UbeonTWvOcFCp7v
uDIeEQA/waFfd+HLgPv2FbMwPxVf0q5FaOZCVJtkkvqJTYpXxhIBXpP+5QTWXY1R
ApGzhW5pW6du3hb/ndxW0pDfagyfwXm41IyeS/pyB2rp+wI8ZQe3PadIv12cCLEf
aD8nrkiaW7PM+mgeith4aKlLy3hs5n3lLrGIyqOW2b/pwSzV90PAqea+qdOSkxYd
3pm3C3WljftjPSAnOpkvQHSQHem5ZkaniQnM5elffG6urtYyJ5b+577SIxZcokH/
D7kLzX0yhR9RyF85eb9G4RrerU438pO7Y2pXsMGC8qg0uEDGTeDvKYqGdW1brIbZ
Zm88LIAcGmpKY7MdHH+8E+AjsOk0bjiNA2deJzE+Sc+sOFPSD3rLqTxQvV7z9HA+
oHv7Vx+5WVhGr5asDyWx1u3y9bZpeuDKmbZFMJljYPq4sEuH4dSHUaaT5aLL4W7v
VjmDkLylBROTtzjLJzNGPAwM+I+hixPoLYDuacn8c9hsjng0xOkBQzpuDt9dQqL9
i5JEcreoX9eG2UaP4OQfeY98HQXWyGaE8utdG74tlNuQQYYOcaqGrUxm941wroJN
6yIbrsvV1jsGBCjUAStX4HXtp3vH3M6Rpm281S1NFxKjcLruX2kGzuI1pe3jVyeb
MS4TcHwglhI07Hrcz6HTj6MDgO76nCbuZmEAU+mVL6QeQWF8qAl6NsaHcxOQ5e/J
e/PmQrug9fXLkHGew29Py/57D6V26Bog5oWT5G2FcgqLscyaeMA2sKRhzeepEXxW
Qj3ORvEBziWKNeB66Mxg1q8HHlMGpJIn05FOKElzGTufgRDy1RvVJR15W7LQKrVQ
fhtO4a74zCX8m4hjC/26ewP/AWOq3F9FI1rhnpsDbXats59avNe2XNE4bxbaZDVV
k8OeG9h76rDN5PxejjWsDAh6hCzGmTtMZHwz6Yv3OTS+66mtOM5kYvZED9cDXgv+
jbTqu5rDk6N1vzAa3tR+A8ZDKe1yKU/qR0gmxGZF+dYAXG+FjiOgCgJoZ5ij3SOV
XnMhltYPn2+T4rHBcSTV0qjg0kPsuY+N7I1O5H3yU2wpIQp/vj3L/6eMes3eTHQp
rJ9NlaDlfPuooW9qzIRKTEbUQV32qvvxHvPxn3SJ9Z5chcKTPkiPi/uEuQPRM4Ma
guHrd1LkTWW9na0KavhVD1qmya5tmwcQ87/4Ufcl8lQM65mJNjvdjLhyqu5k+WfH
Xt8b7UOl3qmirHpH1fTmVBcaXxLRsJ8Jr3Z1PmxaRh3/USH5p2U42ATHo7W/poL8
OkSDilA4FWBrwaNEBtZwf70Eg4EqQq1/2LRgmAqeBV2CCtAJPxzcif1pBTb+wknD
1j8pN6ObB8Y6XH3OICU9UjgHsz2xZyn9G1qSv4ka26ThlQxKv92WwIGFi0V73c8q
aW43J5MkrShi2vQegsctGB/JDqLFBaVQio7HP8Kj6cqXBSd7MbKu33H4+dyqgyQh
6Tewv5uuhdUVFmj0jnwHrl3xsfB1pGrXjihMAOv7slKxRJRieXIgcHXUQPR8AQQV
c4NoOcISOXsHtiMMextrqqVZ5pFK6/wo7kxiJIOjzfn/ZTriNb0aAK093TtnH6hm
xd6TAQg7k6aJRP0Tig2g/VpqPQDbYAC/LK+QOgee4W8afxupYf5YIA8S9sePcj1V
6IdZ+p58YHDh2vY9P1be3lTgm5JkH2tK25ifX7whnSJ/qOYEOkM1T0td86sQXG/I
qsLZWapzHAeHlx2bP5x+NCh0Fs0AfQjPCIJxiQEl3gvSN8gdb6yj+0/cs8flojUC
1qHUrgjGquGv5ZOVAItRy/jrmUn2DTJoyxZMln4lBk3VJeoHuPmptpkVgiatufFX
OhpozsLNOuemTa0YttvhceiJXD6YT2bURMufejOIYQrnInT6P9Ed38Pyxzos80jU
EdbFvhGE2xuDU8/kGERjk4T4+0mQAjzAUGItpRDASvlf5Kx8S3H//dd2wKA7zz/h
wN4bqWlFOlbmYdbfQ0Rhvg5f/q5r1NrSZH1qI/7p+S8TsY86QiTtHq2xZ0c1lyga
7fXWhfwP5L9mAR+Iux6afuDuttaQTP2WLYWcM6g95JJPjcgDH0a+WJTUyghK41P+
gAWOdwPCz5a2bHsmy3GXnfPkZIT0l8UgzhxZLzsX52xUsUqRjzAJUrcEvr7S+JNj
WNTL1HSOdOwGTrKgAJrsSDDYATc2VqlM4Ol5UtV3Q9HFH6e68a4ETMfWD5NwUev5
lFVnajFh04yX9tCO6egatUbss49rwSUk5KHZB+PK0HltyY68SuCm6w7LcV+ibSRT
B83BoGdAqesAmP0p9lXZb/Rd+iuxnD0kQW5liyd6sXQ8PmWFJBHR0+kcVGMCz5sJ
L5PZcPcQXvXMo8hNdxto+afJp8LVmAAxA5XQzvUNt+POCFjE4WBEdJV9ZMkPFf2Y
rDoSlteq9RVttU53Py3M79lRz4DiCVYds4iQw6M932r+jslhhwD3NqAhxPRX0pv4
JLi6iX3qUrYuQTU7ckCtkdwqjyoyioVqEQ7PQ1XYeChAujPM/J7xkGNUogvZfeYX
qIDt6fT/b1XgJImqIoOZqpL/mvnLb4Akbns4NmEyws9FBTgqqXveBqMKBdYBXe/R
ADlScXzzP5xp/28yZUH+JaBisP+hJWA2HFvc7NgfNKZcktyNiHEkwZpL5SmcBNl9
wY30z3/nCtjGpALYjTHp8QN2tYCmy2msZaaLamEfv/NzJMms3oJrPqu5t+8PVzXN
gf8kkwZ9WQyTH1gtbFeeNXLsfhyUpo4Im8eKse/gIW+ITqTyLwrJ1oavAstvMH2K
epvcp30Ohh98EQQfYb8QMLdq0tvgL9YluuiE9eZ0xriwKujtT35SHHwAvq6W7QEq
ylMhr5rdvysvZdpQ7NOI9CCC2lPhpitfEenFaTgDs0PxJ9q5BVwHzlxofe1ecsLk
ECiibRtKaVhO/l0Wv6yHAw88N5cTFZfnSnKnzUwtpEREiusZYWhfDM1B8AtHc6wN
HwAuyhVgYW+fhpUsH1HnHnnvcMQnSUvQTqGh3kt0abwj7TLL+1XHYvzJNz1oPeoN
peu970YCQyiSosjrvA1GpM90FCPq9F+X6wlutDLwyDof0LvXtT8ZkhU2gQmcxdYr
MYZ2kWoUFwOY/HeuIdqmccEg8UhPTNDOKJU6HSFWpVjXZH/8DrKjdcCFKoG858PX
AHuuj19mHLHr1uQznEHCl0e/NoV9cp8/yRUnGubYzKV3X2jiA6zLeTkG0kUDnBae
7clLboNcXfFyQUejn2/eGMqDSJqzBb+79pYJz8Qe8mhEJ9aP8cOS3K+Bb8HEyd29
nUaCxDYOs/zP9591SXaaBM1xReFXpRwXR25L7drW7DmWBKvmqDmrDmSpZSxGZH89
+6p42ivtf+P4Ga2tBp2cFv8ZaJuv1s4oIYgh3IohuYAjhoU6IJwozr1C2sX/GzPK
HJ3X1BhBe7pSuM/hDjBKEGQVCB47EmwFr4ta5BN+Q2AELZSAhOsmz7xFRZRHzoJt
qMolngkBIVF/rliXjYzwHb7s5UzeVC/BLtLIG4Pjhj8sWhuNfYfAVBp0jU4nje4n
EBw5Oukf009l4txUHplKfDOEaxeD0eZ4mgZMuCcHF/R3V7P/M8DFTAj5zA+P2Qqr
F+13p7BddrgrH9sGenSqErwWJxih/Wi43T4xFZMmNEeJFlirj8qN4239du/nV0og
3t5Zyqa8Lpq/EtucwjdWMTUG8tZ0rA7v+7ATalwOyIcu9SkdRV/zthLGKK7mOG8f
Mtv7EfMP61rnLKb7g0Rvli9NmSMYC/0bIWqQ3To46U0Ix5DjmAGd7TUiqz7GDOCo
BcTHpPFXzcFRnHiz4p+jUIl9CVMMUXJO/oYxCxYDvNbr+Tg82erBas1+Uxf0ZZ7A
t4GyYzWSzVAWg0M30/W72cS2X3eDcz+m+i6zJygapOABcC+DHw52wCJ8uoFQBfph
lSQvcrIMQm++FoDqcPLZpL5/KNgcL4X0z/LFK41SysQTt34z7wdZ3EBP9NRvVV36
zBaNLOCB6kbhMJvNMYhgAQ4m50kKYli5kxTYrfrQQBpFfRM9wAMf4dFkTGo9IW6V
m8SnTFTDbdV9q4Ju5QXGmFDSE3qfwfTkj/wgxMA+U07+tvTYP8ppLNlk/8hhlycc
IIaS2094S3ow509rEahQ1Ny3GeHNKmbxBvQFMwHX59hSnU+7Vu2Cp06ziuaz5GFA
8VMH7KyJuXk8/K50/zTBIUWasgFAEgTKkzO8DygQafROpX6nASTrBdSdstvwm+Cj
BF3KMvSZfOhkiuemlCOYKXcJdfewavTDp3bIKEdyABqoVPnpH3DQo3xNWUtJ7q30
i5/zEJhS8kIn/I2Pqpw2J44n0XZ4WeEmw3UK/r1t7eXYAy8Qwnbfec+LM1D/F7vB
MLyjECtsaxbJJlRG7jSs5EHgSMtj9NQmfawAwjOiiAZOohw39rch7tT2iCDg8Ngn
IKx+8AV75zz425JrqdyLn4fM7eoPrOf9Cbnb33UFved56XWKy58paw2oydCG28b3
7KGDueUDIOPd84SOEOA2zVYNy+SkExm76IFVfPiZF5/7+DDfpAqfme6gNTHKBF8o
+tJ1MB2qZeiV6pc45G8mzrP8qzAJ9E/XRF5eEICrPnKiWUxmQlrurBRPI3KLrohn
917N8f46KuTXS2DIr8nMOSyVdDKM8Kr++nyL75vjS+quIwjIhm5yw31nP/x3yce+
UjglQ0UIwg4prnF95U8cWepkeJmj4cVV3jmehB6GcnX7JDEnCzryFWG2P1zMn821
+Hum7xCPy1isBrZgBIR2egNn9jgqSb7PHXF7Z5u7vqheh8aSyaMDU6tqdTjD3uO1
L+jBg2LndlKfK5uyxOBdRxgFmKwThs+GJmtV3pX1DrjPEK8M8PpKC8X39qIoZT0s
VeytjA6aF8QccOqNjOIHn0U5t7s1QQ/pSZ5TezCM6IE2zJslgBIol4WZpFyjeQPT
VDAqCQjFYBWsPh1KC32SpWZ27vtC8MI9xyLO9QGfbl3B/6GfeVldYduhS6s7Cr9U
hkfcbXELUBPiKe0JQPtqKmUhQ3ymu3V6uC9RC1GvArfBjNJikLjIBQPUpGgxlHyN
0tdFe4rDLBmO/oNw8JMso1qQgiz+cn4lHYgpWl6KA72qp5e04vQo8LB+2kBztB3n
tHxciUMoUXzRdYQ0RcbOAunNnv/fXheoSgnzin4PZEOHKSiOD1s9ERZoK3up8c5a
dDwevlwmqdO6pLGdYGz7vbIboMx6S/IXyVy7nam99e0IRwVKR6ibat4l4Y1qJqGJ
Nj9taZ6wCpYoxEWPIjel9+xsNOr1P8boYouTrZKUJqS+xn8FYBF+r+S8NoVFr5HI
V3fnehyrdeipTh2q/1Pkiscv7kscv0RcdQXOqcdv1f7gfbdstveJBYsyqYskQD05
0Uky4mH3lOFZWcXGcVcud1BVug2lrfCDCL6rWdCZk/0OfqwUQnkHcBJuYt4E+E4l
wmjcAbi5vEuxDkjP2UwgEE2dMCDPh/RCWcZj6JdzJDiGGomCYL7SiRKpv3Ahh8/d
/E/Jc2vV8j9KsKNOc33ths4UE2fvFMRpWOraTQPzCFl3AYmcwSb3yoNtFX0rmHhn
f4+WNqo+5JCpSBYvU7cPJJBdQhiB7+AeWV2vV0j05de8Jdyz7KUWAFb/BCm4+7qg
w/3Ynbtg4m6HL4IHGOgMmG5MoJ15KxZ84xTWz2OX4Dqk5chXiz+iU1gFiep9rjY+
Vd3UtJ//MnP31ueByqlQBXAIHYAdPQi+1ABgGMtUADsh2Wow+V9zZu2eszFZsOxz
bTgZxeYScUS/xv1tyLL22LRLX3/IEFGDOZDBo4d1EsOKmX5yntIm/xl1O7cXrtHi
8s/wz4DRc2yUdjnBmbqeZLnsVLB8mCU4zCTnFzvhU1kcyv0eSsnXuFiHiDxZycDz
Mo6Lg0fIghBRUCrDvJFzisvO1FKgmHaCDUXXkmtIMYf4bL/J3LGv49+4xMvSisLW
hH9MZt8ZMCHB5kPNCoDXp3QhjvCHBBM1v08eZSkD/5t3xxs2jh5EWXM/BbwkbDw9
DjWBL8PkCxvdpSMb/rDTVMtCHRTLD49Pc7+zAIRcW13xnnj9eJ23xqBp1gPCuxmw
C34SKZYC2Jw0uZ/fqRDFbwQQYHcwQBvCgsN10N3qj9gwFRo1h4dtma/2Z4d1dHs5
mCFHPxPYHPfPgq3KkE0HvDXReSv+C1cLq3jqy4MDFc+Uje1B7ZAq10v4QuBdPppU
+9XNDBqKQJdD31e/uZeKi1M7Q6G+oZh2DjAnbkca3zi3wd9seFCX2bCTNsGsuaL6
f51bd88XqU3Yy/ejgjiiI/aUlJORKlYdBbw+AvsaFA7NWEmERN14jYZVd3DlWL42
Ak4D5P1SjBQb1OL3GlmYpop2qdMmS8dbEbNf4ER/w25G9M/BtFaq1366slpd91pY
4P3aizky3XrqlKeGCFGPoHqIqDVNMqKZBEH4cKfuH6fLA5GIGHL8IzEinAjQm0DP
J2IhpjqW/KqDSaw9Y0nwYtHVmW/qvCM2gu7DQMFsbtupTbPTyOLSfZbBHM4AMdPc
SF8ZEenfV/NJYTNjbnTxfQJEvuw81b1NVmlVB/bR8QrEQQp/Qy8EMaodhnHyvntW
Fc3Mh8F66KMdNaTS6JCaH5nEfYaG3ssTLoYfAEiiRncF5My2hNrj4O6wyMZpOUt4
1kPh0h6Ly6pT9G0RjNMJUbQV6wBXyYdOzU6rV0n/TBWRtHbPvPrv3sLrv6rrXTJs
0GfKSMqmpAU47h4IBuVogVNeVT8uvWVXfe5+Zi4857rC2Z1Jom0nZr/69FjyI2Vm
0h55PTNDpB9xo8lpjIALCUuT+izF/I+IWvy9lGZi4XQAGWsdBtfeccMGI/cZJxnz
sVbTZB3MLgb3/2wWSvR03/13Fwum4Zv1jAFaC34J20mB1GQwRTKlZYrQFpe+8z34
wdo8gjGy5ud8DJH8NnU+xCqAAGA+F+ZyI08CKw7N57fiKb8USLwi7na3Cjrs0AQ7
xbrViR//yhiG9uRpSG5ItpNJfJ4WLXuEZMNKtTGh1LM3aUPs3x12PeNqnpNaYBqu
yK7cG9TY3FDVAHfWyDdd8a1mawYDLvvDjxUszqKoueLsqSR3i04ZX+ckWHU6cU1R
VU1PuMUNDLSZ8XnUIrUHO3uleKu0nC+cXOnQEhjQs6sezTgXjWa+xhJhLYL3+tmk
IoZt+hhZx9KqCepCugJybs0GxtXZ/lQMxdb011LhTaWielOi1KytFWL2wMjvrRnb
OCZtHDRwr+8IWryWkY9MYs/+c3dM0XTjFb4QS6kPjydp7U9XH6F4K/qPmxWBEwSQ
UkCTKKd2Qt+5JPg2Xilamluo+FxjM2HzmqC6ThJXlloUHInvpvNbLy8ALFmWD4oq
9vtFCX9i9DalTlx4E2f8wvrwcGq8lnIV04LA2kAQFxaWyC6QHGwy4W9oY0uM44RL
0kEmB1+l6gUxrGqwBAbTfVEh47GdER6B1SJvGR3IHTatmk+t8fkbp8x9PY0P4Qin
XWr/xXzNgy4laxQDNDf5KGDorKAuDrEfVXEYmWvfsaPQ6JLdgbL82Ohfxs7lh9EX
nmFCnxQ2N06tlmNRZF8lKvsLRbK5QXJBuBmVFcA38v6jCAr9Lazc5rdeURl3PMv/
c2aexkBb206rHxbAP+dEnGOHBOnEBDR55o3YrFn9xJfy1qSlOcNatenEK5yLlIse
5Pqm57Gqmil+3SXU2ueCfDpMZ3qN1PLP/2P9GHuygwF4smRpI8wKY515aXDB4yTc
BUGAJw1Dr9IVbCnqaF+q9rfD0QpcthIb7xffh1tmqhU/p6pcoPocesQER6LmLnmL
16xJe1z9CDeYy2u+/eNuZSmghcjrl3tQJN1RNyyvU7d8OJKOFicDariMP639f0Bc
NBkxXpIZbNc6ljmjBD2VmA5LI1lq5MK8hITuU1pwGcBApetD7SPuwZdCWPfMsa9P
hzLe0AEm34ptv6+zZfymfbINWRRhJS6frwqM7iGtFBvEDgz7nF6abP6vB4uhdErE
dcWCM48XcNJunFEyq5PYuSj7PEF8aBJP2qi/16ZdeySB94CDhpvSjvV4CO3r6n3b
hN0U+vNkB8auZyh732TZnhrD6xuQUPr4R25qhklX4VxHmnUV5BnnlADGK2l4Q6bn
4OBydsuFGH4/1TrLosQWIxdTyQGA5MSI08XQeSodnKnb5SEy2zKQB/6EkG/8BWjI
vxRbELZ7v0vykm8XCAOLFutdekhpDi2SIAF11S5dxlSeS4xjRe5Gztd+zH/p9sEP
5nCRB2UlTLdCPmoq6hPNvHqmdjTIY5iGmF2xHzYIhY8EbdKHc9GKiRKRfxp5wg4R
/sbbkteOPvKMy0LWmpdgOVT9Z8fNCp6jLP01dXdccx/KJhmWknBiCHDOSzSsqy+9
gz7kNmzNrRBYc0giCXwl6Ngz21lcPAAIYunPImAKBSlTMyor1a8+tsTvFN7KmeR0
pSh4K8sNaGQRGbz3sj+KKPE6+4g8r3j1c9RDnEcNI7u7rgD9lLrGGkoHv4GVbmnA
qqgV49A4dV9KnXxJT/qzu0RDSKd3NvGZTLwqo9nOLbbucgp/+FebyMB+1r5b88nY
O3N0GvuNUTf2DIjoXxKeL5X5ndtia15jszb5l3f8kKNQrx2xr8mYG4vVpXczz/Ui
VVRDgb0tlHoJUpZ2GOzUz+auvwdjQLP/yovbLItQT9rFPvgFD0IXCLldSKIBhslz
+0FonAUomsM7sHwMnHfOp+GfjXKEOfwr7/4nkpmTaCVsKh/rqYKz/slLAmv1xZ8j
Miz8s6BWHvZVKd3Vfez74I4Pcdz/+v6ip9mW7cZyHSHldN3bEjSD/YKHYKz2Z62F
cMwyyfwq7RIf7wYV6+JVPdrec3U9GTnbF5K0b4dftDI4M09vXdeq0GVJi30jBccq
aBuOuqlMA+Y9aptr+6XKFdrDqbbct+R63tAiTWhqdNIMDCCpb2TONe4EyoD/Kb3B
0Ph1skq9QeuX98SlZ8B1f9GCOAFFjdKFdyvgxhvXwNL7oqeTqf65w47ZLVueGO9h
9yB8iWICLbs/+M4QtGhGMMGmKigboXoWAzgq1rUMeAarVsq+uWO9By4YUS5xwRRc
px1L4La/0a8OUPNoeZAUgMfgorELxZF6yyiDtc+x5O+RDMoI0D134Bt3AfgmVMMI
hNL51qUtkVmF4d9rI8OUqTVOk501wlRqMQzQxLc1u42uUI7yp8B+urLLqM3fJj42
s3PzlrRS+7pVz8u/04i3CoLM8WrpZ/OSCinHW472FgjTQtoQA4JR42ktO4EjwZkF
8XzkvDP1omxLrTAumEEy4XHie/FAiMAUdP2pbrglGaybL4DbT7N53DXD2Idj3FNu
8rBq6WhDw6yE6Uhq3wTAcpN9nbDk4s9lFodjK9tlcUPm2J+SnahDE5A7xkMtrSW3
n5umR23j677zSQ8+aTBRNKPwPDreoPrr4y4W+1cACAZNJxj8md2Vve9mxvp0TC3J
A+MMFwWqzO9IZseWgLe5c6+3Dh8npCwuny8WYfbgi6BFe/z/2HvUU6ZK1TPl0V56
IKm2Ls/HvUTp0TfLJoEdtgaVAlY50KhBO83hEaSHs7RVPKta4T53EQgLNi7L+4Sj
YSCoaexPvstmj2EwkUFMjdTNy7XznLnDxgm8TQa+sdeJNvXcB5jCHgBiB/xAbhXu
gPhBCIVpb9boKc11WRuZAwUUmWaDcfPhYR6Y5ldEpi3OxMeg9uWgZeDoIaKz4n8p
v5kkHKkSpUjIa/HrBHAvTw6Y/wx/mX91+Iclv69OvaHDN0sxQTfwEAI7VKMbJxEc
NIbUExFEI9JErzenG2YfuW16yIVMQbnIUfHbFmgHoIOjlPigFgNZ3U/mxZyjWs2D
NKA5GL00sPtSW7edJ9+LwD49R9Uqgxb5NzFYXrpxGH+gT1bwYjeyB4S/sdK+FYrC
eBOuaUiaDZwQkSlaHDd8fFenzDKY1/dh8vHUMUmNkWSqid6FLWMwT7xXXbQqw0El
Iq7GtKmZpwIX199j4LYR3zfY6+qiDJXse+1sMpapZ3cXz7rqLH1sk3TQWeQ4qAFP
rO8DdFOMAHAgm7uKT4GprTZSSmuoNRLal1caViy7d2VKBP7lM3/E5TFFQp8Ygv5F
sfvHdkdzaLHh5JSfPNFiWS+avpkjoq0ZeC1rt2lab3HIUINTr9XYkDWeU17NRRwN
REFd4z8fxXSDstdDzB8zxkC49iEgeXWPwqvZJ2kIep5IxQlk7EdsI3Wju4hnVzhs
yA0Z0o6EOY3c1CImx7XmgRliF5ypURKpC7Pwovkb4k0XZIuBk9N2nSL6isK/pFCD
t+mJ904fw2LVrTm7d/68MUdrAqzqsrEVtzCFvJq3xD7ThWrzIWhxPV76j5qGZTLq
DgDhFh4jqvv3vPW/Lme8rkV8HP+YGTAmnKuLg/5n1O3gZ1Ws/ennWeAyOAZVaYPS
JzP3HKrEBdxEeDL+OQBECmZCFDeJAMjzUOIY/MK3OyGMHsXco5x5RlK25H+2O+e+
yCUrF7iEbpMEeApKJHL2FN4+aq13zTcanT2ACQx+iTSFxHFyZMLsF7JhlnFfPZk6
wsxzi1k7sM4Z84LvfOrRH7fAdZVNZH0TMsahtH8jeKsIo9qSulxedWXXeHH8aKtS
U9akeLgLYy4PYgU5aSG2MUaDv6NBGuoAVuujRS2cqXZgcNlizds4n503lguk0U17
037f1k3aErxPH2uLo9TiaAQ0ZPx3aQPYNahS+zh/n0oMKTpAePcoPxxUIPxxUq5+
lYpXrPCSSOzGddn4h9HPnjk8o9onzU9PpmehJb1QwRPnarP7Xv7n4njWfR2xb6WO
GHIG+EMrZ3q9iZICW/QjbiJx1p/m7QARaaq7j1kWiD/BT2zuoL6pcyXcG+ZjDnvj
DYJqf5SJ7yjnOfpZ8ZHhOQd4yOg2BbqfMKs7zzOHulhmBRb6309ePqMY4V//yuXo
fVmH/8rY+lwvEapu9Cn3TzpEZMdN1wp7o+hPxhenkWp527nnyIi5Wy/wQKiQRn2w
bse7FniBuB55L5Qzke3KRrmgJgwbjUsKLIfAwVSy1wOVKoagl7Sk4AqIa0JHUZPU
ailEVdQe7f0PbViMAfyQj4FIEmdM7MTr7WH8oo0fxvCX4jp6F9fokvdnOwvVE9Yl
mdRxuz8iFUzqLsj6XbtSdvKsKay9mp3JCiq+duAZvmqprNOUgBqc20kxdsnOI/ih
6H/v0IJyWZW1n++ktRJrnDE0JD4EzxT7gKiJxGq1zhHoKFdl2POSXDMxK8VAs5XC
9nRA93S0bHTE2Igd2T1Fh9wjlAlztnBtN1nPWOJ8O8TyvBwvMehDBxc0j72t/aqt
KY9OsDPuAK0ZdlHl208mRjQuZpIs8QsrHMXez4F9RujgHWXfmXY7zKV8LsNwyUaY
C0CFD3fq/CcywFP1dqGpdYSGS6+BROdKGDattEA5KIaLTDE1e9DWRFrt3bY8ghWe
Rcl8sXCNwlTe7hrrixMWgsjsWKjsgVG9s6s28OZf+jqZQ7ck1HfQIzpsmDe7wsTK
LV57JIGy3JKVpRjLrSBl16zb9No2nRqJeNphOJcpF3s7JeKHG9WtGg/6m03aP6Z3
Hs8Iqbk7ha9SfzweSYqYXtT1K3XCCFBl/Mo21vapbVMD7ZeUwbXUmuBFthZ6bMlk
oJeXkQMXQzyccWiELWjOTZypE/vXNzfViwsSWxOV1Ny3ThJJ2Q1c1gC/smhOF6TH
cgQOH8t7Yb2lbtnoYywLTqFqLuthfTA/9HDLJ5eHtIvCNLqau8bb+QyK7kKNPSfb
gLdpRwgMxINPYCF+18OnjuguxxfAIe4Q0aA3MwVXhBnQoXiPBDWt5HBitVWCKGCt
dH4p2oZaj8wM9/N5oucOk6BtSxN8bBP4ptQ+RgBTuvJhaGLLfMKUVLuNlnxICv6g
Uo6pg5teFe7N6KZj2PHflfxz3MUxhXIos4tgULkYuJ/KF8XpNnlJQKevHn7TAapb
yFiNR+oOtHN9jSllZdcNvD23FjVqQuQ1DHo/hL/DkcHEfwKxCUNfL7FKHnDIThYS
ggzmXELE0MaSmCPc6yQodpJfPXPUzBsBVYp1TrQmp0cQ8jLFA+2Lwx9uagv2Wsdg
Auk6gzmBNqPz6SKvxTGOy2i7+j/S8KjERfRpKYdcDghZetxQWGzwp1ly2gbgNZeW
CMaV7bzxIi5zmzDiqKm873prIAACcz4ETRJvlW318ie9Pgj8uio9oSPj9E6/ionB
KBNxfhVyVNxt176z9k6EXjfyfypWM88VrLfHB7yxd5yQliBpj1bUgC88JFQDEOcT
8t8V9w/ZHaSB0YrrT5f5kpuMyArPiHs/vFppg4lgOpCbXfQpZeReosmUw+GvV4KB
HyeLf1liWpC2OU+C2XC3LcoFD/Hat2ZqpbyQBMmpxLwxOV3eeYE9da9hoYT7goAD
ztoJSbSkfaaG3c2UZChjYOVwARepM/5irwHHT79sIdpVBlG6VSo7ZIpm/8K4SVEq
909KCTXqSaBzjMIyi8uuQPbQ1eWdlLR01mL6+06Vt5qRJl4kidgeiCx0yUljbCDC
zoEcxTpZS6I7/oxW8rgGMJCYkLgtuPkESaBWbaDL9hpqgZ5roEc0b7XtvlU2rpMt
53+Y/ut00vnNUfWTjWESmXfG8i2D5X0kB19DHhpDw8qU1BsBfSbepFIOdsuamc/Z
Oy7svqqxNX4NqZcqlJtJh+QR10GUOwJyqiW/0pyZzWATl8UZdfY7m6VAenZknzL8
xBMQgtNwenFuoGWoybb9svWI52s2wViG8bw2soJFkQgPiRne5UQugaHnl/OWJ3xK
Bc3nKtnAlSzq+o01kUKYeem1IktL3/sUU37dyonEprRqjhoNgJN+uJcGHEoLy0rM
DbuXb8b+9Mqz/XoehrvAuXDZy+KRBqmZpGfSXAmDjo9P4J6QMQsh9KGFkyAQ9sYs
rbKkSN8r73l1pzLvbWF9qN+6CdrxN3TmG9up/jfXYf0TphU6kJNt26hi3h/4H10U
6hHQxxQznVHfewwzfjSHNZSgYnzDB0cIX3Mrfx1lwS4CY++2wGY2vYxmHzicdRxA
wIq+xgPa3YZozVduGbCKvHoyOH/HetuQxaYA81On4BxcaYjdFBTjmD+yUSvwHT3H
3mrSqL8iMtgof+/LXPQ7WUkj/p38q78BfnJQAEVcU0IAWMZO/Q3Ze9x61esvovRw
2YiEYwLnMhHICXCgEWM2u9CCSBngvrx4j77ASVlTrRCKHG7WAIJbTfh59x0Rspq2
Z4gY0xHhOV+KT4gpJuV41xZlQLccTHS1OKgaL8k7iGTcIrPFrEwVin/cFW6e+a9Y
Uh0NcEFOQusw+IixIYBR79pIDsGCNRKdvjBYllbgU4rC6rIbb/XWKcvIoJVh2S3I
kPeszKfjZJLk6R/vz8FwZBvs4OZ2V5g6sy7FS0qr1vJMI6OpFqAYL7ejeKKZMcEj
0tiMfSt4v2OvkSDMmW8sMU2MJmCLm3zGe//Y26VF1THSEGh9yh4V0DRwk5T7RdC0
1+O7Vi0k3n3LKRSZgsDh6JCbdnYU1ZVRQGJHpwH6Z6v2wH0acJAGglc+BN3o6KNE
Uao+CmUV+JgcakqCMACmCcwwm8Ilek3/MDd4Ot66cjA3ZQjAnfEqdzIh6NR1sS3P
Vd+kD5GcsNVH7WchADc4gY0rqq5fVGtVUHHXfj4GHpnwvxjJYGoHqLl4jvNJwhgX
urqQdvNkR6hskrRayM/hK6k4XD4nfP3C9uLcKafU698wo5HXhTSY+ekctg3yfWC5
Wo9wOhODg2LZGTph2XHcrw/YxreMMF7MdFLbrE/jiyP2wG0RoMhqbNMhbxWY3Ok6
gd0uefOBO56pmgoy659rJe6wat7JcYDe71BFDyZB+Ek5TJPdm0h+E43NGYvv5ag1
40UE6Z/SYdturN3yI/mYY9wEkwASVgpwwNoFqQUzwzonQEI1eLyw77SfCJIPNpsp
Mz6zz53SIA0ptyNuhY4ASBRFvFnDVM8wvfen3G/xKB2XOUdUQH5UpTfOwca/A20S
B7H1+smk5BztKDLPG+cZbKXYR9wUuV945Vyfjz4WNfHBe67e0k1PHmRg54XIJoo4
FKQ9um0lTkNMuThw2nYT8xADBtBDzFdMoqMv50kBi4vC7koLfWwS9P3ff5LfzQkV
PD+wzIpbYgEEuZzIE5IGdLjrVdYLE5IQ13noDaR/6Hz//meeyazypxrQvSpMuMLH
sHejDswkeYAcmLR8BspkuEV1mQUkx4hGN3ttp3Je4EqJxy2Dg4tQvDpgnUx8Zht9
Le13SS7/xXKDXnoBGVK+G/tdcbYYNP/AILkZ4GBz9xCPpLhz/x3i7ZdTioXnFU4X
/bG7fZYjjFS2EWMPaE4Bk9yhDQiBOJDCTIPkSBrRd9eEzRi7u4FB3e9pcn0x2Dk2
zCOep5D6WSxFx9SSx2U/D68vOqBBduvv3Mpl14qM82LxTlt0uLTnT3OJyTKsx295
U8Ed4U4p5C6/fk0X3A+CNIZLqLucCt8yDWVmP/rZJK1Lppm1hdlEOzf9g/F4sqqq
5I0CHjJ0T4CYxktt1OhGAQXZV9zHUaWw7GwhFzk++QX6Aim/TF/JTe9E4/n+q2a2
Ij0HzbNzekZbOA/RsxjZqjqWARXuC4Gzn6kjxZm/LTuflWd1ii9yX1+wDEKwi7zQ
5opk2G+4llPNGIOweQleGi1nsVW3Io8NSXiNX5mnajJpAwutASHoOOsqnPCcQDng
Yx2J7ByNOZOcHCKNYP1lWqJLNM4XD9Autei0Z1YY0m2h6FdMm3dsmnEoSr8ug2+Z
20y6/YGFSRXn1WxRMC15BJqLhCyC+LdlRbMQ4+hw61OzFa8H6Cs/5FudxdATlx24
3Aa0yGmrrcR7vzjLQLGx9hem5zWsEGf2QPPGgB9CS06bmHzIlK35yVaOhc6qtAzQ
mQygxHhDwUq3J+H0f9vOwWtlEpBVZ5tinlVUkbmLRHSAhm6J3xuE7lrCxkjc+0Pz
g7fZAb7ipIwJbngIvlgxzLyYE/JmdVmVs8TaUAnMn9qBuFaKL6wC9uDpAX7tlc8C
2xSEuCqSr6mCYQCX82vpCzxvw34qTOi0u8R9eGaQh8NQ/uhvylcBcHBpX1fs8mA4
fNwZVeDnPAsIKe4KwyYmYru8kAPBit3QPBdKzRkXA/C0MDoi8Qy3FR7KcZ2V7z7v
MO68V8uWta+WJX7a/U3y9yZIhnbWgcnybFFsC4mCZU/CtXPtQYQ0FxejFwUdH1P4
0U9ZXtkU5G09CcB63TQwHIQw9vYTTqIPfrTK31RiOQM/jd30+paroYrjgWkMlfDM
gWug1EhmCinme/1mjcy8B/7UgiZ/PT7u35ym6U+/BAAx1JyE8v1ZoBseUxfaHEhz
MQXNRfWGpb8HOdX+PoQ2CtT8odfTq4jm0DPd7cbbcLxrDagOn81iyFxcESKT2GlN
4TCcwE4nV+6CWLFTtEQGBhvzJb0ZV5Ii8OVL2iP+fdMoml3rgwfnTH+pwJynr1l5
3W11/UH2p1dcl5vwT+fHFdSIZ6MhQDySlBOcz2enFq5uzW8BCaadifXdXHJZk7AU
S9EQbuPiRLre/v3AaVK7tpMrjtQ0enhjAhVfOGaTJ4sW9tSCTUNF0s8Y33JcXCFC
0VO92h9g8652hkhUnAGHx8ryn2U3jViZAbebs/yaGCBn9RuGH53DE0p5CyrBtgXT
0MRk9sM2KjEskmnKsYyX0NvkyBjEfmFTh753qdtOcw0TWIcbOyUdY7EdD7gcIh7j
sgRDKhJui4pfmmbT4hlRf/4aBsCvZyzGvcf/vSAXk5q0elU3haLiJWDFne0KiQJn
WIqKNXRp4YhWc6/vQnqtfuycLR/zTQoTH6UPpFoAu08X+YtfBiqyjQpbGqZy4BSo
66BnKVrfLMiKuC9kLm/6mpOKlFSTrLJHbX4QfwPLLsoqhisupSftvnUP3aBreNy2
BN4ilixinX2uleBZ038oaYnuvMTmSOk2PT5G2n2MzDrTjVya+wOFrVFLbEjk0OSH
abHVoUdv88RFQk+l2DXSU22w0VuqkEcutTsw6mTooE5koMDnD8/3MQnahoz0Hszv
/N/Skkke2VT55aD6VYEWgB84QgiLfLUn91uIxcrlWNpkvr3sxmBDlOaYrNqTkIsr
nzG6bBgVh9ydkBnuGb+x+owciJH8cTFZJWPdYsaESb7ySt3I6AqK9tWNslyaQELL
Jany3QVpRe8L29HXPGX1k/A+oWcaUyg+KaTAWn0hX0Bo8sLDggkcAjZi5FFYU15F
vqeEeXYLiI4ro7g8lAAb+4tf7lI5yrOHmzNLP/U/PcQUFKFt7t5LVc/fpb5jXRlW
6dopiSG7tB0SN66nKhTiQ4gnSbDOFcPmfPVJY03mMInff+mrwi4uJSq0sKxDB8W2
9Ez6KxhC7ZxmSxjOhWpFW8lhF54tw6Q7w/Ijyp81VdGffkcgF6O2wUZuXxnzY/4t
XDCjoPxqR6z2dER0vrZWmRYu+dlJ7Z7gQXYU7Ia+w2cvETLutV/DtMawWSVu0467
oumyCX8c8p8Cu7zDVZs9qIOQsgfNnioEyNpAO3a4duzMszwrBOY68be6rChSangP
13tnAoAF9QfvVuz4phUnT/CDEWVk3EQLTZ/ZT6UPIYO6K9TBDVRfBI8rvBm4BC/X
j6xjqmnZ15rhb0+97iILzG+hVtkdIUEIm0TIpNc/dEg0JB+ueYJrPB1BXujAvcpz
11xerFmQUa719mho7WKxEY9KYKoGHo5/wQbIFqonSJpH3+gWk5EKW8LdW8p3mtwx
vJ/hr2JxX4qtzqcsl8DQz3sW5Y2akHXwaSeT4ab865upcSf0VfRF/tRTvub824xg
FIkFYiUw7KGLh05/zoBPL5VLlU5YLzjuvQSdo8AwiFoOSXPzt56KkgNrlURlyPgL
5ROShwYpvmry6OfT6upor0CwoWrdYVG0BNehukjWtoGy88ZdRd6unZRKyjpDq+OO
NEYmqHT2oPk8eL2yEcM6kp/MXnlAT1fohqDOI5S6/FjrK5tvahhTelvwnKERAC8Z
gAPFGi+HS9zV5jj9297Jp+E5d/K0NYb6IWc7bvu8nxNk0xMahSvh6C7Iux5cs3uB
oJE5+HJd3/XHNhqi8hwS7ybOVqF8vqaIb7tedzARhUFvUUmo1JdJ0si1CE1gnx1e
XVi6ibRVPJw0dDSA8jsM9O2gVSOhvqRW/yhfNusy3KaOCKuiSi2FQi562FBZgl+P
hZlU7bwqiUj1pFS7aSWOJEpMUTIfJEtPqUekJPfdMEgiJmMqExPZk0SB93nqNUCJ
en8dAOsNoQEfRMSZzvdwQ/OWyomgnfls+CRmDEj4oCKoNLa+m3cybZ67ot3aYWwy
iq3Ks4YDPWcW2mMaLJ6lFWzGysr9MNjq7Tz/VBUJeh7Y3feEANk3FsmFK023fFe6
WsYTNBpSzVIncXNHxDI9QntClus63uOd7F+UHUD9+e0QchfKkQpdB1+qHgOVxUrq
mitDPR2jCpeGIju6btd96lNCuPoU6d/r/aYDKVwXPlq5T8ziTCPxxKtm5YYQ3I+5
coiDBh5+BLlUIyDQzhisPV575Qznh0KHatbI+QYF+eLIgbHcV0pwhKma1p9kMmOM
McoBijlVcNYbpptYusQFhNP7H8x5xpwOW2p5fUFAtxSuN4NVNllisVb5c5DN8KgC
9UGi/URFXZGvy1pElJW3fkjrmz0y2Muk/+2nwuig+U160wspJgxClYIHmBYPdkf+
oKUhdkIFy+jtWSMSqC3QGXrYg+jfu3aAOmMlJPi4isGIWVu6+HIMrnydNKyrFP4n
rHYxFrj7sLWAIe5hOsK81CqaXujffedJHY8HRfhRAqN+dCEqr28jMtGO3WsOMLpT
uEIYXEYS3lslb8QSSVHiVF6QU7YF1gdum+mef+b7F5wXDClEMdH4loyTldowVCWS
R8mkkhqhN47s7D0m83TzuUmliAH6XpSJBiSPKP9cevuw4SjGsHlbWu2KgXqtAuNT
h/eYhQ7Oe2dNFZoewxbjtAxBAvAfXw+p4z96Tw1VQGjgT7IUhHqr2GJ7slBq6+lQ
VjF/oNcxdiTHiVAZ3Pc3oc7eeu/s6E9rTcrKdPDsNYXvEnRJFSVGCYpy4RhmUyCA
1zFMS1WpipUlgABFc4dE/FWU5cJBz+8tHoNVBm/ZsmCC+8ozQ/CqT0naxKXkJjEt
gJSfyT5FTXyDiQsawYEIYzbxATSHdJfI9tgHoLK3QB5qxMSEMbGMrQwV9HGugWbr
h2lucRxemK8E/qTyWTzQtY6z4Fa5YRt4hS9SiACHuOJo+UMcihHxaY7+mfc6D83K
wI/nL1me682mQg5QrLwm4OVOhmgtdSI/wJMgkf2PWCe9MyngWw9Nd9MttBATWzom
qd7+P5ZQsjbuOf7P6SVpIYO384bJeIbWHjbALKs+GzOTo2CVSsDzErB3qAjBkjXe
5hYr5xMVmFeSawhi8Vifq3p9U9J+zauPLp+a1I76tm0TLQ9WCl5t1VRjF+lkSkKW
2h64voA2Zp8rO0mwMlRAyW/V1A9aXAW7Tb1/DhpoowsHG7lK01XPxbx77odLeBlE
SrdNtBOtYWOcSFKG6nxCbk1Msj5W5ZpsUmevqkBH5VKbC2bIPVh3o/1CFFx4bg5u
JaPOr3s53oMQi3nO4p/vrbXVwsIntC6abfF2g0ufL90cHxBLYTsPE2rBLi11y+32
7TOlVgIOlsjQ7Z+cGbJ3tdCfsi7NFn/BMRIHOw94YtHnO/DQwcDUzFvm2DkvDkyu
B9bEChoWQVFYTi4fW+EX26jL8rCT1nClSYl1sWYZhxJJuYWLYUWrks/by45ih3NV
9P18zgMCc5mqtsYRVWYeVJhvH2qUCz3Hm0TQ/v4wtz6JRMT4th/Sx8MK+Bp8asa/
tukDNlAf5kS0tvt9e/4J7EwAN3MktBnIgmnMP6khyKtt+CnSfaSBzc2hc/GDsycf
thLanvXqAQGHCYcdJI1cdR2vQg9a/X+iW9yfO6kaiC171JiVuBOHHiruL6dmgoX+
eZx2MTN/K6XN/D4SY52U/V9Egp5aF2LFEWIxXPAUYkcDl7b/51i3O6JxS6CfiIjC
qlS/knjTvmgJtbMMC94evj3r6PsSDhYB9GKmNu3wWP87uYNM0tLfZl6OddbyWjMm
r0TJTdoOYtDGV+mi+nnxxvOYHuB9SlGkqxTB7pz+U1pSYKzSsbAIMFR7ZMw950lI
FiPA+Pb4B2xDNmNv+q6btWEhrDLW1iSvFhSLzj3i6F4zXsqFK8YmjxflKMTGUPx7
AprEqtEHppDwNsZowfoJNCwEjamVIZ0xJpNEP7LZvIPF+TBn74xwzF6PUlxdxOMH
g2i/ox5bSnGot+TqzpkRxAJDxjoz4OJoDcpbKSp3ykpu8V8YqNmG/WRuJ9/l1DU+
b39K3HyC485Crn1v/UB1nmNT6ngMG+3iJpFqwTplClyXpPBuSk6yBXSuh6b0H1mt
S7/1xPjg5mJeEAo72MxLCCn/78Bu2FkAJQB3A5i2fkXLyNYDtYFPJfX3yCBrQ5Kq
gOe94ArA6yu9MLGPI0ZXSPln7Qi1W/kewpMZdLuyUuu1GH/RR8K58Ag/GPipiURo
1Pm4bpKOb0wAaa+NgvUZJ+IDULYZDsvwHsBtlcfWvBaJUcgIE+iPHPmptZ02Nk/B
YAX1PkaxgNfYlB8FRdxgv1tFSL3nwBzPYFZE82rtwTZXjezgI/filNNkn9MUaHlD
b9KzNIuM0FpocuERFtCtHylMyY7+Vkyh3U5Ni8kTSQPOd39nsu4DYu1Ye6qPysTd
bC+Vj7SBbsfuFafWWDFFfWt79K9XR7Z0zTxSjDQqJjFSAygFykSprX1U4fzygY+5
wGYwxETf+I8b3nZnDwsVAQmLHKqT2ty8MW8+aiEwycgYgPB0JH8dYtXYx0KaNrC1
LnHrDQbhtEyt2628jyyhdOSVsFF75TXdvDOhw6vrOHjV9sdeLbr+74uWiJj+Zf67
icVZANlsUU81yQArHpeLs7lqt69Io1ZNSPgPraV8nJlV7J95IPwi6KIGpQeK6QVe
xzidF/Ot2ta/TbCMvktbhw0wKRSDBjcVq8zkHDokyHKDj+A6MSayFiefEk4bU2n6
2U90ZdWYSu58oEEUsH/dk9J7Cx/iEXIMD2BGebVs442ANaUCSjyd+zP2UZNAnOtP
tlqVn5O9rdhrKArGLn9FYO3SqUNqxi2srcWXcJC6YPozhMomCPkZaxiZXfeNNhbu
wiJixVIjPflHbh3ESENbQ7oI3uxlOlWg7C2v/KcBOfaMm/j26Ndme4SceMesDnSj
4OO/0dGeacKEMb8mWW+Ysv6girIDheOEB7skT8Yw61/AJ4uoe9TTOugJzhOefE+H
SIguk9hgmoiuqhimR5LybaFAFGnb5FdZv3L2S6LsSrNmYRO83fz+LR9qWeHWUnFB
4b7eAWZOTYPaYUDboYC0JMjUnpXhDkujLTNxkrzQoxJO/iKotcJtToqfTRt2mfkx
ry1CHhDikezuJm0xZN77VHNVitU6JwgqxUuiH/uIzgxDYJrhxbTBSvRqbwQYak8q
tTU0efTvNNtAFrg160uk7B16o/jG6pOztJzpEjTHGWajUGLDMh+SR+BlXeAn8Sng
JEbq97j49MrUHSwLxVFuK/c1q56lpHZfJFBDI3K8SOKgkCqgXgqB6Id5SRuiC+0p
EQWCz5xmBZLCPDWfqEL7FXiwPHh3eB6YVp5v5GNm92oxDPX0sQ+21AIUWXbvAgvJ
SVralD1VXHDWSZ098+nMSy9kVD//pJZs/xAjX9rtfnStN/X+xrNPkoI2CNjP1Etl
E9EJLZeApOoyDkkmGGgo+qxgLk9BziwFa4Wo19TJHpxjLyIRpddM30laiDf07MNO
ncJtacAvDQiPaXZUy3WwxKB3LwK8cr77f1db6jb8o7Ts50LSwd35nGF49WklwfXI
hr2MmB6U8iyzXAv4IdCGZSm5jn4245giaMdIWtXeR7DAmnYaZMljtBPR/dz8Koe8
SWLqCS4Xyw+StEvHZcDaWRzBJyoHgthZ7wySkYoT5IEnqI3TF5zCcQN5LrV9GWgV
Rj0SwHswW6Wckz+HftQl8LwUaG6CWDRvbmTnPtMuT1ZVt4S4HeVvhnZtOIyDZt8y
qYpACPcsoWpJvlXGQuqJEIDdDqwXNz6CWm/71s/PfR2Nxi1TxBvcmbS8FGlQ+w+s
qRjhFIU0KLLtuzGz6wPmPnKaDkzgiGK/69Ti+duNVP5X1Sy+P8aEc00ISa6uYjrt
SOXBBzw4atwLlGt85YwUuL7WsRC0XefWSFqo5GK7Kq3YaY3g5Vi/qE+GKpzzsh3K
fv14xpUn+Iw4Q82TWHoM900Fe4yD+C3fkiSF6Qn/7+iGgxCcXPA/k/0F2GipyH0v
L8coFuGMAVUiCdinaDh8Re+0OP04n2p1HvA0IQgP1R8u5FMnSAxm1I6G//SCxpwe
JIB/k70WdkqzcIjLL1RQ94akvD6uQ8EXLflpnnDwAp4b+7bKFK30+LZ7ryRUX+Tl
Xvo8Ce1mWCURiqpa0sAL+5Bix/BUL98XYbV1AwtbZVRMl9nM9zwH5s0r5zptVxLP
ANY6YtpRiaLO4SJ9yQjVNCLiXgDuNk5DiO6a2s18/Bz6vuFOpDWTgLX6SW8ifSXB
u2cOaKuCJ2IxNGK4KL/rVRTaPUrxrw/VCN/N+orAsSbX4gMygTkc0BthHnANVC4D
zWE6Ap4QO5L5LTWv38ExhB6QOOBuCS5H+J0IQfSqxgK/wNpRsge0V3Vs7ST4N+s1
ZOXlr5HY61/1jzGSepz9GBeTLSRhCDNO8NUhEnxOYzAiNXlL7y/G8g9gypoTvN7P
K6ujuu4Ui/4tct7n2AY3e8k8uRvvVPYm+rPRNIfU/M+kJ0T2k+kwpMctowwtKjUY
OKhpALC+eY7l9BYZYKoDspIAlVEwnatTjG4NvNS8/2unhswrXVNJcl7NdfTrTIUz
ctxhoCw5H0EW7wCawlTiyPGxVUKmRf66rY/Coomr/aYG1gHMumPUliD/RjSLfjyz
Nb2FKWwvPWy6PYaCRXb/41Msm+zmUhVedEG+vNiaY0/J04aw9BgrrM974mxlcd7z
s7gkQsyg8UV+CI/qMMwiWOaVRoaGTbwf3Q7Dd8Tr6mhutYkygSaq/xLGjXP5eAUW
CHnOo+aREewnrPikoZzNQfyU39Wp04/4Z1pI5qFMXjsq3hO4xx/orT1qOSeVfkXU
sje7hTvXGebOpZbSOSTsoP9ln/2FsmC+rgQ8BNoDKpVRLKWZ/Yg4WPjFYsseFiIy
fGZN/B6D4PusaM/irOCC953vDPF3o8+fIdtLUpHhNpdAC/oYa8LElpK1MiWMPFY/
RUqtkBx8cyTls0wtpIo9z9jHsr9Zpy0EXfm/oN6sNvzXJL2+5kivRUl2YPEQ9nDt
0jCq88UgZmZpEs/QUeRGxEAoDYUYF+asBq9MN8rvrUG3Dj6p2C08UJa2kyAGL11N
hKssOqI28BWncx5rYk9SEiDg0mtudQOwjAsYg1xG5WxmqMZGCEEhhCJsh0HDNaW2
YkvPjsKE7bKNRGaT9bSzyJFTA88PAzHL/2PBrR4hoxCdSMemNvK4XRUlTdWoaIaN
ECGTkvUCaLMQ20wTxZzD9dAliX4uDN5NLXusV0o6YgoJQ4ZEDdwf2Bwe0tE8ti/l
gubG+D6tFQfNREEhhRo71ItZg5s93u5Z+ckoHPy+gN++PtTBoOpsOfUfHCGXp4KZ
DxA+7g2NIYfvaurVlR/zOsUC7UKDQxL975g0O6v1eJbrYzBfjJcv9jMVOpLD53dz
pCBblEHOMKJlVDlLd29oD1PqHQxM0zqOjMjF18DEBIiJhOUvxDfWz1jEfJZvwdYO
JEJ64WpulwM0PHsD+q6/RdL8RhB13/4rPJXsEAKO9lwD8mF648zMmjOUNrxEvvQa
ilAVv5ke+StQBTzIznI26jv3Pcopz54B5hPmtkKLg1NNOfTYTHADiD0xPM+Wqqg8
T6WhodPKXv0h8EA3ieyWyJi3UT68Ub0IwurhH3Yppblcd/EOtJ27s81UHTzFQjTm
D3FIDbhGeGGsOjVbHLQ5KJ1t0j1cXK/RheabTEW36XDG/hkFPeXbyjaN226UAmzG
+QrxqXh9lpyQwAuIWrinqft+XxGFqOaUm9eMQ2ES/nyjS30+QwKTn5yo4FDV+iCp
GP2ovW3qhLhKc+6gqfvlzQIdGeJ3FchN4tqusDqFczF3sPcDaGyIqleju+qBMBsP
yOWRdCK5sQ+hYMGg2cSATDYmf7Tajqkn2iWehv9UJugjfnI2HvMuXCv8g49YUj8U
Y3IhIiFMlquZW8m3e5SZqE2aczmsufg/k9e2L0AIjMxsPtrZ9HotJx+7nsVVsSQW
fuB85J2r7A46ofSKK5TGEiZxr9feupXf+4UqpRGDrJLrelgUfNSgVxfDExO6UYAR
5ac4B5YsfIQkm7KmBzw+r5+vu0PotIdsvdPiX0FTACjTl2kheEM77Oeo4g0Pu7D1
DzDxW8abMJ/2hPenUThS3lcAo9+nYX5sw+9CJWJt/BJghemwVxgMOKXn16JGo0gp
Pu/G+X7L0+kWbZvOEmKAS3Mk9lQbhswoVZmkte5IcFoZLPEbLQyd0ZTdmslmj0g1
P6y2aHWzQ2hWGrG63+R0Z5sU4XtEXXTidP4SJe3HAzwI9h/vjidU2zVA5DaaannJ
cqpttqojEPqdd2ZExU57ydSjuBy2UTxo9x3d0nSBO3cNMrfJ38SnSam7eaWxHc2B
5WyDsMe70fL8455WvLU8UKpZQ//Yl7AhWqrK1hOboFGjmgqyS15e3iCTH8piwMOF
dm6FQRkjrbdPUBlO0khlvPwtZLwjYg71yZE+6r3ft/DIEsdd2ePaKF25sMBikmP7
1O7QBurZhlg7I6dRHN8H7cwVd881OyP8oc56AEc6YLt3pPZlHcUT9CGDIj/tYfK3
Uc2QS3HgrOofFJwCqOi2KYw61cBYq3i7TksriY1AoIHbK9D3nRfORjTh6jkcpjVz
e9D43bpv+W+8pabEbdQ1/Su7zkXybeB1fF2rTi8Q/vPhR5vvpfA8tusGUes2fkYR
t/KOnVksPAbF/olIzcyWQnezDVMvwIZnxaYCi+BBJdbZxALz2nfiFO57WkwoH1Ik
Hz17z0cX0Itp9pmhME+mggZKT3QkL9z+6y6f4nRRwKivwaC47IgOOMXNCkkFm4gv
d0KztqI2nu/AdIHvhgz2wYCyffmDXAokbJvEI2LHj3lRNjYmZoWq4QQtHsbRl8fi
hCGdkQaOQiIg1IyGFIYBvDLDuvby6hXAPyS7HFeR9ViIegV0WaHaaUZcfmvxSwZE
cp+K86vjloAAAFg1ytzThaCesMpP7ioCjrQUD2udsOWeNMBUAwA6R5fSLq/SVvFs
Y57EgGP2NtqLFyh/SiM59louNSuvtXIGZdD9bYOKcHdLMLT3aH12auIbdHrcBP3a
+Pc/pAGldJZLFtPCDZOVk3ko/R1NfeMDU66PyuLAy8xI5Cr9oRlDjABjnYTpF4Fv
BhdbZb5Z2NnOwjc2TLPViYalPUaZ3XPIYSuchOUgRR5HTfrQG5nXajeZk4Mmd75X
At4rs/17zi1cox4KSe0BC9Ok/Dr0oggX3zctkMEPNRb/YtKxGbVpED3QZvmdJner
/7N7qFbrr4vtMAMjTZrqpoNyRAovbQMZj/OVousah0CJdROoC+bA46HB8nH/Zpxj
l6jlzNq7Zji3YPfOG57c7VzjK6H/+agpH8EdnJbHQgNLmzeHCCqEVnGFzJ64CMdI
no5SJh1qw05biZonnWe5qT6OnYdJS1vSU3TNx7jzXpXsJZgaAmRTkyVTAsTB1cX8
EY+uG2E1gkixd1LDIFZwvpgIagmXdkMfXWWqMmqtqSXj1ya0sPmISluGlgx4tyT6
edNdkMakwX/P1oBdXGb0phkanVQZh8mZ3+UdDS4vQG/CYJbENBCjfNXriOIjFsSM
2mJQqDOT08Nj/oo9j2mHb4rCiKqXME0y3rjdIm9bfi1JV7tWgWbmIwS5jE3ubMQQ
qI08Zq2en3Jsg9NDXOWQUxoV8pNsJThTnIDT7G5CvRKaB7o3i5GYR140ItPJtOMe
5mvC7+plrmBQjZmGprwfJ35Gzgjeg+MWyHm9LtFY3qCysa9LLm/qzdc1CoC/rM6C
7bWgUAOZ3WHc8nrVxMBc7FjOS4fDbCmHlRxXcFacM9qIdFwpB+Dq8PcRtFX+R2tF
wpXwZ45dJSKZNZ39aBgWPAwPSg5HfupiOOLfzpx2CtBLmMWSGJn7ZSVCJIuJuvrM
zrV20kJfP8VyXGKXRkcw768q0tA+3eZFgaBjz0HU8F7wyzS7SjGw0Xwv+lG6wuW4
BjUaJuTwphsgO5sPH3utGYNw1LPE5b6fUkG5/IT808sbQhME85xpVSNZuVuOjWIe
1v0pMRqQfirfmWJpciKEzXg06hEFkzWKPy3uFJ7jJ9+HToCegKX4Adln/ccY/FhJ
W6a9dgMijVG7xy83nxz3i4Ja0ckJvgcNULjMe5Sr7pnI+/DsXNkQ8jaAyN5y13c0
ESg+y1SRYso4vhlwe1Gx+KjpL583kE8myeA0tKFjYFkTyoBoQeWxsQZOdetHGwpx
2Mb8/9/THYwaCPNL4RzRZXU0zke+Dye3FLqfMvePFRyr3AcpbyJqWzVfrUD1cEJ0
r4LFwwopsXXcpNcaw3fGSwkNLKDm13qROafDZZM034I/eghIAiywzfmcEGIyUkol
37PFnX2hysNaweNiQQICcnVw+5dG48RuM601LkkGPw9QY4peHta9kMHiv+KLRA8/
LYNjktZvPtyhcdamMEoOTXwUsXWcztLJ0zDbU3QdDcCdxFTRkKOPr10+9owx4OK2
GqOevZbi6cXco57N90E68TbWit+0B0wzUhyfsz0vGTK1uZ1TAOOPpiae98FDkV5/
W0K2uRE0zPkTbHBIOg5jPAZxBHLd14CIaZrMu2Hk76VvZJYThFYP976/6iGNN6X4
5tdyUpJwVy0VG2g4GkvzHGiWYEWmaq1zyXKMoHBzRf6/stG7Kw1wl1jwlrn1Ub29
VEnBGzq7y1f++sgES0p/ZyU/l2MmJ0gXjNiT+lo3+ZG+HIV7AA0oxByx2sRqp0uA
MjL8eKMdNhFonOgGjeXVeWxYyWc0v1y7ySKeyU2j2JlPRuqaWCXBCAR3xA6mh2Sg
Gv8/3IIj4NWPS/Wo1z8lfmosKXYy2zSTr0jMW6PIz20D51ESDIYdoOCg7gbphpA2
vM2Wk/axYrTF4Kjg2aZUZYZRbhbA9Mg9xvqyaFZaWOA+tTsKTvThOTtIWV6makYj
89QFrT9V/Ej6+20C3XR7o/cc+1/cXZhMZJj+WcGI0jn5WlszgwfBZ1FuoWvdvrUd
OkTgF5Oi2CaUzNUN62rCzUgAk8kBhX0T95biQoS75nN2mywy04w1/d00nd0MoAs8
Xn/dugKa7Tajz1ebJocvpTkWMiqhjJfK+DL3v1L648T4wx/qtNo36sQbPb8QppT2
lV2No6evXJEQgl/2w+P/uwJ0oflvmq+ExbzuOKaQBPIBiJAJekQecZaZ05HQpy7o
SveWDykqkLUNk2sOE1Rq6N2vfdNlzeVCgG1LHgmkyGZniD6bZHxN46Pv+dUci5E3
7P0Xbi3uxGfjRB+VtXQCpxlSv+4ejg+goZGACkh0VNuU527AZWXC3/IFumIFtZdA
cJj1XLrzhwD3xEQskiLcg9DiTY2m7hK7wfqTS6U3mBBHTgK4L1PDQToLJtl3U1et
iNQgyai62js6qnrIfGrVnLC7LzTLnJoNwkHLYa8Tw4ApGIRe0h7BjvtRrzA0tBtZ
KCt1fMvMNk2NP1er9Kk9f+Dqd3FGvOsmpYXs3mjwIVI8uURqXwbjXWITpZEmp4fW
5dTSGjny2hFXfkpZXa6QeUIruTF2ErjrSiG3AygpDlrxhC585Q0LIMBkizVvth95
vbgxtlmPhmyTGyCd0JEilT7XkxQCYMM/bMhgEYGfebgW4hzVibXUAYjXPSxvMzCc
5fKHSKHtJprIcvrYJTEKl2qIkZ5Cn36tQWp4r5sUR6oQ7JDPFOoj9Ki2fosqNpNP
JbUXEJj6K0NRbyjRbuWoAGbUOfWQQiIU6o88Od8J+3DoIQJqUFj7XIrr1kyCk7/z
EwVFLywzq/a5Wg8ABqcoODot2fwr0s9o5y6ePNgi21lPDnO+l6GUD7ZSrbYwT4bv
P0HqTcRcvpq7wG6m3W/BbtvYhwxVIkpfdY0bPziCakYGwRFxkKu8V7ScHImIzK/E
wczpxyHRH6lWP241zKEwWJYLI0WxEXkOIE+IaJAePaN0TMVZf+MF7bmNrKd6vyTH
DB53HIVAYt0pBeeTB4RrduqklcH2FON54SMoUpdj5Lwhn4Jj0WnWxqgPLBliOEB9
1mOP0k3tdsddGn8b1EzIO3Sl5cumi7KM/+a55RCfzki+ku1R4OSSXnGNaZVWsDuX
MQ87vLBFk8nsTCIoxF4YBQhg/UrQVrjitU0WDr+eedwrllAxSC1MMT4NeykCEAmD
FvbzWRb6370QdquL89z2elfxwUI/vsYJNWoSV4pgH+ZHRUNJiIz79Ihch2pqfORz
NQlik+9+JdjpuhRnFCQ063a2XKoDakRYm/aZA0pZX/ghrW52s2VpCKEjm94/uFbx
ipp9VgASyDjaU9bYn1v1lGbFOib2y2lnv5zLpSqaIto3I4tVGXm61vntIHmzdZlc
9kCYVoOwz+u8JgNmsTsv9fYCjroIdEEeNJdz7r/2+CLpLPBx2zVINVeatswFmVcl
NEIkwRXBdREyQ1C55P84e4xmRjenXF1GSgLO/pJiqiWpCfAzeGTkaIptM++gIdMl
AvtVBAH3HLckGAJ/X/tth8Lfw7wpu4HOB7Jh5QYqbA487SOoso3teCiD8VY/XcqC
HAtXTuTNMvOUOJLnfz3oBlUQyyeD0xQtpJhZfm7lK3hxfyd1957In9a8KC88WZB2
nYcwKQJ05U4zr+ZzvYsvuc6v5TP47GxyU74ANnp49rmkrCORuxXWjGvmdbWdcpd6
cs4rKQv/LQdedb2Xlp5VwiI9NF5m25PqH8HA9Axvu5hVqfvtnNVGxQC6sPY2/LBO
vSYQ4BUeNzzkwiiZCXSKW02JbiQNDIMqvy6LWoPg70tyx/PoT8bi5a5DrKNVjPk7
Uqz8cDbp1hV8tFB+kiziFonKYy6dj+ECNIBzk1mKM2HFDhALsjM0i0ke765xI8be
TqaXgU6wNYEps1xdY4tzBUvEtOQeHK6gTmmi8JARB+vpg97AyzndZe/s2IEFCY7b
muh0OBVTrS10ueemAimsNacmRXCGRb/y7GxOKTe3WrXUblgbY2hy3B0Plzkgnw3e
0sjnNfAKKpSME1KdUYG+QDq8eV7n7voZThgVtwYjijjS4TzveDJGdkteUQzmdHcg
xelFnzXg6Y2QT3zM4b83E8ETQRwKTAdq8e6V4KAdNrb6UHBYk0oYHKPw82W+tNdD
DEjJveuYXFXPbqUOu/5dBMDvbY8Qqb8ZwNfm7Uzy/Bambm+EPxFlATe8cjzZegxa
G5IOsrwQgeXJVG8ZTflSQhX/8jEeTUOtuESVJOwOTC9FdXAUjTrQiwFfmjAWq/cf
Dx5GMdNK0qS6n8QJ4lFgM6htYoPhKJpGbxrgwFuyd0m0bJGrGx6B4XpBDD4x7w1Y
t//B+ItGxWS5CuYo6/KJs3aZvFLB8NWpLA5G6ic74p4plIW+iDoJ/nb8ACfWs3mh
w4QJARYNtRlnMpHqh6GDtdDFdsgFh0DR+TOcAY/juWzwl46I/chFEZLWyWhvilo2
wjYqnVHkxTll2+cLKapi2EiJCsv1g43TW83OIlszGVANcjvsPzXEAJWZiRFD6uAX
l+WVZvXrU+SDtWLpC57plHIdMKJvWhYuf9nfDquPta3bN0hRImBTBPuPdSwKV80L
ZTg8O9CCH+jm4bt+VjgnITrhU8wj6D0jRQhz6i9GocEGlj04pXa0TR3iUMackUUG
Od/LrFgqSCEBGVkGVcJ4gp8GBZlAsZRD29+QEZQ/GdSVWF3nji6XK41kkpZFxRIJ
FaZygBLJuldQpcpuBVImAhU1HdU8STEDj1/rlbV/hSra8z3kodbGz7WbgWtPQOZk
LHe+HUxF1GqAbsk9Y4Tz3LJ8SVvApFgRbmNUu+7Lt4QaAwnCgUhKuDy8KBgxB+a2
wKN91a9zKhLNxFInRTFiK3Q/C9HX5mR183y8ugZfBmNQuvqjDWSd+ydrvFUkC+qM
uauWbYXXcIMxkdQpCR3PU6S9euYpEKfdp3H8EpxCFZYcsgeRoVIWxYBpH5kk2VUv
moryvpNvD6TrnF+PJnLrW9vrpgDNcdNHHuKKHt2evs1UgkTaupFAvvNUFCliQrN7
e0adRBNsMQW2bcPx+K5kbsXxQgX4AGZN7aslKtKuAMCbBes/Nu5bA7b3SbJ1LfvK
I0xj0tN7j6u7R2bH0fDMKlI9v8DhTMsKjp86qmMxe1848K7dFFB4Lm4U+Qr+nW9b
/n60N5HoPTD03wswi0zdx80thHXoPKRLTtebnPBl1lewBzqgPkzZPik3xsaniwt7
MHX/KhYpJr/s8aKjSzvzPVpvahqW1SUA25beS/SH4J4+vgnvmKulGrVt9Wj1B5QR
FKq84yzmrHVdKtVHh/gVpNF+Kcgsc3sczTXF75lV0XwKUoaFx7N/JcfQoWTvI5q6
O7qhS+O8FQ3MUz8pHAPJVHHFJcTrgM2DS9WYMWq73HdhiiPU9S0LBdtXHH5wvYOc
czSkfMIHOlo2Sad0uhQOoJ7ZHcIaxV92m0UHZ8M3uVnn2SdrBcwHe68JtIthZaS4
D9LWaZhsqv1p1THgmZ446W3vRrG8XDJsgiupOOA2BllOgSbgXKYwOCWcyNyCP+oz
m4UdWV2xboZT4iYdJxC5ib+LmyoVeqyGFKsiKyWqunj2WBP+8x4qBbwmTlX8y8U/
feK5mHMjlXm6YgVZKCpaSP+P1Oz4J7FxuTzzcn+zXnKTg30dC8cFZ2QWMK/yC3L/
UWAZqrs8h4+Ij22me5sUkurH/riCHwuAj34TekPQQTqrJFLCfRXOfNjQqRkKXmCm
XR85VFGMBF9K55dLnHjrt0/SYtHcewIX4s9OnMC83Uc8ABcKOG6aJ0CtjkvG9JkY
fx9EhINDGAoBvTrRINLzgriRwHG3zaoIxQ//ahGXoZkeMd2GN1qJFKMrT+JxuuhU
PE/2TIcg+87jWNGQkHG6vyY76GnSGh7NBLUzPmyCN+12H0oijz1XYrL3U+U8mezC
ZqFNLUiIAowrrh/G9n1NZq4Akw8Tn4oPJ0Ifag7EnxHp+4GvGoNb7OpBv+g1WZLx
lnAbw7SVg3tJGlxcjhPiuCUltR8pShZD0xHVKoYJX/bpEC/BkQg7hoIXcMaiHMLd
KuCiPx+G39dFo50ct0akeN07p73QGnpfXiUkstdmiyhtjGgPK1DNV9loij0WeDlQ
4a8/iuH3gqaFbqABp7rVXYPFI315ohqeP23jXLyPUWmcP06OD1O1zPayBVr6H/n5
ecy+ORh3PP5qcpcHf4D7aYVwhUjvf9kks53fIbvRKAHgqB9z/iaRi1CKIJNs1cfZ
aF1vpBzjwZph1fvCz7Ra7kBTIqIo1iIBsTw3w/JeRrlM04o/CLH7J5Swm7pAwBF9
XZ0aXyQXYymhWyPAi5f5i7x9qb7o056g6ypP+DWUfA/HSC8l42qaLtuwaMK7PDgV
H0XkZ1sSlIUqLLsq+UJRCRPVL2sAn51fuX6gn4/IyEPEwp/mrvNubaUloeqrc6Tu
S9WLM4ZDBkUha+kArMBRgtx1FzGPr5iwqgDvnDaGz3jxgLbRPdA7N2cnBEHsAj86
V15ueMTqHu0+evwHFCPwaozNdelIxVwcGm4lLle/0o8rqJ1SjuCLswrXx2T6nNDH
qrqcugSBqyeEZ6TZ5rxPnkhJr13eMuK441IWtyLVbDPI0HYy3D6KyXTe+a/RDVwq
fhXEsV8PtFyt9rVUdXGksqh1FBIcJ9rFmTHoQm8QqhzXPwz1ejexzrkf964ak6MG
RZbU2KLMsbODfIrmrklrfxmlNS6/n2wcl00qNmj66yxWQ4t0iJJRP/5JRQ8MaTYB
nKa8hVwt9KRaQQw7PhMcVTVKTTUCGDqli0kXHg9VK+qOQoDAVXRFbE5uTmwpA7O2
RMxBVvmrqfMKdJsI3Yy82WF2Og+ZwFal3blNlmrBs41alBGXYNtuzmSVivtTuuti
CFED9Rg3ziq7X3ZePfFDJtah4iXmwvi7G8aSQJgLyQT9DmGDfxSNafFN8yWfTF8V
lckuKxPuILBH/Nv5iEhEOrzJlcSAK/NsutTVLH2yaQJ5bpla+XAYgGdm/GFZQv0M
3L9qIewfSOl6CMgvZb6F8wBT7AtpAxdqoXa+GZoJYcUGEe0IOPqY04t77ef0TXMz
p4HycnW2aatA4/zALQAnPeGUQXbebfIlaKxcKyFzlHcvK9U7pDglr3HcUg6U6kcx
j3xp45MzhMV4iNnOPKWzjQ7sK9FczF3A2VH4ShRnu/7UOKsJ37wfBE9f9W5z8sbD
/+iHq64sseJip6BfUaO6Zmn+bdMprfYVTPXe06XRhlcP7j8Qxqv82YspmJ2UEaQg
Oh3UKxqupxLyQvx8Hrk00yI1kN4GzC8eDQLxTPxANDxlQBE84h2Ia97LD/6ZKTQR
4/GXKjfls2Fm2wySlGQdseKgieCmb/FPMrhG+DHZIY87FvVcF1yZ1MsGu5Q8TwK4
ZzFEcFB2mrrH2hgcNzfrmBj/Vk9OSIqevbx4rPT8dHzBXaBP7gnVvhyZpv495cQ/
uDlMrNtWLqy3qFsPAw18Bw0gGa7JMABmVUtektnqYFt8XAIl2+25KCtnhICSFCEn
9XPW8lBCRJmk0+Vsev9QjjyUBPNJrl0CpsnTqiKC1I7GgsqTlbfyA21ZrRdDGoWz
syvuOqTc2eZPlcZbC64bFNsfGcFGciROb7LNKrB//6sKN+4rGjiXk5wlkXnb/eN9
r2oBmlTtCQrU0gQzB9f4mS4BmDOh0OAGjL78HnQrTK1ifbc1TBPQlqeEcaWWlheA
7MGGjqCRhGEfd9SHtVKLAVmp29QYBvBddoePr+lxZuf6LsYnXoeq+NEAmXCVwgV7
521Q2HwMlOhZg634GVWRPO4mzwmUKW2EKS+oXyqY8vPrrptrzoFxdmfXOw13P/th
EgO8fsY3h1Pnc1cQXhlneBa3KIXL0JrUryvamNOtnp414PbTHk2j17+Bi6U5UjCI
2rbI0O8MWtFA2lMJe9W7/M2Ebwd+a2sFAr/ASajo9X/XjT4VAQLMmLB7F+KWSoN2
/c4rz/QhyPchN0hyexA4BlIctIYjeHbPstF4izpKWRxacxC62N/WkrjcKgzSo2XB
jra1BczlcdzOa1bjCkquMmfEP3oDaBeh+j6+8LJzfDVuJ657V3XC5/hc5qT4r6Ff
0V3WjiD7rPHssFnd/dETGgek+K0glkeHRj/Llm9D0Pjl3EZjSKR0JO4LfXP+x+GD
SsAi3MBR9dQTXLglL81WQ304SdNYZ7JN94RiGNaoBhwllPGhZ6wuWxQKce/jMqRL
XW8mKInKMV8GCn+aaF2oZwcM9/SJoZG98Z6+vSEAIGr3uWiBgn2vNBMPdoD/9QI5
QxpZF2qi+BNGNttJRTSDdrpFon0/ewiEgyNKBK1rIDchWds5gTNT8ePYSVg++8Z2
+Ibln3bAYZ6bA/zSy5XGQzBYEX5QIscw5AmFohNsjFbjWKvdBudajvErYXvgjvXO
wQjuH5v+8V3SnyGO8seKYPDNwZwJIeuXeL8VURlR1bA3rIo3HbS8tRYuvjjk6Xce
C83IQvfnsER/IJbDM1cvU0UupX2QfTyLGGQkQpBqHEtw8eMlZNdpv3ucjlSopH6i
dSoMrnc7CggKZ+JQzqjNqRaX+Hgs6h8Hj9BCuJVDNgGKEwd6vBfxI2+gAN4Phh4R
NKANJLPH60drpM98jQ7kbdkH9mCpkYcMZ8Nt9gguyWaAyZSOFBsJmxwcRzdrttfF
QVRkQYXoEZ6KKZbZUpvPkJ2/1wXyBT2/5ZLhkd/vbQ+qCHukATnLOfTQck8oZZL7
FTUFRYDpeOcTqIcllHHEouUG/nSz6h997w4lQvrxrxj3SEwKwbwxA/qYGhVLK8gV
CazgSUWEhTAfp3uYtqdx1bZ4P2NI0fgiPMw+lFXEVZwy6JC3Zh1BKiu9noagmBUL
JD0cuNLZqLK+Y5wG6TrEK0PRBjkq0dP9y+eVaLBy2uBnihb+XUduXOBDJ7AdRs1f
syM/FZK+H2c12P7W793zxX/rzw9NlLQRK14Wy4oUP3fmjSWKkubt3jJhd/7TPUJu
19gTr+7sTQztNyBHvE6k0RZ55b2f6z+BrRH8HL/tEWpp8YcmsVc/ZOr07dW/JWOk
cxPDqxa3lbZMmA7S+Gd0uNJAfcpOGI54bEyI6i/o6ZkYiAq27FO7unXLNjc8/Ekn
pBGnLprYLsM+4rtvqLv60MkOPDrGH4+IzPVmjNMEoIKw6A39gTZO51WJMNT+cJep
dBHspz8NTc9x4vgSZ4Viab9Czj99YjBb6IUX9T/rurU5ippBXPU79hW+BafCfZJ5
zoCRLn9uidtqBzTKFBZmuStSxiayH/JLUTHaf0vPCpoh6cE3tY+uXBmXBvdjq0rX
Rp9HsMwTRqwmrU7Yj69fjeTrbjqThn/edVnhY/kBknz/Amv8JGblTORIKdU+7gAc
03VeT1z5GVD9z4X8cmWYVgCLLRHRNE8De2H+eQxhhXWqiq7kcMXgeZ4fCDCLg/nh
TJkLZoHtfk9jzMuilXAMA5J3gkUX3R6H47R7k6lwuQR2LcPDXmKLDkj2HBOuNLCU
RFfUgzUbYt82bzBiOOyBnuK20VvUJxLvOtsYPFiVG0px0xYERoUAb0BJdF32qsLY
mGRn89//RjpyheW69ZJmG8ew+eXc/mqHHZBNTlMRsGVazpzCdyQRZgZJv7eufYF3
wg+b1Lx+TZvV0Ds299qZlO2QD82k8bi74Sr1JFU18PlMzWVqgK1zoP9DwkY2GDAb
ljF7kbvUmOOiPaJvmCaN+fJJIITjRxLCZ4L9k7ej3OuYqdxsrmZZEMGsDK4ze7lj
7F4t9GMxQAakK6BMCYBs5SB1tJFNfQKgvsdJoQkEwN6w8emXRSREFb4PiuOslhEi
l0083v54n3JhVwqZHRwqh1dy0zpwm7AWvs6TzZsOGFO6T/6dTkOBdCeCGFWpuAug
f8UGCKV8oK9nGVmQFOTgA/wdNKhk474R8bCvaHCt2Y7rkrb1ou7worQN2HoOb4IC
a7xhp8r8+yz49UglAWlhtObpaNVu+u6HfO+RLlz9Lgl1XRFq7ggsTKYTlAn9yEVx
fytGlcCoMesdY47XErEobFJQra+Y6885ePdaY7mJkUaWj+lRyOcqupqIzWzrj51J
Z5Q2+NFw8/terE6/OMKj14kXCw8Eq5V+J52wtuM4F9xi9J2X9z7UW2Tvvf28SxgH
QFz78/FAy6p8PSvCLfbr66XNJ2HMs/7jJRdE96cwhtbuiwUh2o7ebdV9TC6wh89m
Z1og39ZkOnA4pwq13J9v81YV0zzVZS12NWVkK7oyb19Jbvx7GgnvcnMbvb3t0BA2
bJxUCSVe6OVKXN5skA+k7ilnxW07hdYxpi/av+oEAgShe5bhg/APeC+peMhemtxL
J+wlendT1lZ+WP+ac+N2KAsLS9kF1pgB7eYR1RkYqOdnRv7KE9yotbKf4spWXIw7
fSkA2oveFz+qerZZ8IBEaAUFxh2e+1EozhGCuRuJrgnCFi/MsoygyUc3a3gbCpDd
MNmaAiYztXsjxRpLRK6sUZh6Iq3RPNZYq0kmG3+qXbrJevJgsgVo/e/frAd57bqk
no2e0D+ji7AGgtwQ8PbXjYfrYX5NT/WHrdIuHcRdZposyjJNuOmin6/PTGLfC+6f
SBuQcrdJ/V1ol2EP2Agv7Y6+iZzXdxmpPtN+BOHPoW1/ecgGkks+l3uPYoh9cf9a
GhUGm9RmMYIDvmnVH7IiUQNgRSj0c1ls6FfxB/DAtttgrbegSRTW9Ucn/XSahk35
cs4njuDEeC9yqxalJcd8Z4hoInPCWBnaQGekb5HWF0dmPiWUOhBTqNkW97zeIhqf
G8+n+yle8FiHhGHzC63G90XHZePJXi2KTZ6GeS8PmFbq3nPoeNQGkY2CY/RNUsh0
CDCj/9VbaD3fTSZlukuNpHy3vKnJnxqDbgz64D/bIGne4aCn4Xy5zQ0enERZWiUB
SsgoCn+oXRZbhlKI78KCBkN5/j61Wf6MkKJCoJPY9OVOQfgqTtau+fidAZTlWXJT
UE5Odyejzb7K2wMh7prkg5kbfEDtN7gvc38oqU4VCI5XhDtStACggdv80Trkvjgv
G/oklvy0f2NFqPTgk97hIA9sVPI5pFr3BI4SqhKC9GEPgN11OMEJjrE3E66tjVF3
djGxVhS3a0J0U1X6Fsez1cmtxhOFE7oUcc4LL0KBWsHRt05SYN6juAt0P58L/voO
mZl6kZURljlvNsb40Nu7ABWVO6+ngj6ZcPin4BVFJnBV26ByVsk/BUEkQVO/WSU7
NrUaMH0yilLEuzmU+X/xG+elHHUPdlPZYOy3b17uC2HTWalgxSnGVUCrVGlO1UER
VHYFVqNbVf2jzjmSu2ycv8/7Q6C7sbbSBcdixX8acZy6E06oCzF5WMSlDMZhbxKX
VaTUB6s2FAidKKATAFnXZq8uT/DjLiHMrdjE/nUxdS4yy/bS7KW3XCa18jHk2nef
vdGEQcWIPi0FYYI4eKVuUTnbdAH6j2E8rENtSu5S7NaZIE1VeJ6MO0JxDKcGVCJL
/CflObO4MPJBrjZaQOGDgcoIA56JSeJm8eVfxeqyermsVnnPLzmE69C9oD625DrI
1U55sPGNzC56axg9SD2ixU0UOZ9gCX2lLduzbJhyoi6sPUruMLm3TqZlHGIVICxc
eJRE0rjZ+VhsnJqYaBZdBuSuCbqlfp50hpkEog0o/IOZ6qRDdTffDURpQQkEbqIb
XRaQ4PcW5JHkscODEoFuKbv6IFJIusE83hnGp07MQ9XYDQrX2tj/Y63oaJNZ3qEm
mi8QVuYzBA4HgWEs1gfTcBVCN/iH7/qX7wr6p7ccVlr25QpiWb3vTeDbIsGvPAAC
Ho6zadqUUtXTixeZMpYjatvgyhpeD2aGrEW6QQ5xgVAyMkKWtOCcqj5J8oW0/1/e
ILtd8988YuNxLix287cqVtKWctlhpX6oEKtPtWcwxm9wamxVAbYew9HJw8Yt9nG2
4EBi645W18aUpp2ZcxLh3ROMCbYJA/+lA35XRko5Wo8oYAtx2/0lc7sjZC9XJc2E
b0FCKZIWMrp2vWlDXFYzRVbp5dphwbetJ9om7l5pWchiIyDP78Kp/jhdVR1CnS/5
ejKCyXd5ABgMKXrxPP5qGgTtgWy/2OvllljFI5o4UbYdmydi6LKStyIJzt0YCu5V
n/KcrchgyJxA+x7lmTglaSvtXW6gP8C7IVlb46lIfQ4YfwUuVBw4YN1FlKL4+yF/
WKlMUhDB3hJgtMVP13tZJXK4XGgii1l96Aev1bAm0mbwFkT14czvtBwqueKLgiHA
LRbD5zzTDfKz5srzvs13QwH+YjN1muI+YwEpMC7AnTwM8sTHHVe3QQHHki6V/yLY
xQaBIhvg7JPcSm7jjgMde5QjcxNB8aOH7mgmakEXk8VXRw3+FxdY3dd/hWY1Ohhf
nYnQOIKdAYp50GNxcGbS+pSdamIHkMjCW7uKc8TakfWtZ544Q+ZFQnERd/UuXbPN
X8Q40CP6K2dAmucRWBYXNcsZsueI80LjH9yH3cpg+jImBtOSiWGva+eqbZRlbkI/
yMxZBE6lgw+unWDctCJQN5018dzd68y/UKZ/VNQ0F66MEL24lv2mSwf6B+fsOJZR
Z7OMkeCdyboJ+Mpdkb9h8MplLIfMI+cVd8Afaa39RU0I57lxoRqK/xxe2d/YVG+O
9ugjQPSa8kaKedwI6kSO0XkHuVQDPkexbWrWZ7w1Y1qEyP0luYB0r8XnLN0xwn/T
HV3i+slTAxpYQc8IlHQNaY3PvIkWkymZIt4YTkSH52JRmZiiqLcS6INrqhBrOxEB
ijLeGnJtuqG+nEYqJokwaXaE4mxc8cB7GAjSlFg+kwMKex+baNqQtf0mtqGLlmqM
EI7SRfisP9ddjUS3XyXbYsgJe711jCo65jRixQku6xfRzBHekg2G6362mg4pxW28
QYVwm89Wnwwp7pL7uCAHfD+z/f70FeBXupHVZYhG1VWgWNbTjBdMbEwLlEyNwRnF
86bwDyG/7iTeeggLZ+ylI4RtgXqT2ujJkAX4UoLAXDhXd8Bg+AKU5kBYQmd5XtPf
1dYJKV9c2Nge6YVZmARIdfyq1x3+98rUm22SJUaGac1OrVf5E2/E/G9QbPam6mvV
HHp/Si0Ya9NA1adUNgJ+uZSoU1DN3ONvDD63gl1Jhm3fVxMNUmcif9UVZR9KXxfn
wo6vtBpPrfJtQLoIS8Cg7SW0sCQ+HFUIgtvuHmfMLSQilTuZMBSDEv3MEAzgQGOj
kdKEWYeZlG9uPpjIYPJoPuhTWI8md0G5INx00PAwq4L1w4H+jOXr301qiPwS6qsU
7NOUi+CkzbVvzVKc+xnkKSFStx2s0cHdQAWZWBhsoLZa73ZOh88FWsGqJLie+QRT
S3cuf4nc+8SetYT5Hc7z+kE0CLfnyryBrBe6VcphH0zMehvlD6HMPFA/jbH/Rh9C
q61GtdxJ8Q2sa5bH6HuFbg+YVbXPWBd9ly4Z8GOs1VDj+6DF6hSCyLdnFPjTXxkp
ZhzjRj7dupIVtdfJ3kxnyr8xHTgmIsdZlOvJxz9GQWmWUWO0ixtpTYDTeN+qMTYT
StUKPJYqD2CXEns48Mq+lm8yB2T7jhiF3IcRi99Cl5zWl/LhdhOj5/CG3fsYM28T
YOh7WSmvBy5XR5XyLm6I1NA7QuwfKl/RO/wV0QYF9JKKkftgKvsjzOu7PU/fBnj8
jCPiWpPnlgk/3jkytjv8o5ySpBTiepiZSF0T6oKkQ7Xnk5677RdhmTeBnjLctdOK
KtBn5YG+EmxNh+gBneL/K6inTgoH+IRp9NhAHLIdNY+E2cr1Gy06+Sy7q6Ei1f/c
KbJTOVO+CSMFrk0QQMsrhmCWcF8z4Ca3qwl+ZefsISElFFimPhPfmrFSiGLj96hp
YlFnnnm6fvMiPbVHItdRfEXW7rNzaRKhedyosyX5lW9nWhKQp7Ylz8urwhDVV3Uo
J24vsn+baOrRj+xCFMHq2GDcZaZW/VOSRQuTv3pkg0ITdI0oP8JYDtwNSDBZ8SN+
4879P+KTEQ2tyxFU8f7+bhlJJ/ssTJ0JGN5LGMV2nCoD0boRaplTvcZtMd7xCAgL
N67p4KykQl0DossfFlKTRG3HMJ9c2ee02MXi1Vrw2HxTjxSdvL1nDuzIzfaUUwT4
YdC7rvq5BMCPnjHifDKa5ELqN0ESjkjATMe4KNa4oDGSyR9CUbB5urNcxzkJ7YcW
CDJpfKEpde8vCXyrLAzaUEZgQ9jJdoMYGy5xbOGvqtIaKrUtnPBx+V8TSkvf8RGX
s8CJGWufoivpMcwefraOwV7ETZzT88B7+mUs9ON8cZYpQ0QeS3ki6OyemNaqq59S
fV766tQ0sTtpAbWpwnww685CcphoF9hWnZ5kGXd6OBkwCZvJXGH9oRcM9lg7TKAH
UEyyY75qrSwRth4D1f2HIj+ikqX5rEebo9L/ExwhoYQ1B9RERMLkwCmcVMryEKWD
CiWhheS7i3wBWw78HEwURZg6o8SsxMU8iLO0PnSWgdFbE9mQy5dYP8HhUW7QVEDZ
cufiO5eSVtvnhEBYiQgIBO//f4DYns6VYQrI93fj3iPWIFYmrf0dRS2Iy+t9/9Wl
r3QE7zSSFEpsfPFCUUEyCtdbu2K0DahZCTI5Tkh48CntHryNn9IZxIP1H4LNwgIt
txOtKOhJ55xD1afyqYosvwgcgJ/uf8wQfWg9LyuLSE5XdKHJ7yOhB3BhNbGtH1Iu
YbGqiATEI4HaNNMGY1jkGzeW6KrQM17R1aOs8TneUNSb61oqDkgvKPokd6b92zl0
R441UZIkFu2Dtv5NPsWNxFAXb8vA2zLbYLt7in0dezKRjZ3S+DNUVHUHeDFdoi1r
TxBvxyzsMKze40Gu2GWNuuGWsT5CBVpr7LzJ72XhuQHKgd0HcIZkPabNwUnuJGyT
dnxPDMsrsCtzv7KBgn1l8e8EEyrT7gFmBacUOlXied0/H8cav9i6TqbyQwdMKuR3
2iPu7l++5wMsnchiRVlXzg+j9Pj7Ld+vX+wnIPf7L/mJrBiiSepjJcPQ5oHstXK5
HcZxvJ42c3+FJ6V+8OKwrYEkybE3l3Q9ML8dk333j67P9bO7//jMMJgAPuzHPEFx
bR5aCeRx7yJhtJfgn3qVnyRpw25GglWpwRI7zyFjO2Gu5xNLrOubvs7X7DerQM8A
l1l90ZLjhcBQ1LV0jljgKc/psI1aFZ6lC4PVPPRwsdv7y8QhI5JT6SfVU7gfh8XF
gY47UvabqJUT+JnqfhyGhsGYFeij1tQU7a4r9jrf9oKNMORugdTrYsZYWUTg2N/W
y15j7inMlUqgyr3II7GwCVqrBLS5hMkpOYcz0LPiQlkpjnwh7Yx0eT4B3N0VpL+L
CYBtwhcYQmYmlDjX7xCGfWGoKo6CrhNyeTs2bfQ6BfyTEno0Jez48fipFxr8ZX9m
C1TzdfNxAUtsABqmg7tY2x7PfTsU86z6fHdDHbR1XnDGk99ojuts/XWbXEcfXkEt
m6aQRLmW9LI+hc3OPxiRxTmUcipLGLD++BX1cw64RUv7sYoSWyLqkI6qY2gikhQL
c7lGsBP+HVkrl+Sp9fUBdYU0ZEMADAXrHGFM1UY+aH/+kZjvOANizidy8qPQlp4d
00C5DwSJ04/nqMMss+Pm1XeB/bZ0MIkkLIamx4TYFqRl3bi4TrA85QrjZIbw4FAb
49AWQncC4xaPt5JzsGDQUyKRWIDaQqeK4qYdMmayk2TiPDUjFvXIBl/invzWTk9o
13K7GyzXXje9X4XWkSbqWi5g5W6Bvdfh0Wv5KNmg1KE/UwGHzEqXsgFuNjFlAbtD
9LoaEyaqdcRkxEQRNgS5+/0UhQVMfbTDlE/H1D8bpH/sbOz2CHen07YV7wEtSQ9F
2NMjHLh1oYuNdCnD6A8MkhfaRmnheKe/1n+jm5tiEBfXQ69xIddxpxeAaiI2+aB6
YZ0oNZlXmyNWpRjKPyy6jNSk32xlDhGGnVxtHQlATD5dKXV4yM4nxB8Ige5NXXo8
CMGWsdZa1arOCHzjCSsdCU3G/oZxIO1yA1FswHsyfAOP8nsbDytJ9QQPUHxHEGQV
1oD9orKW3jw9qkSI29fKBoa/bPsn/OzjLYDynDttFYaShHyOwZj9xI3N06ucFcV1
rK2ERst94m7gRhvOBNuwjEa3buklxkuaYrPRbHtykg6l5932+UbnxU7RSvjOtbOb
QRHRQ2afpyamLt/547cFvuKYODgmWuEeLYIV2PouykZ3DTwRN47hdwmWzcbqdiPV
crkPLvvh7Fq9LTohyuWv4XggH2JuDBLvLr7N2HauHIm8nm5cZVNzXTRU5jOFZZmO
lkLa1cHh6LW9lxomE0sxQl+8Ti1v3sgxVDPK6dFXE/DmNaOv7fPnGkV/Ud7E7u79
krOUQ7Szj6PO7W6QCsLh+uoO3qJkZXFNsLyg9r4UMjJxQBdv3oGZiXE4KGEMikJS
Mw30c/ATNq+lietGrBw/BBEgVjd0wSzTRPFa+clqhCW25omEjKAze3Lu24o7xOhv
gk7NMsEDHR8lmTfcDJF2Zwi0sw7nLxF+ULCFyWK5ioTPToYWKeppgkEZbIA43+kg
4grJkeD2AjPar/rdmjp6p19h7cC2HB1rehwrY0/Wi+lTi9NmkJ5eEhcKjIAzxt3Q
sw7AfkP2yBob2xeiCsRg1cux1EgME5MfSk+RCx5ICnffZJaNDXG4JCN6lIhkyEtp
Aa9xPWPsKg1uzp86bEovDCnRJbCq9bnSOsIRceUDQ5prltR6OSYgQz68+LiqVPd8
lEtgO/duh+D9ZJ1wjlsH6/rb7HogzPOdqvYsA9gR/QrkGChHkdVPLVgfbC+8FtPm
yABfO5i8cmkxLtEmVaK44j5qZNVUPu6o8mcpXrybhJpBDMN1U836TguMdbiz1OB1
AUVLNHtfqfVevByHPL9YSpkUY8JfoJRzOL0FWw11zyFAY5xJwW7wdKPGWuwg01HM
/5LFCfzIs1aIumjgu7tLrXZwPP3fe/nI01aj/TQuRxIGpePy9OnTVY/B6uxw+Dyr
CsgXAjsO9i+IUoGfCEaoglVNLhGq/Bt8rtiqgzxu78WsBcr5VL1ZQuHgoUxh/uK3
qEsWjqeslmHuMGRhL5Mn12YaKm347CVU2cyLDNNDNllZhoA8Ljf3MP64akwi9y3R
S+JhpBXidp1aABOdqVsdf6ZesbLTmsaNNdVCBPm+G+9tQa35UkgOEfwgrJvp9tSU
9XZGmpiy5WFOZG8SVWHbKkHawHZiFL/qpIOsYvawRehgQBu7mPqSndgTCiX6kUxc
kBNUiBm0OgACXSlYgYYJpFP0twacVJ9ZcB5kYiyqWa/zHtWY6XHZgjBOvGrm8Gcu
GJEdeSdS/QdD324cSHncbhdZEbAS485w9GyZE+Z0BbwxEkvikXArGM8Uueskbw8X
lEGmzSBuL+dzoRh/YNxBwx8ZR86rdUVo1NafUVs5WOXKhkKkZq2DkIvYg+kUdlz+
f1wVZOYkdgV6bFU0cQilCtLttJPPBmFYXuzC+xR0UVTWHaz9qTW3zwvybVzTD8JV
fz1yA6KNl1RRWZaAAGYwrTyzkOeC0RWkbv363LXjXAKtSiViCiy09Yl9O7Qs2MBH
tRYtWvfqa1pjuJF3GYu7GtqT1CnCGSLNC+324T86qSJrv/ZvjGA8Q0H4AFOPKcvh
Q3tU6Qiu9PNNMV3GXELsPvMzRKONDjj+gPnfzeIZhIVxxRyk7xJAKFv6bzTCj2NH
IJ44ycXHLTjlAplQan8j14xvcTaI8tS04Wy5CUhmVzwK/ARPXeFUmYzSRCmmJeDS
cdH+w4ovYZXGn4DAWtMoKI9kqWGq1gq6Iu7Q/k5bE6yS7BYq72tyC7OR2+xwCCD9
KA3zoG2/X4bdd3OqHCwdmKQqpaNuhcK2vQsM6JWsvtnDDh8x/DcGAmv1MO2jaEqd
xxHEfaBTGj9MdWbrpumyZvoykTP8Z+PQtPRuFN6M57chBFwY5VuSLoUBjbaFSeVT
iLEzMAjrLjXKB3AZSZWKK+cKSQ+vNTPKzS+MBhkzE8Daat6m8+NCl9Rbg6UHbqN4
YmBn8TlK5otSGXF6TgNeQ6H8H52oEQfzx49yqqb688ISjhBfKNTKdRbXbmJ4Ea1j
zi0+ghCA8Lp6kSwVdTGNOSsdJUOaVCVrNgneqxVkiNT4vqYt2AiLquXQPyAIbrUb
FU24sdBQSgHCiRQRFxDGi9BXrxIhSXUUegAobsFdp/PEQcl+U8c/E9kFqhiGAxiC
4ugNmPHRsvV3PJ8m1sv53Pydj50YpzyDSaPLarHEd8blJybmBgRQqnV3vPVGW+J3
41lZEpY5pB5VQF9r/TuyO4kRG4OPPOUpBlIEhvrbKJv+UnGwcSVQn7VzbkEVUD53
02+bE0yTK7vIgi9Bjw1AxNpFriwooFLFS7+Aq5ybu+hoZM6baCfzwxWF+Ls1aqjp
SqTHCe6O6Cz8af/65C/nDDNaO4h2EfK2rT3gQzxwGQMLUw4qDwePRu16rzGmdGBo
/lbgHeALArTBNEvYnuTbTgeRtyluf0d6EdfWlVfEtukn7C/pxEurUbS2uiLLb56P
QzpdR4sl5l8qhoziVfWo/Q53bn1KugIUo88YJfCiROfyIS/JyzxGFK5RujuFKCF6
BoMx79mc2dnjh3DdVtjF8ZwvCe8nQXuKosb1Wr9CYJpFZYV8PVSsntXJndKBevn6
7g1BnySmX6x0sSiX+pOm3h81yjY4TQh0scAtj2x3BqAB0VZjlIh0UDPvZB2zU57z
fOHsmBvfOztzPe3ZQvp0tbZiz2YwvL7qkTEW2JDam3XrHqeuMlQiKGelcCE7ct/v
apPJymfNqYWo0uxwzB53pqEH2r7dgbEJOWz7EhdDKMhblNkN7ddKwkH8gYx0N7Bd
UATjE4vt/Vg4QFc+e7k9aaKmH0TP4vnoWC7UBY8PdjyuVrVqxABdx9mwXB52db4v
/1nxAgaP0U/YeTOjGQcgJ5EV+A9Rq03AaFQgazruKv0vdn9AIPbOjlHyipaiwq1w
8MmQPfezQanwWy+f98n4RFVaNmckhWV2L2vgwFWnTOqZ4200+tshYtM+Cqeh1RoA
UJcrR2QVkIgDNbMYGhXiCDcJa5EGVGGKZQv2QNEAilDIwNLAGS5xlXmoLHcqVZPC
2PK/EvZ8SfBvXw8LzEFV1KogVxeVCyP89d7OC7ZZav7kaiKT8ogZUrRWboBBhEj0
XGiNEftOADnEm83UU9OpTxFZXHE7mc7dkboL6ORa3n79rby5W+jb8xpj1+DsdBve
DiCQQDCNIGeI/u/smRxpObrJofNqSkFkolHxBECdYSwvP1g/BcRMEH75SkcGdAXx
gqLEgwyHSRfuPxBtEVjtMKrRDLUSP22aRdIywhIn0ZPG1vM38Zv7iDb4BoXQYizN
l+oOPZhOANhQNywJeVrj3kpye4FxrgbZzjK55iRUV6Otp9WyNoeI1Yh3uafwPDZb
iVX9h1GJt0+tqHr6zc1m01lWNV+m79WT9ViLDbRJ6ia0DC9UBF1NeQupOxwF0V6t
RnGlNeBGHWlvq59QJSHWF0y3x02zhnpUtr5Pi8w8eRssFjVvlMN+3xk7jUM9ZAaM
ZzrgiKWg65DtamTlO9MxKwTxR4S9eUmMCCJMjrjSO2ImIxcPsXKEdU929X1kFewz
nYB2NwhwOM03YV3vBJVMjvsbh/ljyQud3jD2LCsUByRTPKN66xZVWr+MAR2/5Bre
WIZ0joEuBzR2GZsyAms8HC26Ss1y+yOPTJ+1dC/wu2hCpcJXg8+A5fHyknR8PcZz
kwglBIsQfZc9K3ciYCG3c+UBINOcO1q4ajKihZa14wm/O88LgzPjWWGfDlT3Dl7e
D45aMBxKjsG+12uixuzujyEAFxWj5ENWWi6VcUpWz32pf/1Gd/tQVbyx6o7WqFl0
10+sXye7rDKaMjsyYQDzHBlNMDm6D3xZSQmPxtltbOnnCtEr3oktSN7MMI+Cf+ro
GPPrTOb2ahwLFaFP56HB53vZ7BzeHfSWxpXL8AlkeEZNk/QXKzdPqi5Kq0JTU8gb
/bZ4/EMeBt4B6Tz8yODR2kHZvnLCAWpbqNyNZoYC5rKcsBebUTEZCLQKP9F29Gjt
SxwqM5tHFL4YJDR5A7++NM+xDZ+Fy6Zf07yK0LjCTjTIHztNqJD9mubMNfElCAtp
Bm2awPlPFQFjX5ZXl2vMItgKaonhM+41W4NUQsz2dYR44AZIHCM8YSDQ5qCm36OI
e2XiQFCKEYH9Y5rGASIKz7nhu343kg5Xs6N4pzgJA0OPXyYvn/6Dp9yrKjbKZgIV
6X2RlPec+UWZPap8szFPoNAwTNgOsSH/dKcPOdczf9CfNTxv9MQbc6yPvUIA3gKm
xMhOdXFgpfpguUJc7bhVivA0Bug6QLZyVP1ypm4XviMKf//h/EvNBXOXwSEKC8/v
QBdwKQJs+M6Bt9E+aDgk6UZhcbKyyx0c5QOtYTyaINgv6r8t5RmlvWjQCfVpVMYA
/qVrD7cqqqP3btFA0qKnBMYYuaoKhn9dXikV5H4ByJm3z68o2JHa4wZC2oObEDl9
q6RSCS/BrHhHTlVIOvzlvXtjX6WM7kpmE31V/g4dOQkXcu17t0xEFA09YXnvWYRL
fRPVVRr81Z8m4923JLeNyAN6O6+QA4IRuAHbJ4rVigoBU74sS40O7AZgYr0WyUVN
3GikrYkFVAmKsFcGcdsx4v8B2rqKpeXkUQSWfWSvlTK34UDlNzX0bZQfxgBuIgKY
+OEVmnLGzftYmCnJaYNW09nLU3nP5try9mW8T8+mOh5+9uoy/JJm9F6TPBXBDoYa
r+a/Y+Hw6KqCC4UIUfDdfHOOcLoQnmgq/lptLQJah1gqVRGWA1aI93Mbpm3hki1t
pqaSvlZdrvMo5C2dztAwBHGVdEwJ/viHucf6JSCoucnFdLMSGl1Upymykj5hyGrM
U6QzF7FbyqAcSI8sFiWTdPD8iB9NCfJZ4WyZPXKFsk37pxPf8fAxF1bePiFoHrdI
cSLUY7F/eB+Fq64RXjc8WAusHkWNW75NyezcfeDx+ToQTqotIFHLi5k7ujyc8rz1
F8NVqXfdEYqzh9t4AoSCt29rTKZmTUz1Wr4pfypXMRT4/Tzahc+aXkemVwLYX8VV
FeQtM+xquNHGgRAkrs96MaYm864WLgusxXp7YOI7GspgYGtL/UURk3oIxP2A8vNi
out/7tfEcF3qYVG+Tm0SZVEQvTvkueWikLp+YuuBBna3YQaJTMuyXJWzoUn5i9e3
6woicN4Xnxj6SIcMi8Vj6gFbjw3ItL4cfQ/aHHQIjVXIPfBeD3Y5KoId5eN+HVk6
mIkCK+0B9CkUbJ2OwWFFFJfzUNiz/vOsAjSC70d1TXxoZjwk3AE0M/JLJTtlraWy
KF0nodzLt3rmZiMCv+9u7wxIi4xErq7X2nrDWatB0Kn1Z4zcbVeAzHQgKcA0uEi2
45aOSVrSewYHa1T121VW8hrjoF/UQImE9I5eYPsXC5zBTs0jzow5g8joxD87Kv/6
cOib9JggQNlI4zrTZPCUGyzZhcOFh8OF3hHBsvKBUjwXs+OFZRP9PT6ZB21uaQxJ
2j1ylrC/mhsyCcvQoGo51lzBsyo763sNITmnk3LHmATHtLl2ochnrh2US6qSor2c
+bExw5l+zqoZ6/0JietduCbH87jKGjzOXGsOLR1pdEkb5S4mw+GK1JfbDnT2IR5r
C+WLDCoka6uRUIqNgJbby3CNL3CN/kXYm//+PbZ1z7nGsgZuV0BC/NDKgDDct4PK
seR1TN0Oi5VExxDmFLO3eH1Fil0GcCPZkBVN35pHvV/bd99lF8hk/uF03Ie5OIzO
qeH26JNasoA0bMfX3wj3QGCsX2AEw88jcqVJzMjHuCexl1kMiV18ooBSGVlyy/B/
Th9y9hYFq7B+6FK7V8gGdfuri1YAQiHTIHRo2QlJ+rAJcPEbglwqaj5qdVwPNuVM
nQWhlM3b/BR4CWXeub+qPiPzWz/oKmHOp/oaPmRK0b6BstlnARI6/qUS9lChCoH7
h4D0/nKLGqG6YMwYj2qbX2pT6bGSQ33r7RlYod3uEZ2wsX8MWEm888rEVsorRZ74
bRN3iqD99Lj+bIiKGOsCZFc9OB0uZrUGZjBCfRWobZm9XK0WOQBcc6cZ7QbnQwjw
Tv8pMfTAQMLGTPRfWnZyW8/UYNa1iarOZvTzAoG1LK8p47aAiuVCg/xLzExt2E3q
/vgCcdbWnWvekDomlqD+GJOPybnZWX02WF4iXIBuukIdjV7OOkXz2DhkRl+r35NL
qJzzZTZ+29KQg2bTLV239g75ORiB3pX59iR2iGv4F2K6UGmqXc9/dBR7Kor1H75T
m75P8GqjtzTSFYEm3t+QK2lPwStoXyCYaUw6jfWoLnc2v9ieA64PI3JHadyqEWsg
FDfu0aunIEWVc9IuarLAD+e4THaa3H/6QHJgp+V4SsSJHl19InjqgHukhCeJsqfI
5HUFDCdjYrSK0Kv8LdKsWH6VUBB7+zf9xEdNQ7ol9+bk683c5kaUQPUcpH4Dnuvd
arCMvih0obogBfcRvRJ6ieFqAeSK4fs792/RQOis5lYsDrlEwSVg1OzeRrVCzpYT
EY6B/pBCYmb/87RWDV1YsSr6fhYOX3YWh7gwFeo5M/FfJOdSOuDmp6k41ew2Pw+P
6/mlHB+8l0PrL6kMGVhnGjH8tL16SSI1c18oVc9uqGcNMhxf1X/xkqkiL7NzENM9
yqLew45WDhwTpNhGYluKOJVZdY12CV3BVtM/Hm7AKVaUTfTmIOhMAoNIuDefOSR6
UeuD6rYblMdWc2xpPieyLAe0QUaRpJHuUASDDhUJtiHZaug4gt9G84kECzA4AKbr
671zdRx1kDAQjCa2tyd2/jzuGUw2rgOgWNI4KRxbyehj0Xkmwl+sV5xx0KQa6DOU
vp8JjlJvnfdpxj2jRwh9sKxLuqaeyOUx+D+lkRQf8Q+babrFvFZAydppWgfrGD26
wih83ebfZ9ZZHLtl68TvMkLqnDeZDd8FAQ0d904sphzEQdCoSmgqsQAwBOSCAJ+3
XZd69z+mF5bkzMi9KcLpaegyY42k+bZooZRpeXv3th56I7gZi8hMm2Hok6kwmqnf
dHb1fLd8Qd3P+gxFK8rjvuZ+5LS8Os4VlaSYyJeV1lG8uMrQepa/OF7TUIITM6lM
jf7GYewQ+XG4V9uWt5jPD2Ma15zcXxslU5rq/FNIb7dQ6Nh5kZNZL27L/Is/PO55
uC/vtIlVpPBmKTB07LorS03BKFNFRO4dRaQOhjWVhEF43st9wTYNZH8/FiBaZkzZ
n05x5cNj9PrW+xsinF/ZgbL1hvCwWk953/u48mTslHPPZdllnx7Ysiy78GSKLW4L
VCdLD1v1EqPGJakI2U2jqdoRMYtC5QKS9k35Ydl4iiFCPu6hmyTswa2ll9Wmn5Tf
ELtlv1Hh6zEeyHW1Xdiy//EN175KEeGAFLRf3SgboEhXobO3U0Sb34OtYZRM4ObW
q8FkYgNGeODiogOqDfr0nhXn/Zbp5hwyp3vP62Ov6VQ0OqWrL2X8kJaNFxef3lYO
i48KbJPhsPKQhZzRJxLi13E+jQ1o0nfdbsPZOOGEdM/6cYiLvSMrKA0yVJKKANxI
oDRym4vROUrkSj0gT4NMlZDqxuovshS+/pvYExw//TDImy2c9WcrjLxjVj1lWEac
QDZFVR10eZYSbVn1sbDAsN7IzfTBbXuk9ZUPNGoy0vrfBo2jqqZH3WrgrpmGEzfp
Jcew/+DkO1xU62V5WtuNCy23Uyl4/oXQOjGR/dCQCeR3ndN0uD7GbSldd9LYBWVn
dnh9orei+dLoQBQGd6Voh04FllTP8YaQ0FKd7OAWhQk7D8K88iBrKAm5YtG72Drf
EnkoxGO+WCeAgAktyMoMMcgNh9JMyUBrGwKowwRCHWvVAHTyZSGXum6lDaY8OpTG
qQTj6ZGRrBcsgyR6O7sNUkZQWL8D2qCKj9+9Y1VuggT+BctITfXNXXyBru9IcmIH
/QoPVtpaHbQrQNayCwCoAmBvZ/dSdeB6mBgpZd+qx0GVKYESnLMAomKBd/KgTnMO
S2o3fAw9OzmS5mqaeur91L9QFPwNU6YBlCtXUgHWWYUP+YWJwIKQ4h0XOdXps+nz
MDR+kKmC8h3Ws3e2lyE0fZOX2tT5Y1quVr/z/41SboDzhZIEsDFlij8LfyCrBQmB
jVp0yZBQ47j6e56E+CBVxuk/BiyJpCol2OZKH3kzIRozSz45VdQeB46K7s9ykISY
8LpPOcfqMVqp+AoW97Wt4w4F761yeVdIRnXV9BKVNjozu/P/VvwQITQZprQzXkj8
hpfISQiN3P2Bh2pI2snVp1g0H66ZCcM4QkOKewFM3hPCqAqNCe7faGDoewlB2dn8
sx1dMeB47Fnqv+qqsLwbiJUya0D/tcTmCzFywqloyx6EAc4vLZ+mqyamcGFS3xaf
/GHhS59/5KEXBfxY0mi8JuQnLbx5htWyHvwEdTTHo3vpDOn5C9E4gf26vDPNDRSh
6dQvr8c47u3sGdj4GDGDchAg8MguC6F1kFy0GnNbhUR+WPpTDZR6RySBFS+z6ilL
k//BwmKUwWIxfyUwuN1tfd3TktiMjnjO6vuJvS6bcSgJyrGPThdduELF9DJ3apMz
UiR13RjIxwYlcnr6yO3hFMVLCyohQVF0eHu/aaiHnH0uAuyxsb2Cm1x95ZNrDs1b
RvnUqsONsYWTFwR0GQCJMrD7yqOGm+AtamDTlhfAtJF6He91QLi73nXvOHKo5g06
03qidObF6XUOVe8h5BHwp4bCvwfJ7wipXRnFMNt19zCbXn7gdQvEnNg2pTOjEo0E
5Te3+tBVr9/2OAB9SQIvbLSVOWqpIyk52WjqguPP9LNqRb5Tnj+0NZifjSf2ratn
dcObp8EGJxLXcoxhz4raiBhZK31wGeKMhLqmWHiyYaP5uV/LW2pGmQ632zhkOM5c
kc+Pm3uAjhFl5OH4D3S1xVLQCloGlJ6DGMMcxmzErsFR/q5aShaRqWit0KSfRhEB
LZdIxn9oL0LpaF2PGlxgU4JzuLoEBux+MqLaDHWBnQPiBZjgPVF6eEqVBAtAkLMm
jRc+KH331sPQ3e+YMj5kP4Zv44P4IAi93DhFntYZbLIY8mHgHiUEHiixutrQh48q
l/wRrYNLUcVLKR/VgdQmC37m82hWYAx+PeYe60nEF4VqYiNayKMVy8cl1eEcM0VT
flahk0k86lnU4Jt7Ax49qCd/sW6BM8u/6SfW+HZGqZROirqyBaIJwJb6Cnh6QVfa
DvtsQcjKzNsx4Y7askYOcOudskBD91oLL+1jlu0FyofZlPyDjJN5/oBJ3pN1cBdz
HQXGyn2NVRLs0KtLnLVoDfe1U5YZf/udpplv9yvOTgFt+sBV7AYiOoGk8dhTIs3m
Abv9s2oiJ9Uwm8v/a/jkPLxlu6/zmJ7JWqnppS6WNPHUZZCeNqLa9AqPjUFNpndd
3oyHXOCt1B2DJqhj7lWmX/QM6vAbmRhaN0CZSUzr3np2Bf1ZbPzkMbtEXjrlr9dd
FMPQQ6i+ScD2hLcZ4BYiQbAuI5X5EAGPsHWVM3SZFBx06nTsT4kqNHToevokUtQR
HVs/h0zm/MKtEOYZuAvRvQ2wu4dCN8SN3O6q7kixi4Y1EYnK0ndFVAYTFdm/VwzZ
Fd0en0oyjM7OLzpEURaK6EXFnFk4ad2dVSunsHAhFo54EZnLfC866fL5Onjit+eP
MyiTwESw0zXetmykgomgvtT7tLuWmgcrtrKvvEv/MKOCu2thsGJdjvqp9ouutiZa
Is5ImpWx9wq17Gs0gqcuhK9cEtpretMEOd5AfXTj7yVLCUTZeiDIaRX1+yYFYl0C
ZFSb+PklHWKc/jZRifPaa0r3u70IJJOXgqDy/v2pdZ34MxRt9m6Ce2s8gyLPkf+j
wMy4M3JXt5tb2iPZLpEjsbgrWSqZtAXuc8Iuk3LS8dGHsMbynC1VQ/tCbycPvK8N
d6fHQqQoTLU5T1kMnj0q/TUnnNI0CYpw8D8bStPGtnYr2K+RC6GSq9Oozb9YIDuw
yL6v5iCP2YOP24LX1g9wim9CUkBSOCRE4sN29N7sMrSGytpwYY4+i5FwuVly71+I
rmj/pzUeAMlEcNhFQqSwSKhwM+jM2B+i/AfcXQGYagfsFqOiw7ZNJFpF90SACw/W
FjllGOL1cJdyH1bmqX/+dkf/PgrbyKVXXYZe+NZzJQCugeqDrL088z8oIF+Tc0lk
ttr7jVP91jW3LWco39+ne7RyZV06CCMPxTj92+CuL5H80xRKk0Fcq7meclnNsB/V
PknBDXYjQ8qDUk5VttR8H3mkLqDX+4URdypJCDnu4ep8qML1luEeSO6QbzIudxvl
za3r6+Qh3q5T2Q4KBNAlHcayPJV8WTzEB8P4/L1qH+rpzWs8NGQiOUvvHyMfjy9j
HWOpzEOvZzB6E9Wp8H6hufn5DxUFnk8PRFqI89gIH/sx6NpADDLUbSCpi5xR4AYm
revSlsOaTDnVjM+iLzHvkFQ8iwo2afXzZAJlq2A84UNjcudHvJFNWhYmvktOZUme
HANpHnxuLzGCkXJp69T81hSrXeMSHIqZRNCKEjLEkeDS+Mp2I4Oe2OkJfrG6nEty
Aw0kYanFv+dLl1hr+7hdqibMrQbtUysFgv9/gm1fOryHMjLjztopVKkI+IcZCTqg
TMAPDPZnqgOAMkRVwl/1cGpdOjk21dkoKGyaLjM7RLx2rPd8/1eALca15f39j6Nk
qDRt7pzhn0aAYViveJnSH2/4CLcs4HlH6iE13HxCj6eFlcUwwlFIfkr1MJznYolJ
uCI5B0pLSfEFvquByP012LUySIMdxSSU+cJMaGeVTq3U8pEhMt//5uCLiAS/AEsR
l1TKUjHklAPLO2TKmQXNZuFjVT+a4xylyrJzqkDezdXijhATs3zOON3MqO0sTbGa
stHXE8dsnYwikJofyIXKOkJv/B0XFRoC5dSVgXuEa2cSKuWWhiMssQ6xp9lJh5Bk
HukVTuI2kl5z2W2boc2lbL0wcc4wqhPXl1rxHYEz+VcDofrJiQ3dLAPjIgRkueca
EtY5KCEjHic+ZHPGOdHCdn7oPxiWDqbHp68zoKHd5e1LA3LnWBhOJLMCnKVPpyRq
MdPARFATTQEo3+MO4wSl6PO0Iyk4TkxDC2vXfsMGsRvnri0gRCmqFOuFGUbUyHZo
f3b85BpdJ2YjxtU71wKmj60VQXiXVGaFKdas6YUESJMXM1lxjaa3TRLmQxfxmjIu
IVg/n6U6d9C+3cvC1i7XQzHBVvxZoqFsIBguAZHw7/flmZERbbrcq6ptczmqRlfG
XX5hfYag7bbR6DHyO4uUmOsPXt3PZsm1G5imElN+pULasM/DrPsiamiR+upAmg+Z
ySll32N2V83S4NGjxySxi8na829XM2o2rTdgi0D+WhrvQFnqsk5H/6l+VICoezFa
JaQx3vm1EJKcs0rbDNF+Cd1/z5mf1Q+CYoaion8KiVk6UBNYoOfoDS7zmHt1Bz5v
AsYF85FwZSXsXUbc+g5dEQdL0Yq3kSZ6m2NkuXM6sxpb8k4VBr0nGgUmw1Zf7xsm
R1JNRw+bw39hoEhKCEZIu9HocUE8/A4sh4oZcrXuu33khhFmlLBovdyv0ihRR511
xfvSR9xAEK5Y7W6nJMb4vaiwsS0IKWvT5kcG4fBy8dkKXD5bJHCj3SsTXBtyuRic
lVARyOIiKXoawubLJhWBlSpw6PkzSOSesC0rJtKZZuUJ/4m78WHT/MQK5C7QgXHU
b9k1MEOy8O34jZOjLTvow93RFu3AeMEBXEGLVjyov3NAghV2uY7I2IbFdy/DYgC7
W1q9WpFWgbcf97Z0O2Xqzbu3bdWrYjGp5re/qcocl3oZIAtzXl3u1Vol0o6FN1B/
ugpxpkCJq74dWQfI35NDYmXx5rJ99TB/MqLAoAlsN3OdJ1QaMPA+xVgrKkfgMU3x
HYbtp9gzif3ehaySnAeRVxz9Ab3NGCR5Ve+gycd0iLb4JdNWKl+m5e7Zn18gLWOD
EHQofz1hsLeC9fN/93SGmLonDK1NiuiaLW6nsknLwAHEW9TkTcD+Zh9xYiBb6yNF
fi2xei2+rUuamH2bTSMbwnp5ixkbJTZJPrB90QPODUqVz2W2yYajPBpZj2vC5zab
queX/0PwKS72TJ50TLIWO3Q7hhn6TBL5OC+VdO/DdPcbIkF4gvm7vwGXlhwJYhm2
pcILjBOM6bGfC9csjqF0qun7Uf/kQ0Denyt2Ozt/ZL9KKMsho3/w8sisvEKBp/w6
UlChYH0ASqs7r7E+mSKACNU/snz20qy3rvN2Shs0pW7f0U+jFoCOcwY9vyybclbT
WKtfVCqgm7ZpiyheKvmxbkkT9OV70N3a04MU5d/p5qXdQgP5XpX493xU7tSJQI0R
iL08WhSoitz9P3h6DoB1BZTawC34+YuBgThg6qEIqYQHzhj290Gsru7PwR3dMCyH
jtidr6SLDnzpIXDPC4TqULjUVtcwTz3mCvOkRP02L+YA0M13ozPfs57tumq3Whrs
A7quhWNsOUfbmkrqdOD/gszWWBaPasM40GdgRVQ2JJu8vDiQRs2g80YTE+X1Do2p
3eJXeOi4NPNeB9Iyl6+WzwwI8aj4+TYZ7i/U7RUzXiEhvWXVX8TtdlTowTjv8lZ+
QGzvqKYV0Q6rUxVjToyeESIymwZu8kCMijJXtzzRO13T5STgY6W9NFRnH2ppPNVl
UVncxWZ4KWnXYvUEIvJvi8MCr6etfMYzHKuWVRkbSUbln8DPEsSUyyyMFZpPV7nb
zHTPcwRJcRDL81it4If0+iaHmKVl2Ftxm7pwzxmObvSgEoyaIJHBlCTmt5vhh7z1
L0OIjfWdS/Zu3cJiG7rsiP3S8h+a+RzM+pRFWUtZuOsPfKlvrA2iB8vnIV7WD5UH
TSUoBF1Nau4+gaR1o6ONShdQQJ4ujr14M7jLPoBgsh1RbQglalLNloEgJ3pzkoVW
hLJYWo11b7nh21jSQaExJQdnQNZ35JAYA/cgeHuuFZd8CuohVHdnVeu5Eyf0hJhF
bfvjszbK45SPDDQtMtpXvg0NxQHpYIcBblbJsXzjHaSXBfYfEQIp08GXJhNEsJx+
PRr47o86XmbJv0qraA7i3bEGayiv4+d1lRf7WA2A3ScWE9P1gfHY3HPgqEBvKWNK
6UmSVl8YfvdcoQ98YT9Wl/PFGZNinrpUgMk7KOIab9oCwcpfMCabqWtQY3ZqiaZJ
P1l7in/I2ruCMmvOUgdxlTTA+cYSdthf+TITsNTI3fOI3GTt7/YZ1IGMmKiMwuSl
nSK5EikvsWU2FQElJcN6xsxfp8GvXfB3mgpGZp603c8Ka3UvdR/AkVccG71Uym4b
4VOLSq6gFfX7LKNh1ssZUjf0ivVq1r2uJgFhpVWLY8DSp5ALon3RWIOer49fzxyE
oaXW25K6ZKXlThagWaGTUMEMskwucQPBoMh1OetAs/ubPbYUDZQ+Y7AXhISEdD4U
GZjKji6lEanj0d0zvE5kcK3WTwwZx6b/v4VLZz2lOtQC9gXYGslyODof9nivfw8Y
9ywywFAbCxfFwECobvG4lYI2OLpb4NpRnTvE37HPX+kSPUPQ1CW5qydhNn5PEBGa
Mb9CuMNTpwZ/A0KCfuu5rjWeFlSpOrerI7TIlmrjSE5N6tbf3xhvT8JBhdnggh/w
lxN/mcc30H3xmCrmJ4w3V/DOWHIWXEFKe4imaKXzCIL0tTzk4JpfsM8kQi2yhdlS
RNRFk2XZF0NWIjS8w4RPlWPwiK/SKXx2zhDwADSjy6OK64zY/vSOyv7a1/funIFX
xr7iT9Uid0SbLMCbBpX/XtnOtQ/EtarCuP1eUIWHJizIb/GLff0WY5cUYIUN7GFD
96vF5JdiSCvQuh9V8qf/5o30miOvwroRVNBDrvWiBkFs+5Xuthh+TQga9cKigW3M
sywJwhriXmhez50HUexrG1kpU1KjYDIB+kANlfhYj9nj2fWZpo57qpPOiYLtlOEI
/Y9VRpScDncH1VeNk1B1AZp3xV3BQ7daitw+NDGJuvBXGU6+YwcWRWybEeQ33qJa
/alcUHs69niul8vTi1xVx66xagyEofDkr3FZAXkUYx9ULML9FZid+SrG/9U2d4bb
rZUlNfKAgGy5+5wR4H6ss0mcKkYHtocE4lszwWQDuLRYXmxTuG8sllyF/xwsOemi
6VnbZsnejYWt0oIuVMH/jnMHlrVZiX0BjqX1imVS2tE+zLd67/C/v0whqvc+VGSg
DgW6GDOHCLETtRLS6oiLz6NHJYRArH6XBbhjlK+w3dAzvhV9hKDcA56djpQfjCFy
RgcWq0ts2oIOgJUKYB1/INmvXT9BR2eyEg3IJKFF7P2AnNVi/a+0xQWLBM9ylnIT
LMf647pzP9c4LfTkFBH/Cj2pag5mAZSWx04HFeFDVkY7PlHCiNUm+9MCW5dD4XE9
U2Q2xAf5ePHZRP2OfWWanlU5mpWMVbRc+Ahj8lQpA6apTfi60nGPWxWlkMgSl12E
qPUldrgZOXB1q+WlJaYDH8gMXXKGV5T0I6VhAAqtPXjP9flkh7LlyaAlwcGsduuJ
xEPeWR+gKmd+kY81tPRJ21R6yrYuwHysFEHKpO6tfN3AJpZa09ogyORPp5t7sAvb
LRMrv6K415V9lb6qp57DWyrlThjbnSkC9CvagrcFaExW+5+lRvGbQKDS2+q6SBKN
AR4guzMzSaflZ9z7zHLzG9u+ZYbQZarKWAthslAQ0kJePagfCYDRNejKT2HARuTM
nB7/CzqOmekHVj6hX5qAMPgV/8TkHxMNmsoOULioT8v6PWMMmgRcBYSAvA00a6fS
kVrmjjYHUsHaJ/y4Fw2UzScddrZvRCQOHTWtu3NzeKy7dvRjEgFxP1AeXSwO7LPJ
3J9f/fHSbS8gYIdTLL381jtrbIJLeeQ5BU67O5vrDxxNE8TnwNRLugIr0sWjGFyT
QvbK05arNiSFAOPOUUMGLMs1NVlOFWMoMyCg3TJ1ZMp1FAVSk/UwgbgY1Ri2LqQv
lfItmdjtiT2bCIuDDwe+ncwl9O6nVJa1ASjv+Y7jHUyTdic4WeH2D5ZoFB6fPBBz
XAyug3HgYnkRFyjt5w1lvqNVEKaBY7tQ4fj3B/JBEU+G2+dWZaA9bQKbKWKLY6Mz
7oHF8PR5lWkacXMbGRY2Y9YG7EohYOQiyYALyQxkSjUXDimI4Bl/Gx4Y1PKKrkpa
PdZcnncTD7VzVftvpuEI2Aw+AmKsHtqd2ygihQuMeLlPcOkZjpv7rD99xXEr3AJx
iv7GzAmHttDDYUpyy5mEcZj3/kBcVfZVk6ka9CCQbATpxQ1B4icE7cdFPFBaLrzV
LC69fIbLf9sKUIjUO+hkdVdlvlMkpuzp/sr/lGFStX/abFKKbQ+iF5p49X8rPjY6
rN2CJ2DAVXqPheesWq87TzJwxxOX9d1wiisq15yA5GumI7DqiB7YcWbVXM1Klp89
okl0OvLPpqM2mJuv/anypRuriEX0x+aiLCNvdG88w9jf/vB86NtM1n6b7VboUKyA
kRup1CZO1680mzTRX5xSQdm4+/J/d3C6lwJrh8jnwy0Xg/ZFNgKKhZc/9AlxIZou
LEk0GQfweWFmiaZUfoQul3R/GIU9m/xS7TzeV4w5qd/OKPERYkbPm1plZEoPn26T
KF0pCTOdJDknnOmp6U87XJvmk0Q+XpNPhIlRyUo9WRz7LUVuj9Wp4CjMi5Pd+zky
zGwvigf35LBorJbbOTL0xFPZnlY5xPlU9BsAcpSvqScVxlqAfcKRggn1RXUe3Xu5
ZkOsk/Esnmv6JhCxXVgVMMDIKAvRy7uOjHhLjhsT+EdHeY95tSFTWwCFsHn/7Ua0
jMRqeAP+aKyP00ETnA/J4gGFMyKeho0Pd247t28Q6hWxqVpmAXrRU1nRz6M9EEMd
xnnf5esbVAcpH8T3YmtbxMkQ7pNFAWMiduyCmJcrLry3WPX854Gw8Ri44AbCJljZ
n6pnNV043Z4/UaSauDqphsWGpbl9pvpX1saA3cT2/SJpsTHQtz8PrEPps+nr7/bN
Gmr3/fo+vU9pJ0FaEfxQXsQh8plfTt456hEuyjlNhJn9ZsKOZnv/XEBF/moZRf+F
HTUhZVYgHjOGZWcputgGl4zMsZWGk6Et0E77WzcLtfrmKdaTedoAVTJonoR4hIOg
s+lf/i392nAu6W8gbe+IbgfVoXFWwC14aou6chHaOG9MpzKnPUu335sbvrG38ThG
K5Y4+BsMiCetXJjHWdpLMnrV3WBQsjdS5ZTLY38E1hJQNDkrlYjfxra5PdFAl+bT
mLYoxeRX2Dj2EbWRWmDdjlbkKsjiD46Tm4m7aTOnlpflwAPCMmaV6d0p99Rd8V53
PH6LB2UgZWHMCXSc0p1Za9M8ZSCc6INzx3r7w/6hljZXGzuQlr2Ol6LZBPauNs6e
fbOPby3Ukd7IYtgJ58L9eScfyN8uZFbomB2YF+cSg9hcJsAb3ZKwpy8zVhNqzfa5
r8yJ4TOqJee2y9EYohy7l9fYPkKVWcTwCG8fRqW8xDbLDySnbQ6ojDqgp2/OND5+
9MZv0mnnKMYZAneHlEw02YjJXtupaeVjn/MOxsokXnCiIvkZIQO5wVQYr45aqD0t
//2GcgmuujAtF1cIBopfUY+8xqeQG8dKelR1ZGfrhrSmaD+CeVCvJBumyX3MrHp/
Le0wDsvvW81n+ET71Ndd7Mlm9NwgFbAo5vyzEdO03PQio5rJSuC6ueAEjZFL10Qz
oYanix+SaUb2x82wz7MPKAUQEUb6ABVnNAy6xVs9c/NklNBeeEooTotc+AMUowGI
zqjBhyAmsblkunhpk6nmbS4sDPWAWVYS4ECekob09sYrlk52Nikbu5ulM246kCXH
Tipd7ZDiipQJyDEE67jGNwm1G1WLhbSKuJG2j0qB7vdwAe/azW+U9WcphkGFO2Yv
9AaIQ7sJkcegD1nz22EpeBxgakDrwNyeV3wdUQCQWShasDuvYZydKtkuQw19kTMy
vAqkjtYvtdzO+Ityv9iGle8ERhrePezPvb0EXtfpjK0tZlShFRqNkYmMHRpaX5Y3
F1KSI+PeHvqHxq02o5DjpEAco3gwY+LPsP5d+MG+UMvBAupNLdWcJ0KSVBVYXOpA
vPsqqvjRmp5E4qi+/6i91xV0p6EqYWGSrtv69P/WyVH/rootSAUteipFNVQOx/C9
QSqxso1d7m6vMHR1IzkNW4Ft0dfr24Q0xB+h4q4glNfBEej+HYP56sih8fK4+4kc
qAp13fQmgO2vIad8PuDiiWHSQiROS+DCZtd9Ok5l7QldRBsHZnCzXM/2GQxbZQnt
93r8x7ZtBQsAyD6f9Xk15qYumyW7pr5wRi2U/O5qybdThe0B0GrRu0P8Is4FLReB
9WBvcQKUUhf00lfaCIp/zVSSARjnh8hsGTf61w2zJ/caR0RluAkhZnrWCidN0Y4a
TQRaLMV9H9SXdas9pLk4JUGPQCfFDoVUv8ZofHnfKouvUoAkqUfueDpEJDTLE6Pm
3DBVA/Qpm16h/RVSlhOq9jTxo8orx/OyF6is/xzqoRJMjAtTxWpklW/7NP69tgi6
iChhPMxp7iH48BsOnXpyQBeNSKwDoxTOD0NLCGY4AC/466YddpWb+ja/t4btNkfw
e4kBWbkwZ2BndRRj0DT9yg5wx3ohdgWjhXGSqlOpKLOF/R/Pn3GJ+60BhjQhYhvW
R7Hxtwo43G7nPqa9uNNtagEKwI5n9UcLTDE7pcLc1hw54MZ51JhSmR29PDpSjw6f
kyzPOupspCkPZc6aJ17jXlw9926K+VfUf45qS92smqysFf/X0kru+M3kfmJ441ho
/oBfKmzEuXSGmI3BGumeswUVp/UNSObUbnFcaaBZUzvKQ6GmkeT6oPfl7E9mzMm9
80C9HL7vLnV29BUCzDO8SvfBN/NAMgidLg99fhzzBgYkYYaCGrRKxI1jrWTyk9Z+
fZzS9I/hH95lT9bRHCD0yuWle0wFdZW99hV540Uz/3dj6I/+wZhLV085PnQbxchr
eV3YMS2EWLx20WAJ6BZm36VBQOi7QnjkHkWb+l5j8NrPc17U/cHcfHoqnJ9fTKd+
jIQvQ1mnbksIoXsoOMNfqKdB/cxMJq4B47aixya7g6IrU14WrHDEyxuwgrhUWS40
c9SXjEvNbTrFkNu8b4nEbhZruqkJyObWTeVXAaP1YMKOoM4CgouD24QBWj3jbKch
CNGmIiN4dLa0B7s3lgmnpeJRFQve2Kw80ku9khL+QUpIfO89sfv77/ySK3+oyq0T
5T8xH1v5a5TIA9mcPVvgVi/UjiiV9Y95muTvuEkch3YWQGS70ZRBneVdLOsctLlO
ll0QFGhPC83LXAts7AQw79L+KYOvE+zryQ8d5esizTpzBE8piQrbgBNnyIUYKP30
lyjD3mDHN7Tp5d/e0yE0YCseQPn+xFO5tW4Jv9Snda6DWnul9vMj6rgXA+ZfdjCH
Z10s3RMrkhFrB/AQz4jdMAiyaD6hYNycyDbgSS3yo2TXPpOismfQpEmq6Hh5N2Lz
RP/2mfkgbRWXkLB4PK2s6H15sUeWba+CmLA+n3caTffRp44a7oQJU5kpUDhW5zqS
If2EsuhTu278w1x2gAyUZgtpD0N3Caakcnt5dCL1X1CfY2loqkVbTnw6l0tTNyKH
GopkCrKqlP65gf2LtWc9OCHQnJN6NAaL+Ph9iFXdpIk6RWxgbqSQkkFkOMAFeEib
4Ol7xalgwXFJKjm3BqvWd5EpcHzkljVN8nucGMSVr82//f+L7kISRqGTtWmAXrRN
Zp11v574vakIL/QOF8VrTOlRCsqChh+XU4cxSikC37QMUrcAUJOUjPz+sxWAMDZ8
oR/D1VgKbdJX1Y4fcw3IH6QvaxCm4v8NdzY4Zj0sbZmXrA0RrPmQfW5VNI0c5MY7
+aldbPQl8S/t++XZlSMKxngL2zH4/stT7btmAUBUdOhPZDVYJ2+4xDJoKpgfNcSI
CjR22omMXfb8OM7NjVosZw1mqserwJhZEAauZJPpF+7W9bIDJR657qW7KlUx0y/y
Dofh4xuE7oi0ZVFOFFfVS3xHlkAUafHZzE4jzeSVFYGvrjgO0z9a2t18of5n8FAk
HR9bUktaXRHoOWunYXzb1BogrbIQN4s5pnvUDadtncPeWPa+GwUQNtVyONND4Pdo
1j9EG2RkyGPsPlkUUOZnZqnpQRrdbSWXjIVUlVUPEC75i0t7+XtBdWV7RqoqCg3s
kOdBEzrNWrrzJlUtMdx3hwo3kmSpivxGPB8ZbkbJGhm62xWRt8e0VZxQOeOnibr9
dddSPwshKuCS+RepG7n9mEr8qI5r5EjuWuzPnshs78/DHQLb++I3oyWKNib6mCBk
H0TxYEbFUgfXtt16BtdyZWB4PBKMcRdajW6Mx3qll5AWqNXQDNoenGOBoAmbtvA9
YJgtbCdZ4/vRu+3n1TBB4WBziT4s22kFgKEAY6+ZSsyB6FG2V4GrQGiqvdv0ver1
hZUMMATuFZTnpmeX7eixwTHK/m251Pm9t/SmK0EC0KDSXYoMTGiSa73wsQtCXRnO
JWoqI9iNWOCaho9S4GoIo/+wc/JSJoxxO9hNRyBTNX8jC1L4UomtaXLcY+M0fFF7
+VMPydH2PvfloOHPnlR0KWGWUr/ApvZTdc1GiOc5OaBnLA4gsR9YrLcNRhcX0uTJ
699Fvj15rHWIqPeS4Fa8k1y0CGICLD36kSv0xFHPZCmyDiy5USDne+BMcnU7dd60
HG7Hz1bPZRzMMvOt0BLIdqXxlVhDRnWcl/ajsJe2M6ZnJZr5QFNjcFc1WB72Xp4k
JpkxVePRDBBTsvCsfa7NKq4SU4G2PYSmQMlVuphvnuXQvyRX1pUinp/jN4D/Pi2g
Z8CMePO2rA1oDHgoxqzLK9+n6bFe6qaJ2yy2MQp0uwEw0pWZCG5fI3OgIThJK/uO
YTm5J1ZqmZQi9RbUn/E3rtyDTFMENaXbyJrUgSMj0lZ4LRpdOqcoDuVL3b7BQkOu
BWxQjDyRF5OmLtXKnJYd2aGpFqduxCZoWnNKKXi4088R6D1ml7k30z76ndnaj+S+
eJn/u0H5DMZyhs0EQDX1A7EV4Uv2LP2POH8mAu3mMZC3ch6sdQDtv6CbjEIrJrPy
XAwKm//UvMyUn2S/wXqFanXWskQalUQY0tZHdgfnakRLyHYOIaB+J0kUa3PAS7ol
LzR5QgiUrcF1d9s2jE1s8DltL0JNlo4RD/SkxHXulWcW2WdeJCaD24OguvJcCaZ9
uEZ0dNkhhgpYYEHtGg42rWnZdaFv1FCGT4WTjAye1iYPLkn4Joaf4j86XIKt3dWn
j7KonvQvDxLE+RVRUsEYE1wPJ438Z2+gEKGVZyHd76UmihpMbCxhCCJ8VwtfD9Md
kdKsPq/4SefCo4QW3YE7atXqrrOt+vZpFqE2luDkAPa7QqrseDikTfUpwiEM0vwR
ulJrDROoctUcIqjspjeDqzrU+O1RD+9cqZzBdaqz1jtC/2Y7QKF/Ai9NI5iQV4qD
2zo/HeU/utekVUWAiJj0U4bUSOQ71Xjnz8/W5heqjo4yJAXfxpI2HbO7Kcu7Bz1Y
/oVe62aMDv54C5qLkIu0J3JoAyH/xp8un13EHYXLKWsL86wYsO5QIYiEjgPIR2W9
LA/U8+0GXiKA+T1eakJM4B7ij8rbjFeNZiKbtQ8NF1Wppkw3OYU9mIosC2fz1ISU
lQr6AcAjSYAuCtnZ+672nz3ldJS4vHThGb5mZ1G3KS6tOs5LQFVv7GEQbUTLW7ib
PJYOw8t51cltsJmJD/Mra3iPX6kkGW8/uIwAMrOvrtBB7PGQXgXUsad4UcdPUfxr
YBKzkHywyErjXIRWavZXmgUoak++SOoFvv8ZeF1b6OhEZOGJ5ifeWqhb/4AGW3vH
ts1QFEpXqIwQFb83nvryM3Jhmwo5rw1ZmtkUDKQpddRjOZjEY9YTj4TS833NoBd/
QtMqCghXG3jetGY4GlSInVv6Seun0JgUKP9w+bkM+efXYGrQHBu62gpeLnzqbUKm
qU1YeDCQEjTYeUk8V4RUYYaybB7tPz70GNcd9pkFA8yQPgmZQ1LwkzPHN1Ah0Sa0
CO7LcC+3/lWs3xKlC8KRGj9W0dowkYZbMRzR0mfuxSN9SSA5ycd/eTqKiJfbZ6Yn
3wPiBAcb96s+Eemdjej/wcIV34WPi5czjMCje+KkqiPUg89j6/QjvpUIwYg+aYB9
VxuHBu8Ngd1/zuHnIp79uSZ89Wi+Woz1f9QeW/QrixpgVjziBlnHXXmqQkmTIcMX
yQzHCg8xh3NzJVVsyleRk6noZI7ImQf9frYSCurzBxLQL/Fs7y8mLItA9tizSsL4
qT+/fOLMROUCB8vnYbvn2ww4UMZwJXnTIICvJFazVwi/Wo6xaTg2LSS/E/utkyK/
ndCh9WubdUyCgaYdh4l/vfECpGj7ir9XMXor3+Rjl/c6J24/lMRYgEApupBfPOiT
uFelpXPGlaoN2eWcoAOdwD2OUxjbx5UiENUh4rg9HPBNQ/yexixhrA/9sllYvBt1
6xli4e6dEbZ9ALFd9G15noOLiJ4bm+DzMeXnpUm4Ol1ujqqijqH4pmHH9LPwRx0s
fbUZV5flpEAGxiyLJlKlUpnfzHyCYglAp8vx7tri70dtEpOm4PkVw27wxYqzRrHn
wPSa2heEQXVJrHLYFXMYvSjkD6uGM2D0+CodtVgTsaVV9Hp2v1I0Z9aNkWqioFZ6
LAEjVfWwhRC1tCQ7n/VYKevpE+2JYOGzpeq+Ge1HYC9uHbbYLWGOhAr+kNoZ4UfS
kn4T4p+rBD1syAA9TL+RX4oWaTRbRV0sgM+W0zL1MMmX1HyI8Qh/dq9DDid+57yu
LU6CJcRQCtxb3HCLLvvhQE5PiRl67HJxGOAwlv63iVC3Xc2PcIRdz5TeebguBvdn
Nqi96y+eroD3RR68K9aTMPp5f/gDXgHB/fVzsyrT1d/IPWgW6ew6e4+mMgY3AB2+
By4MHA/UnDDxT8dVAdMjARVqs/OK6Dm9c5zP7VsDUwNi4qdonQ0nylf3IEAuG1n+
yHP+P5ajjjuMBZ0jn4ZanoUQswsD3uYuWaHBN/AeqQzU36xuGVxUvTKmEzdYsYlP
g7P268r8o8kf1yeRVVXDyjHkFQ9vC4VW8BgNWfq0b9iyKQJCRkIloj7LNkUQrdLZ
rsaG+gImtw6yiuFh6UVi/Qxdig0eAFiL4Tq+qExKpD0uffvBbX9jvPP+pjHSSn6l
gKofZMwCsGotlF9tdQbxb17ZNU7wjr+DDrS9FyXXajQ0Z/MlxZTfr/sggWnnEMXh
wLFjmzmaG01hP2OMA5WBaU/i90JAlPmoDAHqAiyylsGwKJySryS6eP08msvSzKiF
6+bHJvG3RpAQNIfRIK6mNxpOrfEoADiTJFh18mEUfm7FiiDwyyiqQVY9a7yarkRH
h84Rx1rUEV27k8Q3aYbZCvrYAMBbq3F6QHePiZ1PTimt8RkQX9V+fn6m4XFPa0J2
JKSlNEXOdwJ278QN+rFg48WvrGNIbvC6NRaSYGVa4ezJJiNedtHxOZuNqS/Kck2m
Fo+XfwHlL96Kv8WIU++VhCWXrqimQrlX/i0iJYujyS+izkiWcJk6w8y/saiti9GO
NWo54Cv847XLSb6OQkWD7m5CaofytQjlW+JjaY4D11sk+nIeZ34lsmb2P5R2dHSK
AlAfMy55RyDrgKKVg18S9G7LldU0VIMSpYMQUtVEo6Tq8rSLPa1JMVmVBM+gzC+f
QqfzmiN0LVuI2wMajRUJht3k7g+ZxCRBr7QrcLBmby303Fdg2SdwkxoDoxN8nMAL
FTZYErQ+RvK5nhLq1+InPpAd+sGLwucPwX1mWOyUFBQgWHtmZ900WrI4RjOTw3wF
6WzdjlaLQqDvirVad9z5BaVg4PXJHrgg9YOJFbCzu2nahHv2EJ3QEEJG+qX4hQ/a
ukV7TSTnpFiEPDzsLk532o6cO3IPb2AXCqbQXGf+yeB0Efb5XrQkv8jQ3dS3Cd7m
GIskwHAbpkewBa1wn+UDvQpl/4cWsPbeQxyavU8DF68cdPVxH7rTooX7QgwFCqf6
QB42k5OIWdSbrxycQFvwOtPvKg0IjgCf/EUmSt4ka9rjIhtPi1ACsncyS9zEw2YU
zWMJnJvPu7l7+Q65IxC2Mx09OiDWCBT04tWgCEneGb2QAlMX3fGCRjAxWQL2beHd
Wg1O8nXHN9RLlRut+IsJ0LU0HKdcMghGKgxitzIP940UMyf1JD1AfYUHTZDv3BtY
3bC7VPtAHM954y5zbzzD5OzVzjAn+xPkK6zZvJEacD2c8WXM5PmYXts9Yao5tiAm
zJWWGMa9qu8cftN69VvEyJ5qKHHqK/oyXXLV0SFVpvrNTbswk+5sZZGD4YSHv0nt
mROgzGquuqYrBuuXKFSgyz5OQTqaPH8c7276WJmoLanTTRj5ObjB75WerPCT0+Js
ZnAxWU8BCEqFFUzWkXKzBWvfMeDCQGPSSeyDIufIZXLAoKgIMZ5eU/RqyMlvzO0y
mnypjdcp3GoZ6ArDvouynJULZeHgmuJGOT73MUBlqJfRN0N6ZMZkQ5d8M26W3Uhm
fO5rxAS0hekwb1D5wG9/G5fDtrXuE+woSuBz6YGVCESXoLvtgJRBVNf9RZp/1pfU
ksraP6UTDlkA0F4IYtoDN8qIR5/g1xgGr2u6jMDMIiMx9DBUJGPsyMCoSx8V4Fqb
uv0dhnCtSEgrYQQiSDo8pGnv0WP//1E64AAaIqD+pXLEuuNuARjySsKei/07Mv2H
065iRlkTwIrPW3cyiktMybWuv5F0uaaG2Z3uoPst18bv3qXep6fvfG5QVJ/ab7Wd
PTn07XeNkq5AcBwCp9Hi4eW0wd6beUY8i2KAe+bC1r1dLppUp8arQOVOAzZPuABt
6GbFqIU9Dq+/inRoLk8LZlkg/NF/C7FIKlh8B0O2o8u3wo6S+SUv7CWrXs4xxbgJ
MCX3qI7GOgP1seLbsfAt2nO1VnippE/OEQMCoZo/erdXPk6KOhZG+Db0xiRDhNEP
HzCCTM3mVkwp36+IWfFp60nlEjl1pzKtIKRpYPdwLRTYlPNaHJUz3ukUFvJqDy4E
eny0u5vdlCZUsUQ7QQt7XEPyEvzYydw4f3p530i4tqlq8oQf4k0oVeAFk1GZHjvq
Gqlsk1OCHQoJZyHsxClGiTlM9kF1q4pbd2GDb+/5jYnSgVvYwImu5uXlxG4W6/7A
dAiYw06/RoDLU8T8itCdILEww4hxEwI0i76dwSIIBIFaC51quI7M/AkEhaCEj8GX
Y8zMyKoDGZFsXbDL4rIa3zKREzAEZr+xHKceuQMJDUd9pl23l21FaNKI+/I52PEo
nNVNZQKXR/5OUIVdrylH+SmENeDDeUDpCeA7S07khAdVuUHQCQEzD9lEwS6bHcON
1Kf7FPLdBOM3W8ZR1IpsDd+A9E4feXq9FQ8TtNtRJv7Fdu3QEbeBDyTOGY3nYWty
/2ShmuJLXBS0iLWXzq5/DpSKEMQy+iFtGyIdw/SU4/G/IIc517gW084ktqOs5JK2
nC40HgxlU7YClnIo9kiJySMLRi8tDv69PEm3k7Xntja6zjHYH3hVIhD8ILXsawct
J8RaTWxCT5PGgCSaE5pOGawpUdJr4PAMzfFmKiYq1knxE2XPgU00mBgtPZCr+J1W
07PjZtZHsr2G4oImq2KUzRIOkqRT3u6AOiVHs42q94h9arkPHAPYe/fE/VXRq0Ps
YQUZWq94f6tyAwVINKQ8reNaIkJ3h+PXifOUXqEmiVgOgEmP/+ijvFHVTQjannN/
gtM7NjeCU4cIT8IiVZ4CJJ69Fy9CqRw5IAfc4EvWOYtxx77B7N0FjkwoMpec1zqW
d6odnMSfQ7GEet/7ktUQQGCRJq8Cr+KYlhrIoe2+u4Mf3jjmnQkGCJRCg9Cs8yA+
dDz7VQjqsqKQULoPQLvVjbLWw5U2aIMRjoUYynGCttERU7YNOTCZu/yvUSaPXUMh
TpWV4bp0gvRpJNWRJHlL5vwn1PLSsDfUZM0Yn3BpouI7J/q+Ok1vZ4ouOsIp5y2R
qO9N5ev6dFTkgU+6lT59XXQYVG4YZYfWQkBoimxYWSfdohBpS+/o2DlgkEInY0sN
YZshKdVLVZ6wRmV0J3IPdt5i6duL19hUhUacD5DJXRJEYOIrkHiMT2wSyQtyVMco
C21/oJXx3rCcmzrS+fbtI5rP+exqFf3QMyHk7uPzgQLgPtnnRJcsM/FUiUrv97IQ
tj24Z0wCro9vaDuhHXBLlaS1y4QQzX3HHPFIZ6LvLXNxRl4MBCibZ3B9LLQr9fvf
NooPUunQvKfcwerSXP7bceSFbfVWEVrtBVOMWsQUwVOeMMNa2jevP4JffZ8q//R4
TapPJfFq4UDQ2tM6HIKsZgCzHqMFxr9dYptS/bXK95PNQUxtX71ysg3KmMUg8PFo
nHxLLdZFiWHafaS/W4mMcstEetZZ08QtOU4GDLgXV3e2nXcXsSYq/M3pdtOzWml5
vtX4qiU6rwiKMp/6zyPBMlqhEHaLwENdftxcZqfuP7Jy1zrBIBA9jaoAmrDMd8X3
HMBjeydQofdJjSAniw9rA7iV6KMOpkHqBB1OR9w1U7x+xNJEZ2wG3V444m2qH5H4
Of84PFDuMkQ9JK9vM1r31wVbFPx5AkCXPl7hD5Y/pgpx7EENHfiM5f0HtIPeOVBH
7UWgUM6ymDQSxqUcOadT0xu1WWFsK7rTBTWyvf2898niMH6saqA52PLEO4LzL7FW
MJO/ySaKEcYLMchNoi3DsTObxQtYqNw+xHeYTSeLmESlJPDOydL3k+T3B3z7Lq6L
Opb9yG5e8dflKlb9F482c2R3kOjkwjNRqbw9Wgf1uXHQ7O2XPSgBY58rI//E+tc1
Xxl3dqp6imuSLyr6h2wrBG3r2MiGT6IfrS+61GmvqHDSQpt1X15Io6y90B9VN7gb
DYKu/+zpAOrPie4uzwurF36fdpOAOEWTSJwLzfHI/mVnpMahffm1JwIBNFkWJaEv
4io9VwCzL9YTlc7yuNRkdfcPTpqMC09jIoRy0abIoaqonVMa7GqAziRypLFsRZC2
++QwHwrEismdV/4B6uEAILm8AvFYCtLVEwOrtkR2X4gu9aLhImEXDLLkbXlscfeX
sEt+PqAIhtY04uaKiU9iTvU1iocPhe6uZpG2LHlmcuh1JKxhb/vS91+96Jb5YKcM
MUXluHOSwLUFc6CNxeLdUPskxw6xee2oleBqyZJ8guZny4iLiBf/J02vRXJW8Fqd
Ep55O1B8rP9uDwsrVe6vE9Rxp6Oy2rccJcXhehbX5uGVLixUal9rPvmClT0STs6G
JUNNq/g2Arz8pkBzrTRV93Vol0YMX55yN93W/4lqbU7Yx8hJ8kFGYHg2Lq/Wy+ut
pXNfgpLwzD6BPJqQG/rF+J0JNBlelF9D85yei7LFeXFbNjrSOSoFbdL40ch2z/PJ
9Wsy3XeRQFVb09B5aP9PU54arOgKz1nYmGuWpSGF8ySXftDBUPGH3dokNEPGDyuh
Kv9ClZIhqkSC3w7ENkKIlytnxMmxi7VwQEPYfyGZWnxAW4UKdx84JNpfqg3o68/S
kzkkWWKEQvqLd451XktpmgVLut5rHsZ19/AiwxsiRzlLLYdVy6/FQztat2z6fdYG
/CGbSnOi+ydS3vcO+1hjNbdtxJr8kEhj96GEnskI/yefuvBYvfqq+YeX1u7gJr83
AXuGcLUTU3MeNQBkIzZ+1alPXsa4OjOO3NgiumyukiqY5QQtGr8OlBl3o/4NLUVv
jcYgLyDdgIFn7gx9PPsHeDTbt1ML902bBni5uDXWGa9QY/XyrbUOBd8trKqVgWu3
PEuNvA23s1GoKDWuY6d2GOCHJjtMYZwdnChJthh42Ul3/QCZp5pOnRPrYEMiCpXi
nsCdw91dXx+vmiqTnTDxrnOkhKoziIzks1wQ0Io0xm8aWPkMPBXzu388ztHoyFg/
N9BSsCgsP+YoBpGFiosyp9WXhz3TgadI8sHiMgRj2qpbL2b+G0pAK9mKlc+dotLU
CDZRPRKQhbYNhAnF//bCtWtjQzLk/JDNhaWGjTwq+p0uhduLQXMrSafJVePSQPfS
WOYQ1je2ABXxgl3II9HS2tlcl/6vCbuQFta76i6bACUi384hT7Vkfwkln+gbNwHO
eNR1Jsjsby8OB4HK6agl8JuP7TTWOc+GvAcIr7VV6090nmvbrparIIjMElKsAPLY
bfTSGgR5TV807BawdYpbee22x39I07sQSvZ/skzYabX42XGbHBwTk4EP602oKwS9
rtw4IcnoGzZGr8hYoFfEhiTnzxMwnscoQ/+3xYD2MMKof/HvdTXtcX8aBrXd8YyW
OQwdwBifgGQfs7fQZPRPVEZqHXSi+RebtT/OGKcewKk/8OmiT1O+v6K4NolRYvwi
lZ89M2DgbBcOA1/ousSn1YBNuXfNyMjWZbhBVKHT0lLne6vsj2nMGzJK80Kmvd4m
KkmRbAoEf43fSGpOjua50mtKZCo6xCOQGt2ggxCCGcX71R/kqW1Ehx+3xAAOFnB3
qal55VnqJbwCB/kSMu48HE+xFq5chmNPrhdNmSci7x/lf4Y68mPMlmTGEFurLUuC
t85VsemMHMI9YF8uanfsoFT4G5l0eKgDJ2mWFo9HXM0CYrcP/TUc0TmSlC1jAptm
LaNcPCkf1SYu+T+GWUYzKWnjBUKDjLRX7K+EeV9t0b1vf0BBC/R5HhwPFSXqQGKx
/Mvyk4FAjuLD4VCd3Naf2LpNjWtdPzWuRHhu+kDawY+V6G8/VIUrygTh7k96johI
8/KnEUf/80i12NzWFyNSArcLaz4i0Ur6R6S4idz+vP7F0KjRKvC0AhMUOFGnBxOK
V+aify7lUSQal5ngUdaYxWUtjtreSrmibC/lUJOKd+G+Er4EdjSNu/R5qpA1HI46
CMtanB3ow5A86hhr+m9FbDTvBIMcRxgCUQSoerNXKgVuIjflgIyzgEoP+pLVu76O
+HMJwLHAsNDQX1MNYrHcEoL/NsCjLLHcU2TfDElA3l9l2tf9Zf2LUA9IknChE9J9
nBmKJdXmUK456mrOSp0W1zuHTfG+dAleVyQ8aknQhucEle2Ry4WSrTBmbKLzYJQO
XVr0vefMVlSiXoFf1J4adfpxTwECjV8Pc1q0N/940jyhK50Ki8Ibqac8HRm24Ihz
3es13Q84tYQ29hgwQA6JX6R0sDWRdw/dZs9PiiT6xsDRhDJZw6cJncWG9NCEgTcM
z227345whJbvkxuA2n9pM2GoJ+flhjXrCtg50ybmCCx+PaCbus0Oix+XvMqRjeU/
ayBNt2gz3txKyDBkXcGUsV9pb8ZU1u0XQyxPVOu5PbKogVQfRpKmpTr4x9ep6Fku
fkfjVV06yEBOHvqtK0nJ1Yp55Y+5XPwWnTXhodKn+snvH1f+WsOOYREOfESczV4y
bQeKPWPKB1Rd6t0r5wpMvANP1gT7Psw9ktKYRLlfgk53+ggSIbW0ZVrm0FVSs0gY
g9Um8BEyVh9rXzkjAlYypI1gNzrMq1eMu46NHB5BheqUTrXTnnGgRO7+E9TaZY89
zcDnMvzjSW+WQGGSAdvnt/Z+kT5SwEZEJzLsqavUbRuywLs94PT+D7D5gKVcpZmP
t0sO0ZsgnVZJnzDfXDfB431PCMu1QsA3Z3fLGmDs++pM5K+9rVYgYucze+qIyQr7
HZ3U64CydARN/gRhNT4Tp7cf8NCziECJmG3bvC1Pab+E4vcdUdxx/FTaGnntxI6l
8unj9u+K62JUnO1Dpk0tktSwEROWNVUlTD1oGwCLPjT3xzq1ZCjjeqoDJHWpaCrW
glXdtEvo1WzEOureh9XQ2DGdLbjODuym2kZdU7Khbg9YHSP5iajqYkz5aACkx2PJ
Bp5E6L75v8+vivrwBUjR+n1rIaA5RBi10YO9co2qqE55uIi9QJWwoi9Eny4rdmmi
aoi5Abc/HTJBJ1ueMwIfk0ig6N4Y0m/5cV7e6fdUY+g848+hnjLFgiGTbplzo5BM
7kM/b4onbD0Dy5H5WKFlmwuZ42/yAPFxOa0Ac4LRaUTUKi9ZcK0Fz6OLYxzG81dy
ZxUWhlPNHv7FFosr5plzkpxgTsMgKv+TXSbzJ5khAgeqJSdSIbDfa2d7E6SZNXo9
tykf82Hig0+nA19YKeEkpNFOzP4JSKFxMT63Omy4igs9q/2CMPEeleD+x6cO/op6
4+Iv3KGioKLV8gHnH+nyVfvc+J4i6D5gJf1CE4ygCfA8020BeuQGPGdWLoqXrj9S
JF7H1IPDLpYBXcUhaux3yueqzSvHVXGm9aTz1E9JWjRMISKfDpfESJ/ZBS8Hx7F2
+T4rypvGMNVEXu7JHPRkqa208MywMuO5SD7LygtJOxdTRQfEvdF0UQxORXVHUS/9
q6dfRzR0q7Bq4QXRhwPMjYg490F8ed/zkGa6sUSsOZ/37Fs3ETw2TTE/DbRO6rjY
3tLrpugpz7wfXbGEYCHutEApdIV8fNz4J+5BcML93quIpI1vNCgiyCJNgiqYHTRe
kc8NHGrIgngaGZbV3iyGz+RXDnR0tWr59DIJDj8FydCMwQeNYsYy8rN/DFJGh2XW
uvOGtDU9JrJTU+XslERdTlhQzndrIZb2opRCCzeoMuWa+76Lvm5J2pMHVawgRL3N
CVzCNaFgC0fbpIqE0MvHCmgs5yMhAmhRl4a1FqtCapwJn3X9S6FaCUYQYZAvMuC4
srarW82OOs13F69ycCY5BqDifKAmquZhfwFGCTlwGFIah0tI5nytHWhnIkhnT/A1
+QzTMnIz2acdRnjLsq9BnywbB9Zsjv2yoOtsBGDKyEyqITlA/1dlz0ZxYt0re4JU
/JT2GNsedVrYM8wxycpDDJAfrAIP8K6dtE8uajF8p7O1FwXir2jwhZG4v9lsX9cs
Av8M3D5ymUKJX6xMDSd8it0N1IcZc2M3lbA+Qrz9nHk08dQMM97TiRwHKAvgs/Zd
RMRW9bwJLTm1vyoT8QyP4q8WfYHk5SLGm7i0m+ZjHucTa7ISkJ4CKLs1v3S8T1lg
32eFn0XMmMwHaFlor86pFQB/VtffNADLNyLXWoU+6R3LxeBQhNIIZOiGwkU98Pg9
AQeA9lO4L6QpjIn/OueAjN6BnVyjUhGavyDWOoGjELAq7oeL2rtHPdAEI3n+rT+o
xtapDCWy3Zjk0uMk7iwYHapDRNXAfH5+zr61NwBHADdCLKmQPNAm3AznvwA2Tgd7
6u2/QlNGXFJpgNCc5GuByBqkmNY3ZKhRT+mx6zxRsFGyfpso/yUoM5snUjW2de0w
kZdvZPV266jCXAgl+aGnXhefkM5a4HLtmt+jjL0K4wGFcpgeo8dhMxv/cB4EpHTw
qXMjQQrNJhyLD+rTLgGpCLauZ0jfYuFpXIsQxKltELx5N/0HskwxK30YuhNbVd3E
QFuyFXvFCv4FBvSOiSns+ZvNBpBbeRHnYycA6rdt3e/eUADGLd1u5Oq6Nwsg1FCp
XcR0uq3NBH3gdegeY+hDLNjJbSDVtI8N8vgja8R0tNglnqmjaDMTH4MQIENa+0RI
httNg2fzZM1GjbrgU+SOT0/AAapoYtM1wKJ8/KYvo82Xyar9eIqsde7mf/riJvmC
FgU3EVQ2C7BJjyItRoH35QDZqfQlyIb57HMaYhFM50e1/q9fvZDCImIFzy7FN5UI
8i4O7Feian4JaYZmBLNhz8vUsl4qPQCUmzMKOsbIrGmgnB90S+nx5/uEE7Wl+FIZ
JGhbVymyZvHRoTxsrHIkSyXGrAPiY40+2KjIf7VIRajUQHyeqT73VTRDpsOjFl/3
HRXdxdMw6pFJfiT2D7lPETZGQzXWYMKl8y7yf3vI5lL99XbgX9sRDXJSjOM3HGCs
wcmtFdSZzjao/0P+XgRgQX5FE+MiSvO1c2O2s0f+4v6ZQqGb6JdERhr3YGwceKc9
Sgk0lIevDTZIV2vE3krgB0k2ZMJISoSKf+bodbPxhdHWYOBOlRWsfQvc4ZNDxbHF
wjPHB9sDNCUCHV0TcBHJsY/kqQykjHD2showjKqEqQO6/RyhTDVZVnkSyrmRJaGI
Wc93YKf2TCWwyujKcLjkeSt/LIvE/3Ix7S9tjwlx7NXgyvpyw/BfvTmgOfTw/be/
5velkVEu079R6UsbSHb9QVkh7LL8kBakPOrDrHlthGDylGqdWPUZ1XTCqTKzM8ET
wOTzOo4rWIAtjp7LUM6oSOdLKScm4RvYAvpc4t9w8L5cE6BfaWwmcclTcLG411DE
kzdx3wALI8WmZDO3Tl3AwSqyWDuV8/HpBBF5mz6OufdeDIrOASq+UBqXqfqnsbe2
VwYqratC747mWpK/YunWe0gQQkmbP0GaNk+QSra/agSAYBcKlwbu2/VwXe4VlJ1/
AAtuixgU0NUgFp00LHDfBSKAFhavoHg/wDig0FmaDP7j0L8DS/lmIfZOk7oytIma
OdIPGB/wXULfuTLKLt98N7BGEJohCMJhfNm97pUs/OnFZAODoMcbHW690LscTGOA
yv2YT4cauHkRhpIKOmhCky8Tr11Hw21McFh/HCGQGmum/ROj9kuO8AkTkBpAIC3j
qUWOFHtqSlsl048Bf869IEf0qXJ3Sz9zyjmBrKhAkbubEZFICD1yfCEnybLkGBFC
QYE9diN+wGk96VItsahR7ARG3AtTuDdJpla1gvICJJi9vRxrrho8D89cYcKsjN87
HeouA+cc+q3NNxEdPDwKC58m8aQezrEZxhWtE6IPwvsY7EjNaEh6CQjB7pPOmlPN
5NLcfNU+dsTXQL7MpSItggozMJvfYy4/G5xwETeUFYq3sfiDeg+kk7xbYVWDmZbm
Rbcx0NzOiPyjNl7gG9KazJOoQZ67TT0FMS/+NFRklYp7IDGVWMxaODuIdvYVO/k5
b8VhRZPsmzoyc9ULN7Eu3pSQfs+Ght8xpzLUncyVNHNIA5K/3IjjZS5388n/CscQ
ZdG6ph+JVRC6zB1ap2B/K0YjNf514TcHMC1aJpzEqQGfafWSarLrXEvojqP8JKEV
Gr/xbDalMwsR2haFecV21Yq9njrndDoE0ECxgYwq6YQ0DKgusPw8gkLJwJRHEThI
9/kCI403GCDBvBgnfc4HhmLmd97csvwUcWhgN+Ck5v6WfQ7n8fCwZsIuIHEpMkf9
9sCKtAjS5/sNt+TicYrJjFbDudidQmprIua6wQe57FJSfotyOEwy6XWLeyju3Bnw
2NiNCD/flIYAo6H1DGvInoTerE3Bdq0ez4y3tfqXo0Wh8KZZVXQN8YAsC55SDAO8
32nlDKKD6sGesoX7iRpVZAoC5KdNsUIkdlqplLI1zrI1nsKhoZRGc2mDhha+D4/x
tJipFuLOSxeHlJ4jsPITOFlMqGPgalKsE/UiyqJQJRHTsG4oVGiG60JLyPghSRi5
6B40KgmH9zpYUJK8xgr67xBqQgfPX7LwgbjK0xTtYrlI2w/RXtjvqDa8tDOU1uyC
RbDdhkx6o3HzSREt4g0hHqvlKgppz8UwJBWZS9G4GjnMJEwToD57oLlLiyym+wir
zwCN+dci31z6+wd2tmNIQ3RD+lNNJpH5nWx62Feh6H/Dsgr/78J8tWeSR46ANjEu
PYHGj00pg5ieuzJeBRCRLqzWEDsGl5Vzv+nAkgQO20cLOAQZLEfzCNti5+07qFnJ
xgkmJ98rCp7QSPaLDC0hzjIwstQgrfOSLK63QDCVkInhG5rH+ohKc/c5geKOk3gv
v6kRyGTuqTEOu+gGl7U88nVEdcOss3AxJwvcxzrU8MqhkIISjxkk3cBQwq5Lw2id
U5oXXNi9UuFrNfCIcvk9V2dsyCeMJTduLYLE7uyxUlcRaTO2N790Xj7KVrdgvH7i
0d6nmH6CTrAWUjhYKvNDWSCj5qnPi/Sg3yWmPviWHIXBlze8kqpdB/vmxjU8NcuT
TDGqvdWxZilK6XyFkzKKfSH3DNUT9bI38a2Rf5zs7Kb5bwTDeB3Fik/zh8ulw4Gh
fhQKhjSRHVZcV7ysLrBKzNPedr4yXyPULcWi9h82sekOsfabOlkPufWwVJeJ4XBQ
XaYRaOH1ncyWw7six64bWEsjhEL0TZgtSwSR4WXot6kN/npO5ndW0qdtIrBGpEbI
HFJJ7KrX8AaMKCNY85kdcJmE2+p2FPh5ahKJusflzgtIJW1BpKvQUmU4RPDYy1IG
rcRpLwSyGlzVhZBq6dlyKyzmKFDhl3XJL6FIN4rIU6QxhA+zvdxBB/s4a+hBNiUg
YNjmCZMOeCC1SdqDlPCLDUvv5G7zrWZHW9p3fdUpQqLpo556WuPQnK8mjE1dWr5T
5Y0S+t/7Rswn+u84LKv7S+5xKHXckAoFo6Sptr9sMe48Hzjoxcuasg85YfajM8V1
8J/Ch4LT4SGM9iJAWR2r0MZ8IPEBJp7CIVJj3oDtHQ0YaiQhs2javrV2nxc3oz+r
IqpTDeUJ8g1F+5hvau0vKdRKeVYEQyk8PsbhJvvADKU0JuulEDw+W0kV+b813AmG
nTm3LuQIne97k/sBEUpHRhqu3SGtbHB8sfyjqki1LLdO+DlLNHyEG6DvwPA4fBkN
dRifgCUtR+Ad+36itQBBBfVddU2xjPYp+6L1O3ZWieWkEZeP4Lg4c0twfNQrtNdz
J5COMov4ahE8nUu9ORksZeKP7rhz3AQUvRdTsL8kP+IEdvc0KUcWtfR0+dt1vrSP
VA9WQjcuY4FviYs8DJleyr5PXWnsViG69aDUWKMar75tRLWetvSfl4UdCuN+N6bh
vFLy3vidAvA97W61BeAWtEsQqEjE0Yp3GCt5TFE6rkGphCbPJaGo9ysfLEeQup8/
D1cA+SSaLXrsocIWDhuIPLYNNGpwqcEyyJANvTZzuEzWPa7sLJL3v8wxeVFqk7t6
pL2fwQkHLdSBow8+hB6oIxLtalpl9gxCPXIng2bRLoAdivuRCbIR3g4YZSS0MSy6
ze1XgJTh2anpsXn4qNYOA7ZR+Rnxz5x2xh87l7UEau+3LqQCDYCyPjMCeBeTXC9o
ngbqNE+CWB5GY6+pnsXkqkUkSJUccK+HlSsh+1HNBsE+pvI90ZNrChO+w4k/oDSX
x5NX1sma97mHOHzI5zc5BJdoW9sJUDTZWTuA/fvcyilDhCYVo+0aZtFMy58t643C
FnL+mwB+BpWGAYko6aCcQaiRX5mDcI69XkQNwUYzzAP2EIxy12xFmPU42NOEeoAm
6PPezPyEE1JYQIdpRVarTBdHXxh+f34wt4UHMh7zzdmjhVVRAFVZapM4Gsze7VCN
IgMeW7laajhC4QI+joo5I+o44TpfEhU4aSd5S+qks4jhfZ2lb4uBcvZgm8YcyeOr
e0gf9XqQ+/dyblqinpLhKrcdhVsJnhA5qE0Ha5YNKxygw0azZEW3WgxZnqW+3uSu
O5vfwbLCBNHvZTJixvvudIhIZ5LJCW40tdb+F0lY4khvmNRdKD4mklHd069YPWSY
i7fz3Azdu0DOQicQqkB1WokQsQ0oTCS12SAbgLe7QaLUcIVbpYL+YHHbUVJFTouh
hVRnpWd0fer1EOEJ8XWPYD9mJox/dD2I4T0jVJcvQ9EQzFw8zukn/49Sgq0FOV3N
IPdukeo/A+LHehSFqfpxNQpnAqxdvBsOLsrc7L7mFOytzq3op9xspbSpuoEpCj3y
xcESv3/q1RFpoQ70sBSP24YuoxedjrcQa65SyOxlcpMTS/Un07zBtCF6wzLgG5Yo
zc8NCOymTvO9J29tzInzIfAso1BRveRnP3vK/QN78Pj4iRPxGwktnRZ8xd3u8/YJ
K3GTyKLgoPXh65MmP+2cJau3e4dL8rNc7R7Y6N5yetdsY6mwqfQIwdxYtq83PAaK
Ojb2Kpiu4UC+IZtoZqONDIDi6htaqikshVknS79hzLasmndsaQkzgS6QIFH8DqkP
RjTKdpOqnCpcq92cihPChQxvPpQimDBgVjtJVhG2OQLK/5UxhRwAsbUjbM2t0E5x
itNsnMdlG1d9aojdPUtkekUqZzq2OudGoHfYCPenrV7xwhPM5PacNM2Jub3AMkUW
ZacYITTh8AZplgud0h4geqmLIkz/gXOVB0SPpi2/OPUbE3um2R/+DErDUMhHYHfM
P6+3457J7pUSeVnDka4HFzVgRQsTpuzJ3mnIbfRBUi7kEgu9uMNWVgpixFrMjW9P
9aiMbst4H/2mQeyGCknYvkgIhtyYWcOjM1J69WWeE7deM3HxnGqq9CVovZdujcRC
ouv45KaM+KcUUw8geblYXgpRcvI7czPYQAQMgG66RLDebreNVGAFO9A4Myj79STG
Jgo3FlywTu6/eEn8jvBmgE1dWFcwD+g+2eFnPiovr3RpDcBeHhNAlnrA0u7hfN7U
A1BPpS4XSppyqWwVCHGYdGULIAoYY9LYkJTsPV7TISFoib5AXS0MoV0l8abOGiPL
sWmq+ohrKSAhWiNdm7ZbcfJJzvvWiOH0Xg/aYdIztlCNcHUWfTZ2uTOe0UGL1WZS
ZHPV0VOIptMNAKYx/1MwHiUySiz1KXO4Mu1Gx5tooiOfU8+w7T4v0v1deVqAyhRX
Pk+TUcwnMu9lmcK1avkcm/4rxpk/6BBLsh05EfwmZY8NFMGPSNA+OutzllHbSPiB
eFtnYM3aC0bog2T0U9vSYrb4JuCpldOudZpSq9cprVN8e5v3T/q574e4mYiNdYiF
492tzQIyjVNm0ZW4TucmZH0/oitafZrKwkEFHpIL+8ne3DW5GeLN+H32KagSKbhE
1EDaj/NntzOpQh2IgJNDsUmOz4agmEdfNSItHXh4ae0NwB8flmwePseR0TIKh8tc
XikBlP761aQDRvxmOCXP1UN04fJ1UN1wb1IBRmHU0HkBSlSKcapr71PoARFZnP3n
tHr1dzwISD2gBLQdkfqryjngPJ5HVM+zhzQPh6j+mCsRAuqxPgDusai73BTXBkyo
sRv0wKqQn2mrcll0RYZs5EXlrpdFdeXrpED9XUgPBSvC2Hzsp5ZLY11uGtQpzXBq
s97jz0lcO/m5knxK0R9xY9nqOmNl1GingKlc8O5XeBV8MDWJUq45PjddHmRVxX+K
SiYGvgtVna36IZ1X7LUnEvbiLzSccHl9aTtXL1Dafr/EjYBGol5Iy7rmAMCAv9DS
P6K54333r5CVrjJAaBr5v2a703z4H3zFX2fg4SuMTfOmhMZ808g1BR1PiBSO/9DP
ai0yqDgteP85+Smtkawo2VQCJX2lWun31g8Cwr3qImfrsXhIkT8RZKFitWi/YpiT
rXryuEAJJMKrrGPUzoiuow9a6sD6e5xnRNlN5kYqVcZqPfkHTveRLaASlvTJTF6z
DCJz5cNmDi4hGS5CGcOFU5dbCL+61vBCcUsvCey7z7SSg9HMbD0CrURhNz3zroth
l9oPK38xxaJ+h43BBxIzXouq+E6UvYRhf+18mmXoJ5wgFSNTzQVPIQ30O1OumAtQ
YZFkHnSBmy46SmbMeY6BbTSh/CBlLhMUWSKaYc2iRasbcXg1aqmAQvAA7OojH1rN
UXz98bDD3t8q9tyuFilhPDQNuviQ8RYCdlFcmsQOKfqnkbnuOuTwbDI+khN2tLtH
1aNPy1ZzaPEDHNMuYEsa4Pnvds3FzTNM1Fw71GLbDoR7bJfrzDauYXTGdHniR1mV
86RNChFc1i2gD75P9UN97WZCx+zYa/9xa+09TxgWC6M9CZi3UYKsyPYC/E+XZLuS
LSu2yGDfkwci5dWW4VBmX1sr0eMe8Pv1xR+c2UbnNvoDq1H8mIXfB1v9WIdkhSk3
2BoJgFFSX6ImubSg4+Gr8iONBsR8ZBr8YsbXhEdYPLHHXtIA0JItZ1rOxY8F+nZi
xmN6qdDDHqT+N2RRoO8TTrsWPMgTBgdutla1gMnoC3cNiKtaqKtMXBWKw/Pc1DeW
Sx4ZWbxQegNfalc77GMPE/+9PDJgV9sDIW53DVPSYEYml6JZqrGaax/IfS7GWKSw
qg51EcA4vSWSqft1pAiCS8jvEPwJuXdvsSyFjH4HEb19g+lAgMJhWJ9rEZ+n3igK
Ej/0h/u8folpxWad906WD2rAOanxIOoZMdMr8JQwlHcA8n/jA9sjfYAr39J5dATB
WAJFXwRmUn3xBgC50FHgth3OJ8itncVuhmO0anNE1hyA+/0mIXsit0hdZAajgpuY
9UaN4/tZWbzExNsKSM+J9uRQF69917rdR4jXOmikPFq0gVDrJ5ZlPAcf8Yfp6SGk
FiK+0GnvRFSmoZ3nzo02Q+ZBIn6CCDznOe43l10iu2DULI36F6sNOe+ia9ONrZRD
OnmZ2UY+9YBCuwnNeqeIVgqfe4qXQxko4qc2TmSVLCpKqgBxmmnt97FQlviN7LXt
nzPMDqDTOnhTJ07t9X4WK7GxMh24tWLPq+4kg3bCw2/D9MdPNx5MvhT7XVU2pL3H
tkHeej9xPRf3rrjbPqjh2RAhM92dPfgjwaRhIyXpoG0RhbowZmYBYGMho9YkZwI0
E3Ijx9Er3H+IVe710HBAxtOqMZFqgWJmPVuwlbPF1DlYX5N7as/NtAAoEA8yD2Py
BJfRoltpKIKkVhe/JeHEdP1Mgy4STHuZ0l8Hw/NvbEtvWGFE9WNNz+ZE1QFuWKLM
odXx8xYnGYpeInGaySSTx0hoQuszHO2wuIvc/VZpyTU3qpqQnqGkQJ0jh120aNhV
KEJDjHSTUC3s+ouQtvq1bup9ZUCbaI5ZKmpfBRskMVj4uJSYxvAUA892Lr7iWLrh
FM1abthLMpCQdot0JBpjcL1Aytyu7RxkkCVt28/WAbVAEOw6o01vqyLMgL9baJTe
VmAjeohthiBUi2cSbTtoEV4MFK8sIQf0ybgMWY8Mkb8Pa/rcojTIgvvosf0OvTxd
K5aQ9TNIVH18okCcZQR0PJ7S/SSCt416TCB0Rbrf359Mz8JQ164GqguVWXxsrqj3
U0a7itSmYVQ7SwpR3vHLajL68ggtlyMWMbpOml8Dr9ZT3UxynJLwZAzFgerYqHLn
HWWHZfg/SIO7mYnLVRcjfqbsWEOMV8RpXMYbug7rOxrL6mmQKxWVWPHkrZ0kCX8E
f5dOi/G4IH5kDJ2K+tNHo1U7GWNezp61aT+qYpnsLnLNGDKwuaXOPlGE5RpWTmkG
zVy7/Bl5gQjqW8581JBBUthlA7cFaQdnIN8kUwxk6k6Acb96S7rx3Yh06ZMiYP0X
9+/sy9JskpSfPbAVJl3+SJAe6ML9t8l1U1k+c93QtYchOaKHpWqLfUb1KyDsxrJs
vNcJn6I2GS0/LXxqYa3C0aZjLIWUFyFhB3RghmelfJ2Qdlx2rJ4Ti0+zqlr4y+nU
XqFpXTqmqBhEab9sYELzogqFoJM1JvlWj19e06owPOXyEsBoaXwbjP/1O/Dy5xpB
RFLJsGD1gIkYVGmy3btK8fX2/nu0qWjdzgA1qjS/9BIsXFN88RWaAPLvYBOVEoli
WJtkxJy+P/HVoDn+L92K21y0X4SlJxpG2qdh79oLSmPcCiWWIGXvxPMUbiiPtski
Q4gP7eLW34cu0VcHW+3rv2S04jUXqx+B3ACEU71G5pWemOnx5N8R9zKE09ZLlI3l
FYX3Kmd33quWv5Qpck4RNesj4jFQHK0u/vgGqxcq3KkdlfvfTC51b0mBVGaSGR7b
bYxGFfnD8S7Iz1+MDR0wTCtU3zity5WmVUXJpT8QvMmC8s0+9WBIrE2YiToE7FxZ
VkUR293sCYaRUU1jp+OUjSiOkCcE3OTzYNEHzpl2MYVG0pAHjcJNmb4gMp2qNhS0
2N30DdszwRu6YqoAD61Qnn4K9xlfpxLFKPuomflgpeWJzeqEETdyT/y+Gak3uzcw
HwokaFR6IONT4NQHUFwh0yZbHiJAyqQh0xI+ofrS5ZN94Ax3uDJ2X9FsaeB8Zrd1
phvCWtminyR8A7gq8Ien459dY3YikLtaN7cNK7Okducq2gzvjGHVI1oiKwO0rAQj
X9qs5nssbV/bPNz2IgLbPpVetf+ARLB9bvm3H+juWTQ3jQnQZEfZ6Kx/sBrYzkDm
BGcseorASUaYXEvZMb+Ek+jkSjJX+8OgZnTiYOv5SSaj1vgZjG1hs908jKS2ZKyP
3JR5anYPCStVxSEQ3QnENXhaCi7UKUxq1pVHgouGTyfsnuY2Rn+gjzoIC/FDIE4M
/3O6sWqwm70+yq+f9JJbb8Kqq4Ie2VfFH/ouiJ1enNlDFRJcQ6BXC4R0xZDtQZuS
UXxboNcw5w1wnASEooWbnI2hRKWet5ByRQpl48YHFrYPxzWMikrlCBJ09ouG0KP1
P+hF6CGoDssF/RyQNDUfnhbWTmcM+o0ACKxA64TqjmvvdPXirRz1CvDRUr6vKwHz
sbyTikljhnGcPszDYwt7VuE6ydPQzh+rS1gwXcLbkwR2RmwAr1dUHat7yGZoSpxd
dALkUgI5T2ricxWZmqD5pGZXcxKucNd1ebdZovnbJLJ3PbIRm4/37U4jB/xSIw8q
ZL63kX873nIT2Ny/d/3lTnQ0yhIEiSEuoGYSMwlvDXpsHwg2ZTInsBWv2nTthQpI
SsjdEu/T+bp7FpvofDMYAbu+FtnPTsb30VyCRnZ2Hi1GM9SvpWGhdaShSFhS9q/D
hm2com0Bj+6N0FbBeA/bv8Es+kYl4MT19iHOnZsK2MfclUQ6vscMiG1clucFb4z/
RGE+nQBub7TZm/N3Qc5NbR/3nIzadY2eFCJHTDX/uJtCfdrX9owhGmcGJv84Q84p
KwXkPKU1+yW7QYe9w/cUBlpc1OelxNH2dXopFIKf+LbyQ76yZ88dVXJxx96OYqTY
DdR8Md+G9f3tlcyO1g5XYh3ZJl/huQGP+7UUJ9e3nkyK5P+PrlifjJ0kSj3n7cf4
bduFVbMq4tS/VHuee69bK2AZ86lHoynjMTOZ1HtZakpNY3o0hduEIjGDdDHTatkF
m4Jfn2cPkN8QPWwbZi0gR0A912tTI1mAiE2lkAqKiiBo1MhlSAf90SorkaiHmgnX
cO65xX9alPedFtNvxa9uJDK0rvMWyGT24BmG3e0aUMe66H+O/04Dp/5XzpYzbm8i
Mf3206X7eXZ8bYleN4uxRD09Lh4yGswB8kN+1s4ZIPze2LYav6Za64lPdyrFPKcj
Mt2g+xSgmwysrm/ADynQgVVeOlQKxuZ96febHoV52n83A3REk6JQsXCHAfprL8L6
rs2MM9S37hDCzIRc9dBpqMwQmbRZsw5hDCcLGU7XcfJaLPF2svmic3OJwW5Wb27w
vJEEPXiwRmswwAfe71sj8Zg8rRKksLUHeqkj8+Amv9XrBmImYliN3WwzfN1un9Fg
B9hnHjK8ifaUIr6qpeakbrqlBjmfOPnEHJhVK7NOLJf8Lj1l7mUX/FAVeWAP/NHb
UhGvh7ws7kliBtZ9Y1P5RM5UB9xy3IBi1bAba1RhPzChmnzUReXkWUFZQ6unhOr/
wksm2Q13HLLupRyZxjybIqWomkmkwpGIW9Di7I5kxfOuHEGsabC42hERN59Bn39l
4I2OpIdxUSE7NbrnVHtGin5cmJa9gUrFZVFVXbdn2XAomF1H+vG7Olw1Gf9BfT/1
XLTYuUullGXl/KmC7DgetUT91uII9Ooui4aHq5YYW2jANrHyNOHPb8evT2JioImm
ThHeaLayzFU35QCj6BzYhcxnIisgnBMaxnwma6yiNkGQhUnF7ajFUU9N/Il7lSmX
a14m+Ketf2aOWNPaxan+zAZWwrRKdoDGNJEDNu8kay/Gmx7g68asWTrOi4vflHhp
N3Ll9luB5PFyNXda7MdR101QkpCv0rF/ZYj6GXjNH9EZFVP4t7F4FpbXH2y4C6hE
sfJAR+Pj+BWpmewBir59HjpeUXKmiGJ6o2QogYZ/qcYTLfZrA4b7SF5Hm273zTY4
QqecgzEBtff01szRcvnVxCLkZZPp2ry36QkrIlHsNxBo6DnLIMckb1lPpLO5gLhT
bixC0SkJYhCCHkUQcFG0owQyAlo6NtxWDScHVJ2kW3pyVLr1iRPcSYbisc77SosZ
3SLeu4YKXfwZCsLbP3ubEUy04mZxsxd7C4wYcF3TZlJiOA5cihq7QsIMryFElHLD
AR4cGzTltHYf5Ej0IlRm1x8bI+CEMg10kk5yTyPgqdinvQcVSwbWyDwOLtc7h2Rz
DzX0G50UQJPHw/n7hAjIb8Xdi6aVh17dqJ8CbUp8Yg4p3kgXEea/HppOxEmSX+vG
9bzGXLTqETyR156mW7eCx1Ip4hfeyrH+VzBBXM/NxvRGF+QV6Mcv/8p0OWor4HuM
J1G5mkhl/4JiGXgboxu2vh1NGrZygChmS/ZQiz6vF259/l6XdM0fQ/pG5YO0hABx
oHezk2U0iwW+w7aLvxdtG1m16yC/WwR9hPAHoCGpCwQKqaod3f6UgybDrmpyr0Pt
2h/JPqkapZwPKfDh6LADhxOcCIinWekPqPtLqfl03pvTc3i6ni/L2XheiIWzU5zb
C+ZDb4sfKK4aMpqtOKQw72CbYyOaUpMeqx9+zfa65hXjPFWlRTDRhHh4BuiPszc4
heZAmvWckKn/H3s/ID5EkGoO1dvALSycRyQ4iEPK6zGSBpYYtmfhRlosuLi9QsF6
UjfM6YiOs1OT+fnjIA6d4B35icwk3fsH4l7Sq/iHUAwN52cu3k8nWD5FvhffgJK6
53eu6BTRhGl6eFYPk0ncEblvLdOZQRG+uh8+zQXVeEossWQ2YoZuUece7ZuzDd3o
UbZ1VEjPnGlcvAZAVbg+qI+f8rWYiw2Rnihp5KI0NDU4UaJ2AQspjtgv7HfUoW+X
poAal8/2dkYQv+95qI6yuu5ki9SoEYkyS3+VxsCFCHEeDSgTJvURXM6IFQaSm3bw
JeA7dfqNQfzv6kyqxmy5CM2xy5Rd0ASTlMPY3wcJ3QP4UG9wp2AR3tv1Ax5CkJR3
rwXFUrYcUUP2/r0vWM2hvlFMCQBCLrFCDhXMCyzfXanLMBOMl4odHkcKmn5GF3xx
94UKBv2zsh6YD6ZZBLPe7phqm11+Cy5fHQQwyAzV96NU7bQlfR0cOemxY2r76OKv
zI4+b72PtFdYRCIkFYe4AeicWWPXSyaFrWV6J+Hmv2JlbsygIbzCco8x5LI1p/fr
xZTKcd/RycYSvGGurxrglgC1gA2Bz575+R7XwpIo3JT3QzmK11o3r1UJX11bdM2r
x4Oj+PUK/ENa01ikcU5O4+2FGsDps1kZfCxq29IiX0A/90jTRrZTiN7LHB/Ije0a
TeRKIxbtSAkM/BF0AynJ1f/uTQs7Hk2LIj+yfs4awIfwNDSWPn7JB8YINPVm+4vo
Lx9trRfMGNVYXB27i3W/wRwlC25o+6ba4mL5KlDh1LmtYXr4jNku/ssdchrCADwS
lrHNH9WqmdS6bw8WIriAgYQY5DCYW/vz1G9wpz7z5bNNwtcCAlhVLSmcjegKy3CC
gUqbmvbuMDoFsybjVowHM+FZLvcc398+/I7y7/5JFoBVi96MMYCAmghGD1nB41gd
U/AvItiA5epsySPCUyEJd8fIdd97hfR2Vr+9+jGRlhX9M5SGjZxr8EKWg7mar+84
wP/yTmbS0GqRlAr49abnMdagl35gXltWi7Jt6NkSEpdtHttI8jTLETCNXEDowmIp
tfxA9+wbiu8IBqhgduNY8AxQNDbuVURx8f4fliSmmJAurC3NbC54FY+kRGlyMvED
WCy7AQR9Fl/1G/D4oE1o7yy1vf0jcAHeg6RBNQNJ0A+ov8Pi+owIuqGirFLvhsKl
NpEoZVSeISxwhCRwMnvP4xPnsYbilPFZ6Dw/em2AYpS/nxO22+slyNKKWpoCw8kb
ncqKcs6wNuKznEaMfMpfRaNO7PEBL8c7QZkvdFIa25dcbtbmaXPWHH4RGnfP89Vo
Z4CRgk0LPHNplDGj8yh0TLI627+Z8UEN8otcTUxSK9rC1aFO2B2YqkfzrmZ2B4vK
1OTraATz6T5o/wkcfNOmPznR+Wal//KBoo4VF8jm+LDd0IJ/G0h2NJb0lIHk1OIS
ji6TdunfXBdF0ZqgGyFhh5FeRHpMMvF8cWYR32Is9+N5s85QI2iZ3+3Fq74XNmlB
ULomSqDt2Ig73eMGn4MOGO+ROjYBD4nlbxb3bhJqGn/Y9cMAleNO4tRADMCP+MIR
0w0glnaliG7yHrlK3fNvTcJnesHDA0NRdDndjJhWc9euIwEBSDaIdwq+d8dSRKup
jGRpigvDJTEKlehRY0/jMRG4twR6WnKcEdK2shL/rxMiCLkJFYcC7I6ScC2vnibS
9onXEZvXRwEmJeozs/fj8wWi6Vx62iqj5/KMCNALQovjf6Maw1h1cY1cfg5M0l8d
HIEgxHAZIsQVbi/XHbTYkg3T6o7yun6oz7+YjWPtTuCRb9ikNttZ+xfR7S45I84h
O3X9wfXcmUYmAXfcE3aQo2R/KKmRRFDsXGThloMzhjhMvdrhrJz7vcUcObtfI6r9
pLhrpKANWO3F56n1pOZEj6nju+J0rgKcDAtBuoEtB/yBHb2KY1Qr/cs+WkJvBXff
HUgXoKqjegkjIIhzDPCI8jXer0VpvLQsD4tDMVAataXY68EIIAb7ykbNLqdcAtS7
+5jqbqIVzav2K6NpgqSmGQTtFfpXTYyf1KMRE+0VqcYLx02ukoPxNWdtD0JYb0tC
gP8yYSMnEeZunRnPMcF15S1NWI6yy6xmYUKfAmXPExRG+8pBgKfayfTkj9EcG6Ni
CF2YY/rDglR44xoIxK9m/r0ZrwqVzRYtUqtLswLRAQAeZ3Qbhoe1xMkwAZbW6yL4
kWXFRMa2ceQS3nDzPJTRcYPxmcso4WLNyNUsCCRHGD3ui+SPuMW2SJ91x/ttf9/B
g91AKU2YwQ5mO+JW0JluDcZtyVUW7ucJePpsP/YIRf8GRwLXRDU6XZMNyXLEysQk
EIwovXmTae55KWdll01UFE9VcuhXO87LAUnTFQzTpCvuqKkGEI6MQFf99OtC3Ht+
bSu6AuVamBx6gEbpzA9E83Yakdz3N/WwXE5SzDZoEBkVeVzWslw5tXkM++0ye/OC
W41FJSZwtsNx/qCuWr/9n1jVx5CkJ+KRZ0MOebe9POycteI3Wdm67HgQDcY9UCfz
D5bLyX/1emgriiSm9yRn0Z0dC079mixta1MY5NvdK46zP0Q+tOsicqOodd/gHHq5
hJlEfEMnvnJK6F249KQLgJfXn/BjhycaHbvcDdSHZrhPGb04GVFpeue/g15hznzx
QUV5Plz2+34kVMPkzFZVAQxfTDWsxL6d2CtuSk9rQIPLW8shpnPFsKhEN2wcriR9
RiN5HueUAs2i+M3TEXyh+14Gmp120CMV+6c/jdhdWbFswi/PV89xnOq3ndOr+mP4
I2mrsKEk9dEZUsNIMAcPWjSyssPfcd41W6z9Ls2fRoUm9lrqNDJQOJowuhkcX/wy
2AFJpqBjfQOmB/2kkVtrWlN0LKwdtR3ByXtPBlcNKo5HtxYGSHt1XxkSn4AwiCTb
YcqmCNJoiwjBfxD+TS7emMOZHzqb65LeynwYYPTgkKLs+Mo39cF5s2LUgOJZ0s43
OXqLspC4ZNi8VNtA4ANuAV8WhWXkiaBV6WjGJms3h8cOsvZl67O95vhVx28xQ6ex
AgjyTeXycn/NbV9yf5hGyLk0oeskUP7COQP/cizjcUUlTt9L8f6AU1eo1S/SKNck
rXddZYXajni8+4C3tQNm9rdHT4V/+Zk0qv02fYUHNw9dmNbNP0Q1nUBu0xpFGnZ7
K5uf0B6q9pEBzaWe3iuE6OPzcJWdJd9nj1Kim18+Z/23MVs2PB4h2J9ifmRwuMFM
aD+kKRGO1oecEi9g6XaFPjY4hQ2X42B+EmiollIrikBXEhV37w8RtLMefOdyq4gU
kkYiWsy9ndkCuuotRNYIUAyiR3tw0MO6StiC/5sez2C5v/Ns5fnwcajdrzpQ/6jG
v8v9BFkoBZb2NdoA7Bxn1fvQp6Q7P6YXM+1iI5lt/WW6G9df+aLIJjeiXHFhZYYc
tNLYwTvMtXuGrHrBZlA5nrbJcJcUIpjpZ7unejowvrrwrnmHCDJI10ZHzKG2ms8u
wMrsAfmitwAjkTns8e5dkpS0mMbloJwGcoQB4jDAfkvgp9RvFunYRgVydnBX8LwY
dGONSp85xi/QkxGUkD8zRO1lIBgpW5HDby7HluXu8CzwZK7ruhVlU/v46Nu9bDVU
LsGYyEjvqCXFK0JA0AxHgQV1W7RpmZWhjesEk5CXKC5SMNilwDp+6dhGEHi2E+8W
ltfSdovqyKirFenO1MTdfueoR7IHbAt/rv81oc/LX7iE95ediOO8JsmQmXEKNrcz
MYUe5QyKwhJtrOk3V6ycJLL4rYEsI2le+uBWmHA+/kmhHe0TJXueG5L2Rwxkuc/G
V+fBAyVly15RpkuNC77CLHuecjLxh1e9XcUo492semVu3lANr1j5uNPMKCTXUKjm
/PQFKhjPTcDaJUoOFXuo9WSlGXNmhT32RWGd/sS6hGJ5MMkhu2CpSCI7E7oZJ9tu
Axvmo2YxHOHupaMDX4x6XRtkRZ6w3lUdDHh1RezUFLucgwpg3fECgxUTJjGrgI79
tgXQDASivl1DlLsHgFyUVxVy55G2T28tnnRnNufZbdrwQ1iGK/PIXF8d6mN8LsMX
CIYQR+cmRJfiy2DrEeHSrQQ7R2KJn/aKyBGK+QGiSdn7ujOgfH/kW/n6+sojoKmu
u/i55ti+msDuJnCdFz9YvpBb85vpt37MiUfxI7kiR9gYEaRcY+aoHWLXUaX2Cqbx
epYiwiETNriHJn+faUjPcb7GV2b1s69lzO9gQOXVi7fsOFU7VMttrVDaLQrxbv2r
UK0Qc9tf4o04UQRNHy4ZYEl86Hlc/tUBEZNEtU3uxM6aNqOgAGq+pY0KUeUW2DFk
J3ZRgLTzx0faVe6Ex35lJkt4kW2MlN5jE3bE+iP5tOO8NVM4D/RNsbH1hDCm4d0Y
khpch972yx0+G4X4EWuwFeauTfGHqQZddSCVNJ6QhwPiDPtr7yt7i2xNZ8X3RE2c
KgMnstLf2USFFoIRVr0mN6+TVvUf8phrpGh3YSj+6Btkwv5NNTTbsaVVuzie2KiA
fnVuFKI4xbPyV1cDuOd1IqdDZffsq70mnmrZ8gOQA/8BCoJEkaQCctQVBesB0B0P
dL9vfxsU/+FEVrx0Tmsd7i3UXSYjiecX277d3dYRZrRhrmzBjy5W1/L6GkuFzk7M
pLS76vjxNGxNYfOL2eVKyEnNKtCWtvoda6iWE3DqatcYzgzTpt7adyUe1R+I8Udt
vxzrAHfo6370a3x1/AhAU9QQldvI0hfX2/xpzNVHpdZbp5HHJtaGxKX6AQtcAS+E
q9DZDLjwe741NIoae1suWO6/1vvp5ZgMxccHwZeSX58RF7SPw3PaF7zmrzbfRhCv
qyfJVMpdsbyvWpSOXoNDxFuggNonX35Vv27lPs8hF0RyrmSGBGXp7zV8ENZCeMfb
fL9r/G4PBCjXATpZ/gd3Ig0Zd0lvZdWnk9GbB1qE0vcWt9cke/4WgC0wOFCYFlc1
6eUcRGorBuL7f9TlKajWH0Rfk+DVv6hjJup5APehevmNdWZpr8Y4WfN29fM9w52H
1pWmiLOplHrN6hpOoo+UKCUeK+1jvM0FTMBZ0MAd2G7NIbwynjJXmLs2c4eUksgP
Z/7d6B01fSb6M4E+1QBlazfJo+uZEUoGU/zEgedYI4jmggYbjRV3zCXrrCp81YxA
WJceMemGFR8/emMQUVOv2RYhdjjz4X2IwEMcQNyA7szFlPcIwpnnWxKmkFsbxPov
nLJSXTgmr0uPUGSM6c1bhsZMCfPoyd3oB2Wid4n0J4GNoousiqSllPSUFWQA3Qpl
OoAv/6xT6zDBl0EFjj1H7QFaTNUcKGS3n3Bdalx7duCvXhPncFtLfCJLqbbWQ0UP
bcLuI2hFLHXXKeOZ1S7fw5Q2RG+eON4SMgUw5iZ4d1ywhiAXDP7bnLFd7K3+jG4q
hmGNi/of5CwPB2RnvIPnZsp85E1kMctKFTIRq/04tpkV3K3VERV1bTV0O3eGwps2
ZIpRPqQyu95T670RyErCaXWKICf55xLiBLSOHavw/56F555qyAYl+Po02HjEyJuT
zs4BrlVyW+LmgCsLoVRV/viR8RlWVGyt7XITcgpfvfHhovB9McX0I2pMM3dSsBlM
9Hjj9lhJyZuhDZ2rfGGyE0pts1/jEGTGqx01lA4CDTCbU+PHy9UeOB7HT+UB503u
lWwSjwIBh8VZALRVw0FmaWzrv35QrzLeBZpl/Za7YvQTYAn9hjutNsoA5z0ITE9k
iumI7H3pa6H6Gh5JEqPytzhjdUMjtjZDm6LdgvoSqcWe3irSkVsnJvcLuXPqTA6d
s9NlZeNlzL1jDcnGDpCNxbyjZkYPXLHyVqNrZKefRcDuepJI4N0utvf+2SVQeoeF
qawb9Wuqtce5R55N3ifBnk5AY2AKoe3DtzybPeDc+V0Os2vMTZgFjHqx+VpQicdp
0mn4OIUtPzCtd87P8HrXq2Zzj5PZ0s0wcsPrNpyDLZlMkpv8+sQ4Ccizf7w7pBTe
zqm1TAAzACTe1kDW/rd/nfrK67VB6IiRMUqB1PUasxcgroLq8E3RUmnimV4qyJmR
WV9qis388/FcZ03NoN/VeP/Whd4c4gDDXDnNDsEyY2Vg4jcIUbcvRJRzNKeNoNNm
rLn4oJm9hg0eIBsCMKcm7/ek+X4EJinWtYxbOxbmLUIVfNfz83SggKie2gP/HSg8
/vEPjjrSKKNSYC2sVnqZOkKRIARcB0X8PipCo5niQVlg8id5T5VPfMhaXE2HdB7v
hCL+UNzUVnoayN7QInKO0GNR9zwP2iD9+/LGa0DxvSjk/hUn3Hf+DtLDvIvznuTs
hVPBIXWXUoFhEJ5OkfuZTd0NRQc3l4GFsb9qx3qpYc2h6Ooajh1RJhnebk/ts2fZ
TDRfHSfuGHMRaKjnHlZKhGUbgPLTH14SdvJTHw4yaoM8QwNuNN4buKG+TWTWt+fa
UccJv5dpxsIh9QPd4DeyAapiQrYxH3W5e/wwY7Yi0G65Ngv+QvYEnNhDIZeTAEZ+
+h3WKUxsM+YEfk2/kWZ4TY7P6Iyk9cIGfN52l2WClozP8+DLsPgUEHl6UB8JGQas
RxdzBv1nNG6ynrX0S3jl9axU2/Cj3yU9tpAsQoXL+BpPrnrV13MBzbKLQ2fkzeND
I2fMIL8G2NRsCWGfqSP0xWXP8+oaEU8GvqPmfrRj5tbug4pSWbT5daEubL8sgy6m
SNBaxsYoJ39qgNdbTXG1Z391GexZq3+MHulIcSSaYZ9+7uQOENfwz8pIxSQhisf8
CXsVAmvnpF4cknpwf8JPzR/pFIYSXLdtnVVS3Sf1825VO1/nilaGyLP12eo05e/2
LOILdL3y/sJJecTJla+8xB3DWcSoK1k5Xj7huyC21/5N1Z3sbwNjw9jbPW/jLmx/
FlxJ5nJT2Z8a6gHw7mSZG9Goo/BL8HgF4y7Y8em3XllUuL9dT9bINGcoMQ2J1rZX
WLWJoi3zxGck5yHPl2ZLfX+uTyywdinm0rqZ/BkDdo7Lhiao4ZoTtDcgpZ/PZcpx
1eu9v6kfysgZPh3mKWhKCpAgXzHXp6YQs6wckef38uAv/7K45z8HwIWKU8MuHBxt
jErDsdxGMQ5o3uDQhju7J9ToIO16yUJsmMs8wa+fwSnn2rqo7iqszwHYNhpFto6b
u8J9eIDyCIecnacx6YLrEvhUTWYkhDtPOwCOYIzLDCwIQ9EU1J/Me1nAckCdVuRe
Mvrert7n3Oe5YKEXO1PL2uz9v/LiZAJc2K96IlJe6Wz3Lvx+UXc0DmgUu8Vtj9gb
k0x396qeEb6TGQXDee57yme7VJzIUHATtvxX/DCQOJKhAI83w5Yf1XmYoADZIHsA
ACz9g80nPiJJdgmxoOgxC89cAm0+oo4j6LHdMhFlAdxxmpkEGx46JbE9YE/ODxR1
gdZL7HL2HnxbMGF+C9prw3PDo9H43qQsTKr7j+GxR/Mv1li/4008+YNBxeRSfKsy
gAooEb2oC/4kbpPYonyBVEtV+vPQTMZIKBJDvkKG7sAOkIbtALNtwV4ITyg21FoB
LfMNkJh//NEMloycjTYFPUIN4demsG3zYDuASmFW7MbuzHwTzzEOtOBFrf3JvQq9
8GswVRDM7evh/7tOuRrM4NDDwGUjHIQRSl21mFdHQhlRuiUDCO/caAFvzGGvIwS6
7JeaYcJfiO5kodSwQRns+RQnH3UqOffd7kORaZkFsETj+SendItQHBOR9Ep8ZBAb
P2D5cQPAGykE9voBm+aZFe00BMhF9uLB9XRlJuw5W4zqrh1uVPlPOBRnjNlkROrv
WphMQFBhQlXvdL4eSbb1QcYoZE47ZUe+VCCfyqvWJT4keP++19XAb0USY3nTdCVF
GqZUzxoerfM2xtk365IsjkSvb46uRRCoTwmHxwqsQc5FBNqB1euaa8HZEVFNfTRr
sv4Op84WFVJHGE70Mg8+iXDOST/F0ddm4vmD10dvhQrYO9CsXtgGO6EPP5eYLzl+
nvNZtbOHzAH1Jcxmk4/HVZ82YpsPxsu40X1wHqENvIevbupdCuf+F+YA+u7L0ri4
a12ZKO5gjXj7ujGcAHLIktbzuCHmkr0IILIf7K1FDNwhhT/ywmOmI6ufrRkeqBoJ
Rbv+4z38av6fjA3KK3hW6qEo9aXfK4G2Y3IjLJukrMTMpukm4qRMJ0FXLlRD1apn
CdCQ/mFIW6HF8NP3gpV3+TOjkH8za9tBF41b9QTVWQOSwcJb9s1vHvHtccRsvMTe
GeZxLLx5DJ4bahtqfjtjBdJPvtEjDTYFV6/nUfA2E27dDQELKNqr5PpgRow3Ztb3
ir15M2zpHdJmCvKUZm+Om5OmdzjcV7+hbVzuefQ4K+NnRoFYWv+tf/hDahqE18bu
7z4h6DwaLI/Pj1cwYYqlufIecnFuQrILUq/4lbp8g1amcWC8D6ywOnhqVEONDRfc
3ABOCL0Jetue48keKNA7C4f2tcdsKRRgWOiqn2YHNl2WieBIYkvMWdF2PJUfGVag
sZR2Z/KLp0tl3SAdPYmIrQhHBkegKo0VAt/UcsNuu0bd5Ow2453U2MTJlYEoyJ6u
AQ4Blp6AErfACUtRwwpS4d2w8D7YD6VoubhCrOV8mT+W4BDCSnBXFQsJre3IC8b5
coQf8mixoqCdVHaEUTdZW8zcPkz8GkYSOvJfpp8OI09SkdEqhWvO39vW6X2b9NqZ
PGxtozPWHoej01WQhRrcAH5fV0LexnDPdltSj+lLVYgXOMap5lD2UeYoyTv2XHw2
SayZoMgQuX2sE3Qxlg40cky74VF8Vx4SPlN/9BMPEnnXS3iKN23kttT8rEElIr1Z
/SRHuB7iNzrMzuZPRx0Qb15CbSb0fwAQB+7FPCyQvCiQBigfSVQP3qeKscS1R4Cp
dTtgsCBT1zqgJxfESYmErFXvsDQZ2hozMrZeKHBN01TRoUx1plUN20px9lMWs426
myJHw2QhF1uz4xLOMpXAE1HuCxnGtBPrVbnYOGauoIhyOtsOUHOKOexIYgmTwHye
3ghPEpe+H8EP2UuOsQiQwTXHZ5ApHNVXrUZJqdC2SjPWce+5OqVSmAw92iO/jorl
DMkRkGCUxbDE0WjxTJ3ywMlcQ3+hofo71ZW+Q0F8nnzFRIc6K6kmGSJZz+3bC8b1
WOehNdtAQ2RY5DcCzMz0XbnsesDN020J4Mhf3/6Wn2cXBiUffp0sqp3F7NnikIFB
hPKczV8Bhi5aU2dMCs9AtHasa6T6qqX8zceW3kAe9CBwC52Dqvl8cU/ugw2Yd+kt
4iTAMiwrFU4Ga/vjm4XJslS/h3CvA4ZpSythStZGa2I8QEO4wFIzjmvc8fR2I2oY
Rtw61JlZnV9Jn6z5Kg1jAyjAU7i4e2kjXkkmiMjXJx5KFDzCgNGexiP80UXc1fdv
bdlLnpBAuwgsQoGF1cTFV81oPDPytVBQ+2GwagPnHPFdlXxU8AoSx0XEkREorfyj
opVpOEBSVuMnpdiy2q5Wp0/296yAO37sB8Gdrub+JZVPyjnBcNKmD/3aAwjfWPL/
AL3iWChjS5UcWBvzPaEiLq92c1ISDIqYOkzkoRVqRST33NjomHWadpYnLaHIcj0g
5whAx6u4c8PZuaTAaDJqa4x/pb3et+r+NeXnzK1C8Y3E4CFD6RUEVZeuQ/rdMvLV
qZ/dF6qx+dASh3ozNjkkrljuscWQi2SNaVpcDy6Cu3vNGNcuwQ4ZtsluhlzGKqWb
JK/k+Z3S1CZ2uMZYyq94zw/tekacFPGdx+qtUULhtzmj+1ac5RxdtXPAUhyCrzqs
IYejpISgszyHVjmsCSVt4PV58B4+p3XjWo2ZFp0E5wocKf5yFuu/Q+S/dLZg/Slc
B7m4tWYWVNicWUaewJREyZbJ8+BUMqeYgaS67ZzepP2FSIj+pd/YX1iD6knTfat3
CVTMMNMRqZngYY3Yz8mOlA4Bm8O+1MtOjoaVpru7GP9W6Coy3Jo9idH1FA0QqKfp
CK2oxH4XxIsto6O7+1f5VPZcOVXCX5F41s451Rthq2H30Zcd6fkCYRYB03BO4WVM
GHFItsqQ6Z8P+SusbXTAqZMNZCV0pjfZnIwLCejiLBjIQnvyb7ZksyDaXPZvMQRe
dlMemy51ni/u9orycVZZg71D0XoxQ3sai1aw8krgZUHzqYivpHrZzpRlxlTil0js
y7Ah2gtcINpAY/Bn5cOGw24Aqe2VasAtzRFrMjQq0z3hsBjM283OxijjrrNbI31Z
58rj5J0xhaY4bEWbTXYZditMmDGK+GrrCizaGptIAsfutqsAqdL7PIaArM48bRde
57ARNoqcB0dpksrC3JCOYOrAHrpJX1O6iplS1h2x3RWCTuLS30tsrwKSlNC1bhFd
bvhLsOganR5i70oiwIWbgdwdxQFRdxg0TFgX9gwv0MD61qyL72xVvTermbOrRrrG
OXwWVnf1DNhVJfRGTsD/KeMstDfM3t39Sa3XbR1h/cxv7bIObtQISkGN8zt3GYgQ
h+DHG5Y2fKXC4x0yMksOO649ZE6AiyYc4Dh+dwG30/3eewNG2RclaGslPw8WiuLa
aLSTTaVpdNjLjh0zTPrTBlOjnWGdPfrIJC8aNN+m5lTuWxMU1FswCI26N+WEk3Rd
h/N/alQ45u6WB1ztntwdL+RLc6tPwsIIrlE5HqUCyPLAD/S0fWqOx82EtVT+cIJH
choJwRsKrDCFwuRIARGKKBKZ5ht4LEEK03jwDhFm9XsD3XnvL1kWQHHQKnBxN32O
Hg+J5IoWNP7AR/xG3BimKcizf5CwxchfF5wGGQ/QV6umrPWyIxNiruTjKxn4XN3o
kaigKLg5cqd6OANOUYwyIQhZL+QPcpkxpYXvOViWH95IeG/m+G5vqe8pbSKPmvq9
J+s1+uF0WFwCckd5OBCCecBpJRXoqDM6u877jlgOeyezVrISMe3UtsZj1D3pGG/9
W0PMXSKpDsfokVq92H4sqPuMO+clbAS3GZhDiD/+hk2GBaEkxYTUYe0BJPlx5YWj
Ueo7pQBQiAutyTYN/oRbBgsRmESEkxlU9XVTFT731q2rxY77CsW358D0R991jixW
WADzPbqEx+famaTZF9CCogr7CxTkjnvYIe8B/ImXXm05Qwcy2ZXdzJl/3jPwS6UM
6WwE48bbFOx8d+lEV6mVaxto53L/qBp2jta+I2sEnvoY046TQ2y8mycCqZZ+96+N
Pr50zLwQEb/gMpwqA6lhNAtLe3SkP0n8MNBMjM6gCenJF8O/rZvtJg9xwYEHjB1B
pUDU4grw5VXZjiH//94Ll15nEiBvcK4HIr5Jp39oyH8o+YME0ZkQL+dDNOZkkRMr
+qg1AqUcF5SgFiP4TThmuF0/iKoQJFW91G2k0qURZlGgfg+jZDMpMmhi1ijw8zjy
oT1CS9PjL2UsAQX0T8iZIkqb2dxV+VatnhanxlbmFRirSb6MR/q/1qI5s8RtRKwu
jwVXgSbOaqgGEUeQJeWHXkmOpkyMKFw/E5D7X2NfvA3UvtJuApLoQkmQdP3LNXU1
KtBqNyCnU8uzG54ZjtzCjBAH1xoUCe97SXPAK5l3lJ/opqIcD2GZnXRI6fZzgBbo
9/M5ri10HxmUp0oJ6jEHFECLI9KMG6Jjmv2/JAQv3pJ77INi5z3nApAlZEIlodtS
kQ6L0DTrlcYhMKcGtSnvqcH4IzCT4oAd9ODSICNQ/CKNNTjNCQitf8lhOwrQr6Lj
kUyBRIGskgvnKqa8Ywl9oE1UTOrGNivG9i6P5ZiHHshhTsp4rphA3N1YoMVr3Pj1
QeZLGEvp8H36rLOW+P8Nz63OV9qyE76IUPhObvatb8HEos3n/tXSM+OnoyNu3u90
mHmxoabjFH1G1Vz0C+g12ZNWlnBTh32FZnlVbpwJQi+YIIvktPQrjz4cUTIq/e0+
9M8rWcyq3L0VL+29O373symzCQ4nhWBdTujZrJ978vWGE5WwSlMwUN0nARZpR8lX
sypQHSZ72B0OjcyjUkdzI58aNzI/kgGgEbIYyN6VQOH5ZDAwlHy8B5SYtm3O2KkC
Ax1Oxor9u4bJusvaMtn76B8SfcFTYYh/ZIU21UXfrpHG74Mh6hBxDjh/Wdqcyxtf
YzofUOd/wVM4/jvP7epRY0IlCpCZNmejroGhDWJ8wX9IE5XI7qlHw92LYfeKIBqt
s9uSvro/taZXlTSoop+S0Yj3TMkDc5x1fdl5lVgZ2Wn3xySFWsPpCktkYkAZzd31
pOYpYRGHbLkHLmrojtaFQD2nj/jD8a6l+7ZF7bOcW9GpMOLEf3+ijNavCunNo69m
6FfFgf4iEHtLbVCeZTqt48p4FSHc2Ws4O6LOdJeGdsvoP56wlxUxYWMe0d8JLLwk
DUnUEf8yVrgbXRmNcE9rEiaQBaqn8222uMUNnaCvQ6p+JXYmsU1moBRL89igT4a/
icxFymrezJ1CIzvI+a8uHTTzqixmOf4WZ0zHgBsVYFXLiYa4OMnSvRBqIUNPFW+Z
ubkoU+t0fyY7+CpN0f+CSoV2QtDpz2RZf2+7iqCkhCo8NrR7D/kyYaFXUKE3W+8c
GHi1GAZOgxWl5HNWEHNGmgyzB1j0N9n3k4Vh9b7+E5vJAtV2U4X9UJmeQt36Er8B
SH6lR7J5/DU0Qqf9HrJVZQiG8YCCdYz1J/AjZAYskpO89yZIzrCJ6vtlEJOp0veg
AuodQDdn8d0+Z0nYW86gi1Q8j+kRY+crR4u/SISK69vrGafS0ov+xLUUFFDaM7AQ
edoPout2UCn+LqPTLO/Nj5AFBuT6ki+RoO14GgdS226oAKHtg20hLnQii2thKzxn
ukOqLbIi0k36QVFjYeWAOREklSpnVe8rNnaWSIvSAwLbnpV7jS9QPqEexNhuGp48
Ne3SjPZHyLM7j2byLmOOuClRk2zrpp3/oOTibaMV0ZpAHXfEoNg83yFCKmKLsY6/
liN2YffSzQrdgzGglMwNGp/mlru39mqsacIWcuTyhzoNafYMQ0clleFoLp79bz9G
5m0YDJJkWoZFnGFhHsSthsi+S8TdFEnc/oc9f1i725TDLqDkNs2AUqRdZ0kqHvy3
KHvVFIi2VksRSUHqvHtIsQcQJoCzfoA58++2bcuSkpQPi82rAT+o8J+BdHu7UKEy
vmHTMDER+VAHnMPhHR9X3A5qArbVBkwt61rptI1j0RLOFgeZTTWgUvALYLyxwD8C
q44HsKFszWNfOAcllvx3TSquByFJ09y3ZzbPjtcVPtGqz6Ljf/Cb/XHiqUe4nNPR
W2fSjRtaSU+/VNZvuppLo6zgKwUJqV2TdW1qFDxlBE2yACuX9IPV8PJITO+D1fJw
vfzmANiCGNmIXVC1A1gyEa+pwzho76jBPQtpU2P1HEoIEfdgNHvLskQ7QGmFdCQP
hRxoGAchFWa04+ZI2WyX+Vw4LEJ/Oz1bDLK8XjUr7dpwTDvHaKOL/tkb2aanqsIf
fowuoxT+Pugqsb0HcigCtHB/utiUGWpxMJwTMFRUeQdEsJ7EJqN7Yrx/HOPMwwQW
Z9uQwjlRGjXk1j5HIQE6bWZfphAwxmTd/IZy+uVUfEbwA6jp9uuD3T+PolyctpXI
4xfMSRsfzJPxl3SDim+emT5H5vHBhYTiRuGuFNwX8EjeVWnBpUOvKzaVUn+aYVSo
LosOrbos4M5sr+xFAgPWb1fQO878ZqI5/4DYB5nfNQOUpKGR38EIdQwgGpmPjQEK
/jYreCQjN3lE6hnoDbpmHj7OF/9c4l8WEPo47p9KWqtIgSefTr5Zhdux+q2Ef1Un
UirVz7SJ06psHe5VPEL4jjbxHPloCXa+3FufIyTp5Th0oXK/dbkv64pTn90lS+AG
9F4hxJhJc0LnTu/S/ORyLclZa7ryAvE9/4IiuBiEM9nZxd/bHxYseAYNruRDWHF3
Fj2InhGj5kxB5dGd9BThZ4o/9lRVNIZOYhdvVcx6Q32wWcF4SzE5pzHzURUtCUE3
UQxQDXD5v70Ca03D2L3AQ/h3qB8qkAzUYVAt6hWyvuSIN03WjQg/KgvHcNeY0eOF
wbsROfaYsb9g8ghQzsHNZCPmmfeBF8nOAEf2gP9JSBwjJNMULah2okrtOg+zkeJr
f1TFh+8x4oYaqIN7JE3Va18+Spo8Oh7RolUALQCdqM51LY0tOcr9Wnu/d4/HLUn3
6Nhp1yLfJCPWSn0MCxrCd2ynyY2HyvgOctdmJKKlBe7B3agFRgikhSKQZ+J17F5z
75hxs8PD64LvdH7ZeWwj2o6xjjm1xQ+iLlovK5CRRtosP+JvFBjK4j7kcckdfkBC
TeQhzt0MBDNpa/PaMFpTXcY8f7+z6bkt8bMLfUeIP3u7CYaCHTLnorEUgIsQRyXH
GLL5STU9NaB1rRANZdA3HWIIzhbazh30sPD0hv9suIQF2vxh8azV2YhMi2FCRyNh
DzQjy7TG2DQqVDtdtP4qj817ROEECSNOsgGXpNwD7YH2OGCw1Qik0n1G8D4ZVFcS
ubQlel1oyHqITakN5+ZqRFPLADkJhqRx4/aahMkJMyNfrEVoZjwmixeITL5KdlaL
lgtvGJnYwIUKRcf4EZldLRfc6ni0SJBEAKA6EI5vqiPFEe1cXn+eMZb3kOYffkt1
ntiLzuBdmr3qdtdkiZTfpfWtc76O86grzPrXM11WOFjVtOna5frD6ZnM8MmsV+S7
47eixFXw8GyvhaMmgMxFPiB/ksfzeNNE3AC6azDLAZpffm6p0kK5c/KcmKGb/FSu
pnOXBtnJhV+8hQsi9nQOk3WP5ZVqn0A90OnXmAfbxLcUDJ4bklRmBrUf8V1dgZdq
K4WeHYLMkIyPbQPHu/c3GWCoZLu3dy96/wbdU4hs0YvR1a2xkgf+II3K4OkFgQv8
CSrmZlU9kZgaGIJwi0fvivLw9T8nETEuArewEBdA5Dbx1dTGHb7iJPcbtp1kZT52
eFc7U5SPNd0S0nN44CFvL8L2H0sqMD33C/dnxRP5YwsxlnS9btwap84ZfxLRlTaD
g7oHUlPu9xVM/MeTKyb/XZyTQNdCSBbXo4onoWuF2LdIhkU+sC6MNTYsPhvVdDlE
Lhw1XrU42HjiN5XBIhwMyz5nB9phSAkDZPmgJQme2s2iVEDHpoRaWxrCw+J9U1Fd
GV9hYE5rEvv5G6N/DfPx4CrlSSBUM9+AEq+KGFC1yFHRChdlArU1mqhBpGC6t9Ol
LHCdtPK2ltQvGeUoSdhqztI7G5eOv0n6uV+vn24qlzegolwvbB1aIIVTH5AsV84l
2dD2Zt+JczLUFo2Q4Zy0An+ljPpWiore/OpoAw7T88cOGq2uQcMs16dvnxtCBaBi
Gw8o/Ei7kHScNxOlPGL22dxuPDdRy5Sxq5eVJf3PWwHi+T4NOswLJIR5gNweDt0A
kCBLwezboq+uTf9DA2RQeE4Hbm8P4fy/lKfqMXpzDz+WvYdbMFl9wi/DXh8dAPNG
4+qA8GVkaezEZFWc4Zu+40/cFIANhR3ehBb32FNm+mLY8D6x8BxxjtKEqPxIkDre
lw+Cysz7qZC+x0vLCJhbpV8inbhos9Z4V6fMJoaDJPxQiL/zXuxBuWMogAO1smcm
hqNW2W1XDlxgTnnpOsnKn44XwtqbjXTNJAnf6g/0XYUoGP629kVwkaJaLozMzPnM
wErJw9iRbvI61Ic1nJy5mMbts9j+VVuFvc+WYheddT0aZqI9uX//tkX8j3boWBwc
VmvQ7fw2/BNX81JTP7K4aKiwboi6TElzeErq0ByEVZAsOJw9JbodYty4oYLFE/D6
3QA/8bYFMcBulo9QN8L2gpPl64e4SwnB+Waj8VDAy3PQ3IdYH9noIIvRAJFrBAhQ
ZqJ1nqR/53hyM4DQr7XWhmTf4MMtbmAyLwr6O5/MXrrikMYmt7n0E8TmtyyKqBrh
Vt92GBJxss45K+giDLJNrqVTsnZkjHrJif7lLITLDWDbGvZa1GQL/ibmFq+XR2zn
wymtYxF5boCAxPoXv1Oppo6alz1P5KbzfSHhvhkC+1wQQM/GFlpY/IBJCYL6lHXC
enxz6epOtW5g7pWD2S9YRo7witSTyBjJN3221ACdrb2gaE4lDYSj3/Ao9OvGFRA+
fA/tP7KowmQ9M1maY2jXjSEvxdatjkebvrN9OOMHVhAhQOFEUoHQ/to36k6ofhK0
Khmob2nHDfRMdfeNJNpUzeH64piJjftHQNIluPCnuHIboEsax5ya7nbAVz+uMcKT
9thM2otc7hK644965boyMQhbdwlQKvIVtVoRRQlvhoUCHmizywHEIQc6gRP073Oc
BLw79l1tqq6ox/Vf442FsU1jqFf3mEOSF+vmcAPX5UvuYKRUGMd3Y3w7IAdPVtng
StCmtylZD0JtC5SXvqCDAqaMGNRJq7wj1NLgfc3bKL0ZzkQJePM0Tv1hClSNXwV/
iRj3itouJe4r+qdvcUfz260+Fz+FgaqVGewWXFSc7JBlavbxnsFwA1ABunWqpvaT
o5OTYL+AOcooCHY5SjGWGOzDLF0yZ8xFxo24VtyR02WvIV+I51yzaiGJ/eNYu7QF
5pGX5sLUaGEnNbWDTJGo+uvGmhmtcUZgGapPSE/9OmYtTDfW0E98HjyfvSZ2l7nD
aRilX1O5XVy2y8LHuWcHv8qGv4qh07DqGHcaquhLsHIzw5hi3gPM6p/ukbZmUObS
IejJt6F3bnK8lLIc5zu3x8tFq0PNX0AaB32wBObdFK/75kyBlyUm1mCZKpuTiRxX
A1zBZAm/WNKoqNKUYqJw6KP5WI2ekbivjJ/izvfnMNbjpgF2b93YnHPcWDzh1+Fm
y5/8Skw/gcEJ3pgCB4f1vwqFtDLeo/WPo9MCsw7ePnLLZocGGilpu1Ht17f0Kuyo
LqA65UQmq9cQGn2WgjSX7Jub1/pFHD3VexZIT49slJlWTM2DFF3nCaBm9vbWy20M
v/Cen7iNGEYyxjz+AqTN+z6BJViYkxfFj/FTQZ2wzUKG7xKGdReAr7Kxm3YAw9s0
fOKHjnWQ4VMdeYqxbTGcjlSn02yCMPPZv16tF1zDuS75yy+TEEHJF8i3JN8X+11d
WqCjzMtAlW941QM0Fv6dkbwSSkF7DKbQ6bJ5ACSr6tGNpWitZ8dVCXqqrpmcKBt+
vOxI6CUtxvJrRS6sdrC1Ok/HgYXiuROwPUhDpFvcDI/ejfVEO2J5arR09XLdG+Wn
drQd6Xw487ugSdyFcoJ/eRXbf7KVQQlcO0s1PWf0xX52ZYBUeubBqMyp/+NDhWsl
6yCywOlspGe+Akz4hgL0yrucM8H7kUb2SawujvruHZBMx/dojwpevO1aSTXEMXra
N4Q64UHWoWhp4CwO7T4HdIiDALcZF1ArKeVqGv8+RdPVwlAJe3PrR6uYY+SJOlD9
OtvaoGJ7QevwDjdYCMY4d5CrQoSFWmF2juTbgtdN5BFVjQnDlVg1e7djye91Uu+Y
BaYAyralpPuc4YR+C2H4HAzBBvRRTw0EIsOSwZFJ2jcne7Mvn/0bBgPINk/X4D/5
oqpgEnXT9YmqvrFICWU0EP3DbRjbtED16NxOUsMh+UdiF5yLQD450tAk74F8d3kS
36nIm93D/1rimKSsW/3aU+rOuZCVFX2TOq6YArM7HSeILbgs4J27xG+mhj1uJ3fc
AaXvfrfobkkJat5jz+o7bX3SLd660DITX/kDrvbMnMrzfDFszjYy3++FujUm/5j6
CI0BXPSQV57s1KXdUPthK5DthZ5BlMpGsmgFLqZ50UVY9bFfUQuYtYAC8RE9dCvs
D8z6YctMiq786aAFmE672qQYWWORCaScPho2iuoorR9MiAFui6zNYqfSMSjkh3Jr
4J8qjr/dcFIv2+gyAv0foR4ikPQQi2Jo8j94BuOx71kEtCk31duPDN0WnkFirc1d
QqLjlVOU7J8/3ogDi/DvtkskUK8EACRWt9Ochia3W4+yPzbTN1I7d7kvu+s7hWRl
fzanrUjy0OisC/0h0nLCq6KaZBOHJ/k8hTtbLDbhp5cy5X+/ei4juHJhVjEB5CWW
GMp6Et5DHWEbw8HyTg0ethyMLXdVKYi3tUiUGIf2887UUOtSYA64uB4D6vrSJb5n
+jN4JRv8EpBOcnJLXDmDuItzFFHDvUwslbVfP4FXbBR582LxH6xM3g2nEnH23nCU
ZhEykXSARyEZzioACYrSWFeod4/skKFUZun6eE4HCzBfzrDVeZgonb/0ZhDamMOq
gFD9JN7Lbj7y9aZRy3sUMUCvx19dDPDZXRc1G7g+3XrujWmkQYVtiRmfWsChqZQW
HaTfES1OFY7BIe9i3Gss3iAlvQdRLJEahTABG8fLXdzZJf6L899sH4KIWp3vdLMy
p/eVcAVuyfW4wBTuQvSSV7iaZcpZaK5Rqpw3+OqtXrMfyFSEifF3OPmzZdCNsv0H
6065mhNDC/iOlDrSsXzKkBUAA9ABG4aJAMoreCOSAGOSn2FnNecurR7rSPatWnqv
CVvprJey8QBo16ubH/nGvw1F/8sChmrzOIR44AqqbFnAB4+vhDXu8a4nGSwSpWBr
xUTNqY32JaWjLcVJBxbVnUgAzn5Rr89DMIWUA0yqgUPrSUDXLn1mvMvGKacRIeH2
54+UbqBge7Fd3x09RWtXhdiFvhbK27IZed8DqqJdgRU3NNRhPaWmfm7oCEqTaoLh
fu+ivlWsuZ1jFr4O+jBBFdysfizAWe4qhSVlLOYedIVKB/0y2KNsk1FPiKjzkegy
P8F4Iu241qff3uYMdQ2miyByHwk/erNIbrIsej+pZzZebpEOyQw6Oa1lprmehcMQ
d07knuJdLgPzBk9ufwiaulGn+O6RtOc7T+KpLnNnfNPN5hWZ1ywAMptPm96Ix2Hr
hHT3SF6WtQOLx++zYe00BLT/HLjQwadu2syq6AccWBZcea9dqO8KJ8jBnZHZdcoN
K2pQcW7EhREyv4fLMs4lbWcWrvSn+u9y3McgweOLrAkqgB48dDeKrmcKb8oQsE/3
VczVyEfYVH6iz9bQqCUK0IDZonFnUW/FoSa9qh7MWk+fubQdTmhZtncXv4BoFH3t
w6bmXy/vrrppYauFFFf50R0HgI9vQEISN7ltLX75hs63gha37syw/f1Bzwyd0TUj
2h3LMb4EmxU9yJci0ncJ25FyL452CESmkrzgSXr6nvApLKpWIkEtfikHTKZhXJyg
4eCuuvUYogwffqLfiqdwU9Fi/EukXF0hcpqTA33Cup3bcY6wMbZzc4NCStJFISvK
T76UuJUN87C/nq19QyEPqwpSAuhtIpLImJAkRLfzG1VW3Q6qyhl+8mSU1YdGzyro
SIvRwKAaMihwKKCBL0PSFMKVRdIAmVmFfoWCvOq+Pud7vDEhgShdjtuPd1wj1otm
uoLCy1RKelXtNQt2XT5vhCQF4AaNLwMFketaTJb1/koPFdBg871BTW4lfbabm4Nh
kss3zBU59vJADdTehkSnvqFRLeJbKiddymqSLhsxNaQjXi7jYlxOg0if/zcYDO1T
WcpMb84gf6xbGT4p6TVvMb3UyOIN9AXo/9tz2BHYAfhwgyfTw4R43HTZuHY1IiLV
hV7I6/m1h5VFtQ+J4oQeGNFsK4R4Aa/Cim/AwAUPI8DjFDEyPzKEU7rPhx9sBnKU
RsbePWjqepj9eAcHVPgMCIbtpspi9ttQFdxSae61ZbZ8xMx+1T0nXnmq90ysjjBl
jjlQlMXNYQwt9Ap5xVbfRcstMcSYFdtkZc8+0oVwpDRk+zSpdzmyHtgFrcVSntMV
1wuyXogQH44m4A1dRVWojWZB3lXfmL5G5/yc489xLLWuZT6xoTmC7y10filMZ209
KiP6AKHpAVS6qcUw8akMCH8K2iq/49ihI5hlzZrtsKcOwC7IIDhtHmHte17bFXhM
T4WJSazPPi/yJkooPTtkEhJY6+n6VdlRQ4vxYgiTVRS9nArKKnDYvOd3CrkNmulJ
VPOGyLYe6djEFeIMEQP0e02o6Z3ObnP1q2bhRyMo0wtwHZWWRt1xKmfZnhMT3xTC
mriOlSSkoh/PkalH5o5wV7fOq7ScXTCbyi/NJXBicEWsBa4vbOoSKmq6QtZemu76
5L7iZfQ5TJ+o2l7+Q35Kwd6FWnMNa9SfPibL09EDjnEWZ4SrKdSzz8clHIcwwmR1
3Z0viLbrC8hOZGYue/dPvsKbkeiPsZaSsMHAg/2rJuYMDVy2jOTOhQCO2RpctzE3
OXQ+SbuBpZ1W2T2KSOtF5x4njgdLMl2diTzDQeqfx8Ovo/170tpghHgVwr+pmyYQ
EV1S6ll1PhxncdqIq0JNEZyeLbTZrF5RO4GN5bgpZ0YtaFctEHmHW3I0vZMs6FeA
Jn5XCkYoFFw/qKX9NHjn9vqQ7ur20QbgjY5a47lUq5G30KzkLptUkjdDvTYgBPTo
+6ht5HGLCHqtL+mqgHyK8YESP8DheNyiTyUZSWxhWkvmKdRINzv6tCbheunQEk8b
H8i73wd9DI8Fa7qrEEOufrMR5cEG8YcCiHqSagj48l1ZOc1QopvdWovcaUYHozLC
6aTrDm9hg8pEIfB3dyUuA14x8qSD8fJCCg1pllDWMCZMa8EZSDgw3jB5crkBlMdB
3QES7aIX6DqVQzH8hQPxKUnJOr20HMHpwl9A+VhGTWHuJvrR3ZTfguUuGSM88x3z
opZiFZjeKjwwb42oq1Agas2/6xxVADNqdI6Cj+LeJ1bVo+rer2JymnbV0r4nh279
ZdPb224/iXMWdpDJAhrxwhQzxviFKYezNcxQNOcwCgRjNTxTRjA0Hf0blmIHuTwP
cuLcTfPScf+0NGG/7HnH4fBKbPupjT4Fdoge1Tm6B1yIlYN6LxO2yjiIvPlD/Tvg
fklAuCFtchsrYKnhy3B759TIjJNEThyCGbLk1GSshYwx140RdiAIw9vI3je+bRq7
JMvv6dlW88u0zSR1lWQCrokvdzX9SZ/DTBdfnzZImZt7Ujqmq5dcT03z4Vbx98Fn
p12l9KtMASM5BCUmdweOn2SPyKP0diGp9rOfVywD6KzqwtQWr5Ta6OBRgCu/aWF2
0Lm21QNHCbSOfmauEghDFzlDWv5AHMkkIg69pZLKDk9mLudXNqnZugPEsLquntJ3
/ze1lo80D/M6SN8NjRGZXDKIXrrGX/UY03dKONwa5DlBSwzbt7AusZhDLTwl90Xh
Ru+R44VXiNGQc/znn0fP5+nqE4Z1AHXTQJHiHFanUCc/c9MUUqhLk6w5M0aqTg2s
u6eqzVsBLFGxJI64RQlItetxq3tzT2pjff7uTX84XYjuIg68x/IFZoGXzc9OeV4x
Kp1mOGD7Dyz/SRXvbSX7q9ez6juvuuZrRbvtU8ovXt0U33yBsWRmrbJVg4bevR9V
MY285uXtR+Iv4NcYMgui0nbWXAtJ4frnuD7aE9MxY6LOJfU+wxNolxMfR3HHRgUs
NJE4qR6ek39aIQp3h3bPto9nAnEa6zQVDYWuQM0bcsQK87nVzfyrZnqCHvBBG0jt
7ngtlrmRt/BTQqs7cVGWqeiu8eeV6/Gsln67eCh/l1FJlGa0HfUP50B1SdthTfiM
8/ps3Vj8k+1xqVNhwOX3RF+ZIdy7jR2vkMA3I2TKC3N1O018g3igDiITYHbLt4rQ
OhlKVPCprroWS480l9SVo3dNx4yuiGpO2B52I1piYHtB8dJFqpJgkFvYj+GkiDGF
Y/Qe+iv9oZLxnTZHnnTPSVNq6G76YKgNmOA2ULjTcuZEbLIUhpIa67WjJR+1T+GA
jktoLwuNi0ENve0adt6RtNuu4cxR/M0BISlxXYXL+F9bDQp+SA+0Lji8PtyJV/jh
w3zKFI6dk/8GOQbL1CcpCKuiqEbyAzXk6ySCB0psFK2N6lc6eaWa6w/PbYm+ZaLx
78rgVbWowEE8hWKVSTY9Bawdxxp9rSQ043Era19h1YzTQIGrk/2gKaXWxAwSdr9P
8Ss7r62+5615WpBh2utWSLX7t0RjNzwVOorUY7b/dolq1dfVc174npwr2MfCLW3P
ppAAEV1pvzNbuIawCYDlwgB/MCQglFaTSyTKjaQyTLR/nqL00sFSS9zY3trgFpng
SV3lRfQ20+Zo6bb87dDmUXTrAhJXKJuXxMJwuAWlcQzJ1xb2L/0pyjx3yx+WdPdu
ZpNYvVyrdTuMtLLhGzd/A26VZUSU2E3Xr2manjFzuS/yn45iaTYvVXIwnltBz5ta
Gd1kDMW+lDJP7rn6hCelLmr/M3pzTpXeuVlgG/AW4NSrejp4eC1zwKjbsL75h5/S
QqNZsodvZt28I/mEaCqFT2ZyorREABCOYJmUxlDxTX70gkMvRp2QhPgI2sUAnOCD
+GvUFcKysJpMBsd+iq2eABP1hVSNnY44G+XHr5wt+FveLCdsn3xgfN4a1X79fj3h
8YFnyMHfAOsZXiOaZUXVdmq4kKzlMCD33Wny55haK17Xmob96iNCS8r7ywMvia3n
rnMDtUQdllxMgf4ngHaJ1R5GuG36dwA6BnDAjlOaIxscvpvVZ55TZrxRGO0vAio/
o54rIx1zWJhEB0uujF/PRadz4gEL2qn9zsdSYuCydObzqI12kbi8ln+jE5pnMSrH
OpZJ4Lxr6Qo9kruICPlQlgbKtWPIU651ohB2zK3omGqfEc2OwtDcIQDTv8U7Wwfm
juW3om6qRA2mNUOcu9piSGItlWjwiz3KSeeX8qWxl7jtvfEVUzTvBn06u7ID6IF4
sHJs1FO76CSRktkmXuWEpsvNNifXPkooMOZb9m3KzsVl/gyZAmWIROhNB2jHFpGD
LBFPGtDUybpp9Fqbxzv1R3i22Lgy+fVCOgXdLXbh1zzCKSx7ut6xl+E48DH3gQe5
Qqra57YeSGpwa8ym3WNkJxmuYFO6+C89u+y6VHQolVDmWPq0RQrGQ/uK4XAegA7J
Q0kgUVSk5Zaa+yuOaeyegYcYGz5BEhmPJMjWpiavr8/BLR3WO1cyOMrch0LHmaVr
AJ5c6BkOqzBx3Z5MFoi+/9Em5JYn7+3ixyQth1bfinSbLCbfxy2ay4lFgDTHvY5g
uy8G5tNhHQpXqAwA/gTregECe1bwdz9Kant+k76zC+ubeeeKxseq8k6L3mEwMZqg
AYO+7T4N/LevN21f88bsxQIqqCKiOVgI5UCbeIWV59ftqKKJ5tS858mkE1Xq2bQD
WSxtauwUkMAVHoFPUJTGwBA19dRGIxz90S4mrWRNMJPHoIp6NnAmZf4JSfAL2CFc
uSmICZMsYX3H3eCD9QNSwMMFaokH7gOaeTDJZCxzZ/oreTuOmgzuj/Q0B+QVQJPX
YYrP5LWyM7zuSpDdYsOjs3IQrWmASx+zHJNn4JOo2M/QaoZPvrVpBjYCESV8IZm0
qOcejKJ42LP6AWa9UI+yryXudJCGiDZn4sBc6h5lp5tKxv0bxmgRS9uMik/fhZAi
INoRG+vMdKzlATUhUYLL6pXPHj3wHKBqGwPFcOshFcd2bKUNc02fnZO1mUKhXENR
1Hl0Y9O41IbdSxpxuDZ26n4z5OR0gWLLYfjX9SeRjbTq5jHUnuimO3mcrhOWjMtf
12cwDzJdpL3dCvYBDlBYtQ/B3Rb4w8W0XtgSzzGA+1xBKhMmiI1MXBvZz0Q48JWj
FTtUC8qkB67AsPJ1YFAy/aZ/0Kkd8whk1q4+MBL9GWBp5bL63VObnW8m2h7gcUnE
sjLpw2r+QniYkM+6gMbSxk87ixE8jlx1pUf7M2kdYBVi0ksC8bjZFCSFB5doKJ6k
8mIakkl7+awP4d3xaJzcjqPFv1+P+yTigDC/70xEs2Dkl7PsTYuzZTuEeDGCW7yF
ik0cv7aXGOjhSYziwCdrMOqBui9U9AolRA05/5XR/HglCrSzxtm54ZWKEF1kZSp/
cU4S60oBctgPFmVPDVnCfR2/T95kGTcGT6kbIwv4/2UrV4iIsDp0SYM4mz+OzrNG
G/r4aZV+2eM9PIiLSv8aJaMqWiiMAhPqIs3rY/9CYbQSpxpL1W7t2hy6bXx9gyeh
IlH2Pz9AdWzbD4pa1WL6HRR3K48Zs2orlgdf3NeyIr5rkZm8NsIfLzcBY5sjAIRv
OHe3/JEC945wDGH7b/3zR+tmKqa9LkYN2O8OVpxrlMOyp862/75eQfQ4pjJtsV8t
Fec++r9kbpSXCfM2LEN3d0HPGyC4PVnx1TxVU6BacC1mTDgxxixO+XpS9gN5mhYL
fB/yfeMLAufPpe/WekyG4vfGYuGPAVdv4k2XBFdtVqVuNJNK+4T0b0MWGHNWKCD6
YiJWA1wuXhi6z6FyWA1NvD+fcOhhMnlxC5aU+08C0LDjrgu+1YbCKLKfWYEiw+ig
JmTymnX2e491cPE4zLIbIAh+lbz2y5+Iv1gOFNft09uguen3tCSLg43b9HXbbbTk
6iWCDUiedzHhJbtwnbLJDwtirtpF4/0YpPl8HNvyFsO23nMFzCA9M+p3c5ThUUCg
suTfwhavNuYeRe9J5d6tRAj4yBE0qmSFuu897OZ/yP78OjXaLwPQol9JDHbWxxOA
rU/JVPgLNNBSUOheEuqweV/HvtIWL0U7kRfl8kC4bFmynW7q+9kZdcC02s8DDjHJ
rgQbvemV5eN8Dj5/j4PQ9pHjPu5zWTJQjV/1AE15oETn5kecCiI2qICD2P2iwkcz
w0j0aqOjDAzelLl05zqeboWj6QUXwMlEVbkq1Nlyt2qZMwKOovnSlKkhOyriF1Kt
YRkxAHuXcN8PBFTqh67bRLFY6lE99AuIaIzjG01oDYs/1vdmE5gfojcBUM5IVoV/
BFXszq2eN5iSueWMPMlVx3E6X3tzKDyI4JSEb3oTyxk2v8QVyj94pbwuzSDIpqju
Y1tPZVxgAml9dD1qrr9KA/HZhoyfEeumNCJ0FxI0tVnqKF8fREyxm1mQrAYXOw9W
jOC/2Mx2Boco6ndGak3t0z11Q7LFYD7bdazxy21MaIdzUl6LYr+S6QBeSao9VsOt
f5NIYBCtpd5cO1KKdfb5oKufbT5VDVQR+cjcvndzxYboliWAmd6QX3O/ns0Kiefq
xU7iHTi1PKFkYNkLL6H12jxABwd4J5m5pe+6HuyWjflpoCf7ecC8YimRGRdaheqD
t0Xzae4fakIOTxLnX3HNzeReWW1UXpX6mIJdWtDJhVFdocQMWVpB2JGbQ8RKu3ZU
fKnAAqpI7Dh6usYdLi4tBM6gpo8DQ+GCo78Io0o8ktu1p0c3l8KToWXsUhIq+K+W
hzs1az6tYjUAEWayW1NVoW0/Y+18yjLxYChKBys/Sj++mJyEjO2IXoa/qkP1sGjp
AdyuHFv2q7MU1E2QXZNGp8bY0DQLjiDER8GvUpZnkCjEsvJ7PlS3wdS01vg8rul5
hn5eUmf9er7s6hQNW/AbQFCw6tllUZ/m1N4mX/xW16V04InIreIv5oV6SWGFkhqk
GUPdFtdvKjx1/yvOnvaI5m4A6f7hRM1E45/oIv2ut5kfJfxNDm8O9v6KpRYEFXxu
DbmAfzXvts3Oq05d8imonS1wW9ahn6vQkVDZo8E9LpInQokJSDrido/Ix1sFsfAw
T4z8hKZEZHXTu/BNjH8pQDj5v7L9HAKewyezy2JOaP+/msDSRoLSFV+cdj9FJf+3
waJ7WW2FoTCLOB6ncFeojakmYW+fD6FTyE58oVhaNMms6yuYsnkj5DKjXGtRa73F
sx8Zx+vY3PY44xc6dtojzBc+d2GbQRy3GdxvGUAlFEFWzMR7W92/OyJNF1+TDzqL
RX3L8E6fBVBPDLUkdYokU5wY/bPIajBZ2+ghgoZFCrKDR5vnEyWnPjEBosnNchRQ
Wq6ms9m/YON++VM87eOFX4GFbf500RQScJ5JoG3Urdd5T2o1sjwz8ZnF6JWtGw/i
SU0JhOO7xyivWV3FV73uidi3E3vgZE+qDgdq8HFn8tg+YVzp8PyS3OpswDSKfePd
lcJheJG9GJ3/8H1rsC1Y8Mre8Jy79oUHVNm07dSzefVcFE75IkQlCbUTIzbaV7DH
pi+4v3QhQVDlnOOcwYpNCLD7MTf6vgE/Fi4wU07CdtfhWrIoJ2+bQPjq7FQVoa/E
KtX2n6aoDahSzQ72JiGP9oBlwWgDWkC7ZTwT2I+k62ifuDVBNcd4sEUaiAwh1f7h
2UYmrmsDCjUwQDpiZWze97fWQ9R2WnVhpmxKiioncbxSveQAUpuzUPA0eJy/44Eq
BZaGprMA6eePOyCvDwXNSxG+RlUPQRUKtA0f8D+WXJiz5HKTwmi9Hk2EfjT0HB1R
U7+sBz5NRnUt3UgffvTFwWcx8R0/lCh1Bl5z6+ViUV8Q6yFRu157D+Xa3Q0N6Q/G
FD3OHYgBBtPFRxxFalCSXVBfOSIL7d4DHlClrfHoLBZomlxwLRRl4saGO+B1ONOM
Eq2t5v85W2GpHZuJK3Q9IYETFwUxAcBqlD1zFD9/tQbSAIWmkEXggPEVjQZQ1oQf
qhXJh+pI59AJVkRscEyGQqkjJZ6NAfihCkQ+V0bFtyfwdaaQIoLR/selzNYnrFgj
ZgRTJUrwI4s3Qz9I/QPJ1zI3fXqRrWkyx3tgDEZZfEhPcvakmZtKLiIqoBJ4UY96
rY+vbJKgc7WEqMsGtIkj1GD6D2s7RWilUuve0c3HkdFPJiHdDHh/vDS3HgUIErPa
B2+jMAM0bOqjyPOMNtoTpMc+cGzmOG4YL3dEin3yu2vlfsPgkQYWgas8i/VOGaba
cgAMRSR9HfYQxF8Ac9w5W6aOdj1/inD/DEpOT2atnKTGu+VG+rEj81VXxrQyjdW4
sQ8zKbqF2w6oz6kXrxxys9ah/e/OrqHQVotGuGi3dBkdGDw+NNtQCfqBLogxgu7s
Cr+UDOhTe8Z9bRB6XvRCULo7f2l8j9bcEqq/YkJL8mbcEO4nmFXvM2BY/dQSnLRK
Uh9lmkVTtkpG3ZTqm4rLxXp0zoDfXqEXDhYf72Rv72cmbLnS3YKNvBSnq34BpaJR
HuYexUqP0Fyn+Uj9CA1U3ubogbPzYSFdN5C7tJFh/Gx3BsFivE5dFbpYer8DfWoQ
z4VTv4bU4/A2uV1ppgfeHNlnU9YOcx8FQo+wpnddO1YTyrK2uThVXb8rw9Ca8VUT
CZSgN7s4qNT3tfsqXO7NipNC7ZMSxa3ktccaP3ynVRF7iP2r9MZSStbWCHBZn7fZ
EW2LwLmPudZYins2jpVHg6OP7hccaH1cv5SmNEtlW4BZUlfE231htKou2Y8Y4cV4
H+8Rqil4X0iBrmfA3Ui8QvOVrH62paMvvq08uMVAZ/Z+mKY8KSi9fuFIgavXtxzr
7b2dkfypNgo8M+lJKxUlGuB97d3/yDrxLBFLw5G8m04RMR9p2P8oDgYA0fNzZHN2
/RafJAf3aTve8TmbZGVNy5+vG5bIENqKN74zpZMKZWETn+HbDPfYroUQ6JP+hI3X
b0NaClBAKjGNdh/H7SAb9mSnrtvZLXgWbZQL3ddJDLVg44VZWhScJzs4PdcHi7Tg
sdAvhb54AXKTaajr3yvqs2B7Q+HKcmb9wQBE7ijOdv3uEdqkW+u0biMGafoqE4bo
L8h+BzqfMOirOlgXy8ZH/aJT+S8KBLZyVpIHCQIaNwSJisTzYKxhtkL0ilAksHla
gjOIH7FgqDGDc3HVwIoZlNT+i+v8o1lDaCJE9069oKRMBNvOw6kxmIpYB+9MskP9
wTmrc3WMknmUevsE8tDoJNC82uOMxKMRSSxhHHjUycUeT4SRDX8vJ48Ba66CjHNp
YgevNbk0tinMhITohu3Kci9kBihou7QAdEPkBCNYSj36q31R0JmIIkyDnEQ/tsjE
OBHbeDx/GZUbXeKK/Ld0xEFvftPrdeFzv4nXMm7E/FpErSJsNtqF25+/YnGeNat6
ao+BFIZv4Qaw390WL+WqQDNLAATJ5RLQpuiwcMrHLatFY6/1Ob8HLy3ClUQIVMwt
xTy+YVIgSwTXgHmG/ZOoPR6n4sv/AOK8pt/d4I8NE+IjAQVTlHuw8ZOOM3ISwYBX
agwaU7OohgJBYFWrjwiwxewZ4afFCs9bVR4ttQ975+6IF23n+WjHDNJo/c1T9ctq
tkLfJHEYr+9llOL4v0IXiVgPydvpLK1Gu9w1JRWyYN1NWGc+Sm5tIT28ddbebFcB
8TvoLjGbw7jD2Ja3kcMtJ6dzfeY3mO8f2AhgAtCmNy2VxhScQV2JxtJDr68PmEIZ
5ehRcCI++TtWtSgoc7OnV5i4YFaojGuHhhwrVK+kn2n7dPXm3PenDkpBJ7/3FpYv
eSqStLLEwpL4iqWNSnE/c3t+elCX8cm9ClbAmGXi2MfQ5zFfKWTbUMns8AiVzjRb
1Ethjikec052xnLgnNDiplr8t+IBrKyGbPvi0Qrd4A+5qpyCjG0VX4S59Xcmdfdc
2oHHacVGPXEGZvy81JnJr2Jpy2OynyKvkjtMX3+Qb21hFKGsDEX8p562p9AvT0rk
tZ52ITl4673MtPQoJLxfe5jsrXkQ8LrHjiLnj3Bj8oyq4Ee5jvllvQ34K5k5UENH
1yXoTtk2TKWhIbar2inZFuFPbLJJ/QQlBZWmuQkwvzCG5L7xYm0oN/2ZgqPg4krt
MXmCSTm8i6vg2KtY2wAI7uj16lwolWmO94r178zpalJE/ZJSYvy0whifpcKYy8v/
Kyey6EE/xVcK3HhKTI/yFf7EsA8kI3hFaK/99XOv4uS9Ip6v/cClmA+eHxPLVHlH
z3ah44p4CGRCeXriObKDdbf9leDyMg5b5R1MLNzd8uzK9wEJmzsSJHzdXuH8eEkq
HiQDwtT4fbcm4xn6pHQavjVxCyLC4UJEVKf09Z4DYCCBjD+4j53X/QaYdfURzDzy
sa5IhltvM83Gk8bZn55SMANNkKFKg0rQvEvOuwPMwAH/HY6FS7hoD/s4B/cgKqTz
9tGPdconRWaJZqWEKxEJ4w9fcA078awjv427zzBCHLZZLOmEtf2Sbaoadi0YjGRC
RrJZdIP7/tZ2u+9BWp5euHI9w4u5wqsYHCmrvqr5CAshOt/kXzYqfUOSypocF17v
JlszbfcnuXTivgCMHPNsKb6QzIPMPqezzFl+8Ot1W9m8yD9O97A8DP2Zf01ieP03
T2bC3zPCNqnef2bjVPvPFsrJgZJHmUnRNZzWOVvhYsgsYs8VnJbiglscpuTnVUV9
1S4YOEF+h4x5VGA/RKtoj+RMYRqmHpYmZmE6ayv5wD6fkFOGLN82RogmFOpagExe
pEY7T7xtLmpEcLMvzWI5CXsNtzbt5iC7kB9df/rZlt28tb+HamJBdwKcFuWAwjG3
JhXS8QFmqMlulsemRT8pm5NvpTFq2tZp5pl+upl0HTFeA/I76sj985hajByP1Jm/
aQt2Lu3FcrrWl/vaNiUvj0QQcAlY4MRAM+MYgie99ssVthWAPwAnaHhrFFF6TXqd
9TyIP3iJ6zc/D/U3VDfYGMg5YZIqkYMSbpUzuyidGoQNFAL/m+inbQV+6dssEhYO
HDMzcI0u8yg12iBi2WlUkGJWJiLrhssZCFs0sNSxv5YGEz+phIJ1LS0J8VQ9jnQx
lcurmyNVBivPs0jOe1EqeyQz61DQxu0c98j5nBtokb/RFBAz1aOzUDVHg2VA9b6/
uKnUZmp0lT3BqTr/oJK64cwml/wD4C4sgx4G8CiOX0Zo4DCJVn+xl1sIb6Q1WPUi
2NDEw1N0WwuBKLeXeMF84GPVTuaPGM4WIsYTGTL8Lo4rs9ZdeWAsKyy1KsPNpaC6
sBCjTKISKWuxFhQ5NIsHsQynuKxqYpzPlzZa6J2Hp1w+SpjejcgTFLkumqUIDuSa
9cGw0IgLqHiWwlsklygtyk7v2ixDZ5bK+cn0JOes2FvkAFkxHsOgzOL9DB5HUvqj
tP1MuvhCPraNmpIGl5+2FgKzUZA+sRo7tzCgVIHlpdJJZMJuwfXzbkkJWZn9mylR
aGSbdDBxmEgR6PJb0GHwYAQgGZ4DclxguhxTHnz1b4nzGIYDRYoo4dwWeyh7jlJS
0j4yJ9xALeYHk9HLudN968diZ0HDXTj42S3Qnoakk1syJFqmANssyuwpvK/xbUqf
7hr0zohpjevd5Zvr/KFzWcrZR7N4gnauDAZl+fWxunXPz1h1C4oitUNOi/9ocq0n
wSrdX7Mrl+6C3nykh9vJsFo83db65oCMgBj6rTRc6k7qB4l0PPzMAxpcRdea/75a
Tjay9aXxQM4+8JKS7JdJDoZYvnwqqskcIPFvY53JZg80Bjf2MLB15Hw+ANe7BkLH
GYUQ6v81IQfETzBRGWj+bWuPb0f/Xcs422czFf0FUJeSvHl69z+T0DFlBafgP5AP
bY2CuQDCI+rj1z1dBkk6SqcoN5Z+srTZKvt5cE92DAKKDki1WOta8jlwJTQmqVLi
0cPO+7iEuXx2t9GzORkunoieL9Y5jslAEJsNJIY/+I0MrVea4c9LnySVxVfAmwhL
RHEI2Zflu8KNC5Gg92hF+Va2VZtgcGhgwLzPWv/FqKOuoUnAMhrFGsfZlgw/tWWe
QYreMvo928x6j4k7DqOZkj2gaV+P7yn7i3S5ocYr2Y4i9OfxTSpa82f3GMEmuw3g
MvKNwJ1dmFbr1DU2jLHnih42QoB9gSy95fZrbdog8tjGI3HrKMMHiIIRUpRO81WH
XKX7Iyh6TP/BShNIwy4e7Yl97TAbN5YSzLq1TUGEdxlk6bj4XEKvoEPXf0yJIp27
cfCCcXezgVxO4MhSoCXiuMUwOk3MjPN8EwuzVFvKHrNvNz3/Dne5+mHWwlxeBWwY
U4yT5dV+80zUt6sfmD/ivx7EVO37gM8+bgIsHGGHm97au5QIkMsTSySf2IDCK0RM
e6yiHOicpQaxjdn7yBY3Xcojl19jXy1pf/WegEYLfWjS6JyRjepVpeCY8f36pk0V
eTWR47t6AECz2FnWezHaR8GYEaXKvWsJKf0VjNh+NYOc0EoLG8xIDOfRwAO/TmO/
50nI2E2IMF3QR5/9Sx65ksVgXd3YHDDvjuh9y0boOW3WTPHI+ZFD+c1n2UFg4OJv
RVIEeM20kr6BjbAukPszvvMZLZmBJkv2rZvz1lz+Rvj44JL6cpYFhUgN9zmwg1ow
giLWDnUnk8PPsQB/udWLbc+8ePWQsDAMgRkjfKmqxSDow2Lqauu1aCge8RW+ZDgY
Sqd52ASc70BxWG1I0sorLjgvujj9Z/3l6hU5y1jId2KcATbEFtf+BT5+AO40/seM
oa9bCOyjO9PIsgN4brwwTddcVVRE8r4oxo8zf5oH+wMUzywyWuHSYelFjBaNOX/k
f+dHo3awGf/UAXOKqeyWfiDLOCGsK+85WlwgSZSHNyAhKi9NslBMCm1hj6sNx+QD
asnIG7R3nXEbsEYsaRGCOQdz7qgjMDnbExY3fhFdxTbj+pj/ROgKMmndIMHttZqE
aMYgXb7CKRVOrrYWl+9z/Pw6IHFHqZIJ95rT1c1Mw8O719eVrP1ONNRz9mZe2Kdo
nb2eb948vUhuBigG3t2NnQwD1+RHRxeK+4v9qUGoEEnpsQIjTCOxIKOqcnamUCJT
ifr0VyghqMpUcYo7l/2D6Ugu1HWN07r74jDh8ez8fANR6KQh2U3cfx8G5SfQDOZq
9DJwDOGHHewNGE9WQC9G+vZ9TSEDBsuKfh8eNltxsaLaYVo/IOCRyuufV00nZJy2
Tz0drO+SFcDE42UHc+rQx8DnXTakr+ExweIC6xPWcja7aiy6gigAimoi7a5AxVkD
WPzAhXTQ+u4WQU2EcedHU7jYQpDWa7ajMDhpcw4dQErV2cGcSPWvIhyLyVR4YVXY
Fh3bJ6DemqJ9O6+1LBTHDd7c/u6dw9sPG6B7V8pErapEC/zPdJ+L4YklhB5v2ZqV
Jnub/viOYZukm/OeWvIKaSbR1VQzJbOa8BETX+yfyF1xqIoAR/icB5kXryjnS0t5
lFID+1NuJMxbYHmUfUJl+VFcseuQ3VCQOmF3AYd1cVKpcr1RekMJnR2vdDVU5nB5
49UIOJWuLCHJ5qtmdiGH6lqyFSDrOOHEnfzNetK2fVLHySN6MRq+HIr/iIFHZN+S
XCrAQAX0aX2YiBLxZOLxM9sDG8Ob397i1wi72YZSFeE+tjI9mjCZrMO+731fx/GE
hiYecqIXwnciPS0Xl3SN02UXOUhZ+CfdEgjem/GMzSVtn7CMIy+A1yQPn5JI1foy
XNaRAgndZwUmHLWf4KC1DFbac1DKczmjXQF7YJsBlYGbL9PsCi7jLQfTGktOzW+8
8qu1aDNOl3JdYA21ckrdSZQRacMQ+bpWB4NnSk1zA/LtWcT1UKzep7HGro5/Vbzf
rIRrlFwq+H4GiDVqzHI/iWLnZvp1BFchdZty5hGz6S+Bh83OoXoRh6dANhJ5YqCm
7HjoIIV+ula8Wpch9NSpwZgFA0JZSO9dyJZ+vYbJihF6g5VVXiJCgkbmbl/3/0yE
7hkb8tW2Pc8+7bOLUIp+OGL00bzxTYjb+aPUOZiDFah6OdIADm+Bh4zGNnJUBoiE
ufUEsE0ufqiSUC9R5UuK0GcEY0Wqieu5RpSYijXVX95fZjZNOJqMiS16sWAlEW9j
9rlfwMmHJoQ7BLx74qQaqLbS7Cml6oiTDjFchwwZP/2MEun1QZaqEhiaCKpmMmc1
NeYYjxGzVN7+jWF7TVsb8vC/rua1Y7tBx3i1fjl+tewH9bGyf6UbOu3Dj7k7inUx
4vAcm0ppBJG3CMf3qOoHYHU75qW2yQ3V7EYRfMEKaPp1lw5oRzbKiOkPsloyuM7Q
6kDsA7PDOHndmz9NuWEfZwC/kenrJ1RR+IG6Kfw7p5670b7FJ5lL+F2Q315fxe+I
Kb7lG/+14EDbuFDdLah5I779RVxkYY29xZv4Dkqk6QflTUKkbeejbEWd5jhuEoDp
S/PPqTS0RyxlnWZHrKivT5xrcng2BXNYiF23q9j2gY2qCCbb+GMGD2H0ZcC0yBT5
xMPXCEn2ySlsCyQwj22h9IaXtOgctWvZG63Ib3mxAs0/Bx5xvVWH/XQcDYMR6Fyf
Z47Hz/Enrx0KeULGZLoAOKAE5Xr99Eqn2jNCp8I09P2q53LLan65BwPo4y4KAOYp
xt5FfhDQ2nmkg+KXv7d0FgtwSMNrG/+OT9XWlrA23CfRIyvDn60tU8rAQCBVftfl
jLZw+ww3Oa3bi6WoW8/BsGil7fu2EblAG4XGoTJUXc7ZYWgoic2/xb23XOIYBnIl
6q1C1bYsvzeGMgFUMVQBClWEzZ2cfqqFhrfc1gVguLxWXhSWP2xRoT+gUZi2VBsg
TNBroHLeNIed2IEueYeutQwED9MFWBP2FkcqPRD/7nbdMGk7O2KWeAL7zrzqnluv
PNua2N9mn25OutpCHz8kFhXHo6zOh9FQ2qYcPdGWnVwwx3wYvlppE2INGrDPfrw4
Rzjf8ZRzVNqfyd0hZt/9ZPCGYfJYEFnMB+gXESPcDFBTPC4uuaWWOQihHq+0lxcM
SA1ckbnXzef+KxU6289OQKE7NjR7J6pi7Htv5WGjCm+apSeAMehtaOCoaDCAlym/
n2pKiwYfTn6S0EV5BNwHArQVz/ojglA91Yw6C3tEwvA4wYI+4NPpj4COVX8Kgu1x
xgcZ4ea9qP1rAE+9TMVL+7sNmNGWRtWONsaTCmMpcCaUa6/oUXJcGoHTPqdqJHSX
Kd2vlpazM6RvgIhg67/pzOSimdAGiqzSt8nsvevpNZn5PFrYh/jGvFJ5IrPIJhMS
hgljiEnYjJNqFo5PP+ebUqZh0wgf0P7dUjhRYYpjibQbipjriZJButxDq/vy63UC
T38zVomg2xSck/8AIOGcDYqM2s7J5LycHnveS7TBigwJxSfdJ1OrBWFNRiKhxiWe
CnP3PToMRkt49Ye0dcVZpENBkWuj5nQMuwd/tvmyai9nnLeNT1i9c8CgrjrW+xq5
4a8oPD7Ei9Q+bA8xg6cIB9PAbajH2bFVMjBPnkUJRrgaXAjQ4zdwYUZzeaMow15S
Z5TLLicZtBZsSeDUEi/sZ6BhqLVMEHJbycQOcIaC8ZR2FtvmbaUj0tQ3Rd7xDYbm
4VRpJn5aOcB+6OTHr/HnmKOzHWt64mGSGvQhXN/dxT7li6ltuKCUPS6k4vzj4/+I
WZbcnRHdhcVAErPZ3sMEnTxqei8wYvjjJwWMCOBmQ+GyEPFVI4ZfP68SoN5UzvlJ
oPkXxillX6pJlMV9GngE3A0wrUywGkJSrpFhSNBIcQezvjwNENeilQRry5E/SdA5
MRzeslcqM0DEXxIFvSsyrXVNSFb1T47ZZL/9C6CSvVzzQLKfU5aXo1wXG+/fvpB5
pSYpcnaFgo4u4Nl3bJXDQKppVsATKpS/1UNYAvjW6xtfG7m7XCWfoKq5aIFCcuNH
ptLwPMzx8AzrMpcZ3psTOgHSaBLinC29TqAdHlQoH2hyZClFCJeaaOVKVmCXROaN
7vDt+caYyuqF3fEtdZX3OmFe1WYuuQWPsYa1suAMc9vqmzTVhXUNNN+fi76D006s
TTDWcEdydD3JrObM4tm4p/HrZwLUvAGwilyuqZwtHlWrfaUXonCUZtjwQwggOKYP
CHWS5vwdUgQbMDjW7vqn9e2tC0jlNy34zmBpdjQ7AL45EudbzLUeJgQSaVpsNbKx
h1AwGbyrhBSUCoHQm3g6+RJpaBR8efpVDr1x7pUyFQUMG7NzDMkOalyEWUk45gST
IZJZvcYn1RPeS7bCAhU0lJCPLaeN5XSCoGmIQ+K6MqdR4TQF1HdlNL8FEO4Mu02U
+eQTQg9o29lnu3CuK5MbQArsmaBmV0XCGX971so7NU2sGVJOWJuPfquxCVgvjHAa
vIoRbVuQUUKGhwEbEnCHxsA/NlWJh0Tto2zGS7PhFu/WQLkCfl4TsNzjCU62xqQN
fNINiIi5TWU0GvxzGntQBF3xDuucp7NTVnmrYVTTqQNzzPsITup9qpQYYBa0UZAg
fzieIRPnWcq+yafVcfWCptyPPqes93B03MPfyC7/r3libDzAJAL0pw4WnEKuMVqU
bpzRn9RiaT3EOMrGIZVOImYOvBtkrmScaswjXYwkn2EV/Ocu2QE8YLktfdVRX+vX
VHMDKfJeMDXugYLpHEHqRJuSXC6S2Dw53vXoOhyIJFk36GZV/rL4rSAwWAXN41zx
ukzWoSgLtIxx5QRzglrDzKCUh6SnqFE9+O12JxnGclI9xI6tPudBoGnYtclm/4TE
6ATvdgMi8HcPsjgqAu6UthHcAdj1L55O/rWh+tMpfTCnIQOpurBhuHpdm58vh6VH
3NnGtRzkdack0ZDiOTmd3RQ8xlx0BVW5YiAMJ1tVRuRPYN8i4V8ZYAd0t8qHSxex
GKdxfCNP+h6FtulEWEGl2Z0VCxghdAfKb76VYzdTcOg7bZLkSr+Oq3zjQyld2knm
PHB+ITiYxSnkFIvVnAey1E8/6nUw7Cp2TttUMdGh9SJsFG/UulECzNq/zLCNoTW8
g3ZnDEyYD1eRuYJ0BZfAHY3hzdoI1ayiNGLrUMJyYVcB80J3yYLFHWkAiskwlKlM
2s4wiv4j8Gyy3q48+g55EQ91YuGly9P0VzIm8gnLNw5tN15JWyhtFOoI8WEEwJZM
8gNpR4H4rRh2JTiadIA7NDUxqDweg06FfdhvXCZIo+RqxJ2QvUQl/EnRg7VENu/t
gHqNThvNgYozFGJIseQl4HBL/5NFnls/tYUb/JtMxDSh1b3c+Y5wTK1nBWUWxdpw
BzgOrOvrlS5mjwtevBGEwpKiBitXeiJxAFyZEPwEyqoySWhUrUIwW6AmRY4DtCEq
WiHFG6s22VpL9pNJVKocmwFTUp9tSZJvYD6aQeik4BKKEzT2/+gDTJobdDUpMrxf
Nvf8vt0XtYbdgBe2tZBjTe8rjtaA+ksljyNS1eyzYAz+enY4f0svdYPGie13G6vV
UH3r3/TrZUz54dzfxmJPWtHf3Pjsd7E8o5BzAorkPlXb2O27ZgeSa1BVNp/0580D
pCPTTBMck1RiPqB4l6T3jEbc3rMTHh3lghK5vA0b7GJE+xpHYa3ArWW8JyOlVBSG
SN/zGUNH12hKh4SDYmWORmlP9TV+z4/9fmoPzhLqE1NiLMRda7fd/KbFtEdzI3EN
zT6tXxMTWjK/1kgoN3iLPN13/2It4gwpZwQb5uH/uZQj79AnsV+3Z+vOzPD35W9M
7yg5+XF5MwvL8ihb0AnNBHT7tPDB8Wgdq/mlEQtYjleiCnko5fYGMmShXLLoXENb
+NJD/Ex849NT8g9D93NgyXWtSkoL0/rvGSe+wA6MjcKiEhRuQPeZljGHuMhL0QSu
rpnTHWnsclmeIzPTMiG/yMDMpeCmnjJFck6QQmbWSmTRXt/QFinyC/oMvw0lMEHH
Ji5J2EHoFkIEV1473s7R4Y3qfwza/ztJMrRqLA2KociIyBiw4TzNsk0DrMiPdJ6+
wuA5vEGQq0WwBBGoCNuLDrIB9Z2XQzONS8OWf4UJZZ3SE3b3wnZiTbLHyLJlVvzh
mrQqCyfMY7u9yEIOO+sCdlD6/YcV7FHJb+BawOIFoiCFa1mrRRStQZOqx+qPrOAB
1qU6NmGcLkjDO7ajJSNlImHY2eAxfJa3PZaxQj8ylIAvVBgyT53u3htrfTd6bzeE
nMMizMM+8dbOtJtJtIBEA/8rtWxC+t9HoaYpyOHDItCc5Gx3vOUqg7n6RNyGbZdK
3MPqQUFiXJuGwi2uL+rW7PUpxbgQ4xO+Lo2whSxFsrReJpBFqA3FB8CKS38++Z4q
0loMI5u2YVY1xQVy7d9FqA5r2fAHPhJm4uAdDASzFteg5Vf/vp7f37kTZP3pDLk9
MhafhEEWfInXm2nkroGVS/k8jxgNxcEnSq+K0EI2TA545k7WBXZP8vJczWb9EvS2
FNkbYCoEP1e+2TE8O/KgRvSUPyAK6xMMbUWM0PdQDnOwkouR49kvrHfxJRW2QCv2
tguUcJPc8ne2+y1NlfDmn+vmfLV6gIhZQHPGuGAKOVB+vgYq6lwd4hlsv/it9sh3
vMcLsZngoydGi7TswERPUWj5rx473pVI9RKU5eUnn7dPbORynSfj9xfWb8F/KoZy
ubnPMBhDDk0i0qgN8wd+m2ZAkzYUKp3aS2kAxtpR+27s8kPhsQGxd4nAgeQspL4O
Mqd9f+a19bEVZ9DhHVXebCRrLkDc2DcE4Ieuehq47dXA2AMKdqUmYCECKkCVdX5z
JbuA2watklWWxBkEsEiwC3RWJw1Das38FIOSX/FEf/Q8DkZWDRC+ZazkodRJqsb5
HJCu4ZI8nxhEOvuhtvY73PrvcfuBBgLhNkG8sNcu0KKctH4g/jMtL9qVgyVPNWJb
wKyoaGZz7bg2za/i+jO07PiM7ojmPiBm+jHe8I6hmCEXA5pXhCR8kaAH8tSvhVQ7
thmDNt7ZbqnNhiyYSNps7yYPdF88R3NbSNU5ZRn8yr0unG3lWe+Ggk/wsodgqNLc
XnpZdynZWH4NjqlRVm0wzGCJGbeZg7JFsy6/fGVAAcpDhwH0qWrEnrYarsAxE1E7
wP4+DQhHwYj9flFB6R5bMi4ZwqMovBiJ6RXSM5J/cm4LhtMr3cHysTWvjOAV07Py
XqIo/6jwQ9FB36I+JjVwJ04JpWIr6oDcfWIgFLQE19mDXB/Wik2v4KQB8I9B7pqN
csAIwXaDam8emt1TDIUyVzca5t9GxACouR1zmw+CeP8ZzXE3aIlszlJ8Ao3jLEB0
v1rFJ/27ErHA80WPWJ1DlBu4DIAhGFylTSsfKIol9j8+/c1ug5CVoA/d4C3Cr0i0
/ERUGWmP0HGa64MwMWcNbw4FskIkGQVAn6SRod83+cNeZlFoWda7MTY/qMa+qMnp
pFnJyIFbKL+mkLly1qPV0KCKxukjezA3IgHxvEyDMNPUAzLQeNfPvPL+cXO6nC7+
nJSHG8d+EKxnwcX6pKA0s1PFXoYp5lOM0Y8fsSVg7uZYadsDebt9IdInRWfXP2oD
ccuIframyPop6tM8O3P7T7mfNnVMiO+YJlYWDUfaXzX9/npFu5lVE+VITZQgHZBG
FQfVl+K6T512E0KPedDYle3kMP1Oc7Xn39SeTSqMXUicSq+hggh0rmcDiq7sf0Tx
z8o7KcFKw/E+MfETUvySqMRbTgCMJPjdfvSsAVNNG4J5Dm8/5/eLTSfeUx6Z6+gh
b8nKdorxInUCmsX3ePQFmS91xJ49X8Q/BK5zG3fiHrUerjtbx7twbPrQMhLhk4b+
A5sU848+tBb/+UeLG29eWl/URaujfifQ6LkB22bcsXxOs4L/srfxotsUGoksrxoh
XjSf9Ui1VnnDPTKtqhNxz+3g7HGgClxZAtsxKrAG/ignxsIspOwtBLFAbPA1JrGK
aYZ5uM/UuvM5CyPTpdMQph1fFDUEHk1JXcGrzs0BzQ8FAdxxsk2jpkMFjgiLX/K4
bQEgxtLDyF+41qySTH8ntThm693A8YMihi71pptQF6tCYkHY1wDVx9hUoKURu7PU
4sA5RjX0R6nCiBM5mmcTd3IfmPjVfrYygIuFetqprH1OFVmjyQX7GIKKQ2MFe3Xn
GIax5GtyWbEgqEOF8l4Z6vQTTH/d4nV1lg5V1gorcEVH21adSLXPnq15ClHqE/Hd
nuNm58+06w5RkhMzXiz3FUSBhGuoDNaxoHC3GuOXS7EQlea3hO+3f6l4XR+cOiYC
KarBjqxirxnABXReZISSluesga1/Me5RrcUY4hSyG1liwKS8hGy6hjZHZ5pm3LHN
ZQxtk8m9QDlvxxeFLyqIQctrjIgQG2UNy0hI4XiSoQeKbSLpoHTomS9B+EuCDOuL
OkGHlBrCAxw+NYBWom5KWVsUuG8KZ+90h44SENy/ig/fKRBbd0mSsO7d8rzu0tb5
x0jyYLQ0thgeMUHdcI7e5NdJhh+BvVYslDEEOrP18OvoHno1iHS4/bwFZU12I+DW
oZWOsxNutBgipOlK3jUjS0SrMdLaovQZP0qpbYYO3Ks9h7kMf7t1IVDjFG0fSqOg
3gbsRw/p0u6GwYdfQD+KlXK9+YR1fsaJa0dZDcdpkC0KHCAD3Uss7IM3fvknWf4F
GJ+jSn8tWpOYDxbffIDpZFsOMgrPFfBmQU10oAN/OBStIcB/D1lhZXBUH9QRF625
EwC292aOnI9NiN+ZPiCUmIYIBtud04HFnQVgrlDdEGGolAm6HmjM4RpClx/Gxt18
3PnjDTngfwvc0STzdxATsIeWIyF+y2tMfrZNeq4RiyDhSK37sdicCim4QIGJZ/jf
RMBK3s9biWSsxKl+xMQ48AjHsSMN7TLzZ9m7RpuiDXRmlPPvgmm5CWyssULROG/L
75qazj6aYArcXj1ggoyOnqJv/hY2bh8Lww4FQrRVbFzR6+O/YtPrs1UNjkMNIPOD
UQhg2dfD/FynQKQICRFNn7oW9T0YWK8tUhQJR9iDnc5YgcR848SO6ejEdUd+GQtM
cGsjPaDlTzOd0vHoStcDJzR/yZHTD/pmcCFkqcCLp/j/YLYt818mCkO4fJ84+mUh
qu0P1LVZgtddeBODz2qQm3Mhx+Z4LBSmH+a9V2V1+MwTy6EJIhJbZnbuQLwSto+w
8xHArfz/5uG49LkygdJwHpVWjWow83wSwA8Z/6duDJavx7wOQ9yt0/veHRPTL7WX
CXY1HTB4btXRjAHTUfiKvfqZJek7eEh5cArZHubw8pb9siZeaDHrKoVsaWUqBbwj
IANCTbYJhrLPNfDVMcCNkIRy55ZqRALcddZ2UFmPKpiyeOAHGJ3Z62x80F3zi2jJ
g9jzMBKbeFhpmWXLkZdQtY0V9paoU+PEmHfhsKbXxMmAHF9Wj9YRfPBsweDkdpr4
GHqex/GdO0dbMxCd+ukaaqe1fVYv96hpdZAnKJPDLX9RumO6v7kVDamujALcEvGy
7WsYGAatqnTXXuWZGCfNtWnJgzn1ch2OfbZG6DX26veWca0y4K1lz/TWg9rYsg7H
KIGbmCQJz48vRyZ3etBBtwxyMswFnCZ/OCUJZrGomYF2JtVOO20WYPSx38h/cTkD
wdcLfOOla2QOsQW78+4Nf1ad7sOK66jI1dWc4TNl6C9iD62i6Q8sFzuwELIfHybc
IiRAJenYbTJeA0rDswUCHN+bdgjs6/gjF4D4nu0gYxcIA3ekND4q1SBg8xtR7TVU
pAGR75niNIL/ArgBAPPXma3yfHMtKRZREVb8mXdjW1Cf8nNp6befPoWJce5z28L7
COjXFMlCPRVgQ+5shEnOynAcdGDR77GolclRLIRUGiTKREcQursBuhiB+VO3PB8D
eI1GS9o5fNMEAYGtAUTIixWcE8ovUGbYnKj9j9rw11anR2FZinic+wN7hxFmdWO+
06AbkHjRwWC3pk9yjsy7psnL6pwBsnGGDB6cHwIxqmZ5CS6y5LVHOoTwYtKJPFlR
QvfTuZC/MLW0hNMHmjkD2KIRhWz05Vq86gUZqnYY6asKg+NRU59db2ajdWJtShAb
1FxdvaGUDoQOb2ngYUnwAx+2Pqh8KArRETOpBSM4DjmDAVjqmQXkIU4++907ERVl
+gVDLNk4IYIQN+6+kgcJeVqZniltWPKg///o2InyeM9RLBPAdW9fX3RanPrXFX5I
ef9JIl9i4d2oXltpxK47k3HtDO0px0USc9BySsdGBR2GNIj+cMPEbz39poAwEcOW
MTawyjxF+t98tKp311jgDssyRv7D4hYeCcb63SvMuF8KW52o2xav7hQlC27Hn3hj
QaPeSl0LucF5tqZJxEBmZLWNW2V3Je7OfzlBSlI538CYo24cqLyWXPeN+9KHdiy+
MbaSrCvohD/15gErpld4AW2v+qwFDr7XSGweic5gvMpk8dLG8edQs0LLVZksjnV6
rvvlOJGQreocjb06qFYKjvG8U5PlYyakHJI+wCPwkuq1OFIJ3C1ItYkPVzfF65vV
g5nRNNjwLGyiuYLUZ4pPngRnqAczHr7ArPPT4RNbaxBZ4AFrfIEGlvy/FKRU6+LX
ZX7WdYZGGuVbFQVoHA7zOydunvQgJFxsMsyT3bAAdewdQAsp7AeE36A0YX4iJN74
g7G1WaZQ0qzKUE82kwyYcO1byowsGHgYVKrdygVqniWEEnsbdJDJMDFIZFj66pFA
8sSXIAVVKCMDCkK6M5RdW9VHnrVlWnKQ5NTBOBJvdVuYwxpsqNaPEpJMUFRo+/bI
nDAZcAIAETEYUR1LPlDxWA1KMZclTLclJ+hwpPx3GiS7J1Fzh5fkEvGKFQq7jD4R
LmOz2jC9pl4vKVBXUuHbm4M7VQHQIR0g3Ah8MXhDgxjOXBsShzN596BQ/CC88hoN
+dUVc6CPA0BIUS7I1Ed2+EXp9D57eYYJBXnc5z2ml1M+Zh5BHKgmeVq/7nkHXhXE
0BN6c77Z1wydSvl9O2qvju0HlJRhpYA/0+6naQogZ6G7glL/24zYhP6CHPRlLCTy
cX9Uh/bMlHmcFwwBEYES/o+lYt30Wt2FqQslb3kd6aL2XHNvtSu5z0D0Rf4BxrSN
mBTYVwotZhvHmxqL93EcpM/a9AlEvc+RmjC/3JBfcu4M1+iIM2VtkohfK5VGBFXe
/3yOwpyZrNvgMRip4P4LEkf8Xz3kUkMQzWiRPru2MykRThgUdL6CuC+2HVOrzR+5
9Qbd4k0wF7zS76p+myYQPqtsShV3xwnLy3aIf/Q6UX2sUSHMYWGdZMuIde8sidVU
j9+RBXQOa8Rbf2XPCBnUv2xbOlINkm1Fft+x7/adbIejo8rJ6FiIBfNxAVfez8Qq
BTHMG35b9piboXtL1DuuSymXkQ8NHJm/qAvWGFGBmdtPI19QulYeoSxjFzrvu2Vv
yZR/wABzGNO0gCSirAFVsWz7wTXi0/P0+b5eFaSe66E6FXAlb3egbKApTkivuKxa
DO9cj8Kg2+tqz+mO0hVgxkkBf3x/exr3PtHQcC6sLb4SqCg53ClWzj1UFb1058pI
5Y93tgxgmCYO6PnbB71gFNQirAHKGLqn64ixz85+AhY7JdiB7rI/hytiTUUjkIPa
zcibmNFFJeJ7JIkIcrOwUiLGnfwtaDdRmso04xY6wYJZQUdZ5BukGHeEwPljfV7I
mJKW5MC9aZqM/BLimQ6uF9U1VAKdmhdeVwmkKlEVwTQ8A3Tg7j3Mv6oy0elLsMX8
oqXkH9iapk6Zb6aQvtle1wTaXKJiJXWLzlaqDm3CIDvXCtVhBRO5Lvamqv/jzpGK
m503KyS3fL6VlpwGnSDzAIQhvMMon8+fDTR5xX9Qn+GLjnwyicaaujqxTdj5xPLS
N4DnsKHV63JZ4421NoLcgqiGizOCpDQnlVM23knL2tppvtU2BtL+FKYR87xJF6e9
G9xLaHVdt6ISDYyrhr/OChUPX6EDju6O8gzdIHMcBgn9It0DIOJSw7XQLofx9uj3
jd0mu3gfj0JRoyaAGFgZhq0/IGI9IaFPcmN6XA3NjQNRg2XQQkJOmWkthK2ygpGE
yhRboeO+6CT/BcC+GpOnyMnXMPAb79twq/qfBYdgL1nbxri5O8ebXeQN2wLn19In
3/LH9v/7ysnJGQ+egdO03Afy1N49coVj/S9Y7qlRGWehUUprdMO2zTUMmlNTcVAi
N9H4oXaxPmL7S5QXDDACoxYP0CtSKHbBwZZfsBLp88HXDNojqS1Kb+6/UYlNxGhM
VIS0339KQWYDraCq7My1BKzTcgHTaEQAl1kSGQlVY4XCO0EGkDCTRo37QFcw+KyF
GzuAq7E+pTiL9SJdU6RFiel6mVosl1nAha2Kgsn6huIN6bkFReW5HxZsFhOwUsy5
Is/OT32MLBIhfqnOs0FjYhR7Qw56ReGUbHAfSYdOc8iM/0Hek5/4lcBBGlpSuK87
BTg3A3sxcqG+4lj1hz29cJEFIfdgjlDTWFEwtO5XRPmCwsrrbZq9R1epozSRAwuI
ipkULGezwMe2skxyD+ZlibQaO9Fs3MC6qY3HeUhG+tgcmyiZpbch0V7qd04LqA+u
T6boKYCq1hxkMY9hdt0E8/n4daK7YN/VUud52anCCItl8GoKPQE0eW8S2clNLMrh
bP/wpnvEDLAwIXKycLwveGaaa6DoMzOZLwpk85UHMaEcYQcobGsZLGiw/FEyKqmx
Fedqq2cFIPzR07edFQ4qVIvCiBBRcNG6d7VMYSJLTY0uuxzZhem9ei54/pF42cKH
UjCe4NZvGhlSkByYGOJt/Xu80LdpCPxzcvAMunVnHsQc6PJ6kfdLbdjY6EaF2YP3
ZyyjvjYcpkpIxcO+WvQSLe9YwJgVp9Pcnk37+0cAAGXSupbAfeRLVQugAfmeCnfw
42KcT5PKa6729ggz1iPt9sULCxS4/gl/tQ2K8XmtwayTVgXzfaeIUDLYiRXkqo9z
wveKf/hdRAi9pTIB48Cxl2QY56Q2/KfL7KtzMpe5sS/TKLLRrrLTgH5knsd452ED
tST/lOsg+bbSV/3lZvcATRp1mFLAXKKgJ0wOzKsyZsJHQwj7cDV6/vxlM/0f4qXJ
6yRjmMNDmz9iQbvKd5mODFtVkKEG3j/0kA3t4tdHU5vHRUKQtk45trLs04ffYohJ
bEbohSEXOKWkG68iw4YT3IuOj0d+NyMBY3MqExhqo9o3ERuMd7Nto47F1VMTkY3N
FWnnoE91mG0dfZYoJOMnhYTTo9M4GP+cib4aCbZgB9nEJYwiFzKCRl4fWvIuBfaG
XVwGngl4kQAoIhUkISzzHpuFsFKNX5rAyiJX2XJABANJuIMh/I54CJcxcxxPZYVZ
WLvCvOXySQqJ5nSRNU2gnxTbG8nr9NOe1IaNn0v0mBKSsv/P+rB+ERIIhic17PMS
YY3vSU2B1KutAlSwLVVr7Mw+Myxxx1TcZLnfgKDEik5maz2FxGnT9w4zF2GA+gkh
OXBxpWt4F8MJFE+fYF4T+fooxj9thC0yPtZSpw+P2t5a+rCIwlA8IX8NV/KgBiGF
EAeQGaMeVFGGExh+COjn8oMXEbwHz8BJnSyC3FXcTRWC6kc3xTJo7cCOv6bByYjx
i6qo6ukPm4Ld5RcP5Gegp9olD2iO3f9IDeVt6nrWDSxMkZovBHi9iVdbhQ++Xvqs
7I3wu8gOFTVoaH9To6nBFByoQiPNiN3Nkx/ASrEhsvh3sJSl1xLiP12KUqphaMec
x0MjtxGDNs/OBszgRriRm1R4I5IgUVsh5dW8BRVxQDpD2DecyyqmTBUE6lggIF5S
XSbhF0v5sQ1WNDEX54mll0CtNvnanLjSHRYj2pZy0AsTOpEhbTv3SDiEY7yZ7FSl
r9ZcNYRxvGUA5kgRAuwh8bhr5GyP8VpQIg5B/6fq1k6SRfivdjORseTpNw0ySvk8
V5kC0SmuQrH2S7MnmsRcAvOttgKkhMak/6GKasmt6WriGyDhyvpMc0PoZqBNIFUc
E+M7eLPStG9iNdPNO011FbGUZ8XxqebXa9fss0+m/Gj1mL5aB5ZA4wJRc7DDQo/1
0V3wtM1M34/yacNYpwkz2FKdTFS15RXxLQ4splEKxllY5W7k/8axXSdGu6UnAhr7
nMTczeWEZj2BgkElGOHhNO9yxb8S+vgcd8zOyZE4ZenVkJX4d0p8cP5g74G5Rn/6
sl5M5Nua77nEKMlq/bUyMzWKmBto4MCA5roxwBnMf6Xu6XkSRByIp5S4QKKqsLNS
9jglgRy1NjdDMPub0EtngC1nILyMBBUOvhmlO327RH/c4wA8JiQMKrRbu443Rh8H
nhxC7rXFgRVtPPUTSRSAqM1AxrNd+mkhPseOllZWKEXkpgUlTG7TPewhwDhajKFF
jPwFEwAAwog/xnS+LXr0PQT7eop/TMKp1az7lMlLRP/e+RBQLr/PFSz5qpf2pNPs
GaTry2O1UAuZNFjUiOO9RahE15Sb9f2q9bphiV6p6LvgSWCa3TvOeXAvXXwsj1X1
IquXa/UKpxEFtGG0KlfRyxzjNohFwheSJIrUhjgupuv16sXrRXhA6ugHpdzZ9UYn
+CZ25LHEgzJC8yBhSM5MPQxkiVaEgJf2zVCWd7s2QuA97A2SKCnmM3WjZUV8uhKa
ZLpL6QQiz3Mo6Qi6DIQj7niAhrUjma9Kc1/J2LrL3q6l2psO0C1OyJU+0+Hf1Y2Z
zRVfdYsHCIdt0Vab2VoyuQwxsBCkNjc+/CW6XjlIisrgmCweS+2Qx94Ft2K1cR2d
vbDRN/gJOPz1acXnmC04fhTnPbt1zqgjqzltvZL3XEKynSIuGWUX0iT3B4712tkn
g4h9AqlEdyO9YmKgWMQvYGBeCz5WCZnmmCPVFECDQcaU8sk3zmnD+xue6uhjyuxB
X0uaid85XR9i0CM+zipeVfOhOF5VI5WDIMiLJaCOeMn7ltgqoUBrs0hthWgLzui4
81UaGkut8ZegZG4Q/S7q8AFVO1cg+byICcO9B/q6JxID4paZypjEuW4RcjptiVpr
1rhpwhh8Juu/8HtC2lYDmAZAIJuzc7hvB63IZf3MzDnT2y0BD/rs28IMiMvVzk7u
sB8+m+qymzAeGw/V2Dve+A5tfSahP4AnxMufcs1tqGKFMjz0WlpOnLbrGU8cNdQc
56oIzEa39w3RwMhg66dsMvHTWfa0TG3+eZo6zZBPbGUPQ8lXWRtRsoYIwTB/KBKV
0HDr/4ukbOwIZuJYVOdDdO4yk1Q3G2as9qM8Hvv5xOohVKfePiTSj2/FMdNqeJFC
u1HoWPkhHfASlR2f+c+OHkX3OCI2WQnuqN1nKZQ8jBEdNgEswkM8y3WgyOSdD2TM
/G8nbvUlzOff5i3cms8mmrwcBgkzLRZvdtptayI6NxvPMLSxU3ms5sebe34aDYaa
dZgctzGXGUXZhmlbj1Gqe4isUMUegApbzrQUJZ5p3YhtNiNngteSip/3ngAz7k8G
Jf/z5Fp1O7sGkvUF34y2gI9kDfoOnUaNUqKj3VbwdipXq/SPIfLpnlWQpRDQBwLX
wHwps/JVVBUiXTB77RxbN5UtELnd0s03IxX3q4L8vh7kvyMDIq3JibTztVlkqley
Sd2p1q2nnS7h0CDHaWUH8dB/Sd5I0mzgDumf52+R9LghphaxHURktjPRDQvItlpG
HnKWGsxyoTnlvVM9gpKDg4MXs2dqwfOoWd2Ecc+CDYY3tqfDxQNDWsqlEln4L1BA
miABHYKm1o73+RM7Q0h507Ab2x/lM4Bb483o/b1MtCL2x38l607paO8a2hWu2GZr
TgXMbEcI/nE2S2IirhDJtP2S+1xfJrwxJgvN8vX96ZZOXh6M/6HMXx0+rjN/qo4D
zLS6tI5u4SaycA2eSXOOXksdbhv1+DHQ+hYNWeY7MmkhqhzohOVUwI0MgKC4LFRi
aAmHi+6t+Mpjr0V7kKWiOV+82yIlgEdHBAfd3wcA1D23S6Ppuwxy8KDkXu9zZ8Nx
1usk6xsWfLr0aD+Gf3G3aVJX3U+pO3TKzF04HiXn6QMErw7xLC1qq7ZBbDjn3BKG
j8FnXwRHqKlJHrWDbXmeJjspGUmr0lH8rB8kOAinIV5atV66poTkruijgxQAXK9f
LrVOTmH+m/80Fq/C/Zy0PpAZ7Bcb+iWqsN5gpCaFXPuVrzdr6Jq9fNdGb43+9PEX
l6uP0Ep8JU/hjmVOBZURUbbj+sTYT9F/9iK8kBk57z3Ot58cFp7KRFlzHVbI/LMO
omd/OOuZqFFAyj7f8stFT7LVk0RXzx6ivIagGxNbO27/MkDQsYR5v/NYPFJmEdMH
sY8jd4s8bOLCc0Sh8Ipw+S54FeQ8AOKpvUPlVkrh/MmwOEnePaBO7VFOao8xs5UH
Zkke15dJ4dEn+TBsSuW66itA7fke1GkO+mTrwfcCsJI8KSc/YmJoQKC0+HqRNbyi
ZixqVMwM7AV75tnsZPWrw8zKE1MAEcCJjRGCWrwVy92AloDRmcmFKM7kizBMmS/q
65O6gR5sIdKgvlEUjUtLN24EroUPWlaPNtSJF/vJ/lrgZSlPKYQUMVYgMtTbf4/J
QUWe130YMfT6l1IPaC4pRIJMToERT9yeQ+Yf4fUPfYGZtaUYeaZAJOSi5/7Nykq9
iihB9J2r34GD6h15DUznHrPN9Opx+6MyICFZGWcJXklvGXyIIBchcuTnXhUuhuAb
ELE42jgbCZd/lkZ1uMz/maJO8kCW0LkHfiwnJZzThrSvZT6DgJ+mP4lccewq9Wqq
pignwG4ozL3tux+2sf4NXsaEtNtiy9ZT2YOsgqKLd/w4whk05kadZ6Msubm/BhDB
DtMsdCsLz2em+8tlTRpjVmMH6b5Ztbh44M+hOc/fPVUTNQpBdStstA0czd2n5DzM
benJ4eMf1hIOodjeuafw+AsNj4xfODq5zcGnVnkWBQ9IzKElEOVbKpXZflfgPDtN
aqhxkIqCwdt2ZWg3Nr25X2/lVozK/2gsZ//DTaxu6lz3VNTIitA6ay8VPeUcNdYa
JCXSdFAhL2M+P0Qhi1k6/hEKZFyYdugZ2Sbd+amL6X54y/wDxcBdi8iXuDmslLuP
iLbvZhT61CCQiuQDA+rYV6K7asM8Z56lpoemu6VLessI26ITJrp9UDWMYAftwIOk
Js8feiURVzZviw5mbIdMy5UlmOSvzM4a2Kj6Uw6N7Rwz23ikHhb5hjHrfsUNAY/q
oRr4n2YC2/VEPt0OK9n4xo96Oa49dDzyhgM2wTphVinQmaNZ4FiPde8mHFqZ8g0R
tSY0PAZlvGF0AalvzE6F/DvZuoUqvXb6i2d/u1KTdgBCDfGeOFq7b/9IqEIpYJDp
2tjyw9S14ZNYV0sRAMrvQ4XS5SlZUqqyxJ3ACpp0n1fqsUn9KpzHT5psp9J/gLnr
xehv3fFiQe/jZirdM+P1+KJrBEhDaWJw3TKABmcBHNrEO66PsqFbnJPAx5qHcUaI
FM1f0c2angPn6FlfyxJ+PDFQ8ee/ovTUAaqD7wjlwPtS01hsSXfbrQaFJK4QPMPe
PKo40EYHjYUZJbbXPrjvpu6RB6PfBNVUjuk8Y3cgGUcpGr/2zoO0osqi6FV3rsdf
8loXk1VqlBPSOlcgZ4vxvs0LNxjEzeyNDXe1sL0WNhwl1aUnzYntMpBZmSxc0ntS
B+yYHgLEOECPnC/0kY+/d+B5TgMcxTecgkMnZfuzL/bw8hIOM0QsgDaok2pvhNLl
B2PK5iq7fpj0pMDgLNdO+kA+8oX5XD4GeWda0W1nuStfGy9NmifMGYAzKxEPobWO
3VCebg05PpTK+mXjll7D7sGL+xLUjS2gOde8VrK5Sx6PS+KY6bAOhUmk3evlsSgl
rcYj/le9xcUlLjCYLxzd3C5RWSimffI6RZN/VLhSAC0UztGvszIrViHrzmyyLFyZ
dfeuPl/naVdhwADuG6kDn0JY83f/YNsa0yA3AgQp2OUSi8+HivLMl3rHj94u6qdl
NBBuipGfhXqc2M26wci6Lg9ya7vK/Ey9JhKHBCsuo0HrX8h7kt3ChbJewcR0rZ5v
zYOrJFbjhyCDK2jYYSpHnmNhEH4ev8cyJG7ADwyKdeWz7b+a9axnoCZ6Pl1cQmw2
AZPj4ZBQxcFvj6VCAJCs2tDRFYsTgXfuN8ETFUwR+qJ0D2RdmgFuVfMgYopl/Aqx
TY8dN57jVY2zUviHqU/l4cpnZsLOSDobgBSTFm/afhMSBUZBQKdoT/JBekKCH7hg
iGPwvvMusThqBHJup6OvtjsiidzdhV1Y4Z6ei12nDp1eU7DZL5DD/ifubHt9Py04
YYhyCuCDkY6Qxp01RTlPXPm8kT2D5+Ci4lbS7ecx+fDA9aP3HGJKlcxRFSbnahbW
v6lGY12On54MXbYAFKymAQ3VaOeyp05vC40ftxIKSPyjvwnREA1Dk5CxC1KGvacE
sjF1OIbqv4Ko6XIAH6/po6GpmkhvP2CCf4HWgluT22rX1wdwjOsyMYPJ9Xy/iVPd
Ewfing2DL94W4cvl898+Pv0gUjmGFS7Lyv9xNXnOWoYSvdNVdYyM8G/j4n2KW3iB
a1NGJ5t0mi+AawY8cHmTYv67yuR7PR6t5fHlkwqqUeSmxl+lzShesQM9ca1NqOAH
FJx5YU5FELpt3FOkjFwyz339XCNDbWsfJbVnVypTJTzkXK+VqGrwsFpReMCzc4JU
kiq/71CgYHaabrTzzXI1g/Gf+1j5WQvio2PQVXbxUZyzM1ckpmd8ZZrzgeToy0qH
iCvzuiqxmjn6MOM1kAfDbx3MbLDPKd1Cdm8V/zsxsMLHyGo2a0Qi/Ujcbpa4/Tdh
zxgkeEg7WoQODqzIZA83B0e/wGkUsVzCfEl9IDTx8xfKUTmVqF74duv22/QS4x7U
iR27dZ/Wl2Rx4hKZUOav3Sta207fg01Zk+Qfyh0HADTQgiq382X/koCyKWkWwWpm
elotGzy+nl+2aNfvOrJTzxL4nCUxef5cszmD4iZ1zT6xVxSwsKCJJ0yotbDYdzpG
ZmAk7wiGGO2blCYlmE0SUg0f2hWSZ0xkKyYPz8IOdAtfxaArTK+RBr2PYNLkdrkR
EXcL3SMNDBhZJa6Pa4w7kqThqMufWNCbPr9+lJYJs6RyWvdoi/6amuzWMLS4qeuu
6DqevGhUsa5FMgdxC2HxVzyZqff9MsDaOMoWalADtdgoYI6kqZQzRdB8V1rP0IxC
UvXzSCggB7TTmbNF6ASR2qHynvW6ARM76v7M6qOWbfVoe00l8L4nKy4KTRKkzu9e
EcUD3EX4iOy3izm8mYK3o+xzsWGwKqJVbo4iJ2rCIVcwAIapmxodUapD3O7+dywN
L1j30mGKjgMqjRQjK+n3rbrqPk5GA3xYXoAykHB88XV0n7O+K5W2408Bs7fOFSQW
KrBhNNrmye9zHxT+/1pN6TASS3DD+ZT0/Ei6GXtwHDvelKhlXLfPV1NHXXSx9tmB
zOCt5Sb5LoogeXWXYtQX3nAKnF/kSb5tvDfLk21C17GvDOQrnB2ptMuF7Q9yaZOp
lQmYMD8IpQa4aJ2a1yZQziD9tNLngJV9Vas5iLOs/Ld8cRpOt388ZsJyzMqnsqZF
lNlHGVpeU5FnM0uyh24a2R4vu+lggcNMqVm6P/XyzXHAVRg7qXpI5Jj6F3sZA28T
KBGq0WUs+Nv5ebYzFbisIHxysUzxr9O+b5UusZBG1Zy78QCeuDn5HZ5y3oJkA3pB
D8YeHS3j78MTdJvtP0/CtPsan/acQQRr1kOH129/JI/0HO/ytW2hkYHIOM9Zzxco
ZoiVBVxswtVKXgfql2068rRw/zHSUxFAx5pzZLuBooBK91q5juW2jvkSRySmkF8a
4erApeHhsCqbBullBy7DHYl7th1BNCYs+GMmVD0ZLjgDa+1VwcjNH9hdIq5Y2Lt7
+IzBYp/1r/iSKbLlS3LyOT4t+g/cr6HfgahGUZdOR5E1jNsKBOMBV0F8s1E893PR
sJekDjcTp2U7B2G/HsyBzFNDBHAgmIV4py0MLHmGbI5TAB+avRMRnO0gS94fGrlw
xQWaIJ/u7z+Xc3CTMfjL1Sy7on1+wqz3obdeXdgOCy+fValt2VTa5M+aXu6C55gO
02z8U6QM+V8A+AN6atgtk4Ij7Uy+oM/nbVqFobX1wD7FcRBQeCLnodY3OjcIj+Md
npgqudMj62dWvrCAlxcmYEux41SV7Tga1xb7VwLTZN/Ufql5yo+ZGfyIehn/UhrS
F6BuR5McBxB65kDuGfKJBHavN6o4l+09FW5XRRM9iG9429sj94p26SsmUn2tngns
onDpuO8b/+QFlrrKO1/P+rfqm8fBAW/AWkCXTzaH0lytkLfM5Q5kTIPkJF/rZwMg
UQJogJ4P127eodk/ma2cc4kt4XiyIjoAyocfJcv3Mzl3i1mPwwxEQARg/E0Ng7dN
SegBiYRyByA7fXLZPviNBU24XAp9WRLz9iqAyLaJA+KJHGNsMxk4G/xfY61mXZQr
hALDNA7Q5ZidvUoLAyaYRbYjnc34zps9bhGdWq0PYs92xbyrGbqiu/s/OXKZs3O0
vCEJ8nA+Kh9C6ysVrN/FKK6WGC1LoWzgunY/q2TOgTC3+LwKcvCYqocF5asYTgJQ
aPKYEpwcyJhjw0ynF470VLN/pDxTpvs0Jkncne1vM2VOUyMaZvdw0j4Vu0P3B+Bj
MtCN1vO9LC6BFzLIVjHCk6t6q59lKeTvCPXxnrKz25+Vzv38NxhjsXd6qibk40h0
NmRU42TSqX2Y4IAMjMEolOEzZy4Q2X0LHlwneN4qFRAwv4SRJfqgbN7Ij6AiPFxD
D7428YRI3tLeRBX3aj/ufs+FpmQG8iK1vemON2FAcWUcEdTDyQsCg8Kout1YoYU1
X+c4VrVDeaOm1Eme63Pnzvd7S7gNqgoN74tXDtnlswH90+4e7De3T1JrvzqtYM2T
Y/1dDu9IaguOKJLf/ENkjYRw+4ppAJ3P+OHwAa0vRHQ+Yr2ZGFzwXftBpbB90Z7j
lBN6NC3UhNLzztlJ6WeYOJtS+W3QCRQ1J1tatqVkBsO9m630vn09u1qQVKYZJb1g
09TA9QT686mNfNIUxySc8k/D2FeLFauOeLbmRUS0HrySdLqPOVE6t3AJwRv2DVP5
sLX+eqzBkIrMt70xBLKmnIyea8p9Rdt0MEib6h2q7DQrM9ljXygRukpTEgNV/css
xhrl5rvgwZWIfD6GBnooP8beKxupVQzwfnRIeEJVasH0PtnhMMbUi9MrDkw4JJ0e
9WuAcR8tfuesUBWtIMF9cTjyZ6XIBKR71dyryEJ+yF4dTv8vtBBvvj8DlA/9nflB
yAg7O4Vj76IWecHV9sPJGZ2JB27uQRWPus5PvykRp9R30CzHx+p2nVaNwtf+qaBG
CZErlQAasj+Z3VLLAlScU44Yr52Se8XCtqWf2EqKHMG9/iIVEzvFfJZeS27+aNVx
28WrIB8urkOStByiYbHkqv3stMT/oOunHS0MzBhr/b+lLQshpPc0D9ZmCzBeGr4W
CI8s9YMS0bSNVO5mAKM8SbidBh0GZ79jFnaR1m2v0GTzJKTqlIyyUWb1nlRKP4uf
3AJHOk7698yVF5YfOYbcBXEMzcSGM/Yp/a06xfKQPSu+kIUrGEgLR0DrHNt/wbGZ
TA6tFQ03Nbkwco4Y2Sfb83gqZjh7DdZ2G8xgN7Uz6Ks7HRNCaDfKGDuurWpo1U6S
i3hDR6j805s7pXzLTa63MaqW2icfEziAVkUr6pn3/VMRCA7WTk6L1DtU9LIL6Yuh
wWjNIko+Jn+PxlXJ4ImA5a8PkW9qO7tL9d1R2vxzyjHaQd/OOUdg9DR7urdvyNvo
vBWRhhFxJOjeBs83rU6AlOhNiC5qB3dCtJkXYCnu+YmuiLu0FAtPfWo+1gdl/hcT
8cVZ52erKrxZ930pN9QJ41M6LefhKdemb2IoTu5JL4DpBYe4EAcI6qz+09sgZbex
+LMCiMTSq297oUMnd3H8PfQdQN/pej9wipyjrEkF4tlC4i/INBHq+loyocs9Ooov
V+mteJjJSJALTIHobvkr4AUcvSMaY6T3Obu0tmOaDNRkaeVou4X8PF7SXB7E6o7H
w7Nivu0MrtWzu3DlcXKhnYXA/vmM9/niEZkEaa337PB4fEILDInSMsDZ2Q+M8j/O
xBON31Qd02yR+m0MOZF1Oeby7uUL2SAYQTbP84cPUvaE8g0s9jqSMd/zhf99SPA8
uZwAJL4PUHcTBt23EdkN5fgIswlm8o9g0m7YmfUG0fc+9AvJ0GzXtuRy0E/Qmbsq
j8Yzyhlyfj2d9eIRYPfdLBpRTHI/5OpPf01tAE8eIpensvXe+J+kbqGA+DrmJ2YO
z5hljYLw/e+Jc3ZHYlpDyNTlC7I00WrZ/XIFgAD5OJTEt4JuJYSbga+MkbFm5jZJ
oxABwOodnCfqZ5MchoBMicL/sbW1UEsD5n6UP78BJSoUuJCZxR0X4BqNVCmUY7uL
6Of7bsCtacPVVWAygGzKYU4AMaZXXkonhcIqIAxMQAjZTkjCsdwGqhnmVjq6+Xj5
sG8H9nf3e53We+puXy9gcwobr6NM2sKcnNRcRGXEMHvrC484q+BSguhSsTLKWaw8
Ox/hyCWjmMflLaMfMgQCM9UfYpkKQ1fKjjtTg7bkGXCDrlAVpeiMu0e7Er28LZ/M
EauuCvE242gT+Q9datc9ex8WqKe3V0wFqhLFjoOwgTPgq3F7fefDN0baxN3CuiIF
m8E6hZpeZqkBsd9cKDSoCgqreN574c/e3gBDwo+yKjbb1H1jPStyo1ktXvSQevGh
rQs+vve4NeqxBUSLDB7wpLzHnLp+XV0SF8JMJIlvYMulWgz6oh1J/spP4XwVigVS
iSrKCRBicGayQ5MP5VJV573/eepINX7wO1rXy338roS3PMf/eVwSrcq8PBeNU4JB
04B4+URuvyUSPVsCz1GXdiqw97sIb+FO2v2r6oXoUNjduWov3fFi24vwWs6RWaYa
9yHBv+vL9FeLgV5EdTIQe7d8bJiuUda1ptNpJnzWt4HJXbcdz/kWR1/49ipKoqCw
vWT+wfAo2Z0Tx/LQQLsSuOj2xVwYRGDF9zs4W60UJrBvX6Xa4dXHxW/DhTMxh1Wu
K2c7RMQ/2ZYT9rxFI6BCbjwr0nZqjCrLJvCsdSF0O/vg9ZlrbFQkcZbBwDkpczbF
nd53xzqwZw4gzg8BV14iAQttBbVEza+X3vyR5uXce+k4yTd5pqSUUpAQwShOuG7z
3uhbHLtx4rmirkINowSutI3PALhZfR4jsbgdLN+HAdafbAQjvMfuVP9ae5mJBioh
83U665ZQzroOMWBZqSO7lpsmPaTiuR+RCIhmmbFe7u4kHlo5Vi0OMxvzsGrr7gXS
PZUrrRKggRZzqAlGcslqJR1Wo6Fr4Hbawh3L1kHfJstE6iI52ocB5bc+fn65IBFN
ECUbYaxXu9G2W6EM2iQnyvnJxf0kWVPBhxKHjo2AR4YF0r84oyi67AkJbueqOjDp
uklmu1IeFkAFj2oTh6MiK12v3i8OHzHtjeyRiRkIC0WRm0QMCgx6ueWrrqQBA055
BEOBWK2q5dbBd0ESXlsxNQJ1F0TNeLOKZoPHyCyy8rzQfkid73X/9z5JFb1QD5qs
9H+0ax2Z4enOx7HZHJbqwlBbWnGMJzXjPQ6ZRbeVxwWjpGDlRE54LBWM0cDqwrBn
1sqwRq4ezSN8zJ0v5L0pmJfpttJ7qMxBI0rgkFB+zm6oZM2QIKyUXcsp2mANDXid
7tQySNI9CR8lX5dvwHONomVZcP8ux5AHcAlpQ7VBUKENY6rWMoPBSSVO37D5e3td
ZQGwg6udbrvwNbkSf5D1ZFw+Rm189Zv3l0iLO9ux1jJSKTqEiU8vge+LJ7MZq9Y9
2ZnVT6s1sPqDBHLAwXKyDEseyitqcV2AhYfsw1s+pkw8zR6+VRghiYEppJQQ9yZQ
/inVMV9Ybye+0EScaSYflNHZdzszwNmL9vFzRDfJZPxXiibrzL9qBL37dMYMz2Kh
MqIPE/wIXGrPv1e+UJbO87ha3hD6s6szXdhIOu23AYM5aQxCBTPb6w3fma21Orq0
pcnkxZS0n+1S5NVWctA/YJj4fI2/gZ3N88QTHYvLWPTrGLxa1tOaLsluud8s36Ut
uc1V3a4oRcutbVeP886h+vk0zcpsshSneKaupYeFm/RRlcxP7vZjvFiypWXGLfXQ
brf8liR/mzoK0TObF2C4CJ48dc/KOEus4MbxdA9ZFTv6QF81+d1E/WV5pBt/GyUE
aXqexRAiJWemg+GQ39Sh7y7sOiSjtz1VtF6wicawP87D5Hmetmezwd6fXcoWZZJs
HmT884y8t1nSuXLvTsntodPB4+u6WkNhvgOpQDVlAuy3p6bO09YXIeOFmuWOPyAF
qWcu6Bha/1ISSkF5nA2TvzvvjEH0kMrsPZdTzPsRX9fYmAt1C5jOrx39bJC9b0h7
KJE3XcjDrk1EKF/idCnI3zjhor4g6Iid2LnsBgsx1aCt0j8BRr7litP2DTG835Yq
7df0ymGtKpk6YRkFZ5bxl8ZZFtJpjS3omQezH7JEzOEoNhN0nPajTOYZsVazpbpS
RJs1Py2ymNZTDnMnwrqFKkg74sULC7sQax/Dp4VNx9F10nwAT/c0tmsjT6Aul/PN
WM8aK2qUD6Z5WJqXDVpRlMJwShlqh8fGw6MQUd1fOHb0zvkHZ+aAAsadoGsja2MT
gG5r6gj626CHwH1Nxds40E/H7BLzm2vnSt5GlBy6xJchvR3U0WnyiP7v1JqtAcGp
Rkqz5x5C4dbuITwb+iW+q1yyrAGy56dk3kRwkRzA2fG/qrPGMUCbqqwSdSFcAoNg
DyxWAuYgBK0ylYg7bE7S67JF1RfxpyiJHXLnTvuhCQ8xkpVflL37XeqoC+3AaVei
t8YGBVXnkTklI8TH2cysHKLIaDBPYo1tkCjXWBOjRVHTpu7nWxdm8DzoxEM/9k45
cwEAwqP8Sg0YlsIulkJs1sLdq8j09P6AjfCG73cfx0v7jtLkSbMwxBMe/dYzogx9
BnFCm0l6BCcmVNk5i+YtDAPmTVHP9zuRMjhCPS0gTYKNwn/x1zKcFX8wHT2t83XZ
gmkjv/B3ExwsReNWsvCLu92KYjzGHqK4ycnlbUY1Op0GME6F37G93ehZX9Kqxmqt
iD20ntldr6qSMfx1qArjbeVGv/IvBZ3zoNYZsPRyGiQzldbqDJ9Quevwwu1dTPlp
+xSggO3FlUsirsn1REiQnns0RTgMVXxRUaaLifQ8VYIjdWn6iEBkYWa9FBWj+hE7
86J5KoFjeClqKbxYx7vsMTj3HaxK3DtQ6bPUPSO2lMWmD5qZ9Issk7zAi6I4W2fm
xmvXwYuP4riOFDWSJuZ5YDMabd4iXQNBI8oOkD7iJP77bDHnLXQ9m18em5xPdnup
vYMfWkXwYVh0Mh8jgDgpUXOv0QiwwXCZKhSa54SK+qbNoL/19XGsU8hNlw1xa0E9
G+8gOAgiqt8kMcEuY6QJzc05eV1lr91W8tyZ9ofvjxCsMzN49uoLLjWlpWA/CyjB
nG8duSMOZxckHPp01brCEEYXhNOdvbDM5YqOLJORhBMDbwqXyJ/5oSF7VLCWFKLW
l1HlLIXgLSM2g+uti/9EGZQzuarOQZSGM83+Zuqb1nPwBg/B/2SL02ByjDM2gJPT
tX3ATLz9OrhT0fytvVoy3/K8oSk+Is1Xm9IgTTqxGNdHMywV1fWOkot8OIU0rZTy
LuVB/hy2IIRXOiGhJRLzETZAPOrMvtJgmEyJ/pyNWvfnMtRd8GcWd8uD2rM1fbcp
y1VgWNTxErlWW7QqFlRfB5/pT+w5vBw+Rzpkj8pL7fxj9XgdRGkkEPwNvPi9r7C0
qh8h+DT0wT3zl56Caz/A06uNEVloWmSZZkRFcF5T5/UsDdn0kIvmq9eVRFIw13Ue
0lqxGuXZYKf+Fqf1HSVhViyNBCqGXWjHB8cZlcsWp15LzlLyvPyj1x4dz1XUyT1v
D0w16JxTEz7JCLFcyLz1N+NDCcGbHgqY8HwASudNheZKowIul4GnQ1jotluNnq5d
Yyaj+fkgnmDLalrN/lVr4wQlSy+TNEuSZWjuHuMntDqQKduafpM4Nt2d/Dlg+9xV
GDmROVL5dzcLgtYbkMLSnOFnBkWT8gbbeqDj5UHlefRHCNaq7MMUl/Gr5cemfFWw
QMe5uUbnH6THooF/822lpy0jy7It/ReKTIYy6fYOn2OGw/TIWSmMngiLm+XZOMHE
okRyekoOU/d04+oaD0RMHynXU2Con7ZAar0r3qRPNDu6nyI6690st5AC/Q1yp9Iu
gzgW5/KncfdRlOA78HtcEGm663zruUfgzqs0WIWBLLqPg1YFF2eyHa9ba51pYkNt
QKNd5XjFOv7STsNkkNxCTg2MzKVH9LCgp1fJff+qsAmZXZaCO7L03OnSe/jqPI6G
sk+35AxY1wTw1dYtmSdBEXTTCg8GloPqUO2quciXE51MHxSHKhbobaWQY/Xrm0gx
MsK5d9+lT0fRmtZac+5QI5GxRiEZ3BE1G+KE7UgU1nkQQm2ygSi/EU1AuZP5eS+Q
69Hx5U843AoD/zJetTqc8fyxWnzNZjTWBFkxvhFYysRmJCWvl3KSVi71rK1f9xIr
sj4Zzqd8MGqo1Lm/h1S0YggQWa491RNI0OBpXpn3aGMu+pUkzFRT99Y+Td80whSY
QVUf70ZB/mD2UJaNPQxQsWzDV88e2EHGbuBx8aSHMo2x/pFWiDYs0/dcS0/TtZBg
NHiKM32nhLqlDqXykdujEW3KTBWdDiZPX3ciun0TB8s466s0DTHwjV6Qo4kVdSZ0
t38FS/u+7qHViPftK4q4OjRZfqq4maPUAHU8OL0MlMeot05dpJSYFIon0EB/MLID
/f5yJELmQXHhnjgmh70y7aBR2FLue58AKHBBDI6uvawuWVlg/5OeoKLaspQIRXWM
LS9j5Gq3eFr1eS+/EarJ1R4d42uXoFP0lXzHKl3ddGfYfa/cwmmvrq23HZgYSWAD
+LEia/9PCcUJAZtG3OetiD8CuttflisExdgVnW1TOkNIVW9Ccqn1O2krVHhYTpWw
LDNFnp/XB+eho97MfCahrQe+UcBKCrpvTvTuYsqHC2R3fAVNP6sm8iYJhBjhoqLS
IEGgdwqxPxj4UJEtJV/vJtRNoaVlGFQqYrwInM2MohHCDFcb1/6JUB0n59t0tx6t
wmm1Gf9Jir/Md7VSWeJhIuq1yyrHfk+s/2aWf9cUPU/ext/RRbyFWB3YbDZD4ucE
1zGH1S1JCSZBEPHX61I18abPdNj8ssx9y0jW5vhdYoxlyBysLGOdULSU0SJoF6Cm
rIln9RP1Is8xLvFZu/gueshYkn2PiMpnn2obXtyX25m1fZxTn9J20yQJ42tI1p8F
1c7ptXh/6fI62kEpPP2DC3AGm3OXf3sFTWnDVD1C4KuM1BC7Gm88G/TeNKkcbmm6
m+UotOTmDhne9x7GWWkB0kNJesEpQuQbKmrjwGPP8NYDLwdRGn+BVMyEj1nPE1u9
luG1/Q2W6fIFkeYsr7/CF+GDZoU3FqSfjbNmCDmw3uEvBFjaRWV/CYfGob5xxX09
PW2Bp3mn45TEXfB7vQ+KUumJn2EY8Jeiio78vEm7oiK4j/7O/zdcbTAwXofMBF8B
vxvLxohbqZ6j0uiGBxLp/EcrAxrZoSunZWnYYeLDKBB6G2dSzCjdtk9KPhy1iKLe
f27L0kgkzzRPVAnaBtZ+Mx8GxnmyOu14+EAVRqcmEmMtcZsVgLqCXXxP/C/Lyrdl
ZJjVKn1yh4X2xMfcY/Hh0MsHF94Hxcenq+Q0qjVj7omv07u/NWo/79em1oDmynJv
vmcjn2N2PS56LZxy3teaQ9H2dCR2r9gXU8WZ1ptJV9YDZDblpVHmvDC4PpQzLv7X
gJtkmB0bu4ssH3M+NIbcCxpJE2knO8qlZv8+COhe98nr8JNjVkdX9iZWCEyaDWEK
v8BIrHfBD65SqaVPQVAQ8tAjmmntDpoPWzVMzdJghzvF5GRAQoU+5XuUzgwFildj
fCyff/pD/QtnxrRh1dpebo2+7BmFET/UP9r9iTzi1LKd+dtqEPSRVTyIu29aCBbX
m97oiXO+NbSDnPPSqOWbtEJ3V31w6hfXdDKIfqBLizcmGeHyEX4OzSmhB69giNrT
m/ydU+PRzgb5MssPspOg1F+X6uxZalG8ZkniP1Juo2I1t+uTDoGA58kY0lSNaxUz
stOBuF9m3FxMuzbTXcjcZbtEutOj62p6/VKqnJw9fLR+/h+BwKsbobBOvoU1LGq9
p/nMmuK9h87g1v7J19Ep3HOBNtS23+kjGo8fBhC45chPh5VU/9gdb8oq8pd3RmDS
pjDlo2qq2cFVfIjgVMkzF3LJrziM9BnnBYYPKjwiQ/APMYZBBviCHAAhUd0aBDgW
xnlMpFC7SkdYXVKvFI8v3JpANV91Ztok6PX5nn2SPYj2otUTyUC6koyy73BK2Rk0
lDqZVYTyT7MoWUJjXa9amHusyHPRr2lL/jbPg+fA/jLQkTCzFXK4ThC8HnufihTV
vK4hEJOimNyghCneiVn3T0n5G5CFjv+5Nma1oju9DVDfBJxHdnC7QJ913rtc8ATY
XVvJNrN6/LiNmhuQZUdwrl78IPNBLcd57Xs1P2Ft5KEL5vzWerx7DOzpJbTmJiD2
XTx3r+Rm6s4aGd0gIw+vApSP0aJdffGhVrdRbYdzelsbNhjmdZyjAfSKQkUAke7s
xNmTko3su69DDv0r8xAw5KGrzz1KO4XaF7BUShkO0q6kcPpaXnS4P6ax1RZI5cxM
EPZSBSOPjDhunj20gD7D6QGn2P3JW3wZ9cCrhc5SuIUlnkYeF1Fg1ea1vOYMmYz6
sPjL4MrL27oRjKFbjht5UblOKKg04GrYtaPlo4tlC8mkWRRmThWgQc4+Q1MXli/8
N5SHwA1IpgtfVbsYJJiMtnbdQ9H33wXcKsifs9LlO+WiFmdATVC8IwmRfop5r0aw
t6n7p0BPMheF+ypWYf38huNDvgsGnE0B9JNmP8LboWw60rhkFcdpekDlHIfzQggZ
S1SnaVJgvwOKakZ+jMsA4NTHaY2av51LKYgk5roGCLFSGn0/vPYBqnzOAYB1oiHx
o1siI5x0nSC3tEcYMReh9vG2SMpxWAb82lNZNCpkUw1yKYzsxiJN1e6z6sdAyTXN
v3ybA5XdOJDRKvUql+luqxnPicWXedZs9wm+4gd5471ackC7ZX9znzAGKe9dPaaA
6ahVQA/OC1CQAcHvOKwFtYRVItspCeGv2KKOWqoPVI3GpdzLjeFzZDXj/7KDDsEv
w7DPduMpONcZEPB53PsTZ4X6lDY2sKvd0qCmJ4pjXMbmJMyeV79HrRhCwevr2+Uw
BjuvjHQQrBux75u2+Fnx19O5NeaJpaNIEdXSZYB+ELh307eYEYHjLLeawbhZFFF/
4ug8IHXbGZzRUcJcdBT1oIS0MVWMDUYrzc0h7bN3+tgdLRc9mQSrHGOwWYVHPbeU
aV3w2qxv2IkyDjFKKoCp1CLJI/pnEj8V2DdwoHgAMj5E71keuQkI15S6utG2muaH
xmOSbo0MrX2m2O5F3HohgL5KUGVoyQxqOpTzygEhZvvLoLuhJO90BP96aKAPJyYT
fYZCivW5hnT8Kw8aKnn9vJGv5+qIrXsM6MH/SEwkREPaZgGeamv7gidUy/m0ex0e
brBNes+tHLlzDSaFilo/mIog3EpJbrTwwTAxxNHIpuG8TUZrfvQL+Dj8mmZiZCcu
1TDYHAn6kv47GYAF1z3RoU+3iO9chFqDxgyZAwzp6tVu8+WsiVSOrqZ/w+vc3RvP
7p8Tld8/RnIgIhs2JnDs95H8o8JZLaIj8uETF0HJqHkrFWB4wnvVsO5JpjV52LcE
Y+zgfelkUb5a5AWL7prskjuhyU2TH0JH+H4j5cgRcxtYm2k4+D1ad3FxOo9rcwr1
pLhJmNn6e+xtO1CNjcuPHqRtAbRc7wf4aRENDM5SgyQ6elNVq6fgotn8rRREuQiR
XtIS94rIFtGcmGJKClGOMakyf9YioS98L51XumdQ1kG/0UJ11bBJfDQVf/YgLMZc
4DSQwUgYuaaz/v2t31yjbSeET0kjs4+o6uB1yBUBkhrAdZjDDlaNVnepF3JPNuH/
HiA4AOT60hKSdP1ydHO/xX3EI1JQkr76fQ4VV6lGJKtOph3B1Y6F3nL7i1Y4tCIa
QUbr1csuCvFjpsJLV1gS1iAOjaJz9FcRc4mvZTnbwBZiH1D53VAfnVzStkaXHNrz
SYStsJdS2OM1hMsleS0n8/rdC0Sq4UpJwz86FZ1sjjqjBxCkKMqKD380HkQ76GwX
lc58XzO1WgFpOZ02gT1QpcwHJ6rnxvlA08nJ1GddPHofLu0co9D4dZF3JBwsa9AX
O5SZhceJKYVQLFl0Z6YCfecwDhWXxLeLDP3YNrPcxRONFk8Ntd81bnH6yMqAZcSN
LvhvkYP2WaOWGYQ1to8TnclWQyukZxk0ydH+apsbYEnpJvl+Uj8kMFGAAhhIduLO
Jl7rewiEZDYn4cycjtPav6KgpNHHWGo1KBq4Xvi/nwBhk/pu5Qk0VUZ8/8jpBBgB
CjyEMzB/ceTLhAX3b5kfOmiqPsUfERFBCmotMO2ZQ0rpotMbNwCGtIVSWppjF4VN
+0xPZzMajR7IFYN+y0EeJK6JW9p09uhrLkn4FihyCnLp80A96VCD31vt8Q3Otsmm
fpZaouys4H0Sdijvj3fIOsyQoiwtUTwei6WmRDbGj8p7MgMk3bkenLmarREr7py/
2GV62SzlMGC0iIRHNfgYKMH4KN2hHpefOBWxHLTtiQV9jtyUIrENUfU/LdnrAfAr
LG+tB8Y9wao5LesZaoG89j+m/l5CRrZ/vjJ5D5s2tV8vQE9dYAs83wmNMvHozy/C
IMjlHZj7bmwIm0dpByfCX2b+wyPvXYLJOixsGjCPJoHktdds/vLMnTctHSSmQAPI
q6+KIIikDfgdsroQNB7SApUOG60TIfeRJt/q8H7UMczM3Tznt7IisoejLbkgOhLN
hJlq/LZGkkNd0KQAJP8WMaJLlJmKnE+7o3JQ3qhi7mcZdCLpH/RyQdEMOoY4IEVE
JlZj1U3n9/cs3OvBIulOIUk/xHQd+86whzUeZuE2Ixyg21P5mpM7HrlXOeIFslgL
Rrb/6+jIm3XZOgsRBT6B381amP0IiVsnPN/C25T+v93acAj7zB2SQV/YO98cO6qb
CvevosO2IrROiLVpBYEQBJkwVDPsDltfW0/wDahChVk50XdEzgPyFIuRRIggBr3t
x8mFvJsSTyI5wFvkw4iU1CJ8pSH54ONSSDcWpuBWlghXR6QNEOPlF83Xxgl0RjsH
t63NKCFCsEUGziHYOaBsrGE061zpMxubCPKta4eV5ZGk+y10y4mKXkbZEdf/xN6E
qn6jaQBay30f7WEotGfp7F8plGT/4KSxXolhwnwRtAn6mnQUZ7nlsegsbZx/zZW3
6CFDlovKOjopJ3vYloxaFMF8cZPbJNoIm+zSZi6w1IxQFMHR8nBToAYNbR4aQmVL
RrfmR5AO8stqCkYZIhkpMShhp9e8TAntbHB3Ji/EzEVgJSJK4v/Y09vIElgrLddO
keAWPKp/y71KZGk/lXdSFPONxO375nVuK6b/GvsEqODx6T9xXZ0sE24NsmdweIH5
nKMk4Lk3romiFAuL30MPSo5M3L5Lz+B1xaEUen07xUJZ674ILrKJN7/oaMvtZ9LZ
mlGPU/gWTd8t3GstoiTUn515NqkQ+CnIV9NqyEe0ImQ3A+SXnpFzBCLDuj5DFD3p
JrJLuHHYdguxva0ine9xFPTOLlJLxLMDeirMDnrSBkIIr03D7GDKBwFOcpvZWFqo
E0F1gZqXQuOKLURrCgaeBPRJNNF6juhbeMEYnbldVAmWA7UZXLD73fglwRJFOgYo
AjAfiKacknInNOjdRjxK8gbCI+ETvWMBsFGiQTH5/JrRSXhg4uMQVrTz+0kPsmRq
foZl+y658oqW9S44jVV5AI0PjHfyl2T647cxRNmHruViPB71/5dQ2TMPfPUa92eM
XsmR1YKnxgBI78IFTryZiDZQ9rpTVGtILKJNyVd1PMqG3DPfPM3n12Q3LqneZxbk
qIE7s6MhJlUQMv+HHBsma5rQLCFCcqW2LWAjrEB/3TN8NrcYc+HTGg3Hdofwn6Mv
FbCBmqaGY0dALDmzoPGUsGBz5mirsK9zONn2VReOzVCrm4vJ6Bt+AkDVRszf2XiK
6X4Zsm4tBwoaIAJwRaqCwQtBVllJZXy7DMFknN7Wfz7ozRDNM7TDERLFl30V9uUj
BHvAvtj7t3Zsb9HzD0bhTQscRnbu/icT9ksaUfpAU4cxSpWYPkkmi/s/Cq4ZphAn
7w9icwi7zo9EZlkt792q7AacXwyMjTKmL6Sg6mG06LQBvJUx8B0bTQbtGtdv2+wQ
PdNnFJGm+Ptb6ryehD7vYJKBuHPZHUTYwGIqMJcR1LBw2138WYRB+lrBWFkaYulp
TQDBMMJ/X4FtZ7KU1BD8oDIk5ZlbVs/DgTgRHs1xlg99svrs4olUvKValC3Boh9f
NLvk9FzLmMm0NRtzClQC8aeJsfusLBu7A6ANAJuLWMPwbUYCJHzY+/9H6vzelPjY
SDP6qWdTb1OXXCQWIfxNM8qjuQP3xtWNiQeJSuwJ7ztMVS/U/fLTMQn6iwv0NTbE
d+hVh2YdknAATBbUcIp4mIYrZPYkP7x/d6T1UbHeZjVcogoOSeeNBdumNGzPgKvV
m5+ngIgPHkNTVbuR396ZJsgyEhXgJWa1/hyABO9qsZe+ObAbwqEB9agYXoI1BlKq
HBQDn+pqW1xYY2m3BAeIwlgOxheLeuatPt+F7VB4gn051YKj0xaHyFn6EQ5eIqU/
O1pfKheKeoCTcoQ5zWQoNSZIVCk9olvyUeVpxtvYpbW6hPNdVI6Ab0VzonWk3Kvr
Uk8Au3VAbHz2OowdepBG1TGCnDJLqSOUfuc8SurSQrsbVLs2kUGuUGjGAqPpLitg
bFvewELFw7MmHpI05ECMt1aXmigC3bTb7dZkGfsb85/MKDChuwknQ9qaM9NJUQGP
HUN2CFbHdMDgmZ+RO8KvmmiGFS9Kq+rCjbf59Z91RSRIZw87QGTe1GSHgx3EkyCj
J4ibQmWJecZn7m8Zrhu5PJnDQMfv+Zfr4fvA3U4Yinh56QGU6WkX3iOboVh0PCN+
jnwrL560Su7kebcOrwkDccqZakayeztMrO2SoS1rxwn6BT970P+O7pxmG+R8KACh
fgWP5wGDlJjj4qHVodh3szIO5v29JESSgzBwGWB/NTkaESxv4FnrJabUpYAyAHh5
ipe9akw5KM+Vx4PzFk1VEoO2VNr1F8KHZw4/G9CD4vw049WoFqX3grtNkHEhBfPA
LN4XtzDoeIJAnUidgeuixEUY0Gxx4aup7VGPTAolAfnv0DFjkBEGzYf/Pwdw2NO0
wcg7hAzjFpGoKp6XVxjaMCojgOs9zOLoRdfG9yJ8HTCrftVYTaDoYWoukCyt64VK
8ckGz37nhhp1wxd4nR9dOMmmpYWcOq8a/T7LbueTHZXB2V6F7ItG8PgETp5v6Fdg
kSNzr0r1CqNbedEHdar4q1NGEv/vOWr90A5nFNKiun6ukufTRdEDz1BVlxyjwM3l
Sk7FUjgLoh7BkqjtM/QxR87x+O29blMwHvdWrHU7i36tIsFywudclg9UwgCJQLxS
h/y0Ykx0MwuW+DN0jZFB+wYU6876dagtR2zYAGIS9Biu5STnmGKHzrMCh315cbf2
FdC58qOYg4DSlzS5LKPxAzY39rb+OBl5FV9Y1TgUgDeVflN4nDbmIc6FNL8ZUqit
wP9Q//TZop/gBxRZ91d4jVcuMXRG1uIyOdOuvrfWMpoRjiUOsnvxjL3bEotJf35E
OBFMNTyiZtHEfyjN4Okqe2QuNmXFU0XweeRxV8nRdTDLZzbgFzUVy5qsPvcce0oQ
D1KQU5ZD7nL6e82mFUJYoHlGujM33yvF2mdZdLk6NFcqiqiFtMuwSz1iYVdtvi/Y
BwKVjeTS5+wFVns46bN/op+ncLxJuUWhwt4ibmaTHnD4UgKpA4xsqfabrbkQQ4Zx
sYJA22CxFfh8/0ju9ohbSZYckXvoXzy/fODnd6zVvB8ieMEYFIppNBjg1YaksAxt
tAlrrR2spNievuXBd+EiHUgZvTd6JT5brEES+BBn89BaqFGwwBSTFACL47hOyvMw
L3iZ7CrblZQ0RfwIKr58MN6/X7sTnxG89PlGGpkPogdeFSap7vFi86X/pOP/QLHi
DTmf2Ugzgb0ME9nGgiNGV+78++rVbWJo6kHEYiDzW4+tUWrJqyqpdU9spYaaReef
avZEpDdozG7pAobjyqcAZiBhoHsk4+TbVin0Dpi7ypBGt0nTwcgZALHpwDDgwysY
hG4MAkIv4nutTuPF38FCzazk4o+ZXYEBwxmuV+fc2Hy1LTJOckZs3W5wOZDR9eao
aYcxpeJNMvynaLFykFlU5FCEqjG1bJOqzxe0yc9R357cnCvoXVRzfc05JzZqTGSN
WrkrR9KXbuS3hEFrh6Ya+4mf5S2bGNiRP238gN/kE990mRMc9wuDNtv/i2m8prRw
bLdLawkzoOliKlDei15VNeemAMSuOXBOGOSFGivpjCmIPMLJ52fR9KGF2Q68ybqG
VPNXb4JytBpx5AyhdbqHrfiRHy30Gvi3N6jPjme5zZIq7K/HspS9HmbRn2/xlFLC
huPNYRJ6rFGSI7JMhQi5mYtpZmdakhmvOPcMnhnoLsve7qUDbNJleQnrP1BLzvSc
lMsAqGPZ2/bx41iOvuquwY5utXhuhMu0ZY6Z7PjNF9rHH4MCqdu+l2DGO4yy2GAY
vhy5V6W9k/7MAnl574Z7/Bnkp4ETaus99zmRUAvn4+chEtITc8ag7UpucLu/jp3v
2xL693ONDIZlwpqAwzQnuZhS7gKqVME4VnQ0o5/8c4rER4Q37w1oLvPIkkqE/crG
4vdXTuRH00LiQOYIrGGvEl6vvjOjdUbw6khS85bruvKQ+r6nwcOqXEGKACOqfBeM
dsySmLV0RRifWa+rgy1lt06vH4i55t012PuivBnA9eRcTjSaBSJa5yk9ERXrkRWU
aZ8dASL/ydmBHvkBo/S4cexYcv/iNzlG+XyFzsZZ/OOQS18d0qqaiM89Y7TsOTs6
b1HxNv7Oa/nHWiiPITWJx6sHY0LR7KFD4fA0Zif3USE3BtFMYufB9pxXbU9P6RBc
I80uaQhpaVHd9Zj3qDHlWjUyQs7oOssdCGbWnyHd8/0MW0V1fBs6qm08aoFm4dbj
UIQWWUzTYN7NSao3syJF7WqfhTk2TjX3O+gjVJxapH6It4kjz4sb+oCeVrC10AVe
myhq7/k5NwDSyFY1PdWHICo8+yBxGAAQezd+kkN6FVUhuRgYPyh4jMDl64Eq4fO8
8k4nTyyihBe3h/YKEuFhJzYuwi+iKp8I5N/9OWdrnDybIQX12DvbVuZB5gLm+Qb7
WHd3XKRV8gQtP7qogzTfCTXvRSREGpz/kJfFGeH5zTXvGmxRZgV3iu35fgQT8sQs
NLt1+tQGFyOa4gQ6hb1NUvdowGI9SSXiLuQcP4HnHI861TZiBPLbQmgG9LnRRD8o
wE2q8wmyggybOzUkuKTDSdMBJJjjmrtsHkZUfPpAt3L8G4qBhh3BnYAABS4fqIhv
5/eZbf/OmpfU3zvspywrb2g1nz3LMyztf+qMdVOMN5teKf4gppbr1eZXuZCIayTE
4z4mBagan1FTDwgNuxAGqIGpQGangldoxRDE1HYREdlvcfwMzuu/Gln2HmKQL29s
xrBk4oVRd4ZP57BVZNWNjhnPhD7sCnVPMadYe9oOJCDixyr0vsoH/VNPj+gvPUo5
Cji/GERo53JEgcdabyW3OGAFb0Pk9zr3nJT6Jeg98qwXKryTp71FnbCVrQKD0mNc
9+J8bFNFhgAqYH+Vh8sRXSE+0AQHZHLJm+ZiuzsiR3NvE5vOAC6CiWoKyrq8qDAZ
pq4Hdhd0Z232zFieBXXDLKG3tjmONZFyrQDxvhCSzbucP+SjWrL08TgN2LmtZqUH
fRafOV7eW/9t/7mJt09CAw+opN5+qH//Wsz5pGYgJXhC46nXUc5f2m8ZxGNSd1rr
EYfn+fm82jkm7SqmARhwfNVfcJdOCegSelxEPnQ54IeerkdeSqyHtkIck6/O3MV/
2uF/IQalBtpR+LtWdoCO4/+IJ53YjR2ptWWx0ApKpPKm7CW56uKZaFWybcatllvG
TgNue/kTeopyPo93yvHJe0wXudjkRM38+y1MVczZn6erfjx2FDLNqx+Jj8fbZuhE
eWEdlRUJTNjFPVExVfN3CduId/vzVJE3iTyGUuI0zzb1aTeBGJ5pgzBdgNTXvJ3A
eX5CNIFbnEQyeZqZH3A3hwPrhNU0BMTPgnottWDs+8eE+ZNSpHOjLBvM89ID5/18
4n+FYkvWXiHWfTKGCTDpByLOhcfck5OZL9oEpKvaXQQsyLmJicT7Cn3kcDo6q531
lwol6HJPcu84KFaVNty22qW9B0GNw5MA0UgmLsbEZH0+Y6U5+QNjDzK/GBIGIXVR
DEcbTe9KyJ1tXo/l5LVB21U+wINiRGw4evhJxhSwCfecNmU8wteM+TMH9vjXXTok
WRB/LseUv6lAOpIPDS5QcJEft9If1OvPoJ+GkFQ0izGTYvwoNDKhXyKak+FPaiud
nPCB2xe/heGobcji90pwzeQjZlZr/C8EQcayTn6Ys9zGMdrW6UUScFn2hbjmgSlR
SU1soZNBQ2/iMOujvsKrRODTK+GtKpqvFHzHBFN0dVkcxAWP3RBJzFYEotAWkZSO
MjDkpnCmXXMw500ZACpH2FYf4ba/eoxzlA/whOxXFtExUVuk0O5OCIm3WqkmVI1M
HWwpB/84lTrYUq/TPYRgZhDJrPRHgfQOvbxaLgOcks9Zu79w3Mc3Cvh1K+8BKdq/
HUjqivRCQZPFRDEvjSkMZn8BPh7DqFCa6sjgEwxgAtazFZ04Ubn4SvcIIye82z0W
Kuy5i0D7FDCZDzI9j/qreJ/jCZwC7C/aKYnzlYaFDLKQPKx3Y89Y4sZYVzbOO+h1
P56YCacAMCQQ6rcwXqeWF6b7V3cfSim6KnroS79Y5H6HfwPIn1I/BocP+uuvdnea
L14v7BiNmMMmDb3wDRFZowsdG75luVTJC6QnYPxBE1Xk+XUIsKJn2J4Spb3K0bu5
v2MevumLXYK28tujlMCVCT7YU1MC9PWdhocjGTAZjQxsXrNH1Oiqq6lgwyqM7RJL
4ck7kiDEB/XXUMvuTw75dAM2vJfJzLF5IvcqqeLppUuz6AV7PfA3KP4R3Fm21zGA
xiGw33gB6PdPSyPHR/C60rEsiuaP+vVTWrSImLWWLwMIIAxw6SH+NQZ9azvB6zb6
KxU8duHzbxfxvz4Az0fnaNoFm88h/xtI++cw+LDcbGyKzjeD4coLYGp42ByJoP5y
EK8rq8TnBuL2Akl6qndf3H5jyf3Sv68WaxfhDHzH/MVlcPrO9G6w511HijeZePsd
xaaghxYJmrdOTxZXD3YJ5wEUs7P5o/Zl3WzzdaKH72m2f3VlejL1OWEoy7OusG4i
g2891fjyJPilMNsB+Md3KTLwxqiuJzNzYqbYk4XQsUF/XtMyEXt5dspbDEzxcPZu
Cm8STVgxZwk+artm5WTG6RsPbZNZcLpsX1DSClo4i9OnK8i2dPCBqG2snoi2XWaL
yMrrGOb+LiD5Fh3j2T4SvRfXvwj/d8VqSs5Ibb07GXNpaJQvO/gpVVGbMiPi005n
hySlC+9OgE1DAP58YCKCEbWk7f1owFDeMryBjMPEAfLHO+kZ97KMF5npkVjFqN4b
ZBb8lRMv7+GvCBehgPoVxAKFsMG/Dy5u5BR2g3qK3yHgSKCkCfI9RLfUYWbXpFqd
iT2YZtT92v1n3XO85cPilKUtXNnDisS89AzV2bZKX19wHVOk8lUPnYLQt8mAYPoe
3eYuVj5ZZd6309krmqG439bwE/TyawM51bcM9p0HxDFNEWhvOw7U2R8b1U0x5Foy
5XI4/LaFOnI7rThTjN3MsNv5DjcG8M94jXJHfeRJIq/AeroDSDKkAU5yNd07j1Tc
/hV4dyMBpxU+zUqiY9Gkojdp0Umg5IaJo8Po9zZnoh7r1QMA8RTtUSEeyFMBjKPB
DWJd1WiXcYwJLfBojyQZLUz1qlmWHbZWH7RjHxwS++DBjUTeVrKbVeHxlMWJIV6x
l59gsCOa5JuoAIOsr75KSBRVeNuA8+FIFyNiUTXiPEcX7Fc1uQpX8dHtq7XGJnsS
Ux3JkRzC75eSB8lWhBNkkpBHQUVeihETkycJs81D/KwjTFBMZMV3aq3DGAYTxrBh
2Q7quzKj+3cXDTw8xl7IxQxtXfl1OvE/KgA0tWqzjPg5jeeTrE5UJTjonipvFGVO
oSxNcnA06BMF2JeGVQNFFVopvPaT8Taa6+MzRwM+Frm/JBNNxz6XoFqhy8AN7VH/
1UZ4F6MeuDzaGVZXQ0uZ12wK1flZjYGkBKeM+G0frw6OZnam5UpuMTAqJo1MYdzZ
EPkzJ3TcwGKLo3S3ILMNQeBtp146CluXjhbhQyl/i5HeRkNxnzyHVE5h3d4cqOcm
R6ecoYuW41stSSuRo9/QK4QDM72IQLxIULLkUPlbsafSYwIBbRXo0YLIYcheMfYj
+ATSkSMOUW/tpQMl2Ae78JN7d1Gxr6ownPIEeALQbTGnRaPkHJ6SB8yHuTaVOZ4a
2pdHWcw0tI2s02mh+7Z8JAdWKP4SrQNZC3r2qs9yNCKXd3Swp73wWtPmwWHzW1SM
y9W0RTenxiOUvI7bv2WU6YjQRjNXVo0tVOThPppoRq7FL+ziz6/ViRANg4rZTdcS
M07YpUt4Q7AwnoxxbkCYiqBU1/khTCry8sniYvj1ZJHdPLqBqHqH9DnryUJNjIk9
TNEI3kSm8D+/WhMClSyNfnCp6UQMExNGpgtx5G8TID4zgdDltseu8C98tBrgfXjn
QG0FWwxTul/Sz+LWJmPsMp3G4quYNfRmfZGanka1td3tylATYWJiCOulcLpP+GRu
QgZqhgj61HyWo/Vh6bm9M/OyiTvOW6cR7SdLMZ1Fgpocj+ia2Bp0IT8uWdaR7F52
/RbeUvfvfTogjBvPyt0rfO3cUhFQfOELrc1PNk9OI2tMEfWx4U1XQkTlYJ8X47Sf
B1SSsK50WPHIuWNwYgLjDGHqhyPActeCv2sU6t39sMTQzzg9uXP6Pafi0g8bkx/Z
GXZsBQvbpiSKQnAVSQISPyLpjOMiZbQZ1H/Pl6G2oIy35orWMtOjhQYfMMZaSwi6
mtWotB6rEkaNLo47ULgo+DV6Fchi1PkPEKklp5ytVJk8b57dtCAvtgxsQPzsqEZW
WRow9HN5CycnYk/681bbQkjCxwS6PB3dxVnb6Z6nFwe0AnQ1d9lK7kgmVZ18ojjU
wKh+Iwv4O6b8xdnOatS517LItlHlMy1PkQCSkpEMwoGRbcS/qAJfoWd4bKLKEsfa
SAIHixZF4hx3kmw/rE+Q21BqlnSOI2jntf0C/ZtgWjBAyOJl5EqlfYThkpLLdJRh
2dsh/2h7kpRAkr1AIxFQ6l76O0maeI8DI+JDMKkAzB+tPiHNuCKnPQx5xTUspL2O
cvfpdZCBVwZx7tvV9/17gjrX+aPm6cJ4M+r/Y1J+ZY2jIGpW5uXtFzlA2AzJBMIz
9EkoHXtd40HPFdOFnQCpRsq3/QmvPZ1SKRH66UFF4M+DYRHAmIgwflXVk8XDZGFK
mwGoBvD+6vJTt89VP4emxK2tHQGTx/lEQy/j1Q2JvPgxk/pN/IZp3a58I1773dtB
4xSSFgfrz6fGL6bN1Lyat/Wd6KT17TGggUZ8ePfjUjcGputB/dMkYYDWM82xuTVs
/UjJrtfedLMIbcS46DqWWGPPOJf53noa/BEr7ghayKxsI1/vQQnreSkXfACAYKii
3Ls+dgIAy7lDKFqRPE6CHuGTUeMOey4tp1NEFP56HXY4OI6G5y5p5blGA6bW44oR
CbIjUe5LjiZgVqzesjv1fyq94uWJ8I/wohDwJfDp8slgF1BPnT/qzoD183yjB3fk
RsaLWq1P0uchJN7jIWXhgGskwm2PIQNonoOWiuLqGBS6kpsGJkBgJyB2SpTPATrk
ZmsyaStoc2E+1GLpVlTU8FkrDv/bGTlbOcjSO43SL0ZrVLafbKgcczgRi1vtzRHd
nwBiN2bwYGWS2/BlAQVjZVZ1J690duA8ez8wY2Lc4/Br7jBBaEMnLAS8hbaO7YpM
J1TTF+fh7187qAoX80y9Ra2Q137BlQ8sZVO1JiQjcCWbcqNN7KJlDfLEFCxkyg6J
hz1smnhqv6wQ7JOZswyB5FsFkyBDq0I6s3SZoYEaXMuMnXdxIfInTcHOSj5ALQbF
WcaYs9x1vCRxHH1ptMLe5CbxIBzha1Hd9taehYY9bdkHj39K51KfGnngM+Jk9iu4
yxLMUgYcsFZJVOecOCJv1RI7KhXHjh5NLvf9mLW/eJb52J37Syz9eqEQ0BvOUN20
8AQ2Hr+JHN88XySYx0QDmSfcAQjs+xwyw+pRxA52UuiDea26cxMQcZlfdmVwxd6K
MQqwTwaTxkSy+c+yjkT154a6wzVJLKQKFiTP/NOxNOIZoqFvLJo45VX32+75LW+N
F1h4VC+84mbjBG0lZyPqYHjt95RoC/TJ7+to8szQoPx4V7+/XmxXOaUPyo0DeAzf
S4T9K60wCjypaxAk7055ebeldi0xnlk8eGgd6f9MCBEDKdIsrRtHEgwe6Qq3fFl2
yeFYTB7GmcKenyvL7Uvz6jYPc6CvMnXLQSUPF8adXsjac3otQTaKRmzF60Bd1QqD
pujyO8OafuyIf9Y8KliNBSqlEggOK0RiXOHe+CDhhpSAfaO2TOuWgVQzdrtdrlKH
m3H7VfGBZyi8t9/lMqzTUuM2pn45TrWT5PwHkeaGyVifgttWsWQ99dcLDEzON3Wd
/1bCnbr3YFWEWhIEfyTdugo9bgTrVfNdYwXvfGHgkf0Op4kbTUPCIG359+OK9CvG
G6gMDdvCMmItqbKy3KV8GpPN3XAAzRBps5HyZtwPrN9beFyV4siuyYagkU6MEeWT
tnpDnxGGSZCm8m1m1YV+d3mffdOvsn5hjAIToqJJD8ivpLCc7BI3J1F3Psc9gIba
OhIato0fOl8imRM5AY8RahoE+xDPnEE0bE4HuycLf5wwFrKY9Qx8PE5It19CJC4e
jorxOaq3y9zNH62LHmrByHjruvdci1aC1jkn6O0f88pAoFEJPQMX3TBfHoaMqq88
PZAqe/+B4BEXgZbqSOnvcfPYVpX6HKTLgraAgNB+6aKPMFYUuZ9RYfC8xxir1KjS
DVDCWZv1xU2qPRrKL3q91uqEOY/XyVQue7l9HleZPZAQjsJpKZT0b9rU4K2mZj7W
YlQuxzsNAFEC6zNmavFDK+IjHRf3HeflFqWu1mYtAYb+EEL3+94YyqXamDtDJ8lh
D58LB9BHFcBBvi2ik+IEfLwa+2/SNxAMnLeaCjEDYtNmIwPbZY8Q/2jlK8SoMgV1
nOvM7Y+5aXdvxPnxIDBJulQL3LrDfAPwZpuF7wfkFXiS0Udp0W9tcSrM1vLZBcB7
QRnGAUW9SChn8673Uz7pYB0DV5Svb2FpEpkyh8WNWVb4YseEeWVlad7v7V/8xWu8
BjJXEvAtk/7p91Kp7DWHnLTOQXqnZsMcdshQf1ldd1asKKMCSkW64QvC6INsxuz1
H/7M/KpXKPrtH+OaLQLJu/e1c/ZlaU/hRYDqaOMq5kRnT15VXvaP0eF1OYCcbbh9
Qdmk/LhIKPBLRX32oY1Q7pY65UhP8oEu0Q9M1mmXC1eOApEGG1Tqu1TUoyu7prf0
NDAq4CLTq6R/+B/fcrZbUg65cS0qok9aD2b6axrVyH4W1njU4NwgWjvWk74dzMdT
V3peTbruJ3Vcvlkm+51pcQWXS9rYUkokDZ3yyQmmbsFKei3GPfmoCYQbnwR2X3Hg
ibQ2KamKoc7OIkvmYVBnhS+XFV3O2os99ynT1w/XsIEMTW2X7hdDVo3lapiW6d/r
FwHc7qeIoMHMi08pTPSWvxc7L67VDPc7P8RR2S3jXGWUVwUihBw2yRuXS25lSQPj
nSym60prjjS7XNfXg9WueLMlsO/mlSBjOED3bM6QLLXrYF00Nm6Xd7GxVoqEb0pL
6TFad/W1wqj4LPyVOWYJSa4KcsU+LlMpaX8+BvE4mN5eXUb+OBtzHahg5And0uad
MoJGuwHEzUeLMxUuaHHzpgFei9lB+VgyrK6HLxuTrDTHJtzMjXx/A5Y9U2S8r1uP
2ncuBXY9REvvaJiU3qN7RRaR2oN+K6BVSJ6ALh0eVuLf6q6vjlb/XWO4aWq5G9LJ
JRpXSc/XrBr+aw46p+PGSqcYf6VKl1OYDTGgxvG/FUu83NpQIVHthvBu+0XEnKCt
Wh4+2+ZUrG5Jsoe/kG5mbXqVQJAvgmXeRNOqkYPY4f2pi4+7LvEmJ0WeXLfs3fsz
3Av8T9qM/IFMb5NvwDmpHlqVLkgtBIgvTuZqDtrz5CXAO4DxdAk7I3vJpzd1wBwv
1eKKn47HTHM4SOnVQBgXuG8LOYaGhYcsw0VGzv26buTpXXlkqHqu+E6nXgRV3ifw
bvV4hdVfV7JAk35YuqOOLubl1EcWZXzxBQgKNlLLSGmi2N5iJpHz8lpgSvS6PUfK
IaSCEZ7m0QLTXqPWbh8v0Nr/9YPrylHhQ6BPDoQVRknzBbrnw9Fi/soC+JAVzUiP
irD/R8LHgOX6go7QEPT/NNpx5ySeWxsoH33FMEiQ6F/k4SPEujTaGi/l2G72LI2q
C+IFf7e0HEh0wfI5vANLkEEiq7HfGafNE0bPOy8wfxtfVPuZg2baqA17cUQA+paK
036dPF1fosKzKqZvVPY/gvD0a4QMkkN5T5OwiJtNWUnSva5sWE6QiEJpgmeOP2bt
lwyuj/kIzP+xXd72QzBFFRUiN/mXnTd7EmzYsG532yA21gqYEFYbrDUastEvnrdV
OrUtVUfCczsXWKiekDhLIJfxc75wgCLTeUi2jFu0xtNKnIVpamIA4BaJUXBphSFM
sIMNGczYp2E+3MxGnS2JSJozr+uFFQuXhGPUFevKgasWMfb4xNwnP3hLwM35hkA5
Pc7oWY9F+x7gD9WraPs5N9KfocGQjSMCPrCgennfaduwPZfwYoBVG9kr5F2Qgnti
6j8xmdH7v4MYOf+uZeVtV5YmQERxTQoUc++L4WQ1opVDbDthhWSWoI5D60GcACkS
fLDAvb/vF5yzT8uU2gd4EfaLH9rg8qdciYq4m5cCqRWuwxxIH4fhSWURkYH7TrTJ
URdc+UqFJWEpEfE2x9OBz1KUfvFxhZpxpGvI6RiwC5U8tEHQTTqpe5m1hJqns+kD
qGKbSOQSEuEy4RNnfclKgs3/xHzIekGEmsFmV94sQKSiviYayS2cvuhsgmZ21yzO
E8PN/E1e7AUC9AuxuRPsIqU2IUIGWvbGz9paXg/PzoTlaRY51W9sm5PiVOwNNPDu
QplWX/qOux/C/I17qyjKncwo2w9AU8w2Oz6ai/ZHuFPHoE+HEjWIxfaBWKr8K1Ts
KhFBMxWr/WIu+JXJcHf65kjFMilmw0ECP1WKK9SuY5nMpzUuKBAdCXZMaENy47R6
Mmd6ZbF+8eI8MVUCuXtc50rLt8UHh8OlQnEoYTlTFA/mtHkzLOv2bbx2yrtef0JK
+1Nv2FtxEIolquE4cpba308Lfy3NYidzicE/WF0HKGAiBcOXC8xwedHfTLnWxyKn
aql4htI0PmXMdMhwKMphEZ6TGFKEZEPJT4/cfc94WZbKKMCfL6as/qA1D/8fxwxR
EC63xrjNQAQy0IUc30+tCG6my+bnvTosBlXRAXs5nKSPn+EqI6Sxp0AVr6JldRCR
DVJ69sAXYaVi3x10Idi+Vqzb3QycEaRRnqMgcApXc/+S37rYtyPRlKo4jifEZcKU
bjl+xh27eTxIpIccPwWx0itC8h/IlZhbKDM1wqM+hvPRl3LpB2YPxuDp+0GRZDH8
2auFTlH9OUNtc+kWCwXY7/GH/4BFNMubAQyvaIOL3dR1MjOJ0cHmmuAwuRYd6/b/
S1Jpeb7dXwaByMP4N4dnilRb6QmzKkTTy/fFQWHB6LCD8iPCALsMMOnF9NHV/+Dd
0+bYO0MyEzmRvLLeg6EU6pqQWH04/KlWLG6zQRsxOEjuY/eX/PVB/WUWKxFNw468
eulsLbPyzZfMhEuxfpEPx3HIli8eL6sjAJ8NU35rwWEQcisZbAubTOYB3GPEE/op
r5o4DGTyDAEaFPctRX6782W74j+e6NZ9d6SAQvj0HzrENWLlfDdwCiFbYOmKS5xh
SqYb2eGkiTR/1Pa2//WFFSdo9IqCdhnyJpQD1SpnuZogF7dhKwxjeXhiT/Otm9+k
nd3Xf/atERuR4WTTi7fP/O/bDqYAg6X1S2N0j1Fs/A+FkIai//IEr3OUgdW4xeL8
V0xzJNVuP19RN+woUY67Zo7nGr1SUYb0oHt2ZOwmJQTNhE1ij7ViyNDy2s/F01sN
W2LqoqCXQpgJRDApPOemS7c3DH9HXwcKzQbdCcMYHNCdki8wEEWuEL/20UhUa0kl
0GOeVwvRCr2gF51rrWxX+fALEmEqillQw3BoAPci1IXY0WFdhBcAZW22xwK+pswT
C1yIuv5YthhCz/9xxMvG3NQoXNxiYPvKCKxM05cakzV1Ky6BSMD+diqEK7stynVl
ZU5hFN7Peschuf95YXAK9AlD/uqN8pLiPZV85ELvjv1mU1Xgdqb8RD5EPpx/cuva
RKyUx8VqmPRhgIR0BpHq1TyyJbFS+m+UKHXlju0ghkBYCJNyBN8qyojWSP9cJxOy
McWDQTlDPxb8wjDJpc0mJFGXS7hmL73JeCGNaGM42rEGBv2YNek5NMkm6ii7e7fD
NyrzFmRwTG5JVN0bZSohiooQJzolV+ZP4uH7/F8bzK1by35FqInU6WFtcuHkF3a/
mMd2WMi/oLUoNAuZs2W/+9RTtZbjJrs6OCVOytpvgLpqk98lemQe6r8BDjdqvjBQ
CLjNbj28mBDig2eY3uQPMOFxV//2aKIvTalNplA+4dQSeKz+oPTWYaDAo8ijKeyN
RkVysRMUx7v8N4FObUPskkEZK8yhulctHsj4aAaRLamXCUbfhQ1UqdHLa3shS1cm
htxq3ZuqJ4ERZz4glFT1ts8e/jLjXafLttEjMj5hxM93wx2mV8IiG8XWJ6LU5+pd
fyCFGaU+cJD1UlfwqcBY4h6Gm4kUsScZbdFo3pOT3+0P5PmEJecU1o5P+n8oHA4C
aa0RfS9oY9eXJqTIt++OY6/NnO7ilPpCTx0eoO5CWJLc1hv64gLE08EjNwXbOT2u
nxh8wCzr7hpDt/bHmfIwlk83wCi+tg+bBzhYEIfkITD14o0KveD2kWmAbG8IlmDr
LehhnqteMzIqpnWtXWgXBaGfGyj8fUOrdnLkcgfAa3fk8OilVOsNOe9++2VMvWXb
sgHRJHAyAeO6TqZBwqtG8T9lsEx9v4QtGTU4zPvlWuHjnMkB3rJN7i/ktC5FLr/I
IeNFX8X44x6b1pmDOSy6DrTOmSg1OzoV+Tc0j/pJfLonAiRFUlCgbkI1TsHNnork
WqdcsmIRf1pHZSA14wvY2bFuckvwAIPhaLgUvQdNwSv/JV8D/L288MnB9LmBWE8X
m/UyBexQQhlVOlV1PBYqJdUt/eJwzIpv1QqkojZNupv0uuHPjZtuXerumkkSFAwB
VV/W8nH+8ISod5hIDC8vmyZ3lj+DZXf3+fJ//L96wPgrcl9RiMLaprBHwL3rLoP1
he0cwIlpDeSbo4JErvVmFA14qdQ42kAbrMtIVIl69N4BO2jcrjuXkQUazcTNEey2
refURguhj3CokbhYZdyLKIcJBGSmiKXDl/Ev3wNjjBtbTFfiVi1EYOK1yDF+VDL5
q9K+TChAIbdWbSIgu5ViqkdVrPNH483dIKauv2fn1DqxKFLOsHiStpieKw+4BeAf
nw8pr/UzBPUqOp+GIHAhdUNgjU9oJ+LadxuvJpcWBWwEjuGDwyjDUaCxBnM9vnb1
Au7Wh4+Z0EodriryTAg/1YWnET/SOPTLBxgiAq71oujuqzHL5X2+w7PfbT+X+dQ6
YVe7HEJI8g3g7+SaA3FZnik4JJ/otLm91/vlszosc7DoVVmmFFHrHF+5rfljlGFe
ayVoceQLkf/GlmHotGFHas5iWP1zUJPHFj1/LnLc4pStLXxXc2X0lcFBU/DUsjzD
9fA2ZSjqj4t42Qv3vlMcZ9IHwGMzQZDmmzFIdWqy77ha/sXM9pU4uWmUC8qoLEkM
HzvQ6Vx5X7uniAddLLov5PlQvHQ4WkhfYYwMTmNqOZ/2tDtLI5n6lu9JOq+TMRa+
v4MR5sjHpX9yLQ/XWf98NCp+qnyH5vLDRmnNgGKnpW/MtqNvvgGYD4V5Z3XSXgxe
AxLzgz2AHHs/8m0OyD+p44T0AJP5vkxpxKlu2ZOxWordsvmvKBbUH/mbPc8GvpwM
5o8HqWL0d/eQTcNlUG9AZaE/CWIZ6tj0Sx1mtLa5Ka8n33ag7U5m6YsVJpDy0ZhT
KtFC3Jxyyj5WlOBnQqCg3tZIuoXM+RPuI83D10rlJ+sLq4nj6OTayXqjk6zAFxho
f+3O8hDnZGoGdF3k4uLfxNfDSeQBV5TXVNdxj38+PuIYlQ+4dzg5KyPg3QzHwhkp
U7pSYW6itr/rcHo75RqOMXs0/vVNfsQWt1ui7ZVQF+/Se9dGvGIlSSU0BYXxr/bm
erajTe7jtU0GdIT1bLFullHko8FAw2xx69C36YJVebf1DoUKPfLzXJ2yYY/4UXEN
SI3yuA3bxbE3cJikOPB9QPNbElWuugPy86dURjI1TrqTnf1Vebq4c+LN0Y+mkgto
wiOKA4HZ68o0Mk7qu9MByW4+wYxSns5hcZcTRxoVIy4gKarSxSVNhu7NmZBIBclj
N6qJJdegVOQcks5MFc10QUo/n6FhcsXJSq9I4W4znXnkTR43Sst/d9bEXzGkxptk
gLmm7+EBsOHV9mO7vsENIyWFZu/k20S/wDNPN8IH+tEw90wu7YwuXvOARB5k+Hik
PIuEU7+jlf85v7N/lmfibIZamgUBtYBfBVIYfvrRnp9UBx5RrdVdXr4gdVwBSeHF
6u8BymrNVq1yDBlSfZ+fbQC3DlPsoCPsBTk00MecxRPHzNlQFqrpb95VnENbzv6j
rhh/Pj1F55VoPTSixRrSSNMnCdcYPyAD9jerXmeg6X6INlRZzck8G6WxPFkDM/S0
rcpj4956+YftNT25bA8YqGogm7f9DINo13Hqbj+sY7CxNrn7tBPYki1p9iZqGpLL
caMy/ajezZ+lmpQdd32m24vR8p27CITYE1VFr46oo9TRtlsgQ3Y4Ax2uEskQCWwU
d72vvUVc/cBzMJr1+98u34ovudfJ7ZhX7NoV0B5QkOit97zNt2v+c5HMwGztmTou
ruutF9zH8FHOLgT7vHQltSHyrx8Y/eJHpqDd/YXNZxvZHxA08Hh5GvLlg6INNfWf
ERNC1/fUbRAvmwf76+T6EP8sChUcYXyg2k6O40jYaSg5uYag74qFPtKMC/7HsLGr
QEzDCi5cub4OCyDlxSIak4C6wiEOMYLh33Kbvy/oEzHjaQeHOf/ycdQ3EBC/1kQA
YMagxJL/WccQVg77SdNceLF0NBlTIsXtUrDndqbrTbBDtFq9NPpQctfPiqnZQtiQ
Xzjlx5CWoQqUday7EkG6oX6qF3MCm6sFGoflSRSGS2crjLImCPNkW6yLAt7gDfth
ieSGqQIVyNUBqruGmB3yMH6sunHkJiya20Ngw+KVGHuPt8hQtE7l12iOXPvDcJo2
/BvG9mqziqVr2ZRFjycm4t6w4SKhOe/XzJ85vOf0u8vo3HY7k1IDf33V5IeRPJ+C
uURtTPWxnI5xnU7KZaoZJVaBQFkI8ZHcLJ/XxU8HukmI7c3ZyMJuQveQsUAZ5PKs
xc1YhZLMuVg1P9RXdMCSdhpegXAIVm47IV03JpfBNIUdRXkpminQunfYn6D2vvZa
DEdF32Fxlo2MsHBRqT8a+TfGdT/q5OK/s/jE9loNVvVMQ11pd5Qpg4oFVhZRjaFL
AccCr616VFw7/Zok1Dvxh89mmHj9vNSQ1OG+c2QajY6SUXy20JYXMYVynZQChYAo
eEUr/IF7Uau2yqMu4F/iKorTEhwFjw7ojgtcWzUUQoY1vyxB8cB5Cts94I7CYO6N
iSoIzhbdF+BxsjEhzMo6QZ5ZktODgLMs4j9J6d4E6vgOEnIjPZV7o9QjmMc465ox
g+YD65hNHixxQZNkP7K8YXWipj6fhQ5w+EeHog+ZQgzZMX2IpVPE6bemF5+SqJ8N
VbzVcuo0D6pFmQpR9S/fysfDpAUn3AOgDITD+FgW9/Kybwj4ECM2OTrDRvFsXHrD
ZXHzzu/Pc7lF+ImylbuD+WxiVd3xM4J2xfiXSVDVsm1Mwd+ogR7Lj1abudjRnOA2
0ZoQX7aH/Zc+YyTDSqypE+8uYIFm5JluUl/wGhwKNmfeQBx8VEf6yvxh33LMFOty
bLirhvAgM6tFf31ZQXumgbxh1LMb2CxCLGp/j6RVZzSB6gJ2qto3LfvmyapKFjQX
AeReD1JqkmkvPlh4EZ21yFwT+0c5PP2MnpyTi3r3syrfC/0xNr8wnPNe18/740SB
obNdhj+1hQzID3g9yxIJsNg4zcQL/ZwnFivgGpM/zm6LsFGTQMKt0MvJvOpGMAuQ
GbLTQQTx7jVxQNFqQQhQ8qwFwBmLReheRUi3UjAJAqvlluBTTTPHdOZIU8MzSPFD
e65Z5SOJ1BbfE6b3gQiWidvGc7IL8dd54NFgoRuPbo+QAutwEV8ego9iyhwLddT6
bUC6bDdMFfUjvaHXzwdCB+k8kxz+BJxK64UBSB7RGQC2l0w7m+OS7+LAwOvjk8fQ
RWldJWaBfN5xnXocYRty1aJEv1AVaoa85i1K085Nl8eh2jE56PR5Hg1v8rfybMf8
xXcEau1VMkvJwOFQ29siP+s+++AtYvpKX5P4Z9sJ4BSL9G4rTdxO0f3ilLvXi6Gt
sMxODYAumRi3iAJz4vw9fsv5DAWeIVm9Y4wXltpdW4oupzk/y0MpHkz4w/racDic
G+9tX/TFSoiG/Ov3P2HMtjpq4r7xraFRaRFWpAdG6LM7cK9UI6d8CdSxKmJbSpab
ecuHgMz/zA0SQT/XUxNGB73Ops6OPqKu38AvD3wrVr4yaXQTc2rXYnXXMrA2hnUD
IhDKsL8eo5LDZG8LrrfzVUUkVhpRASIfPtngQo5JclsJk/2oRbPuxBmXdAborM3X
DNDe25f+1WScXnvE9chVk7tPw5lgsFB6S/E+S+KLVODtuTGnAiu/kRQt/ijEBXoH
KIqnAo3c4qdbyY8k74W9Qy5ZLVqK/9e+mbAIDvpwEovPkMOH6MUuc9+QCnKKUesH
nMtUsfNsdg/sby7BjoUFiieIxDIpdKQjVgJC9DqtQsz0pQRoAK26C4nzAkJQXC4F
yBwXMfhC8VcE9sdCduQvzjODVI4kVrfamWjbwtGPRAkK0sDKXD0m+t1UbFLzcbN0
VCYnoqmhsGNzsu7PAEJGlzSLBK/0MfRZfKBStnE9wbo9CJ7IH5ZJFIHgJcx7DF6b
4IkP5sQPuYsM+2w1/XsTEsbeoV/Ybi8kP3n1XRm4oOEIAS7G8IB+WZq3A+4hPWcW
px6xFMB17a53kIBkiir5PKOpEFznvVcKE6BKh7ThEmsBwBPaLEYJSkGfMSkqgSKh
nVgSQBR7r4Xe2qcF/2OQsMFiokRfz0tRzFzm9vseL7+gu4uQPkL6l/o9kAe+rVbj
uMDY6rLSsJ7o9W/A2LAeLtsByRFlr4qw4xLMf0Sa2615OdJUKmxzpuFSnuxcHiRI
WudFz5hX+T4RoJH9zNUVyrQGX5TEFgVQeOsK0LvsZYmceq+Ol+f2paBY51bUOHic
mDbbtXcDVa/lDdj1jFnv56TfessNYO5fQotI9CDC/ErsUY6XXuEAEDNQ/wi5IOIK
bgOvcXi8xzwjNMYIJFKXLZUihBQufD1NqGYWl+H/WDn1C0BxRUe5eVgwPu27YruF
zv6ejRa5VX68zDiEZPxF7nsTEqZ2UcQE1JrEIX7J+esYb8/uEACAD13ytqKLlxS9
5OuC1mN+NO4LjHK+iibrodof+du4ya5ZA2umRjpZwXaUCB/DnWKReP1RHq+91UiW
HpUAWwP7uEoEum/7Pp1QfLb7VPqjz8tsc/oT+dgxUsgGXhVwIMh50wRJYLbRuA4Z
60Zvb8fQ3msuADmZHLKP9QvkKC849FvucKRZhSgGQFsVo4807W5nkxdf6STbzhtI
lCAv4VL9bicxtfOKXNhYMPc1XyleZMx+9df77aAMGf7EbRWA1Exo0vWh0wF/2V6I
W1GVGoO4Ptb2MgNrEDyKT88gjAy/qMrdT/CJH7Y7NQdG15aPEnSSs4Keg9tKAo4S
eTt2EreeY1oqDzAGQkQYN80sISy6AYDORA+xDs+ZefEw6iZN747WOlotS3yKDNQg
qkfsgOHibaRP8U8KhTmvvTjMbCro4DV4mh7NXhwy0ZgAHq+KY1Xs9hfdHIwhLzMD
XoY2fBBX2Nyi5reODVF636yio1zlIDREzmJkCfQwIKLFD4y7riv4SKijKpUd/+61
srfrWeaxf2hmX600ONWBhySz8CQf91dQhBGSzYZHsHJoSx5E2fUeF1DlVpQL+3YN
W6isSmCPCL9CZBYGDd6Zt4KngXN6RxdJ+XSSKbGsrVeVL7C3Wwon9zfhyW/OlvFy
LgQHref07PPpTtjWWmBz2jlW7vj0S2LxrPAm7aY/8J08J+1jAtWIs4Pq9+3qTwwe
aNCZOIGfB9HfLA+gDbDGg4zWGy02M+UVzQZqDzJznawgUArAtzYf8BmiRXDYTgWc
nLkYhqhF9V+AsnDoqt4b4yT+BZrBkGyF7FovMUALZ8Zrycbnf8+6eo7VFKFtDXfw
rN5tFYbZsdTzIEZHgXZoFILxdV8Bl1jV9yvh/zhK2yuAAHs8hb20LL/jJdKviq3I
avlzPGDZ0r7kWSIpnKc4Uzwxy0na3ctM4uFwIrGntAtEEqM6xzdskck69+rDqCpg
Yks10juol8ttmxpakoHAcRH2Q3GkEo+aBYu/XGd98tvx4mtj6MGYHvTCcFn1e0I5
HElS+PI2RTq4wRZZWWhSwaMI+8pe09UAL4zRd1G0/rqLflUctWLotyQDc3BWSa5M
0EkOYETZCvkgEFVP9VqWU6DolD0qc4to7cGZiItTXHCUPROCHqsfPLFB987rCpAd
wopy6nwA4Bcoz+zeRUATlc3J1TEraPXA63EgqaqdqM+2rC6H6OeXJSarpCHK2yCf
ySupMXRIBAASp/atF+RQ9xsBl4Fpif1hrXoJ2gq8WpO4yeo9JyBqEdVEaGGETAaL
9wPEFhv6+NKMZWtKmmNKAhqL9kY8HI6MPAMwhXO0D3M9SUWZUfwHNiWbGlnnODFH
p58swTSkBPCSw1kSm24xqKXfIlq0EkIOtNLE1FfEuRC7oeQnrEaa6+98YhiK6r9k
ZLhr6WYrkty6nIPKwc6A62gi8SGin5ApXPmSm1Js7MMWZv+ZLtFgoSkUjE1NA+qJ
cGRVD0sePXAJShZ3FyLlykvtI4x665LQh9BpHttDQm4nR47FuakHhe0pFek+4JVe
8PO/B4JKnSo3nPIAj7TGMUjRr7b+dKs4WDzZw9eiRLBeV2M60vA4L4BG200W5dLw
wx8X8onfCD8ywNrE/nJlpolZVyjZAx7DjSc0tfkfy0S0Mz3VCdBXIN2S5ofY6ivN
tKQuCeXKiC+GY56Asv8LcTRxAZorRXuUuI9+87iUsn2a+yAyY4ECAmqsyB5J8UnX
Y+hMmjb0Qu0XcN97njqdCm5zfiW9kZfyaThNR3bFmUawlCaH8NJztJc9ZQojn1rf
KJS/6BTngibfxsSnMU641HpgqCIX+poric59HOTW/Bwo6UonCviDdKC5gd7SNcTw
/soTqicYmMubJH5CJr2cAo+r2HzZESjmzoEp39lC+t7iHxCgcaJmk26CjRUPyFFp
e3ZH1I99/u75+ySxm+/9cqU0pN/khv7w40V99M6+Rf7EW2HnxuqI6PqwSFz6Flna
aYdA/UTMFOT63Of65ZN2ruknuwFu2mzftMriWnfl7GETyTcaJ2mMrsDnhqhleqf/
2FCt2krj/J8OIinKI46HZJB8z8dToYWKt55eyvwRWwUqcUEhRJvHXp+Ag080UoKw
MCKIlHpW32HJv9r3yApp+KkO49Wz+jQuKU9FZt8RWFJrywswDdeUEqnlXmLwMEwS
ylgpV7DnTbkZTxwABxdn9yRewbyFOjzaowDq9RCEca3X7oJP2sdSKMhogLUwYPfb
DqfsnKjddngjjy4/cQe0cmSTaGTG438zdRPuHo8MKlKOtuvokfZA+x/JVNNcT9id
/7bTatcLcjRgAujeHo2uLFREbtqcTxb2MWcswsPN21srBwHQ0JjD03ZVSvum4Kgz
uunGZHPZ11CkgtPYXc5R6Kf9sU2wRsNYAo02H7113bUkqcGZCMPf2nuykEPeqVv3
cbl2cPISzYbxlmPRj8u2GfXcaOMHXyU0FMj8LvFSQzCe+IZhiLfngula34LnJR2e
eHxFSWVd/i7WCgLlyNxIsMBL1ftdhpUaFQFYTehzsl4SfHjfIxnP46nIznbmUyuo
ydjjKLDTcYeJjRDFsUMAzS/2JnNBzB3SReFF00YkTHnRq3HmqwYWRdFE8+ioc8/b
Vjh8f8pzYeR1ONJ063kruvXoBdiYWt224yGhY3CJZSintMtvIICGJi3LSa/4sf5T
JPCH7SSscri5nuNkDPN7y2byx73/PFB/ZqhjiCIz/WTJXr8zNfdUvRnvSkhZzRbP
LurSWs1eaTjpEo/DCE1DQTk83Z+fgokhVj6SizKZZtZCeRfoPIpNnoVXQKPGqvwV
RWjWIuhUX2TuN01guUy6ujZZ0txL2S51NMR598iiX1U19qWE08DzFMu7AFa7KSge
buB0RgM0c23WW29RPduZIZw94BqzBn3XEOw9UTD0eSfKS9AivIHbblP5T7zXjXUg
iNXRZX09K4yYGWIbt+xFy5UZ1toGOHtb3wWPhEJFdRQDUX4EdEsS1OIVwmldWQ6U
yVu77I+aXxIinodes5UN2lvGe85XlkNclGtc8y7Wc0qOKQUoH+L+GAUHVt64P1Sy
nTrJ4mdQSFz2NlxMBNXtrIN8QTXDevQE9VrFGina987FK3J7qphNuQCiQWy0zaUu
D7EsIPFWYIpxGT9qVLsJrmEsjN5jYK0anrAki52YDKREs9Rf4A34FvGW2I6ipT1p
UPAouYtRLxJHxBr41NUUSdbxBdrqR2yFe40k6VZ/3UKby38bKPRlic1m5U776UXI
cClBpBYIpNyV4KQUZBtom4vSWfdb0esBwhsGV/PwyFn3ReLpQfWJH6xb8/Vp/W8a
a7dfRDfnMSBO5W+iCx71Ymv7akd1thnjoAEvNwqXY+CIyV1JuTO/26u0nIDDHroy
TT5hWFoj/smN3lH78Us7JS6aHARxfUvzd3n+qUnR18GxmOAdZrGVblBuq8rb2g3H
4xE16jlZU7q0vUc5Lz+Oiq/vfI73krEaFSs9tKybeYXvBnnxHW2Cl8+MPfl59Jmj
9op3xUaFA4Z35y8liIV6XCw4nq/z4eFEiv0CIB1DHKsSP28siFSb5hWLZPBWpocM
cu273MxF5PH0x8D7ONPrxArSB1O1UM/NuPh54uJtkb5G9FPY/0YaBewStPQLDUfg
IfSxnH7G952e9j9n7P9VEW4x+aNZdliwnRWKho/xHPmcwW1CSJe1eCGcQl9ah2yY
0iTx54aOWX4XGY+nce5+BX/rsY3XkZBle2WafRzcyzy5o2kBEYtlITyowm9jw/1d
CZW6rHZgcqe5VDA2Hi8G41fFfdCH9ain1aCwf6kOagl858l7rT6HI6nxncKDMAqF
jKXWLeEOJ76bTk1hhL1KA0N5eji+yL5Q0nz14eUZdJg3dtuhfCl0+WtEMyLrjICe
laiVgIyiQwo3TucCdAJjL1o6UdzNpYOBezw+xJVJdpX5D+Bfz+V/3qprsYDOvB+Z
EgsIL4V2qJ8130MAhi6I0o72k98L0rYCLkrb859fA/g65/EArMXmvPQzaILBW2Ek
2hX814Wlihf+MgqQKclbtQkNKt7jrR1BcrxTFu4d2HF8Bz68ztRLTI1kVGu0ZpYd
gRvAnXvRZGVPI/JaZwagTmkrEzHnfn1YqLHv9rM9lNtZPE0LXsk+D2E5lzVBN37v
XeYgkwHxFkU00pSy9IP3o0VVl9GtrZUqilFdtxl5F1RvLr0yjX6cIbTvIuXUOA2g
FBXs8pMIxX4Vhz44x0hSrsuBo03nVV12BrAx4bV7q45Zq034+7HIP4s6Zpw2x3XH
BuCBgz8Qz766UnNrIZlccZkzkizPF3iOLidTjg0ke2HWpeRUBWtgmYFtprm8KY9A
/8s7EsrM2g1vqRjG4cnMkhGSuPGrNg4ePCFqJy+4jcvfjp+Borg8SjqNR17AsVVS
Ine405PrGx8sNbLBatXcKdIH7H762BZAUC/0Q6Jlw8S2XaOKhiYii+u9WieaZ06O
wFWjlMA5a4Q8Dl/rcC4Z7tZA6R03scWG6kFYzMtmMmBGdql/qbcxsD5+4eeOBwJ6
MU4xvxem3AaRyEkdIL8s1yQW3XpKSbKiVnKoFMiGcMqgZXK5h2b5XWkgevT4jvKY
VnrTp4FPMWoHe//9HJwP1MuDAGqDb9m7q9aR3Jnhs0SU8OImNmJHIKAU5lW+BjIz
EwpR6NALL+wOrpdTAgZa1uTSvDOWq3+dcZMskPEYeH06HG8YWNz/u8Acn1lckx47
A4a+sieRP9eLoc/YuJGJeorsgH1VVV/HtHnOfpYpGrz+niS5xx73L6ZsAvmhtHz+
NkefW0zDBKujHPw56m5yFhzHsddj9gfLcs5mEA/NpWANYPeSlnFHVv/xTjDt3yvn
kHys5ynrJ/8hPJq7dDuAJ7rFRzBVZvWbAy4f0Iipr4eAYf+5MMFDFsGYZH2Zc5lx
qEbmbj439P24iBRVsG5xogWWz1tey9y4cv/Y0wrQF0KDR/i3ewmCjulXSF1qog7D
Xe4TjNSQcR/39qumEIXPiofs3EbzbeQQjX4gybY79uvelDDWCloypQNqE3xnC0xZ
LyfYrenVHxgahEkdR8nCfRpq26VlPyO4EQB5mgjsIU2G6UAF/g/IH1aCrzeUITRr
554cc8TsjLwTXYeeJk6a/fmOB7qvj/i2neDszoyoqCvIXmkDtH2mVu/dESPfDotW
pFnNRGBmJgqJVgBcOjj96O88EGxiRw/sX2vSQFfm7UE1V2aMjVJolWw8NUjbZ9UY
OrEEOcvrwffzs2ZYuQzP4ag/f8NMOBER8b24T3FUYTODs0whrzzpinTBArTzQDHs
EEcXelS/HI52UKfmSgk5gHT3RsMiHZnpAGZ2RK1Xt+4KzNIiAVIRi6W5e50XobM/
tbwMxRiAqcGAmIhDnkoBRabXKv4T2pqwT+bMquXo7Yh30AxXIqwiUbZvmbtyj1gZ
YnsmsJQ5FVIr9p73fL7q3X1Bg8VVUL6T+/axy/s+FATVxiyWTXBCSuFvZh+J2Ciz
gs5JggYwJ3Mm9ndw+/EMLi9f57Kh0GRAFtN8qG8zHKjc13ZwScdJrixqKeAT45No
Xcw1sRij2IClWMyngmvffA/weGziofM1nd74AyVmpEZGmkwHp76PVm8BT3hWebh/
vN1pxSTgcGcMhETLMNCKL/Klu1m/t6PHMtEFtcWAouWC7uHrtwBpJYM/ic6NSxnb
Q8eVReanKRr2O1w+GqGGrO3ZZy3xriwLzZHc2HZeShbgMvKyRkbT1evRpBT5lw8P
xga1TO3ZJDY4SXFyZE6dQCGIUVhbJnZ10YpJYldvHzjMUP4FXWS9ouTBl2YfJwOZ
X9ps85lC79v3+VUy61ebw23Myn0Ko3Yo0kuGaYHS6jm0F9liMS5j/g1betJwlf8O
38dJ1othRH330khIq9bOTKm/qdOPckSgNq5vfGyrYpL7E0aQAKhB24ovsIrn0/ho
xfNpdZV2RYF21G7peOlpaWSl5P6dzaemRt9RuOqXpeadg+ajKKiMSsbZAopRiP93
u/zT1A8S8VyuTKM1cGYcNxIdUvBzzVoQ8ckTJacY1r30Qb+Z8IRltewpCPaeImSw
ocfr60XaIOsAMWwj6t6aj5riHEE8zMV9yHrldY1KouPm6xei4l6FYchY2NcFxjDx
YgyoRzfssYlCEw8fCCRsCqFVXxEynClA4sCqIsbB4I/QWqu+FS5E3Ks+WzhxC/EA
nqA2kTB6TQlhJiIpYsHXaMDAMc2jjCtYp9vU1rQ9rxRJrK/xVJwo/Wtv7oUvYQ51
7C7G+VKz27nT94NFwUL9wlnCJ9imRtU21q7WjpgTpn05rl6GqROv1q2dR1TnpCAN
TUm7lmBiAoiDHxLdyyaf5m8/pr+nRG3OKBpirGNskSRKe8Lb4E1QiTls8p4sO1ih
LxYQ1KwVc5btKuWgN24tMkNAwrY317rlL/j8kAoqdhM6hHq7XyJrr4PSwSrv0or0
MZfluFBz/ydytpuUsKIkSKVFtwHpp4CuDA7vFIcyjU2od1g32j+dCqwW2BRS3ym2
K8H5TPqejMAbj5vOgmRawURb4TuJ006xBhqFmyh4t87L/crWLSPtJ0kEAvAvnX+u
KUQsyuPKqynsY8jV6ThoCxeZOlzh4ONLAuSXbWJj3Yq8tnaL2eDiDRml3DP3ES39
5AJQw7KjULk1OLg0ErpCmWh1cTXBoIJqv8GS+8tEUMriFJG7L1VpJXqt0zHCyYk/
xRjX7+vNFIotMGRyL+0EUqNmX6n+6mXMpv96nWyOeTSg0wNFuXKzvNG9ico2gA4x
pzjFaW9pQgvFC1fk29oLVclraWd1J571TKWZ5WLT7mEBdInnTfddiChjw6LQ4rc3
fuyWPDAYWN9FiUNG45Q3qnhFadMaAABxaoYv27WSbJOHzishM3wk3xi/3dl/DoH7
S3md8iWKvtAAJ9WDBtUNWNVJ94widW2OCecsIF48qHuyoNH63JtTORnSU5WxVqgA
r4DKgVrdlhLHhqshQZMrCcMLurQei0jCL4gMWYCdK5lQ+zr5Z6+BUQO0CWhiEVs6
PVv9IPSnYytWfyEPZjumu9eK8yZ+NBPPx/CNfuAB+YQ4Z6Jv8xwf2xN0mgJjT3se
EcWzxCTBildTu0zX5Py5hVFuJaE5Ra6jBjrNK6dfMRY/MKFWjhEhFCt07SdxyM7S
EOKzrV5nNZo6tTzAxFHjKbkFOibReewxqqlS1a0NQ/O3DP7iZh/YpRolQotBaSza
bvwZidEE+SJR4MGO86LWKQFYXh8atTduQHIYyc7R2loNjklZw52Ph/UuyK4eSkt5
8qvFXQAGEio/AhrzyOtW+RQeKgUawS6eUpNKCTqQ7pgQRLrAN4ofB4ecYgLNnPGr
a9d49zH8bMj8XS2Ydd31F+5pyggBzQycwq385QajX5b1Og+nZufVl8HewCNsJCgk
tCP36ydLPz0M99vodLS2tWVJMD4qtUQZPSn/VydqKOR2du/vyqkbH2x5HT1YlGs9
mN0rpDyBL8+clqq7i3wELSJFjpsGgcSiav4CH87K0E8SVkGr/Ms2XY4Y7kVPZxMc
0ig7erVjBTVcGrXksQ/B9nVkaC5vBYroewvRLJMq+dKrnpoPEih+GbgkUzWtm5NE
Rk9w8wH9aNOQVISD/mJADtILKyiuxhNFVAZExB542FEIojQJE7x87ysf78gcGelw
3N5yp0Tc2RzwBIW2ESHAq8nS3ZkLKeEFd2+8J9sYndn/FgdykSjWsFdeHJozLUk4
EtSAF31kErkRVJQQzGuKJXq3QfWq6ri+im52SszGKM43/WrLhQk4c309nJlrrMjD
Q5gYhP6KsUf+3twqYw5QZd+oCyB1Jj2Dkwlu6gvn8wgPl92K9wOXVbbQpiQ+zqvS
cKFGuzkGRkALp9GxEbwq6pNhjCGfzj+o29PyMmQpcOYuexmOwd/uGYkLFMGM3Tzs
r8MyIA2Wq/pbuwaLV1ycgbIPoAnWbsbaWaqWVJzfcXSHEt1guHGBxX5Z8BDyVREc
r4ZH+4m5zbsNOVxSTJOUvRWhpPccwVfJQM4BbYI+fW3YEppAsST5iQX2VwLJjDDe
H/JhY3dngAzOa5pJLQZxGjumw0t8i4vsu22cDLce/Irb2pNkokZ264npuJj7X8EG
79jIdQLl6f4RC0j/4m5QZBCB8QBRn3ZMGsD+gNgbfigGbxrnBwx+9iAYLjvvfgti
BjR9SoQODs4TSMweAgZIWRZznVqDpnNqhLpbicD3X35TgredmSyx9+FkKw716Cts
IZA/jreTtdaZhvcMhOWZbI7d+sNaC0Jw/IxggiZbXcrxge83ZtjhNcWuRUGDAtb6
WNyj2vBs7h4WBcjYsWLgXZhIKOBeIQ3o8j7gA6QEsrzVjE/MquEYiuVMJRkl2ewQ
S9/q2TqiInv/kWlCoL5CDA07vy2sBT3wCYlZlTsTaZLBwnw1tJJFkB4pZFK0hkCr
xVrjVkl/+3ADRq4Xa3duzhZ5P77aHunz2bBUUPuSld4opbzPai/VYa1OepyX/owp
CUMP3gd6bOdTT4Lt8eMzPFZFoz4YAm9AZ4XG7HyJs/QyX8oPKvWTZe0xLm0VgQRu
rznj4Bb2b8tO+O1WlZafT5/flR6wy9nINmS6nuIdeWPTRcO9uh8+m2wbLZrqiqrn
fWQmNdMs7bAIqfLf+LpsUj45nk6CZW4wwUnDI9eP70ls62MjCq4ho5y6QOEwiR9E
HFYVpzuKMggKq2e88JbRDPqk4U9clewM99T4bhio7j8LBsRd0x7MbO496K65bOaf
KtXdxZxD8OcfR797o/ej+WROKZe0aq4ee7pwN1+UYKIBL17C1S74NVdE1ME1n0qa
rPssdhGK0fU3jodnUVeeTidBYLFfkiog388iml26neaijIbTqyf0k8Bv+WDgsK4S
NORhgXnWgF8Mkv08HLHjA/6FuTr4Dq+VyXlZVchrXNYLmLQ9jdSRowjWotkimOaR
5ITxkMVxy2B0pJjGFZ1Si/pxYb0wbLdIUeG46GcLUfDdQ/FLTN8AYzJieqvJLIAP
veHdipRlHJ+T/nowJQ73+AXaXsZ4wquhIQGahNBFXQnVQcO9R9+bEPUjNrJgGRCB
RgYXbICSY1zJkVMEpcIjsoodLZU0LvwM3ku5Ad549mLo4hrK2H+YtApNxPmD7BQN
PVDwLGn7fMBey2LahDNkTZVnHg/mUqu+hQyJasSgCuDF8llpCJlpNnMLS+9tAKnd
8kSNHZX8TNFfmYm1gkqBc0FzS/NiWju1s3X9P8XwUyZKY1AbJ74KAwWxK80+zBaI
HnNoM8B7CvUgCwMSuW9sfuvKhsJps/rLTIXX6XUJtvXdJpZEQAMRiusMqtsvoBSu
WRHW1uc13juPR8QfvSmSHN2caWMkbv23MkI26MO10d7hkhrRxvLnFROaz1MgQPi2
8sL09+s6GFM+152O2td56Ch356IieBtWxXQXBMnRdweYlpxrdWVBLdhAPoJbl3uG
FN/sfc8JSkIHlcpjmHN41lgCO6VVOr1l3IcI2A7Q4nFUqSkJjK1RDz/zQ3UPd1my
U3ESKxm3pqsWvZvjNER+H5ltyMml4XRnTqCXfvk5Nr7T45AI6Bcj/yexHiJuxA/q
qrFsI2AKGrKog37MsADn44NrjFuEro52/eLJ/ICFWECYHnyQqp8pwqs/IY255dIY
i+GOgwHX7DF6n0C/mEjDJXoM7xWYMtNjk+YOJQ0hsCMKf7mkwxykfd0Gm95Hbj5/
JnpDIK/KmbiwSex0fNNlJ4g+U9PXCzF1Zw9qIwnE8/oPBN29BtGUh1frfulXictQ
tei6PA/6DRcnPAv/BYjYijMFhf0tw5QUmuppJMODmwgLdLuqZxI7+27192oyeblk
sYb/7ZkznTazqgPvnYNhSmFBrSFaea6MYyPC6X1CO6X/bSD1bBu7+JJii6hHQv89
7VkK980wjbJHFSo1lK8wMAdnw648IYMT1PxaiVZ/wj4VNNfhGdL79pTk/3LRC0tE
ohSui3a+c41XI5ewL4KPKH6YsY9WCrDRdfRkGwMFBDldEYoZq5J+l9VoIW3IjZNI
G4qyx1xLmsfCZWkOxFCDIiRUv5YUM+21YS3xtrBZHn94ZeOpgvGXf20XfwVzfpig
kYQqKlCofPKauv/T9yKK3e4n1Hb2EEj3j0I6odPjpIg2yUwClj7wP32lV8XCnbSh
MUdficZO/EB008PcVMqaN7TYnJjMTHF0Df4jbJIied+XapmSMv85y7L9XhNbRONk
6PHsepbu/yPurQc2n7P5VVBH4fhuNddQyHDAMg7tjqSu3JUi+nbwdrXKDKDsSpER
/0uKcMG0/JGf+EZebyY3lKeFK0Vhnvcr3pKtr3BrFKxxJ2JeF6ufUvzb7DFAvdgC
RkzPBHnajuyJiFrU6fqQvWNObh1BKPecZ8h6HueZQM41OVzBvNsc/4XRikZTb3Xg
9VBbVNksVm0BnDASpfFd4BdXE23J86DbLUoUDc3TT+liTfkuRrpsdf3M99JPWCzX
C/pwwZqUqWVzbF+xpy20a3YIzypy/i1dXRuDzzSaOhsKHUkaHXLQ+yzSzFtMp05d
WdOKP0Vg+t5ttOE585gkBzm1oTd+vnglAZaLcQqP3qIhkITpDizaVCi+o1RyrouT
WVgbpyKLqhnaHCkby3kAk11thZ5mSiNYp9SUgc9BVm7fPasiLXeVg/d7M7YJGX6F
XCbz1hA7Qkk3ErNb6PYyd1GIAW4KMbkirnja39J5xOnyqgdWXGI8Xq6MiDl/2FGr
JCkkp7dxQJE/2Zt2TS6vs6wsH+CxYRNPqZXbq0WcVWvB1e/3M/5ZS3P0Q7VRVg/j
RMLObgdfwVVMAYTgCtRBo33wGzu+DuYwD4GOR7tujT527fYyUvTF8rN48+urF9io
fluAYpX0u/YDB7GwJQ2BRiuR+xnaNQIbNQpujsZ1IDuB2oUv06m/+kaeiU5iDlz7
NYNBKR1zG0knrNrYK3uPiKFPUMkDuSGsp6HKlDhULeLeQ0FAIr27zPGYekPcT68B
n+LiZA1e5fOEV7QyLdwqxm+JYVA5/qeXmTV9+n60FMXdg4medatThhuC3vPL7fy8
F35lkbVS0VaZLNMFmlEFlxjbwUJL0mPYtnrIWbBfP2q+NFkSjm8BcKbm1PNSPUVK
Qz67DhdatdhzZ0Uf5PLWLip97c8nQ/P5gwpRrel2ZoHWrwkhRdeDTUmFzSvDwH5F
CAOsmN7/5umaHlhDBjX+f/tpr7QDZfFOC5fm+CIXQY3xDgzjDKawT4eqPS84JzOK
aJ+p1A/Ac2G6Rsq9KyEYSWFfjDhyXRoPPGY6g7NgroV3YROzKZFCvbOWwUiw4vyd
ERSOYY0T/JrI0nIwZNrFd/RdqYHetJpVjqogXq52+D+JlRZWgoalBNUQUQEsFPku
J9eLQcTO/QJjahRdOtXyF/8IC6MJB320gJjWVxdBn5mN96R9kVZrq+YbQakpo2rl
rSNpmp+cqQizmIvjpJSVV2Fs1p/jLNXNyTxFNMSRCqret6sVn66yaIGOYiHwwwiM
bBO/6vCsst4J+glESMej80SiUfGbCRSw9HvZ+4HPq0URPAD+3iDI21iffTU2Osbx
zTWQvAgFymw/e6dO/KYFgS10W5mP3GX83ZtqLGOhfVRc5MKDNBMdQHK8a3oTsCzx
AijJ7VbzRQ/2cy5Wq2WvUq0f2dnBpOYlw+xEmwEe4IspiK3ISzSW0AO/6C8NKFka
UiQS6Xuh5iyvArjesTEnPkVyNWUwpyrLqRVfAD181jNXxSsTrE64NLIqAZHIVniY
cr52zpml5vLVADzU2HJSrdcXqXTt44v9sjS9gP37WTPvO2EbolKtj7EGy3BgXbvW
lOHYzvbmZ39e+7URBGwgYUwDf9823tqgMSbzt/t9dbHsLmUY4YAJ63FzxP9QUdYE
Komgag0aCkTdsVXyqW+cNoSQvrQoe/WqCWlveDFBTtC/A1ltemyimK/mG7aJhBLX
cO1ByEQjGrSCIhhXPPhT0LZSSPTNmm36Smdi89aD5AZLNwX1S0WzLKNBXytKokuk
XcynxqLbWfA59MwotsyaQzjmLM2SPNLnoKzUjgZONJ/oFZXXUMuYVjVcOZfPIJ1+
NL/MqrDAB5S3ULmbE+Ed/AUPAnGZR/9fVs4Ka73Zex6yzaFDRovnA67+dcpMc01x
KV4jGuSk5X/8Mdq7E8Xm4iw0L2BMfZlOuICjKYjtynNkA2YF4cEkxgjqw0TiqDG1
LvMzYPBCQv/DpbhQJj9tb2h4/lrexs7ylG4iTkMIY/cXqiWRQkfYxEDChWtIQM/S
9GZWp/R3lKeW4WuJzja1iqlbo1LDKkrvCNqaVY9YseRuYX/IpSKXT9hqYqWKTlMb
qF4PhxCut3cfKxrNOpfaZX2MdvPKyzMzgddhtmlAMZ1qPND7UJ1lBzLzqlJuaPg5
OevXYLrxxyezpCB+4aKUchUGW9x5QZzRi+kklxysDDAtzezb6LBjF2i0W1uKLBx8
Frc6s+xy96E5FbRezMvsUDZbGNWGYG0kotsRfUTRhBWAOiMGjlM/VZxh3+v2qnNV
abIcx/1h1Gu8SwiHYV87JqrpPHWPbYAXAEhix9fcvrB3CG6m2byLWJKzaXgabSVE
uC7PsHVGjcGj9hOgn4DmxWnrkfITM5BXpiaWgImCf7NboCNuwy+oq+XZT1P5ii85
FHyiOlWgxy9+wIf8MWXx3I6zY4L950D47ehmJmbcx5MDv0dqODdedqdTrpSdMsSi
ztiJHZgkM/m1M9+VXchLuMwNfUIsl94yq4OIIqR3VDDDjxYpMj9K45s+XlBTQw5r
Qv/BK9lPdX+Ty/e0nVgg7JiWdi3rnUt27T/GsWN4fiyjnCbJBpTpI87dTkHla2ZW
rx7SmK5tlbJcd0Ddlup9sbfdXMmdslzTvcNny7L1lSzOxigvyG9bXJvNfCxaUO7B
4Flw38gW/IJZPZqdEznWj0Y+w0yhtT/fa8abgDWQVTxDuTbcnR6PGtRsUOOZNv+r
4tUqv/xenLWQFS/T7br8a1UkvlADLKRPYbd9gIITrsI3xjvVshEwIfTI74LtvBkM
mCaqkplWnBmYllUCdpiU3HEXzjPIoO9AyYpigyzkOwS/tLXm5uKK6hN+7Q8da2Wq
s2YVsDKulYpeA/jHN8ievQjeVGk3xR4ViS6L+rooV30cAoCotfvSESF8tCH3F1c0
hkaqEq8t/7XvZdL7nQnOSmsDeZqIXickk+Jfn/ykfuvfQO0pV6v04ng5OvDO8QoO
FnN2Ojc/u/bs0G9r2E5yWOmN41i1d5suL4ujfqFCK/zWhOLKe4AeQLGZNOPDxspj
BH1nv1/+gKM1JNygqaCxkN1Nts0HRQe2TiYr3laN5YFpY2YUypeLvwV09y/xihy1
OtDF9676iOARNycne1KtyvhbT/joiPvFfRuQzlQZjCbqOjqmIxxyxCoF+MzR5SeB
Kzfm3RdX1DpEMkYlg1chL4CtotFyM9N0t12WHfhoI+nugLiLsmIPDsmhGZF0XbaO
225/I1+MZiIGVI7aOY+wgr6Ox4FdHRzJczC9CaBq+uWmPNhxZ3PvFkMa7ZTmGynw
Ah/CPh7Zunbv7APeXrzIlGB8sa/2ShSsMs5domLGEHVUXmC4Is7aDd3jAHt9BCaO
th3j3Ee3Ms+Ry3z+JwGKyS6eh38uPERXpBl0vbg+DHd/OxWMI7nMBtjN/YTfkJSH
XC0E4XEeu/c0LyrbqiFZhb3JVEUK9jYby78ppQBLMXJIvsHjNCJmoRw3Olg1ZUdQ
cyXTfoa5FBgqOlSAKHYzI+KTrNiG2AUIQkOeVJM2ud+7BocvkmQeXs4tTfrys5UO
n3NF/aijWQk/VRzOd8kCUV+mN7VF7ot7fkd66ytFFD8afNAp/Hg/P0aRelkZdAOF
0tHPO/0+U3DLic+NgbknfiDaW5xSdB4kul4SbDXTP/rReBh+eFNMuo2ZG6qKqIIy
ZCLG9GCE89XUVZpEIvqR2UZspCl4sF0HiC+wBjP/mKqft6KevuGhl/nNOpstfwxB
f4gWJRZ3YnC5nYImqd3cIMsKv5JkJBKESPk/RSyolacgjD0WluFX98QfAHG0Bvdw
N2Uhnc/p2Se5khyHGsAIZttUPMaLFgwSWMPyOj3jCtuKYHwQ3sO4TlP8K4gRtaUK
tIucbF98Etkw9GjTJ+g8Uc5xQlga+dV/DbPxmZEjMsl2RfB+jGYBYjqMz8D4CKgv
zi1nhi4WqfjMIMd9j04podhLor6Fy3nH6joiCs4JR5gR9L/vBzlzdeNEvHuuOk9/
0MDxfuH7RKnMaeCHonIiE18yufkGkA4mWotDn76KTaHxcIJ/hWVFZPdTqJTUw+4h
ey5Jt7+0xdhw69khh0sO5RaAlXIN9PMCfskc2GeL1ykKEm/r7i0aDDBJ3F0FvVfY
A6UAM+WWr/5meAARUntGipg91eEK99bzDUxcZIZbLugn2UAKX6hX9voDVET9Yovq
H92O8D8rWn0wxfcpZhQLvcwoxvKcKIkwVKQ8LmuiMfUmfMWciUqDclUzfcmSLM6d
x1nZTewvEbacMUWKTqHG+I7cmwoV0zhODK81217LgkGul0BTV+MZMj6RVqbAwvQg
XgL1K6iHhfUYygwXtUPNMV7k+XOc+6CuE7Q3mDBfk0bOB6LZhhIfaj0t9GcdWxxU
hBseXHBGYMQEHwCoo3Xc/Yioh/nySHyJpXeJzqhcdCdQUYYQUhC92Zs8aTRea9xT
/vu3C0IyN/jvDt4odRy1ZxurIWOGmrHJmJrZF+CKiBXMizE14qroQKiW1C+DcnUR
FRRUHGFejGqxAVrieprWN5coWxOST251Cg/YR9RisJse3H1Tew5QTWRqqcsMWZUw
67yvlFXcy7+2ji2gw5jnTYVBS62XiFIAUpvve6Kn9GszTxTrAb9vEb8v82bIRs9z
0mro4ZJsj17oHcgsw94vTfy1GUgwFNkrvI+0H9v4VKcYzaKCAM/F7eTUfd+WZJyN
e17GfS//D//PERDcOrBHBGosXl7ASyyl+E4Px8DMkzOZ4ScZmE9vuHQwuB91y3Sg
7dSwGQESlFAfLrG39Q8ZfPeNQAcTB4rgTDl7zgn0vf8Cm5d/8ENdVpxUL4zNgqUN
T05+N2HOeYB9yhzBvXpfvkYulWQt9KPtAEudixRPnl/lk0l+RHZ0pdxxRO/7WUaL
rcY6dxfnJlCotGo9sBKgzXdEWrCiRfq57PJvYVDlB9PtKlDGd2xMR5u+UHWuHzTe
bzOiZd0CXq7uPnBQHdMHJQ8zPqBypFKL1feAVs7YrCznSxaJs4LVIIB+TBqeebbY
fwCoIsfbtHjgByhIB0l6zNoHZFNRSfJaq5CZMMM+V9qJ8s3i1kRT07CiSaEUyFxC
gGexv4QTFJBrlXePdw/4X9emfgdpeodcgDGvVE3HnKc5xluRiVaNq2KYufftXJll
Fp3eaFTeMSrefaZfwxyV3NsAL4FF7oXdsnfZFpWRzCBCIKgYcZQdXOHGWuNzB269
8cnYq4mvlqH/s5RpCrLflUomcUHwrBKWT04IIW9qC72wOhx9uWmJeirGP4MGSkLO
ZrzG400gFoo67Ft/ojoOZFGKTIFWY9V/zRK7LubsCRTFH99ib55gQT4BUJCbeGIE
F7TSsNJp+O9RC3xlurSMC3tDBcxpJWi6+NTlgs3VhlOKsk/YdvklQz3+BOIv2CKN
CBislLmCj/SzS5s9tYmRWf1o9yK+NP/Mdru/t+c1r5mV9HBFEQxZzNuB/IE9MMpG
9Y437cBTJaCRMPJGA+Nx4HoL0+o4XJ9U+/3xY4YSIHyGe+lgTwqCuAeB0o0f93/9
g2p4Q/dj4sUT1C30MxE9YEDFu05Hb2kxn3GwOFRhgEmPGcUHZ5Su58FG+hKW1nw7
3D0ftLAO2xaqRlS7gwX+mMJu6j2Smhrq2OwTD5NYHcaSHldyUAXT1n8TJgx1WLad
LI+MRyferbg8JDuicsgxXOj4Cb9sTX3f+PyTYFVVFH9j8zXJ90+k3rdW/L4REJCY
TRwolYw1dVWbmR6Q+4LDLzX9uiH5MOEepm7kARl+EdXCtfm0rFo33GtmGXDixMl0
4PtHqrU/C6Yn8rrFxGsLLS5shmNi3LCDrNCxCxd6w5fHvd6jGiD+yUAbJz1Pwrop
I/2LhKLcuiEj8suGRbHayP4cWTwEbIoinYt/b0PV44yyEziCDd/Ip4WvHsV9986J
5W2tB+Q1Ff6eHadKPh2a/jRmBkf/Js6zJ+lNmowMKU2V+c+M68Gu7t+btd62Dd5Q
Uz1/pLurDCE46t7crrtz7A/SRHW/MiS6WMqerOt8Z9/CzzNcZJ4dVfLMotmwsgjI
iZ/zqutxDogs2CRQhKZ+oFBh5SSMZJiGnRnK6JULfSX+KBoDbXJPrwaug5R5lNdW
iTDBJwfwtPtkcSkoQhEg5pFJcYZLzh/a0V28NlgRTK09I3wpvZWjfPAKTytrMexL
ubrQFaZB42IgJLuWDPOzmMxgY/Qf4Gkq2mCpp+xI2Ag0P0laG7syhs8YbKiYAlPs
bDRMDZi6ZOSuEQoo0BT9tfFxvlLZIiVW9oRO9lLaiF7MxCm8+UpxzYEH7QM0T+xA
jyLqr0mAbzLzMSvx73OXEmu/uBNKPqAll9OyG+Ekk51jBm0TiuYlUrB+Z66deEsq
ezNBrucdnv/GdO890DlUSrcwZvcR3iax8NbzUjce9Fnn93M2/ger8seL5YWSvRf/
afLqH8wU8AeOej3Xeb3FldyHV/kRunDutdtZJv1xkiiHhBsRVKBBA4Z6atwLwlvP
yuQVeMYrM62PKt1M853+6ukUiKrj3JOoRtAHtwgbMGQ7qAQQx/Y1HKRUr3Z61jhY
x0eAAUnKg7GWS6rRBdfiR8PGWb7gmDgsV/g7lZv8Yw/v/KP2+sqXXDKqg+loEM4h
GSs4h0gzWo5gUmNkJe4EoWX0SzHA/p7zSJqJJIbUnqx7xheLQQpjSFOfGWD4kf6j
eICgdiWN1fo4ToKnGN73vUU90b0l4CMQqKge3SCIuErDPMegegNGT+YSjKoadutH
ua9YsJP81R11DCtjbwLMv5sw9B0Tcbm7hmzMMeRhXFd6UJgEaYEOSNFUW9jrFOnv
asjU4uF1Vvr+KDzLDsWnMc2VUWpPI2vhJlcScBBK5yIeTwwRnr8kTeqNllZcdYlI
hzT2LzmUIXXfmhjUOIqVun/w7EK6CHmv7Bnp2S+V4m6PKgmknK/J39I8y3cT14GX
9Vthuq54IPXpmAOTKuR8jrzHfPAadh3qOtwxfTT+EP+NzejwTD+W9iXowoVleFU3
RuKOw50Z4ZlCGhWUlkvLPeHdnQNC9xVAayTdAfb37jD9Soi47ntmO7AupbLotHjk
KprfcFPNhXDVmsGIogOsQ3Ja2EJE2SDmtQaD9mMyxXcJt6MmLnSwUnNmsSTvpmJx
CBM3sv/0nllKYv0+P0+cI4lrN12e/RgPSW81OfMeuH1/GvNyV/LVBJs8DKW+ixf0
w6y8xJoa9MDi8AI9/+FCl/G8eLOcpQsSDeRnNQifTLt79MZQjFSTMCVkQVkWWvKC
W4Muek91JnP+G3Jpa2SaGpcERVG2cxKubZdbO3QtAiGSSTEFe9DP3Y0qnYWguQDY
kCtSRLKzmmXQtzhR3YGD70SO9zPr7pse4OKh0ZIV99fCUh9uXNQV6RwcMIc2mQm+
kmn5ob2FHarKCFmpBysnQVcLcAb0Dv0qGNIATsAQkshYwSd7JQam0zkWjxSqVAkr
o4bF7wsbOxLdYV7lYiDg7DCO4o9eQbi/89NXpEUUj3unnKgbwmXVTAoDcLxJdRm7
1EvT8+nJyh6/Bu/iIq37pgBEkYZ1LDmXOOyACaaF3Xzx2vZpJpUappWqXQRDvIkq
G4EqQDNi0FxomiIJn+KCC47nEunE3qkYfxJTm8gF0jXtvVFs6dCiQTxIQLtVk5LC
d2OIkhxrOBmyZiAXHGmQy6L2+evOLRBrbQRPQKgNgNj4Sgh/T8FPyuAOnhEUADYx
36FnabnJ4CxG0sAUAk2x+5iEQMYE76j/EiKYBmnEI3ncHr2T1AFBp5/1mXXNnnRa
SGwnwzxkwGgmMjQBS7Hu++a0DGxj9EeYY5r55mfCsds1vU6qDnaEAKgNpXB+/Sf2
xaQIRME/lBPCAdjcomdkxvVQGTmTkrbZdm5LE2HpFGs/r7cUeEr97YnEgIID748z
9IiuD3nk8EEmCck6pFgCAl0fBjn+5JTKXu/R/topHEGsalv0NWsRHWJkHiOrHCXN
L99Wp7Pbpg9FqFgJKFKL6Cp5LrIn7kkbwFgnwGf3bppzwpyXlf3HQO7FAK6C9u3o
z0rtew9gcteCpyWyX/0mZ+KlOHYU2mnPr6nQMNU9NQkt2W4LZeHmAW+9lEifaaRj
8k2FI2EdOTGrK7xQtWeUvx/ws2Kl9xkITY/bn/SJaYCEdeIUkksJ1pSB2c6iExL/
D6AwyOetWWRGMWHswiB3sVNs4nNwL3PxW3XgnUj2RCKXkDM6AQHbTbczvqCxnxxU
izjwaFgNg+N9tsPokU1t2vQCqJ+7p2Zk9D+XHmnbkqv16/zxVDFDVpy6qD3w9j6r
zxo3PPifRTLL062L5D8M6F1iL5TZKqlPIr27sDD1IsxN/U0xi/mdic9b2qDi0auQ
KLX85W/io62XqM0v/2Q3XDO3+UyXdoqs0Hhu6Xk95g9hGMPH/J9TK9BSSHXZlZXZ
NMLR4d7rdFpPEtAtsQSD0GGE1EBg4PKI5A7C8CVWyW79SyOommFWfK0oQi4Aiprr
+fMCzlTVOQp1XJX5Rl7IKZ4KIupt89QZpCscI1TlLcL/9jUf+dBgz5+ZLrMWMWb1
wgfcSDJ8sTksTkd1lr1WA4qlDv/18HogFLYJxFZfja0sJVlR8yFuZxlneBW4j+it
LtBAqWj0hxswd8yccpNbU2T1l1yRahLpIs90Zdgvao91QEdTEWo1qBDUKTvE7Etx
Jj8MzxO6ZZTd26McKABuhXlrK1GPPEUOQHAEwTn4MUuPjGv3DsvVaaoDDJo6t1jQ
BEi8s+rrpLgkE2wNoSZIYUUJw2t2Vn8cb/1ELAGPiXIZR0RWAR61hTRODlDEkILP
RTLvQfoYp39ZrTENnTGMKZ8ZLvgKH6h+2ac9Gr0+RSO231Y4nO8/fhPRF7n3ig6R
ZUZyKwmcDSSQd4LgqAh/GPPQvUFTya4iIWaQR5RLnlXF4nkvJrfadc+Hb89eouit
jNxedpXXylK0nidYIdR4E4SA3gA683XlvwjVn2cL4t1nemLPbM3iUCSM66a5VAdc
x7HQ0quivGUgFSVzKhjmljS+KWFXyzNWRwtN0atZ+YLUO42jrYzlz/yJLLKyZ8fZ
Psy1nto+GNSU+tMxTe0jBgUiyCgnc4DJ8iffE/+kDGkpUR651cR9uxnod11oKDIT
xoVMgP5EOvmaVfdElZX8PXJGgRnmKA+eF+nWZVnmY9PUl7vgYU5U7/B/uwHIPNHk
cHJstRuKqVU2EEURSNnro2Qybu/SaeOxUrM1uLMUuXuGnKxSsZ2fPdFFds1jiQj1
x1mnol41bs6Zes2hDYSgy3jMcfqgvTNJJ+2TzQVHLxoMW/vjUbZuE8KGMYFvAOPH
Mm/DDrEGfWj5ysDFHmgs8wvViEMeh9fLEHRhRFs1rO/9NH+p2VW1NSUC9BecTJhp
2wBZrlHSvatpywmRhIg2cWHc250IEWja8VahFVdtSzxF4PRdQMtBk+VZWPEisRP1
9hTBz/U9rO+p9wwsJe6DlMzN6sttwgbtbgP/q9t5khA9o67XLvij+gpkO26MH8n9
EH9vOsSF8iH9K7NyXPNhThVtFmV1oyHwOc5c8qcub24FSYTyZJVkENxqVHCJP1+q
KjngS5/0yTiVh6k5XcXlGGhQKoRv6FGHpTJxnP7ftcoOfxbqsvhzNpiRr8H94R1u
4840+kI9gU9DCmTMjw44l5SSbgI/wmkLp7VRzr3wqs05m8aARFURJKFOGR1nZEsq
WxOmoOtvNkW92Z6Z1yDy/V8a8RTiHLOKMu5WFd5u0PeMRIJkL2Q7UhCP3drMgVIb
fC8mqBqNdFMRp4Y0z+BFx9lvedwl119zbEQ3nBm/Uf4LGLEndHDRw7stCZcEhfDd
dehQGNA+Hh2MUBEAkQ9pglNjZoe1gBIZoW/JgTe3lXmS0zsT1UKkARf0o/WAggDU
GoG39xrA26ErwkrBxfpOX6lR/RAf+49w2AXEoGo3Wc0CCdRWj6wa7iMel20AzfNX
ABP2cx7yA36jln448ky8QX8jowhmng1xhUg3wInXPU6FPNHk3SV5XQgIWKJGYsNL
a7JoRimhdCXm97vs9By1CL0vFtL4EaId98IBCw7Jsuhx7wTasJCODxmSuAKbiyJH
6+yE74BsJwT69CjFoor1qIDM2BHdBT4iYxV69qot9pRu2woBJyUCcTUPYrhKuKb2
rfftPjxhKMpeKy4IRtdujOewkpyzBOm4oKoC1CNSLT+O16cVhXZOB8aR4Rb5wC6X
PQfq0pgTeDkeMbxp8lJArTA4GZs7z1leshtuAdd21WAODgEqNWoEyEu6jLl9s9NI
+ftYrvCG8gPw79Jzem16SztlRx/Y5tyKrwxIMopmxBWmM4GCnDlQKktPVU8vqwXR
szXX4tBwouWz2R8ja5o17EZdZ+JKSavxjzSJgSmK3Qf/CVLJvS4xAT267O7ghr/A
RSZAVGt3JhrHbTkjbygNe6MQ+/KLmPOwmFGLCuSfKhNQC6hFrvkoDU2P9hopW5AV
+dqfvPfuAPOESiTyIG1KhRA1kkI8f+HR0X1FVVAvVW4yeMiLJBryrYh9I3nYwXa6
BqpyYgjZzIhN4mqD56LNHb3WsicXJLA4NjBjLuUrD01THUNHhE81e9DmVtnM8MCb
Pt2Bs58L1NbbSQG1mv+u52vYjfYgC76HU4AyEPfiyII2Eaj00M1JrSdNqnvqB/7A
i50/sSEGl0oKAQazITgrnd6C5nFPbJX/BBN0rYWEVPNIGzh93httNt20ew6zsTuj
H7dSozfA//9LePoM4VrtOaj2581PG1SYYlBabJ1BCIh93EQjtDZZqy0YAI/UNvI8
nQUaxiTIWa5RD/zM7A4n9lQbnZa2EqcdDyxZGj2afNkthCzZXseiF+smX2s7l2q6
JLs225Vb+DOxtYjw7BnybGDdQCFI/vjbRL30fVP81eO/X5qxWYyitW2nkvxcP8J2
CFltYQhZMKAY5AtYqeT41YL8RL7+KDC2etyR6L0d3zOV2p+Zv1FDYj0c/ysnXPrz
vniFVT8lsOCxoPl3MCXNoaJHkK6pqAwi5y29wjhF3ZMv0LYoVyq9QqxMPEz02e92
FuJNO4EEDEhGY/NpG3v20B/J4BzeiQj+Jr9p317qAttNjhi/sUUSYaI5705348gC
cYVARk/ztlPG8+zRXUOo1IWMEb0XCD6j9WL99BlCAkmng9gBGDbEClFwgUAuPpac
r4irrQKvT8fjH+VlauBPPBLmP0TiHrSfX2PNu7mPZ0rksG6uvmaC7jBBl++8fACA
QU8ziM+Wofz//PZw86XAjKpaBJRhXzajNnEPS81G+SaB67LVz6XOTI/qvhQLG2ze
RdPNMf94UTY+H2LIcDnsIPWKHSV/cOjXLeC8jnjOm/mtqfNJIExMLn12qSiLtZpu
PaH3yfGfDoBeL51Wn4ckWFKBZETDDKi2KTRlkfIfiNRZdYR4dohXhN97bBkdfRwG
WGKn15RpTObWQfiBtUik4Mee4z4E2cAlZIMMkgPfFG6WYM7FpqftqGvt/InNlS7I
DLzi9CnxiGFvXrrwrIUP0CP9t5wZX+EnWwpChB9hm9W/3V089K02Rf8GN0WUCjNQ
QWl2bqOyB2x27RzuJgHZ8HX74dRo9LSCqmKGNPfFe/pCv1Z9z6qVcPldh/aW8fSp
NweVqu0hZQJAvvNg0Ljfwhu1VUScnzR2KjOIQC5me6EeGdykXlS1u3lST6CdnCZc
wkyEseTBtfnERnQpEFn5A0/TybHT5LumoIzMiBYZI+Iy5fyfALBgNL1CP9s+RlkY
XDwXtbbpc97fSWV83WL0yA3E7X2IuLIWuvg4W8DNljW3zPEA5aE0Hyjdrsqec9/0
EBWh11r5rtvMdWNAl+f4rbm0ap7Hej/uSJjYyl5vkUz1f4G8rBh4S6zXrg8ZRlnE
USrmcANieJ9ssZss3b/reoJWAsX9ztm7jubS/VC0OBCdKNMZeBQZ/5gRACFfW0ps
rsMBU+q8UaEAaPh3R44EB4luEvbPDcC5vE54QPVe1oCE8fPn9NHvYUcWve1OxBt/
JknOc+YGs/w+wUVqRhDf4geksAkkNvNIHMLzvsLmNb3AdkqzPICaaFD+31OSdsTq
cOQ1kceP1RfXPGjxB69xztSCiPESatKZdbM1NECUo/n9P02AXGJQdKMZdtXD0Ekm
UJ4RWKR/8ppV7LMpfuaXdDdCKAFQ4ld8N43wmVaH+tb331SPWQjXktsayEBBXQQU
PLkHySWZGxgdbffNWCtAyxc6i1pzFUk+g0jBQYplPr+okvuZvsOZKnIvBqG0yvK5
RURyMykOll/zhVCRupZSyBb08rOsAKgoCOg7BFOAy7JhrcyaeLkzi0OhOOKj6XpM
Drh7p68ZGchbCjUIyYjAe7obJO9zEn6tcKamI1GxAONI77f57RfKpchYm5iyRux0
JjrkRkhi7L+XajWt8pdBsI4fopBp+v7myDHg5Z7phoErTxBUnRZcP1ynG1JoUEGU
9oZpimbV5wdnatxQJqvPTJiMN/ASswQQn9dxaX8NqFInLHCXGaR3BmBZHoklW5g+
TuHBjRwfp/84iZr+E552nyCHYlY2Dz/2v9oKM0tNtfz58jmKs41gKJroYTjs+XG2
/qY1Dz+n6aH0kpFP9cVyA50tQXeKFcS1FfzjMrkixYM2Cnj5qbuNrNgsxBzsrLQr
p19om1EoAwI6Ai1EoG36NqLR5g9x4tv8Wg0HBbltL5KN5YVZbTM/XdT6jeUbb30U
q1yqgil2/rnDdwUrnVTq1edjrMzTkVo94rw6+0X0TuIoT7969PKBqA0OEMQPNKwU
Rcz+ejwvFaNPaPcR5AH1wtiJ+FGXMZ8Svp9l9U03FsnRMq+IW55ybYzyd+qydQwa
PM8+JarKLCln4AASZsV/uKW4OhCv9p9BGat+h4/cH0Rts+t60LDrwWmIIlkAUC1V
Anl6FR08rjuRlVZs2XRohPqF+HnpHWxnsDuAF1YUmTtCaAzZ/W54cOzd5bAY9rBY
3wEpIu9xa6udrNlm0CWvJIYl0z3qlW6RjD9UdrSLcmqI4njEimaSs8Z8jH4QhwME
xENSSr+D+ppiZB8EPbkscIoIuBGGhtqSGRL6H7f793sZIA6f2GtuPyZICb3hDRTn
RfnmTW6qCc/ILgJ7t/fbgdudLIU4Q3fMBGoTGayIioGYuCi7heYFp8FcfJnJL+6D
FwuIlwzxXQqQGOqiE0+OsfRSjz97Q9iykId7NI+hay3ZywzWPM0bWIrcw+08XaXi
3sN117scoWEZiCnLMiML1wcXBd1m+GyDh2oT08nN7EXT4KMlY5PU+T4tYMX5ycBq
xsYx0lprrn8d/pGRf73Iw50j7vkXUSjYPOaYfcfP6pwYE0EXHt/veBcInno29N49
DbC5vaHAhkWzKfxzjktH6qxCqkhLFxSxeCiH+/ay73wEXOjLHIA00vRu5UHol5wN
FJ2sSxMWhwBaLaCvDBBM5GtmJscUx6w1hVl3vIaUc1Oc1jUidgHWXtZh8uzPyZwN
RVQsBKdBQoK1FJ0l3iVEIv6yOLFqfvsRQu0CKRz8Mw2djYwgVgxWgPq2LiV7qUN3
0zKZZmNvT2yuaJnhJpM12kjzMyv6Ty/Yp+TAz3BKpufGdxmmd9UfM9bHTgrdWvGe
29J471FL1GAOlIz/e+rJkUReeRhXMfgCXywHLZWKP7OmpIZ/Ti0PbqRxz2I7+0Qd
OEqCuTlJZY6+ALXfx0n5XSU8BX96Vu6uhp2MZjXG/JXM5TtnarpqwUZThymI88C3
nP03PIzUb42EbKkD/idE0ZQ+6SPK3fs3moVZHJtRYF7z+Z09HMPzsfzNlW7G9Tow
wL/IaGbSx2mbAC0f91kLAvTqolhorFT0+ZLgXcji1L20H4yoOSJar+bczKJBkdEM
jdzbJT7HyOcZnlyty5l/4Mln65G78TWbsEpgVQp6T1xnfn6zGYVNEKRq3SNwMoAq
xco+yQfBDTUERB9kYhLLizTpx6I7sj6KXmeKBiF3gmlFHmXqmolrnfJU1PrATEdV
NMP1gtjlZDi2pRaY6rzrVu0j/MtqMD5MNAy5HpFJAKilzfI8gSr7vgUxo9P3dN3Y
i8NqTPtrkrKmSsVAQB9VLo7GxCvIkbEzMlHOR3290fKM56qWJN+k+H779KeJhpAR
n+qZrSmIvPnKkUb3pCRHiihQ69+cTiWi7uXBCi4HLZoKGh6er9Rw1NduUe0slrVB
O+/ilJuBzuLsu6FAqopClmfOTK6NEj3kWSjR3WfzvPP6SAnW/TUMUCyrUOKBnW8P
kjOD1J40FcH101JTvEmqLlEyU2l8t4vjaexYdGLMvgeoxXJr7vAmyhU1FgQBd8TL
qAnyTYHSyhXvDDMjZm7Nlxiia6TMI57AsJnBeGiYnS1FEPOTGv6ojoeYjtDTlHSj
cKLxqO/OGcyOVSlmt3RNXztvt88fhPJzN4eNOtrfA9zmOcBgcYflLIzXkQmzSuMR
5R0JRIu0H/nRZfXbv9AqoO1kAVWbMgo3xlUR2KoHLncTiFfBVZrkN8YQlr/S9Qj+
5wnH+GqW4hHS9O4yzclpW1vSM39+wjiffjEV5eaIdIosziSUZhrD1qcY1NuFJyhm
3ZoDIXjzLf5hMLVv4nR+TsI99kMHSiHdOgRyhgsqqNmD5KhRDUOCN64ufZvv2A6S
dTFUGbW9C5fzBd+YiV8qbVZgJqAi4CwKToNYotCJEDc3nl9n+E0kbHQTmPtQEz56
qTi9lwRMLpanWKvaerTxHEV46TUWyszrrBOiKThn8xf/t4/RMs4IetBGBVOexjAv
G2Uiz6KK+Ph73n/2eJRnrzeDEmP4YBOI4WRfgx5ZQe1bs0i3v3aOJ6Yw/EY42kwx
saIV/wXLSuS/GdV1Vwdw/j7OPQMLI3fVsmj0oM0J7iJgY8ZiIplT4DaLtHTZLi5Y
BU3gR/tA6JEozg4KVEMz3t0/ISQYjGhIptX5FSGnPD2c/rBNSf+V6nvG+9Y9THR9
DCuJAvxMK22yW0uCIv24LJOGqF8yWiyU7wrd0XSQdVNpVu52cN+Hg9wpvdppCmcB
L/4LBZJlv1B26dEx9iVk5tP1Ihj+tCn/N1T2w6r9VVRDI3IJ85GPmk5wop8sgB3g
vm10Hg5DIhTz0xj6MqgOOs5xRDQzyRky7j0+8jStOsoRQabRBv7a2EbiPRkTYz23
2/A3kOfjCiOB7+bihkSBGiJbt+4+PCNmepPxa/TaGP+eLmE6l70Wekwvo5TxQsAL
eMZ9kLyFaJvA9TICx/iNLQxui3YOMeZz1DwOzjoZSvq7iRR0I/PsNaGJkQfI6/6o
1ULGZs8FoarrI7RpPAwxk+frXIECO9DePGWb4cGKGmdiK8sT03egdhXKYsECKPQ4
LEsXh0/QnW9yggBl+hrGFWR7DqE/eoQMHPyivTznmDpwD1epMzYC0Hasqvj4uNkT
aTxWDCYZMEmGj9deoAE1qbyquRf4/Fe8TXXzFdS1wSYXS3PsdYbrMR9cVM4+qg6Q
G+qBbbatGIk/ulFqs7p4ASOL28qgkq70zVQwoBv9Q6Sm8diTssF6+KOnHEw0fmDb
vX0oBzhEDyHxDlPodJTQ/azIvYB2M1B74Iui+w7AeGkMmipT5L8NHU4qio43tFN1
PXbjFYmIaPx6+mWYAY7CCw0i4hDE/z7MG9Yvji4gIF2nKOSv9aLdhnum8GJ5Deva
txgik+hMNLOtRZNdpdmI0+fKQaKpIoMiDtoOdT7QRZT2ADJK2GXL0Y61n5rWvqsu
mSGQ9tuNd5NA8BOy0cCO+JGVw9DQ3E6VzwStwZuhbIdLs7VPqk+FZr52zlI6EQXF
1xSLsu8sX5lsXKizhpvs4ozMxzs4z//OXGJaHqFCpz/havMfG563E3UBG16ZopbU
AhGBio1wUs76PpOeCoglK0AoXPc/tpcE9AwXhxM8eI11KGKTFYDfTeZUEeDLvvIM
QbKVbfpNDcpWVACdPDpar0g4CtG9y1ey0/dvR/2oKBUGoWr+FHE93zaT3DgYaPWS
sflGBjmn35tRrfSqeReIwU3Yvjh9z57akRpxVyY+tB6QcORSDYjqEbpeFa3Xov8Y
JaLUxrlqAYxpTDBYRnolWkodVTF3uVds8DhMrRRiCNSnGcyKen6w0VMKqlAY4Lvw
Ky4AeMJV93VhFEazIVn2ZmqHTZugsLJvOCBt7/sqnykapE3LfZaMg/y6IuaUVpCw
81orkdGjU9OzY2h9q4IjcTlFwwBRhtJLTbYYhhslz0pxfjpcI1Rx5wr9SMqxlOIk
wvTSC60uURA2dX4g9DON3GpmGK5dY29oMJfsngMGk+Jf6ITgvXQIgTIOcnNUo3vX
G47Et+wIOA/wKbs1fDVT7JBfO4QMCSl9MpT1N62gUp17rMN2ytzi42tSvXE6QgUD
BlVzwLKeo0Aq3XWe87G/vNhzg459HrJhGOADuN+kBDwRfKGxmFWOy+EnKIvAF/Wc
sY6ksiFV+FOK09+t81LJUg/OSGpPuhF8xabA4eduZXkUNCCm6VH2lTybbzeUdiD/
vEetUqKDyLlsmwA27kI2utz7V0CTS4dB2SkZ+igmgq5sMAxNHGfJqVtEAliPI5Jh
htJmt8ukUOvzrPcF9ltXjBtyH2EhDgt4Y8tMUS7BKSficnLiYHDqmh8rjVG2NqHL
k6RG0U1Igones7KZVVYvHRCn6FUq7winYwPglL6AXl95HOKeWjW1sBYqqgg75rZn
BHNvDWzw+zq5U1/LfTpNNJN69TiZpFSS9n4CQ5DnzcLMbrSCTlz605q7PbwHeax2
2bztYaLDRmhAvHIMlv989kBbmORI5Z7N7F/2Jvmhh4bPFcHzqph8Yeabjxqe8k9G
8kRXXql9+OeNLuPxIuyZgEXG34ksJzBWOXixOV3dIVpQlPk+n84otMofr4viQaso
tzb64L+4XO3qf32TGZPmo39pRnPQ61082AmBBqKoE8t4Xrs1d8tPEI4vivCt+80P
hKKG4x2EjWgsqfxsBmYcyGW7dqwmBWS/6ew1Z0HH8nuwBo1HafDkGcrhgsQXAAcq
qnaqrxOqJqW0yhXa3PM/uTQCdODev1vmXSfdmq4pI5eTPvsPnf4slc9+xlLsoM7h
DUaW43X0l5UAnlZrC6BsiIc5BCzhefK0O0OIbMmi27PLV1g4t/gARJH1ez1fz1XW
y/5QRtvYtJm3VadboRvhKBwLRib0a1mBMV2Zx2aGvAAroYh2D8iEDh0OFkF/ZZot
0vZnukOjjP0+DUtV978lS+MSotSMJDLb4iW5fN/jPTjWGNtfuuf2AUjHPPFdoAGz
zLHm/AW5XWKFDw38MjBz1bI0Kq+kxxYrpT9l4KxHDsvaOZjFsp5Y46YqWZEWgBVd
Yi3RTkRPAXbdRwTVJKyfoBa+NoyMPwTjq/iS9LzKZ0Na4kXjIIhc4AqWUpfvQnzx
olLijh0nZFN7z6stWZny53Yrqal8ZCVF9By/TO9tzlRsjLH3Vbfwwk2/kgilxqt4
vLbg5w3Tc0Kd57zralMHFSMeujEwPc1GBlYzwqjGSr+fNOPSNi/8z4yH6tNf4TDG
qrb9N9yQmJy/sMSNvXq1+b4DDswzZJs5CZjUDzrIvGWyz3AaN1hKSFOl023B9dY5
nTMMdEhszsgHDbfaM4H/5qBrstSDbazqpe1RddUZov0X0ps2l0w5Baf/TNqRetnB
TC7X89iL8ElEqtJGRMn/J6d3Q0R/IkDq+0dKTmgLwgVu3jP3wHt3RkMKoWZANdtC
m9MJGDWB/Mn1JNh4QLaIR2lXMgXrCf1nRdPcHimSWHbojY67X45zKM9LRngbp/v1
UTykbo5Rw0u5L1iUO2XksTmm6jZmGJr9VQEQZKhXuvJTGa0tH0PzmcupgXOgxbFE
Clh4fr/yTTGZo/w8pJ0VI1j4Yho6e2hkYu3X4IOFU7sRfLt2c1y5lR3IrSvVhZNN
24Rl3fO883YwHVTGXQi025NMS3RLzAIbzFxkkf11MQwk6pwZ+/bLTKL5D84PvpZy
wa7tkEz2HmXzfJEAQN7oz4CL+RkXKBY4nmHeNnFgGAP37oOLYFeGfzJvd1oBsvIF
N7Ij3jiBdYKniQidt4KAprMvjg9Xs5k27Cc7piD/XZtnn+20KD4dC3Z7q1nKpAZz
WyKiWWgTP1A483uiEKx4LNWgY84GrXU206q8T61HdJGMNCWFciQi8KSQQ+tkENL2
psA4oNUC4VLyNTaNMT+THfVVKMYtBxBPcRGvv/Ut28i8HyYjp9FFQXuevCZj0+Lp
amdyZRQMNkayZn9L1zILo6Udqj054NPFtpDMAD+RfPgFJlVYpFP1YkWKnu3O/oMj
r+uLHDJoiudxIvEFx+sxlb3pe9BSeEtC7KqQ2T3AkKRVITxAl2zLylaFaYiWiRlK
k+NI7S79gpxzrSMH0eYhaK23ESQuRiegnBlYqg5ADAF59Lwflqza45s2wHV0kD4D
6Owu02LmKdtKMcDVoKwQfWAZIkgwYqk5TbbdAcMjzzOC2CakADueqEgnepBlpVgx
pSK9aG/29UuA4HGSJosW8390B9KaZr3nRl+NQaiF1ppnLIMsKc1Rlv0CLpmvP8kJ
7MZ4RCZpfFsInDfiqt+D5ZUgET4YwRNjjG+QaRohhDpopbekxPvnVXDt/zeOYkHS
3Ac0RSEbqDOjWZvcbthLxkmLEaBhmKZeSnP+P9i7PwMpdaBcfJc7ALtlHuynQVU1
/cKl86AxzJ3QMiu1Zy7k8xCEMa6/llJyNarFtfMA8vHHW5shILSdzUEtg2/oXv17
UfW0Lq2GSMsZ8gKdD0RJh/qY1UpL5PDJpzy9ILm3v7/ZKncVqs5n7bK3pUm9XtSP
74mXDBHO9fSy+isYukAka53TWkD3rcjC0v+ciXII6WlJjcVAxjCeyBOm6N3bsyX8
g/EZd6xRz+fAGliuuv1fnXrdavzejHd/eRqlrZm/ZrTxL8T/9trvVOuam1JU6/lT
2IDQvgaDQmalFqvy1y4fTaA3ncTdH9IVEdx5WIzU+sZ7ED2N4uWFfELX6eu8n7UG
Qf90XaJ1cct781JFrao6LmHa6gyovAfLoS0AutusR+qCF+MRu40JcJBGwPrrJPBc
3+/9sI+b78GoE8ldEB/oZWhe4kIKnlJPt1vnfUTU1uU3EQ6j4X5P3MdHAZsnqwHg
Fzmjh0GK5VOT39yko8jI1wUf6Xo39xby5HmcvHm56Wa1eQ7kfa6/yJd4o4fjPFWW
bc5LJ5LAx2+mQNB03j4R1n/IZY/fwH/mILOFwakECQireef4Kad3VSjOqOXya4sb
PVYqReIYwqHMzvGDgVNn+WK3wEjqJJFKp0TLTyd/ie07MVQPuHVv5BDQnQ3swOiD
RHygH2yzCeyjCqGNCaZH9BVJSmb0cfgbGZEaXMm+Ta47/2YfPwp8EahgeNpqlz+v
jGAaMmQI1AXfdkNezE4tI3ALmntNLFzO5ntIhipWRmCPUzrhhJvt2W6X1H+5momv
HsRDcnK8derjjheQ3HXNWL4wiASwF8egptM64QyRjbr+6Wnh0dBZk4txs9M7DLuO
BoOX6zXpSEWFvEmTPUTaiPu7x3HwbTb7uluVtn/dcEYK/gytNVE9B00dJZb/mh6Z
l9cWuIq/CxoFndXrE3zLmacNcyxibpYVdlV7qxAlJUthuurE6o4kN8KFFANjMsze
umsi3S2tmcK69EyhwqQ1KHuJWMh1O+CnmvsElR/XoMqktBk4bWOiXlejLr170LIE
nYk8QZobGbw1XgJKqFDlFUFYqOLfLmnYMZ+jxYqxsZhIa/at9FVqUkzlXplptSLO
WNss3li0j0k5XXQ27KzJxnbuuMry57WNFmjAe0VjTRay0JxeA4DVKSkoNsnXgZdd
cLrcjOfMOTMTgixqH6lxPY+Sg767nNoj+AvNe2x1zsuTPIrdKGG5UlMGpOfguGyb
P8jlrd4ZxN0PKcxvzCVCk2uZX6RFKiIghslmNubnYL2DVOTXGsFUDZqxgZuu/2hd
hSdEczU0mYEjx0lkjCgmA1HCgLt9Szu+9ra3QqTFAby2OoHCfKFBCYP/nAHn3hFK
NPsT6yoqWTkQ3DwjbzMhF4gWPDV70BAMoNGFY7wX6r/LwHYevwCi1YDSnKcA7WHk
OlBM0OGOU6a0N0HoKMU9YBwpxoMIj2oM7FiRfl3Xr1M3mOp9eVHGMIsJOYBtn2kN
/wiNgHa+wU5JTdUocnkojNt5BnnkA+6XVe85vDtcSZQeAGn/nUBVG5whyDqCY8AF
dUBB4Uld46qFxGZlSB5VijJJUrJ2ttaamm1crN6vQRxd6PJbjJ7fY4nRu6xnz3aY
OlzflThRM9AMTGXyDX7/mdtBi9jC6unVktnGgtX9sVnAMdezX3PqkuqTm3KxPWSn
KiCHKijvAyVz4z8imLcQ7zHsdPeYlMyQ4ayYQMgKcHa3kpLcwovp1mNaEOF4gmtz
0Nosn1wtmbmLIPiM7Fe39lVV3ezkubt/829kHZX7XU21Dexh96N/BXzgqNF7xSjH
gF6lhfCysjsZSlhzOm3gueFbw+aFYwHSHi8Qh7RzswHD1mIjIILQIfnHRm2KDXwo
4YE6212SsXF0bzX7Er4FANUZBRLZ4G6QC6csV9DkV5xYWtIsPWlzNeCQymJPJvSO
PwyYNM9aAOZAtsrnOuqLJ3B6nMdstja9W2oKGa7TdGeP1rruIvYvR071ykQq9Wph
iBEG5Vg0nbKlp+297Iih/OVv3E7WW7sfvVO8Y87j5BZqkFfbikT8G9RdBEzwNVcX
V4R41qw/XevgDEdhFlbTtNH1knY6mNEtnmuOLe9eu0KbpcmhCUqFFII5f1k2SuOp
NzVyv/B51Mac0HuvvEtv+nFSHy3QGzbdlxkha+sBmnyj1dHRp+sFN3ocJ2r5O0Cp
pIDBgxlc2wR5AfV8BdJIoIJF/J+b5/OK0dRap+IRRXnYs9SmYOEEHnf+TT2AM6pD
1UKONiWTRe0++ngRbvzPFKPSsdubKvkTvt9AfsPTC4qq6hG0we7N432zxLffpqK/
tEe6bc/YPoisReugVIU7FnMzx47U957pb6Frm2zrjpoPCL4h5lW0aSdOE1dogumz
Wu/+YcqhsZHauc9h0E8FYCE1yTKdVBZuWCcjLty5/HECV1VZn5T09m8JOsi2M1nR
NFNklsFpzGpDixKXHjKV5cSx/xqHxSbB4K7KRU5z8QKDdYdyV2ac4LQgxWvZPSA6
OzmBHxjVb7wR4WMCKwmOhqMbxR46U4aHpzxMdv6ys8pSFTQvM3sxmteJQwLYvoRG
uwBbzG6amfh30nbGxlFppAdmBbN6rOYLFrnM4+G0Ei0W/4SvOWuXfvfgRG043KOr
W075DORmhOWzhOhaLKYGRUBsAAbP6OfjiGN6zYc/CvHRJ44l0EFqYBmejgWYmR8d
v2+tQYbGBn0albfX+EAYHB0V7vddUWfxZPoarHC9hTzAdG3+dUmp/VmTJdIxrsCI
JnEzT0lHOP8E39kWdaYPJurNy7NCVwoQFqiVPxo2EL5uOaTWnttt4d2U/FbS00ca
Od4JdxIbc+Tb9SBZwb6gIg+e1Zp6ktQ1yr25hTbRID7Cg4T782+DnghNXlN/VGbI
nJhfs0Y0Xyn/uVRShacOWpkgDvX7oYAImGKJX7rwzijf8Q67BaalVwsS5cXsAl1U
m0TvFFSE9mMuMyRx8vx50HA+o/ZEoqUKuinqQQnSwYDJu2wVELHaJfOQxP3UYGfv
B1qq8gvHfq5I35Nk4gNLREcD7UVyUTNZvkqKPh6Qf/HnFHACNW8m9/NSX1Xld08A
bjboiP491FpTGGU+gKNTLexjCTTD5QZvWCBcVNKqsZL0GbyI7dMJ30atbBgPr7mj
QKWyMCGsr9v6HQhdgsZUzMufAyD59m2WYIAZDBo6Y9/GRUBMgKG7XMTY3QyEHMjW
yeMPsBU/dQlnfOuTfoVy9LwafhKYqMPH78fQw1dA3jKJXp0pM61/HMj6SSNxXqXw
77TymA27JRaKBz7bzWzeuBtck0Pn2TXEVjuP8TMlau5mGxNoF7BLKnl1SDiS5e4+
Vki0wBfRUa6uejCqChPRnMlYOPPskl8m8ZPvTIPqKYVXi+fqXg1jB39Rv0wogLoB
s4jl5M2x1qcLy5bOD4WoUjD6D44Qjnhpj+w2CJhX/2v6V4BhaIiqeNlBKgAoFjO5
8gQ5UoDPgNNiRDVoWlulV6Kazp6B8D39vkYWROc76EkGIRRMojgYt9WO264DGgwn
wkMHW9gnZIzAbKi+jcTSoK9wROpojqmdt84XQ2O6DuVfAHXsVxmZ6sKgXS83CI0n
i+HtHoh5YttxeRpRp36kXo9KT2IGm+Nn+u7TVh6Vlfxtg0ZGeVetxLKxGUkPlmlJ
mn1B4CtjDEZ6PWToPG7u6ggjbkCKY/SnBsA9oSxrO8yAFzS/digUztQQruPJVQZ+
uMRPayGpmg0Up6mv20N7YA4Tb/SFaRylMIdVw5zroMfWMIdLKxJuTvwwJp2QmogJ
orFbvEmpsj/7xD7SZlQJpvGQhg3bpEGa0qraivEZh9QeUF5yyjTIejw81oobg4r7
z2ZaNIUjnx2vACC2RGibWPymFqdY/y0l6Uyn4tr+Wz/kvsPBgRnozYzX+ImZ6E+b
I6J1hIVNaihznvSas5I1JpbjjDqH/ac6070TJjiQJlczswrYS+OtAwL24KL2bpbY
27AV2NM+d2s9fgwEHtUOgT5bzZj7Q0pf0rt7Gv+45CmMUZFyCi/LxfjZSCHagyP/
ccboM8Fh/WTezH95nrS+eJNeZvx4WtnquTho63fhUruh/2N8CL+sJLrf4cx5F0T6
rpjnm8o9d59kGE/yvm55hE2adOpO8Ky/ZRt7W0Z320gostM85xsXNkdfdD4Bn3S7
IhQNmciWms7EKqN3hcfgmn3xk1+YJRnkwsgf6W0STI7D1lB0Cv/P57arZ08T73iF
1twMuzJQ0TcNup8nUCww0MkGFSREAH0E0c93kWE99OWFYH6Gu7RezWEq2UWeOu6r
JdveL+uv5ctGO/UE3VcmbUZRsSAfcDdbUSB1mHtr768oTzaAEr3z3hM0h+YQrsyM
MxV6JtdTL0Fg1XMC49tgaoUMeyJgtEMNyX8OGPfBg9ZyznwWbzqQrEhA+jw/KCMz
LvIVDhv6eKjjjycmDC5nZCr2tE8Kf8MD95Q+4ANcSDUeSjaVdeHauvFD+U4hDK7Y
RmLRvqKUWU0w87Nn+GiyjEybW5uZUG2icwciKipjJ/dr0AjlG2xQTnQNNPufViAK
U4qGg9zl7Us2vIRcWw5EXhPBLMnY7RZboqOCxRrU+YFLJC2viH/VrEcTIl9TmP6M
3t5bXvJNFlJH8fSJRkGuV1ywR/s8TD/fL3o9fT+4AvYHaU25KcHlaFJ96HRLxGIP
xOpNLnzwe9+D7qqtW+NIkhulF2Zh1DYKlY/JOZQrOcGrS1suDOMzqKrxBDK5hvkM
pfj4IiQbn13DNnFPnoQUWJamyT73Ib4X2cJCtaFa0vWtyoQ+93NNTXVuDYnpvQLO
If2bIoD6IwGoSn+mWEv0Khr4l+l/mCPCp7IjVlXAFEVIoqKsKXToE/gONJ/gFk25
/l1Z21a8FUqHyJHxkJK3Fw7waqxGY0Hk9h85Om1fnOKCiQIpWW7MvOJFojIvb0k1
6eMs3OO1m1MfgVWt/+bxoXbDj3BbuNkXJGF71FmXXBpxF7665rv+IR4/guDi4QuM
aigdqtHCzSWZmfccaW0T3Ps0w5xVTUa1S2uQBc3eIKTf4rmt1sTH50wrfhM1MI0T
nneFgb9bjH0wCNKIf0JIsVnrUEyS6vBvQW8X06Xe7bf4TQY9fOcNQWhDqBb3tcUd
x63gGIeACBNbuZZ/LrItllIBt/rHyVKzHb1Ha1+EBmTByTGf73OnMKRIpMwX9f3h
jITgdx/57vH6XtkkvO2Am7ZWj1MRe+1hoYbg3JdElsxCzSnTEVp2E1CEw7QL16uN
XonEEqKnUrBmWMmkSvJ3OReZ1E/P+srmSaBv8sAXJquo/d6mIjgV3QFC80+IjDP1
8q8/WMX4hJagtheGZmc+86cOBPU948ci8WaKtv3P/OsF7kGSijNemsXmlfmBr0V/
6p9RfnOflTzlk6kh4l3D8hr5DcJ50Ota29CZSBgz+eSWeF8UheOgR5lHqco/jI+V
muXFsRtU77Z08St1Po6VlGPFNFfR+YPayJMk3xmJk4eUygZairxhMKOcDqSH4L/V
HBSOfnzN+U54K86/ag+sWu5xCV2s29pGRmB1jKB1IFUaqhAo6Zq7yz4RdHaOdtVj
Ys7mD0U9h8ceh6rYtzraxjoVpugdVJBPo3YY22KDIW4wagMLoLHzsepL9DrP7dDN
plpaIotoTXuu2tHqJITrrZ7BigzV6OoaYc2OFZ3clkeyQqaima5P4YGDBd4oa3rL
HZ4omI0pda8sJAk9Cq9y5E1ChdlXSN++FKthrNFwrSg3LBtzv80Z0RE5F1hcmOY0
Vhh3DEokNTd3ODB7X9DAAeukxSmHAt378vMePIkOqeb43M5zoo7heeIDjSKXfytC
WN8IF8PxIlpWFRQWONXjjPXIvOCRBLKblEvN81dnQOpNITpdxlmxvZ3WfED3lBGv
TozoON/nUtOexPjzM7VRX81Jed0bGK+ZdM/bZi5ppbX9nU1oYTRoa+mzfuiVBom/
w6mu+OnFPimre31IcOXfGC/tPz6Rkk8T1dB/93reQ5vUrpLLZz+ucz1vvYR5KurT
7oxTzOTz0yGDEjf24+/saJMHDSiejR5075IIQvyJABu5ngd44lHZ6biJXdCNvdwN
WJFhCjSQSmEVgIr8c4TBHSQfs9PFZSLxbUn023ASAh15qdFHZ/eULlsg83jL6el1
VxncuHsKmeIqMd2oy7zT7GygQs/tkQPpFPLfRJYLjCLQapQgPg9Za+yjWwVhS9ol
YuUMpvqhberFBM3ux2w8iBFBzbMz2buvCBa0Njtr5n1E00tuEPgCWuatY56CXAwD
C75NAVzhKK4BxIfbEN4Ot5teJhVsRq3n2se81y0VVcMDfIJDwerItgIP7o0caFqr
9HopVr32mRc2F9MTooJ/yMK3jWmSqaORESC0Mx9w2dcQ4kW3mImFMfO8i+3Rr+Yc
7nCR7PZTK+UUG09Xrf5Iq54BILy25QShHTolOasjHG1CJ/7AheO7QDkRVn6arNZq
wUZ0vobn+rW2avDOZ7qjmdeoGGTKxuIBVLvSJE27d3F1i0keFAF7IgtQ2dieFBMq
oS7a/npMA2uvY8dK5MnU6+yx9RBn3SuNn+QUsuZER5q72mXpc6qMUye6WNcmibUG
ZcBpabdiSWMacwVUeAqx1LbQnfafGGu4EvIid0szUYJlA0VEljuEiNvitNOAzrYP
0stoFKvL3LCZ0aGQ/K1OQEGGu/mA6FkUvzP2lvKkPWFlsjcmLu2g9BqDEqOJkMsZ
PvSs3yAOL4n4EpQdhM50UG2VgraE3xt8vNB70+SgF3jf6IldS6YTuLlfYaYpoR9u
bEzrbbtJxXsXV8ddAZaDRWosAY+ElPLUUC5jLvQ0N9ROLLRZnjgQkHWX7np309PT
UcFWJrK+t83jjBWUAUQ2WXfl+g3HLPIvMb+uZO43+aKgeTc4bPR9PONYgEZc4Vfm
HR7U/0WiUjI6myFv45qcA64G/UOzSECKIw8pZF9rWhXgPaO26/psBOGDzV5gB0Ew
6A6rIY8UKlGafy/2uMGqxbwA/YI1IstXJlF6fCA3hsQDTxr1VE3SRb5X4DgCQaxW
VjVIUedcNu26W/sWZZ8dRc3tHauOGIBKVrgGua792ZSzg8fH0/BM+So62oJOgpfO
gkXZV4sCuUPxV0i5irzjdVTpIZ5VHrBJkkteFSv7ArZrIE6Qvg/ko8Kz3dO6vBn2
xHF4P85liAhkjFDp0w3lXG0n6++60AaresPWkh50DJomqUVZL/yFzGuCjaB7eSlD
p54+cp0+uCxDSTwrvXjhZSPleEe5TVkGFXAFuNMGDgCP5ehHJ7iiPAZ+Udl5vmW1
OWZcvt7pwxz8nu5nvY3567kUitVBHFVT0zqyDSVorDbsx1f/FJwGlESy0GSvJ/fh
sPxWXijQxu8BFP3buMS2QeN/K2Zq07WQFmpMe7bztmmwTcdRcnEKnh9LCLX0bkmX
8eTYhUw9vZ4mv0vTt3v2RPKNJzHrb3rEvUZx4BVn5fYyJ1sO2y32NsK0OJdAvYMn
d7bmkoMbXDjqMv4sQsZl5Jr1QqnR9FZXW+yyPoAROgGEuNvGplt/acfWtbv5ZjMo
/w7WZXruJe6MZfSVuXwfjTzKS76roXVr0vkfegfgCJBevvaLK8+TF3z+tNNZRX+M
IdsrKD7Dpvrf6jbAzCZg1hR40sZQS8hJVpZqFw6lD8O8EZI6biN2qmYRkVDig+j1
YFM8DKy3gxjs6mOMH4BWlqNbShCZcy2fdvR7kw0mPEStnXbg16TSVJsTDT2GhEG2
DcYl65/78VCyofDv+NMezzZp/sU+I6HKCTxr5FWQWvAwaA5UaL5BpmQ/jCx9cAkN
CshC9dwRnTmQmI8esiivaxSnWJpWvOJh3RBgTTF1fCGDu52e1SgLT1YBq3LxX8YF
pvHdvvq0nTqS4hqmlvrrJkNbTUmHEp7Jg9Qt/xDVCRBbbIwTNRKbPQ3h4xkycKNL
7D8yud2gl2l627rUh4eATYr0k5h5W2JSLb0m2VGxEwNlR2nNCISqk3dLQjdsHI0p
p2wgLHYBeCbxIY/cK1AmSnH2z28gX4H3uhDHQT030JZV+AAlmYtc6f5yKLbV/2tr
0wPHR2jIzGMcVGsz+SxFx9O1s7zt0N0gc3BVHJlpksktm9uQhrfSRcmEb6jY8vLf
8XLJNx/wnp8zBlEmW2Pc1HabWu1gzSBIQC+gvlXwlkbIWjbboLnvGFz2fC+4MIuL
/TP/lHRq7W0DcgY5YtPp/POvjpuJFe1iNuNwLtGu098hSqH+cP11b/hCpWGRDlQh
N5ciNjw9ZTKzxbS7NBCXaoHd/hFe19L2Bnf/A9nusOTYQJWNJw0glIjMH+hEk+7O
S/7nSFOKPLAW9iSlzUlTPBPAwN7YqJ0lBFOn9aLfJbpbfUMlPMEL+lljZ/OeUqzm
2182ur9XFNhdrWJRz+SLxbj7YKpbHnJxrKv/hVzZXYfT+xIFpFP5ksLIHUmrgLET
u6ylZJyAfZCkilMUrmxoLPRe/o7F3nTTqUpOKPm/fMGZsfrj9qL1tbO1sC8XDYye
4vfyyBlHQ3N8MJVjI1E/b7reBKw1uQ+JtxHBvkG20YDO5IfDiJb5Yq6cv4u1JhKX
Cc7HyD5TjHOSIXtH5mbGdJXjQAxw20niY2q1Ezgj8G3W+/j0/cidpnarPzYOzymX
11ttLRHJdQS5IXvpPPD7WHZCtMmDiQbv48Ulog2GI1gYImt8GtRLyi9tv0/rDMyT
ZeNa7JStK+PZaAVqmOc5yzDQwhS0uYCit4PoJ4dmt+CnXYmcIHBM0ntq5NscMtxV
aL/JlquvTFu0crrNaL48P6HdXqafBkePZ2c1OLcVlNEmtzMHmQzEJXMNrtlCTMyL
vHnvbZlq2z3RM9HAoTmObaGTFpG340qqQitfPzxjrBzCIMH36z4k+H846Nlweaeh
ii3sUleYVM3YtL7jw/4seiq97YczG+9C9yJhlh7LMMft0j5HnhQFZ2ihPSHEB3Mc
IJDDH+RnBiMdxM3QkpeLyyqt5Z1oXVa3SlVKT8VoA88S6IzF+qXKrOcAfpr1aC+M
xJUKx7xlWoyklM1wG5QaKrFi1hjxq680czgEh1a2MXCHcO8Xa9QblP6lrju2D/CK
aEmb+o9WVld3iqOYhHVSnCNm9I9y71Vpr/FB0cJlxXxD3m9n36QRGCB1QygTJ/UU
p5U1GCKTfW2siFhdfo44gF9NWca8+ilW2moiew6EyCybFKJAsOlQlanz7TZTJCfB
Gb+xN1tiiW9iWMadN/WocgHXJq5O7sNipPGgBBHJgPzC7aCku+AghiXBqbyA/HEG
I/4c9Bmz1YsscCZTS+TYErZJKqhye/rru/Lp/2sc2IvqTnxqutEXQCpe2G+Race+
u1VvJAYW527w9E3jRP88FIx3oCIwDCEyNHk0Xz+DoArFLY0gs3NgaEOF83UmD4b6
jGcllH2meTGBCgGXKko0J1bFNCP6Q968StwETGUyM3b8TOBtKKzKAKrr2sI+pOOo
4qWOaQ96wuzBksF2hlVDaNbym62J2kpqh/lc5vtsQUSBUhIAv/FFe+U62E/d4Wqn
Os0M3bI5B/0KL3gxQjmp70bHGwSePgiCjXgn0IljRQXcZ1I9LiIAcur1FQ5BILXG
gdqAFDDnh7jRRg5iV5It+MsD9zn7iI8fiYnZUbQDbekyJB71k5v5xs/RCct2wwbF
+WzSHgw8TVN3IzyEmIT6Y467CypaooLa9fA0ve5MGtOGV2MQdMP1Jph2h3+J+4T0
39lYDb9nXsnhRtBpBwnt+Ugtl5CrIYaYSWd7ttTADt2S7h/wOI7js9pWVyBlOCkc
+1xcI5fnxhs/kJTod62TW7c7QqGrVOheD8F6yFQG63dTyt0+iiW23EgXxRf43lMy
f0kgJZtVMGYAeETaXn5CZloXQYwgg+pX/DHOYWQCauKOF3yfco98sIK9+xCoSaSn
+wGnCK/uWSxoDGLD0Srv5KF/CAOPqwz50dMsuJVq3+uX0OvANXs7SQJdacXC++NE
cNJ9jxhQ4zQO0bJea+qhYQa476K2X4skh/Q4wCnGgmlAhZrDbqOL7CBqc11ndXTO
32+cWYhKFNBRvhlkbI5XwB7i248tX4pC10xZ4Hj+59/HIRU9YrwagEkENpuEqNWY
q4snVb/2zXPfe61sL14f7YXEu/S35kSr7zg2E97Qa5HiU6bs4GoK9ok06IAAd16Z
BxMUZmoDMVNMqT5WQ/i/jjD6sS6yi+Dps1odLsOc16tCN9OyuS+78zxBAO2/0DJP
i18IH6wbqivAO9m5GIJzupLO0YxE3fzawRMQwRzNRJ7fArjVN1hEmYs/FHj31OBG
Auw1qydDyxexgmXiikQVcrpemeAi70IuTa3zKEsyfd+vS4ws+7ewY/2ddxvjKcPZ
B+JhLmLLxR0YY6groUO1Adg8s4zjeoqhO9+OhPjeIPMIO+bOU7ymsAkSb9NRFknC
L5ohJQdDElDu1xnmEr7IsjddLM+mUz+FVrmVaWxS3ywB4KF009x3k2hryJOl57m9
forxuwU5599b7qpt1vHNZ69UpxnYjGd42+G8Zpp/Pyuf3kWetgB1tmqf+SNYUjWj
wfrmldrnR7a/ZJYGm4yGd7Yx3VwtIOAwIRFWdLquyrBRHcmq8i17ErhYlmNk++zm
g2pRzqi2PWjqq+oY8TJbPYrwDVHDyzrceP3D/nAWDqES4+64k4QD02npIxhUViVK
mbNJ1WlhU5KCvc41skCFdU6trpk28Y7MVcf660qlrtBOPqsHIrRtKo00qyEEWkDW
MbwxuseY1Io2mmCNjnLqBiKHo/HIP6c3Q23i7q6FFMU7jb/CEH41Ux5MCScWz1xX
dsxHeC7cHCx75Sa0JMlm038Eqg+b6MSJmcoKqj7SSS7JNZnKKIVVN7LZluTx72ne
uWiRBOo9S0wQoDTzY9RSGFFQRbFLN6FOB8Oe3B+Oo7LWatvqpEoSbHQIsAn99EjW
dIi/JWY7Of2AzvkD/e5HGNxUYEmLuH0LbXZETacT+zyutHNmfHFfVzVJZviPhsRj
scHi+dw6yUmz9kSGAjMKpomGDyPvsTEL/ZOrOHtXkQueLE+Pa3LBF3uRrInzONFj
yTfJO2aBytnZYBNwV5UV5wQTVoQNcAphIsVbErvMdMnwr+OBKrfSYk23+CcSfoAT
IVtLxpt41rnSZmABr55s8tC0dANr2cAMdZCYY8J4Bo6QLXcGdNBYVah0FpWfq8nZ
4BMCRuiyZMAQpZi41iswHBXvAsCv5SJPTTpNCf634f2f61sfsscTrpG845EAnZS9
7MGAhq3YRKjN5t3o5pPsVMALzM73vrYMFbKFLPrBk8OyUECs355zU94x0mS939J4
UX1SgXR6aPA30tUtuA1vG5uBhpkZMaBFs7wz0fktmWzyVYd9I2ktprKfySlgTL7Z
kKiMVTl359pq4E1qeeio/YuZNp+1tKu65KLd0Nzi5Z0ZfQOkvX6ZQ3xWNE2+aPq3
7nlxwZ8B9ha7DKndpu0YyBxVEG1x+OQXk1ALf6aNs/LuJxxWlqrRbPlA9s8d1GPo
8JkG5jZ8UY+rA1tJMcVviTuSJshAhXU9DFNetsoFKlbXjPptm/U7efhw9BbGrjmj
+h8djISOQG9CAjQsi6mmM4rN9ZGpo0+4lu54Aw9Zg9hOj684W2LUebhlXxzto6QO
JOj2Q1K4QDSUt12sfsRAP+m02orLbA/nuSTZurptvllWwrwbpkCZbyTyNzwlfykV
OICM6GU8OfLVT27KdTDjO76AgP8a7Akh8MidavK6014PkYardIunnkgFHZ54dezi
gE1sq34Ei8DK4Z7rs1/OuupeNcDSjYyHzgJy4nmhYHPsAWbwrGcYud4jSm4gIubc
m6rlc+Mr7dAT6OpOig64Yz6OzpijbeBnarYKH/QGvf/mDBUOoQRUWeVxT0JCG/Ru
6xaI73pnPyXTuIprgaOyQc71T57Wi7b/PmTnuCC/zhJntu4M1Ln5S7seR8es7LMI
SYziz0eed//bYZBSkSyDSkG7reyAkYLErAGsUjPYboTHYJokCCcn6DM7vNiucpTo
Qck9Q6VRvA42l9pKr1XTNu9ow+yBRPRyjiPnir7CfRtz+KSxor/+GG/oH6opLksG
ewWfxXvfLlOOEljUVZnY5RJA3gxze6a0ya5X1ebARX67MDn8Im7H4PVZ+r+rMfee
g7F3nHeGQ7LZb369Xr3TVMlq+ZI4yIVRjM1WWjMkcR73hHyvLscVUyAKYh7CQgZg
gxkgGEvkPtF7UQJk6ZbylcRFAeiZAGjev/8dRYq2TVLwf5xZDI4Q58I/BO9eFCIw
TNfpEfxt013MRaHKhhSdjszLVLEqkCINDTcUr1qa2r0xupKEspHmd7ZUW0rGNZ4w
TLv7DYMDwc9FlYUyvTK5a1VelFs5AO54recMh3dBHEgEJ8FZV5ytMCR8L6HQ3Hsr
DUODRktLi0iBHS2o0eOdqvMNlzpv7PHkNQFAJyfdi5TBxOtvcdtzkLhGlxprxH/0
rFmf8u/RHomrZwefdgF53VMV0oxXIwqZ4ns9Hcp4h601RahZ3JZqQU+g6ZlUIQjE
d+hlNBQ7LWwueIMFLvUPxrnoztu+ZBprcQD9T4E26bsr8mHkKwWdFxpesonw2SPr
FYxoN7LkVzKLXOP9qBumGtgQH5qCuP1dIcQOw6IDXRTHcfWIDd6BW0WEb0obKLAz
9ZoCQBQFrHpxGkWHbMT4z6LJXh6MrW5boEqb52kFzSHdjFs+6roAlSrv9ILiTBf4
1fubqqJ9rv6NJT0zAIoqNjdNrckbqRKqXZDLOojzMf4Qt4Xi4Qh3UpgPP0DbejRr
5cmmXSnaq5G1lDoiLqz4oNyUryXDiKFcs0L0g/4qrHEMGZBAbNS+zxqBfSEyA7L8
AsYtXOoBKfBI9PbBrhjAbn7AdPe/izWR4DQVrEX0/KiUqJw96o4aqjCRxjG7EGjd
D+KPT/u6vPvTnRrvDTw8ZSg0j7T4tbifIoW3QpGvvJGMfRS4VBcps32g4j5nJ6mt
FLxQKvwMN/6SFWt9062hrUTpZfeDCG0qxtCMgt7+WzZ6wGSzANna8pLzUHfz9R3h
4d+qS3eV/iZEjIb0aXjPCIEfiUMnsA0RlenViRep3k9+tencH7eQE8ss7+n1D8yW
Qp3t2pbigMJNF0rBaM6s1cnLf9GTk+IVrlXOjB6LiZU57M4A49WheyjgwrmQ3+p2
ZKPfHSFjn5usTizmbBENEgyvVkztPKGBWCFPoYAysdIkYxH+5TCxOIr5TJaHMU0N
EAGmltn1+KGU4uyLyYF+rdYzlyiwvQABy/ITarYYijI8a3fFEGBYTlaUsJOxMXCj
VHJi/JObjfQX7PQ/IQnMDy59zH+dOgYaycZIlZWhcXpkrvzoirGGywsRyYZ9tUJx
9xxycPNtgeTmZz2XMKOwQSr6fImzELsHRZaTBsiX10Hn/d5umc7aeb68+gqE9i0J
bF1dDG3UTtuYRo3kNXSj5zLAJvvSClbjOk5SqPwC1gTe/S/8Ipzx89VvuvqXZyYg
ckXWD9XVqpEkU38qIukT3oTPNt6HRoG/r3R7gM8DaK7nxxmLekmn1KcJyFUzWwEG
dOpLmJ9wE0CQlQd6fr+6MHU4dFe/7pxHFCxUCDOk4cTiFQ2+2/CdpDWA+DZCzI77
1cxyk/WTbbTFCGLImEIMjUt1Dle38LbAh4dW9sca4vatJISqdHipKfjUk2ETToq2
qCf9FxXr22DCI28+Ca0+O15TtCVk/yg3gYZ9BDhA/d/EO1a6zAqquBj5dP4+Cr/h
6ri1HLOHM0L/zYk+CV7DKFaiMQInxzZRemAn9SiAmpN7JgqkCKuLt6Kwus2Kxa69
eeHLsmWrw7dS0LyKozzCINMA4dyTn8BgCJxKV6iumyPZnZ4uiRYeUyi3/TaAvf+b
6NUYx5bUt22+uYhNuWED29XzPvGkxrvvmkQeoIix3xvzHHQ+I9ugBk4bTm2FxaSf
z/3IWnssLxBPYRu0s2ozhbAR12LTMZjO2iJzFgRRF8mk4mCL5y5ph50jaYjLG3id
3/cVccG9TI5b+e1w1augMBUsBbAUuEnSt0ZcYF67iiDsCJlsfubE/MFypeZ1mQgJ
zVvovtcNclcJxIlKWwYj113dxtWBSiAgpIBuwdqOcVymFvQd90+a4nndOijbfbhT
7X30u3nr7eVd1TvArDBCd4r4xSo+4bIVfYfg1mnYC07K1DEDwJp4q65Wzu73gIlS
+48gxDZd+fQVSB9aAKNpcpn235/JyoWKLeh1hvH1d03H6LS9ZVAaq4A31u9J3aWi
Tf+6rTOBvPGdTXkDm0Va3buBv5gudbYqrR5EqKFxF0sx7IoMkcunb+j9c9PthOHE
JKpuubor8yipr/RV+8RFd5pgDScNe037qKgIhTJoO8pT5xBVmn/wJbpt/gweK2AT
pAw8qFRjm3dBxc/1rXF+w2NSmBmmgKQPy9hmP+k2cgozKLECfgCVWI92rmjsXHO9
A7s2FSN0jA6Mk9bV9tnqEJG4FEKM8b+HLK3E8grsJm3x0boK0ktOUplsVA9L9RfQ
o8sn6fHy1BodkWCeoAxMiFYMwHUrcdqi+7OGDqyBFXSYLhlFvn6Tre4/nhXXzPKj
OyPYcpeT0lAls43OlTZ8jQoxFr7f6V/sdNPuAqXQnNlEJfgPAj39NaK9hvotWS/r
QnVYG+zXZXZdsSYmpicD6NvXL/kcfMuaRi7uLW18t0LuMxv+yxFj1yseHJRaH2u2
A4Xjn8k06+r8/M+A5gh4ALMF6Eg9bk2r5O41N7K5BDLvJQuqGcgqNd1cQRBl0s4h
o4nZZNoOQPxXWYREru+++zMuUp1m6ZAVncKjjqJ+c8/JhCPFbj3TfPZGKMhgqiMu
fxcctkKEw4gK8O/1MB3exU7QOBT3FwCbiLBCK0qJBDkyJqbqBe7nYGPt5kpf8khI
EZ1Tvaksyfb3awpCy4d4IZ+0os0eVMOv2IKug3ipKsepe4foTRlErbd4oEFxk9EH
kKtHVmmJI6lwhcv3VT2cdnliH579mbCIMnJ+Hcaho2X/ywSlapVl5cRW5VRJ2K0r
SRIjxt774QIRxJcZ3X6yl605my46Q3CgcZILUV8JUnBr/TA+5qSlyuFieo3u8wZ7
t7Y8FTsZLNleRXqLdWmf5dO8JTY/UFYfdKdYFntOf7i5c+3iwaoM1Zw3pHKd75z8
1Emiygd8Lv8WEQXdVV0om+54XOkIAEV+O8RPNQXsG7gwW3j8tEQ5bq4KB4cm1puZ
gVv9Np8kJWMOMD1H9J0tTcLDbyCzKUp6VxyKEP3AR6vCa5jyM0JtZo0AGXKUNPR8
PO9kl/NDF6PAAqKRwJKO0Vr+IW3gJ2niQrraIkyA7vXkqQU2Ju5RiLx094QB9g6B
1CYggqiNz7JiudQZPCYdMhg1A48Wlb78y1AD4xr1vYGqx/Lk4uT9cPY5nXWSWK4t
9y3cAyzkoZK3SEkHRbInRkJkqs5kOSMU7HjSkF8GwF1RqeBQXm9Il+OZ9l3FJn5O
6K0snu7/OF5SHNsCfeIOjL+SjAftUjYxs38JesRp/Tfo6wYMVGDDG4f0Ahhond/S
w//ErqbQgj84p3/taBEv/ipKNwJwNoEu3uLmOqHg98t+aCbLVwL9s7vvQBlFlap1
ZeH9HkBgTSLgTrfj+ttXSyDfLo+2408+JjQFBBkRq55+SYvKIwm19ghhVtBvT4bz
9JquHxcd2w34K09oyWWNCzgXajRFFC9dC3PU95KthGxXZpKQlrmp0xqDt1gCDM2Y
yCmVo4l6Kc0jdSUZuk+bEA0wlQJX7ybybzu64ZTf+nrVCSbjnbdb7u23myReg1R6
VgeBZROA1i7hrQU19hE5F/7rAkJKf1xspUMCWi6nHsMBJTzH6s4XhKdI01XuLDNU
sNR7QD/VQOajDgrWn01F26IQD2V94U6Bkn22lwMQM+P+wPtUjFJ5p8pMUuhrz0b2
jYkMRCGl1GW59sMYgYUMqwG7Fjwgn6oiXeWHDVbgU5vlDec6jgdO7vCz+Y/uF38p
Fb/lluAj9+HK7PldzKGCmb+j1NlBVeyiiFD3wDGK/neiKlpEN0cUnEoQYA6QEZBH
srviyuuGno5EM8oCH+LnarW7cVPXuxXF3bYdxHnZz4RXqO+abyleHDaWoQPq1Imo
591AMwhYB5q49RDXZ/GiAoF3f8VNLY0ByiYN9lNH801JxKqEjge0uv5eGpVCjOne
FPNXcuy6w01xPfqN86fpcmSnrf2caOI7FRgGIr1gokfgGQv3T+JqOBZvJBabyiIG
sEzXRq83d/DRWy33CIBZk/vCApgZSSQ3zo+ueTs4WZa9kTKwy5UGDwJ9iLBTMpO1
S2unUG9BNZ+nIwR7KWqfbtFDvgGlIhVZiPQHWYFoaUtNHHEzyy5uQ1dvGSZXrCNZ
91PuQmVdg5vN00Zwm6Ij6vPnter4WkHRge9uY0zdWQj0pQI7fEZgsdOoUj158Psa
YmixzZ9N68I7ZH6jHR+jb2ZrGg/jkS/WTTbnpmnKzxAegnRn4kzS+USvMBh7c+C3
X8PtjoFM5K9XUQ1nUv2W96ji3LuILdREyTZjxI35eiQfBzh4Ar/XM3O5KhNAF8t8
D0v2LA7dF+lNabTo8hswpNMYHWwz4emzryRZ8gcTOu3WfwVk0YISMQJUu/chyrG9
XBqrUHe0YtnHihjxIjgz/LebREK5alAizoO1LdL+MTm495CtvMRtJ6pDypURHEj7
Fs/IIIYc1O4Z+cccZZdOOTH6ZwAH2MntzpJRf/fVd0eEJcu0SJmxrDbBAKSBGEgR
8ibzRCXVFA1w2EV9imF6p65oMO4bGh+OSIEfTCfowmU8w5/MvNrOItA3ibAcxcKm
OctSHszgt6aLprJvzqzGdeMnu61/+zopPbsz5xB6I+BstVsIlRerAJB+bsrIRxzk
0JpvtgZavckqSmr8A6t/bewy32G9plNROlLYnGX1CQaLlJ8y7ovN6oRzqdbLh7As
QW+ZBKyxQvBc3+VPP6dvVHuXgB8Iw24U15/Hu5/ocL2WZt2fREiGA4qNMgRm7aHR
xXgD+M7C5/x5+3WarRMEgBV6JFVP18wOKuOf7wXhdN2yVRe3xniKkd4McttNvfzS
9RHIUT/7o1mMoOvxdO/wLOp74nDPvauvO40TgHby7RzkNI6NLy52Hv2nRbsdomqU
7HYsj6hVbqrFy0j8VKmmodvtL3/7X9mctqiPom5xh2SEm4yg04chyOjQ7mD75Q4k
mQ4rQEsCmssCK6lUVgjdDktd5zubNHTA2xXvo2z/9cSU6SwmBnCTPeiC762BO/zj
cJDR/kTJ6Pk27O0tcsu0wGgIbG8RGfmveH26Y7fA8xeREW8+Zm6UOeHz513X9s76
3kQN37cKXQg508sUlqARmLHpZMGCSXX8/odTU7ziK84/5KcKChH4wUnVbkuomCG4
uZkvBs/RSQISgAs1ic5Jbxj+/DrepDminrIM4Ea26cftMs2qL3mon/1L18p6wUgC
aw4lO/vENXoplyXFM9C6rkKEXNtN5PMR0FCY3K5uO5x/n8J3beX8eh2YMRjT7LHR
p8DEx+QjHpSPbnnE/c3QUTbsbgPdWaqExgYLa1gBVqRF8itYCSHuFjpi7xvH9ip3
HHN/qFh7stCpU1bqeTfKpHXH9H/cosgK2nc/s9rV9GbykE9GXIP4xzHS1vLsW2bu
cNueem8nyY/WoYE1wjAwT2bal3kYOUQOCYqLCnNxjBZU+/8belkekWjEU0QWlk6V
22ibbJWRtR3WUhwzabQZ29OmpW0rHc/VnvREXG+HWYT+MQQZFwFv2w6MALeSS6S8
QQEemJSN4Vls2oxk6b+5uO2Iz8FWtG/s1MQx1eOqjrJOnOQw1kgITaJZSY7k0m0v
UOjrOpfTcfJg8GswX+3b94Rb/sWe/amD0h9x+rC1iB2AvDIHiqWbjDEa0oenPbkC
xnDQAd3t9Kp3dq3Pehkp4KJDFbIeb4/ojw/74zS8tiU35WCOzXS5CNI65CQyL0AQ
OLV4YqJifmIZYyGauHilh+bpeDnM17Yc1R/JdyJs3PMf5+OP0q5vxArVU2ar9G56
8KZwLERs0shhP69g1+V1NAOWpYQFVaKps6Ve8UzIi9aQExU33Ft+PN4jbo4m8OVA
J2+MoUT99OmfWISAQHfoZBAInCCS+MoTBvZYxyOOT3furG24Wc+U3U7bDpX4/VI4
Df2eQIjivg9MSS20kxZAMqu8ZQe1fwDSnIci8kxQgr8A4gX06HsLVNacPRsoeBKm
jI1lIEqOq0TcbXk5E7+K+ag3tYjvjL5Dgm5QVvIJ2qP7N2zssV7abPqIAnQ/5C/3
HpEakFTBk3pB5rCj8PU9HzLAYTaHut6w/Su3/wsr84Erak6gNKbndEwfERjYNQu7
yX3/cWRkUpptTyRTTn9z3dXmuqEtZBD0gFND3PFcfwso+j+E38iOrLEoNDb3DL/J
dsd/v/gCMyZYYkYOF0EDQXCOAI6Hmq0wQySzCXKnAzTOnaG1Hg8H639/rT6mgEPz
3wyi9sivxh4Ijm3ncylBcSp0OIReQ3stKy8HqEH+MXQHAkITtF4i37JI4YV8mFc5
SJCcnY1VQuz8UnbQB5VV7aUJwsuwArMovoIJXjvwK59lUiIFWsWJD5wB6/tPHNSr
vXgqnWTvvfFGioSNj3I1RxgGLYb3KeF6zb7ZLkPjCS1DUefjkfKFQVf8E+gzfDK9
VYAz1W4f7l7BN4DdKS44/LTQlmJ5HDhHtuXXUpjexPe7t+/hng/SXfKU0mGT0qEw
y/waQAPs+M8bA139PjZsds+wRY3QTmOWPybWicR0b1PA7gCqePjGnZdQIGHfS3T9
7zYpTiwS7ZyU/V0O8I6aUl/xxT+AqD460Ia4NY4SBdUTe/aNn2QaMjlgkCqC5VSA
4WU+0feNQ+n0mS9ILJLggijBJwVltOOO08Jg2MuK7LcGoG1neD/rm6vBCRwfwKEy
T2Q8a4RnmCC1wvMTqAOpOgH4dtBSzTgZE40++lmpmR/VqlbxKb/mwa4Z6bRA5NKM
yE5DoNTh1ObDy3ZsghE91dSfgHd2ifGAbT18igjoyxjMK6vZmLsG3wK10yyU0XJ5
NxbmXjzPhlhIIkU4+dPkKIX19jIF8TV+EWG2KRwK9kMYYNfnuGejyuBHHJO1H4OF
71Qh8C32Ae3AHt3dpmfeaZ3QNm/w+7i2jSMKaa3KRBj0X8JgUWoQvkvkq6hjn0zG
IPc7qerLH2pDDOlURGNbFCOaQ4eAaIBNp7MY2Iaf7cg8dy8sxFcPJ42EirW8givD
o373mIJRS0zG7Q9GP4jQCjIZxv8gcnfdK6TZ5LAQGCIzQieVRj02Yg9P+hV9iicc
CPEAtY2FQopATREXFNu5WQHtUrFiCSAg4YT2eXpFb0Nz5YBJVkgWJP2KjjHWA903
8CGp4vx+GkZY6eyfKtNQB3wc2inpr/w6rLj4kvqxrgstwQ088RnwDkH7sTtKTmvv
UqwLpboM3IITvyVm7/6OjkHygU31XNmk9o5r68TtAnf0I46DP7CEq99f27uI6IsI
haQx14azlDdYVgy5Xk4MGLFguR+b4DNeU2aHDoWHTGJc9IJBesHaWWe3itSjs81n
x1Gfmtf95tkIXccK9MdDC+227dAvrflFKYxVAOzWXELUAniTWhaDA5+v0STWrF+H
1lRr1jxeUvVvfp1skB7mdcttzRCNpHDgQRZO0agqxA8mdsDCaj8g1u/v+w5Jz+D4
Rbhkq9cWMIJSppGROQlCHit2oMnuzQTB8zL7Fmd8B+xzb1t/F6S2F3gnVA58WgTm
e3itX9PJcZNXrg5rOuQSWII4M3qeBhpPyQG457/sEm2pPuCYkN9NPAeyCcnD/BrL
IwDJg7SYieDEv1blHh3A+gWxV9zmV+W3dotoibvvcJQSy3iX07gxzMwg4Z5xF7x0
kzNJ4JtrXyUA27MVENkFPc+UMt4IdmyJy3kehkbY9ccs22Tbq0YG2EWZcWF8BBiz
9kHMQ/nnXBZ+7RUbWJvZ7QRt9nY+Q19TtmvG+QEaIy58j9HwosXLXfBwzoMu9rja
/ygQu3SLf9sR0dgTEIsdm56TaJ5p4hFJzGATYsEujY9FjrADtsx5nB3eCkqBmsyR
Sy5RY/Ds59hlrA+3zZVESpcpdrnt5rqrroshSN+niaw4nW9vvn0O8Zsn/ozBzK+9
oflourigCouGIWvIZHNcTnJPPMCsmJpNhYEP3qyoPIGUBvFfCST6YVpjA2jc+/oC
zQiLXShEx4gFV/jmPyRRcPEBSvHXmzDXrKt7/f3bAFlVJqM9SAx7lOkojyfsNDuv
x86Lj/fiQws5qV6lj8rVN8ieOwOSdgwpUrnZPaIiItax3/+WoS2qp+x2DpJj15ew
cEFj2pUAP7GywPIHuyW/KvbGKMeRJDVarlIA6NIZI0OgK08Ja86/eV9USq28/4og
0OiMe3WcqUrrh7v3qI23IkhnVEHipTUOb80qPeUlIFHUtAF0jH+IGA8B+eYDJHFt
HriP/jzQ5R2eHU6cMsvw4Kfd2GtI3khTWAqHP8nsgwrsQZ5r9ED3oW6lFUwkrRIx
Q9tGIT6tGHeQWSxfYn0mMJCgvGj/8a+zbiIHnHaRaa9+6nyVCJHI8/c5TOjW0DEb
3qqztRe4tI6IiebkhrRkbcp0vMaC8WgkO2bGqVTwj92Bk9qt5Q20Gdq0by5Yps12
iUjLGjzsKirv9qa5vie0FRi+xOjMBru/Vxs6Ykb7yyIknAda+RuzMPid9urqimxN
5RpRq8JYHjf/ZkwU8S3jpnpQku0rZJSYStCOV4M0hZcNDeRzPsf2N6DZ8/rIB7M0
KS8BNLyQDQZqYz+JVAI9OALk/hhX7sGAJyMSNPMuTvBXL/iOa5M5ekzj2cerpSWO
stcahhWjvYaap8UOIoTLZvf0+AHs7Hdu1u7EMBtA4R0mW3wwkopChTV86TRtcWCC
d5VYcO74w8r6h5269wav8VUa8ssFeRIQkFbXjr3hTBqazdgj4TRjjS2Zez7hQqic
HKuZXtt4hnGZv6N7sgD09Fkiw1x0EXKjsWnQLXrqbTaTpDZ8licrRi46jWYo6RNl
HZyfzR4V1H59C/PHMbGAR3h8EqV4VvvbslrWreVw8K8awD2v99OxsDIP/JvNO2gz
3g5CWEbq+z9H2449JL/7nbOvlGNAxVAIoav++Wuv/v1yZLfs31dwoBrPXjdQXbc7
h6gdJ/yUBUQxGReCuZc8z9Rk2rrWwOx2aeIbvkqaYetHLNnj6OzwXTL9SbHybSPJ
K2mu1A0un8FYKBpNG58gHC0J7yybAOP+oK/nvwdk6+5KF53on/K/II84vp47tAly
8CQJfw7Tf6Kk37le9R5jH9dOXdn2AMG0PtgErxVfOyfjkkpf9L5jpakLjkJFp2ff
KkGvrp5eYjHNZfLU/WtHTkWYyDEFP3wpTk4rtWPJyorJ3tRSIPamNdV4g8sE+BBN
FuwCZ0J2LroIxw0gC9RoCxbGT2K2fSjykSYWWpbct2uRyhCWKUrNbw6I4uTSIo6z
32OoanetzrogCOakFU++qo9NvYBOHLcoQyzoZWbrfNI2oxsWpW6HtJexQOJkrPUf
kT/8/BNzUuOh7qJJHgVdyVEZ3QNZKhuS1d/TPJtUqHIb9m6+z7E06jGeWhuoSjLg
cTiVqfRcgLx/J2DdfAIG0X/CZGemd+i6iDQzS5hKv2mHQLtuWr9iBfjqITe6IAyc
ULioH0NJ7goc01aMAuXssLT8mLbUAzSf2YISf5G33TET9H+OwnkucYZCCBbjbX4k
/aQ+GvYc53Dl7ijG5Y0WywmMtS4cns3VY2ewj0naQrYh8U0aHHRB6UPinCwyt4z8
uTnS4nekG44Z68T8vqUMVJo9CEd3fOMCld8Vc+T1pU6JrfnrnjpnCauj49kwcT3C
YSKSNrOiYvex5ikDt5HKMkLuFLyfh7DPP375pAEBSIlvL5o9YKg4UkwfDNfTOG41
wycvIHO19Ip4HQXFXkvIqt9+irnMPHuQVi6F7XC3L2wwh2ADXnalG4Qd2qsLddXi
UYZGqVYVCHM8yEiSdI6VaI29Z5RMKh9mNbBzW6cHbG73KIUeWdxEFGgWHLiq4xKN
u8FRzE6v5n+cOLzwtaDRJgCmBAiS+NxdN/YxKJ0UDAz4Pq9okdXmgeglu1O3lQva
xldBdl5V4q9An1x/P4Jlfp2L3DJvZ7OIyyJqvuluR9tUDOOzEkKSKnLBeLZl2smP
oYl8v2kBynkAlBfm+UUGcbGKYeuPLBgJyVK81v6Snr9oe7tfSgLxlKKmOSNo8iek
jKpuCe3cY3GgGxFxcmoJojf11kJQfbKiBtjgYUDVUWL6JAemRJ6Kh61d9er36SRK
aqPQPGTmUDaiXD/zkGcfUU8N6i01ge0bpucDN3RvTFR2zfqwR7p7xB/Jer/C8QJ+
1Ehe2bqg8ykySA3lNn73tL+Y9kq3A1NjBEm6SyqkkJoc86PUA+0HAt2QXadNHaT0
DDVQiIQxUgUQMvpPm/3FfRlXthKIqfYbpjhCO4e/sjguGGCmJgoZaJ8P4KwSi1qH
icFi1Y3JCPVLGnC3R6jkdh4OIo95gRN54qnz1YP5aRbtlhP3FPoh7hcAw8iVyog2
8tz3LZvpnqsQtnS/XnAKkAYCQbXyabPZndXqazHXDl40GLHHAo4WPheiVMs0MhOZ
snCfz3KqHq2X/SlpfQBHB7oqv9tnDr3kpoG6Pt3VLo6xxtObcX1M/MoEtD+G/9WY
OXp+hZekBwdOtgjdqQ4PZ/1vwyXKGfwJAxE8pjM34TUrY3U2YDnBUqHoFy2LBdgQ
f7BRi5IDn5URsMeku/2qYdO/uksJtfkwgacxLkG+KdBOJgqn4dslZA+E+VFBjvt2
yM3nqbQbtf/Nie7YFUqngpecvuar20A3RrviQ5R6VWEFmZoY+278jY+Est7E7xaM
J1JNN2JP7+dmmrhzKQpbCNFK3Xble2zmPBXw6uzSMagmY0qnDzQomxTVnyVLJH/U
BWgRduENfsHRNXrfWLjhKZkROgw46wBzZtNYPY3ZR8SBwedFYl0O2zUoGxJ8yBDl
M78gW3F7HWzYn3MwOB47Ci9QvRqQx0lF4etik+9mliYWfG+bGn3MsS1GR8JYdA6z
9L9FblGryxXfhvygukq0pJEZsLQ7aYHarg42tM/EAwXTq1mwHH3t7x7hjNlu+ceI
Qy8PzZ4xMDmCPTa/tHP8gLEGOMWonQm/ctW38hCENk+loZdgPJIih6eezYtwwMVy
CCyLRxdcCI0qJ3BTplAHhk8yRI/XBkRFZw3D5THTB2BXOls8t4Y5NqIKp0ktns1F
pe/K/tzFb4PVWZ5Zo2kAJYt9dJTJDvFW//moQ1/qlx9Mq9aSEH3OvG15Op/i0evF
h2cvr8kR5VkFF+lc9vs9uJ5PTmpEAqc9zL0uRIrlhJvryjp7i186ltyqm1kJmTA/
aOwUY8JMKGmk40R+iTMYbQm1Ac03upDZbvZzfZTxJfDftVlDNffF58TNHWpI9HOD
0Fr6iCPKBzL+9FfxyjsVv9I44csMRucaZJcxpq+K/FWDUGB0xfPt88mrKWWBfkp1
LteQgygvk8a9F9r58OryX42hutT/MOfCaip22+oYmB3ncQ4dXLuNa7JGQF8QdCAX
lm2sgeLkRFZnCY6zP/8Tfc5DvnaRGWsagLjx874fryuub+4e/byNJG/4nDhB/OkS
cGjViSNdrNQ3DbEACO1Mlz81R8mtXwKhJm7lKjJTt1c/9XwfTrlM6v+926yix/Qp
Fuhb6/0Cvk+3/+M6Ghyi33XEc/tusM5o7lmQZ3gNa3+91yZFQRlY9WrNoiibNKjZ
oLKMQfZAaRHMg/bCGvJydEGVqM3vGcxt3AncwFbIUYW/B49cdp0nFd85TW8OZerS
yzvp8qdtKmxEc+7dnJj+b3A219qv04WsU5fQkbP9apUBtab5vkcynGX1sm8c8NTB
hJzfelOGnmFn0rdCyyUfQXOk1vi15Py9g+WUdUSuutKlVtQO2aMAe8dF0wygvvXy
zu4nQHSStt5SMV86H4RNlDjc4cyJsN6X7+4uQDywQnw26qtvyRZtFx7D6R2H0E1k
98qi1iaaD6feoReIVj8qM4SODBtD33OdltctgS08zsjWjQGUmf3EZvDFSp9byVtr
xAGNkSwj+tKEhmdQlmT26hBY6jB1huKA7xvTry5j1a2xaflZEH9+B0PG+R/Y3xsI
uDNqVdiLKtFvwkm0RA8BGOp2kcVq3IDqgapWlwBt4pPHjP/Mq7lZOV9fge4MG2TC
vJzCxhhLgGFfVq543ob6IQIJaOaXXFAJQuOJ9IjSIRyPMXSxwE90Cw7oszSo+Sbp
lM2nfWwxeL+1fINNX9TlwlYa3AjyaTwCKm2RaPolwd9KpFlHhBf2W1Lahc8cT1Lv
POr/GSAfaer565uAwKg9MowmLdoi3T2IEoMzr0ZIFqn3ALdxQwJFz5prCpSmZiGr
BKtu830eNvNeuN1M49J37D5ud+d0EIBrvQEIiijzuBpWRgLgOwjdj1eUbGaZmlY7
8EZcpv2d7jVsYeZ6fGXkrsmIBcKx+rqd4NC4kqq6U95yRsr1JJnEdp3y2KgBmomY
hkMnkUxZwNEp8g/sxMDYJIuOAr9vK0Se4ncWQ3qC6ze2KNHzemON+HL09iIFztfB
MCPUn6ejJQmzXf/vpA16F9r8o4wBvGVOtJIOYxlGFJVIyc21uwdwYIun8nPvuGxB
b3sQYJdHhYf5chHqoeOOCuQLaTrP/26pkbqiSW90OBpmxGGbkSVuaWdQdq6cO9Xk
VTTu0ZbAZyxOFEnWc3oiSJNUC6eubvey12vN0IY36FxR+i6/Oh6jZgE3jR0912Nl
9bq36fdLWxYJsEuB8HkulUigrpjQUUOKQIZjvTYS0zPhdyNCm2LhKuUsVsZ/Npmp
TSFzFlxVXj/umrzHJKeCczW23cnGNlUkyIFl8D4jJWDD/9449iSYstu4uD3f54l/
RYjKWePz43SCwfYFm+R4BQld1h9qZMXfkRdxLaULc5j15IfOljkxgoEe+k6mXHb7
0rN63rHT+MsgZzkTNzPY3CA8+SzlG2l2rno0tUMAZa2ok8O3tIr+8YlJph4fgvkk
1UDuuGUg68lfjjQU6ebOcvumSF5TTeJ+tXoDUrRred5ta3nnEUxYfBYVwGdpkEGs
2V6PdnSt/iRWRjezKLDjfmoN9amX0OP94u/UrWXgVzJhPm0MJWsX2knNRd0A+j7K
/nU0N4nZtNfBEStsqMw+O0Qj+t90MUBL708eJe/4dd0CVpRmpbuywq+dZru18fDX
9e2FdYPZpI2LX+7Y4dgtPGHyaWkPKK/eY1LJYYwMwMkuCJQbrY1bZNDj3qIy3zRG
CAoOs2Im2yXxAQQTYo+OOkeHJjaxt01H+7O67CbaqxChRjuEcEIP67Ea+o4rIkWW
dY/TG1YRCQ4Rrz85u9FKGV4e+Mw7zv/6Y19ZXUQtTFrDO/iwlAV90yYj4iOCVTSE
dVFkXcI2X77+YNtsofNYdFxVGRtcsw9IvXQWPNeqmBtevfMtf4upuWkBSPPTb2xF
jXut8bmHNrbr5G9BhKHNE5XwXJJRHCaApxRYFwXE7oFNI9R0bBw65DbxMsn0IhGy
Klxb/CudaM3iE3KO6M+H3258vcr/4D8GmG6PQ17/c3hrbJk92cUE6fnResR8unYp
Wo9YSQ4ev8jX2ixDD0vionh3rxQ32Uvs5hNhbZywQRbbINnXe86CKJdgnidA44uZ
mBbwhI1xGt0/BXH8MLDB24pEsLpe9xn/31Bx4dn4mXdJDgtKf0jWzgYEQJc1h1/F
kd7eMU1NJNAW4nG6tjXB6hLbRCRE3rQm+tRwBpX8D7cIWelPGk6qSjt5kfubP7eD
6dqVZAfuJTSfD8875ihUEma53nPXVk2ndjE6URf+ktrsDrMPg+0OrDOMLf8Y+sZB
+xroLqY7XcR9ULEVCCl+1bkGnmfFlUErYsX004NnDHtEp38KSYExCFaX7oZgRKlO
aBsAYRylFMtznQJOVTNqOPst0T4MZwtjZhlrJbe/3sj8FbM8W0EzIFgDyqYjKvyB
ADHcOrdF5WdlOaWPov4ygFvqRFXrE0VBU1HO8dUttwzAUbQA96YONb2KtpTOIZvK
2xK37sYK3igyYzlHXaNQp6jiFrXlJ9oxo6gMcFAkKn1eWzjcKXCFy9EF4RqbdA1w
9FMhYbHEtMFOKYleSVLR2UrsOnP462CQS9QjxIg8EbeLJOeJAx/1AzOdtrbXHY49
przVsGGfqe+P0UQkmtcHPsGCsA1uqQaQ9XrBmfyP8pIHI82l602mVe/dJewTCdRH
YFiA+yY2F5d7JFucS7iRlbYIE7dvY26YFbAAVrikeeN1LL+m6KbecaJ6XUKT8wcq
GEAmZp0ptLfdAWkXPls+xqqnRhceiOrc11/ZYdSHhFQh8ZV7itXWyo51dGzcU4SQ
aWmevbJWJdOhPDP3exl75HA1lY/afBigcIwSnU7PfK8z4WI/KEz27pTAXJ49ngvT
ksUmRIibuEkvjeGkGgw/4uXfIcw2n3+n/Z/QfumbXPRxY9iWpwB1QRjJTxbI90QA
AJsH69KVn0kjJZeDDy6LZi0vax4wtcMAwoK+BJY0n3SReyGHTK01ykZsJ3lMG0/a
yjjcLdmQbOxwPGtE5Ps/d979RKOST0TJGDlUyfTtMx04p3IeJaQHTROhdNNYSEcC
3JT3aO1powIpGShjmRsq03nDMiJQ50lnMAa7tvNjMTBYPBTpvvfLsdSC+8CN6XT+
2d3aaaSjSy+Xd9lvOnSeumRFP8gV+AvsKrq90OKtAMVz8/p9V4ugzuwxhADahafC
C81gABcdnt34xHxpjcEoQPvWKCUK27JB6TAJgdPe/PlCzL+OBi9RGxRA+OKBADDW
KmgFQxJpykZ5WKRb3jEekmAFatFiLG+5SDnRziMlKi7+lcoMnYWrk1X6oafrUjLq
YbE4Id3zPvcxjOUYixmzU0gOG+VVGTMhx/yvWleq3sGj1mGlinLeEkP9vhC6cA4s
jJDHFrUGH90jrYKxj8UbwM6Yti4nuPrFQsJPgK2s1dwb2Wa++XANm//FyFeBvXU8
p1PPSR3jSTDxU299ffF+/pRKYjtFj7kUaH4Mc9S1ZoesphK595SHSW/SFwyHLJ/R
br+iqOfX8NGDxfPH9mg0jTyHCELjysK+IUnUeKVcXOcE/+VsSNIYaomrkiArg1Ip
hYIGV7LlDknFYFdLAHiT5DduR04TR3cW8xKjzkHKG3okX15brviwKrmBmwFnUDs4
fF2ve8eSMGsK2EuZLE5gfgWWardA/6ohfrvrIR+JkdO93BNcZZoEqrjnEV5JiBUc
rP3GyHVUNuC5L72fBdQZn1XuZWNq1ylAhIXQfWsG8AnGmcsSrsrLj+wq/9vn3ok8
HgDZjsRvIwP2VaE029mmrhR1Wup7qmOhr2cc2esLdg8Jw2JwBlJWqPmlbjdQCAY5
3Z6agbT9QUaGudo0hx6TagTK8LMr1AEYWWF6oPsaiX72jsdEPV5cZAJoJukZbroI
VI4/01S34aQ2TcgaTNBpT0onqWHDDKaZNcTBJ6DcD1FD7ca1v7rOQfKB/27dAS4g
wwyZvEsCesk/bZyeSEcbVYKGTGeOng6b3uOfJoJcge1rfMGzcjd5jSe+LqDpWobc
fuAJNXQc9GFtk16o3k1DQJQtGSyXEBe7ERMYkMJpIRzDTCxXBhu+hm7RKR6mp57E
pj6UVnhPUr2OrcwtvIe64GfdNo5A/A9eJFULSfmcCQCcS2qBBJS6JFhV/El3PD9m
t3DKfB5r/eMcz0yeDCWPcctA+0xEjB+mtIeEz8EraNyQxOVQcdXrkXY4AAwV6FLP
vLSM/sgPRaox3ChwnpsDol3+cjxNLBNLPY4lL/c93dun/de4WSnkInTooo65byMA
PPOdNAstWCI86wVH60iYebyVQHNVqL26ILCMTF9Q1+4+Lmas6yjMD7Nc4a5iiL+A
W5sZwGmqDw8x/04cno448akmS3NDAfgQ+TDOm7uO6nNK0tkg5KLc4pHiDUjNnrPR
n3EAnscDfBG780kpuUltgG9tqejTuEJc072NaJl+DRr+mNYiElSCVYX3oU+lLiQE
5ljSVm2FFL4+g1IX9bOkkAcEc2pOdxi5FFXyQKjMprmD3krdiP8HmjxZWL3HGXN3
4aDysghgpGlJkWpimiA6zWMrwE9kyCpTnALk0eK7J5whlI27Y8r7zUcwO8ofKRgZ
wklBYPMYY1+v7ObHf12MzKq6BcdUCs9tI/BjIywx4CNZJoF7F1uIZHd6woDr5/St
o7b6JKJXT1OHTNJ2lZJUGCX3kq+71UkzRLAW2x2M/FgNIGQOq0W93cGDJ18HGPPU
6YdjZF6rq0BqWTKlrSwg8mF55qObDJe9xrnNwWAPTo3cfN0upeAYLmCqbrotIkCp
F6hVPH45hRMvIN4+Sbu+3gsRjJRxVki3+mplQNwD63faPp8awC9xEV/qX5AeSD8K
jwT1hBCwW0eS/C6Eq/n9RB8TNeW8kl+CUOIrfer9zX0plJp/MEHbsi3E8iZWZwMs
Fp7DhDE4gF7bR01tUDAvd3oL+sHTZChcT+kcpMYkGgJjhUWpDwcEKCnDNMDhC0Sc
jOl2VJcClYmwUjvEbzWFPhETFONaQ/GgrJcKUTlux6Qoj9uJHuY8hNq6RlHsq9qs
+uBVvjEe4m4alqE+bYjXz8bge9praKjp219VTQrCFhcMwyRYlQikIRdToGyqvHLA
Pi5EdV6LRW9BaHy5HBslC71uHje3YR9qiC/ebvcV8w1Fb3dSGhQSVYW9hv3vdCNW
mW2X5VLDihv4gBlw0kNfqLp6sKyIRf6ZdhxHTJTQ+zWCO0STKdOmTmTdKq/rw9xI
PuSouVnRhLoKuy+dbfF4/SWayUY2mcukwKq8i4KMQ67geuDfFC18oJERygaYCCdM
gslcXWjkOIswQYmFPxN7lf1jag0YIob3ybulKS/zmKWp/u69aJmNajDRgOWMNJut
P/K5oIXxOFQC3JS2wAam8RSkQMgbnJAj3do6WaYkdfmQ5yL3JEbs3nMq17KddhQO
jCOqsIxnXkdp6Fxzd6dPUTgz2TfW5iAAq1KoCGi32hrRaK74CdT+dxDf+45+PyCd
S+9vSrjgvJ22Fgu9S0O/7jee/IkUJ1mhtXrmQ05SnNY89Jag1nwflhABEhMXGB0V
yG16qbSNc32RI6NH3DQ/j2DFdRAh7HThwyCseyuIlFz/5aDj6Y1IsuPYcQH+YBYN
Bvan8YsPLxXC+JCQRchd6uW/4iVtJppmBxaI6ZE5lc8g47QCKLIsaqbGB3mI210J
j1nn4HXVOz+QrDwsgFl/NCkXqQC/gZELYv638CkpHN5aXcjKermLNn3oQK8ENaYI
qUAUYQvP8a4qs8IWpHbHyr1RwDMDTtw7JkwdTbMMlOaz6BX6IhMqYEcFdhZAUBPg
BANW8zOFzhwJ3NAxv9EGqPpn0Had0cwdKYN+k1rCIyxF5R2U+Ndd9gY9j0gd0sYK
IV+V1jGWV4avrRwVzUV4C5Lrmtzxm0gsTEYrak4RM+47ApIEP/YkzElx8O+QvZ0S
Pm3RgD8KShnXf0EO/yHvWdmij/621vL6TjaI6uZ1iiw3jQmDEQiAG+5S+WjQuK4N
BK3jHEuLgX1VRErFMf/5seG0qjNlMPw3ePVRRPj9MSrhHSnO3w1uRrxKbSjgm58f
8AUGg4u1id/4E5nj7Gk0ZIgWNUzSRFOaI8ynQONN3PmI6vp95A16qF5VE4uPy/Br
5yPQJSB4aJsMZT56DwebNxnve6adIw3banvAwxOhb7Sf1Rfzr1aeD4LCe21MpkZW
av79vfBxfFxKf7Y0oHxIjW5RkPJVDUH+JLmZZ/SObOuu7u0Ik1f4zf/3qWt18J6B
ELG9xpMO2yFMHNWKlU5zXB+9LJ6uEUfaJIvIg/tNmnOUyXYbMIzH3EckLeLbBy4P
UYWGCGkEalJRJHNSfm9FFwbY4fuBHl8LOKG+oD/IDEsVftS0LzAjDt+JleQSFgoO
DjJAvM8AA70CnklSoIQcIj8OUbb1sG4UFB/nnj6E/XbK2Bxq559CWdt5vpk+H+Ik
G5oovW/P44Y2ehYey/oMtyXIZU/abBaT04CXE+IhECzsYmJcF0RVWZwNCigusTa4
RKub60X12r044RZk4TYmJx2+6SmZQ6vIpK2SEmgRU+HL1UKKNS2BxKLzc1VR1B1Z
OIT+H1pglfyqh0QYNaw/YJUeOMmIPlVMpf68JX4s5wfUuFbopht6AsGe2rgoDHCE
sHBqo3C96GkpPdQ4oLs4IUxl6X5A1FsXY7H5Nm7jKgsUsHMJ07Tg7Wul1pcgxJsp
+sq7//IddZKllZRkp6atWIx3uP3wQP+gMmNJMM+f3zymy0LtSa/UhzkCZOumXRIr
bT5tTWIG30AhGGaUwRAv0a0V6t6ICcnMeY7q9qEVpV88SSzf6DqYNYfnnQXitIuQ
EPsnsYnsoYU9Aw/O/HeD4MRPU2hLmTdMqEUPbEvbElNY0xliPORGXLIvGNR2Wr/L
Zv4/1evMQ93GyBilazVQuy9lJ63pXSeKMBDP+yGd5Zy5bJcqYFxp6mnHxj2SSE5g
TKs9XcRhznXveZzgHgXouuO1DNVWZ4YsmoQvBGELQmK+HmNqShtaFDIOv2sgxN7q
a8vIb3Dc67U3oCgknZL9m5cM34wTbWQIfrLo3KoxsfskT4+GpXvxbwsPkOHxT/MQ
ywUSIoFHants/QJMvNEVZCNBrq0hWXlBGwixOZgahFYrxh1+pB6134IJ6+nlRatt
0hdjWpTChysKSVdl9vXpCLbChGFeF3X5Bob3UTG0bGFInyU/0kUqBomOzE4RSa0+
qoXTf+kMJTOPcB2btgAsw0M2OqIe2a4wnRg7DV9M9tvbJ/Fbn1pNoacYbUdC+DFK
vzeW8+xHym6PR4PDWmUuXiKbWW9Zm2bDkU7Ap2804ABoyu3CHLiFcnaT5L07ajOA
XyDdrWBLlbSWg/ZDobaauG/ghvylxpKHTJ3fGWXpjrgXeAQoAxw5tg5iGOM6SRkJ
qIw1DscAjz+H/MYoaTAhVKET+Ewg8lwFNIMojka7Th5bhoIfFOBLblGBPcGHeDQU
Y68xb3buDdqCRLEauaamsDogf0HZufJGtBLWDls3oDB6gXNsP7TIIhsR1CiJmWLU
n0bpQl++Bz6jgq7wiYBg9Mddyb4o0qiVo+HndGEewvP0pmN5omJBD9xeCuXLRr6+
4zB/b6q0t8r9anMt2umxGeJFn99A1hbhmjdnGSRmRxI+/ZuzYb7Pgiv/s4MCSm8k
hkpMy7Y852Fu4mz1La0KEDHui7MaNNmvvf1Uuy9BRsuZAiXbYXt2+U8ggNjOkYyY
wRehpfhmvTqxoeRqokkkj/JS3PrD6P4yLAbRRzaUDM7GaOXS4gCzCfDEK3b0MrR8
dX8wI6DyQY6j0kq7Mb/qF0SRV+UopU4G1kGxpVYUGbxRITCc0MO05hoFCBbQZnkt
NDqW07SEcY78knJOTLMkI4EmgOJwUc+OiOawr+13WtLcouf5dSUBnTXBCXDQy4NU
HRL6jkUhExAeWQAymHh0dRST9gAqrzIvHQTRKIRMXb69qIxKSJ5drpXFu8qwhi/O
j4DG8UWJ6l204Uo90iA8P7RPMWSN9L8KLOnlhEAXCVtuvB1uy9smq8A8K1cKO5Kq
1abdbW3XVUieG1rUtk6fXewbl2CCEpZlbxLGBGILEgjMdOSQdntohBDS+9m/C1XR
Rgl1uBEN9iCsJn0PsSKDuhslfW7ZSqVBJWLVYUkdYBFH0BD1T7C6/EVjBMHr4l9t
VptoR7NjJerYKthogHRP3TxLruzX937kDjm5befndyHpAMbP9noytbiIFLC1TG1m
cBzR7+MifrE1Jiiglt3Vv3wpkk3yVeLIC129DSyASPKUbiNe0IdCq3TV9dORvkWg
hrE7/twO85S/Y3fohCBSZ7IIGQbs6T1HOK4ShevXmL2gWz6LCPNwV9V0ppiRsnPa
4Wp1JmGKV+Mk6cLNfzDErzSSpDwz6lc1cBv8Ou+UEZugmp1DTAINmjKKzYZXxs0w
9+Y4v72BJMakcZQYSZBl9ZaTn3871NozVmSJIEAqIPAXLmz0/Rdgg7yBBmPDdgJb
Lhim+bvrGyi6K2vFVZIjX2FdNPciNxIsIJZTIgg6p1O6syxF/w4IrVQpar7t3CLc
xSGqxdUG9mRk8IZptVnei0l1LYtNjQlU7m36Vf2IYNVgREmLiFTcZv+B9ISM/PLG
YRs97jXBYS8P7eAvk+XsQeWtoIbSGAKkKLgd5B8YvmytuL3pIAmDLFoRVN4oZthu
T61UADEdaVOJjFBz8AKx8EtbSu0BDN1cNj2U7kMKHP+M+NXOUp8kiGeSRym0DNh7
/m814Qp0arXZGCsAog2WGGQNRMkqq+84vChiBNCXRXZX4Asx/7NXiv3Tx6KT+mMk
WSVcTBl606G4wieJLlwK189V4eDeH6PsweH/LdfhiS8FymkHPrB0Lf4RPKS3eROu
Zgj7tCKunZ6S+mKeXoRYTRKEyn+CerHf7sOd2N+YAgNPt806DDvZKGnZ9+EyvRsV
b0Ei5jbR3xPxqH89UUEVaHUjgKeYjoXxkAxDEj7mcLFSvnM6/WOtWaBWpgqsM2a8
IrbStNS0nIamS32TTI2GqQopJWEhmFYUusaNl2RaL1iEbn0K1gGppjUP2O5lOL8n
0i+HBUUesg8KJytBOH5K+ZdTsqKiujjmOmj35Bi6TXqUMFZfLtTZomyNIWBSAteh
bhqYq+n45++sYKm8RtTiOAhZTrujxcJqj5uB8f3TfesNB2b3OyzIyrmPLc50qjhQ
G/XCejZL2QpWB83C5K7bGVmO9t/kAuvp3BYBMKYBs6/LM+SBPrECrjgfhWx8s4lw
T5oZuJh6+AscZ7rfuVDaZYx6LgYn9YN/9qGL/olNiJ9rHT8SmOZDT6Z77hNflg7n
7J/IJ+9exyUDbhaH97OwLe7lJTsMdspNAtzx24VABW39VUtTtG/XdFNemqq+NIV4
3cLLxS6Hpfaqse+36rAQPPpO2x8KJahlYmbzKKeRhCERjBvN53/k/fg1J4A6n8fQ
mlWbyJtfX7GPkQUwswpJOzWsWnBk/F9IDcnslPXFEjFuiCN33hPW3pp+Cg0WrooX
RcrfGuX6/oPfP1gm94O4GU7YqYPIA77fCNyl4ZiZxORbilhUA1Mp9+SGI83hOstQ
18imY/6CwkFnYZSEMzI0FBYH1H4CFbhYkkKlyvfQfbT7jQtvsRcMXcEZN26ikiVe
iSFkn34y3DBGia+03gSHqDY6KBguJuAGrOu7UmJ/cyhjRXL0Xpgp6lscHrhFLjWY
dN+0iiU1hwUYIzHcmrmXqfAb9a+T0r62dFZLR93vB5d+mBFArkqnPAP4+f6RD7zT
K9VAlJzxvx2wBit4sCri2CXk3XUORXYnNQLyLGc/mu/qeufUUnuCML1OtKVrsLUZ
nXcjY1HBVuWolw3GfuMkVr6S/RJ1nIB4p9l2qwDqfRmLBV8ghq7oKTpG6HlwkZf9
5t78d7PdVjPQzNEbrENS0Zn0aqTb/au0PTxC74VD5+ueirPFO8RvEeBE7pk2z3GV
/4no0d3djs54th0jx3ZnJL3khUAzjkjOHnmw1xngYflKlzmH7UYdRk6lsoVVPeMW
UyUdt2KMwVD+1z1xtD2ekqq+vrkVbIcjEyA5WkMIKtVUVF7bXLR5yM0huJ5N1tes
P4AwK9VgHLztdJd5BE8FD91rEoPhRY5ijPKfkBcBnEWsfDHcaKKyn+k46a+Jf9XJ
JbSUbBJ4rPgk+/ARLcTrvXNf1UhkCoRGLReVZ31IWC0QbLJ7nahvYusAn9fBkhPy
yiYU5ptuyTG53mbQg8jaNB3YlFSo+u7TC4enRcBxKi60OBtsQLItUNSY3DfwMxzf
QcMr/9drlTcc+POxJSSQZnHYN53vS1LxWcijncHGvyHrT9HwK2tgMjXgDxk7pWCV
r+ftBdbgHSD22Yw3EyoESGLyyYgEPGGMBAhVkrFyUcRXin7vdZSmkUKCInSN8o5b
R7qe4HDSNsVIhnZmMqjBUOizCtzykE3Ok1iz2/5yQ2V7KlyTvLDyA793R6P60PRO
c7PSs2DWq/XBfM0O4wy5Q+BFAd1uar9+a1IgSPGB6sn1sHs0AQNvbaTWKYOZU8Yr
CTEr7968rNb5nWiTK5fjmoxVQ9cp7uOfP8NeI0uWK5jE5qe/bQFiS/5qHKKDGj1P
atZQFy6dVY3yG7I52BeocQVcqaqDG5Cu8b5F91AG46nxKwnH4pDWz8EEmAueHBwR
q9wM+2okcSFED3as7O8GMTmLkKTvNR2WVMcuTcq9jEleyUBYS3tDAzy5agD/53Kf
Ggsj3p42BuyJ3/NH3cdLCy5vbKWV4mND02sTInQMeQGzg+oc1/I1pTS79lW3nune
Fwv+OAGDYfdGvgaVz3qNa//nn12zn1gNN2JmNlxoaF3gVFCnRgN0ZIZ4WZ80/YIu
rhl/DbPxK8v8LJ4zSNffBcBPzkH3Ks6yYOpTXQlvKjcilN1KU9kkXbnIbma/txOy
6+Ea12kapu/UtArqMhxNJeJUYoqRykTADfbp+B9ex8eifKFTr10v/rBM3UuOv4cx
8ZxsUOjtbjmq25jDS0GcP2vgZD+Ck861nvYaIJpK3tzQY/muJ0Gw8PaDbgJkJCV2
a1wRuG4Q3qtBfiikJgHhi+pGQMYNIFLfBp7dvC0L0/W8B4vsazcpnZhJV3xpY96+
xdHVaFIRljSEvCYqxj36buEikKlAqEFYJgjwJFl5u0tDqiqvLSYHAnsxrAFaZcrA
sB0XyGp/tBwI/+irI85zbqdMsnxEXi/7Gjc4koq44sfHk3+4Vh4MFacEYWXvGTnN
ANi/TL9Ht3eNMcgb3yn9pddzMK0BgV6KwcWYGD62CZZWIc7e47nUHRTb0XXkeAPX
6Hxpki5jE4ZlGbd0SeHgEdgLOUPbJ9XR/sdn9uFDfk57zjhLJOR0fCQtVc2jkMh4
P1aSvUDhJXHxs3fQ2sT7+k0/kjm6SR/WsBqz2ZZ10wCs4dITRdEZIPAZmAVu/V+4
TqunqxN2bXZU6zHRUtUJQQsEB407Sfk651Co6HcT3N7b7AZQqHVhohb53BKMnLoC
0cZgzEuA7pt6pHlODw0VojpfZuUXEDtXygDbvPFdxpsWnEYKMwf7WHgTeWHYeIsf
tzqEi2A3I4bDOI+gRMWA5en0N4HSF5AvAfgUGnF4fD/jCOxWZNvEkmHT82H9yru5
VbWIBVtaRmNPZ7DIUjNkluhAiG8Rd2XjiyozEMHTINp5CdgcHWgjlHiW+tr3pGE9
uE7Wn9Qo/9fUWhvK9pYFd4uVgdh1Xd0nshF3kFmXSli9tiQXnzX+oIW4jcZpiMft
lxKWggYUEzdDZO8lH9xKUOQnPE5O0iwRVC8Cj/9KKPW4XJ+JBVo1bD8Wuc9VjS9K
VoGjgzg/PsGF+ft1JkyT/ZP0w0CtxZCfX06PPSt9e/E2a+SF3x5T04A4KCPx79L/
86wTSZEjK+Sq+FiiyzksXTFIFlsEyzb2vI2XwQ65gX9SS6IVJQOmIkIHlvvVokAC
j32nl/YHo9BgEkpR9itza8p/pG4rBCaN5tnm8JBxtDyMDy5E02fKGFeUfWuWU4ah
u98/0mcXm8JpYBqiMVo0Cxnz8gD8lVlnT9CSJmStEp0Cbil/uov/rrETQx9TJMcu
8NiNs6OlQIa+cuYQjxhRVMOmxgq/s+7dO1CAuWBMieY/mtTkjR9rq6WehjomcX6g
f4BeUsUhTmvNIsZBJ2O+JbZ/yWXLrh4Z+th6IXlOyjXcgOYOyOGoiVqLYQQGpQgI
vCMTh+Dj2SPCCmyCaF5oMBmitp5P6GdqeZOzlwH+CCrFCm0CFx+eQ+H1Ut6AkeRN
saWEtNSv73SI5F+Aai8MZeRjfT65ki21BHifocDUo019f7QcWxRNKQfAIMx/dwG0
19VyKRSEYtbt4JYOLq9l8TIY6zesdUt2/hBFXfrqdEdN1yqyfY1j4lzsjrXC9gq2
1R0D+W/0ednRW6Mz382bQPIyERwFg01vCS16wDHCaQqVYnA75R/fhKtXIaFpLGsH
1nrK0CgzFtVtkYZLJ1fOOkRg4oE2zxuq5UWWqmLr8D1wxOJWMHyK/QqethPWNkSO
b36x5Za1PIqvZWWaEgrnfjvjlghk/t+TmCvW8FtHQD9soYbdHvW0qE2bEeCoXcXg
g4YeG7L/ZXL0V8xhOR5KpZZ+JWrqzNIaCejKrq9ICJjuoc3IF2AYAYnhIBGXi+kf
PXgQ1alWcoryYiwpnZbuWOIUGlRNEANOIFzSM2lKYsTiik9u5nHzNguYLN25hS9q
ksAJIpmomrvmyFRn56y8ogf8bAaOEFVwZUXxwdWhc4S4AuQB5qPXqh3VTr9vuBoa
CnArE8xUwhTquhz056KZkOL2VRuoH4FuLpLzFwH6HsYRwTWvhth86tYOrTIxRGo5
imHi8CnpJPONqDcd51XpszuZcWu3BqJSIkyS8getHg3ey4IRGBQCAICX3We4nQk/
AGn2LoKjFKnWMyoKl5bo5RZ0V1ZabdJ3RW8YSvSLtRWHvPMaDlLerTJW2zQM6H2X
vCwmlTyXFAShdG/z+sC37DbVcwF37EZwf86KTOYTAP3yB+jcMbAazz/IPwAdnsFp
vJpKU62empCo/zAaR/fEpRX/Km//baKe10Zh8V3y4k1cid7g/LhTC/7aYbmEcZ5g
hKgjUtgfJomxqhgUQSS8B6G1tbupSzMqbFBMvRdRKZOQGgCHcyaGilniooBkvOQ9
`pragma protect end_protected
