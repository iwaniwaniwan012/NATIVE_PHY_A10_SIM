// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 01:23:56 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WZwCjVoIuupmltL2B3z4Hjshv7FCkiGh+58roNtjZydqjAFdfqgmLh5cq+/5fYV2
c+25bugctqkVLP5+bMKEBiGN8dn2q1Pep2sIpVIrTTXpjVJ1OuSvLGz3GYqSvVKC
URakI2iJakhSpjAg5FjPhQ7gzSaBzwjgAsp3IRbiTNs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5664)
uE6WbxefpRbDmS8IgQXEW3bKdrJmZUN+1Bzl4yblTdQ7zgf+h+pko7RHWiGcwYyz
dMLB3PPnX9NgTRQ1JosFoT+bqFd2rPRhyiwLL/rnQSrvnXcUApQ5KIAdqZADOJ29
sD9N3WaJ8C/QZnjfgzKx4/5jnkZ3ovptiVwOQlSTuEMyeRTj3JDJR+hvqbq3PWY3
VlaKondTTI3hCpDU/fLR0qqqAPfbN928QKI6r2XIpdoHUhLAJcekLfhhNma6EpQ7
1kkEM+8nW0uz1/tSu78mEIkwZWmjZXJH7upVr5fo7W45kyopauOl2g+g+HirvKKx
xZSXYoIpUYxhMTG5fQZmprEHcJkl2GB/6MI+vNYdSYpLeyvQOjHdFad0zJqNXxWq
DcHGFX5t7sYzSx25hRfsNmzz0nNm4RpOcdlN9MtUx/Pg1bmfcncXjC4PQXQgjs4y
P7cf0b+821Mzhb78TMB7F4cZ0P+alEvkMCsWTiiBBFWvOIqKTiecY8YbA+nQtgbe
/dqlUZqmOQTRK8wQZW7ONS6miATnNNPzDT+qHPyQnG0ekDCD2lckvoV/37zOMMZ0
AnKj6zFtk8kfblVXnOnZ9Nnux3bfrn3EYCTlLLUQ1v3S91p5QmJtbPN3ISyJ2CQ9
P8WXrHOShVEKMCNQwhWdpwzSLNeV5YPCMZ1Hwot+GBHrjcPkTdrhOistY4dRPmvW
nFR0wLiB3SMHGl33VZahx0XCSMgSFqY/Yxfx2VWsD0v0HRBgmL6z1Fr92x6yC7GY
oyE4V2nVT5TbrDfvsKKywaTkLU2X2xEc26qn3nPk74nhGSpD7/CkLXjabnIUjNb7
YDd9gzcyild0mvgbZsUKuW0T6YVXhFXByLgMvzYg6Uwvb+V5wtkYwS8oUyd9sxR/
B2YFR9lb9P2njshqIimmyZ3DgaSBiJTTlBIEI6Ej4RnHgfIQOsm6lTEREZiF4Yde
gxAxhibl7ZGFHi9UvNUI/D4DctL+pkdVJ2m00OBfpO9zU/svZaEleLeXTYHB3pz0
ZyGVwUBEy2KWhNHB96IQvTjZfS3hcc34AQ4Vgg8CYbUl7EK/hjQ3RNNbBZ957fPf
WfztpKPgaFSgsr2AA2qPM1r2Mk6FLgWf9mYp6xzVLVPIeNbN3k0BfvRzjt7lq175
H9SCJkCUg8OtLPb9HrzxZOAHjqr/7zA7DgJh50e7PAwjAhs+DfnGsWbZOe/9WElZ
mmoL0dwjr1EPsqBkTxdJjgi/f+LLNPwKocUZ+xcPrl4TaLXcW/QOHeXffXHbsHkr
RyE8bQxC570/z0TH84K4i8lbajQgPBqCq1ZSlbfTIflyOji3lwDwxSHJtIQfr9cu
NinAX3G7O0/PjHfadQox1PmFeAVfhZNp2vwEUh+2ZlNfdofzhGk6DZ7T6MjVICLZ
meaKW2OxXUagCuiDF0xZTUSbLJ5044DFD1n6hJIlbeaYvPl7L0vSuHDmFxXDqVAY
ln1Em/Mf48dMZ/9z9wjjUhySig6HmQxId0m4VsgQJx+EIWMjTK/PhnyCreVleCNg
9Omio/OzPo/IdP8cUGWVdmpvScB0K2QuYwl/abNEm7mkNRcDwnEyMZJxcFboKPfV
a5V7T1JMgy8Jj2nRcInkxHASQoDDosXTnh/JNj2MhyjoVatMnXE5Z2cGzFiocCpb
BVFu1My8vubpwLswguKTuztORbzcNk3twJYZ77TNaF3eDQ7bRaYLvdISezHE+/ux
3A2JvE/NGf3LKvbhOZ0i7skmgenNenQenBcv8CU6aox6v1IGS/PKVf3qA0gvO5yT
SYY6dGRltITvZi/va9V4On/Hej1IHNKVI6AsyZYhMG+HO4Dm+/7yJBivl0SAfOvO
780mMevwM26rDRv7J2qPaWDt+xRufuoG+FRXuN2xYNq0FB3B60jJxASV/P3c4s/2
8V2sgr59QVxvitbRna/ZOPcBkHtQvfR0208f2OTAL/LOq6LRYNCdPkPF8BDexeKZ
kpl7udch8HEdr+dcNGQ7A9cXo/SGF1bE+rJ3y1KmrqbrX5CAKOMPObB6su6NCHLw
vuHgXnDOQwknFnCmkp/oApj9yeIi176MHS1hoDSFCgp2hQqOPLwUrtSgfzlxV5Gz
C31wLB4nXMBVcjONFjhmobIG0InN0JbECvu9G9OKAd3YaJmX8NmtCjGEWW1h7vM+
+wfmd6PZo+bUEoQJe7JTXomYWBSdpS89ft0y4/kCmfa4PzFd6yjeQ1P4wor1m9cs
fyGrjahMdi2IS1l7XM4m48Eifk92+oL8jcTxeteJFvMYG9iTviZlCNRsuepGiu/z
+HLuZbsCS7WhCNVLn/wOs/IwPHjTAgKCnzDqZvJJtiwN6n56G55yeASX2SlAlc5u
tX+ePybPJdE1OJt6oQVW6yfU5rL4CgS5Yd58dTqy087vpmO/GCIT7KGj8xnpfwQw
SSKXeNMNFYHYslb37ELgcA9dshD4TjHH/9tC20zdLH9Sy57o3BOCxrMcfT4VkHiX
mPmW9s9a9ly646FhT/u7J9Xy0d0PpZ9cIkoyYQIrLDDwN3l44YqGJLgoydwq0kOX
stS9purSwTeE6z4aAAQicT6WNkoM2w6Z+iIbeGxUWHqJ7ZTOfDE1JOptJHUXQwXv
HMGiVEXWrieE5mJaAU/L1aawAtl4kCOH4D97GKavhsgOxZDEsQ17NTp2ukWQ3LGU
itO0IqHIy8hdLv2BP19mi+EZ4pxcR8BKD4OX+9beIzBf6wyE2HKUJmS8gY/XFuXB
9fdA5/IUWzU4s0insAEH4DYfYxyEl4ZykYahJM47vyhD7WB/4gzVtT4Rigvk3r92
cU69dP7uBcCS5Xy8WAXqLKAEKA9LsJy31+VLBaK5Y2L4czsFOUag+5hJQYae2DH5
sqX8C61QVoPjpzQ4xOD3wfXkrWlncUOP9ntKdJNIFzUYlgzUmsDjeWu/N6/58wDa
OtXoSyhUG3eHUY4J0R3dPn1MmeVDAJsJt6eUbn1DIYy4MNz8y8gZnL7fG3/6d2OO
s2j73TGAymzBq6ED3ig4gGeELt7DAASCRKRVg+2KWEph0+ADF55Z1ZRHZ28dnKN3
QLDBLpRF3FVu8/vnqx2xfqtMUxkXWpJOLy9hJMTwzzDpu15vqcqLGzIRWtknrRLl
EgfiuEmDxJ8WqdEq9oAGAZI7RbrQKBHfRMHBqDSjpySQ9qSdUFwxgMeg5toMWuiC
0pxRnhFHZeuNhu7hTVJdmH3Y5/1RWMLO1XhfP9pSbKwLDvgKca11kEhekplVMkRr
SwWgFNRDphMvAaaoX9GEscSvDZHzRsKa6YsCfM22E2kFgSq8jrcQY9GkcQeTQZVy
BEsXH4rPK4csMytdyc/bxr9ltMOYYyn+huBxio2RDpHaY5I6+jBCklFvemZb8E4a
g0Ulv8x6ZQeqs7aE/VobWSlW8WUtI6QYHeGkQHrfSXtD//9sh3+DLy7C4OuTn2Cx
fafgPUADkDJUfRJmwvsAhqy3TtEgIDXOFUf/WrtW5KMLa3U5/DFuTpiwERRAizgS
9WfB4z+QSW5+Nkto5T/nrX3jt7cNFY79/cYu7oBGmMQ4oYFMMq2hpaFFebcVuAC4
5RUwEeRrUtT7zvLBv9+6kG6qox0L/I8GHbPVqMyxwPm0QimDFDkYsPgPTN7DtMGM
6Pz7OaNl9nLnn158YWKerOLMwGnaloQcqjGPUJXjzAdaoyybaaP/mnsBIr+ldGi6
/0noSxsf3zjAAzoiEd5+AREOhTYbGfVRJAAOCS1gk70oiShFbhwwQV7gnuuoSwUm
7De3gSz/jyen+sojlNO+LLtJjF7eC7aF6bqztatITXzmVBYfaKg8c2NRzCNQiC/P
GKJvuw0bSZtLFGU1JA2BaJ0eJgKq7y0qI/eCDMHuhHuOGvtkgpnIlN1PxwctOFeI
p83Srv3g/rh+KVvG1JR14wYEqciot/uF4h9y6XIxvNsmBbMOjaZpvLfwB9fSal0k
MXeWT03TJX9EwVUDgiQp3aPjgMiSskXdurtsRajVmq85tg9MAJgUD5dm+dWSzc8f
dndxoEmXWDXXNh1pIn5+YQoeX+E2RWYv+ZUhrogi9H57gNzQ1DUowEnMEfBEyBi0
hhgbpmzbV/RzSWO6AR+bRYpuqpTy6liZHVjBZDzBRh8W/TMGWrP9rv0lHx4vJuGh
P6TimKAu/r+iC6zmqONxdTkRrGhXdqEiddpluewShKeF3SMQp7WzCqYwhht3Xi2j
pUtIXhIjUm8TkzQ2ple2tDP5O0P4ShQFlA10QPxEVWKS3kc/DpDn+mdZTFm3gjED
sobIQOLf2FhQeofh/qjnBlEOr/LIzK2/MHuiZcGYa2i2yPhsyQf86pHCjtYEUMuC
TgM4LigkWfNVLNnsgxssDxRQxIDxg5QtnBZEC065uY2mKyuWE57lkQrW2k7zIPjb
JjOj8g/GOMBSNl1emRVzcT2RQ39rfAT7HsN3+8N5jIsbFyOUnhAjzVlDtyQr60BA
hRhGKkNftKXXPN4ajFb8Jopg7EHPr8Sh9CfaavjCSBVdQ1nXhyEjVTh2qkovv47f
U7YB0ch5jenbRcM90t+ep9cTBAb79YZ0CvM0EXu+lLferNrOeioTbWa0uDhJcyjp
xI4kaMx0KiFNwQfFMdZmMQUzAqj/uKz1Ttoh1WpUdJHWUYfAPPlGJRDL6rSUwy6D
CKwEOfBGWK/XkIrovoW3gtgtiDrgUjL1MfeZLKM5veuPDF+nvS8YU98dkw835A0V
VTnIACcR9tHzWRb1rAkwUbVsvfP6qNGzmS4k1U1/qcEeJfAoS97i6kyksbxTr7j8
/XFSTgAMg1ulduRqhrT2hCJw6jd/s3s9ehHRZW5KVqsHAB6uo+r7QOOLnzRvtheo
0wRaFWub5RIJbZbkO7p1GR7aRDgLdtQ8MMMXgfHstWWB95vSw8XPfHUA1ztCo0T1
rugILhPm/XkW+YHG15/7+qH6Ji2x/SgnoRdbu8NGs23lQlEdlmb6OaWf85RtlFSK
+p5IGGA7ljWf+KqRxARhTV9qlwHjBiCRxkqgsR4pr3kN8Kn72e9gG4//HcAVVRc+
1zFhFHBTQ2JRJgGup9J0peDf0yS1Zmli+3qgDpB8woR3tA3/c9UHMpYVL5VRVg+E
u6NPzXATPZSzrMiYz+SEvbdbE6XhoxWxLKB6VW4Y2RNxCJHxFui5wIKVXpizpFgD
m27AN0CcVT+YEC/sqM2/f9rQGOTUKkI8xhhE8cIj1NMEZnmMNvepWrNX0s9bNlAK
XUG3SXaQX8dIdUdjKIu/SeDG/ibpcV/sGq/4BUAlECePmu8CicE2ztMoOoTrktTC
j813Rz2OJSTCadijsLmtmio8pRJeTTHCEcLgVf7AdMyjF3HDqQrlttXKaSPbwPJa
mAMipSTJG8V/7tWSFv736SMWtyd4bkEKQ4L2m3oFho5g0FAzkmgwNMgOj0umBpfm
9MCop9J/p6DTzPNeBQl6czNaZMHwz+I4joJAhRGX7StE7QWGE36dWsU0lqbdC0yY
XHeV4+QXgO/tPEhPBXuC348I5iMEphITRFtbYvRfntqGdN5NgW27ewtxLUCAVgjo
MXA08OnrxJG5/vjsPLCUGrJ+8ZS+Rpj7nwigzbXlsxUOt4fZu1sTRX58KQy8lzvo
taeGdZOKnUTaHfkIYf7QLu9a67UKOyppWVrAkqiHA2WB8aHmn3gm7hAI5LuZvPHJ
Ybzkm/TslCCsZAztquuC3NIjX5CQhXQMYjzGLjW/YdcuKAkUdn1pm/fFgh1/yWyJ
DcYv2GZo2urdlJ4wNTsRWUQE624JtMu3XH4I3c9o3CGLSNyZgLWY70n/deucuTSH
1sNsI9kDdhCdpI5wYPsq39Jzx+a8yc1rpS9rYtpGDwSPHsf4AehqzIAMWSKrFD8z
IjE2WKIoU42GGHcwi40JQ6ZkT36ZXaxjOZkKqcDqrlS9B6CdI8M74szkhIX37Bba
zmPikZeLobdRXL6DjjVth/bv41VsLgVZL4CJ3H3Wagj3d3GAFol/OrcpmsQLtYSo
et6mo0etzQfcBuzI5Y7N0KMdmgALotip5WA01ePjpRZfZ2n3GDW5D1nmtweIYrQB
njq5F/e4biJnpAZ4FGAg4uU48mAma73hya9xwez30nnutO1z1fBS09x+KFDHgqaj
it3ps++zwlCCy5qYxxy5HSX1FUBHeZFI17Aa6RuCNbbwhGhXZEG7WShddRHk5Z86
kq5oC8RUfmERUcUYitRNp5lIiJOFDjuZqL7/7xn3S23WDHfO514H068JHm5lVUmf
9ZKGzX+u6akxbWsS064AHjEPedWoWozhGJobFl+Nway2uot6Er3sWPTaFTp48fA2
Io4XxbmQ5x5tcTVs0OH23Ye4aslwu5Lbagy2MIiBIeR7wRgPHhpsf6Hvgk9oRnKp
Qp+J5uEvwmOxLtYA+so1Eg/xDuMcumqRLBeY3GtoL7YQGK7knSSqoUReYx1jN/qS
s4A6jKNA91RtQVpWEpS0pi9jLnyRLhiaRdXE/5/ZjoNOxo37w+ZKkUs+cBW14LqR
WOxxpUflTIFP+rlzuxdBrntKSRJWDSxro07q3O8N+0ex3e6wNgPPjD9qQrhiKHQD
l/YjZsVXttfz8BhayLaGLj1qGh3aE3HIs4ekQxG/vcBV9nHLE5v2lH6GBFFzACI7
BkeijVv3gbR/BpREGECUvHKB/OwF9szK7QlQKgPJiCJ0hcF5H5XoUAkDNHYZfXJ5
YzgnMiNfcNjutGHiW6srPlTJ87l7YXl4qmui7ajedgPzKT0GvthMAc9oktL97jMk
Dh2hcNd8tW6NXSci0RbSSqbI1tNUDqjxdKJUbEEikEMZMyeLhr31rZfOayUXiewF
UH7peV+SfN29SfO4kU4vsEjM2/LchXzYWMmhU3i+QRr1yl93NmDSktY8JMNF5PGg
60UMjLdLYiOn3f1HZA7ZiuVww7i8uSlXeb1ODpaBjR58XDf5V6DzsUtEuZHikbg+
1RDJQ6Uv+Tee8+9b1ACkoxw5Lz/ft6JKJ/DVvGYSIucfMI/h2IhAtdcaWLjlwukc
Ad6WsechzbIFcWpp2sqDgqyZX/F2CW9vzlRWK1FprLFcAgWqWWb3oR82xnKLou7F
Qsvu8m7MLjVegEH6O520luBCHeQAPFjjZd+RW7XcqedII4DWcM68sy3cNNSiDLXa
mN2U6kky3FojI4r/XwMsSqEFqO/8NCAH+rmr+8P+1oSpFjE6a83cfkJKFEYCHfBf
9gcJpvFfBz2mlE1DJzNRg8oo2kyp7jMDlwGDyczam/O9CAcZt/zOMn5TMzxwHl16
GYQN1/9WukamYloQ1XL+tnukPTu3zkiS6cPtcYr5gobmxwDvvf1yowrwp63PZH2N
baR2tHUcJre5NcwVRsmpX9D9ceYZ3XZpVjeDWLY3A1svRr6JB/JLOPWHjrvWKq7j
Lt0IWjCPcSa5UPz1UpowVbvtVUTRDbCtAkr3ACT+XUTkHYFi2i4quPO5up8xDStx
e/Y6QJJdlrCK13Sob/eOujGd/YkmRo8kEICZXZSgyQVz61nCuHDO76vooCRwX/K0
`pragma protect end_protected
