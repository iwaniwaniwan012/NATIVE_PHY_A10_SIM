// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 01:23:56 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fuG3zyA0DC+d+DIHecz/V93e8JRQWcRhuauE/J+Jy/KawT04patefoJQtTuPJFB3
nBjTXQFcl1RkmaDDdv/DyLVccxAI7wRV/rKZ11pvvm5cdjYA/0iS8w6z4w2336BS
OcKtE77EPGRatqla8G0wIZXJAM4Xk2gRLpF9W730Xm4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6208)
Fde89w/xaqKBZv0pv7QKzhlRdFoC7USZYRFhb4ZfvwFiaG+Sg7gWaK3uyj3L1tV+
qlqoucAqaBwEcyzq4SSigHp4D3t5AOIH0XFMOgV462TTzAyCrw4OAOeYk3ZNglCT
ypefV3GOXKvMgWcuqdNRw4sHlN4TGioxPNTQrXQuqo53XXRjWyTT9YXL2ul1I26O
1Eb3Vd/BTWyRAu60HuKOli24MnX9ffw0YHQbzlVvMMzHPTUDD3kdLrjvPA86+s2o
Ekq5H9QpiOe31sOsmm8DN8BU5b8P23qLDw0TUi70xECAYWRf+6jXqRFVt8R621aO
ajr95OF8sEn867cyhhUMcyKnoIaIwecuVm9MhRpzJdkPOk+iyr5oAeDBuWG9ryfU
zWSQqcFn5AsJOMd7sg3FUThndHQkbn+xk8i0w03/xo9iGUlwm+v5+HRrnvLqTLG1
/amy5bJa3TGspUsIa2CEcTeKqT93u+joWJJohSU5yeLGUZRN8vm9DMh1DNdFrLbv
UViweU2YHGexr6iFGkw3kmOqnfZht9U0Dfkrt/1RCoDh1xE/Nb8KlO8C17UJ6uMJ
VMoDVbfqHnvHAGUYQayra5j2dQFt2Dl8N3KPVjk5UDZwyxBKmvewXzEC6ajpvOtl
MafMKLyg7iF1nhOC54pTkif3JK6orgxsbSykhB9y0SRyAGpwPCiD+8w4VirBMKNM
LlhUN3bVRubZqTgAVVRVqroUbKLSMz/EHPq+tJEJJPlZwAC85ju0AUg9E5Yq2DUV
H4sqOVygwCqNP9C7nfaGHmLeNbYhnst94MNHWKdayD9jbzfn+4poI5ur3+gRYFBZ
Y+JpsgZAY/CQBevvBLwSU/A5YdYFp+hc82Rdb6HDjLXbkr6h3CFAV/DTlmQmr9Ka
rJbU0oPZy9M5xv7JwtluISo24LBxqRAkcXvVNG/TXXLKjZe9QG//kImuYxS+n5kT
WytLkd8OhWwPhV15MTnMqr1KskY4rNlSKTOC2LuGZaCTyGThTmRO8VGu/SRMPkC5
hK9KmmGNVYlGwY/8Y39vDbWFSUtkZoqhNxnWWjfmf1IJ5bosrHJl6Wm+/rGaTRfg
epgZBAL8QWw2tHuRaV2WacM7wxx03HRK17MS7Tp5dISUuYyJPhOZt0L+G37g7ao9
1lcs5Dyw1+VdY4I6724nYKmj69Ol+pPF5NMUPecWtPNjIYp6lYfEf2kUgKXZmlG/
sl5/ipmGpVU31Rl7vN1T9gSMkunCYy4SM16LX2V9RUCIN9BwF/8djYIrH0bWNj22
67DVWdl2bbmb9IsdmasFv1gaZPiZhsbYsxVxKmPQLHHMvah0P8ntLx8TCplTO6wG
DKqAn2Ig1TvKmx8h0nsPvvMA21/N/+UBDiWkHezvSCv2yMuN/cvZHz+jvp3AJduJ
asGWMQbLEKMshSq/vzPs38Snn2PrdKyvN9/ubUz4C9fa4+7v94rNyrcn88ucQaC3
wSX4q9JCGLzv98C7WFOsSgVNvvqxSLHLzUrJSn2vKycciXMGi84FgMGXSsqHsU2E
0IjrwL4061umf+VCk+MflJHY9xQYLkH126SEPxHuyYzPloLcP5jGkEcjpVjFw/Fj
TviTtGdtZ30OIO7kSkXIwVP0OD6dmIOlhFat/QGtV8t3U7WzuJUc8ks8/YYn2tKa
vtoPezTTmrJWzqg73K4TxELwFRgu/OSX9s1KTS55rxiJtQZITca7yy0AP+7rjN9+
vVZHNsCT+OujtPbaPvcLALKUCeIrGbhy4f4XgjBNIQmgBcctIHNLksH6FUZhvk8R
CLpJSV6ogrKamiP+zlLolpiAjGqWToDfrcxP8ZrxzB5rNsPDtwewdo8fSsVAIjrK
RItpMdgrhGavKnOr+NXMIk02NHkvdi2KOYjq4vHV/zpf5t9yByeBrckmQiolHyiZ
+Ti1NvJM3LlwTPhkh+Aovq4X2a3L/JJ5PR1lMg7oTtv6HgbwGjDNiO+rcdzrDtpn
S0jQJfI9421wnNoKd4jlOKXcydimFbWHp8vaeDiFgn9kergedvdDYhW/1XPoEVQj
gmu9Wk+eORjSQWH3ytt+PIGqXgIwGuxPKMtTq5cJKu69k717Upld24gArnUCLpau
8abnUjAvaFFcp7ahA4klsAWq8Fco0VCMZ/gulFieMLq65UwAoQFygyucXwztj8qh
kAbyCacW0zpqLp04YMRK+nnLUXEDE71BSx9CdegEuaMbqKD8Tdi2oy0PorKvOkuo
XewnnyqmcJudGsCOm2jbPy/L6wFYL0/m2UqY7x46haCEUIEKKkhRa+OeF2sjCppj
dOyiIZs1xK8aaLs0mm8DsRMP4bKVzmJ0RHiz3jYILTrdu1BvRajL/BKdq4Bc9O3/
AZEdHpjJNCPtF00rJOC+3cIw3x1Hre/uYSgH/zqV9frigXOfUBeq3EQJfr3UXTUe
WdceOe2NuE2mQcFy66iuYyax3EM/UfVZImkK8XbjKdRKWjl8lHCLbl0vjfXVowyC
xclad59XRuQMtOZi3LCeHuNOMk4TGq8XMjYeCxi4FYboTIV7bjDzOHF43u+x4gYe
R072Rcs6HrbJhlVQlpOg2jQZCZJluA5Kf8oBDpDwnUgEwFMgtr1FEnRd5Xs0P3cB
zMhIHNGNb8xE/IjKJrnirodkyTv4DkN/R025ZF1YadqPaV1aJQlL1L5v6dGCyhmT
bZRmZRTPTu+wuSIFLqmQn0IRclI6kN0vMyX3eLQPvbQyKXu3DfD8nghZAATr63O2
pbmK5akol1ztbS+af7BAsT5vrGrObJjhQJn7Nv0q2hwoubg5EqddC9jPvOREw/wz
spxDAQGS8Nzx+Yo/srzaTeTuzDeiPOOsW+n9UiWZYFGTz8a5Rjr4EJyAYzdKKenR
JQNlkduG7VK19WHXKsNv7qWSgctubodxgX8MV3u2GajYkF2vuD1pmzm68VGPfoqM
BdnOX6U84sD77G31pnYNQz3jcXeb4AM6Ktg+Mm6ziZ7uDkcJR6v0NP+VV3TWMted
cTAtLffmZKfGactvO5lq3MA+TdFAvmITDTq7KoQZKfzyZMn/EgAZ6RGAeGzNnpwt
MxtwJCuSNut0c3VFxhLvDyecpWnudSEQzjtC60U0tNCJ6+JtI/5rdHOGZmRHzTsP
B7bVPv/VQ7FKnCUQmVuuT7iU6vbDt6whYt/lQTN4ds4m8zw3tMlmeuoNg4TgPMTd
JNCnKwFRpIIc1czCpGOkjNcW2D1RvezynXOLuWnYVf+d1hUOP6uobRj5LPUpLC35
Fp2E1GqIB0cr3MbXbPq1/Eee8gE7IhHY9g8TBAArb2+m+j/NgmH6nmDufLKKGuQd
WEiMKF3enjihDDqOBwWrJGubLw/TqkQN8O6x6phfssMsNBATjMndO7CIvo81Pojv
iuAJ9zosW3qwoB9wyuX1cWAbp6WWl0RL4sINOzMSWFfaSIY8U728Zz50F5qEfmvl
+scIp7YMF2x5bth2IUsOQmXYoLDmOqZpSG2e4G43NW2tODdRlc3+Fc2QgpMoHhyo
Ls/W75inNA0jP1OirbQ9dqNwprjyv+gSJYaMCYiToPzofTq1llAy33E6ggPbG/hI
DNJa3ufhN6e/RxT4Lg56A7moYjGzDT6CH2zo1RsB5hTBx/2ETgI25uDeJmIz9QE4
UyY/mEU0h+pj8dlTbo3fdChZriLgR4uPcOFXHBmZN56dGCbriwD5f8vKgojoX4WL
ErOdRfjPEefXAeArTwB088LWOpJ7HVt1hkjvBI4YkMHUdeuPJuB/9c88Q+ASRYe6
lcJTlLjU6sBsp+/FpV4OJc5xUIh9eOPAMCdml373etpHD1euTs4/LEyVa2p0pVuJ
CMjNXQFGf+css2sSR6p79VqQNJ+fjMuaFcH4Z4JI6fSUbqv1RlNJxK6ls/j4LYDu
THfkvH2pEL8sY3ENaoJvJ7JgMCqdov74bIumMgagRAsSNevQRfqhgQN7K1jaDiWY
wNAZvAQt6PwWlkkhFE/zBWmR9CRGe3LPU5vn/43qyVhvS3qQuVhTGB4p4BZXyyG3
9jNSj8/tTObhIqdRusqFVXOMibaHrzU/ziTkvwcfR7cuwREiuMCpth3ydyP3JOmB
Zuw0eONUhXQerKVDqDVKN+zZT+GKUpk19xPSd0QjLuJ3mU7FNnkTTy+V8PWAVHMk
PvwXDrNu1ELq95g/kI9qnXKD4RpqvdbUbDx+by8FWHr/hib7ArD3T7E5B1wb86SC
KzBbUCbRHqDtqjMldtCzJXRpcCMrksy9fTa5okIbsRuAqbY7xD2x/FDyC21GY35d
m2yKtr7ByhH9fBkbmiIWvh7zcUZq/e4EPQUE9vBzlxXkiTnAGxYvI4jM6kxXEEpA
IH8eJFDzbLwCcSupxtGUsD3waDOWS7ivFwSlSzPWn35fsTvZsIBzyw2360kXkjhT
2CbK6uLLAttyOpyfQIiYHMTZtLQO0dLKfKqkRvOk1ISFLwDJKti7TUuKQRDg35i5
aOu0r4avT7efu+oAyxAyP7RPaGenslNHDAssbHogkzTUXrD1xQ16aASkxi8c57sW
bnkP8DOqFjQ0b2P8KKIJziR+psO+7P2HR3bv3yamcyz/RjWrq6+ohCXjQC0nau1M
HVhQjx12sL1XyaKuWF9SesSv0gf0+8mcI895NTAE4K4vZvaUdpDNCKWQ281pFoe4
3fVMEguzS1Vwt7dKHv4mzBtOZVyr8wqscYjJUVu7sXKJt+3J+vXf/9xG4AdOtu0r
4JbeoJ2RDMu2v4/zxGclkGYRVIkhKCF0qJNtpfv2drKOOpOw2yw307gHAkr/+ZGC
x+MYX46wetDIPV6zpMQXCAa/46wMSqKvUlIlN7EiEF/62WASjxkWcyEQ5iVIJwq2
K7z4aq3NS77mVGj1a6bbpvv/6jpJFaEHaBL3PhBfN1MeFQzU2RJhWwi2QlH5Bigb
E3xD+wuAJS1H4BPN/piX0jIVMIivFasWDCPVLv708c0kt+JJgeSD9d+JHbkdXRJX
K6m15Z8E4AEkeYVOJ6Tap/dfLX9biYr7Thps87YYcPmJi0rK2ux8qsuYC26Kqh44
R27Y3uZxhTCiIbu5cpUKelEQq9BKHqohjeS63uu6UBk5JCTcN3//2j6NfD4EOJg+
ccwHnL1l40/0FvoZnsWxFd7KTMqkSSJUsAwQEfDzyvi89XaPcmO2qwBNi5GacqX5
nH04KqRKftnW9NUiQPzcDIu/V2n9qf/c4vTkkEcJTERQP/SQwQz8bJkK4hiTMKD2
41nBPRvugV0rbdt08art9XRjT6FurjszSTWr4iSU8kjSxVA7URs8jEOGYDrp/wwB
AEIIMBfftK/ryBuDwVFWW4qfda5MGcvoTOY8mfqfTUhjHftNtHG5902gEBdkiSjZ
cYpf/INTxhm2cLXq3bJD6dJOIl4U6ghTVYVgq06zRiXndpOnKXUj6g+cK5AXnsx+
BuSL7zXTqk/sIMS5Pb0EL4SygWDVkwOJRpH4UKajMjdy8KmgKcTBBKrbJqchSeBx
6knLb59K3HjXwZKN6BBZ8r8014MYWCG+9RcQtOQ8rvHfCSws11N06hU/gzovgDnF
9GaEqBzs38bGgJziwMTau043WTyQr0xcQkQIddjelFhk2rIfS3boLWLsWknaQp1e
etyb2UtII00TzS5uNhtKFBn4ujE/W9gsZmklna0+6Jdx9y51nI7T3dgwcbtZu5Xr
x34HRGfVZ21K3bFvPvMS+TzvQnInUSZMzndAakvrvnxG2SrVsNs24FvwHjjcgxHP
lAQn4uzn8GYfw30qncbyJkIt8Z9Uka5bw9HsZVNCV891V6qgcC2JIrzIrBvobHb4
o4b4egSu65sMB45nJAO9n3PRotpMtnqvaTaIXJgQ7q6YT3svqLRU5Igxv4L06249
mALNR0OLCJJcZUkHpvGSGNUbCXDGBs18PE4id/Pbe3V8D4PcUMxDCUSeUL/20l5K
gWa0WwRLb1K3v+3TjuvOlMIDbNlPyPcJr39QqU+pdsNGGDbTb+SyyQWxqcoLpO7N
APYg1wLikVmTN3fm1K65B5hBp682SUE00Iwaf9K4Dt2BcaZ0FhvAFAaATfo80Pf/
cvECDBQRsdmLuXVrqpyLhSYl+GJMbL5hG8tVx50pDSTOMDXoC1vqMlcnaDvrdbHv
gAt9MzTphYLwpdZ0e/Y8rrwAUXHXz5bBW5JIiGovykJYNBQWnjHa+b+dBarLT851
rlolJqKZW6t55TpCLZ5BdRB/gTTd9+NxlGrpJ0UW72BL1U/HH+0hv2NPsDlMwjmh
SsrhWTVReL/XoIGh5/B7OI5BHCMswRpoiTCBIll7O9KwaVOpNMBy9T7pLhCdtxKF
dh7N0ouao9Cs6kbfS/8opiRfbHxr6jscehg+EJvANqv9Hy2Aq+AAIGppBqqA4NeM
qtZuR9Di9AEZwTb657lXMBaOS8ZIHgixm2CY1tI2PHmweDYKduO+7Xx7K/0fQh1m
hZYp5pCoPn/XI9kejeSIGHZ52fnPGaoKfMsqt6RzgOu8qwiXMLZPB7nk1y6cb5EQ
ruSySfM5JC8wZFyzZKYWmrKn7dVOe2iNU7wTCSdn8XDFVlvXZfpj8zJqHHN+yfgV
M0VYEVEZAzyY1vQDCNIVrHqARz57ORZ9Et1mGBO3ad54BQYnFTvEMvYgcv9VIMyZ
Mu6hf28iF11MKSwV765e4OZI8X/5rQLYd7gOxIwGeoN6b1EimOyvTG8gNJ4ONEtj
ugHyBjPUnFsakv2Jv07KaQ7aVxUziq0p/D1I23ZdOJs6AyCk5iRrvWE15Wk7ccDd
KUINMIgKa7tDVp7MtjsBkRMuoe50Xn3ne7vlFVLxWEa3e6KSYwReaoxv+0X2lhhg
zhcN1EBDTZdRZlpEfXAENnzESMLsudP6L8PvAnCftb+xE5tiopZBFG64p9sn40fF
n6wTefp63kPuS7k9N9RAe/KF4JmMGnDOrH9O12KVkii/MXF8rCluYgWtWDN2jxBP
kUXnJ4SmhXdMOZpAAssjxEtBdEvbgwRls2ZpeTza4u43Au9+bM6bZb3MseA2/7fC
mzLyBy9h0zU2oABLMXNRv0ymsRfIMpQJfLX5aSNXl1Xu9ZobFBH8+X71PFnn0Cp3
aK344r/e7F7gGVbJhO+frX9XcEJmVlrQ3yGK7UUXIysJg1J4nqtQcIMa8MM48iaq
SoP03O5QSVOObeE/yyVEa3RZlj+Mj5hscbMw13kn6b5mHKsjc6Fbn9RXQJof0tuR
YaWfW8IDzXUCCLS72w7c5vAtL9/5Y5zhiU9BDWUO/zL4cdfwjnntrwUihBO9Eoap
wkwxQVMEjWElkcf5ctpYdHNEQRDvEnVtuzAamR3jgMqeUgfE9xZ17ICNvYvznqvg
rSShRljaHn3aUUnm0ZgcYVJgF7V3ahHU8x5gNe/pybaSSzW4fRSLj0NnbMENDaI7
erCz2DUIfkz1cP+/dmiKgr5GOqj2sJfo9L8jGITQ99EtVdU0y+TYml7Im9FWQnIA
MTObBtjSJEhDZ9HBnSrD+eCfxNWqbDvyN2R6MnsdhaKvRQeM1DokEANubBhHfwd8
xh/q2ogC1gpriok14nbKCdy8/N0XQBKhrtgUNo6+eS5qBhc/lTvsdNpdhNCu0PwW
UZg6l3t9pdkHhWsTnS6HoVWvGhc6oRUiHDs1In5sYvmuz2vPerpEu8jjrHp/PF5f
xv41SOuva/lqKY+RGzJKMabLEjOrvhuIW2NY9vxOntt7lsH9ExOd3eUYdsmimc9P
MY/AAZjUo+3binZF6/6FRxdoeXFNXvu6/ljEltIGIJuVQpySCDUrWHC9UZiXMMEW
s4mYMPNR8U8j7LQwAlIFVz2h1VS2NPv4El1fNi3/92qSmwiWHeEeWb4sXbAlCoSt
jXI82Jd+DaSgM8minJLrQQGQWdj7uzeReOqj0NxJ2pN0MGZXvDUXgLYx1316jSNV
YoFIGAhjAvwSM+yhBL1FttzMkLJxr3C4KcgwtFCo23TV7LP1eCdhi3YpMIgkLaMM
jOKAsCQykA9i6zSUniJOdnRsplnyR8NKXOyIrpLVrw5rBJWc/0ARWUutujiGJFTI
yeL8Hbi2rDM+y1KQPhqORxhe/azUrZ+iWZUQ4+tgihUtifXV2QjH+B3yOcASGmin
VcVniBIuKkrZE+bCjvn3edkW8CnpLmnL+xAp3ui2ZnPLhZ1GwKpUdfGMhK0cdZWv
rMCQ11h5kyd0V/tlSFEsi/Behb9CybvQD/d4QtfuMSnYHBo7/nZ61ktufsh/B6La
sNQmlBXSLey+10srA8et5w==
`pragma protect end_protected
