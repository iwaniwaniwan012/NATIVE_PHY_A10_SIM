// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 01:23:56 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DjJEmhNwJFNswtjkQl3UIiQ/omqzev6gm18sTWojD7Buv2xW2zmKSelEPerzio16
1Ibpu+eX3EOTU3a8WCcFaBZwr+MgrQHCJhYW9a0aAF5XEstxHT0sL3UUmGGt3hnw
dCjc2VZHxxNcNQ8hKUNhTx1Pkpt9v8aggJ4T3mx9aYs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21472)
/LFi5s3OqVnDJBTw0hlxx8SXqomxReo64/sPEcTUIfzBPWHoM9UDcNayG3SsJRql
ZM43wfhk2VUnFbUjqrVvjVfDmCncam+OfQFZieUe2ERNUXTPnC2WvI8Jw7ZxpF2Z
hHyw8M4BKW6sU4CpKaQwLpoLnrMTUZX4F4NDHXyz+FK/1aUeIsNpllSHKCTawSMZ
TyE5ElSDJ+DElw0svyKaNR6Q7Hzz0vHcGAMKRUkInVqTaoDKLibLQlJBQu9U/NYH
Ll7A3ha9ksEmNjSaAGPPmKh04CmVmV2Yp3VPAHXUDzWsykfpYZb2s+nOBEI1KUp/
X7EhFGlWQvJbBSsML9JkY7GJeI2Xp0x+KEjYgKEYtJuEj37cDMdvZ2/9dR6nDwb7
V7GbEfdeEBm41i85GfASV+Wr7YnK5zteVcCtmbUAOY8L269xCeBOpDEyP/z4vVzf
62Ak0yMlnbjwHQysJnRyT/wfhXGJo5Flgv57pMs0TEG55u0KAfmMPxKjogxoZnrM
0SE/oPykaH96ysg+MyyrjDCiv8Kru0RrUXs8HN0pUgzOFldSeWgGK7gwwNA2RPQX
pFKk3PEVjVexXS6Re9u3OznvKU0IfUDBOmRwMFGgn40fL2MBFvfg5l06GDRAW4tU
yGWOkcodkep3qZ/hJFcKK+37MLWopk65hfqlo3eZgAHKEvpQkv2ZRSii0SUZhEzI
71I6TsOhONwnm611XuNKKd2EFxjC1xgyLoLSapRqWiUzJO7/RLvMsKos/q7mpgdH
7ltKEO64tza4KqlYDklwbjSEHcRDABWyLDQ69u4oauASqWA8DZHOvu0zW770tPkP
LRPzVZUMd3fKiiNgJbYVR+hwVYreeKjhblbyVTechM/df1dtWMFpullryn4crQfg
jDyPNAAOofaF8Y+DaCxSLG3L2d+x7fLXf2WDih+5Scp0bEDs6pxCpyM+y9p9sYOY
ynh397fxZaJSmJbscXPkiwB0680EDz/RVQa5E5/0g79uBIDfQK1a8Jovpmz0fOsF
6hv1ZO5B+zTaL2jYQFhsrVcZ6XVF6osfyFYX3tp/8JW7lCG1S2nq28ogEjtT0HL7
LV6Il8+4Gr9WCGqwpwJV1ceg1K57hjOpQ5RvgrNmz5k+qBlagrI5/QmAis9w1HxW
pe9ILAierrgsVT6vOJkHzspYcSAYVMuuyoPcayHBvfwPHUTBCt93/p/5o2plSzP7
DEdKY5XgeR9hmSpK4RpxurmZihUiAd8vMi678VB0T1FVx/E270MPH+4rp/yV4bti
jwrgJWX/xbaam4avLdC/tA+vqZ6RJ9gsYYL6S6B/F48prV2/umGHAl6oMf2DgzSK
kEsDtrEsI6FW0EVg1lTeR+VBDuBtzdvEBY6EtdKOMKdVvQ9KHPnGlTcGStQn9kIS
nBnX/+kysyW2ALmHREnxJYfNzGp21fDJdv2B2SWOuXu/Rp6Q01S0VhbPyA8ZNjHO
CHXgWUX5Uerxe7CZlFeYCevrnZ3DVPu8lSBqH7D/eGGHA+utlJqfQIeO5Ub9EdF+
upNRZbxTk/FcLZejs4NSgPlcyrM+3S1Oc5ImZZOkc+k6E9itjuN1J1TJu4rY4HKO
dFOUwFkkld0GJYfyf7TfTjGztT94A2GLrd0F2OPkYfVsaGj4tZE5wGhNNj0qwPoD
w0LkS+SHs4t+YEw3aHzK//imLv0gifI/ZiSQFojvZKWaYgMmFuBkNyyZ5FwtxI4j
9J7aegjQ4DUp/vGAs4V7ZHKTSIQ77OLMj9CCMscEsTtcJi6pAIUWb0DIraZrrHyJ
foe4SRg/JfS4CEaN9OP8c4atDzliBDHJO3oobDrp/59iX5u9rKI/L52j+n066KrN
vR5yOMzwXRU9gEa6ITdOd7oQ+ljLs7rEWl2iapIKrQ4yGqmR8YpdooV4Sdfl9AeH
8CFr3OJIK8icH0IzFr9uqd95wN4ch3+33KklID39ViENneEONrUsWiaiQhcf1uZt
Vy1kL8DoFJGcUiRgCSioUYJ8U+3XIuSrjKvHFYdERX0PrTj5BPDvZEh6wj4ady7Y
2vrY/wGTACurb4XwJmkLAkvUzjwghEd7DQfcoRMhPjiglXgS0PCaSPLWh0HybHYV
PKhh0xifk0NrHIQK5iStB+ln+wZG1XZAOsyNN9wzyYa3ujJoZEjgItQF+E7GoUVX
gJY4jRwWN+9Z1kKw8KN3lDsUjvdqwOwBiD1F1uJQF3l1h3U9q3P8uhbcMxStiGzd
ii0Hiu6bKxpaYJ8KkknH4hT1KwO7+Zg5n6jZH4bzmgCLdy1xhOYxs+j2n2Y0b4/M
6+IY/9jqEbfk3U0yifp+45WKA+7Oel15M0JXDT6Q24c3ppeZKxWH0LRH9tPgXTC+
tc0UuKN2kwPz/eGzEp8FCQl8EbVeAcipyX0yrjPHi4kku0ZtGsW6WqL0dXrHBYHj
KqcvFujVLalCBN4jYCm8qQe/oKdB1uyWHBNo0zRGwg78JZYeB/PApVWflORBYoGk
gqFy1uIfG35++OJ60CjOSBViefupchyK+dBSkl4Bi8ZVVQZHfnht9Ii37X/F/Rp1
MEiOnxcRsKMieAn6Cv+GQ1udw+lnUoblb14PZK+qVdLIf1O2Kfl6d3enQ0+emt94
HWxrTTDYvSURkAWH3b4CizoBqgIEgM8ZEh5bTdVzCW9PGAEpPi94QZbk5cY+btAE
BvZrIpQW5dbuzu44nRuN8g99P9kfCVFsDSGQBVWEFgEN4lSf1OC+3xoOEtTlVRqT
tvVxRJ+LUo04/VxFhzz3D8iqOjeHkY+yNIiORIAIgpbP8Q7xGFxg7BclBCVGnq1R
qELfcCrZBRSZBFvwAoA3Oow7b4lM5SmSy2Y7cmkQIHqv522RDrp1Fh/k9y9m9zzF
dDCGC5ih7cc8kr3j77zkHf88lcsLuGywZWzRz4OG61Z5ajzl0AaATILBtj6o6DrD
NNcGeDsoGfMp2GC6R9MROtNFJ7MyjzAWuqmyy0C/9pfo6dRSiLYvLUmzRPJIY47B
0y0yCZ3O8DW0xeoEjzHJfSiPf7kguwAq44sDD8cxNUvlJeNSMzKzVUfcc+zb/qQq
L3klAmEmMPGlvAvRf8F8KM9nPjxKo3zURbvC2jODfmdPbAZuyrVzaGDAm+MWrTBf
an/P6OsVY7mTP1kvn6U9dje40ZiPIyY5EsyGFsItmLUjo+20bhCPzETmI4sUpUNe
XfsHAd4KOZN8WzOJSjZjeQfgTQEnwjR7Z4JElfiaaIXN8yZ89iHXWfd1jVXdeFds
pshZymKsvnrSjZmvTY52X731CD6n/VYXXpE3Maj1TqXGTNKCTms+2JwbWxw6lSvj
E/YIkRGPvCUMGt0Ijg6F4PRGsrDW+fjJkkOv733ELkVct9IbZQISEuPUC4wKqM/M
vxeIx12YD5qS8KFMYFC1xwA5riBPrhD03k8P8ejt2V1IFlC3t0aLO3d4qmmGtBvY
3eV1OgiBJ1Hxe2O4L1QK824PbJt/XQ3nsPTdWRdjN83uJalUbkymALiFgz7hZR0S
QlgtRbY2UhGptDRecZId1rOt4Z3dg5jJeYesg/nl23IsIsoqbkzQsUBqsIC5xOd+
pd29fnOe5PbPQ6/6lcyaoI42xqxHGrZ1K184ljm1HD3v+2s5LkTirbyCq+I1KDq5
En08usZIxk1NuUq2kGJBYpUbY0IzZIJe3O362lBSw875GpL3l8h2/PGwWqHZnDga
QSQfvl4aCG+0BoPXgnWEqY8Bz4pAPPmWyuio2h1TmBHxehxUaaLrXJmAhRaPEBPI
5wAo59Z1DNuRBeTSFNzBiP0vElRUbZL85CAYEXtR8QuL8LJhvfc9ikTeMZPZ7qEp
p17fZtFnRpdY2ub0fPTKZ33LDgfGnjlkIuPZB3x+/Fy/hjZSd4AvMRPcuUC5EvKE
R+RWJzkonLpFi+ZdPruPQtTCFMVqA4k6w9nZxEWw3LhBC2ZWbdHCpQBi4QMNTZeC
VQLtA4WD5vtQVDK6qtBlZ8dJTgtiB1Rbg4WRCEpMSVwSweLWhTbuM4tHsnCCscyC
XHOaQ+gx7o0DW8o1vlWfHNEYCL4GrnMdA8lD8G3NaQItUbX4n6jfk4oNw7qCUv9O
dYOpKvao8+7Fl0UDUAqnvcQTt5dxA8bZjE1uwN4Xy6sdskpNJdT3yO4QR1uDNkA9
OHFfza4djMW7OUgFKy5ZDn0a5f72Dx/vXHrj355eYGJ5PE4gU16Bg+7SOYqHoBN3
3MF4495H89Z46fBkLlYbZ8Adslt+W8a9bsStc1kW196Z+frggOp1dcvG1SW/BrL7
xRtenMS3VkSG7meX1CJxJcrNZNsHLNr/7iDaaMwF85kKS3UMJmJKf3pDF55ay+Si
bLiK05wD8A2vGBP9ypnX7uk+/d7C4Fu8+gmg0LeyrXyOx00uwDMUvUDAhREFz1SF
8P71gRJIm+QyRRyMnsKq/yEeAPhB3obOz2pAvxKWAIku74UQzKamoroaCAVLbRTE
NzlYuslWB3S499QFYq0N/6Tki3xb302korj3BjYO9Cm4bIroOr6PjNVsz3ZZb0b6
yObrZsX0+aiG1lFbrMGQlQMTpn4uiQNRsmpP7xyc1eibdHzGIoIoG1ilkUzNkt34
E65Emj73/FrpCWTIPOj6A23xEvk1SEMmPhmHV6XvqvOgNopikgVjabn6u+RedcQU
wSpzJ+qJ7JooLF+vpFKeDPHOz2N8owIDEFnKAZGjJZ15l7uWlxtQhxJyjt/V3vsY
R0/dQr9K/Yww/j8DWDeaGwChdhgL2ZLdQp+QVN1FAIpPlnsIic36Gc3G1XD6hdEN
ScOEyLtCWN6kzuCZcH/ba2hxErmU1h33kG/QC48FJVFyAyQECfA3eN2xduQC0XrW
TiX296Id45OV9a2002lfXeZfJaXXJX5N4EfHc5Wi1fYZO2raAS4gbNM+/3oNjl35
wFASlxpxZM3/PpDBUo71sgL8Z8awqv2/8NbONCtk3mi4f00oDxA2Ct8UH4pld3wQ
pW6P9dhnL3zeo0aj8QEmIrJzgldh3PHoRBxmKZCBQhKKpc0kV1pdPeCYxBMyuNZM
04gauYwRlKW8HXJng6zvGWc0uONRAO9K16S1KqteJNZ7h8FKLZWTor3kvXs94Rak
a6DPSqdJyDJrpW2Q/RxxYCmoMrRUykzEOdLS/t9NooThgYjwKyjuNuR1A4nsJwP3
jPwLlENM4jbQt6DjE1oSCKjyUwOlDlpMGnM/ni4F3zPS/r6MRsQMLVbT5vgOmIrB
7NK9o0FtD/yPs5FNgfr11qgUVeZHypiXnZy4bq7K/GrtnBBFV87B3dfSfW0K/gtN
a+4NAXMBy3JvtT82+JAvxRrJaNl3kzW8eQbIN+spLA/MqPqJ1Y4h9ZOtmLxdxw4n
hwdRCYeAH7/bdxpHNBUydaGgsJUH9SwDve+cHXZHUNutntpZE5gtdhjpO2i4ry/o
0gLUnY+avYC250voW7Y7kzfQn4GmWLo7gFXzG4oU/8MIzfAB4V6f4iQ/o+CfKeft
NW0TqvcKtQXKiMYi8H/5651dZftrx41omJ2FtOICSr1V0F47TNJ1RkRrNdlWjW5G
Kl5MrCvS/xLDdGp/bFzovaEUBg5NQ3aRZ8cTVrKhyF8k+wpjybMZOvgyi3YjIme5
iARW0vcPKz9wm6VNKvWYiaHoqRr0rdiQvADuy8h8gE1jv/snbGYfMoHdGqmtlkef
nqv/x/U/IRItdmD5wA0IDQ4ovSCOZ07F+otYoI2INAkKBrnrvHR5nTV0i0eq5SRC
JxydekJ1Jz3H1FYymrA5FpItOXOdSGeCQh7bi+qpIIwj0QfXav2zVG+BVuC9N4rI
5mv12S/AKkXj9Eo1b0t5EYaftr67B4adubdKX7Oj+cdmj3PtAyPnnGsoR8aGqgGA
MT5lmpHtA/7MZtVzJMaWqp+NuNezj8cL0gCXXAFQYg0XT9EZjUwxc1ZflHWNT4wB
Nk7JQDgR1uRugoldKR6gAP/qvkiYWYLw3J8V/C91mDn0f7qMto3Lr0j2I9B0NdXG
KU7VNP8Ie/bQirEYjXYSe1TLqY9jW/AOYhh1l6153xWNh++/Qelt1UTnk6vvuiMJ
KsOCzBt3AuB1T1m7HYJ0xT2NnJ2harWTBen1Vd7AyykrBNzZlOjJSBHQ3qWjvSNF
NS8hOsIBPEmisrfyt+WdWLMI1gvGQQ87TnZKrEPd9KKipozOYFPMKMfkNAPoAAHl
lTfnB1vdRm1/CzkorQXrurEfID8s4DtBHCP5cDyLz8SUSx8kLArGucfuWwtHSfyp
9YE3Zb/3sOH0fxFlcpwwHZ5hv4yDIgGGamfQzXbJfVZnZQq3J94IcWd7CMsRjWYz
Af+pK6emPAbWo7lujrFoNk3OYt8fXw7gqaX/KzIRvADvgDSJjtd08oy4FG0Y1AKg
GLmZMQs2uzrplyLMe+c5K29RLtLAQiGhyoCRL2UlAtv+ZILiXXAK2kWxrtztrSrr
oYUWKsdeJYnHex9e/DuGFYJ0OJbK84Aj0GaMKwOtJjuIlLS9ZGqwZ1qpc7q/JVNp
f/z6MT9ipBWfOUzpWptUOoEkZfSS4m5QS8JL2a4pysSBwPZudO6xAA5wamcrXmr6
UnWO6aF/9baPK+0mHf/1yrYW+cWQOgeSMUHueJpiHZrO3RDPlrBPfthPo0mNDZGI
NEWTkFhEOW/f2OVjdLET9Qjzst8ykO2JcT20gjA1dBe2JxAtnRZXypgo0Qsh2IuG
9/533KnodwPQWOeN5QcrW9SDetYqh6H5Go8zPRKrBX/56B7yv7eFP8dQdIJMIXb4
Oa4pPI7Y0DKaHyKvIXxHKOf0hWrcM/Z7nQW99lBjWGRyKazUpkTHLXct117U4pYV
PVv2d+/uNLgyg8TJf/Pt5WXAyRxRpQjmkmsZRRocdIPTX1yMbOvBNk4sExH2pa60
rfLaXryMAnkbwAVjxsIR5V6ZYIFtntBkO6VJhMdkYT6JmANOG/hrgMZLcsysMQuG
oPxGZBi3i76S9nTWqSDu15TG7zVb2v8th/c7B43X+BRxS+n2Ii76iJyA51PqZCoF
CZx0hXgB62sCWt/jbQ1oFkyoZNYYfZZiQpI24fndSvl5MCTfhT9lQRr/p9h8DEHI
R4FGIlmP4b0J0vydTMKhFEo/zZrRHxArvUcthogjpGkG1A6+zZzDiVVbtEpT0k/L
gdtt0rn/JHN99M7gG7M5nAFw8bxFM+3EtKolyH1NlI03LyqdFZU3jqdZZbQrOVT4
/DBH/VRq00KuGdCUiy55mSusNQQacIAK1E9UpChfjexD4svgqeufN0A+av59fpFJ
bPjWOLpji1AvpoiSzAJEszcWKKChvCPlgTNPcMNvgpjwzBfSpLQM+MZ6VAewOSyM
iUF96d3rpa1vSVHtPvZ8KykDp/8WEtO2MRiEl2j4BNk5Juwmw7yfgGe+PnW0DjHG
6ltNIF4ST6uFJ5bfSvMj0XebAHteTlnM2ErUE7qJD3A441F8IOA1O99NRjcYKK0f
pT6ZPBbW8Teo1CNEJASrf3ezHQazvoZ/CSveVYG842uLv2sraCXuQXO4kYl28gln
JRQPHKDCesMt8MmXuIXLGMNgGnvf41egX7VHJqRgrikU8t8ghl+ejAAxj7znu4Lb
YqzX6juAERjlGayOo5O+ULVUj/PY7jKh2e+kfMhjJQQjG9ksi08OLoPLsaFbBTfP
Q40xpp7/CUpX2fHIYVwsh82rn6llQzIbKqY1zD6bGlCRO50khqS/wZGDkHL2+6rA
JGb1AhHCv00IE8uyRhk4A363awrVoo/t9oD/a6dinZOQKdXM5irjxz3T5V0FwI36
XuGs8c7QjF3qwOBylYrMCwlW6I0XUEQYb8Wibb+Ooy/Wbs25Bp9fbRTmGUD/xkmP
VPzRupvPtqes7rz8pO60JniMPjVZBuXdcpNbiiWQozSutZbHwVypOW9xYO79Ul0q
aykbtT+IqQHLT47HPUJzqzXp5I2z+Zj4N1bacS0sS5KgQnw4ISVtzLPBwTEoxrxH
q75OJIHoajNrspSbQBXQXUKPiitshCWUWvCkFHAzmwHmsjK1ZJ/Fnd6bVASxjfMv
XvPsE2yoNptdPjDMQLMyeAAyK9OHecT3MXsDGG8PhEc9nibErG/lhXybKCaMxhlQ
Ua3dkRqtcEsTg7JPfagIsqrOXcPxWpYjGVgG96qIuwnRCzeFxuUbf6gafxyhp642
AwsT3b43UMa5xCD/Vu04Oofm1eWDac1xFNuCm2LQiw8jrAhBP65K2MD98VbO0n0h
1/Vd9pXfhONjzKMYvE9kun/aqWqztnH5HMnDokuYGKACY1qtW5gTgkzMdUe368nw
PuA9EmwPqLi2fsxBRfZXbhhwficbuEMjrbI1+23z4x2w31pQUH2Km800CHzmyg5V
cHklNpKKUGs4YzWqVTQR2G6Oadu7x5xfffmBma3UHQlKvWP+CM3ACy4Nb0sclrdW
RKhN+XeDB9Iw/riZAMfzs0FOi8rupb4vUKugGMA0QxleV+egG02XL/3icbncZyeG
+/mgUri+Gdj/gsWjAbAAQs4PAOMXAaKXwJCWif95KAu22pm5CIDhD64D622ny/xw
sqLS/R93UwL+FsBWbeJicqDZlDMKmjegFH+Tpr8a9WRHYdwuIbTHrLWdVTyVegkr
i0qmhxQmTWbEPGTU4iHek9dkpErDvRwPTE3+O6+5gPxgGcssOT80TV4Xqv6JPk3X
ctmIwghGkwLnaSh0o4o+uzxlDY7lo7Ne+yAjXKsjq5snqkestEZjYgLXq3bN3f8N
vTUyj+SqMr+SBZgCCkW2OteiRJ98zHwfE1Nn+PCOJwblYxvi2KRB1pzWwDyuG7k+
simCui0hmsmOmoBlIEXHUsZEzEPsALY1SRguxC5mFjvUR5+oSdrcXH8giu+Capu3
m9Vd2qFjMjdUZ6W4jiSgJNALPkzZZQcgBgeKK8vTaSzsnpq2FE/q29/7I8zTQqcl
AbDHQMkyfVvOwWHWrV6XCe1efsBzdugzD6eGnWJ3wJJrHV1LWIkprBwyXRGs3d8M
DmcZ29eVDirjyh5mEXEiB8TTfIj8q3jw4fZ42wyzuDbOfqd395fdMutqwZy3vc7a
r25/0JLbWbFXqSLCZ1lyeSamWDs9EkzeElavT89FibBpOwIs4T7bqqSYzUiXJmcR
9gGhqxhKp/yDpgJd8X7yl2m6RjlN68qIWbpDfZmzmSIEgCrBDpoNKNU4eR5rnnOV
bdeQobTuE7VsPlVei8eZxJ8jVzqWyq/Lh9GlyY9QCWKGFnhYKQwfLnWdYG9bfb/S
Cs0ov7TG+Gn8eLZS2qqGM0KD6v3aC5tP3AYU2y12udTCJxs8DW4lrCUArTs7pEXn
lP+pKxNvyHg1MBpkMiZzAwqQrSSBSiZ4xO1alyYENGhOYHH3wwolek85sVORDhBw
yNJSnzrjZw/h4cDINaSWyZg57k6NkjGiMaOGz4Tf9KMESYXfCOQb+zh5zPxCOTin
blqcrrmUlD/ddJHKdqBfV1XFI63QWjDp27iQFM3NvqN3YBjOVadggTFwYR0eufCe
uaztx9ygb0PmSrEXss3H1ziZLnqvVEwUagSSNqAZltKOg1R7PJunk2mXqiGO++Ft
3zaes+PgU3APLXfJTFpkJY1jmJb6e8brbVX+Ikj8IBrCehA8cd3herxvCmkKI+V/
pyGhBFJp2yaYA+0Q1foiiCgXD2rsJXWHE/7QHpflxsLKkxcnJZ2EU83ygRVUWJx6
O/PK6Sjd56V2RnJO/rQ+v4HteiB1/LMqIryGNqVIb8iNWgICsqK3HSJ+BzX5GRDA
qo0KZGtlpEJagnr7i08PynKxQvR2jrNZBGaylIMIhL3xDLs1YmwSqn1cJPJeC1N5
/gG71Q70vDdcK8IQLWoahhoZLVbcrzTVYdrw2HzCRjq7ouJ8iRuEtD1tXK0DWAJu
HhXf+mB4x5EC523EPS26jaZ428RHVOLZy9qOpGc2X5yEMuGguiDEXzSvRuphjheI
OnAMVqwNdZyWgMsULCUyfPgjIFeHIjP12u73qrtHu8k/sg5G9QntcgPGNwH8loxQ
0be12t6xsqmgNiMtwEo4QxDt99zxuuuO2Jqz+hUBXVpSrqiXpbg4Okd+uA1MUbUb
ajSQSGPh93x8YydtkKmlGMnqBM/e55n0tAGrJ7CUbVSKywFYhXjxKv7e2DoQKfu0
NRdmvIogGXebwcQ5Ti320204tS0MCoTNSjOS0aN5cYr7q8Xzz79uzggBHe/JFktQ
rSf9/oV3UnR2eKe14d1oBbWtlueNexaTs2mNlSsKNdFV45QX83mRMigert0GzcqX
KhYMA84ZE+XqdNkziSQ5xEqGSO7oCQ5NLvE37FFi7AusPkN6DGTyPdA4wvQj7kPA
ne5sWmpfefKcpV4HEGWy5MFy4kyLsQlzOzD8lwYKHmT1IcdsYaKTLhPGt88mqWLO
50LaMgS2qSUQB4C+n8hOP8vmSRuKDffAL7mvePSUWAfkuIH/nq3Bk8m2Nvz55MnA
S475XgdMU572hXNFBF75RF0yXz4fgOwPIM3dkgH8nExElFd1XXQ6zhzaozwqXSQO
wBiiOzfDWnVD8Y81oWpN5v03TbhzO7K4KDBYanU4ijQ0b8y6/YKbPqZcSqPm79aO
MFZrjScpBPJFFng0Ah6xjqMLZtTi902j5mrPBOycnx9UlFMcN9VQhDpDNj6qYe/w
sIIYnwWHNKOeS6+ZcIXSnuTnpJEWWZ8AsEy2HqErN+Msba4N0U2QFGTm7Zikkmsg
WO+sxpFCLK7oojt+Zi6i0k7VzB/2z1R/9KkHglJfhty4fKOnpLq+O86bZXsB9s6F
rW8+5MM2IbQhTr89+kXVHswAyk2daLPHE08DDjefUQMbvSqQQRBRpECBpEUT3ltv
cpYanbyEeN8kDonhYdyOOyhseW0Xw3OodgFgNUwGPu2ndr2PlyIeNNZZ4FNEeEkL
SzMx8dTEOI2rd/4Qw1mmru+J5oLrXvnpityNUqV/4rfsynzRE7Y+gjy+spDguBTh
Sv+dvrdx6ODXD6VeihWQaTL1zBlQItGivAfwL00vCRiiLcdg+lDTlMWCkJvhuPUx
DjlpOX+Fu0TxmaKDoBK1fqvgaAGcXA0GYh5pCxhS9jJn+xrOmVn59Hdj7EGeNiOf
j4vVgb17cqTg8cCOp3DofRcHwk+K7mGXkuJ0natZ/Xe9QCU1F0IF0JKgoBJKaVH7
IsrE4FWjrnNxH6OJsEErhE99HDSir9ciXkq2V+lewDXueeNBZ8eDvLIFiOGaVDea
2VjRxq/VhOmUY9dhxZ2cOgVVpQp8H7MmApzXw4qXovsi125pjOcvNNLX5FuLJUK/
lSVeKQN3g3SmGpTNKMwmG2kqyFC+u2Zfcaa3HWlvjN+FqidLrzni46im4ERTVmGm
5FUUucuzKyQKdZxzJYE3X9YR8vcV80R5SMvyEC4BYTJ0qKnm4cuNT27nzueYM7C5
2B7mswrJCPaB1plHkXYsHq/Xq7tSyLg3X8kPswwtf8RLmtEd6GKm/YzXmoh2grSl
d+u8iw/hdjSbf68CJJRFh73IKIHQPE0Urbg2fT8NUecRLnlp00dRoR5x8mn88WlF
a5z4SFMxw8tPZNaq4R3z+Jva0gCgThf2vuQIegStEHaqhtTgBBMHYYkd+gCLjCSD
b6yR9sUoHa5oCoqKB7JIC3+EvcPI3/zoED1Lz4qVFf5YReI1IjXini+TVJMktU1V
Nu9wRgvDhZ84jkxpbW7a8lJ7WGakZb8CLYXjjaXTnJulwev95jdyNe0c7TauGgUj
ctrSuspjeBwGBcDeLlWZe6TxuTFnnDCFXtTKtzVj19TKbVRUCKKen5HOHZxvb+im
lr9hxNxTiNz9VUONClWuetCUy4UG3XIR93WHJ5qCErofcvuojWYsFSjXI94a5+hn
nNz4v9p6J+ERGQd0mA4XvzQwNELxeiAvI/PzK6RdykYZIcMZ0sQWuj1sEBWozmMB
PlHEELoKH6tuQwCsDKLe3m2o5fnGgho5WcKMXmkQH2NATaIOCCUrjbY8Ra61xLwL
CuvXrvllwqOCdIdpXhq1ndUd2nM4rFAQNQmF6/LzVZF6h2HnbOLp6AEced2Rk/NL
O+T5IE1wadEPuTYV0JkuMTmXL+IFB/zcxk9+divXXxJyAkLfrzma2GwiVn4NQPIh
31Xtuduq5aKX1d8QMfhUd+JUc0XjTxM52q157LHgGREj7mx8Ni+fKcrECQQ+G/MG
AByFO3j38qZsYYT9LwxnMlJPzOlmKuynJeG44BTezeP86LAefHb9yVWutm1k6gJ4
zgF+p3pofQ/T8dMyodcE2VH/Qn+VQi6WLmmWJo8wxM1jdSvNrxhkt0C+ZCegcF/O
mvM3XUwXQmn49lppRvWNI7rSAgmdT2785ZkYCJ3LBTmnPScLFmgU46AsNFjkqHhr
up8z2aYQE3edxZka2bZH/8BqGDGqZJR3dH7EmjbIaq0MPEhC0lKrajvZn2AhVS/4
FjdbaqT7pR8JN+5kEbvA9v06783uccxm75JmYMAZEES/Ik+bEtzSIMo9nAsdXvFh
kSa81NI044detgOlstvHNF5CrYbkM0Djr4Rtn+asxm9uqqP4iwnHWY1LrU6BUu3J
VerJymLfGWfvF/a94gAxd1pv9Uo9YKQUMW3cwBDHwktalDxHyD0+Vk7eTl5HBCq7
gg0Pj4PBmUlqo8qp0Lm6UEThqvJzY8lcg/Vpf77D0i3zzpnPNJv7pBSG/iKcvXIw
gnY/mK+MmZOy3jR3A1fioIoc/oKqyjYTrzvfxyP4n0Aa9WEQK7xGMfszFNLBa7bJ
op29pw+Inhd7SJhBeVyTCLjomQJeE7pP6qT1hPc+nfYdCpQhUC9I9IrT8hvMA+mq
v9LWXCbHYUzm/qS2yK8GgkKk/sBqbth3ZNk7asUMWa11xelWhc35P+37vNzJ5gKP
9nLB/8GRZKyY138TpeHjc3ueJOZamAaycqA/ywQodzKUwR6TYQai4P0dkiupp08X
zIED5VUitXZ7ZM+M++EIRT5DBXeDxD+QoXfC0jgRsJkLqRZv56VBY/ZrARCly0RK
WBhi+EWytnl+UM/ryYKpGetMpQAN8MXoD/ydaiuySYS1tfkT5mnLuYJHHHPii7Ii
ZK156fRsalr1QsnpewGR+E6jHlwHW0dN1fWCTyYsMEGh8nakLoZDKY4UcD4M6iEp
VYEEwYAe58BvbBywMGgfx3/+39j/Dq6EMU4uxwM6LJh3zXm7KRB70TKucs9LBB45
1WxPfXO3Egft39mUbcxe800UeVYdflHk42YLvtdcpb5wRbuPGIYlkawCdq+m1zoA
MJuZF5SLzHB3dhq8dcXpsbqU/pL6np+NMJ03BmwpoJdg5l1FuAkAPM0k5fQEswiq
ZpacrCbOCxtBn1PtAfSrOThf1p7NIfqydh4lgxhZY123CGgwQ4lDORORNWZexsIw
5X0c77jxEVnPb0pCNIelaxciSiFZQmLqfwviqc3cTa/pdmnyAcxAx5W9uUou20f2
EfHGMe6R/B7a2//xzygIzA6OXVPu55/gFd2EzjAoR6nnCll4QXLsa580CbXRm47K
tI6Nfjjzv9tz3B1MiLoTpU62Giu0gZ7pwEKtihYydl0lvXdvzzGEtLFspdbkEfaN
pbBxpdEyelvMtPG+mQgNSsuoqG0q/R77WSkHUQAZ7K9eXfuZnEsXJTTiWvS7y950
J+D7roCnkSwVD9PLZQfs0KhtBPWY9J7PeT6TLmFSG3UpT3/ZkLdERImwwo+xWqfS
yNCb8WVd+814oGlXBrfGjBrmn3FeiSRJUkXOVi+fHHuHqNym+mgu20Rd/5G1RAHK
FrSfJevO/A7FVynWk6PPqmbL8sQxJJzT1g20rAu1HuEpRsMe/K8FKTqwLUpTJSjT
WmCv9aGaXuA2uUJfNYRNjPlGmkJ0QOJ+qK2AMfP3Cf9dmtj0gLO9L3JtzNl6Z+Z0
afy4TQYrp5qdaUhXklTVWojJoK/M0Xryy+u/IX5/pSMTGB61za3niH+53UhCqxlJ
SYi16NuXXVfemaRHcHNp4+lHh0Jh1pOxT0msUrkF2P+VML9iSGJVhSsDFDPxBM+2
EY/WftqbQXoCKsMH00l7hqxrXG068FWRLhdResmkQVvxp+plO+nPbmGc9JpW6UBU
DQMV2jRptlRT98LvpMPR1b72d/LfQaVMGwbcV7dd56v8byYUOkrqfTCt6i/HKFWy
GK6v7UO1X/h9J04QPQjHJhk0K2XcUfH3dQJ8mj63dLSR3XmlLhCxW8WZuujS+4xz
Mwr2MOZOVb2gl7w61KfZEjmhxMtoMmii9Cg3C9zBNnkIkO7vsU6e3lgKnzbFf+52
AdJknWQ8lN7DHioT0nduxa9lUBCacP65NWdj2M6hSsSoml0DGedKJKpuXWiXfLOf
zpga3FeLRcdzyIDCec19/YltORubTEwCjq3d1fIQ+dZMO03WWbANP/O/lUnxkQr9
9JBYmSdJCpBneU2YFeucbKz05TOlaDqMSwE03k6IulNdUm+WOoUnSvNnxdbTJozE
0Bg3nmq67mb0317hRXYsvp4yySIEtyXYm/WHeB5ig9bBZ3q/tYx1FkeUMVRrBFf4
2GWDp1YCIBOCu7+pCPQprrf7tWLuxsWPbKe9rILPhoaVUXrSmcGUQfDwK1KUSNWL
2tAiv/QFbRXUSIoSOvNRAdBfz+Xm7SrWnncyBoj9Vnr7+G1ERbblfN/fZouQTKSA
W6DG2ebhGsZQ40Xin4bL2XbQWseCZuRaz4qJafNKQpaPgoxkDeKyBRAhHZjDmo2O
l0z2byiORMFzj9F0YSSQX7wvcEClEpKbWnqzN1N6ObNt6XYjq+IGZs8ImFDG1c4x
iixHEcZWgPbeUsJwI1d9KudvKaZ7Vw8dLqGphjUMkHXcHXx14qnfeXIjZI73aCUS
XH0i/3i9+uef3r9Zzv7Z4nwaQIs8Ca+D6029ihHQ/QB6zQIfiidr4DcvTOKSk6N7
Olx1rw1XpjVhppXiGupabdlB9PGxznMFo5O//bae2O6DiHdpAfeLruiRAmD4oUxK
1ZkLg9TEFDfXY6ZntQsiT56SWfWFJ/T0+E/MFEEncLyAx1MljxyS75PrKB7LF+Lm
2pFiIUT0p7QPpEvPyd72sXZ1i/usaI4N2qzZFyz0dOlMV71nrwF+EA4/fIottAuS
h5A1KhyNjaq86GhHTuinJAqJK7x1920I/mcVt63bZX8Hn+rzFu5gBs58sza0myMZ
q2r7B0pe9ehYF5Kr3cC7zli/jE8RVvsNLg5II+Suse72DSTbyC6rr6b9QXwcdb2N
Cf4Bl/n12/U2Q2EhxQoQNw3OQmgxGUvSCgu+Oog5kxAZww5b4k+UmuDb3HFHCXQQ
Wi1unnrRizZSlTRyqDC7MOSoUtIMYfuT19XqZHMw+vBR5fL+FV5uObuWgl1JDEKE
7wEQelwAJbgJu4dS4MnHr8CsLEMX+mBIfKPCHgoYGEZAP0R/Rr/u/t/vhf+eCTIY
/eYYqjF54DLZ6YH5FCZ3/34PWSzfLaJPNplxpDNMkeYpi4r1GDCJzxk4Nn14Aefc
qCq/9TdAOW0C1MfZhO0SGLL95muSbhHbshBHvNUwMfPaJxiAnxfJz+Cew3F5QwgY
4ZnvtutFa0R22BJfm0uu880SrkFAUqnLfDBau0ggS2c+fuGVjP+ba3Sl3RsFbWQ0
3TrNa1Jg+t2PFsA/KJRMyC9CnfDedBKImvbl4HdkqHUD0wlN0j3ISNpqsirelp6N
gxWl+KpekI0iD1SHGmQGUR36foEgxT/3Oj7UXixqRmtbj5XLui3DSXQBlahFv95C
Nj4o869tu835VRUvFsNLbQpHAl6tLArJBwziKqQChdjZKiUB+KmsU3rMNlziO0M7
66cSxvdY0y69IcP4IKhR7w3GG+9dKmcWIKXlnYNiw37jXExmNMVeLNTXUkdSohhQ
dhf6X1xjkLgQzv3eiPJ+MoQLUY/vO4d0DNz6MJhcEX0bp/Vpps/cdFa7NsP3nIVq
s6bOB64Gcd0YpQ28LwsUKWFId+g4owlEoQNawa+c/TSxSxt8fzz/t2KCWTiexSN2
GamSaQSDTVbRSm1wRVazwsEPIqDpAPeztlwfF4OTTtkRX4HcX6J4TT8lJrknaZle
sS9VkSf1hZZRgIOfOI4A5+EJ+3DIXEf6Tr5If5J3oAM5cvqpDXG6bAf7Z0FI/7b8
6PDbRHpVrx6GU7mnIJiwWQWqpD27iamdrXnBqJqxgvEuRylwbmMPe1KUtvRzV0jf
g7BrfOCWZOsmbz6xl2myMaxX/LgB1otvmdrugnjPiytrokjLbUL2ZXrk6X1Gnxt1
FqPWluYzo+/LorEYV73cg3A6RXR8xFkcMmNQc+dLX4huqN8cMqju5dh6a/g2ZZ5u
q6UOfmh17BBmeps+kOrV62sLvoFzU8GbK81Z20WTc88is4miAAwnUzEDlnokW88w
+PV116n6tdQKj8Y4CFT6tmZTf5DVW7ub9rNWDRKq7EygcrPyY1Ei9epwzz06DFD1
8ph4iikR8RKbm/ULiJqMM5FT5qlkgd1DFHQ8bOS43YcGhFnVi/O5TxHXhWQB8lzv
WHRecxFK1VVPJiOTKEP/HoUxgMj3YzSdn1dhWrNLBR7VDHr4lYClKMXetwQwdhlo
Px//AE53OM4A7DKrumOZz7jELXCRY7hDhNWyB76Yd6Mi9PjMHygGWka2l9z6SWZA
k13Cn7mIhQedtf6zK5cb/37aekOKwxijV9dM+L4YA8eSkiuOhhnYmWD0wHfQekCb
sKzU+dvvNjsp504D7z70wX9yn8JDyrZpLc4iYYoRBPho2u3PtXQXeOxaiEW4yCq8
+qzV5zqpZbAw/cMgHxrVt8J141AkB83CP5z7XnPNF15h/kNdO4Q5FJdtw2JO3Nj+
NE6GBtdWSYQ9LkRp+cAg3bRro4il1wL8Zh+EtZCgApMcsnyNBqSS5bCrlRKhQjXx
IP3DqphB951BLBs+NC9kBpSgRJYIdk/beHXwUuk6hSwuOLxqk5kuIyxlnNqTBrpY
OKsDYkK3DbVLOV36dAfqj8jqZNbQEwwnJDlyg6SNUlLdYlNvtRRLmrJME9ILHqJu
7W9oDJr8rQcDmpK9S//200+Fr8BYcUYDkPjPHbWq6nPluCwaCZsIG7u/K8JXnR3W
FexImAbi9wBUScdUd4/qDE2ZzB1B8Of3fDVao3WcdLYeCSCyNNG3i/0R0N9I2x5R
SjJGDzw1BSw6auD/fvAqNi+r5+nAIsb/OOLIbbhYwpOfrEtpyv50LrSJAA9lAbPo
605khRKjliyROh9sfQftDkFyvmAqJO14Mzr/eqGgcuUjmcTm4PxsOF87UMnmbKdc
UymwQQpOcJGxz59UE3O8ZLgYNupz8YZMePkU/8E5MgmGMnhLMuumzCLR6jqsqdea
CWcvujEVwq4N+ImCG4sHAsEmpxBbsef+iQFUAtdaCZr4llzJefpMKlnDP3VmGr/5
Rfsm/IqvbqOWEsU7TyPHhPtuIkk3J50jtLsQqHUU9MQ3I0ZusxNpI3UHMmURJGKM
1K7GCcKx18ikKXffAMQUvRPoAvuEs50x+1RtyasFEyi/nWsFzs/Wh6AeOP7PRT4R
h3D345/E6a25xKIUCLV0e7i3IZDuNDdu8hh7uzpm3KK4lFtjcn/oSg61eB5X+ZZN
i+GCuhck5NhjetkfYwrAG2OESTlsalufFKjx70d1m8Ge+8feK8V4Sbqj+qJG8j9J
EgcHmQwBAoz7hjgYlv0SnpOryNCQxrGVhsUOrlVhE+Kg9XKSigUwRHzdz5c0HDzi
CkK4iG3rFii80fbDhcQGAzuVbo35vruCOevp+zzxiqXr+yWpauuDlZf9Y6tyYIYD
ygoxR+IR81dw1YpvDumejBaMKo9Xj494wOvxvD6qys7N/2sdksclGb3GHuBb+UsX
up4+b2eeZ4mo0tzDj2BE9PN/ESrOlV5PpoSXovDsK7ZP7ErDj1gQeyEhztXCu/Ml
PRQE80m1RBenCmaxXUPjW+7D4QCt7i+SInmyHcfcU4ZO3DdlIykYPeIovBEHTsCC
F1UxpcH/trwwkXoOS4hq5UW2MK5sm61tiVJTs327dTjt7hIG/MvRKd7FGUd19Iwp
Ohoh2mi1fiXeFoieJKKzdJGgy2VNB1cE9POdyFsa4Z1gO7M34yU9JRvmDH8t0Oa0
BG9ZFp0zPhScImo2rlHBvJtnhCWePfi0c/EsK5IJbt8r/MjotJXw2WyK0z9rCitL
CdNG3YuOPCV3ikSkjhJm10QpHhKCZHPkmLOeYwGS+EeuOzNi6aYGYlDnaIrwGWXz
U6uocBpQFS96xY5OrWAZHjpBUsYZLecuo2++IkxvR1UHW6QVJTBtU4YT7VS1Ohp5
xqtbIz7I3P17Uedz3oXq6voHu+fVTKdaoAlHWreCTmJV4rm1gR22rmz3YtibRG4I
D1XAYLsyxVvx56c4vhIKgGYkyUNi4zbFxC+46meX9GLym7j8/AO+pc2K5LEKUV2W
eiyChaklbNrpZ+Htap1GJTx2whcPZmqBQwjbdVvAmu/MCFp//5fnHYODkBpBvc6a
QL49HAY2QUBacST065w4aw7cAfp84vMagKpkjjRydb3SCwsVSS47ukkt9+tKD93c
kcj/i22ntn3R1cNfh9w/HEA8OJEFQlaMsDNLvijCsgxOmHSyXpnTZYanFHdxlViH
lo+/jCY4P+2F9mSTuqBzkaAXqJCHLhn8FwYQl+NIT3xr46rQDxWkmQv3SQKKNHxa
lZfpPJ9j7YP6Sd03lf+1QQwwIRXhRkdWurEqOTUw4D4N7gOA574W/Dn58Ese+/Jb
oXkHQHBxJqq5478DD6ckADOoRiJhyLrdEA1gE3Cj4Yp7YGB+f+Lsn+b3sBj9e6Na
Z39xqUiRMfFBVCu42jII+q24fMhsc+VpdPLZkam3YibfTYKTdBCylBJHZ0YvhOYC
+Mc8lcpoKHHan4Z1tIL2OWgdbJF6pzZCHIYKx9an+sGsD/+UU7ggx6cYS1hnX+VH
rdrmRkegkw3v5vR+uCphAa6ouUKnnJCDS23Zpu+yZHbW/YRzlA9oGgXKDZubP1G2
LTeJvYCdw+kWTvbsRytc/T4UU+JA1q1RSB76xQDGXWR33mElo0yX4yFyF7MUyTnJ
0LCJWivQuOyHlHhF1mnM2CZyg3zbGNmxyZ0oYORNxere+OYCdWowgtoIBY8hCgaQ
tLLuDlBW4bkdJcaNmdTrtiFSYEf7w4cYyH6Eb5lpFr+mNMMJwWIBWeBe0eKMDDFH
QXqx8B6WTLiunRUVYLNF/uMagjvuxWSyUFd4S9tiRL3NI9bt7HdWI5FdcvChnLc5
nklfYQoraM1oKZ4yUSzncV3nX2Vep8DnQWiSANooGLh1EzSXZFm9BrD+fA0lvk0S
fM66GMGtOJWnRukovRIwACrQvwwSSpeERORgpnKNhssF6xTnnUJaM34+7jvXJANa
Mn4bZIg+ZJgW+ZqNhrPB2KLmrAGHSxkqtfGqol1siUvtAmX+/wOmBbLlLQ4x9R1q
oIIfd0OHeRszUPRlT5Wi2oEwOb1KaLwIkZtSPOTdlKc3JlsI5Zhaech1XCk3ZbNn
tNnBJMKTPxeTIRXEqoNiGHakTYah7stjcxlEaGEg/LOBHTX4ddUARgDG/I4oCKm2
tDFXAec0MKdV+h/Rj4A3aQ7MVXIgVt+uCr5E5F6d1gw7H5Ery3yBprHEx3g0lLrQ
Dqp4eH/YNboGQESRXEURGhesqbhDsc2R7SjHKjIgVcheKNC0c4zzkgIc9wYsqPKo
CwlXgwO1zryUxSiOhninXcjuOdzVw4vvgbkKKGZVS78LvEBy3d2cafwIeWahKBSh
CRkSw/5RkNPwS53BIsPfVjYdUJmjoxBMLVJ7EKuaGwWgp/vbaAmrNMWqpT2uniQi
4rJNZl2+JFFO1CyHE7EFUEsR/HGxZ+9nd0NcJa/epLjVk2KyL+Q3QPQeDwssnw5A
zhZLCXT7vM6Z+6NW8UDuJQRQM9TivfPcKtBqlAMS/mkqbuZXAEp95Mmmx+f6CXsm
/0fvoqp9R2YEANCpUqY+tZizPDWsUW/zP1l+22NzrcmW/ZLYe+F4ppYcCvvEWvBf
aJ7+0QeBqEWUqTnKV3Kmnq0DZxdoV/JexeAhwi0QayvjXWq8ROBCY491jxRhDeC5
Bw93QnTlKdyFfmGPd4t+UlXokIZkYWax/7e9XxYJEqrSgzejx4Ze5oKVgQIbMpdW
1TrOw+Ypp7RBASfOpZHTn7ywc69KkjE239zKkqM+vuq6S2vbVihEPyWwZ5v1Xs7U
s3xaNgTTiD2JCcfN5lDnr1IBuYN8O0gKlBEkEQMcljIIJ12b2YsoGtuv3Und0J4o
Nl6LS7C2HLacruz1wIOosuNcOv0ygg/t0x4wDmn7CgZN8PDNhTFTB1EyMyNmTGs8
zZxhFmPXhLcGfRDOTE9y4NRF86WiGeZrAjg1TbWkEfuSxLmNEAxaOlqTqbQ6dzls
ZATreIxOj6PCorT8sWGNOog1dRDmgUCvyVTRi/a2XsZW6g1Kwuzs0RKEFZtlnT76
XSlAPHpKYcSJsUVsdU8a6KaV0hbgYu5kOXBVIYgKxWxzTnLYwFTSgnJCiZVeD8nC
CpjZzk0h9/Gfd6KUhU4+hLS1MCMWzeVWvpgeSwpKpggy4Lv/ajuS9Lb3JQuk7Pkt
/81IJY2CM2SmHXN9V40lsdJ4anjVO5g7jO4VP/fwC6KOPa4S0j8P6Y299lgtcmvj
Dd74y0HHI3s1M2KeUL+s+AhI1NlKT4Nu+V533nXpWHaYVk7pwPwplDUWsHrgSZE6
xK/+IjPnNpBfhBzh85s1QI5k8xXbkpNyO0EAAEIqU2XAhGK6WHDysrLpasA9JjWO
iV3wVkdoLROeOczXoTxDxoVhPuDKolGsxU6li1bZjE4kuLgweeh1p2Bq1lqa8Uy8
cE31GlvYc6LkLd9KT2nxFrBs8onJh03NjT3WQjxGHG1fg4wKxLIf/M+WqfUBVKwN
qPevdybFTUeuP+XzSjjgtS8C41Z0rI6tsZ2Us4m0Z2zSRrlNTcUxa/nsyIblRaAn
Pj/6fR415J44RbgwYyMJlwrS0n6hVHKYnThdDZloRAxyb9qOW6Zkbk4HTjKCJyzg
nSy4LNs4D7sWhhRZungwacr5EVH0UnCG+bko1uCMJVR7N+d6Vq2TOIGxn0oxBXgK
Uex8PaFcgnBzSJKXK+Q17oPiDEgJvV+k4JwxZTILj+tChTHfjv1M8aDfmJjJwecf
1Mie8Z8Fw+D6gjYVcVio6o/eGXj0nrNzYiWBxosRwd14g9wR1np8pfPHviN5Gunv
2rqMdCNfKf49J7EAAC24ObipUWkFPVOObECAj5nzGWnndNAZvVMjTl04yW1chSgm
Wkyws6CdKhGDzivkpJa85l0qx9OICdmIxNx6bZPUfea7CrvIKjpvttI7/tUHJK+p
YEk3nGNkyFucXmgSI/ggBtANAniw7RdNTgYaKwTrJtImsNvfOHU+uMM+s5H0mQVv
pJytcjTgB+6H3ErRIZT7Spg8JJMhdR33rB4MI6KijL6sXDr8eZsZvVX7nULr9/bC
YwGrzg5GRCImDDSgNekgXt6HPn6W8k9wBtBQ3gOBQU+wHv5izlPShWZaL3onM1OW
9bgD3nTyzPtaMJUqILIPUWnkER6h7ou/xlmYRdY68vnTz4251iVtnOOuvQagVqKU
N7PEBuXwnvJ9cy16v6CjXe2inYdPTfnpEjbI3I9D59DC8FarRbb/RnV9Sb1ho9E3
+cDBpy9FoH1+WppWnMuUvkIN/pFvmLWgIpkMM8qRkVPGDX2bJWVVpnpggZquN5ae
VNoFTj5ZzGsSix1qlmiaRdIQI1KEr4NxE+MnCZSEctsOPWyzLQNjWORZ9JYpTeoR
7i2yBk+Mf1dNoIAObVRy2r7AX+1dJ9SPD4J+VHgNtaY3A5x1D4Uk72MywF+aopCn
A/GHsjYoZ+wycdWzISsXLUvq8Cbl96ybqEU3R8OlnihYaZAsE4JINrVn8HpSsoNE
v28YWIgLlAMEq2rrJNNbaLVIkck8x/fI6rbdb91w5E/xbnHj0WUf7k+DCQ55LOC1
FqEfBavoc4liEy2iS/15S9E/B1CSxeY2Hi0yF08fmS4dF9ByF21LlrI6ZLtWo8Nr
Hkq9VxN5oEGZB6uEXyvGu8dJj+smpOns+Urc3Xs9Pd4EkjN7AoQvfoWcHypdPqju
L9s0WvEHw0n0CXJkwAG0d/is86tR+RyuXYJcBCzFVqcAkgiT0C2eoUZXsFrh9hgf
RPel+UHwYNiPSxQr4m7kdbeIkQ1ugPy/U0SO5RcJEKKGaUsQ6UYmY/Zxv5Ws7PmE
1Atepz/XiCI0wIDY9O1XdFllnU6uNsHVS5M/RMunIqWJFNXA9m+30w7+eo4Xg672
xchNknRYvPUVpABE+PpAAdz0lYrjFo91jp80RALPZ6c3ci+qMS7bYRjFAokQy6r2
yRH7TnTxpl6S23FxG8QMygx4HtrJPnG2CKoz1y2GAK0q0d1fVh8lIXhfXXSIzUpW
wWFnLaz77rVVo/xwDpCNksmaVsDWpTyGjQEZh5SkJnTQhx2G6/2ez5ywtRIIY64V
zHqTmTgGWhuT9wZ5XMThxBr+3cCY1uuhW4DPoNFRVPQLOmpBrSVLKwrXPzfTzu5K
VbSHYfWAGg2JtbCPk1pmntS4ka9KmAUaqZ2wPV/8a69gYlOErQgYB/3lKJQqbKwZ
+TBM3kcsm2GDTkkxNjXT10LgTmQ7zhdHEpRXtko5xnqNXhrxjIxdGhakqmRO2boa
nOathqrQn/4nILrhloJANtJv29D6mrtiq85afzikGZNTMPKM/K5Cpmgkc9EHXffI
VV6hKacCYMpqg3/R7rj4fGeEXLKgfN/qaeMWMaiYxI4t7I5e06fSC0moprW66s1k
69KgmzuvfJfn4eRSyj6tUqWO4Zzc/lVT1KJIsQGJ6WA7pEUH6Z/efJSuQmD7xBmp
YZOIXY9tutKR097ivZEIylX0IrW+5soW5sbIdnnLj3Oiv0mPIedOgV+cG3DlgI3G
84HWfIqaAzraKnFF6+Hysc5hKK9fSYkLrIVyMeg75rfkQNrP7i3B06gTdgK7vS06
oHvcavLbLHjQ69wc1GjgcTJuDNYcnY8D7F9Bge9JrivNKqBOoN5VJU/e8lf7vYXW
K5e7nsISqUdqMMlXd1Hz6dJhEurw38F3/PfKHQ6U67D7jUfJF6UYAo0G28LwCU/H
pHxgAIuyH3X6FOhlhIdQXJi/r5NA/yEhZ9gW9A4aDpuxuHIxwgHGXVXl2ucVTYe1
9pkK/qjp0kB0wlzs0ia/LxrsiZB38uk+F7WyGU0DuuZx8/oovflLZTJJMDVgaV7b
vTG8tSlAPRTsqP7Yjm3l6Ky0E8+R5N6mLwtmHtEdcitjhc4LH3F2fFKRo0yYUXnL
TgHHCZwz6L12cPTABZ2XKDEvR1VfUH3fcMwjKdJur65vhCp42o5gJHB+1vgl4SfH
iifkqHwrxhMv8qx759rRGV6S8+uqHSqSJ+CCSwjgKj+bt3skuzFQdpuF2gNkBdJ3
sRKJmz6YpG/m6i4SPGP3Y5DoHNHnsaYDhWpwR3vPUnBEvkRjvB+mBKebG3anGub9
nMIeh3F32kngIRkm4gNMj9d+0Zx9nJQ7k5S56jA3ZlpMPg+F2iowej1cB1sfX7fz
f9Wf0QkpDlnOrpS4Rd1DHbzhzTdY83zp04VsVJIGg5pCU/+M4Qn4EC2HInKpBBNb
mzn347Fj1Sf5775ccGoq99pN0NvN9TjhdtmQnz0eoRUjtZGFSWmFWBra3lyuzxK4
BOvppUQUIa+5osbajGS03OytJCZbBK1YT0BXcJPlD1S28wS+YRnDHJC1P9Of1Brb
E1DByWuZcOhvKZ6DGbpXQU5AVCCXDzEcKpgIRB2mVjyyt47ZlQvC18GJgioCIMmp
HsK1HTmurGKrB6ipkk9qENS/6fc41ze3qRTOR95OL7ozBWUc0+Lv8aUw7N2vRW0o
dxfOIWOe3ftFGMqd/wcfG+Lv8A0Cb+wq7fKgeWLaCDOdf0sAUIV88JrdMVgOH6h6
+KzVZbJ4y/FyKTP7FYeVZMB1uhy6q13YouwkARM5EqYiRfAXAVRfDKEujwJko8Yc
3Uq68MUjMPKS/HYkoCQj19mL4WiTxf2XIdT4xHBA7kURARpyw51DWo1vh2xlXtva
qrpBAPefgxaq2mlZLgZSgn0uRq/hwHQa7Gjy6u1d4BAfBMeb8yiscoEb1zpUl5ex
awm/oTqY6LzUpiQNwg75LQGCJ4atUQePvZnvKctLnyTuxavnWEKM6eRy6b7J6kW8
KBKg5AClMOqHnqRixCwRdn2tSD5TxmNNYOMSkN658pdZ/OqgEdcotdJxk/AZLkz2
a4Q1TGSIWqf7ONT41y2a0cghFQm/LuKvTrDy8z2BUhCcJjLOTWtbMdIjmeFQlyqR
K9TYnxSe1GbUPADWcrzQzYXV7OzFGMFOOA8T/ApFyE9VDFvzV6H1PjdmX4sGnOG9
3mybtUBTYiRoy/D2+0A/Vy90ROiGY9zWctTQtZZnhcfLGVpKtSuWIlnGM3JkXvyF
a9Uj1QJ/gP8r5jI0VnJypMO0ho9hyXrZkAYSHzN+drVNSId7TuC+SdnF6mDFb3sW
OxC49bvr2vsEVZx5nYJd0MGlrMOC6dCe/gX0g2hlw84JAoW9B7cbxFjVje69Ivnt
s/2TjV+FBaSitAcq2fHfbhg76JJsxsjLZdYLr+kE801f80KSkk5WTZphCUtLVmE1
P0Ainbm5nk4U2FsQ133dVs/1lQpCnRkkvvyMovIlAupy8o8csuwkg6Bru/2yamxz
Fw3IrXQbs/OcdUUJcnlLCk9EB49o/xI3zwkVRXyXe2ALCWnKcMI/VhCAxdjNRtXp
ODJZH3fdU7i9/R5VoSeXSOktj8KFuB6CebvOa/uJ6SlDGaTR7UQ6VdkYCirzCmEk
zsVTc/G/wVJc/xynbAOYxmmosKDviTw2AOiyAoeGvDK32opqPftcE1Y933ZFi3XL
jG1Ervp5mScjwmvoOE+ODP9uTZdA+lkfCquYVLN2pAPWWBdmYXk7yL6QidHZ+Ww9
7/lY2pR6Kiiraa6lFeslWsFnQ+lXc7w6gRC43pqy/HXymZ9nQmEvJJOBPCkQbCYg
hOgUQ9w/QfR09xzrt4iZJurYesIgUrnXPDg9Hsw9PBqkig8Ymc4NCQXQTGekBAod
pBljH1/7LvoYxlJqDjYacji0u0oZirFWrSZjtr0ddtVCKg0yGEKth8JjWCuaRev5
SApV6tDRY0MI6MfxZeL8Z8Kt/ZQS6vim6GbESElvzOemPD42UZZXcGfY5sFWrDek
DErf4yLJi58Ok67Oo61WWTY4Dc0aaU5IQ6FdMWc+GnourRaC2RkByUO11JJid17a
zsYoe177U1JzJyjhoSBF6cHiQbsI21qM3AdbL4ynBO5YljiH8eCnWlJomKpfFmyc
nwxTTxdMi0bL+EOUQcqynX+iFWFzry8ubp99118cdVym10v4OIWSRFmJ2Uudsxke
rOg//zjRkbi1R22lHAOWEfXx9I6arKRhhXQjbzyjZDUdt6s47eaeezWPzHt8Uels
k3u9KnD1fZP6HS2mUl4lh55Ma/hi7laKw2h03g/6r6/FA5bk1lHRKScnw4dVvno/
B7qjPsK+cBZNYK8nZh+H9wbfZeOx633h2HwrSHpaonTSnJ6zAp4XNPnanQOMAKR/
67z1LeQp8e69+RLwNGwBNbFGIGnKVMJtg722AlU72Ro28IZX1hJLNezLQWyUjI9y
mhvgwPIpMzrF9A+/Syd04vQMbLLlfYyaKedTx0ThIYlCJBRSON30mPUMzYqZxANM
/btL0n/pg4mL+eex9YdIHBQQMp3Dqj27raglvb5rX1sjQbLp7AorRCvMJ9TTXyZt
97wct+ebUYUhObC7lSS4hRKO3JaVvbOU9KCfdpg1evF8DjA08+LVHGBEGo6SWyIA
dFAmGzg9/driBysoTLj+XDOjf4tRrYjD+Qx8jPqYVqvrfEAYeV6PUlXO899B7Mu9
CxjgxwlRwY+OCd4nW5U2uEifrnHL7UT2k7UWryo+EPgd6cPeXMQQc9KMR78LurXO
vtH91iOm9rLZtuFM4jrQxSdXpww1EVF4e7lNlmmZ/gkvJwwLiKOlfkxTVBwUPogZ
cTZDQ7JZHE/weQDkDMtKC3tH1S1apTNx2frgpdK/xJe9/uQ9tQsXAgqXwYve0K+C
/s1/vsIA0npBSWNII2P0GW2LAmOh4Y8wQIBc/dui9bLcXGq0oCqaE6atfr9FCPJ3
5zhu+EvxDkYt7Zo1ubG1iI3FdIXX9kBevxSmpCZefhQIPmDIZCzXxnba+HuOGKrI
moij3wvn2wqcmBvcOdIQybJgNfFBz7CdTm7VH4A1GYE/i1LY7XZxVTfB3oGXuo8U
nMoa5aCYaHVxZwiSOlDtP6p0F3xLMQcw/nDh+zHaz0HYFvv15plgIdAPtP/kATQw
4QsNDWNYr2533gMOr7gHyXdSO07MowezyAto8Z5NDvzgMMB729quhoc/Q0s+/fGs
ZGKNsVcuUtnKW3PoTi8itx5K+XuPqP3esi7CBs7TRYIe3511An5i6zqXrYItOYHt
4apoIFDSXHrNELFQ6EmuUjmgb2F2xqkQRAHjxf8xm1Yt8KByNBXY1K51asIEIGuh
xnqkCJKAQoI2QVac4iAqgVHDUQCKTOYlC5EYxg/p37AD+ZPyqJPSDita5dQ4fNIb
bbmCP9aXNZOgv0uqJQ6VaX5Y3fguCGG/H7V9HHRpNyrtysf54VfQVIVa6/ovw1l6
rEdIgzCk+luGh3m0Xe/l5gpSChUHYDiZrC5QatVCMaWfTLoi7jmmEj7olM1306h0
XmZcf8ipAUpuCYg+xSGHXwIobnDDvdTTvWvNbPM6BWs6sePMljXSlAOkSVDF7u6e
K67wK6mjLverrZ+tDDIvoBLedXO9GPanl+JCWpC7zdGw2T+L4dLuMPnvh6q6Crvp
y6izTYdQIG+M9H3nA56BZBPg4TJKYaQn8BXnd4l7G+inzs+A6LNWLWl/QSv1kEhb
KB8jSFA+64o5ES3cp2tDfFWPIIMjXsS9TGtTIna2ezW38ELKx6RbqwNMShgEFieT
xnuWlhU/iH5LdY+rdM7VAGyr4O+LQXvTFtfetA7id+PapJEgXNglOtJeIokQ9eCQ
gaQSNNZyZx+Q21X3ZaCjzOug4fb5YCXBbK/bd6rNlYkh6SU+fVK59ZgKIHrf8AS1
Nw3ybrF4rmdXL4qE03GF3XAn44EkobM4WAp4E4u4wHVBDhiUlOPj8gG8NB4eumnX
2qW12EAyn5H34bJXK7HD/lMqMM9HbNODrNg0v2qLWTTgAM6x22AKFHV4+UJa6XVl
qVINhecHDPC8S9MKtqjxY7+jKHRiX4Xxx0GQKlxraCP3mbEfauiF0ggxiOC2UZZf
K7VFnfwGYQ1eQ8lnQYS9RAdbh8I+BE38Q208SZ7uxwkg4IvnoUry7hI9TpzvS6/x
mLO8sKaqkekaJnKYwf1MFBHeVkBR0ncQ7vVPBID0zZv4/RtOL4cmcrR86jcGtVsw
geRDq2uOFjWqp3GtRBjCSEbfYqHR4MK2CRjG1fiYg7xSBBvFcBfGciNShi8ebIF0
sWTjcWs4F5BQRjS6EQb0jJcyeWpNBFN69jwZIa3e6zcJtOyFnZX5X9Ic0o0+xL+1
zYK+YdByPDRwS/QVvBVnAB09MNfHLqNw1GcB2IIbtDgxw9fXm0bldc4BhOdtHMPL
w7kEVWV8dMaoF8v50y4NusNeSYCHkQCLfKjGxNJUTaINunwWCyoCq+hV7rshsnkQ
YPFh2tCyilstzYbJdoFSCbil71TCAIB3NkFSR2w4BxPsI4HEH3neKiPZPKZOufgh
n8y7D/ObCRC6AVJF4gnvjbN+os9XTyCIkY7BXIGITFKPFVvdna4ZVNi2yC97VmqQ
PbRJ/EIVbXDSYnftwcTgnKvz2hu4/OP7AI4KdbbKUdZ8Pi6ZSUDD51dK+H1k4QGR
JV2FwLM/nMQk10VkACCekBuSSDxGgdi1zqOK7mgf1e1X797K4PqzNwGXm2ITwoJe
QQbcxQAbMEgv/fWbOsVNzO8n7zf3B8Zb7h5MprzyefzVsr42vDK4LL4ypCVmyprR
17h2T5GhLOGBXWCqP7qlUiCNsuAqkgeMjH/2QBPLeJ6VsmOkWk1jvRy2SeVyjJo2
X9NeIvtXPp83Cr7yqSsiCQk9nD8Sxr8BIlV+P0mQjFjap0cIaEC4kiZ2ZF/h3kWN
wGXNzRZD2bGH9CNfMcb2oicz4V+vxFyM7HYYmgmBPTPtN5604Sk9fOdzVBM3HkNh
ShT5Zy/jDfv9Ni9kn7W3DSIMIXjfVOanXC24EzGQp+FLjTZ1xV02V700155gKMsQ
fr1hLBqPzHdniBL5ZG5RpZ5JnhARAs1ISchrUIlHkDxl/irC+qaeIay4zl3Q4WR5
o/w/VcrUYHNCtUWKnm3BDs6mSRsIs0kb9d0/Qk4neeOkIOY7IEI/zbSuYwmQk/Ui
62WlaycgQ8XwDCqcu8N64v8lq+8FDkI+/CrAJVMhkCXa5F45gXYsTyk+UFogrzg8
W3979mixOs3QD945nwdYWQ==
`pragma protect end_protected
