// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 01:23:58 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
miwofb+2qwruzz4+l+LL5tKP6lotx9ewsBfF9BkLDmeDRaLJGrxZcKJzpccF+iy4
wvD/vN5RtPC6VGmtppsoIZENj3Uuqq47+beVtpW4lQv0vR4hPXMQOI+ilLqWLVgh
yStdG6o1rl0CNgLvXLPMGI1epnO+qYHN2HfyXjDXy2w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31728)
QWW8awep4CEs7MXbQhM16+lEqJ8W+ipS9nzn521t32CjkC3wOGtLwVRpLCGgFlrf
JFbisNlSGBY67i/Fz/ibsBqEi7Ko6j/PXIlrCN9Xcl/N9CRwvg6N3MTizMrAviBd
hc14H4rlbdpwb77qKKM52ti/irvFhbAZSjnm7ghV8tCjYh/0UBwaNgwe3elx3gu5
E4Hntrn6ITdO3GnrCMrXZuZwNhZS9/ntkV4/dBfT64Uc/9cUPjBDdhOUc/Z2ENNn
tYYPd1MyikxtMHCJwSb5qoK4aAtX6nYqPfs2NVolcmpcMdf9rdhUAEmPmcqqdoVL
NKiXQ3BsA+3AeouQFgPvPScQJDvELk5Syu1Reg3Cu5SFBVqPhQRe+t0UtPPRD74z
QMVe1f72LooUninY+Pt9yDzpq7ZoNXPxUatb6x1t4nYcQryEbBzCGhWqzcV6afs1
yPVl6ZCqSelZzJRUHWqqgFwOmMPoXfUeGrwzRViGQaXTI84/TmsWDc2mkcRUDZlS
cJ9WcaJUvLjWMQbqTJFb0nbeS9eRQLGGbzP7+iENZAbOyzrbrJNF5U4AwjtQWcmB
WMRW3W5Jvp6Y0p+iVT1ZZ0sz2bLAWCAnitxmLzz1TBmt7sEXZAMYmbDZVNAfMDAE
p6YT/zS6ntjSbcEfj/u3XW3+o+QcYRh5Qa0SYJflsGKl9TFY4+lYUtm+b4pDpRTU
NZKgMQGvTyOElTP+PHGLgGVbUmU4LbEPbC1KsgWPmqD3K21ojHerH8riMcTsnzbU
rU8jXBIraj012dZeeA8N5vbiA9bNFQu1min4igKodamfaaMrHCI4jgp9E4947Ynw
BXjAYzRJ7T9sh36pQzutBGeXf50W+xgH4jmzHAsMDbs/B012rO/bCAy2FxmHSrfY
vl9gVFgHVzyLGtKrLWu9OpZMp36PntHSeI8O52AuLHl0mivX29Lb1jNKYg0EW8+o
8nIOs1KTZU9XXGGzbpT9OUzaxrGRCxObmZg1sG4VM5ZqHQhB6F7SgxEJILRRMrT/
RBsVASruWLzJDh8rTQXbFNXiNvZQDGlVJ3n/PUGDjM+Oyl+e+a2lmCNS8bfh6YfA
ZqlEjqkHv2dW7mkC6cRDGMXImnQmXhHP0ouwNpBlivolw1DjSzebzGG0vqb6WhaN
TJgWbutbTcQ6XVXK+gCh6wYxBxjjSAiXNk3c27xjz6oVIv0Eat4kqubNCfDyzfvk
Eik1svyinzn5rjfpTI7jXcAPH5XaGzHteWJZ8RN/d0+GsMWqyJjwop5kKu6xhAvD
cwnsmHkfui80dbCoAJp+wtIY1E7mHd+nWM2xSYrdJLEyIiu5IGq7Bdxm22H5TLNc
Ubo5ULvQrrbmlNwTBSYikWExY8cxwo4otJWvpJyMaZQekx3MYj0228ghVVj5RxJE
Xt5AMmkAJ/NzoGrBkChTouhLBt/RgW3dBfpTCuaHKTp2/SeBNSK/AJ9Intx1JKjd
P9wC/0LHFyApRHQAbBX1cdtrkWOE2IGKsonvSzw5AcvjAQconp+j4Cihpljahu0m
9y9cPqiwQTuyTqAT67tiYefRSl/m06D61JY5gvT006SK/hRUUpdiHEmCq33XB/pQ
fHbgFR3Xdu/Xiq/gQHO/sufMxQVc2QcrA4u3rNMiYUEM4SRLHv0zeGjjLW3oXIdE
vgy6ajoFh1RWnFylnV2F5t7lyuUEm7mvoQESfwgvMd5ziL8zQTRhvGxtOmAHt5eF
zhAIiDEv1iXSYmzby4XH7jjpAv0TyKeH08Zz5RbyxmyzsSHFgjM+uiqD7jkqglic
sT7iM2bPdojuhWCSYkUCbqup8ibO6tp/qt3tvZERE3b6ZB5v+vJMa/7hgyuQwuRB
UrgYF8GaC1zQ8XpexTb+umsIzC8OzPOAg8GU8fl8tyzkww6M8z0+JvfEpsOWDc7n
aJe+agqpvR5yYeNRe8NZXxP6tfS6txpKERqJzKwNt+fDJjPbI660fjrUpY0nePEX
+zr7I7YKzSyhEdejJDb8xMdRoBY8zvOv6fhJVHkoqqOy6to+jfkomtFGIHG8quu5
w16DEgO+uoHvSANyLnw2NkqAkkZxpx6dICTEyYnjNexsfFTc1k8fI+NScNnb93/R
bMG1eoNVEPqzvGhMZbdJiL0qN9TzE1mdPPct0DXtgY8cr1MAqux67ZBL2BfF4JDQ
l/fegpkE1BAUnEuznFRR3TisJsSUfMbKZowEZxB9/kxysxuptwxzH9BI/bmMRZza
x82DWIvmE9Nib5lGyq1tJc9dOkfIg1lNvnjW9BcBkRt+GKwOdOVNI3gzRXXyCEqu
JVFwDbiwYVTi54/mvILBc1F5bPQt4Nc4Mx/Nj8TvpAI401Rqw7PPJQZrZlUEtNFR
q7gaCuoCOgaFwc+l5gjaEX3mBYmAzJrEMvzWIe7AhLi4Raa8e919saEvmjo9yOfG
vNdNObdhFRA7hbMqiC7W0mPuDHixX0xUQkgd7SPc4eVQ3gxDZ+CzE+KBtewQhMSC
3s4acF7HAfN6hQBz7pahRXbbUFKBrGLoTemK+I+XeO8Tzv1wD7vUCwvUkjnYIa87
YtffDLZG15s/oikF6ycq3nn+DBfAtA63sDV4bQBBEzgsRlahzlInvWsCQd7oRIYN
i0xM4WoWocR6oaVC4U/xnoRSsqCX69NnkxrsxKQvtW8Us7NqvTrPUCZ7O47cDYyf
698ujb2+94wX/C+aPHxocHrQNMn9qe7wexRiEeJqnW+NsRLUHsbhihfmgFHzj6RV
OoGWSsDCt3IBVQZYfaw9ilIkgzP10gp2c6dFb6/yGeU+wWydFkeQlmNZSipfRCxz
ZoRhivvkekDVPreqReOvIRN+kxptL/sZFySjNjkyKtiobZNqNah7YE2F/7uvKQNu
3wRg7rVTRx1GR6DwsrNmkJg8q/7MCIEL9zr3pb1LDUE3JmUYSJ5wAFPb7AaPPm+t
Jan5k8Spk9lwHWILabMl2G2d5qjCSdMZoTaSVPVyB6T5KwxqsYCMCIYek5LyiEkt
VODVWELg7QsUlqG7CZurWCbUqP/l9KFLXl2egBIhGTL99mBfS6BrKqqGnfwevn6F
/1MEi/gcxLXFZvIpR10xxEi758QcOqsrFD4OX0pdblsv1a3jn0ZrYFh46Q9YXKDe
E5Hl7QqwzbalF0XQhzBg0/lBbpYNajWeLV2vzYjYVaR6vrlRsQbH5JCzCFTzqLWh
y1XRvbtRa+rIBYeHLfeFM4r9MpCAncb5bw6Soo0TPO1yQ4V+6JDxmlH47Y0aAiyC
qsR+mavOJBYxULO6WlboAy3m+jE/4nr2Y28WQPXH+dlamcUXGjMkpiJQFv404STv
DCb2wWGMVinIEnHiEcCrPiM+2ohWg3EixgBNt0ahQlQUQ/h7wvC3FELq2TzF56IM
Emf3ZuqNTkqVlV7SOIrr1PDn2BnjDa8omjVRHiSrIlxTV1SjMRi+7Y6Q/W2coov9
08d1JXQt4c4Njwyz70ABL6LLJ/4+nUy8QlcWXdB7ymiOqDU7wWkg6ZPEv18AOjZh
LZNsvwwn4va4Wv9/VHZaQvjCSiq/UDj4dWnubeebHvrWuFfTJjd5LsZWITomyBzl
lwmYjfkaiVS/ybPAV2oPqMwaYFhpMKm4hQiyc39qAap1+G1tFuMIKW2bDfC1I6VE
a+HkDpUF01GzlP7MitEB9DHZgAagslqHInUeoSIxucGy2iN50PL8ObfeYvlF26U4
FoOsizJ8TaUoToC1xTrkhlqdvEYhuF603MGuA+p2ZxmO0o04Ja99ttEJo6A8LZUM
jZ57oEZWI1vDUzxx/dZKctp2uiWA3TJ/sVShdLmJCwsTzyCErxMgWKosyZ8EpYah
ZDbFE0fg3HLjI5RN3sdJ437v6o//uDIg7Ev2kMjnqnoawVJ1A3wRmunrM/pI6I8H
In6aqbyUPKw2UuR0UpKXnv1wQyedWv4qptQFgnuzPCcQBH245Q2PDueC/zvBRaGj
0b8afVcE1+EDUW6yQGCtHy4MkDxzSWFKSHXr8CLWdf8OkNX9zXt7SpfFoFuYbNLC
Fs+AQxDjhwLUKHppz18AR6PTfPG+U+SQ9gZCbhZ8sTHFbsFCROhxUER7g1dfg3j+
8IdK4Mbg9O/qwOm9kJErXUF+Lv9N9lLsYthlayDbFmmSEktRGxBsCgCTP5JsyRRO
btEVRFDDodyYK0EBEsPAZ4RPQCdFH1ZYZn6ujC4wseqH+dq+K8ZpYyk8+wOE2ndq
m9m/HgyEMzp6mPDcknec/truwY7nMzaswHdEw6vuJkURfmlP7/SfymmY25VuqTEH
jCos8t8SYvuQs7+h9A+Mi5sOT7oEV/xsxcHPSUtQpvS7c4W+7FlKpPxYnYDHrSdh
aLccObiUoz89KD1VTJ7jDonwPNdayucDkDBuaybqdkFzKeBUlXGOYehJNWW4NTvd
tqL5EjTPSu2nYrLI1sJUU176bcOXd/P0VC5TOFw1kTfnaPQWZgE7uGaMfYwwjX/q
YB+AWGoQ5OY09CLddlH71Wbqbn7/wE1rlIZasMrOlA2YafmyDFzUSngJOufKh1bi
ODy5yRab0nBc2bmdDIj4aZedq7eFFsvsLHTvb7eC0J/zO1g0QJpV+axyuI2DCsef
eVX2nZLcyBFFyYCjojiYWZ19WVuwPDt5TZimqnhK3PXkO365X3HKYUIzgWqqSxl7
GpERNRHcm3W/61XD7HtBEgMfWqqxn/o8xvYWiGrNvv0lLaS+cuDXsM7jjHmC45kn
6coqejRFC/NULkHTbmd+qKuqal+tDV1wuONpcpBx/lOipJm8JSBIziVV9muS2A+k
VZSHYvHeNCQf/uSQLLsiZ+1vQlRIpr6w6+wl63W0Z49roEEE+m5mU3A/URz+Y1De
5pRF1KRsjSY4mh/zu7NnkUp2xTi5ei1CBl6eaTE+MFe2a4C7RYP2YFCX9/2tzlBv
6TwonbDCG3vSTzMhqstJVXzV+kxCNvmfZ8uWz/UOq1XUb55QbvR8wgDRtgyBeQef
GKb8RHpy8r24ciggc3iVtmx+SIkOSacGjxwE/mafNF2fiGfwvKH9NbQkQNCWyysZ
zipjx4uVS/oULwDhVCcX9Zszx2SFIhQyYhojAoSW61e7Sl1yF2Fm9j4qx0LLHHnM
2ku5d6JJ3y0qC/X5dzFII1sO23s/ry3U/MxL+p22JnfHtf6a2+XhrvUd7oG+2OzL
o0cHayREEV3T60cEvGjpPnNT5+WoIi/iL6z2Qu+u4rZhxgNniyrYGmQTIc0wL8ns
jH4y4rXVaqYIF/Bw/0QSj/v9xvBt/SaYHiNn0Esw7tWt2lbQwiOgFKr25DZD8LTx
FOJfk9t2wgwX9V9LwyBL5OGDNkeJmzWj3H1I9yKjLxNCtwiR8VpM0KsQi5Gg3rbC
Psf1LB8Jpd1ATbQTGLduHsQ7aqNwBOPwjIY1yRgWzg0mRW/0hlQ6hLHBs82rhb9j
0GZA61zQMzwE158eNkC00/S55utTrBm0n4FkoHZfwEgwomkgUuGolKgVjFADBqwC
YOxsZ5mBXAcm5tPzNoRzv0sPAZoLyJqLraM7GQeDm6dvbvSpE1K27TxFqTRpDrYj
wWwVZ33AKn5cBCL6iG9hcTUpPJ+eltkKCqe04FhLrafZQeBq9h4suE6g9Os+Y0JF
YzGky21xbSR/LnwVXDK+vgB5dDumyTLOuSqcOkEGmo/E9Ov0fiZxCqdqSDnwVBpx
7JRu0RYpzOiJGMWgX6cH23YAKMrpQdrwBELhkfnT2ArGhtTsil55cRe5tWYheiNe
e/bM0msZtx1BpPXqnyHDB/jDMpJxUR5FXeC11usxPm3DD/zZeNrg7olmBXourIwK
zi0KynRslQS0hOpMdL0rnY4UVLMFH+L8yKyPtEedAo1lXwt02OKtGGO5dVDNV2PM
KZ9jirMD8eoDj7EihM3t3wuq7oriHHcwZlQiRdTUnI2MBNcEj43wrCou/5dZJGZX
YtydyfT3FN1KlTIxXSTnX7zRLgrmh+YC+t6c08vuhUSjixgVIcyoiOZkfCxl5ET4
Nik7qcefDOHNeFDGx623bTNZwMBwP4J1E7awyvoTjnatcBvx2lYexWbsiYOEa4KM
HoNgfk/Fz4SHxdSwf/H/MWUOOUmQ01Pa2SYALbOaOXzm9NqGmc1iFpAEJ0FDEZzW
VtYNGKuDUC4cd1hQ3n0CcT5yW5veLkZebd6/0bk/HRHYIF5fQ8/DhQ2vjgbjIg3Q
2pEr0PRjRIPRe+NsTSkBIIxCKiOTqO7EydirnIAcIMg7QYHmvRFj+iP2J1CTJRYZ
5IC5zTxCvwK5LS+19DXQHCCp9DlAr2sv0qMC+1byaY+B3CZ3eHFxgTWyeb9ZQLdg
1SDuU4LQY1CwIv9nBELjQgQ8yNENaIiXl+ui/i8IG752UAy/eQkmWieovd8raj9F
3HsqlU+HAv0WLWU+fCSWivPcHlC9Iowf4vgd4BsCNu3EZBil1H2Rn1OuLFWcWIa6
XQD6rkAJ1rkhIM8lqB7/JKAKvJK+HaTw7yNHuTdzebAgunRyXFunEf7px/QO9s8d
JFYca3UZ773fQ0ufGm6KGXYoTUB37UG+e1Edo3rTAc3iscGE3hcbSrMsxYd2R85r
+7tG9hgSfeUzY/0YM1AGqMZZHj7IWTp3EwcconDjkQ3/YkpRTycgez8AMQBxk6nq
upvxQxKSny2sIb2jKYosPPi3A2op0tSuD6YIV2T8bFIQtsIzNTUHmRS36uNl1Kzm
WFD+srBSh4C3GsAFYFzPhO4egMm49zMvW5qMQcq1uSeKwLcDnQnRbsuFxPX6Mbk6
yj+84KmkbZCHJ108qpsIoQ1MGc6hssT88OMyoRbzvFEcZmC5a0Dhp6TK7kBCQroE
ZPW91qKlZ5MrEg9uzX2rtMqq+GWryY8z+fv6yHttaB23gv/RmK8YxpsUwo1i6gx8
ui38l3ryoAUPtXK1n5PC3TbAQbHRvwLddjbFwh6zBDaPb9QE1PNn9UgFnwuV0zTv
X1uhS97fFj5H/Lgp/eMAHLNgi4AaObYMR6L3ibp2PZdeQaHCUi2qRRvxujBNQl+9
x9Emop9T9fV70hmSBRKOy1sPirLLAOQoFTpxM92G0aR6KLfHARdsSK7zSazJ+B8S
+26QK73INfMXFRMD0g0WgJ1FumxlLDbUV982NuIFas3qGfLZegvrTgVQZWsqgJRG
55aeOvYnZ1oEuVVoD+qqqPZhjk6eEbP5XAzcSzkkaS8jx5sCB70ri0t0z6pyoeeO
qKpKFc+Q5YvfaxRcUrMSYzdFJm8DHEUl70MjwIsmg6R3ovuWRpot0Yn6yuEV+2RA
rBEKudj+0FR6j9ggSWAjlFRLdGCgo99uJCazb3eIigEixs72co/BOFHFteo2DZVk
jLUHU2JZTosztpWXCSdbymIzdDhq+k4tbvkQFEaki/BfZT7z+xWsKIZEtjRyKaFa
bJamUzoTiPGbbC004wHSeaYX/rTLYBKbH7VbPdc75drg7Tf+D2EEQOzIHLMAZDQU
DnQI2Tf45TAa6jQ/K+LxCQJsop8Stv/3Ow6dS/+SyBnL7vxYwLmtqG4PmQunu23s
YlHjpEqCujFoJD5v+Ry1eo+XODPASoTn/hnWpq4JQo1CVHllO0gsmRJhloZZ1mkW
Wk4OdnbV69Nr5Q636ntSEd/TAAI/Twc9JQXSbJ9OyQjJedVel/dKEHBqzLyCXtJg
hfV9xNXh9dkVF0+QpXLMuof2yH3cNgEAkGHvOJslGFy1dDHNaSMXhz5QSFrFXe0Y
IyNqclc5SwrYI7ZZLUQfogNw8Vd6zFc9YiMehnJ2WA67zEdukR/XHKMdqMvJfKgx
zjOa2nzkVCy4Hbni5z22xWwR0IWd0oC612hUoQ8r9EV0F0LG3s5hvrVtc3QhXUpB
rygAupmfAXQgSXNRIdeSr5OY6vmbVSUR8lfTzKs01g3gn3umqfLCEb0gxvnVQ9zL
JH+bulKP1xp/mG9zvaUvFSK6SJ+q4S8cAc9jyptUkTtT+ek9herJHEwjbbP1hxoS
EL6af5Ik0H/3XNLGCFk6bXLeQLp4ja7UDkdHjKeprQZ4yWV3+eRVBHc83bebEVOF
H53T5olBGcmj7bh5wAm7zKzVJendg0N4565I8HXn6k+wh0dDOlJMgNuD3EZcftxz
XxSjtkAc+OlpsKqJlA1HZA2IEk8UqQw4b03L3JkreQWE+YppBcwDmGveGXj565O0
+hCFHpY3x+wZVPVpQM6GrWf1BgIRY58c1Y3WdriV+nkAGuZZVXGWcM00Ck2MPn/s
DAQHsJO9DuKFxr5eOlq++I9gvVS2/OIy6DAXAMTvSvfABhQzckD12UlcitWEt/hi
18YQnSme/Z/DkGwif+eFZoij0h7V+doi+rXBEU7GhGKtGJj0ZQPuS/sqCeJWoyJW
vDbaA1pFh7Cd3bdi7H3SKpmUtp5ixoiaFZ8mlQQRPzeL52H1wT1ex7MRMcF87KSL
godwRuP+581px1zNIOXC4/aZpuvhfemmOntE/+s1Orl6expHV88Dh+wG3t4kg2Am
3X/zqZ6Ai/AAEdcmquvNaHuTw6T9nmmwNXx6uXO/0pLpEI3kisZsyW4wbTThmFhM
K4Gwa1cgJwQfzhLcb9mg5vN1vpIspM+TfTA4RCcR79ldLT6mX4L9dgaJbI9OF/uX
/Wy7mXoq4Z0BKsZNxW/UWfIFdAkkfkoRJ1Tfu96mHfjDiAha69nLECJxbpYkSCsh
CIjI2vOlWDyATdEhdT1Oqu0D/b+te6beERffPZTcoUOvwTVyw+aU+R/+k8HMpWXl
1w6nBQRUqqu1MH7Kfg0Y9COPN/RzYRHQL8cRHgJSzUgEX9coqySuiIIFTxoGxQLN
QdiCcTmMVCKp71RcZ/0tY5SN0idJmuZGepLHfTtdwlDO1Ax66MUXHuBNZbl6F5io
TdOwt8ZY+Pr9+0n9yg0g+CbqB8t42wNfgPMKTimYLWfPg+i6JI+1kfIF+kQp7b/F
+1j5Ta7LhJsAxwr/NBREMjtPKweBTAOTMDdMMGv2jshT9svOmh2UhaTE0nWmoFNj
hcN6yop5TW0+ASnb561baUqEsKs7TK7i245Hna2v66MiFwOT9YT4IUi0wCduuS+H
Ogl3RboqDI12mVT5oipspU0yu5/dNVkRJbAFgLbHChkgWDU1HSVCiY+lXYs6kjUh
vRnhGkCRUtvYJnbMyGYugHxbSieiJdaGUHepUtPmqkxMOvKxgWx9Ip0WEl6YMxJb
zA31D6O/YMMxS6r7zSWGajZ8LHrIavoYqLho2Y5hMm0fmVzNQHw1U4tPgvZ1gzvJ
anPh2jMKR0+tSx/VArFfb2IlxoIBebbvkGxEyGCT1+ihI8iyfK96eGdS16qVFs9e
1nH87PERwkHhgOh2TbCUxou/aTILEUxz7hFPkzaY0hKzwdwZZ0edBIaoaZK83AFX
EOyAkjiXdYm/uHpOybzbmvtRYV2dFQz+mUqk060d5Z2D0svj/B7G88P2njoiB6p6
4La3gCXy1xj954gm1snno3r3G6Fln79PjZL6ZUiPv6BKtvIuyyztr9BBgHFx+xs0
Pj1tR9fomDRucIPALrPw23slEE+B2UEjyVIXxSKT2/gi1/JoVWlJY/gcbJMFXSE/
RSdJrid99mjT9YaYvTpDjodarc2Scwu8vtUS0DV0oxA/lyrTGoQHIM7gJsVG2CcM
ExJKmI7QFMqD31Gv1gHLZ/VPp40uaxCapq3M4A9+7/J++exG0T3QksPDNXPSEyjk
EZ3Wgr0swvzK1KFcO1kjVmTkFVA8wRT75sDQcCPVtOEDsL0lyCRuVbFJGqFJ9xfK
Nc7KYocGm96NlPt3aEMncjGo8ZUzDa+MBKxRCwvHVcFj5rogLRg95Hk3QSaBWiJM
1shRtM032frLRP0v78vwh8n45IwasceHkTzyxKqkYzj04cd3DYpVg9XEdgvHAv8F
KxpjoGj5abj4jIDJxWQFmw8qTCK6Tnpx2YJzFzZAYvrsL9p6pO+ZTVbRh9sgvF5d
7pe1DM4OFEPzNCh9CgjgOhy1AQlF1sMtKwCK6ghBQT2i1a/6VwS3URnun4ceY81k
UioC5Ie/Et1O8ZCvteiPBS6y8HUlk879Y6mOHswtDuuHysyxdmYHOESNhixammfd
UGJCpljUjDTPOsUQwoCwA5NrLVJwF42f2ezkGSq9yYsCBbHJvvDCkcH+GxUK9t1M
1S6AfEsovq1LIrpRBmfin6KM2Y0KsdVEp8jA+v3aj8uNie5rFTGjsH0Zd7XTYx70
se6FoFzGpkzMsm/Hug2i3EuD/5p4F+M05YSJ7Z5OVw72jHh+tWdagv+oKSOY0DQP
cd4hNQHm3Dlv+rSB+At+SqJlckBXb/Ys/zEG445IHQigPpwLHzttRv7M5eIBNP2i
b6wb7PrrcXgVapYfmg0KOa49FtQgbWlRYYTIErJRwFWTml/m3Tu+HOR2QQpTx/Gj
TNDkRquehURG9XYZf0GFDcnz2MjGu6sktadRbaKcrUlu6U64pYd/Rt59LCSSoUEC
VecKGyqIECwBzI8uCxGHSOI2aPPBzObS3OkM5VXvrbyUA8zqPQZhJCcLjMixjqgO
Z9y0n9o/YxGGHhiFFMyLTMbkD1X5u+FTIJEWUieF6pp9B+9e+D7QuL4uuGzleBDU
HRY/Jvojd/bGo4fFFhUc+IYCoCU9a4ySwkUaiOLcUHpXhNry8ahU0aa6vtXTXlqg
B6ZIsSY+StoIlbYtZIn0cU2MdVci1Y6jY4QhE3pSNZXjSHyESExYecQUR9NkcRyD
AURlbYXVJEzymC5zhvdl+Rm61pNVqXwj6M7IM4M7qNsewLefGxIxltHXHjN5Mmvr
eZut+Xdwl+mb0G6JEr7kD56iwuMAJW0YEaDTC20LWLLesoOBUwL8E4T4cLrzRaV9
y/49ScKCne8yL757QY8XlMR4UV4vZ74Pt0WfwrSwUzg8S/CvDMjvFrdJOCkwqdLA
1RRox/xi+jAHBOxUAsz6MTHXKgK9WfjMH3fN1e/9vAm6RI0P+VS+Dy9TVatchRj6
ghos3/TWYekP79ioGDQhiolhffFwhQpBgxsIKDC2ny/npjJnHXqKXxZ5fT9s/iAN
6cty07YBleE6KsKaT5cILdjYjfD3U6OHxDrUqK15W1CxFGrsIVqgLKZ8J4goxt7j
f65rejMgp1GW5YyadyyJcl2er5CijoAJYX8eG1qb3QuV/tnEadv15IbdeFo+KFM1
OhTAtQVhVTDX5CE7Py80MZpD7eLHZmIeE0vbTqrU0fj/CEAC62d2XqIkIQ5DCugF
jXZuq9IlohqOReTxNksHputqN/qPuzrxItG9a7brXLL4wr3LShHeE5XhIEOYSJJB
gTmLDqwfFEuhBEvifGqUSGFS3/vj9hm7Uoqkc8H8CaQOyw/tbh1sSe4WtmLiq8s+
iY5ndEtypYhCWsAfH74FbfkV5r8Fl1Z0OxF9TWrQTX0v4TZLs1VPrP0Tci+qpPxK
FFkLUJu6P1G55GE7FiI3+7KsYoyBYxq/t1TrxVBEuGlmwl6VnMym9RZY0H2M5R6x
DBMAexIHntZFMWJeSIa1/+axcY2X8Zq0uXXS93qIZnIFPy8tdR5fQRy7117eSNEr
/A8VkQXSB391JSlQbpa3Cz090THPzWwFzhWVisyP7z1isxSuD+HGctLEXaxDxzRD
SdUrNI+nJbvB1C7D1+eCvMLC0qgGue8h2WEU+8uh2zBVdEBOpgkYhdjs25Z438az
z0Dkj5zmYL2CrQZ0wj9pZ9I2BfnqLXfUhl9hNA2LOKODFlkjYui78CVD6vvfS2Dq
PdIuVYzp4gLCDengd4wHSDYcXwfjqJPvQ1P6It3Ai73WBND0N6FXpwECnjJdlDdx
YqxhJAo699W4sSiofgj2u74j0xGH0WxizWpoKB+YCBzQ3jlTmd4VP310DYzj7czA
QZg8IxUNrcXhg+u+aWwMKortk7CSC3kS826sSOItwZ2Yb+qyZuwrwVqTXfmC7cpg
gV42YprzD+AsNd38qCUeAYf2MGebngLxaWabbiJ9sC+oA7sQDQHo6brJA9c10Lo7
D0Fxry1jexEzdHDUR80j2bDFDrvGTbU59z6j4qyEsptexnec6eWqkHaONOjA6AHI
arbrj6dGRAINx7PGecA2NEt/PFXua+WSRgjxQT3qgTVb1QnpHrZBRa4NEQCyzjWp
Sp+XYnMm2F0HstA+nKzmNdty2s0c8fYFK39EG1PY5CiGn7s3wViDKWZ8cWMbzW8u
X2oBaXu6+KpXM0B9smxm77nGIkrjpffGd1vRkBNCesK4vEwM8e9nhse0ZMXuJ4Y8
mVJ0jYZGnDWylYqJr6Zq9YoARU/LDr03LiToQwTZSyTiN78G+3DBC7Y8iEACV0/+
QzYl+8SVDss6qNJfTZJBky5DD9oFp1AZ8e1ZhLVdqGrC5AbO0t3/c1prV1kMRPvc
xaMBcTJqtuBWpDmDF29XSYxGG3jR1MHByjaWIC2R05ouD/2UQf4Ad5LA0OLxHKsc
xF8ga/sWz+o1Rz+CXAC4KiU3akpEan9uOToyME1viXHwz0P5L6RANDOWPj43Tsg5
XeVB3BHdm2nNszsur1EaMZ1yegjCyQcdyLlz1fWBffE00us3XuMKhRywofKxlLyj
t5qKRoSukBPxACpYb8GtlmVnGmar9Gvtko9TCs8GeyruhBZ3cSYk+7d5dgYC/VGL
x3s9TDq2hy63rppB1aYDMI6r83jQBdXJDspWhJKdC7LXi5iKK6jKUlQFU14m5nw4
maiJQlujiHT1H9+/CGaakm0Xyb+GLGGeTUyYMTqBhzd6f5VKwUWphgkjYwN3dspb
sNssEkSLxTvcK2Sjsu+x38qnqP08J7SH7w9BokLPvAtclpw9FR5T3AoQjD964SNW
pi7DJpeLWSZtQjNhCqlhpk3An/QXbtdGN3h9sIbJ790cNaksP4UU4iFiEGD3TyPI
3coWY3tEXZYi0bNCDaYcVzo+MTg1U0f6vatp43pt8kl37IiDPXAjzzMP/JhYpm/j
QqXj2eopzc1Blhh5j6o4+dNSNR9MAR8Vs/wJTgqRq2XcsCsJ5M/YeI+Me/mpjXk9
mjfZgnIAlX9YoYCTdXBQdqS7OMu51XooKzt2fJGoDwPHS9a+vQa3U4BbYNN1MwxY
W9Jrr0fyhY9yuXcsQxkim93p1pl/C3VF1pu5vWmar+YLi6o8eGvteScEx5td00Tg
pAvniWAaIuo+nRZXmZL/h2SG+gjHzQqMAN8Vf+ft0BMbTkDJ+X2u/0OQorhXZA/9
TnhayxUvh2wR7HzS52GKW28SV3TbtpXAsSTvfFfoRREVBYy6W3ttYbkcfDkuhwbw
2PmZFzYBVLFotoT/B5NY1l+n7YzdIWd+WpYvLWlZCnSYnZpwNqtUiKtnOyDVh5nZ
zWI+Y+m8qgG8/EuWoUlduyOGd2RfuVjwMxGsW+gUV9ruAyybRZJrizzcI20CLHLP
De4c354ECsW6m7VV5CYhaFf1Fl5y/hFOXsD6yaqbIz++rmrAfphK60ShcMcHQiw3
U68KKQd2yIuMUl+s4gpQ7Fpnhe/OiMnHkEzQu3IC7gYUNhchgRzGmqAO6N0TGLBJ
rRHCBn9+Wd5jxJUPf4o22yRPF6ESnYMeGn2H00un2KR38POSLURFbrHl1BqV3F0q
90e14ZHRLnXgpbKMjhRfP4soBbnsgHH6ILI0OTUHvN/OQn3i33Sscs/rZ3hoMY8d
BN91YaWPmPOwhA+H//48K5CObmLBAATy3wyEPqSjHp13m+ksyRHPGFeXz8QgDUhO
a3CCcT1xocUKRh/YhB+yP6GDVLlak8yVjjXg77cdnJz1YTHRJY4Yh0L4cJRkxhRx
1ugfRUAsPaImeM3dUqEWYDJhNrgKCAVL1m7Os7VIbjDGnM3Bp9NuR5aa/czkLjcO
c0U5yXXYS6ceJGJaCvtkaFAVE6baKfXRsZTu9YmuC5YFoUPGUSzMtxht6PVvHV1F
r469+gVHoYQm+bTmKFJhSPRy2ZzLFW76AuAXVlvz50KMh+kl/NU56W/tJ7QnuhVy
hACsoRNEo2y/cujo8QBdMlpdTwZP90ANKjxxibwCbqIFvFABZdMciEBUsAk9uV49
rrZiLuypb1WuKqPJC38J4MUUtyBFpsi3tOurC6LYSd5/2H1SJQ8M0cNXwcjI8FPs
KCIxiQOLK0wc10P5V1AtDDvtbddtX11G7VYhipBn4wbEZ1/4a/hT8XwMvUqT+I6M
xLZ+9XcF2ftD0zaBbsAIeOm5kIx11x/6gMmJdSgtpvRZY5Er+Y2f0TUgGFsBkFf3
8qmNRk0nGZOKTWK4Oh6TJgV+c810f2mzVAKbEflMDcflQkT39+8TxiYAH1nWKBdp
cvfy68Fv6r/BQl/DHGQ8EifeIWG+eJOeJHpYQs1fsTVyHvqI9yi96hpPQinlzvVm
NT/4HLqCaXLEDlgqn9RaJWhgyzusnlcKq7Sy7kc6UXHBAhS4Wio49/N5GHuB/kDA
j3rFAcRg3ElMLGVvJssXlWpoMr1KjgYDJUkMcA+pUzoPk1R/Vlbk7/mdTJgwYitS
JWrKtMc+GiGiSYyv3mIfneyGwMUITW2jvKt2YK7kwRUP3pPF/tKsQyJIVjKXEabS
0DilxBRuSA99bZLmLb2gBPSSJqnQToxoR0ZAIoaG4edZrFWgsGWSC7BJBGw1u5+k
cGGCV7KBWBXPe9U51mTsfVHP1yVMdPVmaRTY4PfQTthgrt+2tC5+05MItIHG3hZL
kAn34C2y15tzJ0g5EwmvkpVpQXzCuVoA3rEcdlpUgPj9/n7O1Y0JjWQbxDFMB/K2
1T3mbK5dxeT0rTPT08ZDj63LesNylRYuex2kS0FPZwufxhTp6VomhivAPEEoDhxR
BdasNaw4GScdjrr3sDE3uMO+xEUr+R17bRmKKpjOY224qsHOzzvG3Y/R7yHiHg7l
Ninnbsi4mk9xS32qOS3KExdqeq5k/ZBzXi7GR72rkz8HsMNnLuwk4Ywpx/UkXJDD
Vuj7GmzHoHhMEWtgDZYi25+YP27SV7ZujTG2Pus4sp9rmla+mL2f6LWZTdxE66A3
4B7V2BhnJgGGNC9aHHhLHu96axdB97QFhuliPY32PBy3QBD2yPHPfRyW2ZyDb2xh
CjC9g4ezDPt1dtU70FfbYCxHUeGuwOP6W0RbAMwAHOGVzVjw70WFTZa4Qkk2i/4z
8nGJDzyqIGEl8F3jFXrhoxG+zBwsNXVt7guRT+QljeHiSvqSzeDKtfZWWSrxp5bc
p4sQ+EKBl2i1QVJPy7o6Qux93QWFzoHnpl3NsCsR7LeGkkE0UPCVL5H7hDJImfOy
6EJEhv0U3FnTpLttVX4gJbOA2XwmrEcuXadEsEeE2PTYUBXruwLRtKmVPM6MA7qM
SF2JHO+tHKgsxYglc5wQPVq4NvgvnAPHEg4ZGD3HJxPQO10oSoErekPvWgy0L7pY
46AeAeRPHJCSCvEKFzqUraE4EAZD4DqPP41D0df/+yF9ybyYqimirHF11AmS1Lus
eyzci5hxzmy2mEdBc4PeosD/nXc6Pv7OhDwLbZJd1jdPa9lLP5mj0hlT4CcgCOMM
IMsgswhmgIjYwdqWiPHwQbxL8Wjo5KplYrWdhIoAu8W8Rpj7wWyc9DOjoVmbthoZ
/6Yn7kIkjrhjMQOJjTuHwgiXJM0NDXyTPA72UrBfHIljvvtOZ2KFOzmQJg3mHCWt
kSTiHNIy02tOLH2+wfd4MilZkPVpTmEr/M7/QCMisWWo54wkGrCJIF765ku8A+Hd
Adi9CQCzYOnjzKE1A45j6VyQP6dYJWJkV4W5s80zZnqg5mNpxVqesn+RvPzSbor4
2cXSV8wJ8VixoQti8zRO9SA2MMETTHbfiuKVA6vCr036hyJKAm8GVSngWHiZHb40
1Z72XLop6tkrE7k6MvwgUMvs3q33jMfjbs+kjkEQ6ibLWPh/+SLEtIQwF9409kt7
woIjN1jSKpMpivRZ2KkIJAiimrByPjh1GlceEP1B4+lf3LeIt0OLtD9zgrtoY5Md
WmTAPdUogr26mm1ntZ+g2rFsPZieI9Odb8f25r9ian7kkO+UVc7V/YVc6pmvA2GE
fftU3+LSGalUhN6kocgsFYvFcHFcnaxJSkSORPsv6MnBZitQ3w9TNF2t54rgF08v
t+HdeKuQDhULAkknRWybtRDvJwdkRZS/6iJMw2DIM2/5e1e5+rkvw4h4ogqRViLG
SDfLd9rK9JcD2nKRnAIwZvFfPd/OJ2A4jD/U1fLRMnHsVoSo5uLHLo5R3fdnbRDo
DVJNmEl3N0jnkTcp6Zn8lsYDmNY9aOIsdHk5ZnOiCeJKgslhc9rqsY6eNcEx5ymv
3n+bIsVBWdZHTBeA1rOZN9wikNBZqx+NgKQ3Ye2K7s1VF91wNz801jgYeDFNgvXz
boxQPgiK3RzHhqyXYjMzG7Tv4qMSbRQx5z7EOT72j0W6HwambZ4zG2F88dc+7ZyX
qNVpTJOzzHm6C5BwX1I1TvZ4z608Qlm7wbHesgaSU+C8wE9M4c4+2tRrKNH8cf4x
qzoeRD8CDGqZc1vLrfFVAz/wSIxp4FpYxRbflz90l9YLgpqqp9r0/mTkV2PpCspR
e51Oi78Wl2HX+vmS2xJz2lvNLGgdqZBCUu8WJtoQJWiq+db8r+prch6UXGeGRj5H
9acJXzSXu5/fYTrJP1hdyHoITGNQcciv0IgzvSJ3OY8YY5ZBZ6hfxDZjUDJ73M4C
KjJFvyKpsb/u+BzAIuAMRyUdaiQsNKIKvf7rle7rIVmgWgZbjsYSUTLsQmQtkGao
yhjjFoEzVFYEj4Z1d5yU5VCXr7yHlsLuWm9aEePPYXXho6amnissUksmbEckOKpL
yD7EtW78DUI5f5uiiFv/9k5Id31HDyZrordJxoDwoy0rNCziQZAyUgCQN28JwcDG
dGX46uWcab1nyLWlRFgA3sE6nRM4qczwJfnlBpDmWoDbNHmno4ql2wCOgUvFNqdm
XnKWvVFv5ZUqFSQzFUC93Fldxm/2DqZ7N8eS/aDA5b+1jAsN0DcIdtpQEYqYnbr7
+yogiXV7RbPnFk+WVu2yyzdsmYW3r4CXY3yAQLptkZjJqhvWpRW3kon527/XIfRn
vdl7vMOmhc5aNj+KkuZPijWkVojlL5fm3IMk7jVBkPQqjLYqOJN2BFIhXFjUL55Q
GLxOp7R70gQm6MQD2lZt8WjiibzNK35Cxt2CWh9sAeDTl6Eh13OUM5tkxy8THVI8
AVuD3Tddw5sgLVISDIsANIJoX6yJZoX43d9CgdBinKnUdLUIi2rok4izMdnl+/0+
7SjndxYRBjA04UHNd7Hva8wcZ4i83e1n+hkuDo0cJ7SgFEUTsR7ZDu2coI21Av8+
Kkzk/Gzst9ovIomfXgqbnuMJWAEycZE6zNMW7i786iAahOe6CHovw2yiRlMMWpgd
anksZK1NSACVvGLYDW8UXxuTz7s7lr9Mh2iCdN5+oI4s8dvP6i7j+9yvYj1+zyp7
SA+hWQYXPbP/T/7MMlAtnGtjnCbaT8rYH37XV6F3gpcxbwxR868JxvaVUs9nqo1K
dsWuCCgYJ+RM4mNbmx1tFrHyq/EwMmhlybamaw1bTcdX8rokk8lyatmgERNPZJga
2HXu0E8RsZ7SYNZjQBGMR5fqFd/o6wxdoG8dcvgqxIlh7uBNjF2kr49m/+YBwjXb
Ca6tWN/zkIcO0jN4s94Kkt9ze3UNcAMQgM0oaZa4mNOw/fNLAzXGWHHr1iKgR32c
GVEjlHoU57aJ2X8tHmMaPVkQUbyeF0V75soukDT2p00mMjeJlzLhCai8lbk8Tx+Z
jUwewV2Z0a7+VanVyND/K80+13MiSNL9Ukg868WXGkSitZoKOP6hg2IiyuJpOKuq
sFYCRKE3gcpN7dnoM5KAap7Xh5aXQsoICBBqLITvA7P1sFnzxVHHwBpEVcaMWAvh
gNFHYcwWlCHD/9UOqeT4P4veO7pXZ1X4MaM0zHvfYTTpj1va3GKZD6i6QbeQQKU8
X0J13Ify1Er1AFb9I+V+ylCzr/ibEUeozgAbtaVjxwd/D9n7D+7z2hg+9n/zEkwh
Xv9tj8W7LRwbdmPPUdEGOV0AbY3I/4iWtj5KKjAhv8w03t1SuBZUB5UL8BvZErjI
Uy2qKpyi6/j4SonyclnKb9xJNwZGFql5AEuEyvuUrAlP4SBJbuaQ6bm5MX9JnTPC
qEvxaZ34fbp6nCfdGAHqv6lqK424cCjPBpTKbIrTyN1AK92YLo20YoBN0sZAeUE/
m6WkBJa1is1I/YYuOdWfZUPi5l/hjk2srgtBkBVg0kfbWtNQqsKGeOcj7gfvqRux
jRFTv/WgPIUIcReKFKMbM7hji9NOhIiaif0sdPLhZO/HAqmeOjIZy0WpvWi+kj+f
BV4FSKWxwh7PlNN3wbVj5MhT8KLWKTCUu1Ps0QbRxwyAb2EDLsrOpbhcigbsEHkc
SY4ekGusfNf2EElTHY1tOVpio/y5GCLSgn5wExUfag+d/ynczupbfXi9R7eCIBGq
BKcqYWmpH1C0d5WoMbWSAEk5O9NvdCq927kaXZpMYDXRIZJrzmfpHLrX4aOWO2uN
zNYvpIijGRpHOaZS8uxrjSpjwwSjazjk2DC5bYj5UHMDj8PKfo9ucYSotxjgMLuP
r8iV4FFPHeIH59dpvpCvgGnGBHdTS2Yc5HJXdaK26uOk8oqmjv8BJ0Sb7jnicvh/
ttQmrFoCg2/zBGc84yj26I14eJjwAgguXatzD2o+Ct4JKxWxEXSPZ1Dq0RaZKBqk
L1yDdb0E66ryQSrOUSZxbvq3w751LiDb41VxS23SCGzCg7FaYAXvZNHx/sG4R4l5
TLutidECeVHEc2/56gzWqDHTbR/TqkgcgBQX8HMJggsjDS028XvWJljwUNO7BAki
6R3hH2ub85DN36Ts27kjdOiTK2skbwJfqRCelNaRpdndw5jdkBrayoXUxPsbUXj2
Qh3t7JlGQPh5q9iWN0G5UfL4oKHV2A2kOIUXwi/ptoTUMxVbbyGvMIuixeNg5yn0
qqto8cvJTJTbuthGubfwpmUvae18WWa6AedKhG9rxWdi69khmyKWQ9kNITuVTiRb
4f6i/ZEs1CgC/TqjpLcuJ+tKa9pBJF5e/wOhzBvbR9KLi1nVIM5xdlqn8Uz0Dor/
emRI+Tuw0cZduo/UPSN7+JQdQrn18sGtfy6WvwvctEB6oKb555Jr7If9d9Sz0mY6
WCSfpUsgmrPVXirt8JDjS4jDSTE1C1NvyhxJ0O+77neUixhtpkbTG/7hRZHgdfGB
WiLO+7/UncMuFT2NHBzvEK3hRKbEcSVuPP4rrvhlDeIpqDT7EcuNXDD855vRRLqL
DwTpftRR4WWdZ1dw6dX+3JqfKU2fMGcgObrAiD2C1pMVPu5D4q4rUS2t7n7FuDNm
m2WyE4LJnbsTGT6n3TP1CrUy6G11MR+oE0BAMM7yfqhjbHSnYydMKi03AkRBqtaZ
3+5wZGrHPzCRkv9ASdX8IYFA4pPpsMyfVd+k/0GKH0NA2drLg0B1Gi6X0zrbBTmk
zqQJA89/mGsIrnV/4wMSqP4KlLHg/C4LB1E6tt/rBgOKoGZArLgnp2oedml+x+m2
O3WlT6cDHX1c1t7MLhnYz5FRqDv/O+UMfmmJ73gbKlGf1F8CfNV8//bemmRcPXw3
HO8pG4RY3kWsh4R0oCrn8XkxTJTTc/YLkVk/jowGeJc7uD798Uqe9qyc9pxtRIHn
Tcqsl19OjFb8nV2e3xkOSnmm8XD7m48nm+zj1lklc6dOXOZQ90AQEcKkd1HGecIu
qyl3UqZSIppJKicDYZY3sPweuPCZeTaIw0aBDROcchQQ3YkKScqnK1nnQOGhgdiC
vNGgoKPQSiWo9qPlYyH5TU3zq0h07yPNSd8LyY+lQ+ykDo0xmK4p2/k9VreSxZTx
4YYD5sAD9KBQoHPx1Wyb0fmnCvt0hkFqbOWjYqw/a8UXXAIET34/1UDImB6ncwJP
AxEsXaq8cc+OaDfnaHqpkS3FYU3jLNZn8bZCakbGDX+mkMST0ceJYiDsm/726KnR
B+Dn/KbUDi06YbHFuK1TQ6MEmhkFasQEKpHXC6iVv8goobvq/6R+ocA1gzqEOb/Q
kmOmYyVpt2GQmCQj4XLhL9UPCvX51674PG1bx2/rn7MVbCuiZ6rbwneEbhXkt/jT
D5qNQS5G+aa523y9obTdSpK1MHOp1mf8+TeE0hcZJSutOKrOv1LIU7rAWfmWkL42
4I5/BAMFS+VS+6knJ/CWudC8mr9wqZQ/fC7lmubOTSyAZjRZMK25efnDtKgmLkRG
jE9nCei4VReF/NVJ4v7y63QYGUwunM51N9Bi46jbhXgHCKRzZfjvpgO9Y52PqMqb
0Fnr6Luzs+C6JzZ91OxWCBdZ8AfIloAzF6RpS89rNx4Kt1CjmGWBhUY/wp/bylCu
quDF/IwkuhSm+4PKFEG+wL8WFnmye6u4dOEtXh294kAzNjJwE/xi7cDKiYhmepdq
YNnW1ku/XPy00PUB3e0LMwjHx8Sj73/Aw6+TtN4qqC9vmISmLjveP7nCqcdB0VO2
ACGRk7up4ouKQoN07EZjc9OH9l/PlhHoqf4GZsm35Ac0iu6z93bH0ThBd398Zf3T
43SHhvVraxdJO+xQgOuvOO9M019Nwery/GECoc5xdiGl5FpbjFEfiUqodzjooDOQ
H1X0NX9vecAA7GCo6KnSOHQjh+h3K0ZuKdr/R1sG4ZXZTP9W4FnPTyV5vMhU4eU8
7J+i4CecPCSLH5MlxPBcLoZWJKs2X78YGTek9kHn53PxZGf0ygAT6cLAHmMrmKvI
rWmsEphIazP9fNIThnDlqDM5f1EP3k6cEIsweib4Vh+tPG2+E81JY2+Q/e6/DqT2
E62XXReFbc60MvXzzbC1d2s/Z5zxpGLmGXm6TOMa7Qz7YDnzIO0OxBsyt1qjFSvC
XwtUZjdzQJrMVzRUTQnqZvAFHXgC9kdd6ZpSw9GESqoyJube4P9JwoXVnij39mZp
RDYlYv8Pe6Y07lmB8mKIy87+OThgVyX7BfkcX86Dv0KWuIUdmca7NtjZxaHZMvUv
k9NS+B6/z7DBEXCwE2KPnXELS8wtQ3ZzpN6OdNSG1sOxNPepQfURn5FoTqEkgQlE
B8bXR22Py4A7EZudD4+IITFeus7XwIq578S1WIEXM/i7DA6+R5WGuI7/5TE0aYTg
XFhilZW4huHA83EW39EWAV3VWu6hIiuVe9/DNmoOnnYMvFbAwz6Fz+jkvqR3TllZ
wu8rVlfOBnP8Eq6WAOAhbyVmz27gLb/VV0htiuK5zlvhQXY09yBgQ9/MJKVYMz1S
s0YtjeMXl5ijG8oajpXrQJ7+qwPDjYhLMb/I/4YKKDFsjRe0b7/fHFtqwn/WJ0Uo
4yD45W05RXBh2DBKhugPPIndsME4CF9DdVkOHpJ2tf1tiHaNSfyqRpKPGxXA3AcY
uEIdeJAElMTV/M6lO4Va6j6d/2atvYslkx133TVHTF+mJK8H1ASj+5gH+1ioeha5
VG0LBdgCWexihiDca2Pbc3JS8wC/cNq7SXFFilXiVQnBB9pHP56fIyox4HkovL3X
5lK/R9flYrcwCzggfvW9VF8LXFgh6QU0ppYBfGrd+WRFyyohf/uk0xT7RDOWI52y
IpDHn7SXZCmVReA6t82PGTa9vA/nC6/x2wbWJnwDoBwMMNgvs0jdwGLYdxFyf4Fs
W4IWnvmpm1tRrgOqU2MfQCrMlWQw1Xj/juXy56kwXWJuAYmF91rod+dTTwvd/eRT
rQ4c2HFGqtCWVVWcyQK7kYxHQ/yaCL3suw2CzbUgY5VJ41xlk+o2XyQ5VVY/EqVw
+WFZA62rj6+RlLJQpxSLVv0zU/y0zQkc8kWu5pxDvPkus09Dz1IcKgKaKSatDBW7
qCkJs6pPV+DVNCpuWBT9bN18vf1w7Crki4w0MU+UJE88GzFcNwj9YWqloTrZgIkt
fxJFTenyiTO9Hu+mxghT5a99mwYkR4BtkYlfmZIpKtJ+fiWj9gyjSTJqSTCb6qB1
9vwzPW7AscKKZVn9BczMAg05DSkUCFR6kYUDLVGlxVQ2NzwrdLCCd4ai+mElJ+5o
99xuf0yEq6eN/di/ZU+2duM5xd/U3V1MulcV0dXXpUvzZ6ou2yfB6nG4k8sMScRp
Bpj5aSQgat4wlk+NGsQjNQNp9c/XLw6siyYjwCLyhAzpSYi2Du5P+ANHDAr7TIem
3DScr1A88Y83LgY+ZI5T2M3DjsFyekIBU+j+MMhoPxjaKKPJe4RRt4nk+NfJ/vFI
7Qvcu82H3u7bdQnDOkFlBiOppV839Z7jfy391iGvS4XlrZEcbzxzzPp+Kj9eGaD8
dbSJVIIpR+HC3eC/2kipgl4u5kB1ndAd0w7nXaABhINSacjG+O494ax/9q1fnVZN
xZZci5RI7VQw9p0dquLKGsxP2fZ7dwzE8Dq3GvIu/dFG9SnRlY9GEXfgm5fmDnJz
e29XAAB1ZaYBVsTAPmOi5KSrHtnZA6RSl0s8+1befRauATHGEFgCDojCpuTrJYs6
5vGmQ/wY0jPI1flrc6gZI8Vh2YYDHv6xqAY70qKekNVPjciaUJWn4+RTAHnvciVL
A0bbbt83bMFbatwPCNKavQn0j88S+Od2Xd2KXB9X1Ual3aspq4wAsKlMgI1QWoOq
D3W5NOZBs68Sqzpvlbw0xBfNygniKVfvUytxPHPZIFHbmtyni2SYTwM0BksLn+qO
Kp7UMbXPHX+j0PFyBY+Ro86geplZP0U0T/5VBj0YDY64iq1QWlWGiN62H9yRQDFn
F5iZTlSwQpUBeQ64EKccq4xcnVU5cD96mlRtI6M/50ZvRX8/27ZqsOvcUhea/ePE
lerWSfomCrDfTEpl0eGphOmHImvSaWYxS66j/TWCWgg9cDrSykpYeGqE4RLl8qtU
4UPUp+QDtMyAT7MW6Mjfp7qO9Z+ZOzcRXYnKUimd50kQWqLl6/EFUt+0nlJAymbp
YXayUMkkdNxF6w4nzW0fSkIKPcaMcZ9owCe9bXm7THD1iRRnXkRRmb4vS8aikKtK
EzRCgI02NuPwpXttrxI6o51lKwTtprb2rr8iomPjLgHlnbZ0D49llzXT+5D9g7lN
AOvHtUibvxjnji9BfUmVRourlI/XP2NK+fw3oFcAllrqLK0sZB0Y0Bgxf3WEJiDh
JjksGW72O+5qlV2t/3qovoig1ywYy3izqWYCWdloASnfGAjpS41NcNHP8Rb5eZJ3
xssV6rlCbeWc2EYOhote+NH+abFm9b+a38v+QsJTEfEaucyPOqE0tElagmJaQE6u
EEb1irPVLhxxD0Zr25tQqyhKLBQrOww1lGRS8jSO5/aYuNQ2oAccX2BJ9aIjSM5n
YNaTcnjoWMzwAYKrVmzN/ta1Id0lPTnKgAbrcfcrUkiDXjwit5ztiFdRxWJpCTYh
uqwZQh9CP8NTuNwrFgjsLhOfPVE7bPdd2TjKbW187eVh+vjEbyuAQGwhIEi6fFRz
WTxhrx1sZ/hAy8OYKXckOrfvAEmAjprM2B0u0NjXWTi177a7S/m/xaagQYmnF6uQ
d1BFIUFmcSm92q5idqRs78qyL0ceTzsq8cBCXQ4b6t2EOTXryFuriLtYWRz1UoNk
m/vg/KAV5Gl9ZODHlp0SmQQbmX3D9CdC7cyKA2CZcrXk+wT0W4f5S8uwLoev85L9
hT+tMwYUxTWMH05UrmlJXd2bhGqxzHwUTiZfE8h608wGNH52qnGAZMk0nl+EQqlA
93PZFh5ukmmKn7ChDU+y1dEmGe9rrDGWV6FiCXrlD7+7MqykGAcV4tRvahYFLIFP
ycwitzx43e3LoixZpl0uF6InQXpY+u5iiMTIfiMPZ6h/7qNDWHXmIXITjNLxDaIx
XVBODFUHBTvpmQQiyDCNwkkgH83jJE6hR4EHE4tDE5VbYaMtbTLrdw0SeWodRyd3
lPdhF776q2yR0lD9xkUIzYFQIkMs145/Q/D/bMVB7+cfoT3HCJ1+/IytovN5x+WF
Zp1zz6JMXKCShQI5wCBMQZMnlO/BHEJX6crmCRHpIV9fAozmwBo1ommNbFR7ZsoJ
pNQ+1glbeuJqwiqoBIPDFQbJIOR+J7daZNRiGmmRhXJNoxj/Gt3SHhPIaZO6yBlj
YZeMTZ9tcWsL4cv7fqKpwcpdpq6RqYmXR7Bw4mrAVA3Pe7H4l7BFIn0uO3QMsxM6
KRb9UpZHafV8jAKP5eXiBxXPEWp/VQHRWlBkyij6CRHyuX9Z3Zfy4leet4w1FhtG
LhAs0F1yrJMSh4oTdRLTYuRn6+CLPITUtmrYUDcd2pAeCB1ExNPq3q5fCPmRXITx
14fzlTHm1trlXWyVP0SNU7KLfQKAQeDQAk9QeBhCGhycQmXTnogigjSRhzdVyKgH
ojsD5OhoRrUUjOa/2RAxFG4KHa1bEYGPIffqSeC5CJ3cxurLJG9DtJ4gwSpXahFx
RRMpVwsP5j8C3mX3ul/ViWDkEntXgtt6lmkTS8MiEOUNC8j2Is0DU4kCcJzNt4xq
ndI92nL5lVN2fxbAZdnSphc0iQJEUIvncRNEI9KeLMvGpaHmdA9Prn0D9L+lIoiD
/GAS2P3/ElVAqJ0qXGb79kTA0XFhgsBrbEKknMrAo+0kh0uWS0yEZscXMNU7OQCe
2jD8rRuq+x45iqJMRPXVZ4pimv9NuHTiRl/ptPjMlyTXSbImlyhYODgEiEr2nh2q
f/Kqmoc9GYQ6rgDkVtoDOnWpYNKnUcfR2JVWugbKoRebIoyuIOe9btTd1wOQCNPy
AmOIguKkl97ir/hzVtz1pRVtHpZpB77Ng1nj5nec6jdMSNQy9f+0EPk7llzoJs/h
UDcRxapRwrZdb8emFwDVtMdLLSUZ57bej2Q8iPFNpmVKrv3VBU6G2cHfKrjbFl1S
nU2nWuONeq1+bz3mUv6GRz97nN7jV+gKIw3JNxTXtOgZAs9nsgXJrBLKzFZ/fID+
fOjGq0lHM3XuHly9LAfTSyT/Tz9sm9rEDsCPqF3XRG2bsrgFN04w935Vyflzl0Ve
o/mMa6FTb370UPV/JdKxFmSsQN30c7h6n9/2jS8EUk/eh+qSFnztYzQ0t9OJZ3mF
Nlakuq7RzJtgyJ1wOY93cZFJHR7neNzS09FlCHOMe9JHdJdNzYF++E94czlw9/wF
BpZJTIDzq5b+XbGSwUYS3+0+b23dZXNveBVZbSF9e8UIobnlAOEcorH2aE4NUN6q
+nDNse4hmx6wTO0h9EPJsJaGNC/IgL/s/pgM/UIG18DKDJY2+7CrgpvtQoVgClhQ
8CaPIAuA3XkKn3E9/PE+XkDWgGqYnwNPMpRsRbvzOeliZ8EOgslkaKYsBnrOd9wR
s5yaS6O9qyd0yDvKAcWfZ0EBYAeggF7iaR72fJCypoB2wbqnubupaY1hm3rO8VUr
orL2iWwqsuyIfFkHjbPgja/rF3UMsWlmTLM5Cu6wpmL0VXmSusn9xt8fgc7YMlth
fJz3/Hpp2You3Rw+klSbX+PwY2ZwqBktJhgfRT5XXTrkbQek5TKoZenPhx+yTBHt
hoFAZs0Im738/pHSwNnL5FZ523jCaNWtFhCiEnE4Y/+TRO1y06x0Frf5BEski3uI
5OrEwY4Ecx5SucrMc+wKTbucE5yOa6D1HARNxoWvWsIULPcV4t+sBpuOQg/pdN+a
YuaWcVyNn4llpa5k+Nobe4U+9CKpZoufH1FgF8fxlMZ8D95r1IdM9YAL6/XAdiix
EqEbsv1J9HviuqqNAmCZ1/hu+dNcriSoUu902Oe2utrgm5VNJWXTt96NugowH7ry
8dO0KQcFGqhv8iM8RU/KXib7lc1ivKPEZwN4oD+fKEXX3mFG1qrFImhM89ZI4ukA
lvW8ocxqS2jCcSkK5g5NhUR6IG33bOn+oq1hB2glvGbKkjVrVGwmUYocHW1semm1
X4dvnJXoUI5ib5z5Ar5K6T3Kc+xvKkj+fZAjf0tfKx3FYzRqpMF0JXJuHCXMh+J7
3vFC5QZ4gG+fdV8a6YiTaRL5lBnAFzVTh7ghqWXpbPxQmykUKQ4vlXN6tp3Ewm6J
A6suo5eKfdTgcCD1Fb/2Yd4x3WvYL86LQlPxPpOWnh978CCnVV7q8+Qfoo+1f6A9
aF62cCLJUL89Fv9mDmsNR2BRR4J0wXBk2VX3+jE5qAqVwoy/gBYJfWm6pgy7M4y1
11O2CKF1BBcKbDlJZBiHysAdR/vv9/W73Oe9AkIucN3GGDMWFSpoabl6rRAlnUnV
LNLqdrb7vOpxoc0qpPxzWEdZ01HTGDVbqTLRVRaXmz9XDaFyffts49kzQRt+/wg9
S4U8m2qJ3Tbn3mr48mdWCMqsI67qtB2O/rvoe5nfqZKBG48HTH3Jmctcu4/6XtC+
ULsTB2Xuy9bZ3ZsmAelJBmtQ3F2jx76bCV5LyfqCNpTj/zizoIRgKRelumpSWCrI
stN8OG1TRuTpBor5XTKXVPKF0IEqKBMDRAS3WfzmwSEeUeAaQamps64ss+BGoLR8
BCOVw1u+gVk7dfXR4D6RhIMwGTB2M55jmtrZ1epUN+EjAvlel4vXLQ2/B5eUleaB
J9sH+OrX/9ComOKPd9uU0BgHaLgcFTfKtAkwU+91D8mFKZw6lQjPMJ0YDv5opsTF
kxEq/oDEo19QVpq5ntX2MkER5ClABNaozv63V37X9OKini8/RCUfz5EoBNs74e/G
PuQ01lISTW7DXU6FzLNcJZrPtIE7uXYaHJoXOCelaxuQYTyMB4Ub5YlJN74xmZ33
3O68ZYyTcm3SlDWpM/l74FvX3N/ALAnsg3R2IwiEG4e5ZL4P74gmPSMqxsvrHbsT
JzI9QI+iiRKqdWgrAFYD+eExTMBGgHxaPVvFRyQrQwAEJKBhEDr4R/L6EPtMx6rx
hDCV+uLKYkJBcxkU7U9IKuKR9WbsNNWfaduzmf/MuhAwdtNgg1RXBu/gMWE06Das
v+eDLYloJR0ehqwDY6HE1BhHuxMNyRnaqCrqxuyBYq0mLSz8GFbl2Jh40x7WWk9S
URLU9Zo0VCXRN9hMLW7rjhFORB26i796clOlvY2umhYP4P1UpqIgKPimeBpEjYOx
BrVTWGfKGtEEsWhUD/N9wfcIRETHRke9GqscqFWve1bCVqIROvkSjgmx0FOBIijR
nmbZ+NyvVSqaw7hMwMUTtTQLRZf6Je9zauqjLxR1ZTsNgiAbIaqY8MCrheleGrls
iu/1ZG0MWbAtnQR8yhpHtrQR5Fgu4e/SLf4dyirgTIpAb1yfK6iGITmi7blULr9J
fDpbuLRvVVB/uoapgPaOJRX4d6jYfV7EttGy7wCrO403PFdudo5WE/R/3od4Hqye
lUXBDIhbhw3RBSTBhhcIKSbsZy5gAdUNY/gSnh05h/hLA5V4hFRKK+huDz/QhlpV
m5Ux3nzr/3snn2B6tTFitvnskQeEOpi887hc/wkd2njS/iAMp+9+dILy2Ut0AtCn
cQ7Vm2bUVDHTvjRdZvuZokTkTiGzKLlYbD1Y4XZgem+5MOlwxGBfFzHHM9d7ZwVw
q0B+LwD9l4TV7IZoqMCSKiwx5ZXJblUibb/1J+JcZJMdWeRetG12cD9+Mbe7sB9D
ML5ydJtteY9IKe+RqGUKe5q3TLhitagejzAHqVwOtTjpQ9UNz/A3dVM1c2iXPssi
rZG3bh3hfM61sweEooSTrp/Xe+pRw66M1XlAO7c7LtloCqHHmgHxYVJF5l4quE8R
Ym5OifoezVh4r4bilh0XpytPdL8XVZg9iUX8we4Hu+blDvbOZ1xqjcCQ74JK8TZd
jzboSXeJL3wDEZB1xj9U/eZzQA3niG8XZGqILz2hk84OrgUure8jWimHSbjr12Fq
63BYAwOJ4x2WcgxGVgrAltn0yPTETgY81VdVB7orVmN/5L0EgK2HEoHOPhJHOxT7
DSBWbHxdxtKafcTqWF20bgn2SR8NP31R/GslxgvFqyJesTKemaWDFYbyZOzCqRO0
MTqKz+lKCdaaclwahE8w16xPR6/0QamoUepRTS+wJpPebjX2AAQPBUd7/NbJohvt
l7CzGJMNsCHKxVpaqnfEmMfmND0MASrMyFgjAZav0ODYMRKvO7vnHsA6zAiDhBe2
XNnvQ9HMpHPcK4UsPJr62oM8y+Auyzz3Y4Kj+5pMzDkJTBQBvT0mgzNTJnz9IWo6
IzddjL7g/YPz9Dkw2I8laSqJZ12WOxr9eJGBOc2Wj4oaBpVn71hip2Qt7p1QAAj4
nSQTx5gYXzEuWlVSij41zApMkdmLAxnUKTTqL47LbDtJG68poSUDc+dwEeNP//wo
n0aq66Qre568rMnqtw0Vn666SKGTqhKHesxFr5vf1cdYpAZMaxcNhYEZgbWth/dF
aAxCWwPj4GGNHHeVor5xZgfDEsrPF8/mBDeqb/tUSgBaNGokbwzT9oYfWI7U6Jic
9js1q9+3zSqEe6MhFT/zYWVrst73loB5OZscvgJadvekM92qA5BSCW1FdYvpGFfQ
uKHwH+Z++bf6/CEjRoJpRMvjpzJ8FFLeBU2Kb9cd3OQnSIKP3ReUkOY+cm+aEg5a
3geoOB8qw72axAVFcKgK8/VLBU3E8AZkRhYiR7zos8gAhClRbK0gdAJ0OCZrnwa7
5o7N9ekKLjB03R9h1hEMQZKGhadwRS1w11qVjD3ts+IQsIyTC9D1j5JB8FGGXzuD
3R63BqZJYXLPOF+fPNV0TdEyI85mxYzIyJPEOLANkk40VNg9HxIWD8I6tEApk5nz
yOYkbq0WRumrOd58OMPZ8h8N+AWM61QgAC51mG4wcHEH97EXm6zq1RVrh/UoYw6M
LL/Dy4X6mQBKq+OS7hKMM+lap/TctZthhRPqQmsC9hBp+TuGXPTgd8CrIsx0VfEm
9+N9TVzDO9q4oQfcRhby9vjXjkhUhAsgHx55U5w3cApHvX3k6f3X3SqSJpXEsl7c
seuq4hWjODMODwgHHqTu9l3X8KxW+kGmtpenkhSAsfbYb/i7eHfctfV9bq28Bx7d
iKDezh0M1B8xHL1bcJIK3A7dn6BE0ZCUfPw7lZpQhTYXV64OQXVFVZPbIFZTKNRg
gcpXkrmpuYz/N0mLEEuEqWv5hbqwhNnkG2F0rKI3idFlqGyPTSGyzkiNGaSemdfT
3cWEbfcXTyRxx2ZTwUuk06ngug/RyDDC+7fdMZ6puktPuOUZpuwtvR1GmSLQTNt/
rRZlT/AiikSTRsjzjp//ciCAalbj+N+Gp50TT/ufkEuhpvgb/O1bBszLLhTvzrNv
lO9wJHG3Il9zH8P8c8nMuIwV3baRjWFtWzDjPfSA3OD2womcLe07TAHRo/Le2x+m
XwI3NV5BIAzThTG7StA2b6axvXYLTqizcxY7X4hRZhtBfWCIfP4LET4r2n9vm61n
sxV7AuLObN6/wxldYsgFHp9D837/1UFx21DtF42RY6KgCEMGAKFQVGw0CCEPmVrx
1IeyPRxfyySP7RHdAou2rmxd/gw2wDB3yiD8CjyUq2FY4OPL86cqHXplLfYZnPHn
1Wtn0OMWGAm1WGBayLKZwJ/aPNguMAtW6bD/E46wvTEABHR9qlvuuKMqkcHllnij
YLBGn6Fgx5Yvz7qPhkryWdfUjl5w/akET1BsoiIJFqSJS9OK9lcQ8srsrAcQYbGA
XlySMUaeLHSpFutgbS8vqIHYDMwbWCSXvuKOy2kH2RaE+gNwoHG8mvBgV6m9mzIx
ipq8L1VZ9zG59GDOFPafCN2qtjimA7UOnouNMnEVL2wAaBEDgLahqvBQ9jS7kw8X
rxQxr24r+NPrpVPSV1lCf/f4E3FpAHuUdz5uAuPKhDq8EXgWud6SvPC4TS3MeZf0
83PBu0YeYHXbQhZG0xR9Pb36rnH8lxof/+uxu4ofZ0cfjkYwuvsAgpDzfHwRZ73v
rDtwMGAoujyJO3DgNByh0/noer83MNWUpQzq+lISK2EeR9Ak8X4wTg4j7RyuDU6/
ZTKAuRc5eIrif4O3gCWlCsps9Zge60FrjdmOyWkuRCfwwdWOGIgmqFvmDogu00IU
4Ck44ojsIiTRc/zi0oASZhTAMZFMhWEYFq//ou1tylVt0I3Z6VM5HvSyExoIlHR3
hRZsdRV/jtQECT4/6wzva7reI9wI8t0rQTJAE+Sj+ghE/pSz9KolEV32RHwpY6iq
9k7NC95PoT0F2rtzLZ1OqHVaFqqfwJWHRXsSyfHje7/guQLpHcoGrsrYydAZbQtd
pywKsE3AsXyJp8trBVBXPiWrXyJBAoSP05NV2PQUf4Iic8+pbPxgT5V2Tfue8WNn
PBhvz0aL3bhdSzTzUXyvAnAbttKJTZd4jet4BgtDjf9lf4uV0KNdXmGk9Q93tkmE
zpxw2B0Ka9T1bejgF+jzgxlKYWTxO9yW1Cev99E2z1R+700BAhOHC3og3rRXdHhK
LflcI7GjWtToAe9U0SiEzVf7rNIsbViHYwdBReEoCL85gLa7jd2hZpXuXFFP2IVq
9o2mE/QwFNX7FbK2zC0cc9cymP/dlMIit7Oe9vQcoaai/aqO6DJwkxOFpnlSRctL
lBkw8x+Fd2cOHxPyRiBR1J5uxzqnzcckNeS56+xetivutA7JwrDvz0e41VTVtgfG
uz+2X1MMAc2WTObduVT0ZZVOYLbR0s38bqWTrqnKuLnIl/mx/S9BCxOo4wh3NnUZ
O6Nc9QyDAP4FRcrtgH+DGXuzgA5J6fZbMDQ6s0K/XqGGzcvA04w/WriNdqJ1/0Wx
xP6QtNJcpBvTvUzK4VotWRxyiW6lWjEhdqu+IJywXD5XOWKNsPjZ+o8QMgcNVOvv
pgwGozItpIBqGFVex9V+wrAhe8Hf1zUCzdkhIwrvCzGe2mk8Xu8GI2C+RM3DquQ+
EN4wyyjDURqiOwBJknYkX7LCvmz/pMw9J0AJlUywYsG+iucP1RxbeYNmGsartmU+
YJZ7RbvpRsVGvbHiFvjFzFkNwSNviafgDj38e6LjH+11ZIWFkGcFssWUJXLDXEKt
F2YqaP0jpLIKs5xNf10dZs5tVWk/5KURtnWpxloBDauNWOn2V/V+yzM66JKD5iEz
DDuuz/uT2MGrYxLi7HSKE51HvNAcwOikuO2AHke/LVkOfNglzAjgjfKTr7CV/dDR
EA5KRkhuwo0uIHvDuvQwfKgmZUB7fB7LhFyLlV5N4gUqJmqKdp9SG0DJYgnvqgA2
dRb3Qi73A8L1IU27bRB9bcWwgWa4yAy4OQxDf/wYOdRkxXfwxjeD1xkM8l7noXAd
dn8bX4mxsFncuuWWI1ZS8TNkuslhhuBMnuLJkynhyztRr7mCROdw0u7qPxux+yYD
wLvzLNGXz20BeDo3wYapPpAUxqGcbLhe4JBNlP3swjhNhhprUmTBvDrSm05t6D11
1FFN478PqMqZq9yPqk7B+40Uds1hgcyuktYho1WC8fXX9onNWxjqv5QwhYmyro1m
drjRdkEZ0lK6G1EmHJhFTu4RDOLd8Slbad0ulncQKedtlvMoIAgIWl3Ktu61qHZ7
KurKTp/+E4tuHDopfMrS7kj77jmws3TAlnpk79OvhMZ/ZF2qncrlplH93YZVk3mh
TZ+bTO2vjyaHH72Hmh4wQMeH2Gtl/Cdo/hocS0jfwWCHfk70PkOgWurv0okxX0cm
Y7JCaI1sT/hlNqr/qRWwYxgAWFqtrlF6l3ZfiaCzKbZWuWSKyXIuW05nAyKO23Tj
1YmenzgmMkXMU87F48TEzI2K4XxhijhQtdQB6vafmk7O2wvbCiFI2WZDNsoui894
qduqRS5UBRC2tqHtAImNtdqCazd7YQ25rDjou9N6ECsKbwr6fLGLGvYmQJ3kKrtZ
vPpGlh0nGxV8snqnj/f1ee5xfJn6JUwJ5LwYjl4Re9+s7+96jT54Zjt/DZqyzdA1
GQnZN/a14gNYcnEV3rLU4tU1w5WNEtwU1Y8qiEq+dhFtnYyfZg2ad+VzvQj2Z0Ab
VO2Eqn/bKHpJ/fXU9z0PfRzrqmWDGD0LCwown7+YS4xJsoXcHdCidfnyM5Yr3GGe
9ovBfzDMT2qcJtUEOkQsmIN74Wc1iOSI+jFiM6EdgRRj86wG9uCE2c1y0FzJOLHV
dgEU8L1mSccIzVGuhy+XC4/yC1e1D2PmvWR0BOCEDBMUsR3rVx7eIxfIngcIPcSw
3cKU/TnmM8s1RkkusM7ZE9f8498ofiah1412idYHNwcDa1WXYdEAMvNXJFGnUyYe
yhg7g+I6hMovzxTskLTTEsJSF7qBLAN/eDENwYELOgQA2pFjTPi0g+kCC3dAS40t
rXOmyJuMiSVx8UxzGWoJT/aLWGT8NRrhnLZ20BUUxxgxSlHVG1ZKyaeKKFrhs9Gm
TXMViPPiXG3/wyRbLkI5P7hWV3m4QXqZjbv2pEuqCX57/S4TVQkPFlCzgi5Ar3SY
XLg6asUISNjC2hk+HiUaaIc4qSLxD63aMlhqU5tSU3nWKQOetzp701jePSpQggeb
fNe7cuKegR2o203Q+zIf+MACrPtnFMc9wWvCInJrq8l0sVzn7w9l2NBVKGi8Ym97
uC0gcrbUeSSz6JBrwA5+GegO7ZOhjzDD68GW7ZKTMdykBuSk5sOjmh3umaNCHvEA
w7HEeH2baEu3ZGafGT+C656j7vmUSjDu+PQr6IBz9terdNR6UeLY7rEya7TJMc05
whmC7SaAO/fPcl159UfIck3kFtpTT/4wX8j2+YSFajJ9AU5L8DffuCKmX7BGFsHB
7SUfXOPQBfwhNBLSoZYCGCtJfv2Oe44qd20UWnFCpu6fi15MAYnT+mMNx6hUCVRk
ZPGOOFgnmlRABYXoMPj2jaWYaz7qpvCIxvWeTz69Y+3Q8K0OMNeJJCKmKZgjdaGd
EB4TN0dOFle1h+qdZwJjNgwu6XbZ1RFNDPEIxPAZ25b7bCZvzQSgfNtbkZ7eZOtQ
w4ZwYxOSKAWvN4lXjCfhZgNTGJK418YBiww+Y4XsjD3bTM3ZdzT/hTGNmgLdXhMv
O1TFKcMLD7rxoB+8U4NVjD2E8AVu6o6ZFF+rN6MQc7XmFtmS2ZgWWj0L9HR5e6D0
U7tbRoy5M881o9hK3DtnFpqruXDJqyAU9snO7l8wbaT1Gp1gaWPD5Whqd9kiDYFI
Cx0CyWNZQsW/vmKBSbf6RNf5YT/t4urqiq9aF2i9u7IYJTUz7GN2UspdGVHuZaNw
I7NzQodtKUIQiXHabHUZWOkz9yBjmIgOrXa33t6ngcq2WyJ6NBP0dwK8792qewpY
Dhi9ZtK/9Vad3KIEguDCGQppm8ORK2xxJNpM84+0QO1YD2Ib0CdCztxz1jf4n3x2
a+iohdz27iEHLxWwCUlPT32T/Rd8WaGaObKnz1h0vsahmPoUVkMEfgFRkS2FxGIg
WTBGOsk+TtUlYvVbP7Af3eqXlU/F3sAqD0VDAq04NXBX17+cNLeVWs9ub7NOzIJa
ydV4lWPieP53ehgFJJcwxBrTDI8o6BTxQj5mgYZEen3rIWBf4EDz1x3WtAhm4iHO
R1jS33CeJVVqRM/j96vPQuToXzrt0sLSWb3dxEl4qIW1/dA8RVdpttN8HLTxoB7g
VdCXWOzszvp//0TnXXdCc/nY4qfqmx47PwVgfRtGJ34TTKlvtGJD2Nn3TcGPm9v3
jIWQSRF6O1rWRL7LIFX9ikhmFOgKQpRW7wXdvePNgSaYdnSVk0xvHfKu83Vh9LiZ
V0VObefV4pf4+VxF7eBpj7TO/pPu+165anJYm3r8Wv3Yg6VOG4reqG4cMxLdlhHy
pSiI6WrSHlVfCFNgLO0JZmRrosBGGYkSwvaJTqpOtd5mQTZAOYsH1z/Lp/RFiW9s
kMvaGe5I2UqGxjDzg+8z+7GhlWFLtXzcrgqiz+PF159YlJ5swZ4QpuKp2Lh7UJZF
fJnGxptW5YOutP1Tiky5v4heoeG5+vKs0nsAhhi9xmfeUeUxs0rUzgtnwV7gTqfE
AE1HLuW15xzScYYDDoBkHQjhPyIyLdTNS3hNsjTCm4UBtn6aXuQ2MMDIekN00SSQ
sc1qSZW+szjaWMUeD1mH5FbdAJmcSV0g3fhw2CcV+bavlkjK1z3fQ1FRsYfQsEeq
f0dN5GnIlgpXujSPsP3nsQYzaAM1QbXLz6mrbhfTO5aCZsoN5lOmX22iiSvrGFsf
vIURMienbM+nhCSYunQDNOyK0eA7Z9RSxNht+o865zO5QZ35v236Ds2/nflBp5l9
fGnCPhMEx4rf4NMNWurGFBSZ49V7VM7JZ+SPfhbPwEd4SfvwfZarYuRWid53MafZ
DvaXrufOv5Y4mt2zrDmbp3+Fbw9lVRP270C+jYEKrEDv75dfSvZl1DAVCh8mniw/
wb7Ew/EgV7EN7LjRF4LZ1UJZh0aJOUjMJ/h/ldc3WMlvfd11Jyd5//GOrc1DkDkI
OyQ554/ZdLlz4ye8CEtGGrliTtRdl/uBdp4J/taILCQPYDU5IbJATKbJ43oSX56M
vudpCAfMgJ/pzBuHNrJLVemLnjJgImwFNsFHJXZkanViEUwSZBGLTIkUUQsl2lkY
GioRwJSMzceJkvHK2WOAeC/sx1PS7MiX4s06tc0MLjR0TY3ILS262Lp7OelJ2dkY
TRvqpFxRfs9zM1PGwuFmGFYn1xFI5cJe5YJwpYLeyEHMCzmdAl/UkGfjjznjSgRl
naMDnApQ19eNaVKQdlvXfSupzf1AbQxRVf6xqUkxr6oBS6IA/bR7BAUdMC/XkOOl
mcKJkTst0yQL/fUCqKA8OGZJ+GWSI2ziHy6jth7E+Q1iwg+iUg4SJx17kc5H68mp
EG5o870Idvnp348C7SQu/brHOv1OnQJ8gSFqNVf4xvxL3MNyFnTKJ+zLpE+ZaQr/
wapIXkUSz21EZCbT0AOOACHT+mz40J+LRRCZENdgk8PDIi2OytuUKzC0ZIxQKw36
lI6abGnJlw+hvVGwujU31BFe8rqHVg2lFoSjDU92NJT7IOn7wpay+Z4b2P84Qx4Z
HRSJnPFUd34LXvi/jVsfazd/+84oebSv6IR5OyPUxYGzE9t/xq9xV7UGwFv/kKBq
QcQa6dSdHYB4aV1H4pHg8o6qsVWo2gWRlcqRhdLa7RRBQKXR1+zSdrMJa4R4UU+A
7F/yQGDptduqvXiXfF24gXqgxZsO7R5gYCERbxz/9N9OWQ6b+eTOhsOJIrjC8J3t
DtA92G23ecS25lW5F+g4k5LKgdouILwKiBgSlQL8kkp+lEKxBKDplc2jQyEQkU77
gudn/68QIt4fiPAqnv1ruHOwtflwn78AdNQxaHWxec3WYD3wo1rECjpuEK+9Rstl
Pwgi/zQU4blKg2eYqAljOFTV4jpmmfmI1fNKIRyTrFv2JQVugyxzcCLO/KdJ95X6
vbFJOOSDpGKlKdStRp40kxA3lzk9p5OjrHk6gSIQX+x4OWxt4cESm5htUxgRHxUZ
3lWwRKB+fUHMIJhajo0M0XRSzrIaBOZlgBJrfEC+FnUt8qbPawwHI2GWMYwxoWxW
ee62cGSa+7NcZ/R5ObYp4YWsyvmThXovtWJ8fceTE7ZktjeqbbTRldWvZCaixkMw
R9i7my1gbGnF8xidEVox5SkVubSZWJHucnc2S9LoUlHCwxGEXt4RbeJfvh3iqyb1
O5uF35X1I+moHLGoqbyTXFuLSwCsVq5djMc8Mx7aRPN6LtwRHjLxtHd5ZtRlmO1q
j9DE+pVfK11uqVbABP239v+wGer/flkOODnIucIPPzrsyagt4OfFiV+oCRE/UsE4
QffB02lhwA8CF5LeCHVTz0ObyqBHP/z8InVB4ANqhm5aLiW9sWG8HHPttnkWUH4L
UYCOoOMeL/b4+Gh8AOz5ZKzhYFpmw3F+b7ceMB00uckZqQcok3fDHWvBzN2XVsum
01hIbzOPX8037JTrJaVRlfP2I7eRkBUREW5telOd74MzQV+V/Gr2991k7HnM5Ouw
+YO1LecFzzYygcQCXG0JMMqJE6Sw8gUaMzZdO33r8dHNShw3JFggJ6kG6wEeT75l
57HNz+zqOLYHYjC6Hz/VYyNeZbFnUMlA7DEN9mEpSbTaqhZNb0FwHDkklW97xagD
cgDy7hbHsyxCb2yR3j8O9UO0WH9ndOesbnkkPLOrxR7b2RDk+9HawPegFBvGUQzx
Rvk5ihUOYAp39bsmgirsERvoR8F3Ze66oH+WgFughfBxHnmE8CJXa1rbs57lEEoK
clyPYESjgFLd90BdBNDPEnNhwr4Bx9QHa+tT7Yzae3n4Ym7sZE8QyBhimCh/Z8pV
Bj700rVY7m9UkAeXStDyJ8jU30+F5rWzmZU46HhjiIdMQgd+bywkjHnkNRhjjWvl
MutlsUf5I23DL4nzGTe2OeHOhfuygYXRou3QuXZZT2KNRpbBSM44N8LIP2b9N2Er
8iV2W/9iNRNyb6TItWLrfxBQTEck3lEPW4YTrcr33JHA0tXxRiYrm6QtXzMwEEuL
Ios9S1VUnB453hFZDPwqUYwemjjzDUUGmWkxTwqMQQ9NMm77NMklpu0DTiBBE9/V
Jm3s8gWKBAIkJRGdZx0cwtOZGZ/stHc68VeGethjvrekUB3M8xMqcMPfmk2Vid6b
2QDP5Wq2Qh5Dxq8gU8pAVllJJKEA6EP1cpIDAo7u/HHanaIYiRNXMX4GcO9g/Ihl
A7ir0Xfo1YhFZrVOZiRpSPZTh1YrYu/vAkG4Itly/D4oAWG/lATWkB3+ut3p8PBv
ByZdCbvRHwpPSnMzG9MGI+ggi0Ghp7tDhMZj7GKLBz3/hDoe9NU+oy94/rGLsmwa
QxdRRg+2nUeTNq3Tp7+MUxVDMq4VXAdPjVdUY5UXMkon8M07yZUoHMXSSnG60Qpc
JOC4YtW22tdSgZ6nxiiBjStSB+uwdMv+I3I6MM/cVz+oi/rj5moNSTeXCdiKrNjJ
DPvbL33ERqXM1sNyt/VprFBuZo1T1t9iVNDp3GpZmqAF0XaqqINfya2KygZUTzvh
rS3dgPfSYh/u7nLRGTU9bfV18MutmddkWEhNweOHmnlNVtCoc2nHJs4b83lF0Gbv
xL83I9Licw99hvUsZ6v0EjGqe0dGkI5YnGJuGAO/sW3Brcu6mt3zXLTa8TSH2/Fp
rmtflIbSFLKjrX4vNJIw4KK/xszgy+DYttnfumtcNMVfd8BgjQaR7N2TFCXiy3A9
YUFQctyPP3nzT5LIv6lfObHTKlIAFoGkZCKUKzVS/0eeRHIuXiG8fe7y9qtj6NK0
QT14KNPAPwhjT3neN66DFz6acInJkGXx+KknSnRS6bqZZAJHxD0O3muuGX3GR3qq
WCD2M0gqvUgJghy6erV0xqwSt3yJCcd3pYqMm1278FvGWJLBqh41zW6szrtl82Uk
NdCGlU1Yqjl9jrXlgknjPfB6jnmxGrC2ZfaOk63L/3AnV2O2Sg5vPoIPCbi4xij9
qcOFJvmrKFKLgaSZaVT7XCESRR2on0wMIzZIXxDzBEn2oefLmw7DGolPbbe4zH3b
exxYJFI6QVPSLmsk1M4xzT1Ay5xTRG+KpIfDTScbbXPtHafngbeayBj+mSZHACn7
y3HC8YrnX3DCnj9+GsuvwhuAaudxIPTPnfSVN8kepxUOa0vaD/pVcjuqgtJLahNB
NSa3mgXN7nSJUIoRPulXfxSWcR//acWwrba/N8rGOqm8YNSUeum033Jo+4SOpiE7
jgiXyPoYbeCgCGgFoslvmBAgIV1Tv3dHB3gbG5Lg+Vzo8ORKxIU3TrNz/6jsSd8u
qhAE/rZfd5xb20H8ZzLQQv1gu9R92cXLK052/XAJEHo/pdtNp5+q5w7wNDW8QAWL
DGxabCycA9/8YfkMi5Z6qbu5ir5OHTaWlxv8YZaN6VfXGmEZtSZFeMleqc43+teS
7tRj+WO7unYE466RVryowiL4mFAOrQyckaXMh3FJLdUOTdPDq3mCkRpJO0+bdQT1
P7kCXxczQzhualDK5wEP+cAKe5e3atEYR392Re84Yay1DpehJdnUO3mtnmi74FZ6
JLamWvpuVx/NRxj4xOo6FQxU+iu1oNCwuE/9CAyFIOLCH57qDPeCznmXRRu1wvt4
rlxbK5roJo+9A59QbWb4T4oK881JRaSCFXM5bfIrfxw1GjgkX9aL740OJAs5Ma32
wdbL+hOxwC2VxJO9NjFxSgT2Z7717kZxeiyo/Go8cnOy5zyeSzhXtXJ55ZfCyzFq
IRLOcVW/4WlOYuXiKhuoYPu4VKWEgfDgVbCYkFhjAsivB+poCFMQ4oA/zbL2hF/n
OEHXcHcJydi4QcqedeKYy+NHLh5ThOg+pbRR9RwBIZnegdDtmzrHjEQhrO14OxRI
5MME8kMGV9pFQt65quc7vOmbsEsk/6E4k4QoDSE2+D3p9mbTvgGChSj9cbCvUtN9
M70KdUzyohICNOJVFOO3HNCMzxrD8y62LIQjfm+rQ1rUSP577vGYiWK0AnL2T0qT
ehff89RlaKYEg8lM7S20NZmF/2YtFtVe9UXT0cfnJjte+QM96ZJYDz7zg9U3IwYs
VIkrzCyv+G+EclvBJ0PRZTTo/Ni6MmOekw8Poav990JqE53XO9hfrpp1/sEgn0go
pDkbM17n4HhpqOx2kxQSvyJ2mIcCwETck0JCWpDflkg8wZipKs7s9JM9YHt/HRC4
qupAlsok612YisdeH2rExqAfmisWH1VEZkA/B411kDUGsVmOMVip9pxFF3/1HKqR
i6jsn0387VDz6hHQV+8vqLWv0Pf9rVlDjEJFTbzxmPusIDXIrF0yzSVM0vmmjrjQ
a823AvpuRfBds0YiFqpko1RCxr+ViFwaIXzznxa0/No/y/BO786dzOSwwLsVS4+t
p+nf97GFTjI+7jEby32wuFO0q+3v07TzKcDB22XzSiZxLwl1iVn505P4AbEybtSj
RD1bgFhB3AR+rHTydmyUfs0KjUR48NVTQXW36uCF3ePQF6b7u20CyfcRaJei1ce6
qWSiJd1qLVIrk0kU1q7oSrhMrnBX/WSeQInbcLC+0GDL3n6KkiAavB2eo+x4cp/v
Ye5Yn6bRNXtt6U8m/5vkd4iKEv9tJjM4i0TewRtYEC0EKJwnZq5eWt6AyLHYHmTd
lW09mESIBgVuvRg6iaZXZSyLm0Z+O0BntSiYrh60EVQRu9bvtwnx5T7vPkevuZ8Y
ueoQTKM+lvPWFFAntvIX4Qx8UMC+t4P+8DnIVB73X5mXPq0n46xvlMlIwI44uBlv
RqfALemk/8J3kaCRKXh2g9zLucfcGaXX7fi9dhE/CjGYCBOLcABG+iynN8QLBhc1
GJBT2ly4V1Emrt7wpXOcJejbxidQfemtlm0mvO4PX9Ijx/OhdkGSzJr/u5tywqYF
NiRZuf5fvt7Lng1lLYo/4Lr/rGO6fY0cFVsV4NDZqpfmakW5lJJOaCKLRwNOHo6M
0e3F2u31ArAS0YR73uj1qJ6e/eLW0FQm2KQihfRVbjqYJT+0z9pmqeAZjDq6MS3c
/8dbqXcBNvh7Ql507b/aMLXGJpRYUVr85Nts8Z8sk53BkZEeIYkFIT4/dyf545Pv
saTU9Py4TSYTrvMbzMhhTlH5IXdlQ0CmyiejViq1ZJnsLk8KYfeOJXoN2OmBHYne
s+Lgl2bQm8frqrelbU6NG0fbFsUeDEY3h5ET1tWSH/U0NPL1l0BsuH7Iky2sQZGD
NAfJr3FSoh5AQN5dC338jp7wCsdHybVoJcc2NdmtZjh/9xE1yNJwJhCB21DPLCyV
JwWCAdR8WDhL20wWaWrKDVpnSXHp7ypIbwehQeuR0EQdkQh//vNSC2PuZ+ngQ2GZ
7fg/DblftGFh/fKldT01VM04NJCJhMz1nu9j4UMgavLe8Nv8wglStuf1J0rB6hGo
Ax6k4GK3BL9rQ3kV68aIYRYOYNgkzIiwbJy2zpR1MDi1RcjDp8MbYKJFgpf+KJAP
p3CYFbZsY2ojy+p5puwbz8NWCz4HP+4STLkXAUeMDR+5ABAOJgK91i3WNbfHQtfx
3o5K4+Nl1597dyy6K7ARDBTaZ/YZPm46GXQlO40Pweama+1R8tFWM0fXyHoxVoHO
/QFMLQ8hAl27GBw2JyEzF5BJQUibopdkedfhd9U3zM6gM6F6IiSlrJXJFRtQlx/q
Q0C/huzOO/+O+3sbpbkF12gi+kbgMmgqIxZgdfN7rA/QihqsXG3GZdJ7U/8phTGZ
0cmHr5RfOYXTpqUAK1SR+BcfjZTlswdfcJZgKGJLnVzc8t50hXakSTMsXpnXPyBE
yl6OVSCYuN4Wq7J54uGHrfjL+tYFQzqsc/6fD0+kdVnj1O5pOFU1JfrnEzrmeUBX
wQ43wFpTt1HVi8uSUcqwauvZV5EpC3LXiIUJ/MCh/S0liSeGwV8nMlijNTWzMjWq
4tr46IW6NQkqhaXkYZUBZA3vfiTlpNB8xliqMQf2dzj1Uejdbi9YfUy5w58i7oNh
ZDNoqOWcK7aT4Rn8N7HdcAUwPWzzs7N4+h8pyy1PrIeXgcqDSDQTsa7uZr/GmUvA
fYEKZTfh3XvBpLcvMh4e5YHUHHeLeHohqKLxO/CZ25zL5VE38i4bEo9RSZVfTxC3
d4Ats3a9bHEnayap/XWBYOFDAfM+VaG+s9mFLeHnz5jFnQd+Dt/SVM90qb8Ia7Ke
hIGZprlITt9OulKc1gvqEA+ixy5ToIU0MEa9SYEN2frPs6SO9OUVw4N1W8hF3dNR
Xonl2055wrjymtrG3IYT2tG5/EhIfwYmvwho4zvIltq7GHpQMxycO+Sxtpk6cW7s
xAOdU/Jn2dNkySLdnixMuRmN8zH+MZXtvfsX/SuDyfXRQczFSAuyT1j3Mf9suTqq
urlu16chGCR29ZHrn9QNlWxfV/e/ciuca4BKWOOjJz1j6jiQ6NgEI/1dHvqRdnkg
q4sOrWIXLud8y10id+aHUeoqO+UJL6kp7/HlSyQYfPgHdYQhbaSOVEdN7f6bVs3v
ntClAqfk8WnWLKlpq7d90+jbApU0gQHk9/4vkwEMikYBIaQgGoi13FgoMD3awsxi
MnL3SWa9X0U3LVDEcJKomy9LLHtE8J4/imAb+A7LYpIAIZZM82FTx5OUXoLEcWqS
icNlNTwZZZr77oky4alz+eG1URAaS3qp8Wq9fYFGoOYpGrR+iPc1jlVU51ltnkuu
YkzSKF3JPbYASSrsG2ZeyyzYnbwvaaGsQmjc3FOyG05t4gp9n5Fp5bTsZdQydvYy
YnJ6iZv+RDo5IEBpXxvT1+T6xOqUlWKyHs7QxDX25hQf0qToTlH57Jo+dAuzng1p
IYrloXyQBIt9h+5Agny1hppvCsCtfgopPODDtA6cUy7Tax212fMtmyZPHIfA4lVC
tdeqrfR6DyF6X5c7NPxMHH28nOtuV0jLgdEe7lyftlq4CAqcnxVCL8ge4xLk+T8S
lsvZD18JZ/BXb8sa0ChaO8ViTm8hqBfWBTr+wT2Px7zy+6MieZU+PVbzy7gTOaYU
pTJHCkx8t/OBaDJpyJLCJiWrDuPRxNJ3UhHmrB/NotGhZGeIfej5Dc8zDYJUhXds
rEPve2W5mxqJ86NVtonunKUZGxOHniIKABm+6+k0sB8zK3DEiJRp5wMljJTqc5+6
8EbTbtpO1fcxEXCbs10Dl8aTVBDZsyJSO81KsBUN3m5n7dg4Q88hQ1Vr1T60vvkm
Qd68UgYLb3SLaWG8v2TKp/fqsKJDgRI2MMvtoTLksu7tL7DcLOeZ7ccVYIyWAT6h
QOprla6IB8puzBaPUQwL9tUd4FvCDVqg38AT+WmES8vwbcKnDJpuM0DcwYszvzpL
4d+AJQhbR63WvcDyurCT/SbTuq2q9emPUeTntMW3u0WKCR22gmSLTuftjVZXjDo5
lUFAqs1zp2CJ0o2XxXtr/dsfo0fjL/t6cshgqLD3u7MWt3eTbvSd96tC+ivkQEFj
uswH/3PkxWVjHTemnDOBd200cBhQkUHlKBzPe/sExPj+/LWA1BSHwRaj6rA+3L7+
XQE0MPWoBPRmGVetB5VH30r+bKMKzKBKGpudiRAIuI1tx1Npg9fY+u3jr8GtShII
I83SYizjRY/fwzDE84wG6qBLkeff9AiINMbtvwFbXIHUv0VE2mtVf5bgUIskz5Eu
bSodEeeUjGyhF0LT0qbr6j8eZ406gDlU/UAp9Ilg1aWIBS1HKPPeHXsLD0wGc7fT
KgoFpbAZSzorJqPS8/7/GG+Df5YDF5N+O3DO0c4QnuD6j9LglxzniO6ZHW77WIya
PNEpLJJKKZA7EIOaLHkX/Lv7X1k9hqrG9MZMCSe8vzAogMiYWP7Yd/fjXMZaOVCZ
sIbOQgxcp5a7Of5lIBepRQp3rfrKfexoEx5DAmQ+IlbLyn+XT/cw2GpzSYMW2wNx
`pragma protect end_protected
